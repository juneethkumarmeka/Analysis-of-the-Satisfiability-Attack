module basic_2000_20000_2500_50_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_1554,In_1687);
or U1 (N_1,In_356,In_1478);
and U2 (N_2,In_274,In_1358);
nor U3 (N_3,In_108,In_114);
xnor U4 (N_4,In_1893,In_1461);
nand U5 (N_5,In_1168,In_1569);
and U6 (N_6,In_257,In_307);
and U7 (N_7,In_528,In_566);
nand U8 (N_8,In_1021,In_553);
nor U9 (N_9,In_567,In_426);
nand U10 (N_10,In_315,In_1938);
nor U11 (N_11,In_1263,In_838);
and U12 (N_12,In_1115,In_190);
nor U13 (N_13,In_743,In_632);
and U14 (N_14,In_52,In_164);
xnor U15 (N_15,In_903,In_321);
xor U16 (N_16,In_800,In_950);
nand U17 (N_17,In_996,In_1627);
nand U18 (N_18,In_1108,In_1354);
or U19 (N_19,In_710,In_872);
xor U20 (N_20,In_1646,In_1255);
nor U21 (N_21,In_514,In_1010);
nand U22 (N_22,In_533,In_285);
and U23 (N_23,In_982,In_198);
and U24 (N_24,In_782,In_1279);
nor U25 (N_25,In_694,In_212);
nor U26 (N_26,In_647,In_608);
nand U27 (N_27,In_1248,In_1260);
nand U28 (N_28,In_1735,In_1838);
xnor U29 (N_29,In_1792,In_313);
nor U30 (N_30,In_861,In_1985);
nor U31 (N_31,In_1929,In_447);
or U32 (N_32,In_1340,In_99);
and U33 (N_33,In_1684,In_272);
nor U34 (N_34,In_1356,In_1729);
nor U35 (N_35,In_1455,In_1890);
or U36 (N_36,In_518,In_381);
nand U37 (N_37,In_573,In_833);
and U38 (N_38,In_1922,In_48);
and U39 (N_39,In_1805,In_880);
nand U40 (N_40,In_111,In_168);
nor U41 (N_41,In_1427,In_920);
and U42 (N_42,In_468,In_843);
nor U43 (N_43,In_1976,In_765);
and U44 (N_44,In_1854,In_1239);
or U45 (N_45,In_721,In_1749);
nor U46 (N_46,In_777,In_1326);
nand U47 (N_47,In_1378,In_715);
nor U48 (N_48,In_101,In_396);
and U49 (N_49,In_1299,In_697);
or U50 (N_50,In_1671,In_438);
nor U51 (N_51,In_1547,In_1416);
xnor U52 (N_52,In_373,In_1570);
and U53 (N_53,In_1691,In_532);
nand U54 (N_54,In_417,In_1874);
nand U55 (N_55,In_1001,In_1568);
nor U56 (N_56,In_1351,In_132);
nand U57 (N_57,In_1578,In_901);
nand U58 (N_58,In_46,In_1617);
xnor U59 (N_59,In_702,In_1635);
or U60 (N_60,In_864,In_744);
nor U61 (N_61,In_1429,In_1705);
nor U62 (N_62,In_1144,In_354);
nand U63 (N_63,In_1487,In_1138);
nand U64 (N_64,In_338,In_1209);
nand U65 (N_65,In_590,In_1191);
xor U66 (N_66,In_870,In_1662);
and U67 (N_67,In_1033,In_137);
nand U68 (N_68,In_668,In_625);
nand U69 (N_69,In_1014,In_1589);
and U70 (N_70,In_488,In_975);
or U71 (N_71,In_1469,In_1619);
and U72 (N_72,In_1472,In_399);
or U73 (N_73,In_379,In_1969);
nor U74 (N_74,In_1392,In_1974);
nand U75 (N_75,In_592,In_495);
and U76 (N_76,In_1973,In_95);
nand U77 (N_77,In_287,In_1787);
or U78 (N_78,In_1479,In_1608);
nor U79 (N_79,In_747,In_1188);
nand U80 (N_80,In_205,In_1561);
and U81 (N_81,In_1374,In_1310);
and U82 (N_82,In_1398,In_1539);
and U83 (N_83,In_1225,In_972);
xor U84 (N_84,In_839,In_1748);
xnor U85 (N_85,In_1869,In_1423);
and U86 (N_86,In_502,In_204);
and U87 (N_87,In_857,In_915);
nor U88 (N_88,In_14,In_442);
nor U89 (N_89,In_1099,In_1625);
xnor U90 (N_90,In_772,In_1774);
or U91 (N_91,In_1201,In_1070);
xnor U92 (N_92,In_678,In_623);
nor U93 (N_93,In_1585,In_570);
or U94 (N_94,In_1163,In_371);
or U95 (N_95,In_1576,In_1402);
and U96 (N_96,In_1029,In_49);
nand U97 (N_97,In_21,In_1492);
nor U98 (N_98,In_1196,In_734);
nand U99 (N_99,In_475,In_1294);
xor U100 (N_100,In_703,In_25);
nor U101 (N_101,In_971,In_1549);
nor U102 (N_102,In_12,In_806);
nor U103 (N_103,In_1140,In_1275);
nor U104 (N_104,In_728,In_1361);
nor U105 (N_105,In_1603,In_4);
nand U106 (N_106,In_1680,In_862);
and U107 (N_107,In_1265,In_949);
and U108 (N_108,In_1642,In_117);
or U109 (N_109,In_1877,In_560);
nand U110 (N_110,In_1773,In_1437);
and U111 (N_111,In_1983,In_1330);
nand U112 (N_112,In_700,In_228);
or U113 (N_113,In_785,In_1777);
nor U114 (N_114,In_1271,In_891);
or U115 (N_115,In_946,In_346);
nor U116 (N_116,In_1522,In_635);
and U117 (N_117,In_1040,In_1887);
nor U118 (N_118,In_300,In_1176);
or U119 (N_119,In_989,In_1604);
and U120 (N_120,In_759,In_1540);
nand U121 (N_121,In_1053,In_195);
xnor U122 (N_122,In_677,In_355);
xnor U123 (N_123,In_430,In_751);
or U124 (N_124,In_644,In_58);
nand U125 (N_125,In_1329,In_486);
nor U126 (N_126,In_1000,In_1675);
xor U127 (N_127,In_1210,In_1649);
or U128 (N_128,In_555,In_1319);
nor U129 (N_129,In_1482,In_752);
and U130 (N_130,In_1698,In_701);
and U131 (N_131,In_10,In_1420);
or U132 (N_132,In_1781,In_75);
or U133 (N_133,In_674,In_1285);
and U134 (N_134,In_182,In_1932);
nand U135 (N_135,In_221,In_1657);
xnor U136 (N_136,In_1019,In_1784);
xor U137 (N_137,In_510,In_303);
nand U138 (N_138,In_1071,In_1344);
or U139 (N_139,In_963,In_366);
or U140 (N_140,In_795,In_961);
xor U141 (N_141,In_1371,In_735);
nor U142 (N_142,In_1804,In_568);
or U143 (N_143,In_587,In_1848);
nor U144 (N_144,In_1020,In_1520);
or U145 (N_145,In_1400,In_1776);
or U146 (N_146,In_557,In_1302);
nor U147 (N_147,In_1615,In_150);
nand U148 (N_148,In_144,In_1668);
or U149 (N_149,In_1170,In_1640);
nand U150 (N_150,In_1677,In_217);
nand U151 (N_151,In_325,In_882);
and U152 (N_152,In_478,In_585);
or U153 (N_153,In_1481,In_848);
nor U154 (N_154,In_141,In_40);
nor U155 (N_155,In_1579,In_266);
nor U156 (N_156,In_987,In_1582);
xnor U157 (N_157,In_403,In_384);
or U158 (N_158,In_565,In_1602);
and U159 (N_159,In_1709,In_1676);
nor U160 (N_160,In_1456,In_1104);
nor U161 (N_161,In_1318,In_541);
and U162 (N_162,In_1950,In_1814);
nand U163 (N_163,In_847,In_1583);
or U164 (N_164,In_1352,In_1833);
and U165 (N_165,In_1409,In_337);
xnor U166 (N_166,In_350,In_974);
and U167 (N_167,In_1222,In_1881);
xnor U168 (N_168,In_1686,In_829);
nand U169 (N_169,In_208,In_246);
and U170 (N_170,In_1008,In_1536);
xnor U171 (N_171,In_1900,In_1553);
nor U172 (N_172,In_1391,In_1079);
and U173 (N_173,In_1613,In_1886);
nand U174 (N_174,In_93,In_793);
or U175 (N_175,In_1118,In_1699);
nor U176 (N_176,In_70,In_1550);
or U177 (N_177,In_265,In_72);
nor U178 (N_178,In_521,In_1591);
nand U179 (N_179,In_653,In_762);
nor U180 (N_180,In_1821,In_27);
or U181 (N_181,In_1965,In_411);
xor U182 (N_182,In_875,In_1244);
xor U183 (N_183,In_136,In_226);
xnor U184 (N_184,In_380,In_1797);
and U185 (N_185,In_911,In_1518);
nand U186 (N_186,In_1439,In_1287);
nor U187 (N_187,In_298,In_296);
nor U188 (N_188,In_840,In_1017);
and U189 (N_189,In_1090,In_1931);
or U190 (N_190,In_131,In_695);
nor U191 (N_191,In_167,In_1467);
nand U192 (N_192,In_1884,In_1178);
or U193 (N_193,In_1058,In_509);
xor U194 (N_194,In_273,In_925);
xnor U195 (N_195,In_741,In_714);
and U196 (N_196,In_807,In_1703);
xor U197 (N_197,In_979,In_1379);
xnor U198 (N_198,In_1066,In_600);
xor U199 (N_199,In_1562,In_317);
nor U200 (N_200,In_176,In_1989);
or U201 (N_201,In_1039,In_1510);
or U202 (N_202,In_1241,In_178);
and U203 (N_203,In_873,In_1411);
nor U204 (N_204,In_1112,In_261);
nand U205 (N_205,In_1525,In_1829);
nand U206 (N_206,In_980,In_1663);
nand U207 (N_207,In_1158,In_937);
nand U208 (N_208,In_581,In_1317);
xnor U209 (N_209,In_1270,In_1164);
and U210 (N_210,In_918,In_830);
nand U211 (N_211,In_96,In_1544);
nor U212 (N_212,In_160,In_1055);
nand U213 (N_213,In_1445,In_1304);
or U214 (N_214,In_1665,In_547);
or U215 (N_215,In_1632,In_630);
or U216 (N_216,In_962,In_225);
nand U217 (N_217,In_1390,In_1876);
or U218 (N_218,In_88,In_1867);
xnor U219 (N_219,In_1968,In_1085);
nand U220 (N_220,In_44,In_1949);
nand U221 (N_221,In_73,In_923);
or U222 (N_222,In_955,In_351);
xor U223 (N_223,In_1606,In_1366);
or U224 (N_224,In_110,In_43);
or U225 (N_225,In_152,In_275);
nor U226 (N_226,In_836,In_1529);
or U227 (N_227,In_219,In_473);
nand U228 (N_228,In_153,In_1643);
xor U229 (N_229,In_98,In_1137);
or U230 (N_230,In_1502,In_1045);
and U231 (N_231,In_1855,In_1289);
and U232 (N_232,In_260,In_1558);
or U233 (N_233,In_493,In_1462);
or U234 (N_234,In_1631,In_480);
or U235 (N_235,In_1656,In_402);
nand U236 (N_236,In_1659,In_867);
xor U237 (N_237,In_250,In_649);
nor U238 (N_238,In_174,In_1531);
nand U239 (N_239,In_679,In_1009);
nor U240 (N_240,In_1772,In_1359);
and U241 (N_241,In_766,In_1484);
nand U242 (N_242,In_930,In_732);
and U243 (N_243,In_392,In_866);
or U244 (N_244,In_973,In_462);
nor U245 (N_245,In_1908,In_542);
nor U246 (N_246,In_383,In_1281);
nor U247 (N_247,In_33,In_1921);
xnor U248 (N_248,In_1919,In_1394);
nor U249 (N_249,In_1645,In_1024);
nand U250 (N_250,In_1828,In_673);
or U251 (N_251,In_484,In_1979);
and U252 (N_252,In_1007,In_756);
nand U253 (N_253,In_1430,In_1513);
or U254 (N_254,In_1405,In_1080);
and U255 (N_255,In_531,In_1820);
nor U256 (N_256,In_1722,In_1069);
nand U257 (N_257,In_1088,In_742);
or U258 (N_258,In_846,In_1224);
nor U259 (N_259,In_15,In_753);
nand U260 (N_260,In_804,In_1274);
nor U261 (N_261,In_415,In_1764);
xnor U262 (N_262,In_1283,In_1574);
xor U263 (N_263,In_605,In_767);
nand U264 (N_264,In_1493,In_1559);
xor U265 (N_265,In_459,In_574);
xnor U266 (N_266,In_707,In_1727);
and U267 (N_267,In_1817,In_1597);
nand U268 (N_268,In_22,In_604);
or U269 (N_269,In_1413,In_1217);
nand U270 (N_270,In_1743,In_23);
nor U271 (N_271,In_1381,In_1234);
nor U272 (N_272,In_1667,In_1903);
xnor U273 (N_273,In_85,In_310);
and U274 (N_274,In_1496,In_1059);
xnor U275 (N_275,In_779,In_722);
nand U276 (N_276,In_691,In_1717);
nor U277 (N_277,In_497,In_591);
nand U278 (N_278,In_1514,In_259);
nor U279 (N_279,In_1862,In_1966);
nand U280 (N_280,In_811,In_1997);
nand U281 (N_281,In_237,In_1785);
xnor U282 (N_282,In_413,In_726);
xnor U283 (N_283,In_609,In_1808);
xor U284 (N_284,In_1957,In_1844);
xor U285 (N_285,In_1956,In_1744);
nor U286 (N_286,In_667,In_449);
or U287 (N_287,In_1180,In_1681);
xnor U288 (N_288,In_1946,In_1802);
and U289 (N_289,In_327,In_1690);
or U290 (N_290,In_1702,In_1162);
and U291 (N_291,In_516,In_1031);
xor U292 (N_292,In_1845,In_504);
nand U293 (N_293,In_892,In_349);
nor U294 (N_294,In_935,In_1673);
nor U295 (N_295,In_550,In_1600);
or U296 (N_296,In_684,In_172);
or U297 (N_297,In_1527,In_1948);
and U298 (N_298,In_1713,In_554);
xor U299 (N_299,In_269,In_1827);
xnor U300 (N_300,In_62,In_1043);
nand U301 (N_301,In_494,In_1197);
nand U302 (N_302,In_316,In_29);
xor U303 (N_303,In_1630,In_1511);
or U304 (N_304,In_8,In_1535);
xnor U305 (N_305,In_942,In_1192);
or U306 (N_306,In_1012,In_1288);
nand U307 (N_307,In_666,In_1920);
nor U308 (N_308,In_1565,In_951);
and U309 (N_309,In_1262,In_1725);
nor U310 (N_310,In_1172,In_232);
nand U311 (N_311,In_1276,In_717);
nand U312 (N_312,In_1878,In_1512);
nor U313 (N_313,In_428,In_1801);
or U314 (N_314,In_1422,In_1078);
and U315 (N_315,In_311,In_850);
or U316 (N_316,In_1202,In_1047);
nor U317 (N_317,In_1293,In_572);
nor U318 (N_318,In_420,In_1952);
and U319 (N_319,In_1474,In_1146);
nor U320 (N_320,In_1923,In_1745);
and U321 (N_321,In_227,In_333);
nand U322 (N_322,In_1334,In_1128);
nor U323 (N_323,In_1339,In_1593);
nor U324 (N_324,In_832,In_189);
nand U325 (N_325,In_501,In_1056);
xor U326 (N_326,In_998,In_68);
and U327 (N_327,In_1091,In_844);
and U328 (N_328,In_64,In_387);
and U329 (N_329,In_1834,In_1910);
and U330 (N_330,In_1425,In_1605);
or U331 (N_331,In_357,In_469);
xnor U332 (N_332,In_790,In_1770);
nand U333 (N_333,In_1860,In_258);
or U334 (N_334,In_1182,In_124);
or U335 (N_335,In_485,In_299);
nand U336 (N_336,In_1022,In_1978);
and U337 (N_337,In_1832,In_393);
or U338 (N_338,In_1912,In_601);
nand U339 (N_339,In_279,In_1081);
and U340 (N_340,In_764,In_1489);
nand U341 (N_341,In_578,In_34);
nor U342 (N_342,In_1428,In_1726);
and U343 (N_343,In_890,In_1972);
or U344 (N_344,In_561,In_871);
or U345 (N_345,In_1837,In_1100);
nand U346 (N_346,In_390,In_1719);
and U347 (N_347,In_145,In_1015);
or U348 (N_348,In_1587,In_778);
xnor U349 (N_349,In_738,In_1035);
nand U350 (N_350,In_1737,In_928);
xor U351 (N_351,In_636,In_1842);
nand U352 (N_352,In_1338,In_1084);
and U353 (N_353,In_1799,In_1733);
and U354 (N_354,In_1951,In_1933);
nand U355 (N_355,In_499,In_948);
nand U356 (N_356,In_1121,In_1195);
nand U357 (N_357,In_1120,In_546);
nand U358 (N_358,In_19,In_1365);
or U359 (N_359,In_283,In_1312);
nor U360 (N_360,In_1064,In_1937);
nand U361 (N_361,In_837,In_588);
xor U362 (N_362,In_616,In_1873);
nor U363 (N_363,In_1453,In_1184);
xor U364 (N_364,In_1557,In_1044);
and U365 (N_365,In_1607,In_1232);
and U366 (N_366,In_1152,In_902);
xor U367 (N_367,In_662,In_745);
nand U368 (N_368,In_466,In_686);
nand U369 (N_369,In_1150,In_359);
and U370 (N_370,In_30,In_1618);
xor U371 (N_371,In_1486,In_37);
nor U372 (N_372,In_638,In_483);
and U373 (N_373,In_1147,In_943);
nand U374 (N_374,In_812,In_1200);
nand U375 (N_375,In_1193,In_711);
and U376 (N_376,In_1796,In_16);
nand U377 (N_377,In_1438,In_1507);
nand U378 (N_378,In_1982,In_1145);
or U379 (N_379,In_640,In_1269);
nor U380 (N_380,In_1780,In_612);
nor U381 (N_381,In_977,In_1746);
and U382 (N_382,In_410,In_1468);
xor U383 (N_383,In_125,In_187);
or U384 (N_384,In_1082,In_1227);
nor U385 (N_385,In_78,In_11);
nand U386 (N_386,In_826,In_263);
nand U387 (N_387,In_1305,In_1870);
nor U388 (N_388,In_1650,In_1506);
nand U389 (N_389,In_1614,In_739);
xor U390 (N_390,In_1454,In_1678);
or U391 (N_391,In_687,In_1417);
xor U392 (N_392,In_520,In_924);
nor U393 (N_393,In_817,In_126);
and U394 (N_394,In_1450,In_815);
nand U395 (N_395,In_1537,In_472);
or U396 (N_396,In_723,In_234);
or U397 (N_397,In_539,In_645);
or U398 (N_398,In_1116,In_63);
nand U399 (N_399,In_1523,In_1728);
xnor U400 (N_400,N_47,N_279);
and U401 (N_401,In_1028,N_319);
or U402 (N_402,N_291,In_1755);
nor U403 (N_403,In_435,In_1303);
and U404 (N_404,N_374,N_304);
and U405 (N_405,N_144,In_845);
nand U406 (N_406,In_1707,In_119);
or U407 (N_407,In_1353,In_1219);
nand U408 (N_408,In_1648,N_6);
and U409 (N_409,In_519,N_256);
nor U410 (N_410,In_1223,N_162);
xnor U411 (N_411,In_1516,N_186);
xnor U412 (N_412,In_1363,In_641);
xnor U413 (N_413,In_1521,N_122);
nor U414 (N_414,In_976,N_150);
nand U415 (N_415,In_1712,In_582);
nor U416 (N_416,N_77,In_404);
xor U417 (N_417,In_1812,In_123);
xnor U418 (N_418,In_1331,In_1990);
or U419 (N_419,In_1495,N_180);
and U420 (N_420,In_821,N_311);
and U421 (N_421,In_620,In_1715);
and U422 (N_422,In_1588,In_1532);
nor U423 (N_423,In_1110,In_450);
nand U424 (N_424,In_1231,N_141);
nor U425 (N_425,N_174,In_954);
xnor U426 (N_426,In_985,In_1465);
nor U427 (N_427,N_393,In_945);
nor U428 (N_428,In_1917,In_1988);
and U429 (N_429,N_127,In_1154);
nor U430 (N_430,N_259,N_132);
nand U431 (N_431,In_1769,In_1883);
and U432 (N_432,N_23,In_1068);
xnor U433 (N_433,N_75,In_869);
nor U434 (N_434,In_1199,In_1695);
or U435 (N_435,In_243,In_1315);
or U436 (N_436,In_166,In_1639);
and U437 (N_437,In_1823,N_352);
or U438 (N_438,N_206,N_202);
nand U439 (N_439,N_155,In_244);
nor U440 (N_440,In_319,In_397);
xor U441 (N_441,In_991,In_184);
or U442 (N_442,In_665,In_1925);
xnor U443 (N_443,In_1524,In_584);
or U444 (N_444,In_1272,In_1815);
or U445 (N_445,In_1596,In_798);
xor U446 (N_446,N_195,In_1364);
nor U447 (N_447,In_229,In_128);
xor U448 (N_448,In_1375,In_1296);
nor U449 (N_449,In_1062,N_329);
xnor U450 (N_450,N_307,N_335);
xnor U451 (N_451,In_1789,In_1980);
and U452 (N_452,In_841,N_238);
or U453 (N_453,In_2,N_147);
nand U454 (N_454,In_1237,In_792);
nor U455 (N_455,N_146,N_230);
xnor U456 (N_456,In_939,N_312);
nand U457 (N_457,In_1939,In_322);
nor U458 (N_458,In_787,In_60);
xnor U459 (N_459,In_140,N_268);
or U460 (N_460,N_135,In_146);
nand U461 (N_461,In_398,In_1954);
nor U462 (N_462,In_1380,In_893);
nor U463 (N_463,In_1449,In_1308);
or U464 (N_464,In_1782,In_1864);
and U465 (N_465,In_400,N_191);
nand U466 (N_466,In_1633,In_1824);
or U467 (N_467,In_633,N_118);
nor U468 (N_468,In_831,In_297);
nor U469 (N_469,In_436,In_1267);
xnor U470 (N_470,In_121,In_1894);
and U471 (N_471,In_1016,N_343);
and U472 (N_472,In_209,In_1113);
nor U473 (N_473,N_168,In_1994);
xnor U474 (N_474,In_1940,In_577);
and U475 (N_475,In_352,In_1975);
nand U476 (N_476,In_235,N_249);
nand U477 (N_477,In_718,In_708);
and U478 (N_478,N_139,N_30);
nand U479 (N_479,In_454,In_161);
xor U480 (N_480,In_981,In_552);
and U481 (N_481,N_362,In_642);
nand U482 (N_482,In_1098,In_1386);
nor U483 (N_483,In_1840,In_763);
or U484 (N_484,N_353,N_3);
xnor U485 (N_485,In_341,In_1682);
and U486 (N_486,In_1205,In_1601);
and U487 (N_487,In_1284,In_589);
nor U488 (N_488,In_1984,N_267);
nor U489 (N_489,N_112,In_1914);
nand U490 (N_490,In_158,In_330);
and U491 (N_491,In_1290,In_1830);
nand U492 (N_492,N_61,N_15);
or U493 (N_493,In_1041,In_112);
and U494 (N_494,N_348,In_1609);
and U495 (N_495,In_1882,In_879);
nand U496 (N_496,In_610,N_270);
and U497 (N_497,N_328,In_143);
nor U498 (N_498,In_1011,In_558);
nor U499 (N_499,In_1739,In_881);
xnor U500 (N_500,In_545,In_1337);
nand U501 (N_501,In_1996,In_522);
nand U502 (N_502,N_308,In_758);
and U503 (N_503,N_282,In_432);
or U504 (N_504,In_1042,N_232);
xor U505 (N_505,In_71,In_1075);
nand U506 (N_506,In_1629,N_384);
or U507 (N_507,In_1119,In_1594);
nor U508 (N_508,In_1018,In_912);
nand U509 (N_509,N_0,In_1768);
nand U510 (N_510,In_1448,N_73);
nor U511 (N_511,In_188,In_332);
or U512 (N_512,In_788,N_197);
and U513 (N_513,N_79,N_25);
nand U514 (N_514,In_211,In_768);
nor U515 (N_515,In_1383,In_1157);
or U516 (N_516,In_17,N_379);
nor U517 (N_517,In_1620,In_419);
xor U518 (N_518,In_1775,N_169);
or U519 (N_519,N_383,In_530);
or U520 (N_520,In_1133,N_367);
nor U521 (N_521,In_853,In_1266);
nand U522 (N_522,In_1106,In_1546);
and U523 (N_523,In_293,N_4);
nand U524 (N_524,In_1941,In_223);
and U525 (N_525,In_1509,In_1185);
xnor U526 (N_526,In_1758,In_1385);
and U527 (N_527,In_575,In_548);
and U528 (N_528,N_98,In_906);
or U529 (N_529,In_35,In_1621);
xor U530 (N_530,In_353,N_131);
nor U531 (N_531,In_1177,In_905);
or U532 (N_532,In_1373,N_87);
xor U533 (N_533,In_233,In_54);
nor U534 (N_534,N_51,In_482);
nand U535 (N_535,In_828,N_178);
and U536 (N_536,In_1321,N_171);
nor U537 (N_537,N_136,N_331);
xor U538 (N_538,In_611,N_266);
nor U539 (N_539,In_312,In_1307);
nor U540 (N_540,In_823,N_318);
nor U541 (N_541,N_354,In_544);
xnor U542 (N_542,N_323,In_1166);
or U543 (N_543,In_1572,In_536);
nand U544 (N_544,In_1498,N_363);
nor U545 (N_545,In_1350,In_1250);
nor U546 (N_546,In_1658,In_796);
nand U547 (N_547,In_1335,In_67);
nand U548 (N_548,In_1443,N_176);
nand U549 (N_549,In_425,N_294);
nor U550 (N_550,In_1174,In_369);
or U551 (N_551,N_58,In_1251);
and U552 (N_552,In_1025,In_614);
nor U553 (N_553,N_161,N_83);
xnor U554 (N_554,In_720,In_65);
and U555 (N_555,In_199,In_1533);
xor U556 (N_556,N_37,In_241);
or U557 (N_557,In_1060,In_251);
and U558 (N_558,In_709,In_1491);
and U559 (N_559,N_332,In_1779);
xnor U560 (N_560,In_1661,N_26);
nor U561 (N_561,In_1567,In_1756);
and U562 (N_562,In_1208,In_1738);
nor U563 (N_563,In_422,N_156);
nand U564 (N_564,In_1257,In_1101);
and U565 (N_565,N_188,In_952);
and U566 (N_566,In_268,In_94);
or U567 (N_567,In_267,In_414);
and U568 (N_568,In_142,In_676);
nand U569 (N_569,In_389,In_1751);
or U570 (N_570,In_409,In_130);
or U571 (N_571,In_458,N_365);
nor U572 (N_572,In_277,In_1306);
nor U573 (N_573,In_909,In_1388);
xor U574 (N_574,In_171,N_167);
nand U575 (N_575,In_1918,In_978);
xor U576 (N_576,In_24,In_607);
and U577 (N_577,In_511,In_1072);
and U578 (N_578,In_1880,In_1418);
or U579 (N_579,N_89,In_820);
nand U580 (N_580,In_693,In_1664);
and U581 (N_581,In_162,N_85);
and U582 (N_582,N_315,N_44);
and U583 (N_583,In_452,In_1369);
or U584 (N_584,N_314,In_1825);
nor U585 (N_585,In_1858,N_248);
and U586 (N_586,In_858,In_661);
and U587 (N_587,In_1004,In_1584);
and U588 (N_588,N_301,In_856);
nand U589 (N_589,In_564,In_1074);
nand U590 (N_590,In_1097,In_1406);
xor U591 (N_591,N_94,N_36);
or U592 (N_592,In_443,N_234);
or U593 (N_593,N_149,N_124);
nor U594 (N_594,In_1612,In_1057);
nor U595 (N_595,In_1731,In_907);
or U596 (N_596,N_152,N_305);
or U597 (N_597,In_280,In_1847);
and U598 (N_598,In_18,N_78);
nor U599 (N_599,In_175,In_1054);
and U600 (N_600,N_11,N_320);
nand U601 (N_601,In_1087,In_1345);
nand U602 (N_602,In_685,In_1560);
or U603 (N_603,In_406,In_431);
nand U604 (N_604,N_368,N_41);
nand U605 (N_605,In_80,In_1490);
and U606 (N_606,In_1872,In_97);
and U607 (N_607,In_1971,N_212);
xnor U608 (N_608,In_681,N_59);
nand U609 (N_609,In_773,In_74);
and U610 (N_610,N_253,N_377);
and U611 (N_611,N_338,N_93);
or U612 (N_612,In_1181,N_272);
or U613 (N_613,In_597,In_1541);
xnor U614 (N_614,In_1130,In_1934);
and U615 (N_615,In_712,In_1961);
and U616 (N_616,In_7,In_181);
nand U617 (N_617,In_194,In_1826);
xor U618 (N_618,In_1930,In_1538);
or U619 (N_619,In_1700,In_1076);
or U620 (N_620,In_306,In_586);
and U621 (N_621,In_1794,N_286);
or U622 (N_622,In_26,In_1095);
or U623 (N_623,In_220,In_1641);
nor U624 (N_624,In_1264,In_1238);
or U625 (N_625,In_291,In_215);
nor U626 (N_626,In_1407,In_1636);
or U627 (N_627,In_1839,N_33);
nand U628 (N_628,In_155,In_770);
or U629 (N_629,N_49,N_106);
or U630 (N_630,N_322,In_222);
and U631 (N_631,In_1368,In_537);
xnor U632 (N_632,In_239,In_895);
nand U633 (N_633,N_378,N_182);
xnor U634 (N_634,In_818,In_3);
or U635 (N_635,In_278,In_868);
nand U636 (N_636,In_1328,N_243);
nor U637 (N_637,In_1720,In_1102);
nor U638 (N_638,In_965,In_66);
xnor U639 (N_639,In_1327,In_761);
and U640 (N_640,In_382,In_571);
and U641 (N_641,In_434,In_737);
xnor U642 (N_642,In_1229,In_1526);
xor U643 (N_643,N_326,N_211);
xor U644 (N_644,In_1464,In_1879);
or U645 (N_645,In_1505,In_1947);
xor U646 (N_646,In_388,In_1245);
or U647 (N_647,In_490,In_344);
nor U648 (N_648,N_8,In_904);
or U649 (N_649,In_106,N_34);
nor U650 (N_650,N_290,In_1357);
nand U651 (N_651,In_524,N_67);
nor U652 (N_652,N_210,In_1517);
nand U653 (N_653,In_253,N_70);
xor U654 (N_654,In_646,In_1415);
nand U655 (N_655,In_1136,In_615);
xor U656 (N_656,In_201,In_894);
nand U657 (N_657,In_1314,In_39);
and U658 (N_658,N_104,In_1592);
xnor U659 (N_659,In_1674,In_855);
nor U660 (N_660,N_17,N_275);
or U661 (N_661,N_223,N_71);
xor U662 (N_662,In_1211,In_491);
nor U663 (N_663,In_819,In_1710);
nand U664 (N_664,In_1622,In_1322);
nand U665 (N_665,In_1991,In_538);
and U666 (N_666,N_72,N_336);
nand U667 (N_667,In_1246,In_157);
or U668 (N_668,In_1859,In_1282);
nand U669 (N_669,In_968,N_2);
nand U670 (N_670,In_374,In_1111);
xor U671 (N_671,In_1857,In_1258);
and U672 (N_672,In_1711,In_47);
nor U673 (N_673,In_1865,N_116);
xor U674 (N_674,In_367,In_1911);
nand U675 (N_675,N_260,In_672);
and U676 (N_676,N_91,In_248);
or U677 (N_677,In_87,In_776);
nor U678 (N_678,In_1026,N_265);
nand U679 (N_679,In_1451,In_563);
xor U680 (N_680,N_342,In_84);
nor U681 (N_681,N_54,N_345);
and U682 (N_682,N_208,In_1730);
nand U683 (N_683,N_111,N_349);
or U684 (N_684,N_205,In_757);
or U685 (N_685,In_1444,In_1473);
and U686 (N_686,In_1249,In_783);
nor U687 (N_687,In_1206,N_96);
xnor U688 (N_688,N_346,In_364);
xor U689 (N_689,N_217,In_236);
nor U690 (N_690,N_82,In_281);
or U691 (N_691,N_388,In_675);
and U692 (N_692,N_231,In_1959);
or U693 (N_693,In_1999,In_705);
or U694 (N_694,N_40,In_1548);
nor U695 (N_695,N_296,In_1586);
nor U696 (N_696,N_192,In_1995);
and U697 (N_697,N_65,In_643);
nand U698 (N_698,In_1153,In_127);
nor U699 (N_699,In_683,In_992);
nor U700 (N_700,In_513,In_1555);
nand U701 (N_701,In_729,In_492);
xnor U702 (N_702,N_239,N_154);
nor U703 (N_703,In_81,In_580);
nor U704 (N_704,In_301,In_1093);
xor U705 (N_705,In_1488,In_1885);
and U706 (N_706,In_1595,In_440);
nand U707 (N_707,In_876,N_20);
nand U708 (N_708,In_1372,In_680);
or U709 (N_709,In_1856,In_749);
xor U710 (N_710,In_331,N_107);
or U711 (N_711,N_95,N_157);
or U712 (N_712,N_289,N_263);
and U713 (N_713,In_1117,In_1471);
and U714 (N_714,In_877,In_733);
and U715 (N_715,In_487,N_39);
and U716 (N_716,In_154,In_1986);
or U717 (N_717,In_1944,In_938);
xor U718 (N_718,In_1599,In_1670);
nor U719 (N_719,In_439,In_1367);
or U720 (N_720,N_327,In_1156);
or U721 (N_721,In_594,N_92);
and U722 (N_722,In_814,In_1836);
xnor U723 (N_723,In_42,In_1904);
and U724 (N_724,In_1236,In_328);
or U725 (N_725,In_481,In_0);
nand U726 (N_726,In_1382,In_1803);
or U727 (N_727,In_1907,In_1278);
nor U728 (N_728,In_1822,In_170);
or U729 (N_729,In_416,N_389);
and U730 (N_730,In_929,In_336);
xnor U731 (N_731,In_1300,N_264);
nor U732 (N_732,N_128,N_392);
nor U733 (N_733,In_1556,In_791);
and U734 (N_734,In_824,In_1736);
or U735 (N_735,In_1067,In_897);
nand U736 (N_736,In_286,In_1811);
and U737 (N_737,In_302,In_1926);
or U738 (N_738,In_477,In_489);
or U739 (N_739,In_1653,In_1734);
xnor U740 (N_740,N_119,N_292);
nor U741 (N_741,N_201,In_1377);
xor U742 (N_742,In_746,In_1818);
nand U743 (N_743,In_1905,N_13);
or U744 (N_744,In_599,In_816);
or U745 (N_745,N_261,N_21);
nor U746 (N_746,In_886,In_1142);
or U747 (N_747,In_1252,In_329);
nor U748 (N_748,In_1610,N_244);
nor U749 (N_749,In_365,N_255);
nand U750 (N_750,In_148,In_1767);
and U751 (N_751,In_345,N_369);
nand U752 (N_752,In_1077,In_151);
and U753 (N_753,In_993,In_1404);
nor U754 (N_754,N_218,In_441);
and U755 (N_755,In_1410,N_189);
and U756 (N_756,In_270,In_990);
or U757 (N_757,In_527,N_66);
xor U758 (N_758,In_1628,In_988);
nand U759 (N_759,N_164,In_1408);
xor U760 (N_760,In_1571,In_55);
or U761 (N_761,In_1247,In_1672);
xnor U762 (N_762,In_1807,In_109);
nor U763 (N_763,In_1942,N_262);
xnor U764 (N_764,N_372,In_206);
nor U765 (N_765,In_1970,N_350);
and U766 (N_766,In_865,In_100);
or U767 (N_767,In_360,In_463);
nand U768 (N_768,In_535,N_56);
nor U769 (N_769,In_1762,N_22);
nor U770 (N_770,In_1697,In_983);
and U771 (N_771,In_1623,In_122);
xor U772 (N_772,In_1694,In_207);
and U773 (N_773,In_424,In_427);
nor U774 (N_774,In_878,In_842);
or U775 (N_775,In_1871,In_1611);
xnor U776 (N_776,In_1660,In_1704);
nor U777 (N_777,N_257,In_1819);
nor U778 (N_778,N_298,In_916);
or U779 (N_779,In_997,In_699);
or U780 (N_780,N_113,N_52);
xnor U781 (N_781,In_1309,In_1913);
nand U782 (N_782,N_193,In_1750);
nand U783 (N_783,N_1,N_32);
xor U784 (N_784,In_1515,N_57);
xnor U785 (N_785,In_1159,N_361);
or U786 (N_786,In_1708,N_333);
xnor U787 (N_787,In_1590,In_361);
nand U788 (N_788,In_515,In_451);
xnor U789 (N_789,In_1295,N_181);
or U790 (N_790,In_305,N_269);
nand U791 (N_791,In_401,In_650);
and U792 (N_792,In_1161,In_639);
nand U793 (N_793,In_1167,In_1198);
nor U794 (N_794,N_68,In_1850);
nand U795 (N_795,In_1718,In_179);
nor U796 (N_796,In_340,In_525);
nor U797 (N_797,In_1786,In_1114);
and U798 (N_798,N_24,In_405);
xnor U799 (N_799,In_618,In_498);
or U800 (N_800,N_247,N_334);
and U801 (N_801,N_306,N_121);
nor U802 (N_802,In_1761,In_808);
xor U803 (N_803,N_431,N_697);
or U804 (N_804,In_1125,In_810);
xnor U805 (N_805,In_921,N_518);
xor U806 (N_806,In_1132,N_316);
xor U807 (N_807,N_767,N_752);
nor U808 (N_808,N_596,In_1753);
nand U809 (N_809,In_334,In_372);
and U810 (N_810,N_129,N_541);
nor U811 (N_811,N_741,N_559);
and U812 (N_812,In_1320,In_1494);
xnor U813 (N_813,N_434,In_1909);
and U814 (N_814,In_1534,In_1841);
xor U815 (N_815,N_564,In_249);
xor U816 (N_816,In_736,In_1401);
or U817 (N_817,In_813,In_959);
or U818 (N_818,In_1543,In_347);
nand U819 (N_819,N_528,In_1376);
xnor U820 (N_820,N_782,N_414);
xor U821 (N_821,N_707,In_86);
or U822 (N_822,In_129,N_198);
or U823 (N_823,In_716,N_46);
nor U824 (N_824,In_706,In_147);
nand U825 (N_825,N_371,N_754);
nor U826 (N_826,N_102,In_1129);
and U827 (N_827,In_1655,In_602);
and U828 (N_828,In_1446,N_593);
nor U829 (N_829,N_645,In_245);
xnor U830 (N_830,N_799,N_652);
and U831 (N_831,In_896,In_556);
nand U832 (N_832,N_449,N_12);
nand U833 (N_833,In_231,In_1103);
nor U834 (N_834,In_789,N_591);
or U835 (N_835,In_660,In_1861);
and U836 (N_836,N_717,N_532);
or U837 (N_837,N_420,N_183);
or U838 (N_838,In_28,In_626);
xor U839 (N_839,In_936,N_553);
and U840 (N_840,In_874,In_51);
and U841 (N_841,N_90,In_1049);
xnor U842 (N_842,N_685,In_202);
nor U843 (N_843,In_1452,In_1503);
and U844 (N_844,N_695,In_9);
and U845 (N_845,N_490,N_738);
xor U846 (N_846,N_427,In_1476);
nor U847 (N_847,In_1888,In_689);
xnor U848 (N_848,N_797,In_1654);
and U849 (N_849,In_1143,In_859);
xor U850 (N_850,In_1189,In_57);
nand U851 (N_851,N_638,In_543);
xor U852 (N_852,In_103,N_614);
nand U853 (N_853,N_587,In_944);
nand U854 (N_854,In_1679,N_339);
nor U855 (N_855,In_386,N_482);
or U856 (N_856,N_665,In_698);
nand U857 (N_857,N_778,N_577);
nand U858 (N_858,N_771,N_648);
xnor U859 (N_859,N_565,N_299);
and U860 (N_860,N_403,In_1906);
and U861 (N_861,N_387,N_213);
nand U862 (N_862,N_62,N_590);
or U863 (N_863,In_1253,N_691);
xor U864 (N_864,In_1261,N_798);
xnor U865 (N_865,N_452,In_507);
nand U866 (N_866,N_630,In_1233);
nor U867 (N_867,N_537,In_318);
nand U868 (N_868,N_221,In_113);
nor U869 (N_869,N_84,N_765);
nand U870 (N_870,In_1194,In_1013);
or U871 (N_871,N_373,In_370);
nor U872 (N_872,In_1362,In_1566);
or U873 (N_873,In_453,In_1485);
nand U874 (N_874,In_1897,In_309);
xnor U875 (N_875,In_1348,In_595);
and U876 (N_876,N_220,In_1964);
xor U877 (N_877,In_1421,In_102);
or U878 (N_878,In_1002,In_579);
nand U879 (N_879,In_1003,In_1793);
and U880 (N_880,N_433,In_1298);
or U881 (N_881,In_1073,In_1151);
nor U882 (N_882,N_576,N_254);
nand U883 (N_883,N_200,In_1216);
nor U884 (N_884,In_1096,In_1123);
and U885 (N_885,N_138,In_794);
xor U886 (N_886,In_1259,N_654);
and U887 (N_887,N_612,N_225);
xor U888 (N_888,N_483,N_405);
xor U889 (N_889,N_555,N_525);
and U890 (N_890,N_572,In_1701);
or U891 (N_891,In_79,N_758);
nand U892 (N_892,N_558,In_1992);
and U893 (N_893,N_478,In_1277);
xnor U894 (N_894,N_469,In_1981);
nand U895 (N_895,N_398,In_1268);
nand U896 (N_896,N_423,In_105);
xor U897 (N_897,In_1242,In_1046);
or U898 (N_898,N_250,N_677);
and U899 (N_899,In_289,In_186);
xnor U900 (N_900,In_956,N_520);
or U901 (N_901,N_459,N_592);
or U902 (N_902,In_671,In_41);
and U903 (N_903,In_613,In_966);
or U904 (N_904,In_1752,In_730);
nor U905 (N_905,In_931,N_772);
and U906 (N_906,In_1742,N_487);
xor U907 (N_907,In_1347,In_116);
and U908 (N_908,In_456,In_1431);
nand U909 (N_909,N_701,In_255);
or U910 (N_910,In_1124,N_19);
xor U911 (N_911,In_1441,N_105);
xor U912 (N_912,N_672,N_633);
and U913 (N_913,N_660,N_29);
nand U914 (N_914,N_611,In_1179);
and U915 (N_915,N_498,N_199);
and U916 (N_916,N_309,N_325);
nand U917 (N_917,In_740,N_712);
nor U918 (N_918,In_1849,In_1960);
and U919 (N_919,N_763,In_421);
nand U920 (N_920,In_1563,In_89);
and U921 (N_921,N_461,N_158);
and U922 (N_922,N_747,In_191);
or U923 (N_923,In_780,In_238);
xnor U924 (N_924,In_1169,In_1432);
and U925 (N_925,N_444,N_533);
xor U926 (N_926,In_1036,In_1575);
xor U927 (N_927,N_60,N_664);
xnor U928 (N_928,N_130,In_1754);
nor U929 (N_929,In_1089,In_363);
nor U930 (N_930,In_31,In_512);
and U931 (N_931,In_1778,In_1341);
xnor U932 (N_932,N_675,In_854);
xnor U933 (N_933,N_209,N_616);
nand U934 (N_934,In_192,In_629);
nand U935 (N_935,N_643,N_521);
xor U936 (N_936,N_728,N_115);
nand U937 (N_937,N_538,In_1706);
nor U938 (N_938,N_233,In_1005);
and U939 (N_939,N_400,N_356);
or U940 (N_940,In_56,In_230);
nand U941 (N_941,N_472,In_1360);
nand U942 (N_942,N_535,N_457);
or U943 (N_943,In_696,N_117);
and U944 (N_944,In_323,N_442);
nand U945 (N_945,N_471,N_523);
or U946 (N_946,N_760,In_1798);
xnor U947 (N_947,In_771,N_273);
or U948 (N_948,In_1953,In_1634);
nand U949 (N_949,In_326,N_703);
nand U950 (N_950,In_576,N_284);
and U951 (N_951,N_756,N_271);
or U952 (N_952,N_10,N_456);
or U953 (N_953,In_343,In_1851);
and U954 (N_954,N_390,In_377);
nor U955 (N_955,In_320,N_766);
xor U956 (N_956,N_622,N_506);
xnor U957 (N_957,N_618,In_1724);
nor U958 (N_958,In_664,In_1483);
nand U959 (N_959,In_247,N_28);
nand U960 (N_960,N_170,In_1866);
xnor U961 (N_961,In_1962,In_1254);
xnor U962 (N_962,In_13,In_1757);
nor U963 (N_963,In_682,In_1740);
nand U964 (N_964,N_702,In_1693);
nor U965 (N_965,In_5,In_517);
xnor U966 (N_966,N_364,N_636);
xnor U967 (N_967,N_463,N_793);
xnor U968 (N_968,In_1790,In_476);
and U969 (N_969,N_42,In_264);
or U970 (N_970,N_507,In_1901);
or U971 (N_971,N_435,N_464);
or U972 (N_972,N_503,N_620);
xnor U973 (N_973,In_314,In_1475);
or U974 (N_974,In_688,In_724);
nor U975 (N_975,In_135,N_45);
xnor U976 (N_976,In_1891,N_556);
nor U977 (N_977,In_523,N_549);
or U978 (N_978,In_385,In_1696);
or U979 (N_979,In_964,In_295);
xnor U980 (N_980,In_1434,In_254);
nand U981 (N_981,In_1771,N_495);
nor U982 (N_982,In_1342,N_779);
nor U983 (N_983,N_686,N_745);
xor U984 (N_984,N_588,N_165);
or U985 (N_985,In_549,In_1134);
and U986 (N_986,N_476,In_418);
nand U987 (N_987,In_1349,In_1397);
or U988 (N_988,N_303,N_358);
nand U989 (N_989,In_1426,N_428);
nand U990 (N_990,In_1863,N_35);
nor U991 (N_991,N_794,In_624);
xnor U992 (N_992,In_899,In_801);
nor U993 (N_993,In_408,In_1105);
nand U994 (N_994,N_608,In_713);
or U995 (N_995,In_437,N_458);
nor U996 (N_996,N_406,In_1256);
and U997 (N_997,In_551,In_994);
or U998 (N_998,N_236,N_705);
nand U999 (N_999,N_408,N_748);
and U1000 (N_1000,N_173,In_569);
or U1001 (N_1001,N_768,In_1204);
and U1002 (N_1002,In_1048,N_582);
and U1003 (N_1003,N_450,N_749);
nand U1004 (N_1004,In_900,In_1175);
xnor U1005 (N_1005,N_580,N_775);
xor U1006 (N_1006,N_653,N_784);
nand U1007 (N_1007,N_678,In_1061);
or U1008 (N_1008,N_185,In_750);
nand U1009 (N_1009,In_1109,In_621);
nand U1010 (N_1010,In_725,N_222);
xnor U1011 (N_1011,In_1332,N_120);
nor U1012 (N_1012,N_110,In_1927);
and U1013 (N_1013,N_224,In_1852);
xnor U1014 (N_1014,N_16,In_69);
or U1015 (N_1015,In_1721,In_107);
and U1016 (N_1016,In_781,N_729);
nor U1017 (N_1017,In_1846,In_1765);
nor U1018 (N_1018,N_597,In_834);
xor U1019 (N_1019,In_1027,N_246);
xnor U1020 (N_1020,In_339,In_1542);
nor U1021 (N_1021,N_203,N_578);
and U1022 (N_1022,In_1336,N_789);
nand U1023 (N_1023,N_480,N_351);
nand U1024 (N_1024,N_762,In_1235);
or U1025 (N_1025,In_470,In_1333);
xnor U1026 (N_1026,N_288,In_1967);
nor U1027 (N_1027,N_395,N_531);
and U1028 (N_1028,N_114,In_784);
and U1029 (N_1029,In_1023,In_704);
xnor U1030 (N_1030,In_995,N_674);
nor U1031 (N_1031,In_1977,N_50);
xnor U1032 (N_1032,In_927,In_1215);
or U1033 (N_1033,In_1528,N_391);
nor U1034 (N_1034,In_1038,In_156);
or U1035 (N_1035,N_603,In_1564);
nand U1036 (N_1036,In_290,N_493);
nor U1037 (N_1037,In_288,N_517);
xor U1038 (N_1038,N_477,N_750);
nor U1039 (N_1039,In_252,N_724);
or U1040 (N_1040,N_313,In_598);
xor U1041 (N_1041,N_422,N_623);
nand U1042 (N_1042,In_1092,N_550);
nand U1043 (N_1043,In_1759,N_732);
and U1044 (N_1044,In_82,N_621);
and U1045 (N_1045,N_619,In_1186);
nand U1046 (N_1046,N_787,N_500);
nand U1047 (N_1047,N_631,N_609);
nor U1048 (N_1048,In_1809,In_835);
nand U1049 (N_1049,In_1955,In_1387);
xnor U1050 (N_1050,N_722,In_984);
nor U1051 (N_1051,In_1552,In_1898);
nand U1052 (N_1052,N_505,In_1435);
nand U1053 (N_1053,N_347,In_1160);
or U1054 (N_1054,In_61,In_849);
xnor U1055 (N_1055,N_670,N_481);
xnor U1056 (N_1056,In_658,In_1006);
or U1057 (N_1057,In_1458,N_278);
xnor U1058 (N_1058,N_781,In_92);
nor U1059 (N_1059,In_53,N_466);
or U1060 (N_1060,N_283,N_719);
xnor U1061 (N_1061,In_120,In_529);
xnor U1062 (N_1062,In_461,N_598);
and U1063 (N_1063,In_1800,N_401);
and U1064 (N_1064,In_655,In_1669);
and U1065 (N_1065,N_376,N_492);
nor U1066 (N_1066,In_540,N_690);
nor U1067 (N_1067,N_417,N_63);
or U1068 (N_1068,In_83,In_1683);
or U1069 (N_1069,In_593,N_355);
nand U1070 (N_1070,In_368,In_617);
nor U1071 (N_1071,N_514,N_337);
or U1072 (N_1072,In_1187,N_276);
xnor U1073 (N_1073,In_1230,N_108);
and U1074 (N_1074,N_713,In_77);
xor U1075 (N_1075,N_166,N_126);
and U1076 (N_1076,In_1644,N_100);
nor U1077 (N_1077,In_932,In_1626);
xnor U1078 (N_1078,In_1273,N_667);
xnor U1079 (N_1079,N_693,In_104);
xnor U1080 (N_1080,In_731,N_366);
xor U1081 (N_1081,N_468,N_585);
xor U1082 (N_1082,N_744,In_922);
nor U1083 (N_1083,In_1240,In_1207);
nor U1084 (N_1084,N_467,N_715);
nor U1085 (N_1085,In_1747,In_754);
xor U1086 (N_1086,In_526,N_683);
nand U1087 (N_1087,N_796,N_600);
and U1088 (N_1088,In_1935,In_1624);
xnor U1089 (N_1089,N_226,In_1788);
xor U1090 (N_1090,In_1052,N_563);
nor U1091 (N_1091,In_1813,In_1530);
xor U1092 (N_1092,In_1243,N_411);
xnor U1093 (N_1093,In_1504,N_293);
xnor U1094 (N_1094,N_709,In_183);
xnor U1095 (N_1095,N_776,In_32);
or U1096 (N_1096,In_1325,N_562);
or U1097 (N_1097,In_637,In_1399);
xor U1098 (N_1098,In_91,N_711);
nand U1099 (N_1099,In_1050,In_1436);
or U1100 (N_1100,In_634,In_888);
or U1101 (N_1101,N_682,N_31);
or U1102 (N_1102,In_139,N_219);
or U1103 (N_1103,N_595,In_825);
or U1104 (N_1104,N_634,N_9);
or U1105 (N_1105,N_792,N_274);
or U1106 (N_1106,In_203,N_324);
nor U1107 (N_1107,In_1652,N_661);
or U1108 (N_1108,N_757,N_357);
or U1109 (N_1109,N_625,N_570);
nor U1110 (N_1110,In_619,In_663);
nor U1111 (N_1111,N_557,N_714);
or U1112 (N_1112,N_502,In_1442);
nand U1113 (N_1113,N_718,N_419);
or U1114 (N_1114,In_429,In_1065);
nor U1115 (N_1115,N_81,N_604);
and U1116 (N_1116,In_827,In_1155);
nand U1117 (N_1117,In_1384,In_1616);
xor U1118 (N_1118,In_603,N_773);
nand U1119 (N_1119,In_1875,N_421);
nor U1120 (N_1120,N_241,N_496);
or U1121 (N_1121,In_216,N_737);
and U1122 (N_1122,In_256,N_710);
and U1123 (N_1123,In_1,In_1638);
and U1124 (N_1124,In_970,N_160);
nor U1125 (N_1125,In_335,In_797);
or U1126 (N_1126,N_699,In_852);
or U1127 (N_1127,In_1457,In_1141);
nand U1128 (N_1128,N_429,In_1480);
or U1129 (N_1129,N_242,N_554);
and U1130 (N_1130,N_430,N_453);
and U1131 (N_1131,N_560,In_1810);
and U1132 (N_1132,In_774,In_1637);
xor U1133 (N_1133,In_1419,In_276);
nor U1134 (N_1134,N_359,In_1280);
and U1135 (N_1135,In_479,N_751);
and U1136 (N_1136,In_786,N_386);
nand U1137 (N_1137,N_540,N_510);
or U1138 (N_1138,In_1958,N_74);
nand U1139 (N_1139,N_688,In_45);
xnor U1140 (N_1140,In_464,N_399);
and U1141 (N_1141,In_860,In_654);
and U1142 (N_1142,In_457,N_38);
or U1143 (N_1143,N_321,N_606);
or U1144 (N_1144,In_1899,N_526);
or U1145 (N_1145,N_415,In_467);
or U1146 (N_1146,N_252,N_375);
xor U1147 (N_1147,In_1218,N_679);
xnor U1148 (N_1148,In_727,N_668);
nor U1149 (N_1149,N_669,N_88);
nand U1150 (N_1150,In_809,In_1051);
nor U1151 (N_1151,In_177,In_1501);
nand U1152 (N_1152,N_575,N_494);
or U1153 (N_1153,In_240,N_86);
xor U1154 (N_1154,N_545,N_515);
nand U1155 (N_1155,N_27,In_648);
nor U1156 (N_1156,N_567,N_484);
xor U1157 (N_1157,N_317,In_1666);
xor U1158 (N_1158,In_1689,In_1685);
or U1159 (N_1159,N_640,N_519);
and U1160 (N_1160,In_196,N_485);
and U1161 (N_1161,N_599,N_451);
nor U1162 (N_1162,N_470,In_719);
xor U1163 (N_1163,N_251,In_1466);
xor U1164 (N_1164,In_138,N_237);
and U1165 (N_1165,N_551,N_462);
or U1166 (N_1166,In_38,N_627);
or U1167 (N_1167,N_245,In_465);
nor U1168 (N_1168,N_607,In_210);
nand U1169 (N_1169,In_20,N_370);
nor U1170 (N_1170,In_631,N_465);
nor U1171 (N_1171,N_524,N_175);
nand U1172 (N_1172,N_48,In_1508);
or U1173 (N_1173,In_1723,In_460);
nor U1174 (N_1174,N_441,N_240);
nor U1175 (N_1175,N_646,In_324);
nor U1176 (N_1176,In_1843,In_1716);
nor U1177 (N_1177,N_123,In_534);
or U1178 (N_1178,In_755,In_1551);
nor U1179 (N_1179,In_284,In_622);
nor U1180 (N_1180,In_1499,N_671);
xnor U1181 (N_1181,In_908,In_508);
nand U1182 (N_1182,In_1030,In_214);
and U1183 (N_1183,N_409,In_1139);
xnor U1184 (N_1184,N_742,N_783);
nand U1185 (N_1185,In_1993,In_362);
nor U1186 (N_1186,N_662,N_445);
nand U1187 (N_1187,N_425,In_657);
nand U1188 (N_1188,N_692,In_1732);
nand U1189 (N_1189,N_163,N_380);
or U1190 (N_1190,N_569,N_513);
xnor U1191 (N_1191,In_1497,In_1783);
nand U1192 (N_1192,N_53,In_163);
nor U1193 (N_1193,N_579,N_573);
nand U1194 (N_1194,In_851,In_941);
xor U1195 (N_1195,N_488,N_497);
xnor U1196 (N_1196,N_179,In_1440);
or U1197 (N_1197,In_6,N_137);
or U1198 (N_1198,N_736,N_536);
nand U1199 (N_1199,N_740,In_503);
xnor U1200 (N_1200,N_969,N_1021);
and U1201 (N_1201,N_1131,In_1998);
nand U1202 (N_1202,In_919,N_1111);
or U1203 (N_1203,N_1175,N_864);
nand U1204 (N_1204,N_642,In_1651);
or U1205 (N_1205,N_1009,In_659);
xor U1206 (N_1206,In_90,In_1291);
or U1207 (N_1207,In_1835,N_974);
xor U1208 (N_1208,N_1025,N_658);
nand U1209 (N_1209,N_852,N_940);
nor U1210 (N_1210,N_508,N_1196);
and U1211 (N_1211,In_1083,N_1053);
xor U1212 (N_1212,In_412,N_819);
nor U1213 (N_1213,N_511,N_930);
or U1214 (N_1214,In_395,N_739);
and U1215 (N_1215,N_552,N_1070);
or U1216 (N_1216,N_172,N_285);
nor U1217 (N_1217,N_1084,N_1094);
xor U1218 (N_1218,In_271,N_436);
nor U1219 (N_1219,N_310,N_426);
or U1220 (N_1220,N_190,N_816);
nand U1221 (N_1221,N_412,N_918);
and U1222 (N_1222,N_649,N_1080);
nor U1223 (N_1223,N_1180,N_859);
xnor U1224 (N_1224,N_227,N_952);
and U1225 (N_1225,N_1093,N_1079);
or U1226 (N_1226,N_207,In_1577);
or U1227 (N_1227,N_730,N_1062);
xor U1228 (N_1228,N_982,N_983);
nor U1229 (N_1229,N_946,N_810);
and U1230 (N_1230,In_1063,N_1044);
xor U1231 (N_1231,N_509,N_1082);
nor U1232 (N_1232,N_964,N_601);
or U1233 (N_1233,N_1029,N_1075);
nor U1234 (N_1234,In_1573,In_213);
nand U1235 (N_1235,In_1343,N_999);
and U1236 (N_1236,N_1099,In_1212);
or U1237 (N_1237,N_1127,N_543);
xnor U1238 (N_1238,In_391,N_924);
or U1239 (N_1239,N_840,N_681);
xnor U1240 (N_1240,N_544,N_884);
and U1241 (N_1241,In_1127,N_851);
nor U1242 (N_1242,N_656,N_998);
nand U1243 (N_1243,N_7,N_944);
xor U1244 (N_1244,N_1141,N_786);
nand U1245 (N_1245,N_1121,In_1987);
nor U1246 (N_1246,N_416,In_940);
nor U1247 (N_1247,N_1007,N_1078);
or U1248 (N_1248,N_396,N_805);
xnor U1249 (N_1249,N_454,N_1167);
or U1250 (N_1250,N_655,N_1161);
and U1251 (N_1251,N_103,N_725);
nor U1252 (N_1252,N_1124,N_882);
nand U1253 (N_1253,N_726,N_1182);
nor U1254 (N_1254,N_791,In_1580);
xnor U1255 (N_1255,N_959,N_1152);
or U1256 (N_1256,In_1936,N_888);
and U1257 (N_1257,N_1166,N_843);
or U1258 (N_1258,N_863,In_1286);
nand U1259 (N_1259,In_1760,In_1924);
nor U1260 (N_1260,In_1126,N_953);
nor U1261 (N_1261,In_1853,N_1132);
and U1262 (N_1262,N_424,N_148);
xnor U1263 (N_1263,N_1050,In_1433);
nand U1264 (N_1264,N_929,N_774);
nor U1265 (N_1265,N_684,N_916);
nor U1266 (N_1266,N_432,N_1037);
or U1267 (N_1267,N_881,In_999);
nor U1268 (N_1268,In_1203,N_1155);
and U1269 (N_1269,In_934,N_909);
and U1270 (N_1270,N_910,N_837);
xnor U1271 (N_1271,In_583,N_1150);
xnor U1272 (N_1272,In_1519,N_942);
xor U1273 (N_1273,N_904,N_827);
xor U1274 (N_1274,N_1091,N_76);
and U1275 (N_1275,N_159,N_753);
nor U1276 (N_1276,N_777,N_1011);
nand U1277 (N_1277,N_1140,N_1147);
or U1278 (N_1278,In_1791,N_1012);
and U1279 (N_1279,N_876,In_822);
xor U1280 (N_1280,N_501,N_1162);
and U1281 (N_1281,N_804,N_1085);
nand U1282 (N_1282,N_287,N_955);
nand U1283 (N_1283,N_1103,N_1163);
nor U1284 (N_1284,In_1094,N_1038);
and U1285 (N_1285,N_1164,N_817);
nand U1286 (N_1286,N_770,N_854);
nor U1287 (N_1287,N_1006,N_215);
or U1288 (N_1288,In_1868,In_375);
or U1289 (N_1289,N_694,In_947);
xor U1290 (N_1290,N_404,N_860);
or U1291 (N_1291,N_1005,N_546);
nand U1292 (N_1292,N_1023,N_1031);
nor U1293 (N_1293,N_258,N_1069);
nor U1294 (N_1294,N_1188,N_574);
nor U1295 (N_1295,In_1173,N_1126);
xor U1296 (N_1296,N_610,N_605);
xor U1297 (N_1297,N_1186,N_644);
and U1298 (N_1298,N_1170,N_499);
or U1299 (N_1299,N_584,In_1346);
and U1300 (N_1300,N_1125,In_883);
nand U1301 (N_1301,N_302,N_534);
nand U1302 (N_1302,In_967,N_1119);
or U1303 (N_1303,N_720,N_1059);
or U1304 (N_1304,In_1149,N_639);
nand U1305 (N_1305,In_445,N_184);
nand U1306 (N_1306,In_358,N_1106);
and U1307 (N_1307,N_1173,In_1220);
nand U1308 (N_1308,In_407,N_1081);
or U1309 (N_1309,N_979,In_1292);
nor U1310 (N_1310,N_109,N_101);
or U1311 (N_1311,N_529,N_479);
nand U1312 (N_1312,N_594,N_917);
xnor U1313 (N_1313,In_1183,N_474);
nand U1314 (N_1314,N_385,N_530);
nand U1315 (N_1315,N_1199,In_690);
and U1316 (N_1316,N_1197,N_903);
and U1317 (N_1317,N_841,In_282);
nor U1318 (N_1318,In_562,N_1159);
nor U1319 (N_1319,N_216,In_802);
and U1320 (N_1320,N_177,In_960);
or U1321 (N_1321,N_1022,N_1129);
or U1322 (N_1322,N_986,N_583);
xor U1323 (N_1323,N_280,N_1158);
or U1324 (N_1324,N_1073,N_1143);
or U1325 (N_1325,N_1067,N_1156);
xnor U1326 (N_1326,N_992,N_997);
or U1327 (N_1327,N_1077,In_134);
nor U1328 (N_1328,In_1324,N_489);
xnor U1329 (N_1329,N_721,In_656);
nor U1330 (N_1330,N_780,N_920);
xor U1331 (N_1331,N_1100,N_850);
nand U1332 (N_1332,N_1060,N_1071);
xor U1333 (N_1333,N_1034,N_764);
and U1334 (N_1334,In_1165,N_1168);
nor U1335 (N_1335,N_912,N_1136);
or U1336 (N_1336,N_134,N_1055);
and U1337 (N_1337,N_80,N_125);
or U1338 (N_1338,N_708,N_761);
nand U1339 (N_1339,N_1051,N_948);
xnor U1340 (N_1340,N_1108,In_262);
nor U1341 (N_1341,N_977,N_1015);
nand U1342 (N_1342,N_808,N_987);
nand U1343 (N_1343,N_821,N_1145);
xnor U1344 (N_1344,In_1895,N_1148);
and U1345 (N_1345,N_976,N_602);
nor U1346 (N_1346,N_900,N_885);
or U1347 (N_1347,In_1688,N_1076);
or U1348 (N_1348,N_1104,N_676);
or U1349 (N_1349,N_889,N_1181);
nand U1350 (N_1350,N_696,In_1741);
nand U1351 (N_1351,N_996,In_1943);
nand U1352 (N_1352,N_991,N_69);
and U1353 (N_1353,N_1032,N_950);
and U1354 (N_1354,N_440,N_214);
xor U1355 (N_1355,In_348,N_704);
nand U1356 (N_1356,N_1138,N_866);
nand U1357 (N_1357,In_606,In_1902);
and U1358 (N_1358,N_628,N_800);
and U1359 (N_1359,N_1171,N_921);
or U1360 (N_1360,In_863,N_994);
xor U1361 (N_1361,N_949,In_884);
and U1362 (N_1362,In_889,N_5);
nand U1363 (N_1363,In_1301,N_1153);
or U1364 (N_1364,In_917,N_1184);
and U1365 (N_1365,N_97,N_438);
xor U1366 (N_1366,N_886,N_973);
or U1367 (N_1367,In_1500,In_1581);
xnor U1368 (N_1368,N_689,N_893);
nand U1369 (N_1369,N_872,N_1013);
nand U1370 (N_1370,N_1033,N_947);
and U1371 (N_1371,N_801,N_836);
nand U1372 (N_1372,N_931,N_1185);
nand U1373 (N_1373,N_626,N_919);
xnor U1374 (N_1374,N_960,N_1193);
nor U1375 (N_1375,N_906,N_680);
nor U1376 (N_1376,N_1090,N_522);
nand U1377 (N_1377,N_965,N_1039);
or U1378 (N_1378,N_1010,N_883);
xnor U1379 (N_1379,N_911,In_1714);
xor U1380 (N_1380,N_1117,N_1028);
nor U1381 (N_1381,N_666,In_1226);
and U1382 (N_1382,N_402,N_1183);
nor U1383 (N_1383,N_1146,N_928);
and U1384 (N_1384,In_913,N_941);
nand U1385 (N_1385,N_807,In_59);
or U1386 (N_1386,N_1179,N_1190);
and U1387 (N_1387,In_1032,N_1017);
or U1388 (N_1388,N_895,N_897);
nand U1389 (N_1389,N_1026,N_1118);
xor U1390 (N_1390,N_1110,In_1928);
and U1391 (N_1391,In_308,N_140);
nand U1392 (N_1392,N_1154,N_1096);
nand U1393 (N_1393,N_1174,N_844);
nand U1394 (N_1394,In_1447,In_669);
or U1395 (N_1395,N_943,N_769);
nor U1396 (N_1396,N_790,N_913);
nor U1397 (N_1397,N_1133,N_99);
xor U1398 (N_1398,N_1137,N_868);
nand U1399 (N_1399,N_1043,In_76);
or U1400 (N_1400,N_818,In_500);
and U1401 (N_1401,N_281,N_1097);
or U1402 (N_1402,N_617,In_455);
nand U1403 (N_1403,N_878,In_505);
nor U1404 (N_1404,N_962,In_596);
nand U1405 (N_1405,N_1191,In_197);
nand U1406 (N_1406,N_1194,In_986);
nand U1407 (N_1407,N_647,N_1000);
nand U1408 (N_1408,N_1151,In_1171);
or U1409 (N_1409,N_1101,N_1112);
and U1410 (N_1410,N_814,N_839);
xor U1411 (N_1411,N_812,N_823);
nand U1412 (N_1412,N_894,N_825);
or U1413 (N_1413,N_1018,N_344);
xnor U1414 (N_1414,In_118,In_378);
xnor U1415 (N_1415,N_397,In_304);
xnor U1416 (N_1416,N_1128,In_898);
or U1417 (N_1417,N_615,N_813);
nand U1418 (N_1418,N_802,N_571);
xor U1419 (N_1419,In_803,N_194);
nor U1420 (N_1420,In_471,In_1122);
or U1421 (N_1421,N_629,N_957);
and U1422 (N_1422,N_835,N_1061);
nand U1423 (N_1423,N_659,N_235);
nor U1424 (N_1424,N_899,N_143);
xor U1425 (N_1425,N_539,N_958);
nor U1426 (N_1426,N_858,In_224);
xnor U1427 (N_1427,N_295,In_1131);
nand U1428 (N_1428,N_873,In_748);
nand U1429 (N_1429,N_990,N_809);
nor U1430 (N_1430,In_670,N_410);
and U1431 (N_1431,N_1003,In_1037);
or U1432 (N_1432,N_1134,In_969);
and U1433 (N_1433,N_657,In_1389);
or U1434 (N_1434,N_988,N_1120);
and U1435 (N_1435,N_1068,N_993);
and U1436 (N_1436,N_1123,N_18);
nor U1437 (N_1437,N_985,N_936);
nand U1438 (N_1438,N_228,N_923);
nor U1439 (N_1439,In_1396,In_1313);
xnor U1440 (N_1440,N_795,In_394);
or U1441 (N_1441,N_1114,N_933);
and U1442 (N_1442,N_1072,N_833);
or U1443 (N_1443,In_1647,N_382);
nand U1444 (N_1444,N_55,In_1395);
xnor U1445 (N_1445,In_1470,N_820);
xnor U1446 (N_1446,N_512,In_1228);
nor U1447 (N_1447,In_169,N_1144);
and U1448 (N_1448,In_1213,In_200);
or U1449 (N_1449,N_845,N_448);
nor U1450 (N_1450,N_187,N_151);
or U1451 (N_1451,N_1089,In_376);
and U1452 (N_1452,N_865,N_407);
and U1453 (N_1453,N_862,N_869);
xnor U1454 (N_1454,In_180,N_1054);
nor U1455 (N_1455,N_945,N_1016);
and U1456 (N_1456,N_934,N_64);
nor U1457 (N_1457,In_805,In_1915);
nor U1458 (N_1458,In_1806,In_446);
or U1459 (N_1459,N_890,N_842);
nor U1460 (N_1460,In_448,N_1004);
nor U1461 (N_1461,N_963,N_1169);
nand U1462 (N_1462,In_133,N_828);
or U1463 (N_1463,N_824,In_1412);
and U1464 (N_1464,N_637,N_330);
nand U1465 (N_1465,N_811,N_491);
nor U1466 (N_1466,N_731,N_516);
xnor U1467 (N_1467,N_455,In_926);
or U1468 (N_1468,In_1916,N_1198);
nand U1469 (N_1469,N_204,N_1088);
or U1470 (N_1470,N_142,N_1107);
and U1471 (N_1471,In_193,N_527);
nand U1472 (N_1472,N_650,N_901);
xnor U1473 (N_1473,N_847,N_1001);
xor U1474 (N_1474,In_218,N_907);
nand U1475 (N_1475,N_413,N_1177);
nor U1476 (N_1476,N_831,In_692);
xor U1477 (N_1477,N_1056,N_277);
nor U1478 (N_1478,In_1393,N_815);
and U1479 (N_1479,N_733,N_874);
nand U1480 (N_1480,N_613,N_1087);
nor U1481 (N_1481,N_641,N_848);
nor U1482 (N_1482,N_394,N_1113);
and U1483 (N_1483,N_938,N_635);
or U1484 (N_1484,N_1057,N_1019);
or U1485 (N_1485,N_984,N_743);
nand U1486 (N_1486,In_1214,N_624);
or U1487 (N_1487,In_1034,N_446);
nor U1488 (N_1488,N_651,N_803);
nor U1489 (N_1489,In_1135,N_1109);
nand U1490 (N_1490,N_896,In_1892);
nand U1491 (N_1491,N_785,In_933);
and U1492 (N_1492,N_133,In_559);
nor U1493 (N_1493,N_566,In_1323);
nand U1494 (N_1494,N_935,N_561);
xor U1495 (N_1495,In_474,In_342);
nor U1496 (N_1496,In_910,N_834);
or U1497 (N_1497,N_967,N_1040);
nor U1498 (N_1498,N_856,N_1046);
xor U1499 (N_1499,N_568,N_875);
or U1500 (N_1500,In_149,N_981);
and U1501 (N_1501,N_880,N_486);
nor U1502 (N_1502,N_1142,N_975);
xnor U1503 (N_1503,N_153,N_956);
xnor U1504 (N_1504,N_1024,N_970);
xnor U1505 (N_1505,N_1047,N_1052);
nor U1506 (N_1506,N_788,N_1058);
or U1507 (N_1507,In_433,N_908);
or U1508 (N_1508,N_1095,N_381);
and U1509 (N_1509,In_173,N_846);
and U1510 (N_1510,N_504,N_968);
xor U1511 (N_1511,N_989,N_951);
xor U1512 (N_1512,N_437,N_870);
nor U1513 (N_1513,N_887,N_830);
and U1514 (N_1514,N_914,N_1187);
nor U1515 (N_1515,N_1098,N_297);
nor U1516 (N_1516,In_1460,In_444);
or U1517 (N_1517,In_1190,In_957);
nor U1518 (N_1518,N_1066,In_769);
and U1519 (N_1519,N_1049,N_853);
nand U1520 (N_1520,In_1221,N_1041);
or U1521 (N_1521,In_775,N_898);
or U1522 (N_1522,N_1030,N_1074);
xnor U1523 (N_1523,N_673,N_927);
xor U1524 (N_1524,N_980,N_418);
xor U1525 (N_1525,N_460,N_14);
or U1526 (N_1526,In_292,N_829);
xor U1527 (N_1527,N_1195,In_1459);
and U1528 (N_1528,In_506,In_1477);
nand U1529 (N_1529,N_1122,In_1311);
xnor U1530 (N_1530,N_1139,N_341);
or U1531 (N_1531,N_755,In_1107);
xor U1532 (N_1532,N_1014,In_1795);
and U1533 (N_1533,In_1945,N_932);
and U1534 (N_1534,N_1002,In_651);
nand U1535 (N_1535,In_953,N_939);
nor U1536 (N_1536,N_698,N_1115);
xor U1537 (N_1537,In_885,In_1355);
or U1538 (N_1538,In_799,N_542);
nor U1539 (N_1539,N_832,In_760);
xnor U1540 (N_1540,N_1063,N_475);
nand U1541 (N_1541,In_165,In_1889);
xor U1542 (N_1542,N_838,In_36);
nand U1543 (N_1543,N_1042,N_196);
nor U1544 (N_1544,N_877,N_473);
or U1545 (N_1545,N_915,N_1092);
or U1546 (N_1546,N_1149,In_1086);
and U1547 (N_1547,In_50,N_972);
and U1548 (N_1548,N_1165,N_1105);
or U1549 (N_1549,N_922,In_1598);
xnor U1550 (N_1550,N_954,N_806);
nor U1551 (N_1551,In_627,In_1297);
and U1552 (N_1552,N_902,In_423);
or U1553 (N_1553,N_1027,In_958);
xor U1554 (N_1554,N_1064,In_1414);
nor U1555 (N_1555,In_185,In_1370);
nand U1556 (N_1556,In_652,N_723);
xor U1557 (N_1557,N_229,N_1083);
nor U1558 (N_1558,N_735,N_746);
nor U1559 (N_1559,N_1172,In_1766);
and U1560 (N_1560,N_663,N_822);
and U1561 (N_1561,N_1157,N_43);
nand U1562 (N_1562,N_905,In_1692);
xor U1563 (N_1563,N_1048,N_926);
xnor U1564 (N_1564,N_727,N_700);
nor U1565 (N_1565,N_300,N_849);
nor U1566 (N_1566,N_1176,In_1963);
or U1567 (N_1567,In_115,N_978);
and U1568 (N_1568,N_1135,N_1192);
and U1569 (N_1569,N_1045,N_892);
xnor U1570 (N_1570,N_961,N_1035);
and U1571 (N_1571,N_443,N_1008);
and U1572 (N_1572,N_145,In_914);
and U1573 (N_1573,N_966,In_294);
nor U1574 (N_1574,N_340,In_1763);
or U1575 (N_1575,In_1896,N_447);
and U1576 (N_1576,In_159,N_581);
nor U1577 (N_1577,In_887,N_879);
xnor U1578 (N_1578,N_586,N_826);
and U1579 (N_1579,N_1130,In_1816);
xnor U1580 (N_1580,N_1020,N_716);
xnor U1581 (N_1581,N_706,In_1424);
nor U1582 (N_1582,N_1116,In_1831);
nor U1583 (N_1583,In_1545,N_1036);
xnor U1584 (N_1584,N_855,N_937);
and U1585 (N_1585,N_439,N_971);
nor U1586 (N_1586,In_242,N_995);
nand U1587 (N_1587,N_861,N_548);
nor U1588 (N_1588,In_628,N_925);
nand U1589 (N_1589,N_734,N_687);
xor U1590 (N_1590,In_1316,N_1160);
xnor U1591 (N_1591,In_1463,In_496);
nand U1592 (N_1592,N_589,N_547);
and U1593 (N_1593,N_1102,In_1403);
xnor U1594 (N_1594,N_360,N_759);
and U1595 (N_1595,N_1189,N_871);
and U1596 (N_1596,In_1148,N_867);
nor U1597 (N_1597,N_857,N_1065);
nand U1598 (N_1598,N_1178,N_632);
nand U1599 (N_1599,N_1086,N_891);
nor U1600 (N_1600,N_1482,N_1426);
nor U1601 (N_1601,N_1251,N_1278);
or U1602 (N_1602,N_1562,N_1243);
nor U1603 (N_1603,N_1200,N_1487);
nand U1604 (N_1604,N_1543,N_1512);
xor U1605 (N_1605,N_1254,N_1556);
and U1606 (N_1606,N_1463,N_1210);
nand U1607 (N_1607,N_1334,N_1589);
nor U1608 (N_1608,N_1424,N_1320);
nand U1609 (N_1609,N_1502,N_1402);
nor U1610 (N_1610,N_1412,N_1270);
nand U1611 (N_1611,N_1504,N_1245);
nand U1612 (N_1612,N_1235,N_1291);
nand U1613 (N_1613,N_1574,N_1297);
nand U1614 (N_1614,N_1330,N_1230);
or U1615 (N_1615,N_1385,N_1266);
nor U1616 (N_1616,N_1500,N_1212);
nand U1617 (N_1617,N_1339,N_1441);
and U1618 (N_1618,N_1457,N_1473);
nor U1619 (N_1619,N_1501,N_1440);
xor U1620 (N_1620,N_1211,N_1443);
xnor U1621 (N_1621,N_1526,N_1517);
or U1622 (N_1622,N_1591,N_1445);
xor U1623 (N_1623,N_1413,N_1498);
nor U1624 (N_1624,N_1479,N_1223);
nor U1625 (N_1625,N_1311,N_1359);
and U1626 (N_1626,N_1447,N_1575);
and U1627 (N_1627,N_1471,N_1327);
nor U1628 (N_1628,N_1495,N_1579);
and U1629 (N_1629,N_1345,N_1333);
xnor U1630 (N_1630,N_1290,N_1328);
xor U1631 (N_1631,N_1461,N_1303);
nand U1632 (N_1632,N_1419,N_1532);
and U1633 (N_1633,N_1382,N_1496);
nand U1634 (N_1634,N_1294,N_1552);
nand U1635 (N_1635,N_1475,N_1584);
and U1636 (N_1636,N_1257,N_1312);
nor U1637 (N_1637,N_1576,N_1425);
nand U1638 (N_1638,N_1319,N_1452);
nand U1639 (N_1639,N_1233,N_1302);
nor U1640 (N_1640,N_1340,N_1244);
or U1641 (N_1641,N_1313,N_1565);
and U1642 (N_1642,N_1462,N_1283);
and U1643 (N_1643,N_1555,N_1394);
xnor U1644 (N_1644,N_1459,N_1390);
nand U1645 (N_1645,N_1274,N_1338);
nor U1646 (N_1646,N_1468,N_1590);
xnor U1647 (N_1647,N_1314,N_1224);
nand U1648 (N_1648,N_1400,N_1374);
and U1649 (N_1649,N_1371,N_1241);
xnor U1650 (N_1650,N_1505,N_1350);
or U1651 (N_1651,N_1269,N_1342);
nand U1652 (N_1652,N_1455,N_1393);
and U1653 (N_1653,N_1518,N_1523);
nand U1654 (N_1654,N_1375,N_1279);
nor U1655 (N_1655,N_1355,N_1489);
and U1656 (N_1656,N_1396,N_1260);
nand U1657 (N_1657,N_1222,N_1226);
or U1658 (N_1658,N_1386,N_1264);
nor U1659 (N_1659,N_1407,N_1285);
or U1660 (N_1660,N_1369,N_1595);
nand U1661 (N_1661,N_1531,N_1238);
nand U1662 (N_1662,N_1456,N_1218);
or U1663 (N_1663,N_1207,N_1300);
xnor U1664 (N_1664,N_1356,N_1389);
and U1665 (N_1665,N_1492,N_1446);
nand U1666 (N_1666,N_1414,N_1436);
and U1667 (N_1667,N_1520,N_1524);
xor U1668 (N_1668,N_1304,N_1252);
xnor U1669 (N_1669,N_1561,N_1406);
and U1670 (N_1670,N_1451,N_1401);
and U1671 (N_1671,N_1522,N_1227);
nand U1672 (N_1672,N_1321,N_1301);
or U1673 (N_1673,N_1280,N_1553);
and U1674 (N_1674,N_1521,N_1253);
nand U1675 (N_1675,N_1439,N_1405);
or U1676 (N_1676,N_1219,N_1429);
xnor U1677 (N_1677,N_1315,N_1541);
nor U1678 (N_1678,N_1308,N_1485);
nand U1679 (N_1679,N_1564,N_1507);
and U1680 (N_1680,N_1373,N_1282);
nor U1681 (N_1681,N_1599,N_1409);
nor U1682 (N_1682,N_1347,N_1240);
xor U1683 (N_1683,N_1324,N_1594);
nand U1684 (N_1684,N_1381,N_1516);
and U1685 (N_1685,N_1547,N_1488);
nor U1686 (N_1686,N_1542,N_1215);
nor U1687 (N_1687,N_1351,N_1431);
or U1688 (N_1688,N_1464,N_1548);
xnor U1689 (N_1689,N_1474,N_1387);
nand U1690 (N_1690,N_1566,N_1361);
or U1691 (N_1691,N_1284,N_1325);
xnor U1692 (N_1692,N_1399,N_1203);
xnor U1693 (N_1693,N_1341,N_1236);
or U1694 (N_1694,N_1364,N_1550);
nor U1695 (N_1695,N_1318,N_1449);
xor U1696 (N_1696,N_1398,N_1397);
nand U1697 (N_1697,N_1348,N_1506);
nor U1698 (N_1698,N_1322,N_1513);
and U1699 (N_1699,N_1583,N_1209);
and U1700 (N_1700,N_1433,N_1423);
nand U1701 (N_1701,N_1395,N_1261);
and U1702 (N_1702,N_1585,N_1332);
or U1703 (N_1703,N_1293,N_1289);
nand U1704 (N_1704,N_1343,N_1494);
or U1705 (N_1705,N_1571,N_1588);
and U1706 (N_1706,N_1416,N_1206);
or U1707 (N_1707,N_1448,N_1438);
xnor U1708 (N_1708,N_1596,N_1533);
or U1709 (N_1709,N_1410,N_1377);
and U1710 (N_1710,N_1404,N_1204);
xnor U1711 (N_1711,N_1587,N_1480);
and U1712 (N_1712,N_1572,N_1360);
or U1713 (N_1713,N_1379,N_1503);
nor U1714 (N_1714,N_1296,N_1466);
and U1715 (N_1715,N_1370,N_1357);
and U1716 (N_1716,N_1569,N_1242);
and U1717 (N_1717,N_1559,N_1508);
xor U1718 (N_1718,N_1421,N_1353);
and U1719 (N_1719,N_1510,N_1467);
or U1720 (N_1720,N_1263,N_1490);
or U1721 (N_1721,N_1249,N_1267);
nor U1722 (N_1722,N_1392,N_1256);
nand U1723 (N_1723,N_1337,N_1580);
nand U1724 (N_1724,N_1239,N_1335);
nand U1725 (N_1725,N_1536,N_1491);
nor U1726 (N_1726,N_1530,N_1593);
or U1727 (N_1727,N_1586,N_1465);
nor U1728 (N_1728,N_1331,N_1388);
and U1729 (N_1729,N_1205,N_1567);
or U1730 (N_1730,N_1378,N_1273);
xor U1731 (N_1731,N_1213,N_1568);
nand U1732 (N_1732,N_1525,N_1432);
and U1733 (N_1733,N_1344,N_1558);
nand U1734 (N_1734,N_1298,N_1411);
nor U1735 (N_1735,N_1250,N_1234);
and U1736 (N_1736,N_1287,N_1460);
or U1737 (N_1737,N_1202,N_1478);
nor U1738 (N_1738,N_1201,N_1271);
nor U1739 (N_1739,N_1310,N_1534);
xor U1740 (N_1740,N_1231,N_1476);
xor U1741 (N_1741,N_1577,N_1275);
or U1742 (N_1742,N_1499,N_1365);
or U1743 (N_1743,N_1349,N_1560);
nor U1744 (N_1744,N_1539,N_1288);
xnor U1745 (N_1745,N_1391,N_1481);
or U1746 (N_1746,N_1598,N_1597);
or U1747 (N_1747,N_1228,N_1214);
or U1748 (N_1748,N_1537,N_1352);
nor U1749 (N_1749,N_1535,N_1326);
and U1750 (N_1750,N_1376,N_1509);
or U1751 (N_1751,N_1453,N_1422);
nand U1752 (N_1752,N_1362,N_1458);
or U1753 (N_1753,N_1367,N_1268);
xnor U1754 (N_1754,N_1472,N_1220);
xor U1755 (N_1755,N_1363,N_1528);
nand U1756 (N_1756,N_1538,N_1483);
xor U1757 (N_1757,N_1511,N_1497);
and U1758 (N_1758,N_1435,N_1493);
and U1759 (N_1759,N_1277,N_1225);
or U1760 (N_1760,N_1428,N_1372);
nor U1761 (N_1761,N_1557,N_1259);
nand U1762 (N_1762,N_1316,N_1366);
xnor U1763 (N_1763,N_1295,N_1570);
and U1764 (N_1764,N_1551,N_1380);
nor U1765 (N_1765,N_1276,N_1247);
or U1766 (N_1766,N_1217,N_1323);
or U1767 (N_1767,N_1442,N_1384);
and U1768 (N_1768,N_1563,N_1281);
nor U1769 (N_1769,N_1592,N_1346);
and U1770 (N_1770,N_1258,N_1208);
and U1771 (N_1771,N_1368,N_1358);
xnor U1772 (N_1772,N_1237,N_1515);
nand U1773 (N_1773,N_1444,N_1549);
nor U1774 (N_1774,N_1519,N_1248);
nor U1775 (N_1775,N_1292,N_1329);
or U1776 (N_1776,N_1486,N_1354);
nand U1777 (N_1777,N_1484,N_1546);
and U1778 (N_1778,N_1408,N_1427);
nand U1779 (N_1779,N_1299,N_1415);
nand U1780 (N_1780,N_1454,N_1255);
or U1781 (N_1781,N_1434,N_1229);
nand U1782 (N_1782,N_1383,N_1477);
nand U1783 (N_1783,N_1317,N_1529);
xnor U1784 (N_1784,N_1545,N_1232);
xor U1785 (N_1785,N_1430,N_1470);
xnor U1786 (N_1786,N_1221,N_1336);
or U1787 (N_1787,N_1265,N_1540);
nor U1788 (N_1788,N_1403,N_1417);
or U1789 (N_1789,N_1437,N_1578);
nor U1790 (N_1790,N_1418,N_1514);
or U1791 (N_1791,N_1305,N_1307);
and U1792 (N_1792,N_1544,N_1581);
xnor U1793 (N_1793,N_1573,N_1450);
and U1794 (N_1794,N_1554,N_1469);
nor U1795 (N_1795,N_1246,N_1582);
or U1796 (N_1796,N_1262,N_1216);
and U1797 (N_1797,N_1309,N_1306);
xor U1798 (N_1798,N_1420,N_1286);
nor U1799 (N_1799,N_1527,N_1272);
and U1800 (N_1800,N_1225,N_1517);
and U1801 (N_1801,N_1597,N_1422);
nand U1802 (N_1802,N_1534,N_1338);
and U1803 (N_1803,N_1583,N_1555);
xor U1804 (N_1804,N_1204,N_1241);
or U1805 (N_1805,N_1385,N_1540);
or U1806 (N_1806,N_1449,N_1399);
nor U1807 (N_1807,N_1532,N_1393);
or U1808 (N_1808,N_1419,N_1377);
nand U1809 (N_1809,N_1445,N_1336);
nand U1810 (N_1810,N_1333,N_1245);
and U1811 (N_1811,N_1261,N_1512);
and U1812 (N_1812,N_1584,N_1426);
nand U1813 (N_1813,N_1406,N_1221);
and U1814 (N_1814,N_1426,N_1398);
or U1815 (N_1815,N_1277,N_1212);
or U1816 (N_1816,N_1466,N_1573);
xor U1817 (N_1817,N_1499,N_1492);
and U1818 (N_1818,N_1207,N_1577);
or U1819 (N_1819,N_1577,N_1363);
or U1820 (N_1820,N_1576,N_1247);
or U1821 (N_1821,N_1578,N_1454);
or U1822 (N_1822,N_1563,N_1225);
or U1823 (N_1823,N_1443,N_1501);
xor U1824 (N_1824,N_1446,N_1550);
and U1825 (N_1825,N_1586,N_1500);
and U1826 (N_1826,N_1229,N_1220);
nand U1827 (N_1827,N_1203,N_1537);
nand U1828 (N_1828,N_1371,N_1329);
and U1829 (N_1829,N_1375,N_1472);
or U1830 (N_1830,N_1589,N_1450);
nor U1831 (N_1831,N_1448,N_1458);
nand U1832 (N_1832,N_1217,N_1450);
nor U1833 (N_1833,N_1558,N_1277);
xnor U1834 (N_1834,N_1424,N_1387);
or U1835 (N_1835,N_1518,N_1340);
nand U1836 (N_1836,N_1506,N_1243);
nor U1837 (N_1837,N_1283,N_1290);
nand U1838 (N_1838,N_1375,N_1344);
nor U1839 (N_1839,N_1458,N_1409);
nand U1840 (N_1840,N_1354,N_1304);
nor U1841 (N_1841,N_1313,N_1506);
and U1842 (N_1842,N_1535,N_1269);
xor U1843 (N_1843,N_1506,N_1208);
xnor U1844 (N_1844,N_1251,N_1491);
nor U1845 (N_1845,N_1511,N_1461);
nor U1846 (N_1846,N_1232,N_1309);
nor U1847 (N_1847,N_1413,N_1495);
and U1848 (N_1848,N_1374,N_1538);
and U1849 (N_1849,N_1500,N_1304);
nor U1850 (N_1850,N_1213,N_1230);
nand U1851 (N_1851,N_1506,N_1283);
nand U1852 (N_1852,N_1344,N_1355);
and U1853 (N_1853,N_1229,N_1426);
xnor U1854 (N_1854,N_1264,N_1467);
xnor U1855 (N_1855,N_1204,N_1207);
or U1856 (N_1856,N_1566,N_1504);
nor U1857 (N_1857,N_1249,N_1213);
nand U1858 (N_1858,N_1232,N_1224);
xnor U1859 (N_1859,N_1441,N_1355);
nand U1860 (N_1860,N_1271,N_1449);
or U1861 (N_1861,N_1428,N_1509);
and U1862 (N_1862,N_1440,N_1305);
xnor U1863 (N_1863,N_1383,N_1222);
nand U1864 (N_1864,N_1469,N_1274);
or U1865 (N_1865,N_1300,N_1451);
and U1866 (N_1866,N_1430,N_1428);
nand U1867 (N_1867,N_1363,N_1520);
or U1868 (N_1868,N_1273,N_1388);
or U1869 (N_1869,N_1309,N_1334);
or U1870 (N_1870,N_1391,N_1495);
xnor U1871 (N_1871,N_1306,N_1248);
or U1872 (N_1872,N_1346,N_1377);
nand U1873 (N_1873,N_1500,N_1523);
nor U1874 (N_1874,N_1506,N_1533);
xnor U1875 (N_1875,N_1472,N_1285);
or U1876 (N_1876,N_1527,N_1206);
or U1877 (N_1877,N_1583,N_1527);
nor U1878 (N_1878,N_1350,N_1453);
nand U1879 (N_1879,N_1285,N_1449);
and U1880 (N_1880,N_1279,N_1253);
nand U1881 (N_1881,N_1203,N_1452);
or U1882 (N_1882,N_1462,N_1428);
or U1883 (N_1883,N_1305,N_1422);
nor U1884 (N_1884,N_1594,N_1457);
and U1885 (N_1885,N_1519,N_1485);
nand U1886 (N_1886,N_1254,N_1584);
nand U1887 (N_1887,N_1535,N_1214);
xnor U1888 (N_1888,N_1541,N_1429);
and U1889 (N_1889,N_1222,N_1534);
and U1890 (N_1890,N_1230,N_1440);
nor U1891 (N_1891,N_1299,N_1312);
xnor U1892 (N_1892,N_1341,N_1550);
nor U1893 (N_1893,N_1294,N_1511);
nor U1894 (N_1894,N_1403,N_1402);
xor U1895 (N_1895,N_1448,N_1331);
xor U1896 (N_1896,N_1560,N_1449);
nand U1897 (N_1897,N_1475,N_1411);
or U1898 (N_1898,N_1468,N_1250);
and U1899 (N_1899,N_1550,N_1271);
or U1900 (N_1900,N_1541,N_1294);
nand U1901 (N_1901,N_1392,N_1286);
nor U1902 (N_1902,N_1295,N_1542);
xor U1903 (N_1903,N_1585,N_1221);
or U1904 (N_1904,N_1489,N_1239);
or U1905 (N_1905,N_1511,N_1528);
or U1906 (N_1906,N_1539,N_1500);
nor U1907 (N_1907,N_1552,N_1242);
nor U1908 (N_1908,N_1562,N_1511);
nand U1909 (N_1909,N_1456,N_1572);
or U1910 (N_1910,N_1415,N_1468);
nor U1911 (N_1911,N_1222,N_1552);
nand U1912 (N_1912,N_1429,N_1485);
or U1913 (N_1913,N_1481,N_1467);
xnor U1914 (N_1914,N_1560,N_1363);
xor U1915 (N_1915,N_1419,N_1551);
nor U1916 (N_1916,N_1281,N_1438);
nand U1917 (N_1917,N_1500,N_1295);
nand U1918 (N_1918,N_1346,N_1279);
and U1919 (N_1919,N_1590,N_1239);
xnor U1920 (N_1920,N_1324,N_1256);
and U1921 (N_1921,N_1457,N_1282);
or U1922 (N_1922,N_1592,N_1520);
and U1923 (N_1923,N_1322,N_1591);
and U1924 (N_1924,N_1466,N_1379);
nor U1925 (N_1925,N_1332,N_1317);
xnor U1926 (N_1926,N_1329,N_1342);
xnor U1927 (N_1927,N_1315,N_1514);
xor U1928 (N_1928,N_1583,N_1420);
nor U1929 (N_1929,N_1316,N_1433);
nor U1930 (N_1930,N_1596,N_1327);
nor U1931 (N_1931,N_1588,N_1309);
nand U1932 (N_1932,N_1380,N_1305);
nor U1933 (N_1933,N_1540,N_1472);
and U1934 (N_1934,N_1443,N_1450);
nor U1935 (N_1935,N_1361,N_1352);
and U1936 (N_1936,N_1449,N_1537);
and U1937 (N_1937,N_1278,N_1211);
or U1938 (N_1938,N_1552,N_1541);
nor U1939 (N_1939,N_1488,N_1361);
nand U1940 (N_1940,N_1581,N_1579);
nor U1941 (N_1941,N_1358,N_1281);
or U1942 (N_1942,N_1217,N_1497);
nand U1943 (N_1943,N_1437,N_1548);
nor U1944 (N_1944,N_1342,N_1229);
and U1945 (N_1945,N_1496,N_1300);
and U1946 (N_1946,N_1282,N_1594);
nor U1947 (N_1947,N_1261,N_1420);
or U1948 (N_1948,N_1379,N_1506);
nand U1949 (N_1949,N_1373,N_1236);
xor U1950 (N_1950,N_1434,N_1212);
xor U1951 (N_1951,N_1502,N_1507);
nand U1952 (N_1952,N_1308,N_1427);
nand U1953 (N_1953,N_1421,N_1306);
nor U1954 (N_1954,N_1204,N_1264);
or U1955 (N_1955,N_1334,N_1580);
or U1956 (N_1956,N_1457,N_1428);
and U1957 (N_1957,N_1286,N_1276);
nor U1958 (N_1958,N_1418,N_1538);
or U1959 (N_1959,N_1382,N_1465);
nand U1960 (N_1960,N_1237,N_1512);
nand U1961 (N_1961,N_1550,N_1290);
and U1962 (N_1962,N_1291,N_1395);
nor U1963 (N_1963,N_1588,N_1590);
xnor U1964 (N_1964,N_1511,N_1407);
and U1965 (N_1965,N_1220,N_1233);
nor U1966 (N_1966,N_1254,N_1316);
or U1967 (N_1967,N_1480,N_1238);
nand U1968 (N_1968,N_1418,N_1426);
and U1969 (N_1969,N_1292,N_1267);
or U1970 (N_1970,N_1345,N_1377);
or U1971 (N_1971,N_1280,N_1586);
and U1972 (N_1972,N_1468,N_1376);
nand U1973 (N_1973,N_1474,N_1519);
and U1974 (N_1974,N_1398,N_1335);
xor U1975 (N_1975,N_1396,N_1405);
nor U1976 (N_1976,N_1525,N_1585);
nor U1977 (N_1977,N_1556,N_1256);
nand U1978 (N_1978,N_1513,N_1482);
and U1979 (N_1979,N_1514,N_1548);
nor U1980 (N_1980,N_1258,N_1523);
xnor U1981 (N_1981,N_1525,N_1346);
nor U1982 (N_1982,N_1318,N_1515);
and U1983 (N_1983,N_1427,N_1227);
or U1984 (N_1984,N_1440,N_1219);
nor U1985 (N_1985,N_1414,N_1220);
and U1986 (N_1986,N_1315,N_1416);
and U1987 (N_1987,N_1439,N_1408);
and U1988 (N_1988,N_1535,N_1268);
or U1989 (N_1989,N_1521,N_1336);
xnor U1990 (N_1990,N_1295,N_1381);
xor U1991 (N_1991,N_1234,N_1583);
and U1992 (N_1992,N_1544,N_1259);
xor U1993 (N_1993,N_1346,N_1529);
nand U1994 (N_1994,N_1440,N_1484);
nand U1995 (N_1995,N_1405,N_1530);
and U1996 (N_1996,N_1566,N_1404);
xor U1997 (N_1997,N_1595,N_1428);
nand U1998 (N_1998,N_1492,N_1381);
and U1999 (N_1999,N_1419,N_1412);
nor U2000 (N_2000,N_1621,N_1733);
and U2001 (N_2001,N_1662,N_1893);
nor U2002 (N_2002,N_1661,N_1628);
nor U2003 (N_2003,N_1625,N_1776);
nor U2004 (N_2004,N_1610,N_1999);
nand U2005 (N_2005,N_1886,N_1858);
nor U2006 (N_2006,N_1618,N_1943);
and U2007 (N_2007,N_1729,N_1942);
xnor U2008 (N_2008,N_1809,N_1951);
nand U2009 (N_2009,N_1745,N_1826);
or U2010 (N_2010,N_1975,N_1716);
nor U2011 (N_2011,N_1813,N_1705);
nor U2012 (N_2012,N_1856,N_1931);
or U2013 (N_2013,N_1614,N_1602);
nor U2014 (N_2014,N_1750,N_1773);
xor U2015 (N_2015,N_1781,N_1731);
nor U2016 (N_2016,N_1883,N_1816);
and U2017 (N_2017,N_1712,N_1935);
nor U2018 (N_2018,N_1861,N_1607);
nor U2019 (N_2019,N_1890,N_1604);
xor U2020 (N_2020,N_1896,N_1822);
and U2021 (N_2021,N_1980,N_1634);
xnor U2022 (N_2022,N_1792,N_1910);
nor U2023 (N_2023,N_1635,N_1644);
nor U2024 (N_2024,N_1944,N_1879);
and U2025 (N_2025,N_1674,N_1791);
nor U2026 (N_2026,N_1752,N_1629);
or U2027 (N_2027,N_1912,N_1667);
and U2028 (N_2028,N_1904,N_1627);
or U2029 (N_2029,N_1663,N_1666);
xor U2030 (N_2030,N_1640,N_1723);
xor U2031 (N_2031,N_1703,N_1693);
and U2032 (N_2032,N_1742,N_1649);
or U2033 (N_2033,N_1988,N_1677);
nand U2034 (N_2034,N_1829,N_1786);
or U2035 (N_2035,N_1965,N_1766);
xnor U2036 (N_2036,N_1905,N_1623);
xor U2037 (N_2037,N_1916,N_1737);
or U2038 (N_2038,N_1979,N_1795);
nor U2039 (N_2039,N_1815,N_1747);
xor U2040 (N_2040,N_1682,N_1653);
and U2041 (N_2041,N_1877,N_1976);
nor U2042 (N_2042,N_1963,N_1798);
and U2043 (N_2043,N_1933,N_1639);
or U2044 (N_2044,N_1958,N_1801);
and U2045 (N_2045,N_1721,N_1811);
and U2046 (N_2046,N_1664,N_1962);
nand U2047 (N_2047,N_1995,N_1728);
or U2048 (N_2048,N_1803,N_1997);
nor U2049 (N_2049,N_1631,N_1757);
nand U2050 (N_2050,N_1929,N_1880);
nor U2051 (N_2051,N_1679,N_1884);
nor U2052 (N_2052,N_1642,N_1970);
xor U2053 (N_2053,N_1857,N_1819);
or U2054 (N_2054,N_1800,N_1651);
xor U2055 (N_2055,N_1977,N_1724);
or U2056 (N_2056,N_1866,N_1814);
xor U2057 (N_2057,N_1796,N_1768);
and U2058 (N_2058,N_1810,N_1847);
nor U2059 (N_2059,N_1804,N_1684);
nand U2060 (N_2060,N_1761,N_1996);
and U2061 (N_2061,N_1897,N_1966);
nor U2062 (N_2062,N_1947,N_1820);
xor U2063 (N_2063,N_1992,N_1864);
nor U2064 (N_2064,N_1670,N_1899);
xnor U2065 (N_2065,N_1840,N_1885);
nand U2066 (N_2066,N_1732,N_1675);
and U2067 (N_2067,N_1983,N_1685);
and U2068 (N_2068,N_1941,N_1688);
or U2069 (N_2069,N_1952,N_1789);
and U2070 (N_2070,N_1710,N_1936);
nand U2071 (N_2071,N_1828,N_1671);
nor U2072 (N_2072,N_1709,N_1928);
nand U2073 (N_2073,N_1605,N_1609);
or U2074 (N_2074,N_1878,N_1770);
or U2075 (N_2075,N_1741,N_1799);
and U2076 (N_2076,N_1669,N_1696);
and U2077 (N_2077,N_1626,N_1774);
or U2078 (N_2078,N_1844,N_1643);
nor U2079 (N_2079,N_1895,N_1706);
nand U2080 (N_2080,N_1746,N_1969);
nor U2081 (N_2081,N_1730,N_1638);
and U2082 (N_2082,N_1735,N_1889);
xor U2083 (N_2083,N_1915,N_1823);
xor U2084 (N_2084,N_1641,N_1964);
nand U2085 (N_2085,N_1700,N_1989);
xnor U2086 (N_2086,N_1867,N_1914);
xnor U2087 (N_2087,N_1802,N_1824);
nor U2088 (N_2088,N_1923,N_1955);
nor U2089 (N_2089,N_1849,N_1901);
nand U2090 (N_2090,N_1753,N_1727);
nand U2091 (N_2091,N_1722,N_1718);
nand U2092 (N_2092,N_1658,N_1739);
or U2093 (N_2093,N_1787,N_1848);
xnor U2094 (N_2094,N_1917,N_1755);
and U2095 (N_2095,N_1632,N_1973);
nor U2096 (N_2096,N_1659,N_1719);
xnor U2097 (N_2097,N_1600,N_1873);
and U2098 (N_2098,N_1772,N_1833);
nand U2099 (N_2099,N_1763,N_1838);
or U2100 (N_2100,N_1926,N_1784);
and U2101 (N_2101,N_1665,N_1839);
nand U2102 (N_2102,N_1817,N_1689);
xor U2103 (N_2103,N_1646,N_1940);
nand U2104 (N_2104,N_1862,N_1900);
or U2105 (N_2105,N_1633,N_1603);
nor U2106 (N_2106,N_1701,N_1919);
nand U2107 (N_2107,N_1749,N_1938);
nand U2108 (N_2108,N_1779,N_1624);
or U2109 (N_2109,N_1793,N_1998);
nor U2110 (N_2110,N_1756,N_1985);
nand U2111 (N_2111,N_1612,N_1853);
or U2112 (N_2112,N_1948,N_1961);
nor U2113 (N_2113,N_1830,N_1863);
nand U2114 (N_2114,N_1949,N_1702);
and U2115 (N_2115,N_1695,N_1692);
xor U2116 (N_2116,N_1790,N_1754);
nor U2117 (N_2117,N_1835,N_1846);
or U2118 (N_2118,N_1836,N_1778);
or U2119 (N_2119,N_1868,N_1842);
nor U2120 (N_2120,N_1854,N_1777);
or U2121 (N_2121,N_1619,N_1767);
xnor U2122 (N_2122,N_1882,N_1699);
nand U2123 (N_2123,N_1921,N_1738);
nor U2124 (N_2124,N_1805,N_1872);
or U2125 (N_2125,N_1950,N_1694);
xnor U2126 (N_2126,N_1762,N_1908);
or U2127 (N_2127,N_1825,N_1852);
and U2128 (N_2128,N_1974,N_1794);
and U2129 (N_2129,N_1870,N_1622);
nor U2130 (N_2130,N_1888,N_1945);
or U2131 (N_2131,N_1707,N_1668);
nand U2132 (N_2132,N_1650,N_1617);
or U2133 (N_2133,N_1691,N_1812);
and U2134 (N_2134,N_1930,N_1764);
nand U2135 (N_2135,N_1611,N_1991);
or U2136 (N_2136,N_1608,N_1759);
or U2137 (N_2137,N_1990,N_1720);
or U2138 (N_2138,N_1673,N_1655);
xnor U2139 (N_2139,N_1657,N_1647);
xor U2140 (N_2140,N_1704,N_1913);
xnor U2141 (N_2141,N_1874,N_1807);
nand U2142 (N_2142,N_1937,N_1953);
nor U2143 (N_2143,N_1859,N_1881);
xor U2144 (N_2144,N_1887,N_1934);
nand U2145 (N_2145,N_1954,N_1855);
xnor U2146 (N_2146,N_1765,N_1939);
nand U2147 (N_2147,N_1907,N_1808);
xnor U2148 (N_2148,N_1920,N_1606);
and U2149 (N_2149,N_1748,N_1686);
xnor U2150 (N_2150,N_1831,N_1771);
xor U2151 (N_2151,N_1932,N_1827);
nor U2152 (N_2152,N_1711,N_1637);
and U2153 (N_2153,N_1850,N_1994);
nand U2154 (N_2154,N_1615,N_1865);
xor U2155 (N_2155,N_1783,N_1656);
or U2156 (N_2156,N_1832,N_1845);
xor U2157 (N_2157,N_1697,N_1968);
nand U2158 (N_2158,N_1751,N_1946);
and U2159 (N_2159,N_1906,N_1717);
and U2160 (N_2160,N_1760,N_1978);
xor U2161 (N_2161,N_1841,N_1834);
or U2162 (N_2162,N_1672,N_1981);
or U2163 (N_2163,N_1843,N_1797);
or U2164 (N_2164,N_1708,N_1894);
nor U2165 (N_2165,N_1681,N_1818);
nand U2166 (N_2166,N_1680,N_1869);
xnor U2167 (N_2167,N_1630,N_1924);
nand U2168 (N_2168,N_1744,N_1971);
xnor U2169 (N_2169,N_1715,N_1986);
or U2170 (N_2170,N_1726,N_1851);
nor U2171 (N_2171,N_1875,N_1927);
nor U2172 (N_2172,N_1909,N_1725);
xor U2173 (N_2173,N_1648,N_1959);
nor U2174 (N_2174,N_1758,N_1660);
nor U2175 (N_2175,N_1743,N_1736);
nand U2176 (N_2176,N_1860,N_1698);
nand U2177 (N_2177,N_1982,N_1734);
or U2178 (N_2178,N_1984,N_1782);
xor U2179 (N_2179,N_1876,N_1902);
and U2180 (N_2180,N_1690,N_1918);
xnor U2181 (N_2181,N_1601,N_1620);
or U2182 (N_2182,N_1806,N_1613);
xnor U2183 (N_2183,N_1780,N_1922);
xor U2184 (N_2184,N_1714,N_1616);
or U2185 (N_2185,N_1960,N_1871);
xor U2186 (N_2186,N_1957,N_1676);
xnor U2187 (N_2187,N_1821,N_1713);
nand U2188 (N_2188,N_1652,N_1967);
or U2189 (N_2189,N_1769,N_1925);
or U2190 (N_2190,N_1956,N_1788);
nand U2191 (N_2191,N_1636,N_1740);
nor U2192 (N_2192,N_1892,N_1683);
or U2193 (N_2193,N_1678,N_1903);
xor U2194 (N_2194,N_1911,N_1837);
or U2195 (N_2195,N_1687,N_1993);
nand U2196 (N_2196,N_1987,N_1775);
xnor U2197 (N_2197,N_1972,N_1785);
nand U2198 (N_2198,N_1654,N_1645);
nand U2199 (N_2199,N_1891,N_1898);
nand U2200 (N_2200,N_1607,N_1688);
xor U2201 (N_2201,N_1803,N_1823);
nor U2202 (N_2202,N_1708,N_1858);
nand U2203 (N_2203,N_1727,N_1851);
nand U2204 (N_2204,N_1727,N_1931);
xor U2205 (N_2205,N_1914,N_1992);
xnor U2206 (N_2206,N_1750,N_1847);
or U2207 (N_2207,N_1816,N_1774);
xor U2208 (N_2208,N_1706,N_1732);
nor U2209 (N_2209,N_1835,N_1775);
and U2210 (N_2210,N_1642,N_1854);
nand U2211 (N_2211,N_1759,N_1893);
xnor U2212 (N_2212,N_1761,N_1822);
and U2213 (N_2213,N_1715,N_1859);
or U2214 (N_2214,N_1753,N_1964);
nand U2215 (N_2215,N_1668,N_1738);
or U2216 (N_2216,N_1604,N_1968);
nand U2217 (N_2217,N_1981,N_1866);
or U2218 (N_2218,N_1803,N_1696);
and U2219 (N_2219,N_1871,N_1693);
nand U2220 (N_2220,N_1738,N_1836);
and U2221 (N_2221,N_1701,N_1757);
xnor U2222 (N_2222,N_1607,N_1810);
nor U2223 (N_2223,N_1637,N_1854);
nor U2224 (N_2224,N_1608,N_1816);
xor U2225 (N_2225,N_1989,N_1693);
xor U2226 (N_2226,N_1996,N_1923);
xnor U2227 (N_2227,N_1637,N_1773);
and U2228 (N_2228,N_1816,N_1805);
xor U2229 (N_2229,N_1653,N_1988);
nand U2230 (N_2230,N_1876,N_1930);
and U2231 (N_2231,N_1869,N_1831);
and U2232 (N_2232,N_1810,N_1603);
or U2233 (N_2233,N_1739,N_1614);
or U2234 (N_2234,N_1610,N_1815);
xnor U2235 (N_2235,N_1811,N_1891);
nand U2236 (N_2236,N_1891,N_1636);
nand U2237 (N_2237,N_1907,N_1697);
nand U2238 (N_2238,N_1995,N_1752);
or U2239 (N_2239,N_1694,N_1615);
nor U2240 (N_2240,N_1839,N_1973);
nor U2241 (N_2241,N_1856,N_1916);
xor U2242 (N_2242,N_1857,N_1942);
nor U2243 (N_2243,N_1730,N_1874);
xnor U2244 (N_2244,N_1956,N_1792);
nand U2245 (N_2245,N_1862,N_1870);
nand U2246 (N_2246,N_1792,N_1888);
xnor U2247 (N_2247,N_1888,N_1929);
or U2248 (N_2248,N_1868,N_1736);
xor U2249 (N_2249,N_1646,N_1655);
nand U2250 (N_2250,N_1914,N_1882);
and U2251 (N_2251,N_1968,N_1949);
nor U2252 (N_2252,N_1823,N_1916);
xor U2253 (N_2253,N_1877,N_1959);
and U2254 (N_2254,N_1749,N_1912);
and U2255 (N_2255,N_1850,N_1790);
xnor U2256 (N_2256,N_1964,N_1663);
xor U2257 (N_2257,N_1749,N_1705);
or U2258 (N_2258,N_1660,N_1685);
and U2259 (N_2259,N_1819,N_1936);
xnor U2260 (N_2260,N_1832,N_1910);
or U2261 (N_2261,N_1813,N_1803);
nor U2262 (N_2262,N_1880,N_1736);
and U2263 (N_2263,N_1990,N_1684);
nand U2264 (N_2264,N_1850,N_1630);
nor U2265 (N_2265,N_1685,N_1837);
and U2266 (N_2266,N_1883,N_1976);
and U2267 (N_2267,N_1883,N_1660);
and U2268 (N_2268,N_1713,N_1745);
xor U2269 (N_2269,N_1804,N_1624);
or U2270 (N_2270,N_1913,N_1888);
nand U2271 (N_2271,N_1601,N_1606);
nor U2272 (N_2272,N_1678,N_1890);
nand U2273 (N_2273,N_1831,N_1820);
and U2274 (N_2274,N_1995,N_1644);
xor U2275 (N_2275,N_1788,N_1666);
nand U2276 (N_2276,N_1830,N_1741);
or U2277 (N_2277,N_1795,N_1914);
nor U2278 (N_2278,N_1730,N_1666);
xnor U2279 (N_2279,N_1759,N_1703);
xnor U2280 (N_2280,N_1722,N_1767);
nor U2281 (N_2281,N_1648,N_1844);
nand U2282 (N_2282,N_1827,N_1631);
or U2283 (N_2283,N_1893,N_1616);
or U2284 (N_2284,N_1855,N_1969);
and U2285 (N_2285,N_1701,N_1846);
xor U2286 (N_2286,N_1965,N_1897);
or U2287 (N_2287,N_1646,N_1913);
and U2288 (N_2288,N_1798,N_1993);
nor U2289 (N_2289,N_1852,N_1908);
nand U2290 (N_2290,N_1894,N_1823);
xnor U2291 (N_2291,N_1608,N_1983);
and U2292 (N_2292,N_1601,N_1729);
nor U2293 (N_2293,N_1616,N_1677);
nor U2294 (N_2294,N_1872,N_1926);
nand U2295 (N_2295,N_1908,N_1628);
nor U2296 (N_2296,N_1616,N_1866);
or U2297 (N_2297,N_1800,N_1819);
and U2298 (N_2298,N_1712,N_1907);
xnor U2299 (N_2299,N_1755,N_1615);
nor U2300 (N_2300,N_1967,N_1969);
nor U2301 (N_2301,N_1897,N_1619);
nor U2302 (N_2302,N_1733,N_1851);
nand U2303 (N_2303,N_1630,N_1613);
nor U2304 (N_2304,N_1759,N_1932);
and U2305 (N_2305,N_1606,N_1954);
xor U2306 (N_2306,N_1714,N_1813);
xor U2307 (N_2307,N_1684,N_1677);
nor U2308 (N_2308,N_1689,N_1871);
nor U2309 (N_2309,N_1719,N_1984);
and U2310 (N_2310,N_1836,N_1931);
nor U2311 (N_2311,N_1899,N_1753);
or U2312 (N_2312,N_1864,N_1997);
xnor U2313 (N_2313,N_1929,N_1937);
xnor U2314 (N_2314,N_1778,N_1858);
and U2315 (N_2315,N_1994,N_1663);
or U2316 (N_2316,N_1968,N_1642);
or U2317 (N_2317,N_1885,N_1685);
nand U2318 (N_2318,N_1928,N_1946);
or U2319 (N_2319,N_1603,N_1638);
nor U2320 (N_2320,N_1700,N_1923);
nand U2321 (N_2321,N_1735,N_1782);
or U2322 (N_2322,N_1624,N_1603);
nand U2323 (N_2323,N_1654,N_1731);
or U2324 (N_2324,N_1784,N_1980);
nand U2325 (N_2325,N_1687,N_1866);
nor U2326 (N_2326,N_1914,N_1830);
nand U2327 (N_2327,N_1864,N_1637);
xor U2328 (N_2328,N_1987,N_1812);
and U2329 (N_2329,N_1753,N_1747);
or U2330 (N_2330,N_1795,N_1830);
xnor U2331 (N_2331,N_1665,N_1725);
nand U2332 (N_2332,N_1771,N_1850);
nor U2333 (N_2333,N_1671,N_1872);
xnor U2334 (N_2334,N_1968,N_1998);
and U2335 (N_2335,N_1785,N_1830);
or U2336 (N_2336,N_1834,N_1801);
and U2337 (N_2337,N_1664,N_1683);
nor U2338 (N_2338,N_1869,N_1833);
nand U2339 (N_2339,N_1841,N_1990);
or U2340 (N_2340,N_1826,N_1689);
xnor U2341 (N_2341,N_1868,N_1660);
nand U2342 (N_2342,N_1638,N_1677);
and U2343 (N_2343,N_1906,N_1766);
and U2344 (N_2344,N_1804,N_1828);
nand U2345 (N_2345,N_1703,N_1620);
nand U2346 (N_2346,N_1643,N_1702);
xnor U2347 (N_2347,N_1967,N_1860);
and U2348 (N_2348,N_1645,N_1894);
or U2349 (N_2349,N_1913,N_1785);
xnor U2350 (N_2350,N_1845,N_1939);
or U2351 (N_2351,N_1962,N_1794);
or U2352 (N_2352,N_1714,N_1945);
or U2353 (N_2353,N_1907,N_1973);
and U2354 (N_2354,N_1872,N_1611);
or U2355 (N_2355,N_1856,N_1668);
xor U2356 (N_2356,N_1773,N_1725);
nor U2357 (N_2357,N_1849,N_1600);
xnor U2358 (N_2358,N_1909,N_1829);
nor U2359 (N_2359,N_1703,N_1799);
xor U2360 (N_2360,N_1811,N_1675);
nand U2361 (N_2361,N_1659,N_1933);
nor U2362 (N_2362,N_1931,N_1973);
and U2363 (N_2363,N_1754,N_1851);
xnor U2364 (N_2364,N_1669,N_1838);
nand U2365 (N_2365,N_1604,N_1714);
and U2366 (N_2366,N_1664,N_1770);
nor U2367 (N_2367,N_1893,N_1645);
or U2368 (N_2368,N_1777,N_1661);
xor U2369 (N_2369,N_1613,N_1820);
nor U2370 (N_2370,N_1999,N_1910);
nor U2371 (N_2371,N_1847,N_1720);
nor U2372 (N_2372,N_1861,N_1604);
or U2373 (N_2373,N_1943,N_1834);
xnor U2374 (N_2374,N_1761,N_1613);
or U2375 (N_2375,N_1763,N_1978);
or U2376 (N_2376,N_1965,N_1709);
or U2377 (N_2377,N_1782,N_1917);
nand U2378 (N_2378,N_1629,N_1807);
nor U2379 (N_2379,N_1989,N_1985);
nor U2380 (N_2380,N_1659,N_1869);
or U2381 (N_2381,N_1883,N_1979);
or U2382 (N_2382,N_1936,N_1780);
and U2383 (N_2383,N_1651,N_1950);
and U2384 (N_2384,N_1957,N_1805);
or U2385 (N_2385,N_1806,N_1997);
nor U2386 (N_2386,N_1944,N_1765);
nor U2387 (N_2387,N_1655,N_1789);
and U2388 (N_2388,N_1623,N_1657);
nor U2389 (N_2389,N_1792,N_1946);
and U2390 (N_2390,N_1976,N_1677);
nor U2391 (N_2391,N_1606,N_1979);
xor U2392 (N_2392,N_1957,N_1800);
xor U2393 (N_2393,N_1994,N_1703);
nor U2394 (N_2394,N_1782,N_1936);
nor U2395 (N_2395,N_1901,N_1949);
nand U2396 (N_2396,N_1840,N_1831);
and U2397 (N_2397,N_1674,N_1695);
xnor U2398 (N_2398,N_1792,N_1879);
nand U2399 (N_2399,N_1822,N_1644);
and U2400 (N_2400,N_2109,N_2379);
xor U2401 (N_2401,N_2008,N_2191);
nand U2402 (N_2402,N_2090,N_2286);
nor U2403 (N_2403,N_2304,N_2295);
xnor U2404 (N_2404,N_2234,N_2240);
or U2405 (N_2405,N_2071,N_2118);
xnor U2406 (N_2406,N_2168,N_2365);
xor U2407 (N_2407,N_2194,N_2265);
xor U2408 (N_2408,N_2085,N_2394);
xnor U2409 (N_2409,N_2092,N_2017);
nand U2410 (N_2410,N_2341,N_2167);
nor U2411 (N_2411,N_2364,N_2031);
or U2412 (N_2412,N_2370,N_2289);
xnor U2413 (N_2413,N_2115,N_2223);
and U2414 (N_2414,N_2059,N_2318);
nand U2415 (N_2415,N_2236,N_2328);
and U2416 (N_2416,N_2121,N_2345);
xnor U2417 (N_2417,N_2035,N_2013);
nor U2418 (N_2418,N_2188,N_2074);
nor U2419 (N_2419,N_2348,N_2228);
and U2420 (N_2420,N_2352,N_2076);
or U2421 (N_2421,N_2334,N_2395);
nor U2422 (N_2422,N_2303,N_2149);
nand U2423 (N_2423,N_2276,N_2201);
nand U2424 (N_2424,N_2256,N_2219);
nand U2425 (N_2425,N_2269,N_2292);
and U2426 (N_2426,N_2246,N_2218);
nor U2427 (N_2427,N_2263,N_2018);
xor U2428 (N_2428,N_2380,N_2091);
nand U2429 (N_2429,N_2162,N_2270);
or U2430 (N_2430,N_2125,N_2313);
xnor U2431 (N_2431,N_2081,N_2012);
nor U2432 (N_2432,N_2349,N_2332);
nor U2433 (N_2433,N_2038,N_2355);
nand U2434 (N_2434,N_2089,N_2338);
or U2435 (N_2435,N_2183,N_2116);
xnor U2436 (N_2436,N_2032,N_2268);
xor U2437 (N_2437,N_2039,N_2309);
and U2438 (N_2438,N_2014,N_2235);
xnor U2439 (N_2439,N_2046,N_2232);
xor U2440 (N_2440,N_2158,N_2202);
nand U2441 (N_2441,N_2363,N_2330);
and U2442 (N_2442,N_2140,N_2101);
nand U2443 (N_2443,N_2399,N_2026);
xor U2444 (N_2444,N_2137,N_2391);
nor U2445 (N_2445,N_2048,N_2061);
or U2446 (N_2446,N_2004,N_2015);
and U2447 (N_2447,N_2385,N_2175);
and U2448 (N_2448,N_2337,N_2245);
and U2449 (N_2449,N_2357,N_2233);
and U2450 (N_2450,N_2192,N_2378);
xnor U2451 (N_2451,N_2339,N_2130);
xnor U2452 (N_2452,N_2144,N_2011);
and U2453 (N_2453,N_2152,N_2300);
or U2454 (N_2454,N_2311,N_2104);
xor U2455 (N_2455,N_2325,N_2347);
and U2456 (N_2456,N_2077,N_2197);
and U2457 (N_2457,N_2221,N_2249);
nor U2458 (N_2458,N_2283,N_2056);
or U2459 (N_2459,N_2151,N_2088);
or U2460 (N_2460,N_2262,N_2065);
and U2461 (N_2461,N_2293,N_2244);
xor U2462 (N_2462,N_2258,N_2281);
and U2463 (N_2463,N_2041,N_2000);
nand U2464 (N_2464,N_2297,N_2377);
xnor U2465 (N_2465,N_2095,N_2242);
or U2466 (N_2466,N_2350,N_2374);
xor U2467 (N_2467,N_2062,N_2143);
xnor U2468 (N_2468,N_2139,N_2078);
xor U2469 (N_2469,N_2390,N_2287);
nor U2470 (N_2470,N_2133,N_2306);
xor U2471 (N_2471,N_2190,N_2354);
nor U2472 (N_2472,N_2098,N_2299);
or U2473 (N_2473,N_2171,N_2146);
nand U2474 (N_2474,N_2068,N_2315);
xor U2475 (N_2475,N_2069,N_2119);
or U2476 (N_2476,N_2070,N_2393);
or U2477 (N_2477,N_2298,N_2264);
xor U2478 (N_2478,N_2073,N_2226);
and U2479 (N_2479,N_2185,N_2372);
xnor U2480 (N_2480,N_2215,N_2282);
or U2481 (N_2481,N_2361,N_2216);
or U2482 (N_2482,N_2055,N_2134);
or U2483 (N_2483,N_2271,N_2141);
xor U2484 (N_2484,N_2001,N_2003);
nand U2485 (N_2485,N_2358,N_2019);
or U2486 (N_2486,N_2214,N_2285);
or U2487 (N_2487,N_2186,N_2237);
nand U2488 (N_2488,N_2169,N_2179);
and U2489 (N_2489,N_2272,N_2248);
xnor U2490 (N_2490,N_2336,N_2033);
or U2491 (N_2491,N_2037,N_2198);
nand U2492 (N_2492,N_2398,N_2381);
xor U2493 (N_2493,N_2180,N_2154);
or U2494 (N_2494,N_2320,N_2047);
nor U2495 (N_2495,N_2054,N_2253);
nor U2496 (N_2496,N_2093,N_2166);
nor U2497 (N_2497,N_2369,N_2126);
or U2498 (N_2498,N_2213,N_2099);
nand U2499 (N_2499,N_2057,N_2072);
or U2500 (N_2500,N_2131,N_2049);
and U2501 (N_2501,N_2207,N_2386);
xnor U2502 (N_2502,N_2002,N_2206);
nand U2503 (N_2503,N_2110,N_2294);
and U2504 (N_2504,N_2225,N_2324);
nand U2505 (N_2505,N_2020,N_2028);
nor U2506 (N_2506,N_2148,N_2029);
nand U2507 (N_2507,N_2335,N_2117);
nor U2508 (N_2508,N_2060,N_2333);
nand U2509 (N_2509,N_2243,N_2080);
nand U2510 (N_2510,N_2096,N_2396);
nor U2511 (N_2511,N_2209,N_2160);
or U2512 (N_2512,N_2387,N_2051);
xor U2513 (N_2513,N_2023,N_2277);
xnor U2514 (N_2514,N_2239,N_2120);
xnor U2515 (N_2515,N_2195,N_2040);
or U2516 (N_2516,N_2138,N_2174);
nor U2517 (N_2517,N_2319,N_2321);
or U2518 (N_2518,N_2327,N_2302);
nor U2519 (N_2519,N_2107,N_2278);
nor U2520 (N_2520,N_2288,N_2368);
xnor U2521 (N_2521,N_2156,N_2108);
and U2522 (N_2522,N_2097,N_2280);
and U2523 (N_2523,N_2301,N_2044);
xnor U2524 (N_2524,N_2178,N_2208);
and U2525 (N_2525,N_2229,N_2273);
xor U2526 (N_2526,N_2124,N_2042);
and U2527 (N_2527,N_2022,N_2052);
xnor U2528 (N_2528,N_2314,N_2067);
and U2529 (N_2529,N_2312,N_2153);
or U2530 (N_2530,N_2009,N_2200);
and U2531 (N_2531,N_2142,N_2389);
nor U2532 (N_2532,N_2360,N_2388);
or U2533 (N_2533,N_2122,N_2006);
nand U2534 (N_2534,N_2105,N_2103);
nor U2535 (N_2535,N_2163,N_2100);
and U2536 (N_2536,N_2058,N_2317);
xnor U2537 (N_2537,N_2176,N_2005);
nor U2538 (N_2538,N_2255,N_2045);
nor U2539 (N_2539,N_2343,N_2084);
nand U2540 (N_2540,N_2172,N_2181);
nor U2541 (N_2541,N_2279,N_2284);
xnor U2542 (N_2542,N_2331,N_2274);
nor U2543 (N_2543,N_2063,N_2086);
and U2544 (N_2544,N_2083,N_2193);
nor U2545 (N_2545,N_2127,N_2367);
nand U2546 (N_2546,N_2254,N_2113);
xnor U2547 (N_2547,N_2356,N_2066);
nand U2548 (N_2548,N_2159,N_2353);
nor U2549 (N_2549,N_2267,N_2212);
and U2550 (N_2550,N_2308,N_2373);
nor U2551 (N_2551,N_2307,N_2132);
or U2552 (N_2552,N_2205,N_2251);
or U2553 (N_2553,N_2227,N_2261);
or U2554 (N_2554,N_2164,N_2027);
nand U2555 (N_2555,N_2376,N_2170);
xnor U2556 (N_2556,N_2220,N_2034);
xor U2557 (N_2557,N_2275,N_2252);
nand U2558 (N_2558,N_2161,N_2257);
xnor U2559 (N_2559,N_2383,N_2135);
or U2560 (N_2560,N_2177,N_2259);
nor U2561 (N_2561,N_2310,N_2145);
nor U2562 (N_2562,N_2375,N_2344);
nor U2563 (N_2563,N_2136,N_2222);
nand U2564 (N_2564,N_2021,N_2323);
nor U2565 (N_2565,N_2250,N_2203);
nor U2566 (N_2566,N_2329,N_2184);
and U2567 (N_2567,N_2025,N_2224);
or U2568 (N_2568,N_2316,N_2094);
and U2569 (N_2569,N_2087,N_2291);
and U2570 (N_2570,N_2231,N_2112);
nand U2571 (N_2571,N_2359,N_2016);
xnor U2572 (N_2572,N_2114,N_2157);
nand U2573 (N_2573,N_2173,N_2296);
nor U2574 (N_2574,N_2128,N_2340);
and U2575 (N_2575,N_2305,N_2007);
nor U2576 (N_2576,N_2147,N_2150);
and U2577 (N_2577,N_2326,N_2102);
or U2578 (N_2578,N_2230,N_2199);
and U2579 (N_2579,N_2397,N_2210);
or U2580 (N_2580,N_2082,N_2322);
xnor U2581 (N_2581,N_2075,N_2050);
xor U2582 (N_2582,N_2382,N_2024);
nor U2583 (N_2583,N_2111,N_2366);
nor U2584 (N_2584,N_2106,N_2064);
or U2585 (N_2585,N_2165,N_2079);
nand U2586 (N_2586,N_2129,N_2123);
xnor U2587 (N_2587,N_2241,N_2196);
and U2588 (N_2588,N_2217,N_2010);
and U2589 (N_2589,N_2187,N_2204);
and U2590 (N_2590,N_2043,N_2189);
xnor U2591 (N_2591,N_2392,N_2155);
nand U2592 (N_2592,N_2260,N_2053);
and U2593 (N_2593,N_2238,N_2371);
nor U2594 (N_2594,N_2346,N_2342);
nand U2595 (N_2595,N_2290,N_2384);
xnor U2596 (N_2596,N_2351,N_2362);
xnor U2597 (N_2597,N_2211,N_2247);
and U2598 (N_2598,N_2030,N_2182);
nand U2599 (N_2599,N_2036,N_2266);
nand U2600 (N_2600,N_2087,N_2184);
nand U2601 (N_2601,N_2306,N_2024);
and U2602 (N_2602,N_2137,N_2307);
nor U2603 (N_2603,N_2190,N_2353);
xnor U2604 (N_2604,N_2389,N_2013);
xor U2605 (N_2605,N_2119,N_2115);
nor U2606 (N_2606,N_2163,N_2072);
xor U2607 (N_2607,N_2270,N_2286);
xnor U2608 (N_2608,N_2239,N_2306);
and U2609 (N_2609,N_2254,N_2172);
or U2610 (N_2610,N_2345,N_2183);
and U2611 (N_2611,N_2229,N_2348);
and U2612 (N_2612,N_2250,N_2375);
xnor U2613 (N_2613,N_2245,N_2239);
xor U2614 (N_2614,N_2328,N_2199);
xor U2615 (N_2615,N_2284,N_2388);
nor U2616 (N_2616,N_2180,N_2059);
nand U2617 (N_2617,N_2186,N_2201);
or U2618 (N_2618,N_2093,N_2259);
nand U2619 (N_2619,N_2207,N_2021);
nor U2620 (N_2620,N_2260,N_2269);
nand U2621 (N_2621,N_2037,N_2197);
nand U2622 (N_2622,N_2070,N_2146);
xnor U2623 (N_2623,N_2038,N_2266);
xor U2624 (N_2624,N_2212,N_2361);
and U2625 (N_2625,N_2397,N_2301);
and U2626 (N_2626,N_2356,N_2185);
nor U2627 (N_2627,N_2124,N_2002);
nor U2628 (N_2628,N_2394,N_2052);
and U2629 (N_2629,N_2398,N_2387);
nand U2630 (N_2630,N_2225,N_2142);
and U2631 (N_2631,N_2363,N_2078);
and U2632 (N_2632,N_2210,N_2089);
xor U2633 (N_2633,N_2114,N_2195);
and U2634 (N_2634,N_2207,N_2276);
nand U2635 (N_2635,N_2049,N_2342);
nand U2636 (N_2636,N_2396,N_2139);
or U2637 (N_2637,N_2095,N_2000);
nor U2638 (N_2638,N_2231,N_2012);
nor U2639 (N_2639,N_2381,N_2186);
nor U2640 (N_2640,N_2381,N_2082);
or U2641 (N_2641,N_2151,N_2200);
and U2642 (N_2642,N_2166,N_2001);
nand U2643 (N_2643,N_2332,N_2361);
nand U2644 (N_2644,N_2354,N_2083);
or U2645 (N_2645,N_2126,N_2236);
nand U2646 (N_2646,N_2136,N_2373);
or U2647 (N_2647,N_2266,N_2117);
xor U2648 (N_2648,N_2352,N_2184);
nand U2649 (N_2649,N_2366,N_2230);
nand U2650 (N_2650,N_2304,N_2366);
nor U2651 (N_2651,N_2198,N_2180);
nor U2652 (N_2652,N_2127,N_2357);
and U2653 (N_2653,N_2063,N_2364);
or U2654 (N_2654,N_2257,N_2390);
or U2655 (N_2655,N_2308,N_2329);
nand U2656 (N_2656,N_2184,N_2254);
nand U2657 (N_2657,N_2031,N_2306);
nor U2658 (N_2658,N_2287,N_2239);
or U2659 (N_2659,N_2296,N_2385);
or U2660 (N_2660,N_2336,N_2352);
nor U2661 (N_2661,N_2066,N_2174);
xnor U2662 (N_2662,N_2182,N_2216);
xor U2663 (N_2663,N_2203,N_2125);
nor U2664 (N_2664,N_2327,N_2060);
and U2665 (N_2665,N_2391,N_2162);
or U2666 (N_2666,N_2007,N_2042);
and U2667 (N_2667,N_2231,N_2000);
nand U2668 (N_2668,N_2076,N_2069);
xnor U2669 (N_2669,N_2161,N_2091);
xnor U2670 (N_2670,N_2390,N_2111);
xnor U2671 (N_2671,N_2092,N_2114);
or U2672 (N_2672,N_2388,N_2048);
xnor U2673 (N_2673,N_2306,N_2106);
or U2674 (N_2674,N_2093,N_2209);
nor U2675 (N_2675,N_2242,N_2248);
and U2676 (N_2676,N_2027,N_2276);
nand U2677 (N_2677,N_2108,N_2046);
xnor U2678 (N_2678,N_2118,N_2187);
or U2679 (N_2679,N_2054,N_2132);
xnor U2680 (N_2680,N_2018,N_2043);
xor U2681 (N_2681,N_2208,N_2322);
nor U2682 (N_2682,N_2176,N_2083);
nand U2683 (N_2683,N_2182,N_2399);
or U2684 (N_2684,N_2376,N_2313);
and U2685 (N_2685,N_2213,N_2057);
or U2686 (N_2686,N_2211,N_2370);
nor U2687 (N_2687,N_2197,N_2082);
nor U2688 (N_2688,N_2231,N_2037);
xnor U2689 (N_2689,N_2084,N_2225);
nand U2690 (N_2690,N_2242,N_2319);
and U2691 (N_2691,N_2148,N_2153);
or U2692 (N_2692,N_2180,N_2388);
or U2693 (N_2693,N_2230,N_2143);
xor U2694 (N_2694,N_2011,N_2272);
nand U2695 (N_2695,N_2366,N_2052);
xor U2696 (N_2696,N_2376,N_2325);
and U2697 (N_2697,N_2175,N_2269);
xor U2698 (N_2698,N_2265,N_2118);
and U2699 (N_2699,N_2371,N_2332);
nand U2700 (N_2700,N_2119,N_2073);
and U2701 (N_2701,N_2108,N_2320);
or U2702 (N_2702,N_2081,N_2003);
nor U2703 (N_2703,N_2334,N_2385);
xor U2704 (N_2704,N_2151,N_2111);
nor U2705 (N_2705,N_2285,N_2301);
xnor U2706 (N_2706,N_2135,N_2044);
xor U2707 (N_2707,N_2064,N_2209);
or U2708 (N_2708,N_2129,N_2398);
nand U2709 (N_2709,N_2149,N_2056);
nor U2710 (N_2710,N_2093,N_2086);
and U2711 (N_2711,N_2369,N_2343);
nand U2712 (N_2712,N_2291,N_2216);
nand U2713 (N_2713,N_2390,N_2308);
or U2714 (N_2714,N_2026,N_2380);
or U2715 (N_2715,N_2398,N_2109);
nand U2716 (N_2716,N_2113,N_2147);
nor U2717 (N_2717,N_2108,N_2310);
nor U2718 (N_2718,N_2092,N_2079);
or U2719 (N_2719,N_2266,N_2231);
nor U2720 (N_2720,N_2063,N_2387);
and U2721 (N_2721,N_2100,N_2399);
nor U2722 (N_2722,N_2117,N_2070);
nand U2723 (N_2723,N_2119,N_2382);
and U2724 (N_2724,N_2189,N_2071);
and U2725 (N_2725,N_2276,N_2182);
nand U2726 (N_2726,N_2318,N_2212);
nand U2727 (N_2727,N_2210,N_2399);
xor U2728 (N_2728,N_2002,N_2014);
or U2729 (N_2729,N_2264,N_2379);
or U2730 (N_2730,N_2126,N_2241);
xor U2731 (N_2731,N_2333,N_2187);
or U2732 (N_2732,N_2158,N_2076);
or U2733 (N_2733,N_2275,N_2118);
nor U2734 (N_2734,N_2297,N_2316);
and U2735 (N_2735,N_2119,N_2340);
nand U2736 (N_2736,N_2202,N_2013);
and U2737 (N_2737,N_2271,N_2228);
xor U2738 (N_2738,N_2080,N_2165);
and U2739 (N_2739,N_2113,N_2355);
and U2740 (N_2740,N_2219,N_2076);
xnor U2741 (N_2741,N_2399,N_2251);
or U2742 (N_2742,N_2123,N_2016);
nand U2743 (N_2743,N_2395,N_2085);
xnor U2744 (N_2744,N_2018,N_2266);
nor U2745 (N_2745,N_2125,N_2187);
and U2746 (N_2746,N_2021,N_2232);
or U2747 (N_2747,N_2256,N_2257);
nand U2748 (N_2748,N_2012,N_2286);
xor U2749 (N_2749,N_2205,N_2253);
nor U2750 (N_2750,N_2214,N_2366);
or U2751 (N_2751,N_2300,N_2192);
and U2752 (N_2752,N_2354,N_2042);
nor U2753 (N_2753,N_2275,N_2023);
and U2754 (N_2754,N_2328,N_2150);
or U2755 (N_2755,N_2090,N_2333);
nor U2756 (N_2756,N_2195,N_2178);
and U2757 (N_2757,N_2187,N_2162);
xnor U2758 (N_2758,N_2271,N_2075);
nor U2759 (N_2759,N_2185,N_2353);
or U2760 (N_2760,N_2061,N_2272);
or U2761 (N_2761,N_2006,N_2371);
nand U2762 (N_2762,N_2137,N_2326);
xnor U2763 (N_2763,N_2284,N_2255);
nand U2764 (N_2764,N_2395,N_2325);
nor U2765 (N_2765,N_2075,N_2199);
nand U2766 (N_2766,N_2147,N_2285);
or U2767 (N_2767,N_2386,N_2270);
nor U2768 (N_2768,N_2143,N_2280);
or U2769 (N_2769,N_2382,N_2090);
or U2770 (N_2770,N_2107,N_2039);
or U2771 (N_2771,N_2323,N_2012);
or U2772 (N_2772,N_2112,N_2111);
nor U2773 (N_2773,N_2103,N_2267);
xor U2774 (N_2774,N_2361,N_2057);
nor U2775 (N_2775,N_2231,N_2048);
nor U2776 (N_2776,N_2226,N_2021);
xnor U2777 (N_2777,N_2190,N_2360);
xnor U2778 (N_2778,N_2164,N_2043);
xnor U2779 (N_2779,N_2377,N_2359);
nor U2780 (N_2780,N_2026,N_2278);
nor U2781 (N_2781,N_2111,N_2229);
and U2782 (N_2782,N_2233,N_2197);
or U2783 (N_2783,N_2223,N_2009);
nor U2784 (N_2784,N_2277,N_2264);
nand U2785 (N_2785,N_2194,N_2312);
nand U2786 (N_2786,N_2150,N_2090);
and U2787 (N_2787,N_2049,N_2291);
nand U2788 (N_2788,N_2148,N_2115);
nor U2789 (N_2789,N_2339,N_2273);
nor U2790 (N_2790,N_2078,N_2284);
xor U2791 (N_2791,N_2340,N_2039);
xor U2792 (N_2792,N_2010,N_2256);
nor U2793 (N_2793,N_2062,N_2216);
or U2794 (N_2794,N_2230,N_2214);
nor U2795 (N_2795,N_2354,N_2163);
nand U2796 (N_2796,N_2080,N_2117);
and U2797 (N_2797,N_2298,N_2013);
nand U2798 (N_2798,N_2184,N_2376);
nor U2799 (N_2799,N_2116,N_2270);
nand U2800 (N_2800,N_2702,N_2490);
nand U2801 (N_2801,N_2774,N_2770);
nand U2802 (N_2802,N_2452,N_2788);
xnor U2803 (N_2803,N_2686,N_2672);
or U2804 (N_2804,N_2640,N_2783);
nand U2805 (N_2805,N_2515,N_2603);
or U2806 (N_2806,N_2406,N_2442);
nand U2807 (N_2807,N_2456,N_2411);
nand U2808 (N_2808,N_2520,N_2680);
nor U2809 (N_2809,N_2528,N_2419);
and U2810 (N_2810,N_2580,N_2410);
nor U2811 (N_2811,N_2726,N_2545);
or U2812 (N_2812,N_2633,N_2649);
nand U2813 (N_2813,N_2499,N_2568);
nand U2814 (N_2814,N_2777,N_2542);
xnor U2815 (N_2815,N_2427,N_2594);
nand U2816 (N_2816,N_2500,N_2464);
or U2817 (N_2817,N_2573,N_2479);
or U2818 (N_2818,N_2562,N_2642);
nor U2819 (N_2819,N_2712,N_2740);
nand U2820 (N_2820,N_2448,N_2577);
or U2821 (N_2821,N_2509,N_2635);
nand U2822 (N_2822,N_2721,N_2485);
or U2823 (N_2823,N_2673,N_2742);
xor U2824 (N_2824,N_2625,N_2648);
nand U2825 (N_2825,N_2768,N_2558);
and U2826 (N_2826,N_2763,N_2614);
or U2827 (N_2827,N_2472,N_2478);
and U2828 (N_2828,N_2595,N_2604);
xnor U2829 (N_2829,N_2705,N_2759);
nand U2830 (N_2830,N_2549,N_2799);
nand U2831 (N_2831,N_2547,N_2766);
xnor U2832 (N_2832,N_2772,N_2677);
nor U2833 (N_2833,N_2522,N_2429);
nor U2834 (N_2834,N_2756,N_2486);
and U2835 (N_2835,N_2457,N_2465);
or U2836 (N_2836,N_2707,N_2557);
xor U2837 (N_2837,N_2647,N_2674);
and U2838 (N_2838,N_2591,N_2637);
nand U2839 (N_2839,N_2659,N_2449);
or U2840 (N_2840,N_2527,N_2761);
and U2841 (N_2841,N_2439,N_2598);
nand U2842 (N_2842,N_2618,N_2709);
or U2843 (N_2843,N_2744,N_2495);
or U2844 (N_2844,N_2785,N_2781);
or U2845 (N_2845,N_2664,N_2609);
nor U2846 (N_2846,N_2661,N_2634);
and U2847 (N_2847,N_2584,N_2581);
or U2848 (N_2848,N_2529,N_2590);
xor U2849 (N_2849,N_2616,N_2473);
or U2850 (N_2850,N_2643,N_2621);
xnor U2851 (N_2851,N_2612,N_2511);
nand U2852 (N_2852,N_2422,N_2600);
or U2853 (N_2853,N_2487,N_2698);
nand U2854 (N_2854,N_2446,N_2460);
or U2855 (N_2855,N_2741,N_2592);
or U2856 (N_2856,N_2715,N_2482);
nand U2857 (N_2857,N_2607,N_2402);
nand U2858 (N_2858,N_2583,N_2787);
and U2859 (N_2859,N_2719,N_2670);
nor U2860 (N_2860,N_2639,N_2469);
or U2861 (N_2861,N_2636,N_2501);
nand U2862 (N_2862,N_2694,N_2556);
xnor U2863 (N_2863,N_2574,N_2668);
nand U2864 (N_2864,N_2747,N_2748);
nor U2865 (N_2865,N_2657,N_2569);
and U2866 (N_2866,N_2773,N_2650);
and U2867 (N_2867,N_2714,N_2765);
xor U2868 (N_2868,N_2623,N_2723);
or U2869 (N_2869,N_2463,N_2521);
xor U2870 (N_2870,N_2754,N_2471);
or U2871 (N_2871,N_2455,N_2588);
nand U2872 (N_2872,N_2414,N_2493);
or U2873 (N_2873,N_2602,N_2537);
xor U2874 (N_2874,N_2481,N_2624);
and U2875 (N_2875,N_2572,N_2441);
xor U2876 (N_2876,N_2484,N_2786);
and U2877 (N_2877,N_2717,N_2552);
and U2878 (N_2878,N_2458,N_2738);
and U2879 (N_2879,N_2536,N_2506);
and U2880 (N_2880,N_2498,N_2737);
and U2881 (N_2881,N_2518,N_2587);
nand U2882 (N_2882,N_2666,N_2413);
nand U2883 (N_2883,N_2681,N_2401);
or U2884 (N_2884,N_2758,N_2533);
or U2885 (N_2885,N_2445,N_2760);
or U2886 (N_2886,N_2720,N_2660);
and U2887 (N_2887,N_2795,N_2571);
xnor U2888 (N_2888,N_2746,N_2652);
and U2889 (N_2889,N_2671,N_2412);
xor U2890 (N_2890,N_2767,N_2415);
nor U2891 (N_2891,N_2576,N_2444);
xor U2892 (N_2892,N_2676,N_2638);
nor U2893 (N_2893,N_2578,N_2755);
and U2894 (N_2894,N_2524,N_2693);
or U2895 (N_2895,N_2416,N_2459);
nor U2896 (N_2896,N_2585,N_2733);
or U2897 (N_2897,N_2728,N_2437);
and U2898 (N_2898,N_2778,N_2599);
or U2899 (N_2899,N_2434,N_2407);
or U2900 (N_2900,N_2436,N_2622);
nor U2901 (N_2901,N_2554,N_2409);
nand U2902 (N_2902,N_2789,N_2505);
nand U2903 (N_2903,N_2575,N_2739);
nand U2904 (N_2904,N_2691,N_2779);
nor U2905 (N_2905,N_2601,N_2764);
nand U2906 (N_2906,N_2539,N_2704);
and U2907 (N_2907,N_2752,N_2711);
nor U2908 (N_2908,N_2507,N_2503);
or U2909 (N_2909,N_2513,N_2796);
or U2910 (N_2910,N_2420,N_2532);
nor U2911 (N_2911,N_2404,N_2615);
nor U2912 (N_2912,N_2496,N_2735);
xor U2913 (N_2913,N_2790,N_2403);
nor U2914 (N_2914,N_2605,N_2596);
or U2915 (N_2915,N_2519,N_2468);
nand U2916 (N_2916,N_2516,N_2695);
nand U2917 (N_2917,N_2793,N_2613);
or U2918 (N_2918,N_2725,N_2631);
nand U2919 (N_2919,N_2586,N_2570);
nand U2920 (N_2920,N_2497,N_2757);
and U2921 (N_2921,N_2699,N_2654);
xor U2922 (N_2922,N_2491,N_2494);
and U2923 (N_2923,N_2651,N_2658);
nand U2924 (N_2924,N_2730,N_2476);
and U2925 (N_2925,N_2555,N_2474);
nor U2926 (N_2926,N_2559,N_2426);
nand U2927 (N_2927,N_2477,N_2563);
xnor U2928 (N_2928,N_2431,N_2608);
and U2929 (N_2929,N_2679,N_2645);
nand U2930 (N_2930,N_2492,N_2560);
xnor U2931 (N_2931,N_2689,N_2710);
nand U2932 (N_2932,N_2697,N_2690);
and U2933 (N_2933,N_2462,N_2701);
and U2934 (N_2934,N_2453,N_2762);
xor U2935 (N_2935,N_2713,N_2475);
nor U2936 (N_2936,N_2667,N_2450);
xor U2937 (N_2937,N_2408,N_2632);
nor U2938 (N_2938,N_2530,N_2470);
and U2939 (N_2939,N_2696,N_2687);
and U2940 (N_2940,N_2617,N_2646);
nor U2941 (N_2941,N_2589,N_2467);
nor U2942 (N_2942,N_2610,N_2708);
or U2943 (N_2943,N_2611,N_2619);
nand U2944 (N_2944,N_2579,N_2423);
xnor U2945 (N_2945,N_2743,N_2718);
nand U2946 (N_2946,N_2418,N_2692);
xnor U2947 (N_2947,N_2550,N_2510);
nand U2948 (N_2948,N_2544,N_2685);
and U2949 (N_2949,N_2502,N_2753);
and U2950 (N_2950,N_2797,N_2517);
nor U2951 (N_2951,N_2566,N_2706);
xor U2952 (N_2952,N_2641,N_2512);
nand U2953 (N_2953,N_2700,N_2424);
and U2954 (N_2954,N_2451,N_2428);
nand U2955 (N_2955,N_2421,N_2682);
xnor U2956 (N_2956,N_2736,N_2443);
and U2957 (N_2957,N_2433,N_2716);
nand U2958 (N_2958,N_2489,N_2644);
nand U2959 (N_2959,N_2731,N_2703);
nor U2960 (N_2960,N_2561,N_2724);
nand U2961 (N_2961,N_2483,N_2727);
or U2962 (N_2962,N_2553,N_2769);
or U2963 (N_2963,N_2628,N_2653);
nand U2964 (N_2964,N_2775,N_2734);
nor U2965 (N_2965,N_2488,N_2514);
nor U2966 (N_2966,N_2438,N_2729);
or U2967 (N_2967,N_2627,N_2548);
nand U2968 (N_2968,N_2663,N_2480);
and U2969 (N_2969,N_2523,N_2567);
xnor U2970 (N_2970,N_2425,N_2722);
nor U2971 (N_2971,N_2551,N_2750);
xnor U2972 (N_2972,N_2606,N_2688);
xor U2973 (N_2973,N_2794,N_2432);
nor U2974 (N_2974,N_2684,N_2656);
or U2975 (N_2975,N_2593,N_2626);
and U2976 (N_2976,N_2565,N_2400);
nor U2977 (N_2977,N_2678,N_2541);
and U2978 (N_2978,N_2780,N_2531);
or U2979 (N_2979,N_2798,N_2749);
xnor U2980 (N_2980,N_2461,N_2564);
nor U2981 (N_2981,N_2526,N_2597);
nand U2982 (N_2982,N_2417,N_2751);
xnor U2983 (N_2983,N_2540,N_2466);
nor U2984 (N_2984,N_2630,N_2534);
nor U2985 (N_2985,N_2675,N_2447);
xor U2986 (N_2986,N_2440,N_2538);
xnor U2987 (N_2987,N_2620,N_2535);
xnor U2988 (N_2988,N_2430,N_2504);
or U2989 (N_2989,N_2771,N_2732);
xnor U2990 (N_2990,N_2683,N_2776);
nand U2991 (N_2991,N_2745,N_2782);
xnor U2992 (N_2992,N_2405,N_2669);
xnor U2993 (N_2993,N_2791,N_2435);
nor U2994 (N_2994,N_2525,N_2546);
nand U2995 (N_2995,N_2792,N_2629);
or U2996 (N_2996,N_2665,N_2784);
and U2997 (N_2997,N_2543,N_2508);
xor U2998 (N_2998,N_2454,N_2662);
nand U2999 (N_2999,N_2582,N_2655);
nand U3000 (N_3000,N_2649,N_2673);
xor U3001 (N_3001,N_2567,N_2798);
nor U3002 (N_3002,N_2423,N_2617);
and U3003 (N_3003,N_2620,N_2497);
nand U3004 (N_3004,N_2469,N_2532);
xnor U3005 (N_3005,N_2558,N_2553);
nor U3006 (N_3006,N_2676,N_2791);
or U3007 (N_3007,N_2691,N_2669);
xnor U3008 (N_3008,N_2420,N_2450);
nand U3009 (N_3009,N_2526,N_2640);
or U3010 (N_3010,N_2530,N_2567);
nor U3011 (N_3011,N_2604,N_2597);
nand U3012 (N_3012,N_2442,N_2770);
xnor U3013 (N_3013,N_2545,N_2419);
or U3014 (N_3014,N_2431,N_2490);
or U3015 (N_3015,N_2699,N_2551);
xor U3016 (N_3016,N_2675,N_2427);
or U3017 (N_3017,N_2651,N_2497);
nand U3018 (N_3018,N_2691,N_2639);
or U3019 (N_3019,N_2465,N_2682);
and U3020 (N_3020,N_2744,N_2464);
xnor U3021 (N_3021,N_2733,N_2769);
or U3022 (N_3022,N_2563,N_2787);
nor U3023 (N_3023,N_2654,N_2770);
or U3024 (N_3024,N_2509,N_2484);
nor U3025 (N_3025,N_2481,N_2725);
xor U3026 (N_3026,N_2523,N_2502);
xor U3027 (N_3027,N_2602,N_2661);
xor U3028 (N_3028,N_2559,N_2668);
nand U3029 (N_3029,N_2697,N_2631);
and U3030 (N_3030,N_2779,N_2615);
or U3031 (N_3031,N_2416,N_2701);
xor U3032 (N_3032,N_2726,N_2490);
or U3033 (N_3033,N_2482,N_2471);
or U3034 (N_3034,N_2630,N_2758);
nor U3035 (N_3035,N_2652,N_2592);
or U3036 (N_3036,N_2692,N_2673);
and U3037 (N_3037,N_2777,N_2406);
and U3038 (N_3038,N_2538,N_2424);
nor U3039 (N_3039,N_2643,N_2703);
or U3040 (N_3040,N_2424,N_2632);
and U3041 (N_3041,N_2443,N_2729);
nor U3042 (N_3042,N_2640,N_2592);
nor U3043 (N_3043,N_2572,N_2599);
nor U3044 (N_3044,N_2718,N_2720);
nor U3045 (N_3045,N_2456,N_2655);
nand U3046 (N_3046,N_2795,N_2753);
nor U3047 (N_3047,N_2648,N_2563);
xor U3048 (N_3048,N_2732,N_2463);
nand U3049 (N_3049,N_2661,N_2734);
nor U3050 (N_3050,N_2508,N_2630);
and U3051 (N_3051,N_2655,N_2679);
xor U3052 (N_3052,N_2757,N_2760);
and U3053 (N_3053,N_2659,N_2711);
nand U3054 (N_3054,N_2472,N_2707);
xnor U3055 (N_3055,N_2426,N_2717);
nand U3056 (N_3056,N_2487,N_2542);
nand U3057 (N_3057,N_2510,N_2754);
or U3058 (N_3058,N_2669,N_2566);
nand U3059 (N_3059,N_2425,N_2542);
and U3060 (N_3060,N_2416,N_2778);
nand U3061 (N_3061,N_2711,N_2574);
or U3062 (N_3062,N_2731,N_2655);
nor U3063 (N_3063,N_2549,N_2592);
xnor U3064 (N_3064,N_2728,N_2679);
nand U3065 (N_3065,N_2411,N_2687);
nor U3066 (N_3066,N_2639,N_2544);
nand U3067 (N_3067,N_2736,N_2593);
or U3068 (N_3068,N_2593,N_2482);
nor U3069 (N_3069,N_2658,N_2706);
nand U3070 (N_3070,N_2676,N_2569);
nor U3071 (N_3071,N_2747,N_2704);
and U3072 (N_3072,N_2464,N_2445);
and U3073 (N_3073,N_2417,N_2604);
or U3074 (N_3074,N_2544,N_2612);
nand U3075 (N_3075,N_2610,N_2647);
or U3076 (N_3076,N_2485,N_2525);
xnor U3077 (N_3077,N_2529,N_2433);
xnor U3078 (N_3078,N_2469,N_2789);
nor U3079 (N_3079,N_2661,N_2515);
xnor U3080 (N_3080,N_2421,N_2564);
nand U3081 (N_3081,N_2505,N_2746);
or U3082 (N_3082,N_2639,N_2793);
xnor U3083 (N_3083,N_2777,N_2689);
xor U3084 (N_3084,N_2724,N_2710);
and U3085 (N_3085,N_2447,N_2767);
or U3086 (N_3086,N_2661,N_2470);
and U3087 (N_3087,N_2776,N_2593);
nand U3088 (N_3088,N_2787,N_2577);
and U3089 (N_3089,N_2508,N_2477);
or U3090 (N_3090,N_2550,N_2408);
xnor U3091 (N_3091,N_2655,N_2742);
and U3092 (N_3092,N_2503,N_2652);
and U3093 (N_3093,N_2623,N_2467);
nor U3094 (N_3094,N_2580,N_2683);
nand U3095 (N_3095,N_2747,N_2525);
and U3096 (N_3096,N_2472,N_2494);
nor U3097 (N_3097,N_2438,N_2686);
xor U3098 (N_3098,N_2552,N_2762);
nand U3099 (N_3099,N_2661,N_2773);
and U3100 (N_3100,N_2416,N_2564);
or U3101 (N_3101,N_2665,N_2456);
xor U3102 (N_3102,N_2704,N_2684);
and U3103 (N_3103,N_2410,N_2448);
nor U3104 (N_3104,N_2417,N_2708);
nand U3105 (N_3105,N_2748,N_2496);
xor U3106 (N_3106,N_2636,N_2703);
nand U3107 (N_3107,N_2445,N_2421);
and U3108 (N_3108,N_2779,N_2759);
or U3109 (N_3109,N_2568,N_2550);
and U3110 (N_3110,N_2487,N_2547);
nand U3111 (N_3111,N_2581,N_2432);
nand U3112 (N_3112,N_2414,N_2670);
xor U3113 (N_3113,N_2643,N_2458);
nor U3114 (N_3114,N_2593,N_2502);
nor U3115 (N_3115,N_2627,N_2606);
nand U3116 (N_3116,N_2499,N_2706);
xnor U3117 (N_3117,N_2664,N_2502);
or U3118 (N_3118,N_2517,N_2522);
nand U3119 (N_3119,N_2501,N_2528);
and U3120 (N_3120,N_2561,N_2685);
nor U3121 (N_3121,N_2593,N_2766);
nand U3122 (N_3122,N_2643,N_2566);
or U3123 (N_3123,N_2588,N_2510);
or U3124 (N_3124,N_2520,N_2498);
xor U3125 (N_3125,N_2489,N_2582);
nand U3126 (N_3126,N_2572,N_2702);
nor U3127 (N_3127,N_2465,N_2593);
nand U3128 (N_3128,N_2751,N_2586);
nor U3129 (N_3129,N_2492,N_2411);
nand U3130 (N_3130,N_2467,N_2541);
nand U3131 (N_3131,N_2505,N_2470);
and U3132 (N_3132,N_2727,N_2703);
and U3133 (N_3133,N_2554,N_2726);
or U3134 (N_3134,N_2615,N_2580);
nor U3135 (N_3135,N_2790,N_2672);
nor U3136 (N_3136,N_2689,N_2617);
or U3137 (N_3137,N_2657,N_2777);
xnor U3138 (N_3138,N_2547,N_2522);
xor U3139 (N_3139,N_2601,N_2628);
or U3140 (N_3140,N_2557,N_2406);
nor U3141 (N_3141,N_2416,N_2510);
or U3142 (N_3142,N_2590,N_2420);
and U3143 (N_3143,N_2569,N_2780);
nand U3144 (N_3144,N_2677,N_2605);
or U3145 (N_3145,N_2635,N_2696);
and U3146 (N_3146,N_2544,N_2418);
and U3147 (N_3147,N_2662,N_2530);
nor U3148 (N_3148,N_2680,N_2665);
or U3149 (N_3149,N_2764,N_2568);
xor U3150 (N_3150,N_2688,N_2515);
or U3151 (N_3151,N_2503,N_2647);
and U3152 (N_3152,N_2563,N_2502);
and U3153 (N_3153,N_2625,N_2571);
xor U3154 (N_3154,N_2410,N_2555);
or U3155 (N_3155,N_2718,N_2790);
nor U3156 (N_3156,N_2615,N_2671);
or U3157 (N_3157,N_2579,N_2628);
nand U3158 (N_3158,N_2714,N_2664);
or U3159 (N_3159,N_2780,N_2438);
and U3160 (N_3160,N_2506,N_2758);
nand U3161 (N_3161,N_2566,N_2693);
or U3162 (N_3162,N_2706,N_2581);
nand U3163 (N_3163,N_2579,N_2606);
xnor U3164 (N_3164,N_2611,N_2792);
xnor U3165 (N_3165,N_2786,N_2543);
nand U3166 (N_3166,N_2491,N_2513);
or U3167 (N_3167,N_2632,N_2531);
xor U3168 (N_3168,N_2596,N_2440);
nor U3169 (N_3169,N_2471,N_2432);
and U3170 (N_3170,N_2527,N_2788);
xor U3171 (N_3171,N_2437,N_2681);
or U3172 (N_3172,N_2636,N_2436);
and U3173 (N_3173,N_2715,N_2773);
and U3174 (N_3174,N_2651,N_2590);
and U3175 (N_3175,N_2662,N_2455);
and U3176 (N_3176,N_2796,N_2577);
or U3177 (N_3177,N_2663,N_2791);
and U3178 (N_3178,N_2586,N_2549);
or U3179 (N_3179,N_2655,N_2606);
and U3180 (N_3180,N_2487,N_2662);
nand U3181 (N_3181,N_2793,N_2524);
nand U3182 (N_3182,N_2506,N_2595);
nor U3183 (N_3183,N_2438,N_2401);
and U3184 (N_3184,N_2782,N_2735);
nor U3185 (N_3185,N_2619,N_2773);
nor U3186 (N_3186,N_2702,N_2495);
or U3187 (N_3187,N_2779,N_2731);
xnor U3188 (N_3188,N_2489,N_2400);
and U3189 (N_3189,N_2411,N_2663);
nor U3190 (N_3190,N_2793,N_2440);
nand U3191 (N_3191,N_2767,N_2436);
and U3192 (N_3192,N_2765,N_2766);
nor U3193 (N_3193,N_2769,N_2473);
or U3194 (N_3194,N_2797,N_2515);
nand U3195 (N_3195,N_2465,N_2543);
nor U3196 (N_3196,N_2554,N_2441);
and U3197 (N_3197,N_2753,N_2610);
nand U3198 (N_3198,N_2404,N_2691);
and U3199 (N_3199,N_2645,N_2584);
nand U3200 (N_3200,N_3010,N_2993);
and U3201 (N_3201,N_2909,N_2925);
nor U3202 (N_3202,N_2870,N_3057);
nor U3203 (N_3203,N_2894,N_3086);
xnor U3204 (N_3204,N_3099,N_3176);
and U3205 (N_3205,N_3000,N_3124);
and U3206 (N_3206,N_3035,N_2805);
and U3207 (N_3207,N_2841,N_2918);
xor U3208 (N_3208,N_3115,N_2911);
and U3209 (N_3209,N_2825,N_3062);
and U3210 (N_3210,N_2883,N_3047);
nor U3211 (N_3211,N_3043,N_2972);
xnor U3212 (N_3212,N_3050,N_2992);
or U3213 (N_3213,N_3056,N_2851);
and U3214 (N_3214,N_2952,N_2882);
nand U3215 (N_3215,N_2981,N_2937);
nor U3216 (N_3216,N_3156,N_2818);
or U3217 (N_3217,N_3072,N_3161);
and U3218 (N_3218,N_2812,N_3112);
or U3219 (N_3219,N_2915,N_2906);
nor U3220 (N_3220,N_2847,N_3140);
nand U3221 (N_3221,N_2879,N_3184);
nand U3222 (N_3222,N_3041,N_3085);
and U3223 (N_3223,N_2854,N_3172);
nand U3224 (N_3224,N_2919,N_2916);
nand U3225 (N_3225,N_3132,N_3191);
and U3226 (N_3226,N_2964,N_2904);
nand U3227 (N_3227,N_3053,N_3190);
nor U3228 (N_3228,N_3194,N_2950);
and U3229 (N_3229,N_3147,N_3187);
nand U3230 (N_3230,N_3048,N_3098);
nor U3231 (N_3231,N_3123,N_3101);
nor U3232 (N_3232,N_2913,N_2844);
nor U3233 (N_3233,N_3049,N_2941);
xnor U3234 (N_3234,N_3154,N_3185);
or U3235 (N_3235,N_3145,N_2938);
and U3236 (N_3236,N_2890,N_3074);
nor U3237 (N_3237,N_2803,N_2824);
nor U3238 (N_3238,N_3071,N_3068);
nor U3239 (N_3239,N_2830,N_3116);
xor U3240 (N_3240,N_2876,N_3066);
nor U3241 (N_3241,N_3054,N_2974);
nand U3242 (N_3242,N_2986,N_2936);
or U3243 (N_3243,N_2924,N_3005);
and U3244 (N_3244,N_3080,N_3175);
and U3245 (N_3245,N_3032,N_2880);
nor U3246 (N_3246,N_2802,N_2908);
or U3247 (N_3247,N_3103,N_2998);
nand U3248 (N_3248,N_3177,N_2966);
and U3249 (N_3249,N_2853,N_3199);
nand U3250 (N_3250,N_2875,N_3144);
xor U3251 (N_3251,N_3029,N_3107);
nand U3252 (N_3252,N_2929,N_3059);
and U3253 (N_3253,N_2995,N_3188);
or U3254 (N_3254,N_2867,N_2801);
xnor U3255 (N_3255,N_3164,N_3093);
xnor U3256 (N_3256,N_3195,N_3118);
nor U3257 (N_3257,N_3133,N_3028);
or U3258 (N_3258,N_2943,N_2808);
xnor U3259 (N_3259,N_3170,N_2874);
nand U3260 (N_3260,N_2900,N_3061);
xnor U3261 (N_3261,N_3044,N_3169);
or U3262 (N_3262,N_3090,N_3001);
or U3263 (N_3263,N_3075,N_3127);
nor U3264 (N_3264,N_3137,N_3025);
or U3265 (N_3265,N_3166,N_3129);
nor U3266 (N_3266,N_2817,N_3180);
or U3267 (N_3267,N_2951,N_2862);
or U3268 (N_3268,N_2920,N_2982);
nand U3269 (N_3269,N_2804,N_2921);
and U3270 (N_3270,N_2822,N_2944);
or U3271 (N_3271,N_2816,N_3130);
xor U3272 (N_3272,N_2835,N_3045);
or U3273 (N_3273,N_2831,N_3198);
xor U3274 (N_3274,N_3136,N_3165);
xnor U3275 (N_3275,N_3143,N_2836);
xnor U3276 (N_3276,N_2991,N_3120);
xor U3277 (N_3277,N_3135,N_2852);
nor U3278 (N_3278,N_2806,N_3146);
nor U3279 (N_3279,N_2829,N_2898);
and U3280 (N_3280,N_3018,N_3117);
or U3281 (N_3281,N_3004,N_2839);
xor U3282 (N_3282,N_2815,N_2855);
or U3283 (N_3283,N_3069,N_2869);
nor U3284 (N_3284,N_3158,N_2878);
or U3285 (N_3285,N_2907,N_2859);
nor U3286 (N_3286,N_3014,N_2948);
and U3287 (N_3287,N_2910,N_3163);
and U3288 (N_3288,N_3155,N_2902);
xnor U3289 (N_3289,N_3134,N_3174);
xor U3290 (N_3290,N_3179,N_2845);
or U3291 (N_3291,N_2860,N_3031);
or U3292 (N_3292,N_3036,N_3051);
or U3293 (N_3293,N_3026,N_2927);
xor U3294 (N_3294,N_3017,N_3009);
nor U3295 (N_3295,N_3067,N_2856);
nand U3296 (N_3296,N_2901,N_2984);
nand U3297 (N_3297,N_3173,N_2842);
and U3298 (N_3298,N_3110,N_2871);
nand U3299 (N_3299,N_2857,N_2828);
or U3300 (N_3300,N_2980,N_2814);
xor U3301 (N_3301,N_2926,N_3012);
or U3302 (N_3302,N_2826,N_3015);
nand U3303 (N_3303,N_3021,N_2807);
or U3304 (N_3304,N_2861,N_2858);
and U3305 (N_3305,N_3065,N_2811);
nor U3306 (N_3306,N_3142,N_3019);
nor U3307 (N_3307,N_3058,N_2928);
nand U3308 (N_3308,N_3192,N_2959);
nor U3309 (N_3309,N_3040,N_2810);
and U3310 (N_3310,N_2994,N_2935);
nor U3311 (N_3311,N_3104,N_3092);
nor U3312 (N_3312,N_3183,N_2899);
xor U3313 (N_3313,N_2837,N_2961);
and U3314 (N_3314,N_2989,N_2887);
and U3315 (N_3315,N_3128,N_2958);
nand U3316 (N_3316,N_3039,N_2912);
and U3317 (N_3317,N_3034,N_2983);
nor U3318 (N_3318,N_3149,N_3084);
and U3319 (N_3319,N_2872,N_2973);
or U3320 (N_3320,N_2886,N_3055);
xor U3321 (N_3321,N_3131,N_3159);
and U3322 (N_3322,N_2955,N_2820);
xor U3323 (N_3323,N_2965,N_3087);
xnor U3324 (N_3324,N_2939,N_3076);
nand U3325 (N_3325,N_2968,N_2813);
and U3326 (N_3326,N_2819,N_3020);
nand U3327 (N_3327,N_2963,N_2914);
or U3328 (N_3328,N_2970,N_3095);
nand U3329 (N_3329,N_2840,N_3186);
xor U3330 (N_3330,N_2903,N_2850);
and U3331 (N_3331,N_3013,N_2848);
or U3332 (N_3332,N_3016,N_2843);
and U3333 (N_3333,N_2873,N_2865);
and U3334 (N_3334,N_3168,N_3102);
and U3335 (N_3335,N_2881,N_3091);
and U3336 (N_3336,N_2864,N_2949);
or U3337 (N_3337,N_2891,N_3079);
nand U3338 (N_3338,N_2827,N_3150);
nand U3339 (N_3339,N_3151,N_3027);
nand U3340 (N_3340,N_2846,N_3167);
xor U3341 (N_3341,N_3193,N_2967);
and U3342 (N_3342,N_2885,N_2889);
or U3343 (N_3343,N_2800,N_3042);
nand U3344 (N_3344,N_2947,N_3037);
nand U3345 (N_3345,N_3052,N_2832);
nand U3346 (N_3346,N_3152,N_2996);
xor U3347 (N_3347,N_2834,N_2893);
or U3348 (N_3348,N_2987,N_2821);
and U3349 (N_3349,N_2975,N_3022);
xor U3350 (N_3350,N_3109,N_3106);
nor U3351 (N_3351,N_2990,N_2971);
or U3352 (N_3352,N_3141,N_2884);
and U3353 (N_3353,N_3077,N_3178);
nor U3354 (N_3354,N_3006,N_3023);
and U3355 (N_3355,N_3070,N_3060);
and U3356 (N_3356,N_3063,N_2888);
xor U3357 (N_3357,N_3100,N_2849);
xnor U3358 (N_3358,N_3111,N_3024);
xnor U3359 (N_3359,N_2868,N_2877);
xnor U3360 (N_3360,N_3181,N_3126);
nand U3361 (N_3361,N_3046,N_3094);
nand U3362 (N_3362,N_3113,N_2954);
and U3363 (N_3363,N_2946,N_2896);
xnor U3364 (N_3364,N_3119,N_2962);
xor U3365 (N_3365,N_3038,N_3189);
or U3366 (N_3366,N_3088,N_3073);
nand U3367 (N_3367,N_2978,N_2956);
and U3368 (N_3368,N_2923,N_3002);
nand U3369 (N_3369,N_2940,N_3081);
and U3370 (N_3370,N_2957,N_2931);
nand U3371 (N_3371,N_3033,N_2917);
xor U3372 (N_3372,N_2988,N_3197);
or U3373 (N_3373,N_2833,N_3003);
or U3374 (N_3374,N_2922,N_3139);
nand U3375 (N_3375,N_2895,N_3083);
nand U3376 (N_3376,N_2969,N_2905);
or U3377 (N_3377,N_3030,N_2897);
nand U3378 (N_3378,N_2976,N_2942);
xnor U3379 (N_3379,N_2977,N_3105);
and U3380 (N_3380,N_3011,N_3125);
nor U3381 (N_3381,N_2997,N_3064);
and U3382 (N_3382,N_3008,N_2809);
nand U3383 (N_3383,N_3108,N_2823);
nor U3384 (N_3384,N_2892,N_2933);
or U3385 (N_3385,N_3171,N_3148);
nor U3386 (N_3386,N_2838,N_3007);
nor U3387 (N_3387,N_2953,N_3162);
nand U3388 (N_3388,N_2934,N_2960);
or U3389 (N_3389,N_3114,N_3182);
and U3390 (N_3390,N_3078,N_3121);
nand U3391 (N_3391,N_2932,N_2985);
nand U3392 (N_3392,N_3082,N_3138);
or U3393 (N_3393,N_2930,N_2866);
xor U3394 (N_3394,N_3097,N_3089);
xnor U3395 (N_3395,N_3196,N_2863);
nand U3396 (N_3396,N_2999,N_3153);
xnor U3397 (N_3397,N_2979,N_2945);
or U3398 (N_3398,N_3122,N_3157);
xnor U3399 (N_3399,N_3160,N_3096);
or U3400 (N_3400,N_2815,N_3156);
xnor U3401 (N_3401,N_2827,N_2838);
xor U3402 (N_3402,N_2987,N_2915);
xor U3403 (N_3403,N_2856,N_2907);
or U3404 (N_3404,N_2805,N_2999);
or U3405 (N_3405,N_2912,N_3188);
nor U3406 (N_3406,N_2808,N_3191);
nor U3407 (N_3407,N_2829,N_2918);
xnor U3408 (N_3408,N_2872,N_2975);
xor U3409 (N_3409,N_2969,N_2846);
nand U3410 (N_3410,N_3071,N_2893);
nor U3411 (N_3411,N_3024,N_2995);
xor U3412 (N_3412,N_2963,N_3089);
xor U3413 (N_3413,N_3010,N_3163);
nor U3414 (N_3414,N_2974,N_3025);
and U3415 (N_3415,N_3173,N_3002);
or U3416 (N_3416,N_3145,N_3008);
and U3417 (N_3417,N_2845,N_2819);
nand U3418 (N_3418,N_2919,N_2801);
nand U3419 (N_3419,N_3131,N_2871);
nor U3420 (N_3420,N_2882,N_3036);
and U3421 (N_3421,N_3092,N_2878);
nand U3422 (N_3422,N_3174,N_3077);
or U3423 (N_3423,N_3047,N_2802);
nor U3424 (N_3424,N_3141,N_2800);
or U3425 (N_3425,N_3105,N_3110);
or U3426 (N_3426,N_2993,N_3103);
and U3427 (N_3427,N_2844,N_2806);
xor U3428 (N_3428,N_3064,N_3188);
xor U3429 (N_3429,N_3001,N_2816);
and U3430 (N_3430,N_3088,N_3036);
nand U3431 (N_3431,N_2991,N_3141);
nor U3432 (N_3432,N_3141,N_3105);
xnor U3433 (N_3433,N_3066,N_2885);
and U3434 (N_3434,N_2901,N_3137);
or U3435 (N_3435,N_2889,N_3120);
xnor U3436 (N_3436,N_2821,N_2970);
xor U3437 (N_3437,N_3111,N_2808);
xor U3438 (N_3438,N_3049,N_2827);
nand U3439 (N_3439,N_3154,N_2934);
and U3440 (N_3440,N_2937,N_2835);
and U3441 (N_3441,N_3052,N_2917);
and U3442 (N_3442,N_2891,N_2916);
nor U3443 (N_3443,N_3083,N_3053);
and U3444 (N_3444,N_3182,N_2996);
nor U3445 (N_3445,N_3004,N_3074);
or U3446 (N_3446,N_2987,N_3130);
nor U3447 (N_3447,N_3102,N_3151);
xor U3448 (N_3448,N_2870,N_3133);
nand U3449 (N_3449,N_2914,N_2897);
nand U3450 (N_3450,N_3159,N_2832);
or U3451 (N_3451,N_2860,N_3046);
nand U3452 (N_3452,N_2836,N_2927);
nand U3453 (N_3453,N_2850,N_2908);
or U3454 (N_3454,N_2836,N_3095);
or U3455 (N_3455,N_2992,N_2865);
nor U3456 (N_3456,N_2824,N_2883);
and U3457 (N_3457,N_3143,N_3157);
nor U3458 (N_3458,N_3004,N_2960);
xnor U3459 (N_3459,N_3002,N_2943);
nor U3460 (N_3460,N_3150,N_2910);
or U3461 (N_3461,N_3107,N_2901);
and U3462 (N_3462,N_3177,N_3172);
xor U3463 (N_3463,N_2972,N_2914);
or U3464 (N_3464,N_3049,N_2836);
nand U3465 (N_3465,N_2834,N_2816);
nor U3466 (N_3466,N_2831,N_3109);
xor U3467 (N_3467,N_2888,N_3137);
nand U3468 (N_3468,N_3110,N_3099);
xor U3469 (N_3469,N_3102,N_3040);
and U3470 (N_3470,N_2863,N_2857);
and U3471 (N_3471,N_2871,N_2909);
xnor U3472 (N_3472,N_2997,N_2916);
and U3473 (N_3473,N_2933,N_2921);
or U3474 (N_3474,N_3057,N_2910);
and U3475 (N_3475,N_3022,N_3017);
or U3476 (N_3476,N_3011,N_2885);
nand U3477 (N_3477,N_3052,N_2849);
nor U3478 (N_3478,N_2944,N_3043);
or U3479 (N_3479,N_2832,N_2841);
or U3480 (N_3480,N_3104,N_3147);
or U3481 (N_3481,N_2962,N_3056);
and U3482 (N_3482,N_3007,N_2869);
nor U3483 (N_3483,N_2846,N_2845);
xor U3484 (N_3484,N_2941,N_3183);
nand U3485 (N_3485,N_3070,N_2991);
or U3486 (N_3486,N_2922,N_2967);
nor U3487 (N_3487,N_2893,N_2869);
or U3488 (N_3488,N_2840,N_2820);
and U3489 (N_3489,N_2812,N_3047);
nor U3490 (N_3490,N_3131,N_3078);
and U3491 (N_3491,N_2951,N_2843);
xor U3492 (N_3492,N_2895,N_3126);
and U3493 (N_3493,N_2801,N_3109);
nor U3494 (N_3494,N_2834,N_2900);
xor U3495 (N_3495,N_3156,N_3107);
and U3496 (N_3496,N_3094,N_3148);
or U3497 (N_3497,N_2946,N_3043);
or U3498 (N_3498,N_2958,N_2896);
and U3499 (N_3499,N_2808,N_2881);
xnor U3500 (N_3500,N_2842,N_3116);
nand U3501 (N_3501,N_3104,N_3132);
xor U3502 (N_3502,N_2806,N_2814);
and U3503 (N_3503,N_3013,N_3177);
and U3504 (N_3504,N_3153,N_2843);
xor U3505 (N_3505,N_3083,N_2932);
nand U3506 (N_3506,N_2808,N_2871);
xnor U3507 (N_3507,N_3143,N_2872);
xnor U3508 (N_3508,N_2867,N_2917);
nand U3509 (N_3509,N_3192,N_3053);
nand U3510 (N_3510,N_2997,N_2837);
or U3511 (N_3511,N_3083,N_3179);
nand U3512 (N_3512,N_3043,N_2926);
nand U3513 (N_3513,N_2966,N_2801);
nor U3514 (N_3514,N_3159,N_2956);
or U3515 (N_3515,N_2865,N_2864);
nor U3516 (N_3516,N_2808,N_2945);
and U3517 (N_3517,N_2904,N_2939);
and U3518 (N_3518,N_2813,N_3036);
nor U3519 (N_3519,N_2989,N_2956);
or U3520 (N_3520,N_2829,N_2850);
nor U3521 (N_3521,N_2916,N_2900);
and U3522 (N_3522,N_2875,N_2884);
xor U3523 (N_3523,N_3023,N_3170);
or U3524 (N_3524,N_3095,N_3078);
and U3525 (N_3525,N_3168,N_2862);
and U3526 (N_3526,N_2993,N_3059);
xnor U3527 (N_3527,N_2917,N_2810);
xor U3528 (N_3528,N_2812,N_3062);
nor U3529 (N_3529,N_2964,N_3191);
or U3530 (N_3530,N_2930,N_3136);
nand U3531 (N_3531,N_2943,N_2830);
xor U3532 (N_3532,N_2804,N_2899);
xor U3533 (N_3533,N_2901,N_3115);
nor U3534 (N_3534,N_2986,N_2921);
nor U3535 (N_3535,N_2914,N_3143);
and U3536 (N_3536,N_2989,N_3074);
xnor U3537 (N_3537,N_3075,N_2894);
nor U3538 (N_3538,N_2812,N_3123);
nand U3539 (N_3539,N_2810,N_2842);
and U3540 (N_3540,N_3180,N_2905);
and U3541 (N_3541,N_2951,N_2915);
nand U3542 (N_3542,N_3059,N_3049);
or U3543 (N_3543,N_2969,N_2987);
xor U3544 (N_3544,N_3185,N_3175);
nand U3545 (N_3545,N_3106,N_2887);
nor U3546 (N_3546,N_3090,N_2936);
xor U3547 (N_3547,N_3066,N_3172);
xnor U3548 (N_3548,N_2851,N_2819);
xor U3549 (N_3549,N_3098,N_3190);
and U3550 (N_3550,N_2904,N_3026);
nor U3551 (N_3551,N_3056,N_2804);
nor U3552 (N_3552,N_2887,N_3167);
nor U3553 (N_3553,N_2895,N_3140);
nor U3554 (N_3554,N_2820,N_2967);
xor U3555 (N_3555,N_3124,N_2878);
or U3556 (N_3556,N_3129,N_3033);
xor U3557 (N_3557,N_3182,N_2885);
nand U3558 (N_3558,N_3011,N_3020);
nor U3559 (N_3559,N_2807,N_3153);
and U3560 (N_3560,N_3146,N_3117);
xnor U3561 (N_3561,N_2849,N_3058);
nand U3562 (N_3562,N_3128,N_3077);
nand U3563 (N_3563,N_2944,N_2952);
nor U3564 (N_3564,N_3022,N_3141);
and U3565 (N_3565,N_2977,N_3071);
nor U3566 (N_3566,N_3169,N_2812);
nor U3567 (N_3567,N_3185,N_2928);
nand U3568 (N_3568,N_3080,N_2964);
xnor U3569 (N_3569,N_3174,N_2970);
xnor U3570 (N_3570,N_2902,N_3024);
and U3571 (N_3571,N_3053,N_3172);
nor U3572 (N_3572,N_3128,N_2888);
and U3573 (N_3573,N_3145,N_3126);
nor U3574 (N_3574,N_3037,N_3040);
nor U3575 (N_3575,N_2870,N_3159);
nand U3576 (N_3576,N_3123,N_2803);
nand U3577 (N_3577,N_3038,N_2921);
xor U3578 (N_3578,N_3082,N_2832);
and U3579 (N_3579,N_3036,N_3143);
nor U3580 (N_3580,N_2854,N_3065);
nand U3581 (N_3581,N_2914,N_2953);
nor U3582 (N_3582,N_2825,N_2923);
or U3583 (N_3583,N_3127,N_2894);
and U3584 (N_3584,N_2921,N_3019);
or U3585 (N_3585,N_3008,N_3081);
or U3586 (N_3586,N_2870,N_2934);
nand U3587 (N_3587,N_2911,N_2809);
nor U3588 (N_3588,N_3128,N_3152);
nand U3589 (N_3589,N_2976,N_3077);
and U3590 (N_3590,N_3158,N_3144);
or U3591 (N_3591,N_3026,N_2945);
nand U3592 (N_3592,N_3113,N_3172);
xor U3593 (N_3593,N_3026,N_3192);
nor U3594 (N_3594,N_3074,N_2965);
and U3595 (N_3595,N_3162,N_2806);
nor U3596 (N_3596,N_3032,N_2956);
nor U3597 (N_3597,N_3075,N_3198);
nand U3598 (N_3598,N_2913,N_3175);
xnor U3599 (N_3599,N_3142,N_2808);
or U3600 (N_3600,N_3532,N_3390);
nor U3601 (N_3601,N_3321,N_3435);
and U3602 (N_3602,N_3535,N_3530);
xnor U3603 (N_3603,N_3387,N_3355);
and U3604 (N_3604,N_3445,N_3457);
nand U3605 (N_3605,N_3566,N_3385);
nand U3606 (N_3606,N_3436,N_3254);
xnor U3607 (N_3607,N_3307,N_3556);
xnor U3608 (N_3608,N_3454,N_3523);
or U3609 (N_3609,N_3204,N_3210);
and U3610 (N_3610,N_3518,N_3593);
nor U3611 (N_3611,N_3282,N_3559);
nor U3612 (N_3612,N_3586,N_3304);
or U3613 (N_3613,N_3303,N_3238);
or U3614 (N_3614,N_3400,N_3281);
nand U3615 (N_3615,N_3545,N_3336);
or U3616 (N_3616,N_3524,N_3391);
nand U3617 (N_3617,N_3581,N_3398);
nand U3618 (N_3618,N_3360,N_3473);
and U3619 (N_3619,N_3509,N_3252);
nand U3620 (N_3620,N_3257,N_3534);
nor U3621 (N_3621,N_3533,N_3245);
nor U3622 (N_3622,N_3450,N_3531);
and U3623 (N_3623,N_3225,N_3510);
or U3624 (N_3624,N_3364,N_3213);
xnor U3625 (N_3625,N_3411,N_3280);
nor U3626 (N_3626,N_3367,N_3599);
nand U3627 (N_3627,N_3244,N_3590);
or U3628 (N_3628,N_3591,N_3242);
nor U3629 (N_3629,N_3255,N_3262);
or U3630 (N_3630,N_3372,N_3481);
and U3631 (N_3631,N_3437,N_3350);
and U3632 (N_3632,N_3230,N_3462);
nor U3633 (N_3633,N_3594,N_3301);
nor U3634 (N_3634,N_3577,N_3337);
xor U3635 (N_3635,N_3413,N_3502);
xor U3636 (N_3636,N_3424,N_3451);
and U3637 (N_3637,N_3408,N_3380);
or U3638 (N_3638,N_3389,N_3520);
and U3639 (N_3639,N_3270,N_3206);
or U3640 (N_3640,N_3421,N_3460);
xnor U3641 (N_3641,N_3572,N_3399);
nor U3642 (N_3642,N_3203,N_3375);
xor U3643 (N_3643,N_3538,N_3309);
or U3644 (N_3644,N_3235,N_3563);
and U3645 (N_3645,N_3517,N_3357);
and U3646 (N_3646,N_3542,N_3208);
nand U3647 (N_3647,N_3453,N_3376);
xor U3648 (N_3648,N_3467,N_3278);
nand U3649 (N_3649,N_3403,N_3526);
or U3650 (N_3650,N_3381,N_3305);
or U3651 (N_3651,N_3342,N_3248);
xor U3652 (N_3652,N_3466,N_3491);
nor U3653 (N_3653,N_3271,N_3386);
or U3654 (N_3654,N_3499,N_3539);
and U3655 (N_3655,N_3316,N_3366);
or U3656 (N_3656,N_3211,N_3505);
nand U3657 (N_3657,N_3494,N_3267);
xnor U3658 (N_3658,N_3293,N_3547);
nor U3659 (N_3659,N_3444,N_3319);
xnor U3660 (N_3660,N_3279,N_3332);
nand U3661 (N_3661,N_3562,N_3475);
nand U3662 (N_3662,N_3228,N_3402);
nand U3663 (N_3663,N_3344,N_3504);
xor U3664 (N_3664,N_3277,N_3216);
xor U3665 (N_3665,N_3234,N_3229);
nor U3666 (N_3666,N_3331,N_3354);
xor U3667 (N_3667,N_3565,N_3345);
nand U3668 (N_3668,N_3479,N_3264);
and U3669 (N_3669,N_3485,N_3374);
xor U3670 (N_3670,N_3596,N_3495);
xnor U3671 (N_3671,N_3480,N_3379);
xnor U3672 (N_3672,N_3438,N_3439);
nor U3673 (N_3673,N_3202,N_3430);
xnor U3674 (N_3674,N_3236,N_3584);
or U3675 (N_3675,N_3492,N_3221);
nor U3676 (N_3676,N_3500,N_3231);
nand U3677 (N_3677,N_3348,N_3395);
or U3678 (N_3678,N_3300,N_3410);
xnor U3679 (N_3679,N_3498,N_3318);
xnor U3680 (N_3680,N_3392,N_3340);
or U3681 (N_3681,N_3476,N_3470);
nand U3682 (N_3682,N_3343,N_3256);
nand U3683 (N_3683,N_3461,N_3568);
nand U3684 (N_3684,N_3553,N_3418);
or U3685 (N_3685,N_3579,N_3478);
nor U3686 (N_3686,N_3283,N_3201);
xor U3687 (N_3687,N_3583,N_3570);
and U3688 (N_3688,N_3442,N_3223);
nor U3689 (N_3689,N_3456,N_3573);
xor U3690 (N_3690,N_3434,N_3261);
nand U3691 (N_3691,N_3429,N_3525);
or U3692 (N_3692,N_3263,N_3455);
and U3693 (N_3693,N_3362,N_3292);
nor U3694 (N_3694,N_3288,N_3446);
and U3695 (N_3695,N_3290,N_3295);
nor U3696 (N_3696,N_3541,N_3516);
xnor U3697 (N_3697,N_3401,N_3219);
nand U3698 (N_3698,N_3592,N_3415);
nand U3699 (N_3699,N_3508,N_3598);
and U3700 (N_3700,N_3511,N_3544);
nor U3701 (N_3701,N_3207,N_3515);
or U3702 (N_3702,N_3349,N_3514);
nand U3703 (N_3703,N_3464,N_3550);
xor U3704 (N_3704,N_3260,N_3302);
nand U3705 (N_3705,N_3521,N_3394);
nand U3706 (N_3706,N_3294,N_3370);
xor U3707 (N_3707,N_3320,N_3396);
xor U3708 (N_3708,N_3363,N_3426);
and U3709 (N_3709,N_3585,N_3589);
nand U3710 (N_3710,N_3468,N_3339);
and U3711 (N_3711,N_3503,N_3404);
nor U3712 (N_3712,N_3273,N_3465);
or U3713 (N_3713,N_3459,N_3458);
or U3714 (N_3714,N_3487,N_3449);
xnor U3715 (N_3715,N_3325,N_3406);
and U3716 (N_3716,N_3324,N_3346);
and U3717 (N_3717,N_3315,N_3249);
and U3718 (N_3718,N_3289,N_3486);
nor U3719 (N_3719,N_3285,N_3243);
xor U3720 (N_3720,N_3463,N_3432);
nand U3721 (N_3721,N_3259,N_3549);
nor U3722 (N_3722,N_3306,N_3347);
nor U3723 (N_3723,N_3373,N_3537);
nand U3724 (N_3724,N_3588,N_3443);
xor U3725 (N_3725,N_3308,N_3595);
nand U3726 (N_3726,N_3384,N_3569);
nand U3727 (N_3727,N_3469,N_3352);
or U3728 (N_3728,N_3368,N_3326);
and U3729 (N_3729,N_3507,N_3571);
and U3730 (N_3730,N_3296,N_3351);
xor U3731 (N_3731,N_3597,N_3484);
xor U3732 (N_3732,N_3582,N_3575);
and U3733 (N_3733,N_3226,N_3265);
nand U3734 (N_3734,N_3297,N_3274);
xor U3735 (N_3735,N_3431,N_3323);
nand U3736 (N_3736,N_3237,N_3557);
xor U3737 (N_3737,N_3452,N_3217);
or U3738 (N_3738,N_3209,N_3311);
or U3739 (N_3739,N_3501,N_3253);
nand U3740 (N_3740,N_3338,N_3477);
or U3741 (N_3741,N_3416,N_3382);
nand U3742 (N_3742,N_3528,N_3471);
and U3743 (N_3743,N_3328,N_3548);
xnor U3744 (N_3744,N_3567,N_3212);
and U3745 (N_3745,N_3417,N_3546);
nor U3746 (N_3746,N_3540,N_3286);
nor U3747 (N_3747,N_3555,N_3269);
nand U3748 (N_3748,N_3272,N_3275);
nand U3749 (N_3749,N_3359,N_3383);
xnor U3750 (N_3750,N_3448,N_3215);
and U3751 (N_3751,N_3497,N_3335);
xnor U3752 (N_3752,N_3493,N_3356);
nand U3753 (N_3753,N_3488,N_3353);
and U3754 (N_3754,N_3587,N_3218);
nand U3755 (N_3755,N_3420,N_3365);
and U3756 (N_3756,N_3564,N_3241);
or U3757 (N_3757,N_3371,N_3333);
or U3758 (N_3758,N_3580,N_3251);
and U3759 (N_3759,N_3266,N_3543);
nor U3760 (N_3760,N_3529,N_3258);
nor U3761 (N_3761,N_3239,N_3536);
or U3762 (N_3762,N_3388,N_3397);
nand U3763 (N_3763,N_3522,N_3232);
xnor U3764 (N_3764,N_3405,N_3287);
xnor U3765 (N_3765,N_3327,N_3447);
nor U3766 (N_3766,N_3512,N_3412);
or U3767 (N_3767,N_3276,N_3574);
or U3768 (N_3768,N_3341,N_3233);
nor U3769 (N_3769,N_3322,N_3425);
nor U3770 (N_3770,N_3284,N_3205);
nand U3771 (N_3771,N_3560,N_3489);
xnor U3772 (N_3772,N_3227,N_3299);
xnor U3773 (N_3773,N_3330,N_3378);
xnor U3774 (N_3774,N_3329,N_3558);
nand U3775 (N_3775,N_3291,N_3419);
or U3776 (N_3776,N_3441,N_3561);
xor U3777 (N_3777,N_3409,N_3423);
nor U3778 (N_3778,N_3427,N_3552);
and U3779 (N_3779,N_3268,N_3220);
or U3780 (N_3780,N_3224,N_3472);
xnor U3781 (N_3781,N_3250,N_3474);
and U3782 (N_3782,N_3496,N_3377);
xor U3783 (N_3783,N_3554,N_3310);
or U3784 (N_3784,N_3482,N_3312);
and U3785 (N_3785,N_3422,N_3246);
nand U3786 (N_3786,N_3483,N_3222);
xor U3787 (N_3787,N_3358,N_3576);
and U3788 (N_3788,N_3428,N_3551);
nor U3789 (N_3789,N_3490,N_3519);
and U3790 (N_3790,N_3527,N_3433);
nor U3791 (N_3791,N_3578,N_3298);
xor U3792 (N_3792,N_3513,N_3393);
xor U3793 (N_3793,N_3369,N_3407);
nor U3794 (N_3794,N_3317,N_3414);
nor U3795 (N_3795,N_3440,N_3200);
nor U3796 (N_3796,N_3314,N_3361);
nor U3797 (N_3797,N_3334,N_3506);
and U3798 (N_3798,N_3313,N_3240);
nor U3799 (N_3799,N_3247,N_3214);
and U3800 (N_3800,N_3304,N_3537);
xnor U3801 (N_3801,N_3584,N_3477);
xor U3802 (N_3802,N_3402,N_3595);
nor U3803 (N_3803,N_3253,N_3572);
or U3804 (N_3804,N_3376,N_3225);
nor U3805 (N_3805,N_3347,N_3200);
nor U3806 (N_3806,N_3534,N_3438);
or U3807 (N_3807,N_3419,N_3340);
and U3808 (N_3808,N_3313,N_3320);
or U3809 (N_3809,N_3331,N_3224);
nor U3810 (N_3810,N_3330,N_3553);
nand U3811 (N_3811,N_3272,N_3477);
or U3812 (N_3812,N_3599,N_3436);
or U3813 (N_3813,N_3565,N_3420);
nand U3814 (N_3814,N_3298,N_3273);
nand U3815 (N_3815,N_3267,N_3533);
and U3816 (N_3816,N_3298,N_3347);
and U3817 (N_3817,N_3343,N_3345);
nand U3818 (N_3818,N_3358,N_3508);
nand U3819 (N_3819,N_3374,N_3545);
nand U3820 (N_3820,N_3275,N_3504);
nor U3821 (N_3821,N_3362,N_3428);
nand U3822 (N_3822,N_3375,N_3250);
nand U3823 (N_3823,N_3482,N_3333);
nand U3824 (N_3824,N_3230,N_3479);
xnor U3825 (N_3825,N_3219,N_3492);
or U3826 (N_3826,N_3311,N_3577);
nand U3827 (N_3827,N_3315,N_3358);
or U3828 (N_3828,N_3425,N_3414);
nor U3829 (N_3829,N_3590,N_3463);
and U3830 (N_3830,N_3598,N_3329);
or U3831 (N_3831,N_3551,N_3384);
nand U3832 (N_3832,N_3311,N_3567);
nand U3833 (N_3833,N_3563,N_3297);
nor U3834 (N_3834,N_3219,N_3598);
xor U3835 (N_3835,N_3435,N_3324);
nand U3836 (N_3836,N_3538,N_3393);
xnor U3837 (N_3837,N_3318,N_3333);
and U3838 (N_3838,N_3560,N_3383);
xor U3839 (N_3839,N_3335,N_3593);
or U3840 (N_3840,N_3423,N_3503);
or U3841 (N_3841,N_3534,N_3503);
and U3842 (N_3842,N_3232,N_3207);
and U3843 (N_3843,N_3257,N_3418);
xor U3844 (N_3844,N_3413,N_3208);
nor U3845 (N_3845,N_3392,N_3342);
nand U3846 (N_3846,N_3317,N_3564);
nor U3847 (N_3847,N_3257,N_3412);
nor U3848 (N_3848,N_3553,N_3456);
and U3849 (N_3849,N_3396,N_3577);
nor U3850 (N_3850,N_3591,N_3343);
or U3851 (N_3851,N_3520,N_3223);
and U3852 (N_3852,N_3337,N_3371);
and U3853 (N_3853,N_3279,N_3503);
or U3854 (N_3854,N_3474,N_3452);
or U3855 (N_3855,N_3413,N_3381);
and U3856 (N_3856,N_3552,N_3289);
nand U3857 (N_3857,N_3396,N_3388);
or U3858 (N_3858,N_3290,N_3501);
nand U3859 (N_3859,N_3502,N_3540);
nor U3860 (N_3860,N_3477,N_3553);
nor U3861 (N_3861,N_3402,N_3382);
xnor U3862 (N_3862,N_3530,N_3270);
nand U3863 (N_3863,N_3282,N_3522);
and U3864 (N_3864,N_3304,N_3478);
nand U3865 (N_3865,N_3334,N_3519);
or U3866 (N_3866,N_3328,N_3597);
nor U3867 (N_3867,N_3329,N_3400);
nor U3868 (N_3868,N_3475,N_3571);
and U3869 (N_3869,N_3290,N_3251);
nor U3870 (N_3870,N_3452,N_3328);
or U3871 (N_3871,N_3549,N_3470);
and U3872 (N_3872,N_3302,N_3339);
and U3873 (N_3873,N_3513,N_3358);
nand U3874 (N_3874,N_3434,N_3396);
xor U3875 (N_3875,N_3395,N_3373);
xnor U3876 (N_3876,N_3300,N_3474);
or U3877 (N_3877,N_3258,N_3241);
nor U3878 (N_3878,N_3561,N_3324);
and U3879 (N_3879,N_3585,N_3450);
or U3880 (N_3880,N_3441,N_3342);
or U3881 (N_3881,N_3339,N_3249);
and U3882 (N_3882,N_3484,N_3406);
or U3883 (N_3883,N_3548,N_3477);
nand U3884 (N_3884,N_3201,N_3544);
or U3885 (N_3885,N_3579,N_3339);
nand U3886 (N_3886,N_3520,N_3491);
nand U3887 (N_3887,N_3411,N_3274);
and U3888 (N_3888,N_3547,N_3496);
or U3889 (N_3889,N_3328,N_3503);
nor U3890 (N_3890,N_3279,N_3570);
xnor U3891 (N_3891,N_3240,N_3545);
and U3892 (N_3892,N_3304,N_3265);
and U3893 (N_3893,N_3506,N_3508);
and U3894 (N_3894,N_3428,N_3291);
nand U3895 (N_3895,N_3236,N_3457);
xor U3896 (N_3896,N_3282,N_3214);
or U3897 (N_3897,N_3423,N_3517);
nand U3898 (N_3898,N_3470,N_3495);
and U3899 (N_3899,N_3450,N_3401);
xnor U3900 (N_3900,N_3547,N_3486);
xnor U3901 (N_3901,N_3486,N_3312);
and U3902 (N_3902,N_3569,N_3480);
nor U3903 (N_3903,N_3348,N_3261);
or U3904 (N_3904,N_3416,N_3305);
nor U3905 (N_3905,N_3437,N_3352);
or U3906 (N_3906,N_3236,N_3308);
and U3907 (N_3907,N_3446,N_3238);
or U3908 (N_3908,N_3579,N_3234);
xnor U3909 (N_3909,N_3390,N_3578);
nor U3910 (N_3910,N_3234,N_3283);
nand U3911 (N_3911,N_3214,N_3382);
and U3912 (N_3912,N_3514,N_3393);
and U3913 (N_3913,N_3377,N_3260);
nand U3914 (N_3914,N_3528,N_3487);
and U3915 (N_3915,N_3230,N_3457);
nand U3916 (N_3916,N_3382,N_3353);
or U3917 (N_3917,N_3570,N_3339);
nand U3918 (N_3918,N_3391,N_3450);
nand U3919 (N_3919,N_3309,N_3364);
nor U3920 (N_3920,N_3301,N_3313);
nand U3921 (N_3921,N_3347,N_3589);
or U3922 (N_3922,N_3522,N_3542);
or U3923 (N_3923,N_3540,N_3471);
nand U3924 (N_3924,N_3301,N_3480);
or U3925 (N_3925,N_3484,N_3310);
xor U3926 (N_3926,N_3392,N_3274);
nand U3927 (N_3927,N_3464,N_3486);
nand U3928 (N_3928,N_3410,N_3240);
and U3929 (N_3929,N_3590,N_3410);
nand U3930 (N_3930,N_3399,N_3513);
nand U3931 (N_3931,N_3319,N_3549);
nor U3932 (N_3932,N_3369,N_3475);
nor U3933 (N_3933,N_3566,N_3237);
xor U3934 (N_3934,N_3429,N_3254);
nand U3935 (N_3935,N_3329,N_3211);
xnor U3936 (N_3936,N_3259,N_3458);
nor U3937 (N_3937,N_3503,N_3408);
and U3938 (N_3938,N_3416,N_3242);
nor U3939 (N_3939,N_3397,N_3233);
or U3940 (N_3940,N_3227,N_3485);
nor U3941 (N_3941,N_3384,N_3362);
or U3942 (N_3942,N_3414,N_3565);
and U3943 (N_3943,N_3298,N_3551);
xnor U3944 (N_3944,N_3558,N_3277);
and U3945 (N_3945,N_3244,N_3571);
or U3946 (N_3946,N_3570,N_3519);
nor U3947 (N_3947,N_3488,N_3325);
nand U3948 (N_3948,N_3320,N_3346);
and U3949 (N_3949,N_3219,N_3417);
and U3950 (N_3950,N_3405,N_3334);
nand U3951 (N_3951,N_3511,N_3447);
or U3952 (N_3952,N_3484,N_3264);
xor U3953 (N_3953,N_3401,N_3482);
nand U3954 (N_3954,N_3529,N_3437);
and U3955 (N_3955,N_3464,N_3215);
nand U3956 (N_3956,N_3507,N_3585);
nor U3957 (N_3957,N_3497,N_3426);
nand U3958 (N_3958,N_3551,N_3307);
xnor U3959 (N_3959,N_3287,N_3339);
and U3960 (N_3960,N_3466,N_3404);
nand U3961 (N_3961,N_3326,N_3544);
nand U3962 (N_3962,N_3345,N_3590);
xor U3963 (N_3963,N_3508,N_3545);
nand U3964 (N_3964,N_3464,N_3420);
or U3965 (N_3965,N_3572,N_3219);
and U3966 (N_3966,N_3367,N_3226);
nand U3967 (N_3967,N_3483,N_3354);
or U3968 (N_3968,N_3345,N_3231);
xnor U3969 (N_3969,N_3336,N_3414);
xor U3970 (N_3970,N_3303,N_3272);
nor U3971 (N_3971,N_3291,N_3576);
and U3972 (N_3972,N_3310,N_3415);
and U3973 (N_3973,N_3465,N_3477);
and U3974 (N_3974,N_3470,N_3385);
and U3975 (N_3975,N_3347,N_3204);
nand U3976 (N_3976,N_3334,N_3591);
nand U3977 (N_3977,N_3425,N_3519);
xnor U3978 (N_3978,N_3360,N_3454);
or U3979 (N_3979,N_3206,N_3585);
xor U3980 (N_3980,N_3572,N_3282);
xor U3981 (N_3981,N_3536,N_3521);
xor U3982 (N_3982,N_3355,N_3250);
xnor U3983 (N_3983,N_3333,N_3381);
nand U3984 (N_3984,N_3452,N_3399);
nor U3985 (N_3985,N_3454,N_3527);
xnor U3986 (N_3986,N_3248,N_3349);
or U3987 (N_3987,N_3406,N_3256);
nand U3988 (N_3988,N_3483,N_3331);
or U3989 (N_3989,N_3443,N_3423);
and U3990 (N_3990,N_3214,N_3386);
nor U3991 (N_3991,N_3317,N_3405);
nor U3992 (N_3992,N_3414,N_3207);
xor U3993 (N_3993,N_3356,N_3530);
nor U3994 (N_3994,N_3566,N_3349);
nand U3995 (N_3995,N_3364,N_3593);
or U3996 (N_3996,N_3302,N_3341);
xnor U3997 (N_3997,N_3449,N_3502);
or U3998 (N_3998,N_3577,N_3550);
and U3999 (N_3999,N_3343,N_3389);
and U4000 (N_4000,N_3680,N_3864);
nand U4001 (N_4001,N_3863,N_3622);
xor U4002 (N_4002,N_3613,N_3719);
and U4003 (N_4003,N_3930,N_3875);
nand U4004 (N_4004,N_3760,N_3766);
nand U4005 (N_4005,N_3829,N_3817);
or U4006 (N_4006,N_3689,N_3934);
or U4007 (N_4007,N_3681,N_3605);
nand U4008 (N_4008,N_3634,N_3782);
xor U4009 (N_4009,N_3686,N_3606);
nor U4010 (N_4010,N_3789,N_3882);
or U4011 (N_4011,N_3845,N_3742);
or U4012 (N_4012,N_3933,N_3985);
nor U4013 (N_4013,N_3820,N_3832);
and U4014 (N_4014,N_3923,N_3873);
nor U4015 (N_4015,N_3773,N_3759);
nor U4016 (N_4016,N_3993,N_3772);
xnor U4017 (N_4017,N_3872,N_3885);
or U4018 (N_4018,N_3690,N_3717);
nor U4019 (N_4019,N_3611,N_3748);
xnor U4020 (N_4020,N_3657,N_3836);
nor U4021 (N_4021,N_3931,N_3977);
xnor U4022 (N_4022,N_3627,N_3951);
and U4023 (N_4023,N_3617,N_3929);
or U4024 (N_4024,N_3895,N_3948);
xor U4025 (N_4025,N_3837,N_3816);
nor U4026 (N_4026,N_3917,N_3850);
or U4027 (N_4027,N_3749,N_3721);
xor U4028 (N_4028,N_3735,N_3903);
xnor U4029 (N_4029,N_3950,N_3911);
nand U4030 (N_4030,N_3683,N_3778);
nand U4031 (N_4031,N_3830,N_3849);
nor U4032 (N_4032,N_3747,N_3843);
nand U4033 (N_4033,N_3907,N_3807);
or U4034 (N_4034,N_3635,N_3653);
or U4035 (N_4035,N_3600,N_3664);
or U4036 (N_4036,N_3645,N_3896);
or U4037 (N_4037,N_3608,N_3784);
or U4038 (N_4038,N_3987,N_3765);
or U4039 (N_4039,N_3770,N_3734);
xor U4040 (N_4040,N_3960,N_3607);
or U4041 (N_4041,N_3884,N_3900);
xnor U4042 (N_4042,N_3751,N_3716);
and U4043 (N_4043,N_3745,N_3732);
or U4044 (N_4044,N_3753,N_3965);
or U4045 (N_4045,N_3691,N_3641);
xnor U4046 (N_4046,N_3866,N_3713);
or U4047 (N_4047,N_3706,N_3955);
nor U4048 (N_4048,N_3990,N_3840);
nand U4049 (N_4049,N_3910,N_3636);
xor U4050 (N_4050,N_3906,N_3796);
and U4051 (N_4051,N_3915,N_3610);
xor U4052 (N_4052,N_3647,N_3892);
nand U4053 (N_4053,N_3656,N_3947);
nor U4054 (N_4054,N_3852,N_3808);
and U4055 (N_4055,N_3779,N_3880);
nor U4056 (N_4056,N_3997,N_3661);
and U4057 (N_4057,N_3888,N_3709);
nand U4058 (N_4058,N_3959,N_3899);
and U4059 (N_4059,N_3962,N_3777);
or U4060 (N_4060,N_3640,N_3924);
or U4061 (N_4061,N_3614,N_3637);
xor U4062 (N_4062,N_3769,N_3942);
or U4063 (N_4063,N_3901,N_3730);
nand U4064 (N_4064,N_3788,N_3938);
and U4065 (N_4065,N_3902,N_3795);
nor U4066 (N_4066,N_3806,N_3867);
xnor U4067 (N_4067,N_3886,N_3913);
or U4068 (N_4068,N_3940,N_3722);
nor U4069 (N_4069,N_3620,N_3909);
or U4070 (N_4070,N_3826,N_3660);
or U4071 (N_4071,N_3618,N_3746);
nand U4072 (N_4072,N_3694,N_3665);
nand U4073 (N_4073,N_3804,N_3776);
or U4074 (N_4074,N_3966,N_3976);
nand U4075 (N_4075,N_3714,N_3791);
xnor U4076 (N_4076,N_3961,N_3897);
or U4077 (N_4077,N_3630,N_3983);
xor U4078 (N_4078,N_3964,N_3710);
or U4079 (N_4079,N_3908,N_3616);
nand U4080 (N_4080,N_3720,N_3739);
nor U4081 (N_4081,N_3889,N_3932);
or U4082 (N_4082,N_3674,N_3649);
xnor U4083 (N_4083,N_3844,N_3684);
and U4084 (N_4084,N_3752,N_3705);
nand U4085 (N_4085,N_3638,N_3982);
and U4086 (N_4086,N_3787,N_3954);
and U4087 (N_4087,N_3935,N_3887);
or U4088 (N_4088,N_3673,N_3797);
or U4089 (N_4089,N_3658,N_3652);
or U4090 (N_4090,N_3912,N_3823);
xnor U4091 (N_4091,N_3890,N_3738);
nor U4092 (N_4092,N_3833,N_3898);
nor U4093 (N_4093,N_3715,N_3973);
nor U4094 (N_4094,N_3841,N_3968);
or U4095 (N_4095,N_3718,N_3944);
or U4096 (N_4096,N_3628,N_3857);
xor U4097 (N_4097,N_3891,N_3803);
nor U4098 (N_4098,N_3812,N_3633);
nand U4099 (N_4099,N_3919,N_3644);
and U4100 (N_4100,N_3991,N_3619);
or U4101 (N_4101,N_3838,N_3846);
nand U4102 (N_4102,N_3972,N_3854);
and U4103 (N_4103,N_3624,N_3648);
nor U4104 (N_4104,N_3995,N_3952);
or U4105 (N_4105,N_3802,N_3811);
xor U4106 (N_4106,N_3729,N_3741);
nor U4107 (N_4107,N_3615,N_3655);
or U4108 (N_4108,N_3786,N_3870);
or U4109 (N_4109,N_3904,N_3853);
nand U4110 (N_4110,N_3975,N_3970);
or U4111 (N_4111,N_3632,N_3957);
or U4112 (N_4112,N_3963,N_3956);
nor U4113 (N_4113,N_3663,N_3831);
nand U4114 (N_4114,N_3876,N_3727);
or U4115 (N_4115,N_3785,N_3750);
or U4116 (N_4116,N_3926,N_3743);
or U4117 (N_4117,N_3996,N_3978);
nand U4118 (N_4118,N_3819,N_3601);
nor U4119 (N_4119,N_3783,N_3822);
and U4120 (N_4120,N_3939,N_3894);
and U4121 (N_4121,N_3642,N_3754);
nand U4122 (N_4122,N_3639,N_3825);
nand U4123 (N_4123,N_3775,N_3744);
and U4124 (N_4124,N_3799,N_3669);
or U4125 (N_4125,N_3928,N_3862);
nand U4126 (N_4126,N_3800,N_3893);
nor U4127 (N_4127,N_3941,N_3755);
xnor U4128 (N_4128,N_3723,N_3842);
nor U4129 (N_4129,N_3953,N_3992);
xnor U4130 (N_4130,N_3676,N_3984);
nand U4131 (N_4131,N_3869,N_3974);
or U4132 (N_4132,N_3946,N_3659);
nor U4133 (N_4133,N_3677,N_3967);
nand U4134 (N_4134,N_3767,N_3865);
nand U4135 (N_4135,N_3625,N_3678);
or U4136 (N_4136,N_3654,N_3805);
and U4137 (N_4137,N_3835,N_3626);
nand U4138 (N_4138,N_3927,N_3814);
nand U4139 (N_4139,N_3612,N_3945);
and U4140 (N_4140,N_3700,N_3914);
xnor U4141 (N_4141,N_3604,N_3707);
xnor U4142 (N_4142,N_3859,N_3871);
nand U4143 (N_4143,N_3979,N_3858);
xor U4144 (N_4144,N_3736,N_3781);
nor U4145 (N_4145,N_3603,N_3971);
or U4146 (N_4146,N_3697,N_3667);
or U4147 (N_4147,N_3883,N_3988);
nor U4148 (N_4148,N_3763,N_3916);
or U4149 (N_4149,N_3815,N_3740);
nor U4150 (N_4150,N_3824,N_3695);
nand U4151 (N_4151,N_3925,N_3761);
nand U4152 (N_4152,N_3711,N_3792);
and U4153 (N_4153,N_3687,N_3801);
nor U4154 (N_4154,N_3774,N_3703);
nand U4155 (N_4155,N_3877,N_3969);
nor U4156 (N_4156,N_3981,N_3847);
nand U4157 (N_4157,N_3623,N_3696);
nand U4158 (N_4158,N_3949,N_3794);
or U4159 (N_4159,N_3943,N_3675);
xor U4160 (N_4160,N_3855,N_3834);
or U4161 (N_4161,N_3643,N_3856);
xnor U4162 (N_4162,N_3921,N_3813);
or U4163 (N_4163,N_3768,N_3712);
or U4164 (N_4164,N_3688,N_3671);
nand U4165 (N_4165,N_3685,N_3733);
nor U4166 (N_4166,N_3698,N_3672);
or U4167 (N_4167,N_3980,N_3692);
and U4168 (N_4168,N_3629,N_3994);
and U4169 (N_4169,N_3693,N_3848);
or U4170 (N_4170,N_3918,N_3726);
nand U4171 (N_4171,N_3810,N_3728);
nand U4172 (N_4172,N_3737,N_3851);
and U4173 (N_4173,N_3679,N_3936);
and U4174 (N_4174,N_3874,N_3821);
nand U4175 (N_4175,N_3758,N_3708);
xnor U4176 (N_4176,N_3868,N_3879);
and U4177 (N_4177,N_3651,N_3798);
xor U4178 (N_4178,N_3670,N_3861);
nand U4179 (N_4179,N_3818,N_3937);
or U4180 (N_4180,N_3682,N_3986);
nand U4181 (N_4181,N_3958,N_3780);
or U4182 (N_4182,N_3757,N_3828);
nor U4183 (N_4183,N_3790,N_3602);
or U4184 (N_4184,N_3998,N_3650);
xor U4185 (N_4185,N_3905,N_3662);
or U4186 (N_4186,N_3839,N_3793);
or U4187 (N_4187,N_3704,N_3631);
xnor U4188 (N_4188,N_3922,N_3756);
or U4189 (N_4189,N_3621,N_3878);
and U4190 (N_4190,N_3666,N_3731);
or U4191 (N_4191,N_3702,N_3999);
or U4192 (N_4192,N_3989,N_3762);
nor U4193 (N_4193,N_3860,N_3699);
nand U4194 (N_4194,N_3827,N_3764);
nor U4195 (N_4195,N_3809,N_3668);
nand U4196 (N_4196,N_3609,N_3771);
nand U4197 (N_4197,N_3725,N_3701);
nand U4198 (N_4198,N_3646,N_3881);
and U4199 (N_4199,N_3724,N_3920);
and U4200 (N_4200,N_3640,N_3960);
and U4201 (N_4201,N_3846,N_3678);
or U4202 (N_4202,N_3928,N_3918);
xnor U4203 (N_4203,N_3805,N_3701);
or U4204 (N_4204,N_3717,N_3899);
and U4205 (N_4205,N_3658,N_3847);
xor U4206 (N_4206,N_3674,N_3834);
or U4207 (N_4207,N_3616,N_3638);
or U4208 (N_4208,N_3820,N_3848);
nand U4209 (N_4209,N_3847,N_3860);
nor U4210 (N_4210,N_3854,N_3675);
xnor U4211 (N_4211,N_3965,N_3823);
or U4212 (N_4212,N_3884,N_3899);
or U4213 (N_4213,N_3915,N_3866);
xnor U4214 (N_4214,N_3894,N_3684);
xnor U4215 (N_4215,N_3797,N_3868);
xor U4216 (N_4216,N_3646,N_3820);
and U4217 (N_4217,N_3930,N_3888);
nor U4218 (N_4218,N_3815,N_3738);
xnor U4219 (N_4219,N_3691,N_3628);
nand U4220 (N_4220,N_3890,N_3707);
xnor U4221 (N_4221,N_3839,N_3704);
xor U4222 (N_4222,N_3960,N_3694);
xor U4223 (N_4223,N_3707,N_3726);
or U4224 (N_4224,N_3818,N_3982);
and U4225 (N_4225,N_3724,N_3956);
and U4226 (N_4226,N_3972,N_3713);
nand U4227 (N_4227,N_3737,N_3928);
nor U4228 (N_4228,N_3886,N_3709);
nor U4229 (N_4229,N_3744,N_3705);
xnor U4230 (N_4230,N_3978,N_3745);
xor U4231 (N_4231,N_3865,N_3746);
or U4232 (N_4232,N_3918,N_3729);
or U4233 (N_4233,N_3683,N_3686);
and U4234 (N_4234,N_3765,N_3700);
nand U4235 (N_4235,N_3890,N_3713);
and U4236 (N_4236,N_3749,N_3629);
or U4237 (N_4237,N_3795,N_3629);
or U4238 (N_4238,N_3705,N_3757);
nand U4239 (N_4239,N_3627,N_3875);
or U4240 (N_4240,N_3842,N_3676);
nor U4241 (N_4241,N_3747,N_3943);
nand U4242 (N_4242,N_3713,N_3652);
and U4243 (N_4243,N_3633,N_3668);
nor U4244 (N_4244,N_3731,N_3618);
or U4245 (N_4245,N_3977,N_3965);
nor U4246 (N_4246,N_3962,N_3651);
nor U4247 (N_4247,N_3706,N_3867);
or U4248 (N_4248,N_3623,N_3743);
and U4249 (N_4249,N_3865,N_3948);
xnor U4250 (N_4250,N_3624,N_3674);
and U4251 (N_4251,N_3869,N_3876);
nor U4252 (N_4252,N_3719,N_3747);
and U4253 (N_4253,N_3658,N_3672);
nor U4254 (N_4254,N_3735,N_3822);
nor U4255 (N_4255,N_3646,N_3622);
xor U4256 (N_4256,N_3641,N_3723);
nor U4257 (N_4257,N_3720,N_3689);
xor U4258 (N_4258,N_3696,N_3650);
nor U4259 (N_4259,N_3858,N_3660);
or U4260 (N_4260,N_3879,N_3804);
or U4261 (N_4261,N_3690,N_3669);
nand U4262 (N_4262,N_3760,N_3771);
nor U4263 (N_4263,N_3918,N_3848);
and U4264 (N_4264,N_3829,N_3863);
nor U4265 (N_4265,N_3670,N_3918);
xor U4266 (N_4266,N_3857,N_3675);
or U4267 (N_4267,N_3660,N_3654);
nand U4268 (N_4268,N_3804,N_3634);
xor U4269 (N_4269,N_3972,N_3824);
or U4270 (N_4270,N_3656,N_3883);
xnor U4271 (N_4271,N_3854,N_3887);
and U4272 (N_4272,N_3961,N_3939);
nand U4273 (N_4273,N_3741,N_3780);
nor U4274 (N_4274,N_3811,N_3940);
or U4275 (N_4275,N_3902,N_3861);
nor U4276 (N_4276,N_3985,N_3804);
and U4277 (N_4277,N_3845,N_3780);
and U4278 (N_4278,N_3689,N_3919);
nand U4279 (N_4279,N_3606,N_3793);
nand U4280 (N_4280,N_3650,N_3661);
xor U4281 (N_4281,N_3801,N_3806);
or U4282 (N_4282,N_3766,N_3921);
nand U4283 (N_4283,N_3971,N_3689);
or U4284 (N_4284,N_3639,N_3646);
nor U4285 (N_4285,N_3924,N_3844);
or U4286 (N_4286,N_3776,N_3948);
nor U4287 (N_4287,N_3641,N_3979);
nor U4288 (N_4288,N_3934,N_3794);
xor U4289 (N_4289,N_3996,N_3865);
nand U4290 (N_4290,N_3865,N_3679);
nand U4291 (N_4291,N_3688,N_3676);
xor U4292 (N_4292,N_3658,N_3767);
nor U4293 (N_4293,N_3968,N_3692);
and U4294 (N_4294,N_3747,N_3993);
and U4295 (N_4295,N_3679,N_3856);
or U4296 (N_4296,N_3876,N_3868);
or U4297 (N_4297,N_3721,N_3775);
or U4298 (N_4298,N_3851,N_3621);
nor U4299 (N_4299,N_3642,N_3963);
nor U4300 (N_4300,N_3632,N_3960);
xnor U4301 (N_4301,N_3668,N_3772);
xnor U4302 (N_4302,N_3634,N_3846);
nor U4303 (N_4303,N_3851,N_3653);
nand U4304 (N_4304,N_3740,N_3691);
nor U4305 (N_4305,N_3919,N_3987);
and U4306 (N_4306,N_3834,N_3629);
or U4307 (N_4307,N_3918,N_3903);
nand U4308 (N_4308,N_3783,N_3937);
nand U4309 (N_4309,N_3995,N_3659);
nand U4310 (N_4310,N_3655,N_3916);
or U4311 (N_4311,N_3870,N_3636);
nor U4312 (N_4312,N_3611,N_3675);
nand U4313 (N_4313,N_3686,N_3857);
or U4314 (N_4314,N_3609,N_3923);
nor U4315 (N_4315,N_3654,N_3846);
xnor U4316 (N_4316,N_3774,N_3994);
xnor U4317 (N_4317,N_3814,N_3979);
and U4318 (N_4318,N_3690,N_3897);
or U4319 (N_4319,N_3989,N_3994);
nor U4320 (N_4320,N_3638,N_3735);
nor U4321 (N_4321,N_3641,N_3988);
nor U4322 (N_4322,N_3684,N_3906);
and U4323 (N_4323,N_3653,N_3629);
nor U4324 (N_4324,N_3811,N_3744);
and U4325 (N_4325,N_3891,N_3611);
and U4326 (N_4326,N_3837,N_3903);
and U4327 (N_4327,N_3722,N_3833);
and U4328 (N_4328,N_3742,N_3886);
and U4329 (N_4329,N_3673,N_3791);
or U4330 (N_4330,N_3957,N_3729);
nor U4331 (N_4331,N_3754,N_3730);
xor U4332 (N_4332,N_3755,N_3968);
or U4333 (N_4333,N_3862,N_3660);
xor U4334 (N_4334,N_3722,N_3757);
nor U4335 (N_4335,N_3686,N_3782);
or U4336 (N_4336,N_3601,N_3636);
or U4337 (N_4337,N_3820,N_3856);
or U4338 (N_4338,N_3627,N_3922);
and U4339 (N_4339,N_3614,N_3992);
or U4340 (N_4340,N_3669,N_3910);
and U4341 (N_4341,N_3763,N_3810);
or U4342 (N_4342,N_3811,N_3866);
xnor U4343 (N_4343,N_3780,N_3638);
nand U4344 (N_4344,N_3781,N_3909);
nand U4345 (N_4345,N_3733,N_3989);
and U4346 (N_4346,N_3691,N_3853);
nor U4347 (N_4347,N_3953,N_3624);
nand U4348 (N_4348,N_3934,N_3718);
and U4349 (N_4349,N_3608,N_3897);
or U4350 (N_4350,N_3951,N_3832);
and U4351 (N_4351,N_3658,N_3827);
and U4352 (N_4352,N_3757,N_3939);
nor U4353 (N_4353,N_3675,N_3864);
nor U4354 (N_4354,N_3940,N_3934);
and U4355 (N_4355,N_3848,N_3621);
and U4356 (N_4356,N_3847,N_3669);
nand U4357 (N_4357,N_3801,N_3622);
and U4358 (N_4358,N_3869,N_3652);
or U4359 (N_4359,N_3706,N_3813);
xor U4360 (N_4360,N_3877,N_3652);
nor U4361 (N_4361,N_3734,N_3609);
xnor U4362 (N_4362,N_3976,N_3998);
nand U4363 (N_4363,N_3739,N_3751);
xor U4364 (N_4364,N_3801,N_3726);
xor U4365 (N_4365,N_3953,N_3663);
nand U4366 (N_4366,N_3939,N_3731);
nor U4367 (N_4367,N_3735,N_3805);
nand U4368 (N_4368,N_3720,N_3840);
xnor U4369 (N_4369,N_3671,N_3849);
nand U4370 (N_4370,N_3637,N_3829);
and U4371 (N_4371,N_3995,N_3719);
xnor U4372 (N_4372,N_3937,N_3732);
xor U4373 (N_4373,N_3882,N_3940);
nor U4374 (N_4374,N_3778,N_3670);
xor U4375 (N_4375,N_3968,N_3631);
nor U4376 (N_4376,N_3903,N_3784);
xnor U4377 (N_4377,N_3991,N_3822);
and U4378 (N_4378,N_3673,N_3627);
and U4379 (N_4379,N_3680,N_3612);
xnor U4380 (N_4380,N_3952,N_3755);
or U4381 (N_4381,N_3766,N_3834);
nand U4382 (N_4382,N_3833,N_3837);
and U4383 (N_4383,N_3680,N_3802);
and U4384 (N_4384,N_3644,N_3763);
nor U4385 (N_4385,N_3930,N_3733);
xnor U4386 (N_4386,N_3766,N_3791);
or U4387 (N_4387,N_3761,N_3980);
and U4388 (N_4388,N_3859,N_3745);
xor U4389 (N_4389,N_3688,N_3628);
nand U4390 (N_4390,N_3610,N_3954);
xor U4391 (N_4391,N_3742,N_3787);
nand U4392 (N_4392,N_3777,N_3944);
nand U4393 (N_4393,N_3723,N_3683);
or U4394 (N_4394,N_3720,N_3771);
xor U4395 (N_4395,N_3806,N_3662);
and U4396 (N_4396,N_3949,N_3765);
or U4397 (N_4397,N_3704,N_3942);
xnor U4398 (N_4398,N_3672,N_3887);
xor U4399 (N_4399,N_3634,N_3952);
xor U4400 (N_4400,N_4207,N_4253);
or U4401 (N_4401,N_4112,N_4243);
and U4402 (N_4402,N_4359,N_4300);
and U4403 (N_4403,N_4092,N_4064);
xnor U4404 (N_4404,N_4339,N_4127);
xor U4405 (N_4405,N_4031,N_4372);
nand U4406 (N_4406,N_4148,N_4356);
or U4407 (N_4407,N_4036,N_4371);
nor U4408 (N_4408,N_4061,N_4394);
xor U4409 (N_4409,N_4101,N_4119);
nor U4410 (N_4410,N_4305,N_4073);
nor U4411 (N_4411,N_4156,N_4026);
xnor U4412 (N_4412,N_4290,N_4087);
nor U4413 (N_4413,N_4147,N_4267);
xor U4414 (N_4414,N_4179,N_4353);
or U4415 (N_4415,N_4355,N_4387);
nand U4416 (N_4416,N_4354,N_4192);
nand U4417 (N_4417,N_4367,N_4198);
or U4418 (N_4418,N_4158,N_4130);
xor U4419 (N_4419,N_4074,N_4384);
and U4420 (N_4420,N_4103,N_4399);
nor U4421 (N_4421,N_4320,N_4117);
or U4422 (N_4422,N_4168,N_4204);
nor U4423 (N_4423,N_4197,N_4069);
xnor U4424 (N_4424,N_4319,N_4047);
or U4425 (N_4425,N_4178,N_4196);
and U4426 (N_4426,N_4341,N_4011);
xor U4427 (N_4427,N_4102,N_4262);
nor U4428 (N_4428,N_4208,N_4050);
nor U4429 (N_4429,N_4080,N_4374);
xor U4430 (N_4430,N_4020,N_4019);
or U4431 (N_4431,N_4155,N_4000);
xnor U4432 (N_4432,N_4239,N_4330);
nand U4433 (N_4433,N_4043,N_4125);
nand U4434 (N_4434,N_4212,N_4235);
and U4435 (N_4435,N_4266,N_4039);
and U4436 (N_4436,N_4052,N_4062);
and U4437 (N_4437,N_4346,N_4098);
or U4438 (N_4438,N_4199,N_4307);
and U4439 (N_4439,N_4395,N_4351);
nand U4440 (N_4440,N_4280,N_4210);
nor U4441 (N_4441,N_4077,N_4070);
nor U4442 (N_4442,N_4358,N_4301);
xor U4443 (N_4443,N_4334,N_4076);
nor U4444 (N_4444,N_4265,N_4299);
nand U4445 (N_4445,N_4288,N_4390);
nand U4446 (N_4446,N_4032,N_4397);
nand U4447 (N_4447,N_4206,N_4377);
xnor U4448 (N_4448,N_4063,N_4289);
nor U4449 (N_4449,N_4256,N_4304);
xor U4450 (N_4450,N_4149,N_4398);
or U4451 (N_4451,N_4317,N_4163);
xor U4452 (N_4452,N_4223,N_4093);
nor U4453 (N_4453,N_4051,N_4183);
or U4454 (N_4454,N_4042,N_4392);
xnor U4455 (N_4455,N_4040,N_4217);
or U4456 (N_4456,N_4201,N_4314);
nand U4457 (N_4457,N_4056,N_4246);
or U4458 (N_4458,N_4231,N_4382);
xor U4459 (N_4459,N_4283,N_4129);
nand U4460 (N_4460,N_4181,N_4272);
and U4461 (N_4461,N_4104,N_4139);
xor U4462 (N_4462,N_4228,N_4381);
nand U4463 (N_4463,N_4234,N_4105);
nor U4464 (N_4464,N_4194,N_4275);
or U4465 (N_4465,N_4164,N_4325);
nand U4466 (N_4466,N_4328,N_4251);
or U4467 (N_4467,N_4257,N_4360);
nor U4468 (N_4468,N_4128,N_4009);
xnor U4469 (N_4469,N_4028,N_4295);
nor U4470 (N_4470,N_4068,N_4321);
xor U4471 (N_4471,N_4385,N_4236);
nor U4472 (N_4472,N_4309,N_4244);
xor U4473 (N_4473,N_4143,N_4035);
or U4474 (N_4474,N_4086,N_4136);
nor U4475 (N_4475,N_4135,N_4015);
nand U4476 (N_4476,N_4190,N_4099);
or U4477 (N_4477,N_4344,N_4030);
or U4478 (N_4478,N_4368,N_4270);
nor U4479 (N_4479,N_4150,N_4323);
nand U4480 (N_4480,N_4154,N_4378);
xnor U4481 (N_4481,N_4141,N_4110);
and U4482 (N_4482,N_4193,N_4189);
nand U4483 (N_4483,N_4174,N_4010);
and U4484 (N_4484,N_4124,N_4023);
nor U4485 (N_4485,N_4337,N_4258);
and U4486 (N_4486,N_4348,N_4152);
xnor U4487 (N_4487,N_4297,N_4088);
nand U4488 (N_4488,N_4396,N_4365);
nor U4489 (N_4489,N_4245,N_4233);
nor U4490 (N_4490,N_4188,N_4084);
nor U4491 (N_4491,N_4123,N_4222);
xor U4492 (N_4492,N_4362,N_4095);
nor U4493 (N_4493,N_4140,N_4126);
or U4494 (N_4494,N_4331,N_4302);
nand U4495 (N_4495,N_4044,N_4312);
nand U4496 (N_4496,N_4109,N_4071);
or U4497 (N_4497,N_4191,N_4380);
nor U4498 (N_4498,N_4165,N_4213);
nor U4499 (N_4499,N_4175,N_4389);
or U4500 (N_4500,N_4303,N_4014);
nand U4501 (N_4501,N_4157,N_4350);
xnor U4502 (N_4502,N_4146,N_4249);
nand U4503 (N_4503,N_4027,N_4037);
xor U4504 (N_4504,N_4091,N_4376);
nor U4505 (N_4505,N_4131,N_4315);
and U4506 (N_4506,N_4318,N_4224);
nand U4507 (N_4507,N_4298,N_4038);
nand U4508 (N_4508,N_4293,N_4215);
or U4509 (N_4509,N_4161,N_4016);
or U4510 (N_4510,N_4361,N_4022);
or U4511 (N_4511,N_4151,N_4013);
nand U4512 (N_4512,N_4006,N_4046);
nand U4513 (N_4513,N_4214,N_4169);
nand U4514 (N_4514,N_4226,N_4345);
nor U4515 (N_4515,N_4004,N_4096);
or U4516 (N_4516,N_4232,N_4138);
nor U4517 (N_4517,N_4349,N_4145);
nand U4518 (N_4518,N_4184,N_4211);
xnor U4519 (N_4519,N_4269,N_4058);
xor U4520 (N_4520,N_4282,N_4259);
or U4521 (N_4521,N_4144,N_4291);
nand U4522 (N_4522,N_4343,N_4209);
nor U4523 (N_4523,N_4075,N_4120);
and U4524 (N_4524,N_4336,N_4078);
xor U4525 (N_4525,N_4276,N_4286);
nor U4526 (N_4526,N_4142,N_4048);
xor U4527 (N_4527,N_4260,N_4053);
and U4528 (N_4528,N_4106,N_4254);
nor U4529 (N_4529,N_4153,N_4383);
and U4530 (N_4530,N_4072,N_4271);
or U4531 (N_4531,N_4242,N_4094);
nor U4532 (N_4532,N_4296,N_4121);
nor U4533 (N_4533,N_4114,N_4230);
or U4534 (N_4534,N_4167,N_4264);
nor U4535 (N_4535,N_4067,N_4041);
nor U4536 (N_4536,N_4118,N_4186);
nor U4537 (N_4537,N_4203,N_4310);
nand U4538 (N_4538,N_4170,N_4352);
xnor U4539 (N_4539,N_4066,N_4200);
nor U4540 (N_4540,N_4160,N_4108);
or U4541 (N_4541,N_4116,N_4054);
and U4542 (N_4542,N_4033,N_4247);
or U4543 (N_4543,N_4012,N_4081);
nand U4544 (N_4544,N_4357,N_4187);
xor U4545 (N_4545,N_4391,N_4241);
nor U4546 (N_4546,N_4060,N_4285);
xnor U4547 (N_4547,N_4292,N_4240);
and U4548 (N_4548,N_4219,N_4284);
xor U4549 (N_4549,N_4263,N_4375);
xnor U4550 (N_4550,N_4333,N_4079);
and U4551 (N_4551,N_4185,N_4238);
xnor U4552 (N_4552,N_4133,N_4274);
nand U4553 (N_4553,N_4225,N_4347);
nor U4554 (N_4554,N_4221,N_4055);
nor U4555 (N_4555,N_4082,N_4018);
and U4556 (N_4556,N_4332,N_4273);
nand U4557 (N_4557,N_4342,N_4340);
xor U4558 (N_4558,N_4287,N_4202);
nor U4559 (N_4559,N_4329,N_4227);
nand U4560 (N_4560,N_4237,N_4393);
and U4561 (N_4561,N_4172,N_4364);
nand U4562 (N_4562,N_4326,N_4134);
and U4563 (N_4563,N_4083,N_4316);
nor U4564 (N_4564,N_4388,N_4255);
nor U4565 (N_4565,N_4366,N_4001);
nor U4566 (N_4566,N_4268,N_4065);
or U4567 (N_4567,N_4278,N_4281);
xor U4568 (N_4568,N_4137,N_4308);
xor U4569 (N_4569,N_4279,N_4363);
nand U4570 (N_4570,N_4008,N_4205);
or U4571 (N_4571,N_4049,N_4311);
and U4572 (N_4572,N_4252,N_4057);
and U4573 (N_4573,N_4324,N_4322);
nand U4574 (N_4574,N_4338,N_4100);
nor U4575 (N_4575,N_4306,N_4177);
and U4576 (N_4576,N_4229,N_4373);
and U4577 (N_4577,N_4182,N_4369);
nor U4578 (N_4578,N_4250,N_4111);
xnor U4579 (N_4579,N_4089,N_4034);
or U4580 (N_4580,N_4097,N_4045);
nor U4581 (N_4581,N_4025,N_4327);
nand U4582 (N_4582,N_4166,N_4220);
xor U4583 (N_4583,N_4002,N_4335);
nor U4584 (N_4584,N_4085,N_4159);
nor U4585 (N_4585,N_4180,N_4218);
or U4586 (N_4586,N_4029,N_4003);
and U4587 (N_4587,N_4132,N_4162);
and U4588 (N_4588,N_4024,N_4294);
or U4589 (N_4589,N_4277,N_4248);
and U4590 (N_4590,N_4216,N_4122);
nor U4591 (N_4591,N_4090,N_4113);
xor U4592 (N_4592,N_4059,N_4021);
nand U4593 (N_4593,N_4171,N_4007);
and U4594 (N_4594,N_4107,N_4386);
and U4595 (N_4595,N_4017,N_4173);
xor U4596 (N_4596,N_4195,N_4115);
nand U4597 (N_4597,N_4313,N_4176);
nor U4598 (N_4598,N_4261,N_4370);
xor U4599 (N_4599,N_4005,N_4379);
and U4600 (N_4600,N_4036,N_4030);
nand U4601 (N_4601,N_4259,N_4175);
nor U4602 (N_4602,N_4299,N_4381);
and U4603 (N_4603,N_4275,N_4293);
xor U4604 (N_4604,N_4243,N_4384);
nand U4605 (N_4605,N_4257,N_4140);
nand U4606 (N_4606,N_4102,N_4179);
nand U4607 (N_4607,N_4172,N_4107);
or U4608 (N_4608,N_4016,N_4112);
nand U4609 (N_4609,N_4190,N_4187);
and U4610 (N_4610,N_4366,N_4279);
and U4611 (N_4611,N_4146,N_4078);
nor U4612 (N_4612,N_4002,N_4040);
nor U4613 (N_4613,N_4013,N_4074);
nand U4614 (N_4614,N_4297,N_4241);
or U4615 (N_4615,N_4144,N_4103);
or U4616 (N_4616,N_4152,N_4139);
nor U4617 (N_4617,N_4182,N_4391);
nand U4618 (N_4618,N_4119,N_4345);
or U4619 (N_4619,N_4095,N_4038);
or U4620 (N_4620,N_4279,N_4342);
nand U4621 (N_4621,N_4202,N_4277);
and U4622 (N_4622,N_4019,N_4131);
nand U4623 (N_4623,N_4266,N_4317);
and U4624 (N_4624,N_4025,N_4149);
xor U4625 (N_4625,N_4071,N_4124);
nor U4626 (N_4626,N_4208,N_4317);
or U4627 (N_4627,N_4171,N_4196);
xnor U4628 (N_4628,N_4080,N_4173);
xnor U4629 (N_4629,N_4173,N_4262);
nor U4630 (N_4630,N_4091,N_4121);
xnor U4631 (N_4631,N_4286,N_4018);
and U4632 (N_4632,N_4373,N_4027);
and U4633 (N_4633,N_4040,N_4033);
and U4634 (N_4634,N_4056,N_4072);
nand U4635 (N_4635,N_4127,N_4015);
nor U4636 (N_4636,N_4304,N_4084);
nand U4637 (N_4637,N_4169,N_4298);
or U4638 (N_4638,N_4055,N_4342);
or U4639 (N_4639,N_4395,N_4193);
or U4640 (N_4640,N_4357,N_4002);
or U4641 (N_4641,N_4335,N_4230);
and U4642 (N_4642,N_4133,N_4379);
xor U4643 (N_4643,N_4345,N_4198);
xnor U4644 (N_4644,N_4127,N_4331);
or U4645 (N_4645,N_4007,N_4169);
and U4646 (N_4646,N_4209,N_4394);
or U4647 (N_4647,N_4394,N_4103);
nand U4648 (N_4648,N_4223,N_4310);
nor U4649 (N_4649,N_4106,N_4136);
and U4650 (N_4650,N_4213,N_4217);
or U4651 (N_4651,N_4377,N_4079);
nand U4652 (N_4652,N_4372,N_4330);
xor U4653 (N_4653,N_4288,N_4101);
xor U4654 (N_4654,N_4347,N_4110);
or U4655 (N_4655,N_4037,N_4272);
nand U4656 (N_4656,N_4283,N_4341);
or U4657 (N_4657,N_4067,N_4317);
nor U4658 (N_4658,N_4084,N_4287);
xnor U4659 (N_4659,N_4221,N_4047);
and U4660 (N_4660,N_4034,N_4358);
and U4661 (N_4661,N_4106,N_4208);
nand U4662 (N_4662,N_4107,N_4259);
xnor U4663 (N_4663,N_4110,N_4225);
nor U4664 (N_4664,N_4147,N_4366);
nand U4665 (N_4665,N_4091,N_4347);
xnor U4666 (N_4666,N_4288,N_4112);
and U4667 (N_4667,N_4316,N_4278);
or U4668 (N_4668,N_4014,N_4285);
and U4669 (N_4669,N_4066,N_4208);
or U4670 (N_4670,N_4001,N_4250);
and U4671 (N_4671,N_4218,N_4020);
xor U4672 (N_4672,N_4320,N_4081);
xor U4673 (N_4673,N_4187,N_4353);
xor U4674 (N_4674,N_4183,N_4025);
nand U4675 (N_4675,N_4005,N_4245);
or U4676 (N_4676,N_4047,N_4375);
nand U4677 (N_4677,N_4142,N_4130);
nor U4678 (N_4678,N_4063,N_4009);
nor U4679 (N_4679,N_4265,N_4396);
or U4680 (N_4680,N_4083,N_4121);
or U4681 (N_4681,N_4339,N_4322);
nor U4682 (N_4682,N_4193,N_4296);
and U4683 (N_4683,N_4081,N_4365);
or U4684 (N_4684,N_4115,N_4340);
and U4685 (N_4685,N_4244,N_4154);
nor U4686 (N_4686,N_4174,N_4022);
xnor U4687 (N_4687,N_4127,N_4277);
nor U4688 (N_4688,N_4330,N_4238);
and U4689 (N_4689,N_4296,N_4145);
nor U4690 (N_4690,N_4084,N_4385);
or U4691 (N_4691,N_4247,N_4216);
nor U4692 (N_4692,N_4372,N_4296);
nor U4693 (N_4693,N_4156,N_4109);
or U4694 (N_4694,N_4004,N_4015);
or U4695 (N_4695,N_4364,N_4082);
and U4696 (N_4696,N_4308,N_4377);
nor U4697 (N_4697,N_4318,N_4233);
nor U4698 (N_4698,N_4257,N_4111);
and U4699 (N_4699,N_4019,N_4253);
nor U4700 (N_4700,N_4038,N_4224);
nand U4701 (N_4701,N_4323,N_4136);
and U4702 (N_4702,N_4375,N_4286);
xnor U4703 (N_4703,N_4325,N_4193);
nor U4704 (N_4704,N_4158,N_4221);
and U4705 (N_4705,N_4161,N_4210);
nor U4706 (N_4706,N_4348,N_4182);
and U4707 (N_4707,N_4011,N_4147);
nand U4708 (N_4708,N_4394,N_4154);
nor U4709 (N_4709,N_4058,N_4341);
or U4710 (N_4710,N_4105,N_4104);
or U4711 (N_4711,N_4196,N_4180);
or U4712 (N_4712,N_4295,N_4354);
nor U4713 (N_4713,N_4367,N_4322);
or U4714 (N_4714,N_4168,N_4257);
and U4715 (N_4715,N_4088,N_4171);
or U4716 (N_4716,N_4201,N_4346);
or U4717 (N_4717,N_4229,N_4092);
or U4718 (N_4718,N_4315,N_4390);
and U4719 (N_4719,N_4353,N_4021);
nor U4720 (N_4720,N_4116,N_4379);
or U4721 (N_4721,N_4376,N_4087);
and U4722 (N_4722,N_4398,N_4112);
nor U4723 (N_4723,N_4078,N_4091);
or U4724 (N_4724,N_4272,N_4227);
nand U4725 (N_4725,N_4140,N_4296);
nand U4726 (N_4726,N_4266,N_4230);
xor U4727 (N_4727,N_4033,N_4100);
nor U4728 (N_4728,N_4302,N_4137);
nand U4729 (N_4729,N_4228,N_4288);
xor U4730 (N_4730,N_4067,N_4006);
nor U4731 (N_4731,N_4033,N_4378);
nand U4732 (N_4732,N_4377,N_4333);
xnor U4733 (N_4733,N_4135,N_4226);
xor U4734 (N_4734,N_4322,N_4284);
or U4735 (N_4735,N_4391,N_4282);
or U4736 (N_4736,N_4075,N_4169);
nand U4737 (N_4737,N_4298,N_4164);
nor U4738 (N_4738,N_4302,N_4012);
or U4739 (N_4739,N_4355,N_4139);
xnor U4740 (N_4740,N_4051,N_4199);
nand U4741 (N_4741,N_4203,N_4225);
xnor U4742 (N_4742,N_4361,N_4279);
or U4743 (N_4743,N_4162,N_4365);
and U4744 (N_4744,N_4201,N_4327);
xor U4745 (N_4745,N_4142,N_4184);
nand U4746 (N_4746,N_4055,N_4385);
xor U4747 (N_4747,N_4177,N_4265);
nor U4748 (N_4748,N_4074,N_4342);
xnor U4749 (N_4749,N_4087,N_4068);
nor U4750 (N_4750,N_4307,N_4346);
nor U4751 (N_4751,N_4080,N_4180);
nor U4752 (N_4752,N_4337,N_4391);
and U4753 (N_4753,N_4134,N_4120);
nor U4754 (N_4754,N_4180,N_4117);
nor U4755 (N_4755,N_4154,N_4392);
nor U4756 (N_4756,N_4197,N_4261);
xor U4757 (N_4757,N_4118,N_4152);
or U4758 (N_4758,N_4223,N_4001);
nand U4759 (N_4759,N_4105,N_4269);
and U4760 (N_4760,N_4316,N_4272);
nor U4761 (N_4761,N_4060,N_4136);
or U4762 (N_4762,N_4354,N_4056);
nor U4763 (N_4763,N_4109,N_4310);
nor U4764 (N_4764,N_4257,N_4017);
xnor U4765 (N_4765,N_4209,N_4134);
xnor U4766 (N_4766,N_4095,N_4247);
and U4767 (N_4767,N_4033,N_4396);
and U4768 (N_4768,N_4240,N_4396);
nor U4769 (N_4769,N_4159,N_4237);
or U4770 (N_4770,N_4358,N_4035);
nor U4771 (N_4771,N_4331,N_4387);
nand U4772 (N_4772,N_4205,N_4206);
nor U4773 (N_4773,N_4011,N_4159);
nand U4774 (N_4774,N_4135,N_4225);
xor U4775 (N_4775,N_4127,N_4011);
nand U4776 (N_4776,N_4293,N_4222);
or U4777 (N_4777,N_4293,N_4250);
nand U4778 (N_4778,N_4107,N_4184);
nor U4779 (N_4779,N_4347,N_4211);
xor U4780 (N_4780,N_4150,N_4195);
and U4781 (N_4781,N_4368,N_4281);
or U4782 (N_4782,N_4006,N_4177);
nand U4783 (N_4783,N_4094,N_4122);
and U4784 (N_4784,N_4037,N_4004);
xor U4785 (N_4785,N_4226,N_4333);
xor U4786 (N_4786,N_4066,N_4344);
and U4787 (N_4787,N_4236,N_4372);
or U4788 (N_4788,N_4397,N_4309);
and U4789 (N_4789,N_4116,N_4040);
nor U4790 (N_4790,N_4018,N_4257);
nor U4791 (N_4791,N_4219,N_4084);
nor U4792 (N_4792,N_4324,N_4135);
xnor U4793 (N_4793,N_4205,N_4361);
nand U4794 (N_4794,N_4343,N_4022);
xor U4795 (N_4795,N_4004,N_4135);
nand U4796 (N_4796,N_4107,N_4313);
xor U4797 (N_4797,N_4161,N_4294);
and U4798 (N_4798,N_4289,N_4264);
nor U4799 (N_4799,N_4086,N_4324);
nor U4800 (N_4800,N_4699,N_4478);
or U4801 (N_4801,N_4643,N_4638);
xor U4802 (N_4802,N_4568,N_4526);
and U4803 (N_4803,N_4603,N_4572);
xnor U4804 (N_4804,N_4613,N_4671);
and U4805 (N_4805,N_4628,N_4466);
and U4806 (N_4806,N_4767,N_4609);
or U4807 (N_4807,N_4456,N_4665);
or U4808 (N_4808,N_4780,N_4556);
xor U4809 (N_4809,N_4471,N_4601);
or U4810 (N_4810,N_4632,N_4490);
nor U4811 (N_4811,N_4434,N_4579);
or U4812 (N_4812,N_4753,N_4681);
nor U4813 (N_4813,N_4407,N_4631);
nand U4814 (N_4814,N_4581,N_4797);
or U4815 (N_4815,N_4598,N_4687);
or U4816 (N_4816,N_4716,N_4626);
nor U4817 (N_4817,N_4500,N_4522);
xor U4818 (N_4818,N_4560,N_4589);
nand U4819 (N_4819,N_4439,N_4704);
nand U4820 (N_4820,N_4736,N_4454);
nor U4821 (N_4821,N_4515,N_4529);
and U4822 (N_4822,N_4552,N_4719);
or U4823 (N_4823,N_4667,N_4537);
nor U4824 (N_4824,N_4482,N_4587);
nor U4825 (N_4825,N_4702,N_4447);
xnor U4826 (N_4826,N_4777,N_4615);
nand U4827 (N_4827,N_4683,N_4532);
nor U4828 (N_4828,N_4745,N_4402);
nor U4829 (N_4829,N_4510,N_4694);
xor U4830 (N_4830,N_4645,N_4627);
nor U4831 (N_4831,N_4690,N_4472);
nor U4832 (N_4832,N_4504,N_4404);
nand U4833 (N_4833,N_4507,N_4420);
or U4834 (N_4834,N_4614,N_4610);
xor U4835 (N_4835,N_4557,N_4723);
or U4836 (N_4836,N_4755,N_4486);
or U4837 (N_4837,N_4569,N_4469);
xor U4838 (N_4838,N_4461,N_4750);
or U4839 (N_4839,N_4594,N_4503);
and U4840 (N_4840,N_4756,N_4752);
xor U4841 (N_4841,N_4652,N_4658);
and U4842 (N_4842,N_4676,N_4520);
nor U4843 (N_4843,N_4475,N_4588);
nand U4844 (N_4844,N_4430,N_4514);
or U4845 (N_4845,N_4567,N_4639);
nand U4846 (N_4846,N_4442,N_4707);
xnor U4847 (N_4847,N_4784,N_4661);
and U4848 (N_4848,N_4483,N_4734);
xnor U4849 (N_4849,N_4426,N_4709);
and U4850 (N_4850,N_4728,N_4495);
and U4851 (N_4851,N_4717,N_4738);
nand U4852 (N_4852,N_4769,N_4487);
nand U4853 (N_4853,N_4467,N_4494);
xor U4854 (N_4854,N_4437,N_4751);
xnor U4855 (N_4855,N_4692,N_4528);
or U4856 (N_4856,N_4758,N_4663);
nor U4857 (N_4857,N_4502,N_4629);
or U4858 (N_4858,N_4438,N_4521);
xor U4859 (N_4859,N_4549,N_4480);
nor U4860 (N_4860,N_4673,N_4539);
nor U4861 (N_4861,N_4477,N_4433);
nand U4862 (N_4862,N_4740,N_4536);
and U4863 (N_4863,N_4417,N_4550);
or U4864 (N_4864,N_4633,N_4771);
xor U4865 (N_4865,N_4449,N_4462);
or U4866 (N_4866,N_4443,N_4468);
nand U4867 (N_4867,N_4582,N_4696);
or U4868 (N_4868,N_4703,N_4782);
and U4869 (N_4869,N_4655,N_4656);
nor U4870 (N_4870,N_4714,N_4463);
and U4871 (N_4871,N_4508,N_4511);
and U4872 (N_4872,N_4600,N_4440);
and U4873 (N_4873,N_4516,N_4620);
or U4874 (N_4874,N_4781,N_4741);
or U4875 (N_4875,N_4799,N_4733);
and U4876 (N_4876,N_4698,N_4635);
nand U4877 (N_4877,N_4748,N_4489);
and U4878 (N_4878,N_4743,N_4700);
nor U4879 (N_4879,N_4617,N_4785);
nor U4880 (N_4880,N_4425,N_4649);
nand U4881 (N_4881,N_4608,N_4637);
nand U4882 (N_4882,N_4742,N_4474);
and U4883 (N_4883,N_4435,N_4406);
or U4884 (N_4884,N_4691,N_4686);
nor U4885 (N_4885,N_4693,N_4796);
xor U4886 (N_4886,N_4506,N_4411);
or U4887 (N_4887,N_4416,N_4530);
and U4888 (N_4888,N_4444,N_4583);
and U4889 (N_4889,N_4597,N_4773);
or U4890 (N_4890,N_4721,N_4565);
nand U4891 (N_4891,N_4695,N_4746);
and U4892 (N_4892,N_4445,N_4497);
or U4893 (N_4893,N_4762,N_4405);
nor U4894 (N_4894,N_4423,N_4496);
nor U4895 (N_4895,N_4547,N_4586);
nand U4896 (N_4896,N_4509,N_4523);
xor U4897 (N_4897,N_4418,N_4421);
or U4898 (N_4898,N_4559,N_4488);
xor U4899 (N_4899,N_4524,N_4760);
and U4900 (N_4900,N_4622,N_4754);
nor U4901 (N_4901,N_4621,N_4533);
nor U4902 (N_4902,N_4790,N_4476);
nand U4903 (N_4903,N_4720,N_4465);
nand U4904 (N_4904,N_4660,N_4545);
nor U4905 (N_4905,N_4473,N_4689);
and U4906 (N_4906,N_4562,N_4584);
nor U4907 (N_4907,N_4505,N_4527);
or U4908 (N_4908,N_4670,N_4606);
and U4909 (N_4909,N_4644,N_4427);
nand U4910 (N_4910,N_4446,N_4571);
xnor U4911 (N_4911,N_4759,N_4410);
xor U4912 (N_4912,N_4535,N_4675);
nand U4913 (N_4913,N_4401,N_4607);
and U4914 (N_4914,N_4595,N_4457);
or U4915 (N_4915,N_4715,N_4685);
xnor U4916 (N_4916,N_4677,N_4566);
nor U4917 (N_4917,N_4593,N_4450);
xor U4918 (N_4918,N_4554,N_4636);
xnor U4919 (N_4919,N_4747,N_4558);
and U4920 (N_4920,N_4611,N_4585);
or U4921 (N_4921,N_4612,N_4657);
xor U4922 (N_4922,N_4408,N_4664);
and U4923 (N_4923,N_4541,N_4599);
xnor U4924 (N_4924,N_4538,N_4436);
nand U4925 (N_4925,N_4464,N_4678);
xnor U4926 (N_4926,N_4737,N_4776);
and U4927 (N_4927,N_4653,N_4616);
nor U4928 (N_4928,N_4544,N_4574);
and U4929 (N_4929,N_4744,N_4732);
nand U4930 (N_4930,N_4540,N_4551);
nand U4931 (N_4931,N_4542,N_4592);
xor U4932 (N_4932,N_4646,N_4727);
and U4933 (N_4933,N_4739,N_4580);
and U4934 (N_4934,N_4662,N_4484);
xor U4935 (N_4935,N_4513,N_4789);
nand U4936 (N_4936,N_4798,N_4414);
nand U4937 (N_4937,N_4619,N_4431);
or U4938 (N_4938,N_4725,N_4648);
xor U4939 (N_4939,N_4518,N_4485);
nor U4940 (N_4940,N_4428,N_4705);
or U4941 (N_4941,N_4413,N_4548);
xnor U4942 (N_4942,N_4679,N_4577);
and U4943 (N_4943,N_4791,N_4666);
nand U4944 (N_4944,N_4697,N_4710);
xnor U4945 (N_4945,N_4458,N_4564);
or U4946 (N_4946,N_4561,N_4775);
nand U4947 (N_4947,N_4711,N_4712);
nor U4948 (N_4948,N_4674,N_4688);
or U4949 (N_4949,N_4630,N_4682);
and U4950 (N_4950,N_4591,N_4452);
nor U4951 (N_4951,N_4672,N_4757);
nor U4952 (N_4952,N_4546,N_4492);
xor U4953 (N_4953,N_4726,N_4422);
xnor U4954 (N_4954,N_4761,N_4731);
nor U4955 (N_4955,N_4735,N_4787);
nand U4956 (N_4956,N_4718,N_4634);
and U4957 (N_4957,N_4455,N_4543);
xor U4958 (N_4958,N_4793,N_4788);
and U4959 (N_4959,N_4459,N_4525);
or U4960 (N_4960,N_4623,N_4642);
nor U4961 (N_4961,N_4763,N_4400);
nand U4962 (N_4962,N_4481,N_4684);
and U4963 (N_4963,N_4650,N_4766);
nand U4964 (N_4964,N_4764,N_4654);
and U4965 (N_4965,N_4575,N_4774);
nor U4966 (N_4966,N_4708,N_4605);
nor U4967 (N_4967,N_4722,N_4596);
xnor U4968 (N_4968,N_4460,N_4792);
nor U4969 (N_4969,N_4625,N_4724);
nand U4970 (N_4970,N_4493,N_4429);
xor U4971 (N_4971,N_4453,N_4499);
xor U4972 (N_4972,N_4783,N_4659);
or U4973 (N_4973,N_4602,N_4519);
or U4974 (N_4974,N_4501,N_4498);
nand U4975 (N_4975,N_4534,N_4604);
nor U4976 (N_4976,N_4470,N_4409);
nor U4977 (N_4977,N_4641,N_4578);
nor U4978 (N_4978,N_4778,N_4618);
or U4979 (N_4979,N_4730,N_4770);
nand U4980 (N_4980,N_4651,N_4680);
and U4981 (N_4981,N_4669,N_4768);
or U4982 (N_4982,N_4412,N_4424);
nor U4983 (N_4983,N_4479,N_4576);
and U4984 (N_4984,N_4573,N_4794);
xnor U4985 (N_4985,N_4517,N_4512);
xnor U4986 (N_4986,N_4555,N_4729);
nor U4987 (N_4987,N_4772,N_4624);
nor U4988 (N_4988,N_4419,N_4765);
nand U4989 (N_4989,N_4590,N_4706);
and U4990 (N_4990,N_4668,N_4786);
and U4991 (N_4991,N_4448,N_4563);
nor U4992 (N_4992,N_4570,N_4779);
nand U4993 (N_4993,N_4403,N_4432);
nor U4994 (N_4994,N_4795,N_4531);
xnor U4995 (N_4995,N_4415,N_4553);
xor U4996 (N_4996,N_4451,N_4640);
nand U4997 (N_4997,N_4749,N_4701);
nand U4998 (N_4998,N_4491,N_4441);
or U4999 (N_4999,N_4647,N_4713);
nor U5000 (N_5000,N_4571,N_4556);
nor U5001 (N_5001,N_4581,N_4641);
or U5002 (N_5002,N_4722,N_4659);
or U5003 (N_5003,N_4668,N_4737);
nor U5004 (N_5004,N_4549,N_4794);
and U5005 (N_5005,N_4578,N_4792);
or U5006 (N_5006,N_4415,N_4563);
and U5007 (N_5007,N_4716,N_4635);
and U5008 (N_5008,N_4446,N_4729);
nand U5009 (N_5009,N_4766,N_4547);
and U5010 (N_5010,N_4686,N_4562);
nand U5011 (N_5011,N_4480,N_4492);
and U5012 (N_5012,N_4676,N_4619);
and U5013 (N_5013,N_4634,N_4643);
nor U5014 (N_5014,N_4775,N_4511);
nor U5015 (N_5015,N_4453,N_4670);
nand U5016 (N_5016,N_4512,N_4574);
nand U5017 (N_5017,N_4610,N_4452);
and U5018 (N_5018,N_4560,N_4584);
nor U5019 (N_5019,N_4732,N_4544);
xor U5020 (N_5020,N_4532,N_4684);
xor U5021 (N_5021,N_4693,N_4713);
xnor U5022 (N_5022,N_4460,N_4563);
nand U5023 (N_5023,N_4517,N_4578);
and U5024 (N_5024,N_4569,N_4750);
nand U5025 (N_5025,N_4581,N_4674);
and U5026 (N_5026,N_4665,N_4719);
xnor U5027 (N_5027,N_4433,N_4750);
or U5028 (N_5028,N_4508,N_4527);
nand U5029 (N_5029,N_4719,N_4690);
and U5030 (N_5030,N_4649,N_4682);
nand U5031 (N_5031,N_4434,N_4418);
and U5032 (N_5032,N_4447,N_4647);
and U5033 (N_5033,N_4622,N_4596);
or U5034 (N_5034,N_4472,N_4409);
nor U5035 (N_5035,N_4677,N_4771);
xor U5036 (N_5036,N_4797,N_4734);
xor U5037 (N_5037,N_4490,N_4651);
and U5038 (N_5038,N_4498,N_4414);
or U5039 (N_5039,N_4413,N_4795);
xnor U5040 (N_5040,N_4518,N_4665);
and U5041 (N_5041,N_4600,N_4497);
nor U5042 (N_5042,N_4493,N_4567);
and U5043 (N_5043,N_4651,N_4445);
xor U5044 (N_5044,N_4756,N_4774);
and U5045 (N_5045,N_4584,N_4771);
nor U5046 (N_5046,N_4466,N_4502);
or U5047 (N_5047,N_4726,N_4657);
or U5048 (N_5048,N_4755,N_4528);
nand U5049 (N_5049,N_4607,N_4568);
nand U5050 (N_5050,N_4454,N_4568);
nor U5051 (N_5051,N_4723,N_4669);
xor U5052 (N_5052,N_4509,N_4781);
and U5053 (N_5053,N_4699,N_4732);
nand U5054 (N_5054,N_4723,N_4788);
nand U5055 (N_5055,N_4672,N_4778);
xor U5056 (N_5056,N_4600,N_4565);
and U5057 (N_5057,N_4570,N_4664);
or U5058 (N_5058,N_4572,N_4670);
xnor U5059 (N_5059,N_4768,N_4661);
nor U5060 (N_5060,N_4558,N_4661);
nor U5061 (N_5061,N_4496,N_4796);
xnor U5062 (N_5062,N_4521,N_4473);
nor U5063 (N_5063,N_4729,N_4636);
xnor U5064 (N_5064,N_4526,N_4735);
or U5065 (N_5065,N_4618,N_4571);
or U5066 (N_5066,N_4659,N_4667);
xnor U5067 (N_5067,N_4459,N_4457);
nand U5068 (N_5068,N_4519,N_4505);
xnor U5069 (N_5069,N_4656,N_4414);
nand U5070 (N_5070,N_4689,N_4704);
xor U5071 (N_5071,N_4420,N_4631);
nor U5072 (N_5072,N_4459,N_4442);
or U5073 (N_5073,N_4436,N_4649);
and U5074 (N_5074,N_4795,N_4564);
nand U5075 (N_5075,N_4658,N_4584);
or U5076 (N_5076,N_4487,N_4776);
xnor U5077 (N_5077,N_4578,N_4745);
nor U5078 (N_5078,N_4443,N_4428);
nor U5079 (N_5079,N_4660,N_4589);
and U5080 (N_5080,N_4602,N_4740);
and U5081 (N_5081,N_4766,N_4759);
or U5082 (N_5082,N_4696,N_4553);
or U5083 (N_5083,N_4465,N_4681);
xnor U5084 (N_5084,N_4510,N_4490);
nor U5085 (N_5085,N_4483,N_4670);
nor U5086 (N_5086,N_4445,N_4553);
or U5087 (N_5087,N_4528,N_4479);
or U5088 (N_5088,N_4788,N_4639);
nand U5089 (N_5089,N_4479,N_4670);
xor U5090 (N_5090,N_4712,N_4490);
xnor U5091 (N_5091,N_4720,N_4754);
nor U5092 (N_5092,N_4750,N_4747);
or U5093 (N_5093,N_4673,N_4442);
or U5094 (N_5094,N_4578,N_4779);
and U5095 (N_5095,N_4670,N_4409);
or U5096 (N_5096,N_4693,N_4624);
nor U5097 (N_5097,N_4536,N_4635);
or U5098 (N_5098,N_4712,N_4780);
and U5099 (N_5099,N_4552,N_4611);
xor U5100 (N_5100,N_4788,N_4632);
or U5101 (N_5101,N_4734,N_4414);
nand U5102 (N_5102,N_4668,N_4626);
nor U5103 (N_5103,N_4536,N_4748);
and U5104 (N_5104,N_4799,N_4797);
nand U5105 (N_5105,N_4757,N_4596);
nor U5106 (N_5106,N_4484,N_4791);
xnor U5107 (N_5107,N_4447,N_4617);
nand U5108 (N_5108,N_4468,N_4663);
nor U5109 (N_5109,N_4786,N_4496);
nand U5110 (N_5110,N_4778,N_4751);
nand U5111 (N_5111,N_4439,N_4698);
nand U5112 (N_5112,N_4614,N_4676);
and U5113 (N_5113,N_4671,N_4734);
nor U5114 (N_5114,N_4406,N_4721);
or U5115 (N_5115,N_4615,N_4741);
and U5116 (N_5116,N_4619,N_4760);
nand U5117 (N_5117,N_4603,N_4567);
xnor U5118 (N_5118,N_4402,N_4587);
nand U5119 (N_5119,N_4432,N_4696);
xor U5120 (N_5120,N_4616,N_4757);
and U5121 (N_5121,N_4527,N_4701);
or U5122 (N_5122,N_4544,N_4581);
or U5123 (N_5123,N_4420,N_4707);
nor U5124 (N_5124,N_4749,N_4420);
nand U5125 (N_5125,N_4699,N_4681);
nor U5126 (N_5126,N_4606,N_4576);
xnor U5127 (N_5127,N_4454,N_4505);
xnor U5128 (N_5128,N_4516,N_4517);
nor U5129 (N_5129,N_4452,N_4778);
and U5130 (N_5130,N_4434,N_4669);
nor U5131 (N_5131,N_4429,N_4586);
nor U5132 (N_5132,N_4453,N_4647);
nand U5133 (N_5133,N_4778,N_4568);
nor U5134 (N_5134,N_4429,N_4729);
nor U5135 (N_5135,N_4516,N_4667);
or U5136 (N_5136,N_4730,N_4511);
or U5137 (N_5137,N_4602,N_4495);
nor U5138 (N_5138,N_4612,N_4469);
or U5139 (N_5139,N_4562,N_4542);
xor U5140 (N_5140,N_4524,N_4646);
nand U5141 (N_5141,N_4484,N_4680);
xor U5142 (N_5142,N_4627,N_4672);
nor U5143 (N_5143,N_4633,N_4657);
nand U5144 (N_5144,N_4772,N_4716);
nor U5145 (N_5145,N_4460,N_4644);
nand U5146 (N_5146,N_4439,N_4515);
nor U5147 (N_5147,N_4442,N_4760);
xnor U5148 (N_5148,N_4743,N_4632);
and U5149 (N_5149,N_4777,N_4549);
xnor U5150 (N_5150,N_4787,N_4785);
and U5151 (N_5151,N_4450,N_4527);
or U5152 (N_5152,N_4731,N_4740);
or U5153 (N_5153,N_4634,N_4598);
nor U5154 (N_5154,N_4550,N_4732);
or U5155 (N_5155,N_4609,N_4557);
or U5156 (N_5156,N_4616,N_4625);
xnor U5157 (N_5157,N_4555,N_4770);
or U5158 (N_5158,N_4433,N_4616);
or U5159 (N_5159,N_4586,N_4575);
nand U5160 (N_5160,N_4437,N_4586);
nand U5161 (N_5161,N_4594,N_4640);
nor U5162 (N_5162,N_4624,N_4612);
and U5163 (N_5163,N_4699,N_4566);
or U5164 (N_5164,N_4656,N_4458);
nand U5165 (N_5165,N_4597,N_4513);
or U5166 (N_5166,N_4504,N_4554);
and U5167 (N_5167,N_4714,N_4544);
xnor U5168 (N_5168,N_4412,N_4586);
or U5169 (N_5169,N_4534,N_4782);
and U5170 (N_5170,N_4664,N_4462);
nor U5171 (N_5171,N_4498,N_4434);
nand U5172 (N_5172,N_4483,N_4411);
and U5173 (N_5173,N_4779,N_4410);
nor U5174 (N_5174,N_4739,N_4412);
or U5175 (N_5175,N_4505,N_4534);
and U5176 (N_5176,N_4441,N_4722);
or U5177 (N_5177,N_4784,N_4562);
nor U5178 (N_5178,N_4623,N_4501);
nand U5179 (N_5179,N_4685,N_4408);
xnor U5180 (N_5180,N_4428,N_4759);
xnor U5181 (N_5181,N_4510,N_4664);
nor U5182 (N_5182,N_4550,N_4491);
and U5183 (N_5183,N_4642,N_4755);
or U5184 (N_5184,N_4679,N_4777);
nor U5185 (N_5185,N_4534,N_4645);
and U5186 (N_5186,N_4561,N_4755);
nand U5187 (N_5187,N_4639,N_4779);
or U5188 (N_5188,N_4694,N_4454);
or U5189 (N_5189,N_4766,N_4549);
and U5190 (N_5190,N_4783,N_4668);
nand U5191 (N_5191,N_4714,N_4472);
nor U5192 (N_5192,N_4458,N_4624);
xor U5193 (N_5193,N_4754,N_4440);
nand U5194 (N_5194,N_4659,N_4636);
or U5195 (N_5195,N_4772,N_4509);
xnor U5196 (N_5196,N_4498,N_4420);
nand U5197 (N_5197,N_4637,N_4584);
nor U5198 (N_5198,N_4511,N_4525);
xnor U5199 (N_5199,N_4743,N_4414);
nor U5200 (N_5200,N_4800,N_4815);
nand U5201 (N_5201,N_4884,N_5115);
or U5202 (N_5202,N_5107,N_5082);
nor U5203 (N_5203,N_4877,N_4934);
or U5204 (N_5204,N_5187,N_4924);
nand U5205 (N_5205,N_4976,N_5152);
nor U5206 (N_5206,N_5046,N_5135);
xnor U5207 (N_5207,N_5028,N_4827);
xor U5208 (N_5208,N_5188,N_4835);
or U5209 (N_5209,N_5105,N_4834);
xor U5210 (N_5210,N_5084,N_5104);
xor U5211 (N_5211,N_5142,N_5074);
or U5212 (N_5212,N_4999,N_5090);
and U5213 (N_5213,N_5038,N_5015);
and U5214 (N_5214,N_4845,N_5042);
xor U5215 (N_5215,N_4975,N_5000);
xor U5216 (N_5216,N_5175,N_5009);
nor U5217 (N_5217,N_5071,N_5075);
nor U5218 (N_5218,N_4969,N_5058);
nand U5219 (N_5219,N_5167,N_5100);
xor U5220 (N_5220,N_5036,N_5010);
nor U5221 (N_5221,N_4919,N_4892);
and U5222 (N_5222,N_4961,N_4988);
and U5223 (N_5223,N_5035,N_4809);
xor U5224 (N_5224,N_4942,N_4900);
and U5225 (N_5225,N_4850,N_5013);
nand U5226 (N_5226,N_5153,N_5192);
nor U5227 (N_5227,N_4876,N_5102);
nand U5228 (N_5228,N_4825,N_4996);
xor U5229 (N_5229,N_5161,N_4816);
nor U5230 (N_5230,N_4808,N_4965);
nand U5231 (N_5231,N_5180,N_5016);
nor U5232 (N_5232,N_5120,N_5076);
nand U5233 (N_5233,N_4891,N_4926);
or U5234 (N_5234,N_5198,N_4925);
and U5235 (N_5235,N_4865,N_5119);
xnor U5236 (N_5236,N_5131,N_4970);
xor U5237 (N_5237,N_5037,N_4953);
nand U5238 (N_5238,N_4862,N_4908);
xnor U5239 (N_5239,N_4978,N_5041);
and U5240 (N_5240,N_5024,N_4803);
nor U5241 (N_5241,N_4833,N_4917);
nand U5242 (N_5242,N_5149,N_5044);
xor U5243 (N_5243,N_4895,N_5110);
nand U5244 (N_5244,N_5083,N_4853);
nand U5245 (N_5245,N_4826,N_4915);
nand U5246 (N_5246,N_5116,N_5048);
or U5247 (N_5247,N_4894,N_5095);
nor U5248 (N_5248,N_4913,N_5091);
and U5249 (N_5249,N_5061,N_4974);
nor U5250 (N_5250,N_5113,N_4986);
and U5251 (N_5251,N_5164,N_4812);
xor U5252 (N_5252,N_4998,N_5136);
or U5253 (N_5253,N_5086,N_4859);
nor U5254 (N_5254,N_4964,N_5002);
nor U5255 (N_5255,N_4931,N_5025);
xor U5256 (N_5256,N_4967,N_4977);
nor U5257 (N_5257,N_5063,N_4874);
nand U5258 (N_5258,N_5108,N_5027);
and U5259 (N_5259,N_4904,N_4860);
xor U5260 (N_5260,N_4947,N_5055);
nor U5261 (N_5261,N_4899,N_4930);
or U5262 (N_5262,N_5172,N_5125);
nor U5263 (N_5263,N_4863,N_5069);
or U5264 (N_5264,N_5080,N_5132);
nor U5265 (N_5265,N_5026,N_4937);
nor U5266 (N_5266,N_5174,N_5052);
or U5267 (N_5267,N_5033,N_4940);
nand U5268 (N_5268,N_5158,N_5183);
or U5269 (N_5269,N_4918,N_4910);
or U5270 (N_5270,N_4866,N_4855);
nor U5271 (N_5271,N_4807,N_5007);
nand U5272 (N_5272,N_5062,N_5017);
xnor U5273 (N_5273,N_5134,N_5039);
or U5274 (N_5274,N_4992,N_5157);
and U5275 (N_5275,N_4868,N_4839);
and U5276 (N_5276,N_4932,N_5138);
nand U5277 (N_5277,N_5151,N_4994);
nand U5278 (N_5278,N_5068,N_5099);
nand U5279 (N_5279,N_5056,N_5098);
nand U5280 (N_5280,N_5154,N_4843);
and U5281 (N_5281,N_5111,N_5001);
nand U5282 (N_5282,N_5106,N_4869);
nand U5283 (N_5283,N_5176,N_4841);
nand U5284 (N_5284,N_4979,N_4813);
xor U5285 (N_5285,N_5032,N_5128);
nand U5286 (N_5286,N_5143,N_4956);
xnor U5287 (N_5287,N_4968,N_5011);
nor U5288 (N_5288,N_4963,N_4840);
or U5289 (N_5289,N_4804,N_5191);
or U5290 (N_5290,N_5040,N_4893);
xor U5291 (N_5291,N_5092,N_4820);
nor U5292 (N_5292,N_4989,N_4844);
nor U5293 (N_5293,N_5023,N_5144);
and U5294 (N_5294,N_5081,N_4801);
nand U5295 (N_5295,N_5182,N_5127);
or U5296 (N_5296,N_5112,N_5078);
or U5297 (N_5297,N_5031,N_5193);
and U5298 (N_5298,N_5146,N_5114);
or U5299 (N_5299,N_5005,N_4888);
nand U5300 (N_5300,N_4907,N_5148);
and U5301 (N_5301,N_5050,N_4973);
xor U5302 (N_5302,N_4902,N_4885);
nand U5303 (N_5303,N_5072,N_4896);
and U5304 (N_5304,N_4838,N_4985);
nand U5305 (N_5305,N_5170,N_4922);
or U5306 (N_5306,N_4921,N_4858);
and U5307 (N_5307,N_4912,N_5124);
nor U5308 (N_5308,N_4945,N_5054);
nand U5309 (N_5309,N_5189,N_4957);
and U5310 (N_5310,N_4819,N_5147);
nor U5311 (N_5311,N_5159,N_4870);
or U5312 (N_5312,N_5029,N_5059);
or U5313 (N_5313,N_4948,N_5077);
xor U5314 (N_5314,N_4861,N_5129);
xnor U5315 (N_5315,N_5034,N_5030);
nor U5316 (N_5316,N_5049,N_4920);
nor U5317 (N_5317,N_4901,N_4943);
nor U5318 (N_5318,N_5155,N_5117);
or U5319 (N_5319,N_4854,N_4890);
nand U5320 (N_5320,N_4911,N_5003);
nand U5321 (N_5321,N_4802,N_4950);
or U5322 (N_5322,N_4806,N_5185);
nand U5323 (N_5323,N_4822,N_5150);
and U5324 (N_5324,N_5051,N_4887);
and U5325 (N_5325,N_5012,N_5165);
and U5326 (N_5326,N_5178,N_4847);
nor U5327 (N_5327,N_5181,N_4856);
nor U5328 (N_5328,N_5047,N_4875);
or U5329 (N_5329,N_4980,N_5139);
nor U5330 (N_5330,N_4829,N_4849);
xnor U5331 (N_5331,N_4981,N_4949);
nand U5332 (N_5332,N_4846,N_4960);
and U5333 (N_5333,N_5121,N_4883);
xor U5334 (N_5334,N_4929,N_4886);
or U5335 (N_5335,N_4878,N_5194);
and U5336 (N_5336,N_5085,N_4864);
and U5337 (N_5337,N_5168,N_4962);
nand U5338 (N_5338,N_4941,N_4928);
xor U5339 (N_5339,N_4909,N_5014);
or U5340 (N_5340,N_5073,N_5123);
and U5341 (N_5341,N_4905,N_5089);
or U5342 (N_5342,N_5019,N_4982);
and U5343 (N_5343,N_5197,N_4879);
nand U5344 (N_5344,N_5088,N_5079);
nor U5345 (N_5345,N_5103,N_5021);
nor U5346 (N_5346,N_5130,N_5087);
or U5347 (N_5347,N_5190,N_4837);
nand U5348 (N_5348,N_4971,N_5163);
nand U5349 (N_5349,N_5020,N_4958);
xor U5350 (N_5350,N_4873,N_5140);
nand U5351 (N_5351,N_5196,N_4810);
or U5352 (N_5352,N_5004,N_5067);
nor U5353 (N_5353,N_4898,N_4811);
or U5354 (N_5354,N_4991,N_5070);
nand U5355 (N_5355,N_4954,N_5122);
nand U5356 (N_5356,N_4882,N_4935);
xnor U5357 (N_5357,N_4851,N_5018);
nor U5358 (N_5358,N_5065,N_4990);
nand U5359 (N_5359,N_5126,N_5057);
nand U5360 (N_5360,N_4944,N_5141);
and U5361 (N_5361,N_4871,N_4987);
nand U5362 (N_5362,N_4872,N_5160);
and U5363 (N_5363,N_4916,N_5043);
and U5364 (N_5364,N_4952,N_5064);
xnor U5365 (N_5365,N_4842,N_4983);
xnor U5366 (N_5366,N_4933,N_4848);
and U5367 (N_5367,N_4972,N_4821);
nor U5368 (N_5368,N_4823,N_5184);
xor U5369 (N_5369,N_4881,N_4951);
nor U5370 (N_5370,N_4830,N_4997);
xnor U5371 (N_5371,N_4836,N_4889);
nor U5372 (N_5372,N_5162,N_5145);
and U5373 (N_5373,N_4805,N_4832);
nor U5374 (N_5374,N_5060,N_5008);
xor U5375 (N_5375,N_5177,N_4828);
nand U5376 (N_5376,N_5093,N_4984);
nand U5377 (N_5377,N_5109,N_4959);
nand U5378 (N_5378,N_4995,N_4936);
xor U5379 (N_5379,N_4993,N_5097);
or U5380 (N_5380,N_5171,N_4831);
or U5381 (N_5381,N_5118,N_5094);
nor U5382 (N_5382,N_5022,N_4938);
nor U5383 (N_5383,N_4817,N_4897);
and U5384 (N_5384,N_4903,N_5006);
and U5385 (N_5385,N_5156,N_5101);
or U5386 (N_5386,N_4946,N_5186);
or U5387 (N_5387,N_4867,N_4966);
xnor U5388 (N_5388,N_4927,N_4814);
and U5389 (N_5389,N_5133,N_4824);
or U5390 (N_5390,N_4857,N_5179);
and U5391 (N_5391,N_5137,N_4923);
nand U5392 (N_5392,N_4852,N_5199);
nor U5393 (N_5393,N_4880,N_5166);
nand U5394 (N_5394,N_5169,N_5066);
nand U5395 (N_5395,N_5173,N_4955);
nand U5396 (N_5396,N_4914,N_4939);
xnor U5397 (N_5397,N_4818,N_5096);
nand U5398 (N_5398,N_5045,N_5053);
nand U5399 (N_5399,N_5195,N_4906);
xor U5400 (N_5400,N_4800,N_5161);
or U5401 (N_5401,N_4814,N_4830);
xnor U5402 (N_5402,N_4954,N_4806);
xor U5403 (N_5403,N_4969,N_5066);
nor U5404 (N_5404,N_4814,N_5111);
nand U5405 (N_5405,N_5173,N_5176);
or U5406 (N_5406,N_4966,N_5096);
or U5407 (N_5407,N_4859,N_5040);
xnor U5408 (N_5408,N_5061,N_4911);
xor U5409 (N_5409,N_5144,N_4841);
nor U5410 (N_5410,N_4880,N_4939);
and U5411 (N_5411,N_5006,N_5101);
and U5412 (N_5412,N_4950,N_4852);
and U5413 (N_5413,N_5048,N_5023);
xor U5414 (N_5414,N_4912,N_4813);
xor U5415 (N_5415,N_4918,N_5073);
xnor U5416 (N_5416,N_5039,N_4815);
and U5417 (N_5417,N_5089,N_4976);
and U5418 (N_5418,N_4902,N_4803);
and U5419 (N_5419,N_4994,N_5164);
xnor U5420 (N_5420,N_4987,N_4841);
nand U5421 (N_5421,N_4905,N_4965);
xnor U5422 (N_5422,N_5130,N_5179);
xnor U5423 (N_5423,N_5145,N_5136);
or U5424 (N_5424,N_4806,N_4884);
nor U5425 (N_5425,N_4825,N_4853);
nand U5426 (N_5426,N_4920,N_5037);
or U5427 (N_5427,N_4826,N_5035);
or U5428 (N_5428,N_4840,N_4964);
xnor U5429 (N_5429,N_5114,N_4804);
or U5430 (N_5430,N_4849,N_5033);
or U5431 (N_5431,N_4839,N_5082);
and U5432 (N_5432,N_4944,N_4855);
and U5433 (N_5433,N_5012,N_4954);
nor U5434 (N_5434,N_5050,N_4933);
nand U5435 (N_5435,N_5011,N_4926);
or U5436 (N_5436,N_4896,N_4800);
or U5437 (N_5437,N_5149,N_4968);
or U5438 (N_5438,N_4951,N_4838);
xnor U5439 (N_5439,N_5027,N_4987);
nor U5440 (N_5440,N_4970,N_4813);
and U5441 (N_5441,N_5148,N_5159);
or U5442 (N_5442,N_5027,N_4889);
xnor U5443 (N_5443,N_4949,N_4900);
nor U5444 (N_5444,N_5145,N_5196);
xnor U5445 (N_5445,N_4857,N_5013);
or U5446 (N_5446,N_5060,N_4831);
or U5447 (N_5447,N_4814,N_4870);
or U5448 (N_5448,N_4960,N_4925);
xnor U5449 (N_5449,N_4930,N_5011);
nand U5450 (N_5450,N_5008,N_4905);
xnor U5451 (N_5451,N_5160,N_5154);
nand U5452 (N_5452,N_5110,N_4841);
or U5453 (N_5453,N_4884,N_4818);
xnor U5454 (N_5454,N_4829,N_4966);
or U5455 (N_5455,N_4955,N_5099);
nand U5456 (N_5456,N_5030,N_5156);
and U5457 (N_5457,N_4958,N_4852);
nor U5458 (N_5458,N_4965,N_4955);
or U5459 (N_5459,N_5140,N_5095);
or U5460 (N_5460,N_5150,N_5000);
xor U5461 (N_5461,N_4802,N_5001);
or U5462 (N_5462,N_5187,N_5168);
and U5463 (N_5463,N_5138,N_5017);
nand U5464 (N_5464,N_4878,N_5165);
and U5465 (N_5465,N_4928,N_4930);
xor U5466 (N_5466,N_5179,N_4910);
and U5467 (N_5467,N_5121,N_5013);
nand U5468 (N_5468,N_4953,N_5025);
nand U5469 (N_5469,N_4942,N_5107);
and U5470 (N_5470,N_5031,N_5156);
or U5471 (N_5471,N_5106,N_5027);
and U5472 (N_5472,N_4844,N_5111);
and U5473 (N_5473,N_5056,N_4973);
xnor U5474 (N_5474,N_5085,N_5011);
and U5475 (N_5475,N_4850,N_5037);
xor U5476 (N_5476,N_4819,N_5143);
nand U5477 (N_5477,N_5170,N_4936);
and U5478 (N_5478,N_5006,N_5156);
or U5479 (N_5479,N_5044,N_4818);
xor U5480 (N_5480,N_5090,N_4854);
or U5481 (N_5481,N_4987,N_5063);
nand U5482 (N_5482,N_5000,N_4857);
nand U5483 (N_5483,N_4941,N_4890);
xnor U5484 (N_5484,N_4921,N_5036);
nand U5485 (N_5485,N_5097,N_4958);
nand U5486 (N_5486,N_4937,N_4885);
xor U5487 (N_5487,N_4965,N_4999);
nand U5488 (N_5488,N_4922,N_4874);
nor U5489 (N_5489,N_5017,N_4956);
and U5490 (N_5490,N_4975,N_4848);
and U5491 (N_5491,N_5104,N_4950);
nand U5492 (N_5492,N_4886,N_5161);
nand U5493 (N_5493,N_5159,N_5057);
nand U5494 (N_5494,N_4883,N_5040);
or U5495 (N_5495,N_5143,N_5155);
or U5496 (N_5496,N_5025,N_5037);
nand U5497 (N_5497,N_5077,N_4840);
nor U5498 (N_5498,N_5074,N_5060);
and U5499 (N_5499,N_4863,N_5155);
nand U5500 (N_5500,N_4857,N_4803);
nor U5501 (N_5501,N_4865,N_4920);
and U5502 (N_5502,N_5035,N_5075);
and U5503 (N_5503,N_5137,N_4805);
xnor U5504 (N_5504,N_5154,N_5173);
and U5505 (N_5505,N_4931,N_4804);
xor U5506 (N_5506,N_5158,N_4955);
xnor U5507 (N_5507,N_5062,N_4966);
nor U5508 (N_5508,N_5057,N_5153);
and U5509 (N_5509,N_5170,N_5102);
nor U5510 (N_5510,N_5094,N_5147);
and U5511 (N_5511,N_4944,N_5042);
or U5512 (N_5512,N_5189,N_4829);
and U5513 (N_5513,N_5076,N_5124);
xor U5514 (N_5514,N_4970,N_5169);
nor U5515 (N_5515,N_5115,N_4998);
nor U5516 (N_5516,N_5010,N_5061);
nor U5517 (N_5517,N_4924,N_4852);
and U5518 (N_5518,N_4965,N_5055);
or U5519 (N_5519,N_4909,N_4861);
or U5520 (N_5520,N_4974,N_4911);
nand U5521 (N_5521,N_5181,N_4874);
and U5522 (N_5522,N_4924,N_5112);
nor U5523 (N_5523,N_5117,N_5126);
nor U5524 (N_5524,N_4820,N_5038);
xnor U5525 (N_5525,N_4866,N_4899);
nand U5526 (N_5526,N_5121,N_4998);
or U5527 (N_5527,N_5020,N_5156);
nor U5528 (N_5528,N_4832,N_5024);
nand U5529 (N_5529,N_5041,N_4839);
nand U5530 (N_5530,N_4935,N_4811);
or U5531 (N_5531,N_4922,N_4971);
nor U5532 (N_5532,N_5188,N_4854);
and U5533 (N_5533,N_5063,N_5052);
nor U5534 (N_5534,N_5193,N_4940);
or U5535 (N_5535,N_5197,N_4960);
or U5536 (N_5536,N_4886,N_4813);
or U5537 (N_5537,N_4914,N_4937);
or U5538 (N_5538,N_5172,N_4946);
and U5539 (N_5539,N_5011,N_5069);
nand U5540 (N_5540,N_5109,N_5191);
and U5541 (N_5541,N_5016,N_5149);
xor U5542 (N_5542,N_5120,N_5106);
xnor U5543 (N_5543,N_4805,N_5085);
nor U5544 (N_5544,N_4867,N_4929);
xnor U5545 (N_5545,N_5173,N_5187);
nor U5546 (N_5546,N_5114,N_4923);
or U5547 (N_5547,N_5196,N_4838);
nor U5548 (N_5548,N_5118,N_5108);
nor U5549 (N_5549,N_5094,N_4974);
xor U5550 (N_5550,N_4815,N_5086);
nand U5551 (N_5551,N_5092,N_5128);
nand U5552 (N_5552,N_4902,N_5160);
nand U5553 (N_5553,N_4899,N_4814);
and U5554 (N_5554,N_4866,N_5139);
nor U5555 (N_5555,N_4987,N_4935);
nand U5556 (N_5556,N_4919,N_4862);
nor U5557 (N_5557,N_5090,N_4960);
xnor U5558 (N_5558,N_4824,N_4839);
and U5559 (N_5559,N_5096,N_5005);
or U5560 (N_5560,N_5167,N_4844);
and U5561 (N_5561,N_4828,N_5119);
nand U5562 (N_5562,N_4957,N_4800);
nor U5563 (N_5563,N_4845,N_4918);
xnor U5564 (N_5564,N_5090,N_4880);
nand U5565 (N_5565,N_4887,N_5116);
xnor U5566 (N_5566,N_5027,N_5030);
and U5567 (N_5567,N_4858,N_4800);
or U5568 (N_5568,N_5094,N_4801);
nor U5569 (N_5569,N_5004,N_5028);
nor U5570 (N_5570,N_5187,N_5030);
nor U5571 (N_5571,N_5116,N_4823);
nor U5572 (N_5572,N_4819,N_5094);
xnor U5573 (N_5573,N_5170,N_4921);
or U5574 (N_5574,N_4930,N_4853);
or U5575 (N_5575,N_4843,N_4990);
and U5576 (N_5576,N_5109,N_4808);
or U5577 (N_5577,N_5180,N_4829);
and U5578 (N_5578,N_4827,N_4889);
nand U5579 (N_5579,N_4817,N_4816);
or U5580 (N_5580,N_4904,N_4848);
xnor U5581 (N_5581,N_4889,N_4846);
xor U5582 (N_5582,N_4846,N_4927);
and U5583 (N_5583,N_5097,N_5168);
nand U5584 (N_5584,N_4864,N_5147);
xnor U5585 (N_5585,N_4903,N_4997);
and U5586 (N_5586,N_5044,N_5107);
or U5587 (N_5587,N_4893,N_4831);
xor U5588 (N_5588,N_4858,N_4848);
or U5589 (N_5589,N_5038,N_5095);
or U5590 (N_5590,N_5193,N_4814);
and U5591 (N_5591,N_5172,N_5192);
or U5592 (N_5592,N_4862,N_5079);
or U5593 (N_5593,N_5005,N_4860);
or U5594 (N_5594,N_5127,N_5174);
nand U5595 (N_5595,N_4936,N_4992);
or U5596 (N_5596,N_5171,N_5189);
nor U5597 (N_5597,N_5134,N_5136);
xor U5598 (N_5598,N_4914,N_4996);
nand U5599 (N_5599,N_4868,N_4842);
nand U5600 (N_5600,N_5558,N_5289);
nand U5601 (N_5601,N_5354,N_5459);
nand U5602 (N_5602,N_5335,N_5272);
xnor U5603 (N_5603,N_5291,N_5583);
xnor U5604 (N_5604,N_5487,N_5202);
nor U5605 (N_5605,N_5415,N_5475);
and U5606 (N_5606,N_5267,N_5318);
nor U5607 (N_5607,N_5217,N_5446);
xor U5608 (N_5608,N_5581,N_5441);
or U5609 (N_5609,N_5286,N_5419);
xor U5610 (N_5610,N_5397,N_5316);
and U5611 (N_5611,N_5392,N_5219);
nand U5612 (N_5612,N_5206,N_5511);
nand U5613 (N_5613,N_5435,N_5311);
nor U5614 (N_5614,N_5274,N_5270);
xor U5615 (N_5615,N_5205,N_5571);
and U5616 (N_5616,N_5405,N_5433);
nand U5617 (N_5617,N_5361,N_5221);
nor U5618 (N_5618,N_5516,N_5338);
nand U5619 (N_5619,N_5545,N_5216);
nand U5620 (N_5620,N_5233,N_5380);
and U5621 (N_5621,N_5313,N_5478);
xnor U5622 (N_5622,N_5372,N_5554);
nor U5623 (N_5623,N_5207,N_5237);
nand U5624 (N_5624,N_5301,N_5300);
and U5625 (N_5625,N_5265,N_5327);
and U5626 (N_5626,N_5279,N_5442);
nand U5627 (N_5627,N_5473,N_5412);
nand U5628 (N_5628,N_5462,N_5406);
xor U5629 (N_5629,N_5238,N_5533);
nand U5630 (N_5630,N_5468,N_5578);
nand U5631 (N_5631,N_5251,N_5243);
and U5632 (N_5632,N_5440,N_5388);
and U5633 (N_5633,N_5296,N_5323);
nor U5634 (N_5634,N_5501,N_5261);
nand U5635 (N_5635,N_5496,N_5491);
or U5636 (N_5636,N_5359,N_5390);
and U5637 (N_5637,N_5551,N_5257);
and U5638 (N_5638,N_5467,N_5394);
xnor U5639 (N_5639,N_5585,N_5402);
nor U5640 (N_5640,N_5203,N_5236);
and U5641 (N_5641,N_5444,N_5263);
xnor U5642 (N_5642,N_5593,N_5574);
and U5643 (N_5643,N_5465,N_5396);
or U5644 (N_5644,N_5333,N_5505);
nor U5645 (N_5645,N_5503,N_5398);
xnor U5646 (N_5646,N_5555,N_5549);
or U5647 (N_5647,N_5234,N_5352);
xor U5648 (N_5648,N_5517,N_5422);
nand U5649 (N_5649,N_5411,N_5413);
and U5650 (N_5650,N_5497,N_5370);
nor U5651 (N_5651,N_5480,N_5218);
and U5652 (N_5652,N_5563,N_5389);
and U5653 (N_5653,N_5531,N_5343);
or U5654 (N_5654,N_5375,N_5342);
or U5655 (N_5655,N_5246,N_5524);
xor U5656 (N_5656,N_5292,N_5567);
xor U5657 (N_5657,N_5482,N_5284);
nor U5658 (N_5658,N_5494,N_5573);
nor U5659 (N_5659,N_5509,N_5362);
or U5660 (N_5660,N_5417,N_5229);
xnor U5661 (N_5661,N_5507,N_5429);
nand U5662 (N_5662,N_5543,N_5577);
and U5663 (N_5663,N_5214,N_5317);
nor U5664 (N_5664,N_5499,N_5579);
and U5665 (N_5665,N_5223,N_5331);
or U5666 (N_5666,N_5454,N_5250);
xor U5667 (N_5667,N_5493,N_5366);
nor U5668 (N_5668,N_5588,N_5209);
nor U5669 (N_5669,N_5483,N_5421);
or U5670 (N_5670,N_5456,N_5337);
or U5671 (N_5671,N_5455,N_5576);
nor U5672 (N_5672,N_5285,N_5596);
xnor U5673 (N_5673,N_5303,N_5374);
or U5674 (N_5674,N_5277,N_5283);
xnor U5675 (N_5675,N_5385,N_5535);
or U5676 (N_5676,N_5339,N_5381);
and U5677 (N_5677,N_5213,N_5248);
or U5678 (N_5678,N_5500,N_5249);
xor U5679 (N_5679,N_5458,N_5510);
nor U5680 (N_5680,N_5200,N_5314);
xnor U5681 (N_5681,N_5556,N_5589);
xnor U5682 (N_5682,N_5377,N_5241);
or U5683 (N_5683,N_5294,N_5386);
nor U5684 (N_5684,N_5320,N_5464);
xor U5685 (N_5685,N_5452,N_5239);
and U5686 (N_5686,N_5513,N_5268);
or U5687 (N_5687,N_5340,N_5368);
nand U5688 (N_5688,N_5538,N_5259);
nor U5689 (N_5689,N_5282,N_5230);
xnor U5690 (N_5690,N_5308,N_5439);
or U5691 (N_5691,N_5276,N_5526);
nand U5692 (N_5692,N_5211,N_5378);
xor U5693 (N_5693,N_5575,N_5519);
nor U5694 (N_5694,N_5400,N_5324);
nand U5695 (N_5695,N_5363,N_5280);
and U5696 (N_5696,N_5351,N_5278);
nor U5697 (N_5697,N_5408,N_5434);
nor U5698 (N_5698,N_5321,N_5393);
or U5699 (N_5699,N_5557,N_5334);
xor U5700 (N_5700,N_5445,N_5485);
or U5701 (N_5701,N_5356,N_5245);
nand U5702 (N_5702,N_5548,N_5528);
and U5703 (N_5703,N_5428,N_5404);
nor U5704 (N_5704,N_5382,N_5210);
xnor U5705 (N_5705,N_5477,N_5347);
and U5706 (N_5706,N_5547,N_5522);
xnor U5707 (N_5707,N_5220,N_5472);
xor U5708 (N_5708,N_5532,N_5253);
nand U5709 (N_5709,N_5527,N_5212);
or U5710 (N_5710,N_5287,N_5502);
and U5711 (N_5711,N_5438,N_5569);
or U5712 (N_5712,N_5580,N_5410);
xnor U5713 (N_5713,N_5228,N_5262);
nand U5714 (N_5714,N_5275,N_5420);
xor U5715 (N_5715,N_5360,N_5498);
nor U5716 (N_5716,N_5329,N_5561);
nand U5717 (N_5717,N_5590,N_5369);
and U5718 (N_5718,N_5599,N_5451);
nand U5719 (N_5719,N_5562,N_5495);
nand U5720 (N_5720,N_5231,N_5447);
xor U5721 (N_5721,N_5319,N_5414);
or U5722 (N_5722,N_5346,N_5423);
or U5723 (N_5723,N_5476,N_5479);
xnor U5724 (N_5724,N_5332,N_5432);
and U5725 (N_5725,N_5508,N_5322);
nand U5726 (N_5726,N_5515,N_5348);
and U5727 (N_5727,N_5595,N_5299);
and U5728 (N_5728,N_5568,N_5570);
nand U5729 (N_5729,N_5518,N_5457);
and U5730 (N_5730,N_5376,N_5591);
or U5731 (N_5731,N_5520,N_5325);
xnor U5732 (N_5732,N_5310,N_5357);
or U5733 (N_5733,N_5470,N_5492);
nand U5734 (N_5734,N_5598,N_5537);
or U5735 (N_5735,N_5407,N_5328);
or U5736 (N_5736,N_5312,N_5364);
or U5737 (N_5737,N_5484,N_5358);
or U5738 (N_5738,N_5330,N_5387);
or U5739 (N_5739,N_5403,N_5460);
and U5740 (N_5740,N_5594,N_5232);
or U5741 (N_5741,N_5255,N_5453);
nand U5742 (N_5742,N_5449,N_5553);
nand U5743 (N_5743,N_5371,N_5242);
or U5744 (N_5744,N_5489,N_5584);
or U5745 (N_5745,N_5256,N_5293);
nor U5746 (N_5746,N_5426,N_5281);
and U5747 (N_5747,N_5240,N_5227);
nor U5748 (N_5748,N_5315,N_5399);
or U5749 (N_5749,N_5409,N_5559);
nor U5750 (N_5750,N_5542,N_5416);
and U5751 (N_5751,N_5383,N_5350);
xnor U5752 (N_5752,N_5288,N_5264);
xor U5753 (N_5753,N_5271,N_5297);
nor U5754 (N_5754,N_5306,N_5427);
or U5755 (N_5755,N_5260,N_5525);
nor U5756 (N_5756,N_5430,N_5367);
or U5757 (N_5757,N_5504,N_5349);
nand U5758 (N_5758,N_5506,N_5431);
nor U5759 (N_5759,N_5254,N_5448);
nor U5760 (N_5760,N_5305,N_5541);
and U5761 (N_5761,N_5269,N_5224);
and U5762 (N_5762,N_5521,N_5474);
xnor U5763 (N_5763,N_5443,N_5514);
xnor U5764 (N_5764,N_5326,N_5471);
nor U5765 (N_5765,N_5463,N_5295);
nand U5766 (N_5766,N_5437,N_5488);
nor U5767 (N_5767,N_5466,N_5461);
nand U5768 (N_5768,N_5592,N_5309);
xor U5769 (N_5769,N_5490,N_5597);
nor U5770 (N_5770,N_5436,N_5536);
nand U5771 (N_5771,N_5424,N_5215);
or U5772 (N_5772,N_5247,N_5395);
xor U5773 (N_5773,N_5486,N_5244);
nor U5774 (N_5774,N_5307,N_5336);
and U5775 (N_5775,N_5546,N_5345);
nor U5776 (N_5776,N_5304,N_5258);
and U5777 (N_5777,N_5373,N_5225);
and U5778 (N_5778,N_5222,N_5566);
nand U5779 (N_5779,N_5550,N_5344);
nand U5780 (N_5780,N_5540,N_5290);
xor U5781 (N_5781,N_5273,N_5355);
or U5782 (N_5782,N_5530,N_5572);
or U5783 (N_5783,N_5425,N_5379);
nand U5784 (N_5784,N_5418,N_5302);
or U5785 (N_5785,N_5204,N_5534);
nor U5786 (N_5786,N_5586,N_5391);
or U5787 (N_5787,N_5201,N_5523);
or U5788 (N_5788,N_5587,N_5266);
xor U5789 (N_5789,N_5353,N_5235);
nand U5790 (N_5790,N_5298,N_5450);
and U5791 (N_5791,N_5565,N_5401);
xor U5792 (N_5792,N_5564,N_5365);
nand U5793 (N_5793,N_5539,N_5582);
xor U5794 (N_5794,N_5552,N_5560);
or U5795 (N_5795,N_5469,N_5529);
and U5796 (N_5796,N_5252,N_5481);
or U5797 (N_5797,N_5226,N_5208);
xor U5798 (N_5798,N_5512,N_5384);
nand U5799 (N_5799,N_5341,N_5544);
nand U5800 (N_5800,N_5267,N_5258);
nand U5801 (N_5801,N_5497,N_5526);
or U5802 (N_5802,N_5530,N_5262);
nand U5803 (N_5803,N_5260,N_5484);
nor U5804 (N_5804,N_5247,N_5476);
and U5805 (N_5805,N_5449,N_5501);
nor U5806 (N_5806,N_5298,N_5465);
xnor U5807 (N_5807,N_5356,N_5300);
xor U5808 (N_5808,N_5352,N_5386);
and U5809 (N_5809,N_5401,N_5250);
or U5810 (N_5810,N_5235,N_5479);
nand U5811 (N_5811,N_5313,N_5496);
and U5812 (N_5812,N_5317,N_5212);
and U5813 (N_5813,N_5208,N_5340);
or U5814 (N_5814,N_5278,N_5452);
and U5815 (N_5815,N_5211,N_5261);
and U5816 (N_5816,N_5551,N_5521);
nand U5817 (N_5817,N_5439,N_5347);
nand U5818 (N_5818,N_5351,N_5256);
nor U5819 (N_5819,N_5566,N_5252);
xnor U5820 (N_5820,N_5400,N_5323);
or U5821 (N_5821,N_5529,N_5462);
and U5822 (N_5822,N_5266,N_5321);
or U5823 (N_5823,N_5414,N_5261);
or U5824 (N_5824,N_5359,N_5364);
and U5825 (N_5825,N_5298,N_5491);
nand U5826 (N_5826,N_5344,N_5529);
xor U5827 (N_5827,N_5455,N_5591);
and U5828 (N_5828,N_5554,N_5362);
nor U5829 (N_5829,N_5584,N_5223);
and U5830 (N_5830,N_5507,N_5300);
nand U5831 (N_5831,N_5270,N_5315);
nor U5832 (N_5832,N_5487,N_5557);
and U5833 (N_5833,N_5224,N_5570);
nor U5834 (N_5834,N_5329,N_5594);
xnor U5835 (N_5835,N_5490,N_5383);
nor U5836 (N_5836,N_5382,N_5208);
and U5837 (N_5837,N_5242,N_5459);
or U5838 (N_5838,N_5538,N_5211);
or U5839 (N_5839,N_5440,N_5250);
nor U5840 (N_5840,N_5531,N_5480);
xnor U5841 (N_5841,N_5505,N_5525);
nand U5842 (N_5842,N_5379,N_5375);
or U5843 (N_5843,N_5483,N_5422);
and U5844 (N_5844,N_5515,N_5363);
nor U5845 (N_5845,N_5280,N_5200);
and U5846 (N_5846,N_5305,N_5562);
nand U5847 (N_5847,N_5420,N_5591);
xor U5848 (N_5848,N_5519,N_5504);
xnor U5849 (N_5849,N_5267,N_5550);
xor U5850 (N_5850,N_5354,N_5224);
nand U5851 (N_5851,N_5289,N_5553);
or U5852 (N_5852,N_5414,N_5357);
and U5853 (N_5853,N_5412,N_5529);
xor U5854 (N_5854,N_5256,N_5371);
nand U5855 (N_5855,N_5581,N_5406);
or U5856 (N_5856,N_5454,N_5529);
nor U5857 (N_5857,N_5571,N_5317);
nor U5858 (N_5858,N_5412,N_5525);
nand U5859 (N_5859,N_5369,N_5431);
xor U5860 (N_5860,N_5344,N_5554);
or U5861 (N_5861,N_5283,N_5379);
and U5862 (N_5862,N_5467,N_5444);
xor U5863 (N_5863,N_5368,N_5358);
and U5864 (N_5864,N_5546,N_5210);
and U5865 (N_5865,N_5379,N_5585);
nand U5866 (N_5866,N_5378,N_5457);
nor U5867 (N_5867,N_5537,N_5562);
nand U5868 (N_5868,N_5359,N_5452);
or U5869 (N_5869,N_5525,N_5375);
nand U5870 (N_5870,N_5513,N_5434);
nor U5871 (N_5871,N_5315,N_5324);
xnor U5872 (N_5872,N_5565,N_5448);
nor U5873 (N_5873,N_5429,N_5432);
nand U5874 (N_5874,N_5418,N_5296);
and U5875 (N_5875,N_5362,N_5453);
nand U5876 (N_5876,N_5324,N_5434);
nand U5877 (N_5877,N_5252,N_5323);
and U5878 (N_5878,N_5458,N_5330);
and U5879 (N_5879,N_5336,N_5267);
or U5880 (N_5880,N_5316,N_5483);
nor U5881 (N_5881,N_5229,N_5383);
nor U5882 (N_5882,N_5232,N_5331);
nand U5883 (N_5883,N_5459,N_5283);
and U5884 (N_5884,N_5402,N_5343);
and U5885 (N_5885,N_5284,N_5428);
xnor U5886 (N_5886,N_5502,N_5416);
nand U5887 (N_5887,N_5513,N_5322);
or U5888 (N_5888,N_5230,N_5391);
or U5889 (N_5889,N_5468,N_5272);
xor U5890 (N_5890,N_5507,N_5222);
nor U5891 (N_5891,N_5516,N_5251);
or U5892 (N_5892,N_5450,N_5432);
nand U5893 (N_5893,N_5269,N_5306);
nor U5894 (N_5894,N_5481,N_5338);
and U5895 (N_5895,N_5391,N_5472);
and U5896 (N_5896,N_5293,N_5400);
or U5897 (N_5897,N_5243,N_5218);
nor U5898 (N_5898,N_5212,N_5296);
and U5899 (N_5899,N_5473,N_5323);
xor U5900 (N_5900,N_5201,N_5475);
or U5901 (N_5901,N_5261,N_5564);
xnor U5902 (N_5902,N_5397,N_5490);
nand U5903 (N_5903,N_5554,N_5322);
xor U5904 (N_5904,N_5294,N_5415);
or U5905 (N_5905,N_5281,N_5587);
nor U5906 (N_5906,N_5362,N_5572);
xor U5907 (N_5907,N_5299,N_5409);
and U5908 (N_5908,N_5555,N_5552);
nor U5909 (N_5909,N_5493,N_5387);
or U5910 (N_5910,N_5551,N_5590);
xor U5911 (N_5911,N_5468,N_5367);
nor U5912 (N_5912,N_5463,N_5395);
nand U5913 (N_5913,N_5525,N_5494);
xnor U5914 (N_5914,N_5311,N_5268);
xor U5915 (N_5915,N_5428,N_5259);
or U5916 (N_5916,N_5222,N_5465);
nand U5917 (N_5917,N_5386,N_5490);
nor U5918 (N_5918,N_5437,N_5448);
and U5919 (N_5919,N_5272,N_5285);
nand U5920 (N_5920,N_5239,N_5540);
nor U5921 (N_5921,N_5230,N_5474);
or U5922 (N_5922,N_5516,N_5295);
and U5923 (N_5923,N_5362,N_5414);
xor U5924 (N_5924,N_5554,N_5599);
xor U5925 (N_5925,N_5224,N_5280);
nor U5926 (N_5926,N_5445,N_5591);
nand U5927 (N_5927,N_5300,N_5512);
nor U5928 (N_5928,N_5219,N_5279);
nand U5929 (N_5929,N_5500,N_5338);
nor U5930 (N_5930,N_5358,N_5227);
or U5931 (N_5931,N_5531,N_5327);
nand U5932 (N_5932,N_5325,N_5248);
xnor U5933 (N_5933,N_5473,N_5360);
nand U5934 (N_5934,N_5567,N_5202);
nand U5935 (N_5935,N_5595,N_5273);
nor U5936 (N_5936,N_5491,N_5386);
or U5937 (N_5937,N_5235,N_5200);
and U5938 (N_5938,N_5595,N_5485);
nor U5939 (N_5939,N_5336,N_5264);
nor U5940 (N_5940,N_5258,N_5462);
nand U5941 (N_5941,N_5402,N_5454);
and U5942 (N_5942,N_5245,N_5574);
nand U5943 (N_5943,N_5424,N_5247);
xnor U5944 (N_5944,N_5523,N_5300);
xnor U5945 (N_5945,N_5441,N_5237);
xor U5946 (N_5946,N_5598,N_5487);
xor U5947 (N_5947,N_5421,N_5206);
nand U5948 (N_5948,N_5231,N_5315);
xnor U5949 (N_5949,N_5551,N_5319);
and U5950 (N_5950,N_5439,N_5557);
nand U5951 (N_5951,N_5573,N_5319);
and U5952 (N_5952,N_5318,N_5204);
xnor U5953 (N_5953,N_5268,N_5300);
nor U5954 (N_5954,N_5546,N_5587);
xnor U5955 (N_5955,N_5428,N_5489);
xnor U5956 (N_5956,N_5341,N_5507);
nand U5957 (N_5957,N_5553,N_5344);
nor U5958 (N_5958,N_5242,N_5531);
nand U5959 (N_5959,N_5392,N_5439);
and U5960 (N_5960,N_5516,N_5504);
nor U5961 (N_5961,N_5204,N_5512);
xnor U5962 (N_5962,N_5489,N_5259);
or U5963 (N_5963,N_5255,N_5297);
xor U5964 (N_5964,N_5246,N_5430);
nor U5965 (N_5965,N_5528,N_5509);
or U5966 (N_5966,N_5381,N_5237);
and U5967 (N_5967,N_5282,N_5477);
xor U5968 (N_5968,N_5464,N_5243);
nor U5969 (N_5969,N_5357,N_5214);
nor U5970 (N_5970,N_5319,N_5216);
or U5971 (N_5971,N_5536,N_5214);
nor U5972 (N_5972,N_5412,N_5218);
and U5973 (N_5973,N_5304,N_5451);
nand U5974 (N_5974,N_5556,N_5382);
nand U5975 (N_5975,N_5576,N_5539);
and U5976 (N_5976,N_5570,N_5506);
or U5977 (N_5977,N_5411,N_5362);
nand U5978 (N_5978,N_5400,N_5267);
nor U5979 (N_5979,N_5310,N_5252);
or U5980 (N_5980,N_5395,N_5501);
nand U5981 (N_5981,N_5508,N_5255);
and U5982 (N_5982,N_5285,N_5282);
nand U5983 (N_5983,N_5383,N_5258);
xnor U5984 (N_5984,N_5599,N_5396);
or U5985 (N_5985,N_5236,N_5438);
nor U5986 (N_5986,N_5292,N_5544);
and U5987 (N_5987,N_5497,N_5436);
and U5988 (N_5988,N_5591,N_5312);
or U5989 (N_5989,N_5231,N_5296);
nand U5990 (N_5990,N_5501,N_5463);
xor U5991 (N_5991,N_5320,N_5426);
nor U5992 (N_5992,N_5375,N_5218);
or U5993 (N_5993,N_5383,N_5349);
xnor U5994 (N_5994,N_5495,N_5581);
nand U5995 (N_5995,N_5351,N_5588);
nor U5996 (N_5996,N_5524,N_5230);
xor U5997 (N_5997,N_5410,N_5242);
nor U5998 (N_5998,N_5284,N_5498);
or U5999 (N_5999,N_5561,N_5550);
nor U6000 (N_6000,N_5707,N_5943);
and U6001 (N_6001,N_5618,N_5780);
xnor U6002 (N_6002,N_5837,N_5744);
or U6003 (N_6003,N_5939,N_5658);
nand U6004 (N_6004,N_5906,N_5991);
nor U6005 (N_6005,N_5924,N_5805);
nand U6006 (N_6006,N_5788,N_5617);
or U6007 (N_6007,N_5810,N_5623);
and U6008 (N_6008,N_5801,N_5749);
and U6009 (N_6009,N_5872,N_5789);
or U6010 (N_6010,N_5777,N_5735);
nor U6011 (N_6011,N_5908,N_5818);
and U6012 (N_6012,N_5624,N_5732);
xnor U6013 (N_6013,N_5947,N_5655);
or U6014 (N_6014,N_5697,N_5942);
nor U6015 (N_6015,N_5698,N_5733);
and U6016 (N_6016,N_5742,N_5967);
nand U6017 (N_6017,N_5954,N_5625);
and U6018 (N_6018,N_5798,N_5864);
or U6019 (N_6019,N_5791,N_5806);
nor U6020 (N_6020,N_5687,N_5729);
nand U6021 (N_6021,N_5979,N_5731);
or U6022 (N_6022,N_5686,N_5739);
or U6023 (N_6023,N_5907,N_5769);
nor U6024 (N_6024,N_5946,N_5875);
or U6025 (N_6025,N_5710,N_5711);
xor U6026 (N_6026,N_5845,N_5824);
xnor U6027 (N_6027,N_5935,N_5862);
nor U6028 (N_6028,N_5898,N_5737);
nand U6029 (N_6029,N_5955,N_5610);
and U6030 (N_6030,N_5855,N_5933);
xor U6031 (N_6031,N_5677,N_5870);
or U6032 (N_6032,N_5685,N_5869);
xor U6033 (N_6033,N_5985,N_5636);
and U6034 (N_6034,N_5668,N_5746);
nor U6035 (N_6035,N_5633,N_5866);
nand U6036 (N_6036,N_5682,N_5960);
xnor U6037 (N_6037,N_5723,N_5771);
nand U6038 (N_6038,N_5759,N_5721);
xor U6039 (N_6039,N_5702,N_5832);
and U6040 (N_6040,N_5889,N_5899);
or U6041 (N_6041,N_5650,N_5675);
or U6042 (N_6042,N_5774,N_5603);
and U6043 (N_6043,N_5852,N_5888);
or U6044 (N_6044,N_5911,N_5823);
or U6045 (N_6045,N_5612,N_5948);
or U6046 (N_6046,N_5830,N_5931);
or U6047 (N_6047,N_5868,N_5965);
nand U6048 (N_6048,N_5760,N_5716);
xnor U6049 (N_6049,N_5740,N_5683);
nor U6050 (N_6050,N_5909,N_5662);
nand U6051 (N_6051,N_5886,N_5772);
and U6052 (N_6052,N_5893,N_5792);
nand U6053 (N_6053,N_5797,N_5784);
and U6054 (N_6054,N_5644,N_5993);
nand U6055 (N_6055,N_5807,N_5622);
or U6056 (N_6056,N_5642,N_5666);
nor U6057 (N_6057,N_5902,N_5722);
nor U6058 (N_6058,N_5874,N_5794);
xor U6059 (N_6059,N_5951,N_5853);
xnor U6060 (N_6060,N_5885,N_5724);
and U6061 (N_6061,N_5693,N_5883);
xor U6062 (N_6062,N_5934,N_5843);
nor U6063 (N_6063,N_5858,N_5609);
xnor U6064 (N_6064,N_5753,N_5854);
xor U6065 (N_6065,N_5773,N_5982);
or U6066 (N_6066,N_5957,N_5988);
nor U6067 (N_6067,N_5983,N_5894);
nor U6068 (N_6068,N_5978,N_5826);
or U6069 (N_6069,N_5802,N_5630);
nor U6070 (N_6070,N_5614,N_5763);
xor U6071 (N_6071,N_5691,N_5790);
or U6072 (N_6072,N_5992,N_5660);
xnor U6073 (N_6073,N_5605,N_5775);
nor U6074 (N_6074,N_5767,N_5952);
xnor U6075 (N_6075,N_5646,N_5895);
or U6076 (N_6076,N_5627,N_5996);
and U6077 (N_6077,N_5997,N_5880);
nor U6078 (N_6078,N_5611,N_5913);
nor U6079 (N_6079,N_5674,N_5681);
xnor U6080 (N_6080,N_5847,N_5940);
and U6081 (N_6081,N_5961,N_5816);
or U6082 (N_6082,N_5938,N_5840);
nor U6083 (N_6083,N_5664,N_5941);
xnor U6084 (N_6084,N_5835,N_5704);
xor U6085 (N_6085,N_5833,N_5706);
and U6086 (N_6086,N_5669,N_5928);
or U6087 (N_6087,N_5663,N_5915);
xnor U6088 (N_6088,N_5901,N_5678);
xnor U6089 (N_6089,N_5828,N_5764);
nor U6090 (N_6090,N_5922,N_5918);
xor U6091 (N_6091,N_5844,N_5950);
nor U6092 (N_6092,N_5871,N_5607);
nor U6093 (N_6093,N_5689,N_5796);
or U6094 (N_6094,N_5708,N_5804);
nand U6095 (N_6095,N_5964,N_5857);
nand U6096 (N_6096,N_5989,N_5656);
and U6097 (N_6097,N_5990,N_5652);
nor U6098 (N_6098,N_5638,N_5713);
and U6099 (N_6099,N_5747,N_5719);
or U6100 (N_6100,N_5672,N_5756);
and U6101 (N_6101,N_5972,N_5679);
and U6102 (N_6102,N_5757,N_5766);
and U6103 (N_6103,N_5643,N_5980);
nand U6104 (N_6104,N_5851,N_5831);
xnor U6105 (N_6105,N_5912,N_5932);
or U6106 (N_6106,N_5998,N_5647);
or U6107 (N_6107,N_5970,N_5629);
nor U6108 (N_6108,N_5846,N_5945);
nor U6109 (N_6109,N_5859,N_5755);
nor U6110 (N_6110,N_5842,N_5953);
and U6111 (N_6111,N_5613,N_5999);
nor U6112 (N_6112,N_5606,N_5812);
xor U6113 (N_6113,N_5602,N_5659);
or U6114 (N_6114,N_5878,N_5994);
xor U6115 (N_6115,N_5700,N_5929);
nor U6116 (N_6116,N_5919,N_5717);
nand U6117 (N_6117,N_5782,N_5695);
xnor U6118 (N_6118,N_5971,N_5709);
nand U6119 (N_6119,N_5649,N_5949);
xor U6120 (N_6120,N_5936,N_5921);
or U6121 (N_6121,N_5631,N_5877);
nor U6122 (N_6122,N_5920,N_5986);
xnor U6123 (N_6123,N_5701,N_5822);
nor U6124 (N_6124,N_5838,N_5690);
and U6125 (N_6125,N_5688,N_5849);
xnor U6126 (N_6126,N_5910,N_5861);
xor U6127 (N_6127,N_5973,N_5848);
and U6128 (N_6128,N_5714,N_5778);
nand U6129 (N_6129,N_5968,N_5654);
xnor U6130 (N_6130,N_5754,N_5670);
or U6131 (N_6131,N_5692,N_5665);
nor U6132 (N_6132,N_5696,N_5975);
or U6133 (N_6133,N_5926,N_5632);
nor U6134 (N_6134,N_5839,N_5694);
xor U6135 (N_6135,N_5781,N_5800);
xnor U6136 (N_6136,N_5834,N_5923);
and U6137 (N_6137,N_5730,N_5819);
and U6138 (N_6138,N_5829,N_5863);
nor U6139 (N_6139,N_5745,N_5734);
nand U6140 (N_6140,N_5620,N_5640);
and U6141 (N_6141,N_5751,N_5787);
nand U6142 (N_6142,N_5969,N_5958);
nand U6143 (N_6143,N_5684,N_5616);
xnor U6144 (N_6144,N_5873,N_5601);
xnor U6145 (N_6145,N_5904,N_5628);
nor U6146 (N_6146,N_5977,N_5626);
nand U6147 (N_6147,N_5720,N_5892);
or U6148 (N_6148,N_5715,N_5779);
and U6149 (N_6149,N_5748,N_5813);
nand U6150 (N_6150,N_5884,N_5639);
nand U6151 (N_6151,N_5699,N_5850);
xor U6152 (N_6152,N_5661,N_5887);
and U6153 (N_6153,N_5600,N_5963);
nand U6154 (N_6154,N_5879,N_5765);
xnor U6155 (N_6155,N_5758,N_5761);
nand U6156 (N_6156,N_5783,N_5905);
and U6157 (N_6157,N_5786,N_5750);
xor U6158 (N_6158,N_5836,N_5881);
or U6159 (N_6159,N_5768,N_5741);
nor U6160 (N_6160,N_5811,N_5987);
xor U6161 (N_6161,N_5673,N_5653);
nand U6162 (N_6162,N_5927,N_5841);
nand U6163 (N_6163,N_5762,N_5937);
or U6164 (N_6164,N_5914,N_5785);
nor U6165 (N_6165,N_5814,N_5651);
and U6166 (N_6166,N_5865,N_5728);
nor U6167 (N_6167,N_5743,N_5995);
nand U6168 (N_6168,N_5635,N_5648);
nand U6169 (N_6169,N_5981,N_5817);
or U6170 (N_6170,N_5604,N_5820);
and U6171 (N_6171,N_5776,N_5712);
and U6172 (N_6172,N_5799,N_5671);
nor U6173 (N_6173,N_5821,N_5615);
or U6174 (N_6174,N_5736,N_5956);
nor U6175 (N_6175,N_5803,N_5897);
and U6176 (N_6176,N_5917,N_5856);
nor U6177 (N_6177,N_5641,N_5974);
and U6178 (N_6178,N_5738,N_5916);
nor U6179 (N_6179,N_5726,N_5657);
and U6180 (N_6180,N_5645,N_5680);
and U6181 (N_6181,N_5867,N_5718);
and U6182 (N_6182,N_5795,N_5976);
nor U6183 (N_6183,N_5984,N_5793);
xor U6184 (N_6184,N_5608,N_5703);
nand U6185 (N_6185,N_5966,N_5808);
nand U6186 (N_6186,N_5621,N_5903);
and U6187 (N_6187,N_5752,N_5827);
nor U6188 (N_6188,N_5900,N_5860);
nor U6189 (N_6189,N_5705,N_5809);
or U6190 (N_6190,N_5725,N_5925);
nand U6191 (N_6191,N_5634,N_5959);
nor U6192 (N_6192,N_5876,N_5896);
xnor U6193 (N_6193,N_5637,N_5882);
and U6194 (N_6194,N_5676,N_5770);
xor U6195 (N_6195,N_5825,N_5891);
nand U6196 (N_6196,N_5944,N_5727);
or U6197 (N_6197,N_5890,N_5667);
and U6198 (N_6198,N_5815,N_5930);
and U6199 (N_6199,N_5619,N_5962);
xnor U6200 (N_6200,N_5953,N_5990);
or U6201 (N_6201,N_5692,N_5835);
xnor U6202 (N_6202,N_5977,N_5868);
xnor U6203 (N_6203,N_5640,N_5757);
nand U6204 (N_6204,N_5849,N_5691);
nor U6205 (N_6205,N_5659,N_5828);
or U6206 (N_6206,N_5693,N_5833);
xnor U6207 (N_6207,N_5856,N_5645);
nor U6208 (N_6208,N_5640,N_5629);
xnor U6209 (N_6209,N_5644,N_5839);
or U6210 (N_6210,N_5982,N_5650);
and U6211 (N_6211,N_5719,N_5944);
nor U6212 (N_6212,N_5723,N_5919);
nand U6213 (N_6213,N_5922,N_5854);
nor U6214 (N_6214,N_5866,N_5672);
nand U6215 (N_6215,N_5901,N_5937);
xnor U6216 (N_6216,N_5818,N_5760);
or U6217 (N_6217,N_5981,N_5606);
xnor U6218 (N_6218,N_5772,N_5953);
nand U6219 (N_6219,N_5810,N_5640);
or U6220 (N_6220,N_5894,N_5892);
xor U6221 (N_6221,N_5646,N_5918);
nor U6222 (N_6222,N_5772,N_5712);
xor U6223 (N_6223,N_5686,N_5732);
nand U6224 (N_6224,N_5925,N_5703);
nor U6225 (N_6225,N_5637,N_5910);
nand U6226 (N_6226,N_5922,N_5820);
nand U6227 (N_6227,N_5655,N_5662);
nor U6228 (N_6228,N_5825,N_5724);
nand U6229 (N_6229,N_5853,N_5834);
nand U6230 (N_6230,N_5928,N_5848);
xnor U6231 (N_6231,N_5893,N_5666);
xnor U6232 (N_6232,N_5612,N_5702);
or U6233 (N_6233,N_5839,N_5723);
or U6234 (N_6234,N_5759,N_5694);
and U6235 (N_6235,N_5728,N_5732);
nor U6236 (N_6236,N_5799,N_5871);
nand U6237 (N_6237,N_5649,N_5982);
xnor U6238 (N_6238,N_5872,N_5663);
nand U6239 (N_6239,N_5652,N_5969);
nor U6240 (N_6240,N_5699,N_5620);
or U6241 (N_6241,N_5804,N_5933);
and U6242 (N_6242,N_5983,N_5718);
and U6243 (N_6243,N_5971,N_5730);
xor U6244 (N_6244,N_5883,N_5801);
or U6245 (N_6245,N_5642,N_5719);
nand U6246 (N_6246,N_5885,N_5803);
nand U6247 (N_6247,N_5825,N_5838);
and U6248 (N_6248,N_5843,N_5650);
xnor U6249 (N_6249,N_5797,N_5698);
nor U6250 (N_6250,N_5988,N_5678);
nor U6251 (N_6251,N_5674,N_5856);
nor U6252 (N_6252,N_5836,N_5916);
or U6253 (N_6253,N_5782,N_5755);
nor U6254 (N_6254,N_5999,N_5766);
nor U6255 (N_6255,N_5740,N_5718);
or U6256 (N_6256,N_5601,N_5688);
and U6257 (N_6257,N_5872,N_5800);
and U6258 (N_6258,N_5989,N_5951);
and U6259 (N_6259,N_5658,N_5811);
nand U6260 (N_6260,N_5848,N_5723);
nand U6261 (N_6261,N_5752,N_5758);
and U6262 (N_6262,N_5632,N_5981);
and U6263 (N_6263,N_5733,N_5900);
nor U6264 (N_6264,N_5607,N_5687);
and U6265 (N_6265,N_5614,N_5774);
and U6266 (N_6266,N_5732,N_5706);
nand U6267 (N_6267,N_5732,N_5937);
and U6268 (N_6268,N_5656,N_5900);
and U6269 (N_6269,N_5947,N_5830);
xnor U6270 (N_6270,N_5668,N_5902);
and U6271 (N_6271,N_5727,N_5835);
and U6272 (N_6272,N_5801,N_5751);
nor U6273 (N_6273,N_5957,N_5720);
or U6274 (N_6274,N_5933,N_5772);
or U6275 (N_6275,N_5826,N_5791);
xnor U6276 (N_6276,N_5871,N_5948);
nor U6277 (N_6277,N_5857,N_5886);
nor U6278 (N_6278,N_5833,N_5765);
nor U6279 (N_6279,N_5939,N_5879);
nand U6280 (N_6280,N_5721,N_5745);
or U6281 (N_6281,N_5748,N_5683);
and U6282 (N_6282,N_5694,N_5944);
nand U6283 (N_6283,N_5881,N_5801);
xor U6284 (N_6284,N_5621,N_5972);
nor U6285 (N_6285,N_5893,N_5897);
or U6286 (N_6286,N_5720,N_5698);
or U6287 (N_6287,N_5947,N_5791);
xnor U6288 (N_6288,N_5743,N_5742);
nor U6289 (N_6289,N_5729,N_5830);
or U6290 (N_6290,N_5719,N_5700);
nor U6291 (N_6291,N_5643,N_5730);
or U6292 (N_6292,N_5643,N_5765);
nand U6293 (N_6293,N_5989,N_5808);
xor U6294 (N_6294,N_5995,N_5654);
or U6295 (N_6295,N_5736,N_5791);
xnor U6296 (N_6296,N_5642,N_5876);
nand U6297 (N_6297,N_5817,N_5601);
nand U6298 (N_6298,N_5851,N_5869);
nand U6299 (N_6299,N_5883,N_5942);
or U6300 (N_6300,N_5636,N_5881);
and U6301 (N_6301,N_5774,N_5720);
or U6302 (N_6302,N_5656,N_5973);
nand U6303 (N_6303,N_5607,N_5709);
or U6304 (N_6304,N_5778,N_5930);
and U6305 (N_6305,N_5831,N_5943);
nor U6306 (N_6306,N_5803,N_5889);
xnor U6307 (N_6307,N_5873,N_5991);
xnor U6308 (N_6308,N_5969,N_5644);
or U6309 (N_6309,N_5921,N_5806);
xor U6310 (N_6310,N_5753,N_5696);
xnor U6311 (N_6311,N_5861,N_5937);
nor U6312 (N_6312,N_5698,N_5974);
and U6313 (N_6313,N_5746,N_5952);
nand U6314 (N_6314,N_5851,N_5833);
xor U6315 (N_6315,N_5921,N_5649);
nor U6316 (N_6316,N_5697,N_5916);
and U6317 (N_6317,N_5802,N_5627);
and U6318 (N_6318,N_5964,N_5931);
and U6319 (N_6319,N_5903,N_5923);
xor U6320 (N_6320,N_5750,N_5679);
and U6321 (N_6321,N_5807,N_5918);
and U6322 (N_6322,N_5755,N_5931);
or U6323 (N_6323,N_5852,N_5956);
nor U6324 (N_6324,N_5972,N_5622);
nand U6325 (N_6325,N_5847,N_5795);
nor U6326 (N_6326,N_5918,N_5939);
nor U6327 (N_6327,N_5940,N_5674);
nor U6328 (N_6328,N_5747,N_5788);
nor U6329 (N_6329,N_5718,N_5809);
nor U6330 (N_6330,N_5904,N_5903);
xnor U6331 (N_6331,N_5852,N_5688);
nand U6332 (N_6332,N_5740,N_5870);
and U6333 (N_6333,N_5923,N_5665);
nor U6334 (N_6334,N_5719,N_5813);
nor U6335 (N_6335,N_5690,N_5839);
or U6336 (N_6336,N_5787,N_5961);
nor U6337 (N_6337,N_5911,N_5804);
nor U6338 (N_6338,N_5732,N_5677);
nand U6339 (N_6339,N_5944,N_5783);
xor U6340 (N_6340,N_5782,N_5671);
nand U6341 (N_6341,N_5800,N_5637);
and U6342 (N_6342,N_5984,N_5810);
or U6343 (N_6343,N_5770,N_5778);
nand U6344 (N_6344,N_5755,N_5619);
or U6345 (N_6345,N_5794,N_5991);
nor U6346 (N_6346,N_5666,N_5806);
nor U6347 (N_6347,N_5618,N_5876);
nor U6348 (N_6348,N_5819,N_5825);
xnor U6349 (N_6349,N_5706,N_5728);
xnor U6350 (N_6350,N_5946,N_5879);
nor U6351 (N_6351,N_5909,N_5996);
and U6352 (N_6352,N_5699,N_5701);
nor U6353 (N_6353,N_5990,N_5759);
nand U6354 (N_6354,N_5797,N_5659);
nor U6355 (N_6355,N_5794,N_5906);
nor U6356 (N_6356,N_5635,N_5629);
nand U6357 (N_6357,N_5643,N_5900);
or U6358 (N_6358,N_5646,N_5746);
xor U6359 (N_6359,N_5879,N_5822);
or U6360 (N_6360,N_5763,N_5986);
nor U6361 (N_6361,N_5777,N_5809);
and U6362 (N_6362,N_5662,N_5712);
and U6363 (N_6363,N_5673,N_5824);
nor U6364 (N_6364,N_5786,N_5776);
nor U6365 (N_6365,N_5813,N_5961);
or U6366 (N_6366,N_5665,N_5966);
or U6367 (N_6367,N_5907,N_5603);
or U6368 (N_6368,N_5866,N_5858);
or U6369 (N_6369,N_5895,N_5831);
or U6370 (N_6370,N_5813,N_5835);
or U6371 (N_6371,N_5708,N_5920);
nor U6372 (N_6372,N_5778,N_5816);
xnor U6373 (N_6373,N_5948,N_5873);
and U6374 (N_6374,N_5843,N_5700);
or U6375 (N_6375,N_5935,N_5770);
nor U6376 (N_6376,N_5621,N_5709);
and U6377 (N_6377,N_5950,N_5974);
or U6378 (N_6378,N_5804,N_5903);
nor U6379 (N_6379,N_5838,N_5660);
and U6380 (N_6380,N_5859,N_5685);
nor U6381 (N_6381,N_5649,N_5673);
and U6382 (N_6382,N_5770,N_5846);
and U6383 (N_6383,N_5970,N_5800);
nand U6384 (N_6384,N_5794,N_5642);
nand U6385 (N_6385,N_5667,N_5640);
xor U6386 (N_6386,N_5605,N_5972);
and U6387 (N_6387,N_5733,N_5755);
xor U6388 (N_6388,N_5908,N_5989);
and U6389 (N_6389,N_5650,N_5914);
nand U6390 (N_6390,N_5932,N_5769);
nand U6391 (N_6391,N_5804,N_5939);
nand U6392 (N_6392,N_5896,N_5600);
and U6393 (N_6393,N_5629,N_5649);
or U6394 (N_6394,N_5803,N_5739);
and U6395 (N_6395,N_5903,N_5766);
xor U6396 (N_6396,N_5873,N_5958);
nor U6397 (N_6397,N_5920,N_5786);
and U6398 (N_6398,N_5711,N_5730);
nor U6399 (N_6399,N_5994,N_5803);
nor U6400 (N_6400,N_6036,N_6299);
xnor U6401 (N_6401,N_6298,N_6307);
xnor U6402 (N_6402,N_6341,N_6280);
nor U6403 (N_6403,N_6022,N_6336);
nand U6404 (N_6404,N_6112,N_6084);
nand U6405 (N_6405,N_6044,N_6312);
and U6406 (N_6406,N_6277,N_6079);
and U6407 (N_6407,N_6393,N_6060);
or U6408 (N_6408,N_6353,N_6064);
or U6409 (N_6409,N_6369,N_6134);
and U6410 (N_6410,N_6217,N_6264);
nand U6411 (N_6411,N_6174,N_6290);
nand U6412 (N_6412,N_6103,N_6049);
or U6413 (N_6413,N_6319,N_6200);
nor U6414 (N_6414,N_6287,N_6025);
nand U6415 (N_6415,N_6052,N_6105);
or U6416 (N_6416,N_6096,N_6180);
xor U6417 (N_6417,N_6172,N_6095);
and U6418 (N_6418,N_6254,N_6222);
nand U6419 (N_6419,N_6184,N_6041);
nand U6420 (N_6420,N_6042,N_6219);
or U6421 (N_6421,N_6098,N_6005);
and U6422 (N_6422,N_6032,N_6121);
nand U6423 (N_6423,N_6133,N_6156);
nand U6424 (N_6424,N_6283,N_6035);
and U6425 (N_6425,N_6255,N_6252);
xnor U6426 (N_6426,N_6304,N_6061);
nand U6427 (N_6427,N_6040,N_6232);
nand U6428 (N_6428,N_6395,N_6381);
nand U6429 (N_6429,N_6146,N_6192);
or U6430 (N_6430,N_6224,N_6116);
xor U6431 (N_6431,N_6333,N_6250);
nand U6432 (N_6432,N_6322,N_6068);
nand U6433 (N_6433,N_6015,N_6018);
nand U6434 (N_6434,N_6340,N_6372);
nand U6435 (N_6435,N_6039,N_6202);
and U6436 (N_6436,N_6159,N_6066);
and U6437 (N_6437,N_6392,N_6382);
nand U6438 (N_6438,N_6070,N_6108);
nor U6439 (N_6439,N_6050,N_6379);
xnor U6440 (N_6440,N_6198,N_6242);
nand U6441 (N_6441,N_6002,N_6065);
nor U6442 (N_6442,N_6323,N_6364);
and U6443 (N_6443,N_6339,N_6124);
xnor U6444 (N_6444,N_6157,N_6366);
xnor U6445 (N_6445,N_6263,N_6214);
and U6446 (N_6446,N_6245,N_6031);
and U6447 (N_6447,N_6115,N_6089);
or U6448 (N_6448,N_6361,N_6194);
xnor U6449 (N_6449,N_6123,N_6334);
nand U6450 (N_6450,N_6059,N_6296);
nand U6451 (N_6451,N_6346,N_6310);
and U6452 (N_6452,N_6344,N_6086);
xnor U6453 (N_6453,N_6145,N_6139);
and U6454 (N_6454,N_6099,N_6396);
and U6455 (N_6455,N_6094,N_6291);
and U6456 (N_6456,N_6046,N_6125);
xor U6457 (N_6457,N_6269,N_6024);
nand U6458 (N_6458,N_6003,N_6056);
xnor U6459 (N_6459,N_6072,N_6229);
nor U6460 (N_6460,N_6260,N_6330);
nand U6461 (N_6461,N_6132,N_6249);
and U6462 (N_6462,N_6138,N_6082);
nand U6463 (N_6463,N_6380,N_6142);
nand U6464 (N_6464,N_6211,N_6164);
or U6465 (N_6465,N_6152,N_6228);
nor U6466 (N_6466,N_6129,N_6062);
nor U6467 (N_6467,N_6197,N_6186);
nor U6468 (N_6468,N_6316,N_6216);
nor U6469 (N_6469,N_6267,N_6240);
xnor U6470 (N_6470,N_6092,N_6391);
and U6471 (N_6471,N_6350,N_6016);
xor U6472 (N_6472,N_6160,N_6375);
nor U6473 (N_6473,N_6302,N_6169);
nand U6474 (N_6474,N_6177,N_6276);
and U6475 (N_6475,N_6332,N_6221);
or U6476 (N_6476,N_6102,N_6080);
or U6477 (N_6477,N_6179,N_6397);
nor U6478 (N_6478,N_6203,N_6143);
nand U6479 (N_6479,N_6014,N_6337);
or U6480 (N_6480,N_6338,N_6356);
xor U6481 (N_6481,N_6107,N_6300);
nor U6482 (N_6482,N_6218,N_6207);
or U6483 (N_6483,N_6141,N_6370);
or U6484 (N_6484,N_6258,N_6013);
and U6485 (N_6485,N_6385,N_6342);
or U6486 (N_6486,N_6009,N_6210);
or U6487 (N_6487,N_6351,N_6233);
nand U6488 (N_6488,N_6153,N_6374);
or U6489 (N_6489,N_6308,N_6359);
nand U6490 (N_6490,N_6275,N_6326);
nor U6491 (N_6491,N_6320,N_6347);
nand U6492 (N_6492,N_6256,N_6030);
and U6493 (N_6493,N_6128,N_6273);
nor U6494 (N_6494,N_6193,N_6007);
or U6495 (N_6495,N_6085,N_6286);
or U6496 (N_6496,N_6176,N_6227);
or U6497 (N_6497,N_6166,N_6215);
nand U6498 (N_6498,N_6185,N_6367);
or U6499 (N_6499,N_6043,N_6093);
or U6500 (N_6500,N_6020,N_6029);
nand U6501 (N_6501,N_6243,N_6167);
nand U6502 (N_6502,N_6144,N_6027);
nand U6503 (N_6503,N_6135,N_6209);
xnor U6504 (N_6504,N_6189,N_6331);
xor U6505 (N_6505,N_6305,N_6274);
or U6506 (N_6506,N_6373,N_6165);
nor U6507 (N_6507,N_6151,N_6244);
or U6508 (N_6508,N_6278,N_6109);
nor U6509 (N_6509,N_6051,N_6261);
nand U6510 (N_6510,N_6126,N_6088);
or U6511 (N_6511,N_6309,N_6136);
nand U6512 (N_6512,N_6120,N_6220);
xnor U6513 (N_6513,N_6069,N_6377);
nand U6514 (N_6514,N_6208,N_6268);
xnor U6515 (N_6515,N_6294,N_6101);
nand U6516 (N_6516,N_6033,N_6281);
nor U6517 (N_6517,N_6226,N_6285);
nor U6518 (N_6518,N_6076,N_6137);
and U6519 (N_6519,N_6117,N_6148);
or U6520 (N_6520,N_6368,N_6113);
or U6521 (N_6521,N_6149,N_6329);
xor U6522 (N_6522,N_6131,N_6354);
and U6523 (N_6523,N_6190,N_6259);
nor U6524 (N_6524,N_6012,N_6321);
nand U6525 (N_6525,N_6171,N_6311);
xnor U6526 (N_6526,N_6386,N_6253);
nor U6527 (N_6527,N_6335,N_6362);
xnor U6528 (N_6528,N_6073,N_6114);
and U6529 (N_6529,N_6371,N_6378);
xnor U6530 (N_6530,N_6162,N_6236);
or U6531 (N_6531,N_6057,N_6063);
nor U6532 (N_6532,N_6201,N_6205);
nand U6533 (N_6533,N_6265,N_6071);
nor U6534 (N_6534,N_6325,N_6047);
or U6535 (N_6535,N_6127,N_6075);
or U6536 (N_6536,N_6279,N_6038);
or U6537 (N_6537,N_6158,N_6140);
nand U6538 (N_6538,N_6241,N_6303);
xor U6539 (N_6539,N_6196,N_6223);
and U6540 (N_6540,N_6213,N_6006);
and U6541 (N_6541,N_6122,N_6388);
or U6542 (N_6542,N_6188,N_6376);
nor U6543 (N_6543,N_6343,N_6118);
xnor U6544 (N_6544,N_6357,N_6078);
and U6545 (N_6545,N_6206,N_6204);
and U6546 (N_6546,N_6110,N_6272);
nor U6547 (N_6547,N_6023,N_6314);
xor U6548 (N_6548,N_6284,N_6246);
nor U6549 (N_6549,N_6389,N_6091);
and U6550 (N_6550,N_6363,N_6055);
nor U6551 (N_6551,N_6247,N_6045);
and U6552 (N_6552,N_6081,N_6355);
nor U6553 (N_6553,N_6074,N_6106);
or U6554 (N_6554,N_6001,N_6390);
xnor U6555 (N_6555,N_6383,N_6235);
nor U6556 (N_6556,N_6161,N_6147);
nor U6557 (N_6557,N_6238,N_6349);
xnor U6558 (N_6558,N_6288,N_6191);
xnor U6559 (N_6559,N_6262,N_6225);
and U6560 (N_6560,N_6234,N_6301);
nand U6561 (N_6561,N_6058,N_6028);
xnor U6562 (N_6562,N_6011,N_6348);
nand U6563 (N_6563,N_6239,N_6293);
or U6564 (N_6564,N_6021,N_6195);
nor U6565 (N_6565,N_6119,N_6170);
xnor U6566 (N_6566,N_6178,N_6087);
nand U6567 (N_6567,N_6394,N_6292);
or U6568 (N_6568,N_6212,N_6175);
and U6569 (N_6569,N_6154,N_6270);
xor U6570 (N_6570,N_6352,N_6054);
nand U6571 (N_6571,N_6387,N_6271);
nor U6572 (N_6572,N_6100,N_6317);
nand U6573 (N_6573,N_6248,N_6000);
xnor U6574 (N_6574,N_6199,N_6083);
xor U6575 (N_6575,N_6168,N_6097);
or U6576 (N_6576,N_6318,N_6017);
and U6577 (N_6577,N_6327,N_6282);
xor U6578 (N_6578,N_6399,N_6090);
or U6579 (N_6579,N_6026,N_6004);
xnor U6580 (N_6580,N_6360,N_6365);
xor U6581 (N_6581,N_6173,N_6104);
nand U6582 (N_6582,N_6077,N_6237);
or U6583 (N_6583,N_6297,N_6313);
and U6584 (N_6584,N_6324,N_6019);
and U6585 (N_6585,N_6328,N_6111);
and U6586 (N_6586,N_6306,N_6067);
nor U6587 (N_6587,N_6182,N_6266);
nand U6588 (N_6588,N_6155,N_6231);
xnor U6589 (N_6589,N_6257,N_6037);
or U6590 (N_6590,N_6034,N_6251);
nand U6591 (N_6591,N_6048,N_6130);
nand U6592 (N_6592,N_6295,N_6230);
xor U6593 (N_6593,N_6187,N_6315);
and U6594 (N_6594,N_6183,N_6010);
nand U6595 (N_6595,N_6345,N_6384);
and U6596 (N_6596,N_6053,N_6181);
xnor U6597 (N_6597,N_6163,N_6398);
and U6598 (N_6598,N_6358,N_6008);
xor U6599 (N_6599,N_6289,N_6150);
and U6600 (N_6600,N_6079,N_6219);
nand U6601 (N_6601,N_6303,N_6330);
xor U6602 (N_6602,N_6160,N_6210);
xnor U6603 (N_6603,N_6226,N_6078);
nand U6604 (N_6604,N_6351,N_6164);
xnor U6605 (N_6605,N_6047,N_6050);
or U6606 (N_6606,N_6090,N_6202);
nand U6607 (N_6607,N_6071,N_6348);
or U6608 (N_6608,N_6337,N_6110);
xor U6609 (N_6609,N_6190,N_6084);
nand U6610 (N_6610,N_6018,N_6026);
nor U6611 (N_6611,N_6255,N_6274);
xnor U6612 (N_6612,N_6117,N_6292);
nor U6613 (N_6613,N_6214,N_6310);
nor U6614 (N_6614,N_6355,N_6027);
nand U6615 (N_6615,N_6141,N_6303);
nand U6616 (N_6616,N_6000,N_6225);
xor U6617 (N_6617,N_6369,N_6322);
and U6618 (N_6618,N_6384,N_6132);
nand U6619 (N_6619,N_6110,N_6089);
or U6620 (N_6620,N_6072,N_6144);
nor U6621 (N_6621,N_6056,N_6116);
xnor U6622 (N_6622,N_6163,N_6090);
xor U6623 (N_6623,N_6073,N_6042);
nand U6624 (N_6624,N_6347,N_6177);
and U6625 (N_6625,N_6169,N_6251);
or U6626 (N_6626,N_6163,N_6061);
xnor U6627 (N_6627,N_6024,N_6252);
and U6628 (N_6628,N_6352,N_6225);
xor U6629 (N_6629,N_6144,N_6228);
and U6630 (N_6630,N_6248,N_6258);
or U6631 (N_6631,N_6370,N_6164);
or U6632 (N_6632,N_6298,N_6134);
xnor U6633 (N_6633,N_6130,N_6239);
nand U6634 (N_6634,N_6385,N_6180);
or U6635 (N_6635,N_6061,N_6178);
nand U6636 (N_6636,N_6146,N_6353);
xnor U6637 (N_6637,N_6215,N_6386);
or U6638 (N_6638,N_6005,N_6146);
or U6639 (N_6639,N_6048,N_6080);
nand U6640 (N_6640,N_6294,N_6062);
xnor U6641 (N_6641,N_6119,N_6220);
nand U6642 (N_6642,N_6253,N_6268);
xor U6643 (N_6643,N_6315,N_6358);
nor U6644 (N_6644,N_6108,N_6368);
xor U6645 (N_6645,N_6327,N_6172);
nor U6646 (N_6646,N_6133,N_6279);
xor U6647 (N_6647,N_6191,N_6103);
and U6648 (N_6648,N_6020,N_6304);
nand U6649 (N_6649,N_6219,N_6241);
or U6650 (N_6650,N_6301,N_6000);
and U6651 (N_6651,N_6325,N_6351);
xnor U6652 (N_6652,N_6086,N_6239);
and U6653 (N_6653,N_6300,N_6084);
nand U6654 (N_6654,N_6219,N_6197);
or U6655 (N_6655,N_6292,N_6124);
nor U6656 (N_6656,N_6005,N_6357);
or U6657 (N_6657,N_6195,N_6185);
and U6658 (N_6658,N_6281,N_6298);
and U6659 (N_6659,N_6251,N_6126);
nor U6660 (N_6660,N_6373,N_6147);
and U6661 (N_6661,N_6036,N_6005);
nand U6662 (N_6662,N_6364,N_6109);
xor U6663 (N_6663,N_6368,N_6034);
or U6664 (N_6664,N_6248,N_6107);
nand U6665 (N_6665,N_6060,N_6295);
and U6666 (N_6666,N_6118,N_6004);
or U6667 (N_6667,N_6342,N_6316);
nand U6668 (N_6668,N_6141,N_6322);
nor U6669 (N_6669,N_6210,N_6116);
and U6670 (N_6670,N_6299,N_6351);
xor U6671 (N_6671,N_6307,N_6295);
or U6672 (N_6672,N_6162,N_6093);
xor U6673 (N_6673,N_6249,N_6387);
nor U6674 (N_6674,N_6172,N_6381);
nand U6675 (N_6675,N_6101,N_6381);
xnor U6676 (N_6676,N_6321,N_6268);
nor U6677 (N_6677,N_6356,N_6047);
xnor U6678 (N_6678,N_6026,N_6222);
xnor U6679 (N_6679,N_6056,N_6075);
and U6680 (N_6680,N_6025,N_6034);
nor U6681 (N_6681,N_6352,N_6263);
xor U6682 (N_6682,N_6014,N_6319);
xor U6683 (N_6683,N_6344,N_6251);
xnor U6684 (N_6684,N_6159,N_6081);
nand U6685 (N_6685,N_6044,N_6279);
or U6686 (N_6686,N_6179,N_6181);
or U6687 (N_6687,N_6286,N_6038);
nand U6688 (N_6688,N_6334,N_6283);
nor U6689 (N_6689,N_6291,N_6085);
and U6690 (N_6690,N_6079,N_6054);
and U6691 (N_6691,N_6371,N_6166);
nor U6692 (N_6692,N_6372,N_6173);
nor U6693 (N_6693,N_6037,N_6143);
nor U6694 (N_6694,N_6222,N_6164);
or U6695 (N_6695,N_6034,N_6068);
or U6696 (N_6696,N_6233,N_6178);
nand U6697 (N_6697,N_6298,N_6150);
and U6698 (N_6698,N_6000,N_6148);
and U6699 (N_6699,N_6302,N_6290);
and U6700 (N_6700,N_6319,N_6356);
and U6701 (N_6701,N_6360,N_6280);
and U6702 (N_6702,N_6053,N_6357);
nor U6703 (N_6703,N_6189,N_6236);
and U6704 (N_6704,N_6101,N_6143);
nand U6705 (N_6705,N_6181,N_6266);
nand U6706 (N_6706,N_6257,N_6186);
xor U6707 (N_6707,N_6090,N_6269);
nand U6708 (N_6708,N_6228,N_6048);
or U6709 (N_6709,N_6373,N_6279);
or U6710 (N_6710,N_6016,N_6359);
xnor U6711 (N_6711,N_6059,N_6210);
xor U6712 (N_6712,N_6278,N_6269);
xor U6713 (N_6713,N_6156,N_6058);
nor U6714 (N_6714,N_6223,N_6111);
nand U6715 (N_6715,N_6347,N_6219);
nor U6716 (N_6716,N_6208,N_6138);
nand U6717 (N_6717,N_6142,N_6001);
or U6718 (N_6718,N_6321,N_6219);
and U6719 (N_6719,N_6263,N_6371);
nand U6720 (N_6720,N_6193,N_6004);
nor U6721 (N_6721,N_6033,N_6253);
nor U6722 (N_6722,N_6062,N_6132);
nand U6723 (N_6723,N_6344,N_6275);
and U6724 (N_6724,N_6072,N_6373);
nor U6725 (N_6725,N_6168,N_6309);
nor U6726 (N_6726,N_6153,N_6099);
nand U6727 (N_6727,N_6163,N_6297);
and U6728 (N_6728,N_6207,N_6157);
nor U6729 (N_6729,N_6136,N_6053);
xor U6730 (N_6730,N_6185,N_6029);
or U6731 (N_6731,N_6321,N_6144);
nor U6732 (N_6732,N_6318,N_6110);
and U6733 (N_6733,N_6026,N_6297);
xnor U6734 (N_6734,N_6101,N_6060);
xor U6735 (N_6735,N_6305,N_6368);
or U6736 (N_6736,N_6373,N_6250);
or U6737 (N_6737,N_6138,N_6307);
or U6738 (N_6738,N_6139,N_6192);
xnor U6739 (N_6739,N_6210,N_6013);
nand U6740 (N_6740,N_6399,N_6341);
nand U6741 (N_6741,N_6300,N_6078);
xnor U6742 (N_6742,N_6148,N_6212);
and U6743 (N_6743,N_6123,N_6314);
xor U6744 (N_6744,N_6060,N_6303);
xor U6745 (N_6745,N_6339,N_6323);
and U6746 (N_6746,N_6065,N_6191);
nor U6747 (N_6747,N_6259,N_6124);
and U6748 (N_6748,N_6145,N_6005);
xor U6749 (N_6749,N_6306,N_6381);
and U6750 (N_6750,N_6238,N_6342);
nor U6751 (N_6751,N_6388,N_6037);
xnor U6752 (N_6752,N_6135,N_6221);
nor U6753 (N_6753,N_6340,N_6065);
xnor U6754 (N_6754,N_6034,N_6008);
nand U6755 (N_6755,N_6054,N_6201);
and U6756 (N_6756,N_6352,N_6279);
nand U6757 (N_6757,N_6342,N_6261);
nand U6758 (N_6758,N_6376,N_6115);
or U6759 (N_6759,N_6252,N_6097);
nand U6760 (N_6760,N_6299,N_6084);
and U6761 (N_6761,N_6216,N_6129);
nand U6762 (N_6762,N_6115,N_6043);
xor U6763 (N_6763,N_6304,N_6384);
xnor U6764 (N_6764,N_6250,N_6282);
xor U6765 (N_6765,N_6222,N_6323);
or U6766 (N_6766,N_6036,N_6391);
and U6767 (N_6767,N_6140,N_6237);
and U6768 (N_6768,N_6040,N_6066);
xor U6769 (N_6769,N_6209,N_6091);
nor U6770 (N_6770,N_6074,N_6378);
nor U6771 (N_6771,N_6297,N_6092);
xnor U6772 (N_6772,N_6020,N_6197);
nor U6773 (N_6773,N_6269,N_6370);
and U6774 (N_6774,N_6197,N_6390);
nand U6775 (N_6775,N_6258,N_6032);
and U6776 (N_6776,N_6059,N_6094);
nor U6777 (N_6777,N_6263,N_6223);
and U6778 (N_6778,N_6136,N_6061);
and U6779 (N_6779,N_6014,N_6389);
and U6780 (N_6780,N_6257,N_6202);
or U6781 (N_6781,N_6377,N_6109);
or U6782 (N_6782,N_6048,N_6171);
xor U6783 (N_6783,N_6226,N_6355);
nor U6784 (N_6784,N_6010,N_6230);
nor U6785 (N_6785,N_6188,N_6305);
xor U6786 (N_6786,N_6373,N_6280);
or U6787 (N_6787,N_6065,N_6294);
xor U6788 (N_6788,N_6346,N_6267);
nor U6789 (N_6789,N_6085,N_6319);
nor U6790 (N_6790,N_6341,N_6260);
and U6791 (N_6791,N_6310,N_6303);
or U6792 (N_6792,N_6376,N_6091);
nand U6793 (N_6793,N_6082,N_6064);
or U6794 (N_6794,N_6398,N_6384);
or U6795 (N_6795,N_6324,N_6366);
nand U6796 (N_6796,N_6391,N_6038);
nor U6797 (N_6797,N_6334,N_6080);
or U6798 (N_6798,N_6059,N_6313);
nand U6799 (N_6799,N_6118,N_6033);
and U6800 (N_6800,N_6484,N_6497);
xor U6801 (N_6801,N_6670,N_6663);
xor U6802 (N_6802,N_6400,N_6774);
nor U6803 (N_6803,N_6405,N_6782);
nor U6804 (N_6804,N_6542,N_6417);
or U6805 (N_6805,N_6587,N_6625);
or U6806 (N_6806,N_6713,N_6518);
nor U6807 (N_6807,N_6621,N_6402);
nand U6808 (N_6808,N_6797,N_6596);
and U6809 (N_6809,N_6532,N_6473);
and U6810 (N_6810,N_6488,N_6432);
nand U6811 (N_6811,N_6793,N_6543);
and U6812 (N_6812,N_6748,N_6746);
nand U6813 (N_6813,N_6412,N_6468);
or U6814 (N_6814,N_6766,N_6733);
and U6815 (N_6815,N_6602,N_6641);
nand U6816 (N_6816,N_6667,N_6781);
and U6817 (N_6817,N_6608,N_6716);
and U6818 (N_6818,N_6649,N_6560);
xnor U6819 (N_6819,N_6692,N_6768);
nor U6820 (N_6820,N_6465,N_6493);
or U6821 (N_6821,N_6655,N_6592);
nor U6822 (N_6822,N_6423,N_6654);
xor U6823 (N_6823,N_6720,N_6409);
nor U6824 (N_6824,N_6688,N_6642);
xnor U6825 (N_6825,N_6447,N_6647);
nor U6826 (N_6826,N_6430,N_6666);
nand U6827 (N_6827,N_6433,N_6787);
nor U6828 (N_6828,N_6544,N_6718);
nand U6829 (N_6829,N_6615,N_6722);
and U6830 (N_6830,N_6457,N_6675);
and U6831 (N_6831,N_6777,N_6533);
xor U6832 (N_6832,N_6789,N_6515);
nor U6833 (N_6833,N_6479,N_6730);
nor U6834 (N_6834,N_6694,N_6507);
nand U6835 (N_6835,N_6734,N_6407);
or U6836 (N_6836,N_6579,N_6744);
nand U6837 (N_6837,N_6442,N_6411);
and U6838 (N_6838,N_6697,N_6617);
or U6839 (N_6839,N_6662,N_6652);
and U6840 (N_6840,N_6440,N_6434);
nor U6841 (N_6841,N_6584,N_6699);
xor U6842 (N_6842,N_6547,N_6426);
and U6843 (N_6843,N_6772,N_6645);
and U6844 (N_6844,N_6593,N_6798);
nor U6845 (N_6845,N_6745,N_6478);
or U6846 (N_6846,N_6415,N_6630);
xor U6847 (N_6847,N_6681,N_6472);
xor U6848 (N_6848,N_6622,N_6427);
or U6849 (N_6849,N_6682,N_6672);
nand U6850 (N_6850,N_6685,N_6438);
xor U6851 (N_6851,N_6714,N_6770);
and U6852 (N_6852,N_6595,N_6604);
xor U6853 (N_6853,N_6710,N_6704);
xor U6854 (N_6854,N_6643,N_6562);
nand U6855 (N_6855,N_6453,N_6790);
or U6856 (N_6856,N_6701,N_6657);
or U6857 (N_6857,N_6756,N_6709);
nand U6858 (N_6858,N_6715,N_6421);
nand U6859 (N_6859,N_6413,N_6420);
nand U6860 (N_6860,N_6445,N_6727);
or U6861 (N_6861,N_6758,N_6500);
nand U6862 (N_6862,N_6650,N_6698);
or U6863 (N_6863,N_6546,N_6728);
or U6864 (N_6864,N_6422,N_6762);
and U6865 (N_6865,N_6731,N_6477);
or U6866 (N_6866,N_6742,N_6786);
xnor U6867 (N_6867,N_6678,N_6598);
and U6868 (N_6868,N_6509,N_6606);
and U6869 (N_6869,N_6726,N_6449);
nor U6870 (N_6870,N_6503,N_6429);
and U6871 (N_6871,N_6700,N_6581);
xnor U6872 (N_6872,N_6740,N_6502);
or U6873 (N_6873,N_6609,N_6705);
nor U6874 (N_6874,N_6463,N_6570);
xnor U6875 (N_6875,N_6618,N_6737);
or U6876 (N_6876,N_6516,N_6446);
nand U6877 (N_6877,N_6611,N_6508);
and U6878 (N_6878,N_6640,N_6646);
nand U6879 (N_6879,N_6536,N_6696);
and U6880 (N_6880,N_6776,N_6600);
nand U6881 (N_6881,N_6582,N_6462);
xnor U6882 (N_6882,N_6638,N_6613);
and U6883 (N_6883,N_6464,N_6719);
nor U6884 (N_6884,N_6619,N_6495);
nand U6885 (N_6885,N_6401,N_6486);
and U6886 (N_6886,N_6636,N_6639);
nand U6887 (N_6887,N_6729,N_6741);
nor U6888 (N_6888,N_6751,N_6565);
nor U6889 (N_6889,N_6431,N_6512);
xnor U6890 (N_6890,N_6605,N_6573);
xor U6891 (N_6891,N_6796,N_6632);
and U6892 (N_6892,N_6548,N_6452);
or U6893 (N_6893,N_6563,N_6513);
nand U6894 (N_6894,N_6499,N_6761);
and U6895 (N_6895,N_6626,N_6448);
nand U6896 (N_6896,N_6648,N_6603);
and U6897 (N_6897,N_6491,N_6599);
nand U6898 (N_6898,N_6703,N_6559);
xnor U6899 (N_6899,N_6406,N_6764);
and U6900 (N_6900,N_6580,N_6708);
nand U6901 (N_6901,N_6754,N_6725);
and U6902 (N_6902,N_6634,N_6556);
or U6903 (N_6903,N_6624,N_6467);
or U6904 (N_6904,N_6724,N_6569);
or U6905 (N_6905,N_6674,N_6687);
or U6906 (N_6906,N_6784,N_6437);
nand U6907 (N_6907,N_6738,N_6778);
nand U6908 (N_6908,N_6676,N_6435);
nor U6909 (N_6909,N_6660,N_6444);
nor U6910 (N_6910,N_6476,N_6780);
nor U6911 (N_6911,N_6783,N_6763);
xnor U6912 (N_6912,N_6481,N_6585);
and U6913 (N_6913,N_6590,N_6623);
and U6914 (N_6914,N_6723,N_6506);
or U6915 (N_6915,N_6689,N_6616);
and U6916 (N_6916,N_6656,N_6571);
nor U6917 (N_6917,N_6735,N_6691);
xor U6918 (N_6918,N_6628,N_6671);
nor U6919 (N_6919,N_6436,N_6561);
nor U6920 (N_6920,N_6601,N_6549);
xnor U6921 (N_6921,N_6683,N_6456);
xor U6922 (N_6922,N_6458,N_6529);
xnor U6923 (N_6923,N_6665,N_6574);
xor U6924 (N_6924,N_6530,N_6610);
or U6925 (N_6925,N_6695,N_6554);
and U6926 (N_6926,N_6775,N_6607);
nor U6927 (N_6927,N_6749,N_6767);
xor U6928 (N_6928,N_6588,N_6597);
and U6929 (N_6929,N_6769,N_6760);
or U6930 (N_6930,N_6614,N_6576);
nand U6931 (N_6931,N_6577,N_6717);
nor U6932 (N_6932,N_6519,N_6664);
nor U6933 (N_6933,N_6525,N_6454);
nor U6934 (N_6934,N_6552,N_6589);
nand U6935 (N_6935,N_6788,N_6459);
nand U6936 (N_6936,N_6702,N_6550);
nand U6937 (N_6937,N_6526,N_6673);
and U6938 (N_6938,N_6644,N_6736);
and U6939 (N_6939,N_6586,N_6523);
nand U6940 (N_6940,N_6408,N_6711);
or U6941 (N_6941,N_6498,N_6679);
xnor U6942 (N_6942,N_6575,N_6686);
and U6943 (N_6943,N_6707,N_6537);
nand U6944 (N_6944,N_6633,N_6637);
and U6945 (N_6945,N_6690,N_6653);
nand U6946 (N_6946,N_6558,N_6441);
nand U6947 (N_6947,N_6771,N_6489);
or U6948 (N_6948,N_6651,N_6721);
or U6949 (N_6949,N_6494,N_6669);
or U6950 (N_6950,N_6480,N_6527);
and U6951 (N_6951,N_6572,N_6539);
xnor U6952 (N_6952,N_6794,N_6511);
nor U6953 (N_6953,N_6551,N_6680);
xor U6954 (N_6954,N_6799,N_6568);
or U6955 (N_6955,N_6792,N_6514);
nor U6956 (N_6956,N_6534,N_6424);
or U6957 (N_6957,N_6629,N_6564);
and U6958 (N_6958,N_6583,N_6416);
or U6959 (N_6959,N_6795,N_6578);
or U6960 (N_6960,N_6460,N_6471);
or U6961 (N_6961,N_6466,N_6419);
or U6962 (N_6962,N_6555,N_6779);
nor U6963 (N_6963,N_6684,N_6545);
and U6964 (N_6964,N_6635,N_6553);
or U6965 (N_6965,N_6566,N_6474);
and U6966 (N_6966,N_6404,N_6627);
nor U6967 (N_6967,N_6755,N_6747);
or U6968 (N_6968,N_6661,N_6482);
and U6969 (N_6969,N_6510,N_6418);
and U6970 (N_6970,N_6428,N_6620);
and U6971 (N_6971,N_6492,N_6451);
nor U6972 (N_6972,N_6475,N_6485);
nor U6973 (N_6973,N_6773,N_6414);
or U6974 (N_6974,N_6739,N_6557);
or U6975 (N_6975,N_6706,N_6455);
and U6976 (N_6976,N_6425,N_6757);
nor U6977 (N_6977,N_6791,N_6693);
nand U6978 (N_6978,N_6540,N_6496);
nand U6979 (N_6979,N_6759,N_6522);
and U6980 (N_6980,N_6567,N_6594);
and U6981 (N_6981,N_6677,N_6524);
or U6982 (N_6982,N_6487,N_6535);
nand U6983 (N_6983,N_6450,N_6538);
or U6984 (N_6984,N_6785,N_6541);
nor U6985 (N_6985,N_6668,N_6631);
nand U6986 (N_6986,N_6490,N_6469);
and U6987 (N_6987,N_6517,N_6591);
and U6988 (N_6988,N_6410,N_6612);
xnor U6989 (N_6989,N_6765,N_6521);
nand U6990 (N_6990,N_6505,N_6752);
xor U6991 (N_6991,N_6750,N_6531);
nor U6992 (N_6992,N_6443,N_6461);
and U6993 (N_6993,N_6403,N_6658);
xor U6994 (N_6994,N_6504,N_6483);
xnor U6995 (N_6995,N_6528,N_6743);
nand U6996 (N_6996,N_6659,N_6470);
xnor U6997 (N_6997,N_6753,N_6439);
xnor U6998 (N_6998,N_6520,N_6501);
nor U6999 (N_6999,N_6712,N_6732);
nand U7000 (N_7000,N_6487,N_6775);
nor U7001 (N_7001,N_6650,N_6440);
xor U7002 (N_7002,N_6517,N_6536);
and U7003 (N_7003,N_6526,N_6433);
and U7004 (N_7004,N_6603,N_6759);
nand U7005 (N_7005,N_6750,N_6510);
xnor U7006 (N_7006,N_6739,N_6488);
nand U7007 (N_7007,N_6798,N_6610);
nand U7008 (N_7008,N_6680,N_6409);
and U7009 (N_7009,N_6506,N_6784);
nor U7010 (N_7010,N_6780,N_6438);
xnor U7011 (N_7011,N_6540,N_6544);
nand U7012 (N_7012,N_6664,N_6495);
or U7013 (N_7013,N_6615,N_6635);
xnor U7014 (N_7014,N_6464,N_6566);
or U7015 (N_7015,N_6648,N_6514);
or U7016 (N_7016,N_6404,N_6577);
or U7017 (N_7017,N_6790,N_6681);
and U7018 (N_7018,N_6591,N_6522);
and U7019 (N_7019,N_6528,N_6739);
and U7020 (N_7020,N_6457,N_6664);
and U7021 (N_7021,N_6483,N_6420);
and U7022 (N_7022,N_6692,N_6762);
nor U7023 (N_7023,N_6632,N_6683);
xnor U7024 (N_7024,N_6432,N_6791);
or U7025 (N_7025,N_6619,N_6735);
xor U7026 (N_7026,N_6430,N_6659);
nand U7027 (N_7027,N_6491,N_6598);
nor U7028 (N_7028,N_6541,N_6478);
or U7029 (N_7029,N_6699,N_6773);
nand U7030 (N_7030,N_6615,N_6718);
or U7031 (N_7031,N_6572,N_6427);
and U7032 (N_7032,N_6519,N_6543);
or U7033 (N_7033,N_6643,N_6772);
or U7034 (N_7034,N_6645,N_6796);
xor U7035 (N_7035,N_6705,N_6778);
or U7036 (N_7036,N_6416,N_6660);
xor U7037 (N_7037,N_6446,N_6539);
and U7038 (N_7038,N_6672,N_6742);
nor U7039 (N_7039,N_6462,N_6612);
and U7040 (N_7040,N_6606,N_6631);
and U7041 (N_7041,N_6638,N_6757);
xnor U7042 (N_7042,N_6559,N_6510);
nor U7043 (N_7043,N_6431,N_6616);
and U7044 (N_7044,N_6560,N_6463);
nor U7045 (N_7045,N_6529,N_6774);
xnor U7046 (N_7046,N_6440,N_6656);
or U7047 (N_7047,N_6492,N_6634);
xor U7048 (N_7048,N_6797,N_6430);
or U7049 (N_7049,N_6735,N_6774);
or U7050 (N_7050,N_6674,N_6536);
nor U7051 (N_7051,N_6723,N_6530);
nor U7052 (N_7052,N_6480,N_6611);
or U7053 (N_7053,N_6723,N_6703);
and U7054 (N_7054,N_6490,N_6771);
xnor U7055 (N_7055,N_6585,N_6550);
nand U7056 (N_7056,N_6622,N_6648);
nand U7057 (N_7057,N_6701,N_6777);
nor U7058 (N_7058,N_6431,N_6426);
xnor U7059 (N_7059,N_6499,N_6527);
nand U7060 (N_7060,N_6669,N_6425);
or U7061 (N_7061,N_6604,N_6438);
and U7062 (N_7062,N_6725,N_6790);
or U7063 (N_7063,N_6479,N_6734);
nor U7064 (N_7064,N_6657,N_6791);
or U7065 (N_7065,N_6618,N_6436);
and U7066 (N_7066,N_6457,N_6637);
or U7067 (N_7067,N_6691,N_6712);
or U7068 (N_7068,N_6502,N_6736);
or U7069 (N_7069,N_6407,N_6473);
nor U7070 (N_7070,N_6574,N_6598);
nor U7071 (N_7071,N_6785,N_6584);
or U7072 (N_7072,N_6751,N_6400);
xor U7073 (N_7073,N_6665,N_6432);
nor U7074 (N_7074,N_6688,N_6753);
xnor U7075 (N_7075,N_6791,N_6595);
or U7076 (N_7076,N_6582,N_6729);
nor U7077 (N_7077,N_6436,N_6446);
nand U7078 (N_7078,N_6620,N_6553);
and U7079 (N_7079,N_6781,N_6732);
or U7080 (N_7080,N_6463,N_6665);
and U7081 (N_7081,N_6435,N_6428);
or U7082 (N_7082,N_6794,N_6487);
xnor U7083 (N_7083,N_6513,N_6582);
xor U7084 (N_7084,N_6717,N_6686);
nand U7085 (N_7085,N_6448,N_6561);
or U7086 (N_7086,N_6564,N_6624);
nor U7087 (N_7087,N_6527,N_6728);
and U7088 (N_7088,N_6552,N_6791);
nand U7089 (N_7089,N_6486,N_6722);
and U7090 (N_7090,N_6685,N_6467);
and U7091 (N_7091,N_6542,N_6471);
nor U7092 (N_7092,N_6585,N_6459);
nand U7093 (N_7093,N_6601,N_6433);
xnor U7094 (N_7094,N_6423,N_6777);
nor U7095 (N_7095,N_6524,N_6450);
nor U7096 (N_7096,N_6779,N_6455);
xnor U7097 (N_7097,N_6708,N_6438);
or U7098 (N_7098,N_6567,N_6751);
nand U7099 (N_7099,N_6547,N_6600);
nand U7100 (N_7100,N_6740,N_6742);
xnor U7101 (N_7101,N_6787,N_6634);
or U7102 (N_7102,N_6714,N_6495);
xnor U7103 (N_7103,N_6645,N_6773);
nor U7104 (N_7104,N_6557,N_6553);
nor U7105 (N_7105,N_6615,N_6776);
or U7106 (N_7106,N_6537,N_6670);
nor U7107 (N_7107,N_6575,N_6657);
xnor U7108 (N_7108,N_6679,N_6745);
xor U7109 (N_7109,N_6557,N_6780);
xor U7110 (N_7110,N_6637,N_6542);
nand U7111 (N_7111,N_6754,N_6412);
nand U7112 (N_7112,N_6474,N_6706);
or U7113 (N_7113,N_6515,N_6548);
or U7114 (N_7114,N_6644,N_6774);
and U7115 (N_7115,N_6726,N_6446);
nor U7116 (N_7116,N_6600,N_6748);
nor U7117 (N_7117,N_6655,N_6741);
and U7118 (N_7118,N_6432,N_6718);
nand U7119 (N_7119,N_6749,N_6495);
nor U7120 (N_7120,N_6410,N_6487);
or U7121 (N_7121,N_6486,N_6605);
nand U7122 (N_7122,N_6715,N_6772);
nor U7123 (N_7123,N_6668,N_6418);
xor U7124 (N_7124,N_6430,N_6779);
nand U7125 (N_7125,N_6615,N_6595);
nand U7126 (N_7126,N_6488,N_6625);
nor U7127 (N_7127,N_6661,N_6729);
nor U7128 (N_7128,N_6734,N_6649);
or U7129 (N_7129,N_6718,N_6692);
nor U7130 (N_7130,N_6691,N_6504);
and U7131 (N_7131,N_6463,N_6480);
nand U7132 (N_7132,N_6418,N_6450);
nor U7133 (N_7133,N_6625,N_6402);
xor U7134 (N_7134,N_6506,N_6640);
and U7135 (N_7135,N_6735,N_6623);
xor U7136 (N_7136,N_6640,N_6634);
nand U7137 (N_7137,N_6593,N_6596);
and U7138 (N_7138,N_6596,N_6643);
and U7139 (N_7139,N_6753,N_6790);
or U7140 (N_7140,N_6717,N_6655);
nor U7141 (N_7141,N_6752,N_6409);
nor U7142 (N_7142,N_6546,N_6507);
nor U7143 (N_7143,N_6424,N_6504);
or U7144 (N_7144,N_6490,N_6425);
xor U7145 (N_7145,N_6652,N_6636);
nor U7146 (N_7146,N_6753,N_6461);
nand U7147 (N_7147,N_6771,N_6552);
or U7148 (N_7148,N_6668,N_6470);
xor U7149 (N_7149,N_6727,N_6504);
and U7150 (N_7150,N_6474,N_6699);
nor U7151 (N_7151,N_6739,N_6789);
xor U7152 (N_7152,N_6624,N_6787);
or U7153 (N_7153,N_6708,N_6780);
or U7154 (N_7154,N_6702,N_6574);
or U7155 (N_7155,N_6605,N_6708);
nand U7156 (N_7156,N_6470,N_6524);
nor U7157 (N_7157,N_6660,N_6430);
xnor U7158 (N_7158,N_6419,N_6690);
nand U7159 (N_7159,N_6433,N_6643);
nor U7160 (N_7160,N_6545,N_6783);
or U7161 (N_7161,N_6701,N_6408);
nor U7162 (N_7162,N_6467,N_6625);
and U7163 (N_7163,N_6565,N_6757);
or U7164 (N_7164,N_6446,N_6708);
and U7165 (N_7165,N_6498,N_6547);
nor U7166 (N_7166,N_6790,N_6682);
or U7167 (N_7167,N_6655,N_6721);
nand U7168 (N_7168,N_6484,N_6714);
xor U7169 (N_7169,N_6487,N_6653);
or U7170 (N_7170,N_6404,N_6433);
or U7171 (N_7171,N_6506,N_6690);
xnor U7172 (N_7172,N_6488,N_6777);
nor U7173 (N_7173,N_6494,N_6590);
xnor U7174 (N_7174,N_6584,N_6476);
and U7175 (N_7175,N_6775,N_6595);
or U7176 (N_7176,N_6669,N_6648);
and U7177 (N_7177,N_6407,N_6501);
or U7178 (N_7178,N_6689,N_6495);
xnor U7179 (N_7179,N_6555,N_6425);
or U7180 (N_7180,N_6584,N_6498);
xor U7181 (N_7181,N_6427,N_6585);
nand U7182 (N_7182,N_6723,N_6671);
nor U7183 (N_7183,N_6518,N_6674);
xor U7184 (N_7184,N_6792,N_6422);
or U7185 (N_7185,N_6533,N_6767);
nand U7186 (N_7186,N_6748,N_6649);
xnor U7187 (N_7187,N_6442,N_6718);
nand U7188 (N_7188,N_6560,N_6697);
nor U7189 (N_7189,N_6673,N_6452);
and U7190 (N_7190,N_6673,N_6722);
nor U7191 (N_7191,N_6676,N_6516);
xnor U7192 (N_7192,N_6500,N_6644);
or U7193 (N_7193,N_6475,N_6756);
nor U7194 (N_7194,N_6562,N_6681);
and U7195 (N_7195,N_6712,N_6658);
nor U7196 (N_7196,N_6457,N_6493);
xor U7197 (N_7197,N_6766,N_6698);
or U7198 (N_7198,N_6783,N_6677);
or U7199 (N_7199,N_6633,N_6459);
nand U7200 (N_7200,N_6883,N_7073);
or U7201 (N_7201,N_6854,N_6871);
or U7202 (N_7202,N_6849,N_7195);
xor U7203 (N_7203,N_7144,N_7011);
and U7204 (N_7204,N_7159,N_6879);
nand U7205 (N_7205,N_7179,N_7187);
nand U7206 (N_7206,N_6991,N_7010);
xnor U7207 (N_7207,N_6996,N_7133);
and U7208 (N_7208,N_7130,N_7048);
xor U7209 (N_7209,N_6902,N_6964);
nand U7210 (N_7210,N_7118,N_7165);
nor U7211 (N_7211,N_6842,N_6889);
nand U7212 (N_7212,N_7002,N_6838);
nor U7213 (N_7213,N_6868,N_7197);
xor U7214 (N_7214,N_6853,N_6805);
and U7215 (N_7215,N_6983,N_6888);
nor U7216 (N_7216,N_7193,N_7125);
nor U7217 (N_7217,N_6811,N_6900);
xnor U7218 (N_7218,N_6814,N_7140);
or U7219 (N_7219,N_6926,N_7035);
and U7220 (N_7220,N_6917,N_6828);
nand U7221 (N_7221,N_7062,N_6867);
xnor U7222 (N_7222,N_7168,N_6945);
xnor U7223 (N_7223,N_7163,N_7024);
and U7224 (N_7224,N_6920,N_7131);
xnor U7225 (N_7225,N_6940,N_7136);
nand U7226 (N_7226,N_7094,N_6881);
nand U7227 (N_7227,N_7051,N_6815);
or U7228 (N_7228,N_7107,N_7000);
nand U7229 (N_7229,N_6885,N_6998);
or U7230 (N_7230,N_6872,N_6919);
nor U7231 (N_7231,N_6905,N_6890);
nor U7232 (N_7232,N_7146,N_7007);
or U7233 (N_7233,N_6858,N_7087);
or U7234 (N_7234,N_6812,N_6826);
or U7235 (N_7235,N_7019,N_6984);
or U7236 (N_7236,N_7192,N_7169);
or U7237 (N_7237,N_7040,N_6975);
nor U7238 (N_7238,N_6801,N_6995);
or U7239 (N_7239,N_6957,N_7045);
xnor U7240 (N_7240,N_6891,N_7154);
nand U7241 (N_7241,N_6845,N_6950);
xnor U7242 (N_7242,N_6852,N_7149);
xor U7243 (N_7243,N_7185,N_6808);
or U7244 (N_7244,N_6892,N_6921);
and U7245 (N_7245,N_6873,N_7079);
nor U7246 (N_7246,N_7139,N_7138);
xor U7247 (N_7247,N_7114,N_6869);
xor U7248 (N_7248,N_7120,N_6914);
nor U7249 (N_7249,N_7038,N_7137);
nor U7250 (N_7250,N_7009,N_6912);
and U7251 (N_7251,N_6954,N_6836);
and U7252 (N_7252,N_6972,N_6870);
xor U7253 (N_7253,N_7027,N_6832);
or U7254 (N_7254,N_7116,N_7054);
xor U7255 (N_7255,N_7059,N_6865);
or U7256 (N_7256,N_6857,N_7039);
nand U7257 (N_7257,N_6863,N_7157);
xnor U7258 (N_7258,N_7181,N_7050);
nand U7259 (N_7259,N_7109,N_7156);
or U7260 (N_7260,N_7106,N_6913);
or U7261 (N_7261,N_7098,N_6880);
or U7262 (N_7262,N_6966,N_7003);
xnor U7263 (N_7263,N_6800,N_7173);
and U7264 (N_7264,N_7084,N_6804);
nand U7265 (N_7265,N_7055,N_6882);
and U7266 (N_7266,N_6947,N_7028);
nand U7267 (N_7267,N_7115,N_6990);
nand U7268 (N_7268,N_7162,N_6915);
xor U7269 (N_7269,N_7012,N_6884);
nand U7270 (N_7270,N_6978,N_7014);
and U7271 (N_7271,N_7151,N_7167);
nor U7272 (N_7272,N_6807,N_7170);
nand U7273 (N_7273,N_7015,N_7070);
or U7274 (N_7274,N_6893,N_7194);
and U7275 (N_7275,N_7111,N_7066);
xnor U7276 (N_7276,N_7025,N_7158);
or U7277 (N_7277,N_7126,N_6822);
xnor U7278 (N_7278,N_7102,N_6830);
nor U7279 (N_7279,N_7089,N_6951);
xor U7280 (N_7280,N_6965,N_6819);
xnor U7281 (N_7281,N_6813,N_6887);
nor U7282 (N_7282,N_7005,N_6861);
or U7283 (N_7283,N_6939,N_7046);
nand U7284 (N_7284,N_6925,N_6859);
or U7285 (N_7285,N_7033,N_7152);
xnor U7286 (N_7286,N_7017,N_6907);
xnor U7287 (N_7287,N_6875,N_6855);
and U7288 (N_7288,N_7075,N_7117);
nand U7289 (N_7289,N_6961,N_6993);
xor U7290 (N_7290,N_6904,N_6970);
nand U7291 (N_7291,N_6820,N_6982);
xor U7292 (N_7292,N_7072,N_6924);
nor U7293 (N_7293,N_7036,N_7037);
xnor U7294 (N_7294,N_6897,N_6846);
xnor U7295 (N_7295,N_7099,N_6829);
and U7296 (N_7296,N_6910,N_7123);
nand U7297 (N_7297,N_6909,N_6877);
or U7298 (N_7298,N_7199,N_6840);
or U7299 (N_7299,N_7064,N_6929);
or U7300 (N_7300,N_7177,N_7067);
or U7301 (N_7301,N_6860,N_7143);
nand U7302 (N_7302,N_6806,N_6927);
and U7303 (N_7303,N_6944,N_7128);
nand U7304 (N_7304,N_6974,N_6958);
xnor U7305 (N_7305,N_6994,N_6850);
nor U7306 (N_7306,N_6918,N_6862);
xor U7307 (N_7307,N_6844,N_7078);
or U7308 (N_7308,N_6946,N_7030);
nand U7309 (N_7309,N_7150,N_7020);
and U7310 (N_7310,N_7043,N_6930);
nand U7311 (N_7311,N_6968,N_7122);
nand U7312 (N_7312,N_6816,N_6823);
nor U7313 (N_7313,N_6827,N_6803);
xor U7314 (N_7314,N_6981,N_7093);
nand U7315 (N_7315,N_6878,N_6864);
nand U7316 (N_7316,N_6825,N_7057);
xor U7317 (N_7317,N_6977,N_7182);
nand U7318 (N_7318,N_7108,N_7153);
and U7319 (N_7319,N_7100,N_7077);
xnor U7320 (N_7320,N_6971,N_6931);
and U7321 (N_7321,N_7095,N_6948);
nand U7322 (N_7322,N_7001,N_7056);
and U7323 (N_7323,N_7141,N_6979);
xnor U7324 (N_7324,N_7063,N_7080);
xor U7325 (N_7325,N_6848,N_6980);
xnor U7326 (N_7326,N_6901,N_7082);
or U7327 (N_7327,N_6956,N_6923);
or U7328 (N_7328,N_7161,N_6936);
xor U7329 (N_7329,N_7196,N_6903);
xor U7330 (N_7330,N_6833,N_7147);
or U7331 (N_7331,N_6906,N_6809);
nand U7332 (N_7332,N_7189,N_6999);
nand U7333 (N_7333,N_7006,N_6988);
or U7334 (N_7334,N_7069,N_7041);
and U7335 (N_7335,N_6898,N_6895);
and U7336 (N_7336,N_6989,N_7183);
nand U7337 (N_7337,N_7174,N_7091);
nor U7338 (N_7338,N_7053,N_7191);
and U7339 (N_7339,N_7086,N_6866);
or U7340 (N_7340,N_7121,N_6943);
and U7341 (N_7341,N_6843,N_7112);
and U7342 (N_7342,N_7097,N_7032);
xnor U7343 (N_7343,N_7124,N_6955);
nor U7344 (N_7344,N_7186,N_7119);
and U7345 (N_7345,N_6959,N_6935);
xor U7346 (N_7346,N_7029,N_6886);
xnor U7347 (N_7347,N_6802,N_7088);
or U7348 (N_7348,N_7058,N_7178);
xnor U7349 (N_7349,N_6834,N_7074);
or U7350 (N_7350,N_6942,N_6841);
xor U7351 (N_7351,N_6899,N_7127);
or U7352 (N_7352,N_7184,N_7044);
nand U7353 (N_7353,N_6876,N_6967);
nor U7354 (N_7354,N_7101,N_6952);
nor U7355 (N_7355,N_6831,N_7008);
or U7356 (N_7356,N_6937,N_7188);
or U7357 (N_7357,N_6824,N_6821);
and U7358 (N_7358,N_6856,N_7166);
nand U7359 (N_7359,N_7180,N_7083);
or U7360 (N_7360,N_6992,N_7081);
xor U7361 (N_7361,N_7052,N_6916);
nor U7362 (N_7362,N_6934,N_6938);
nor U7363 (N_7363,N_6969,N_7071);
xnor U7364 (N_7364,N_7004,N_7061);
nor U7365 (N_7365,N_6817,N_7026);
and U7366 (N_7366,N_6894,N_6837);
nand U7367 (N_7367,N_6987,N_7018);
nor U7368 (N_7368,N_6949,N_7103);
xnor U7369 (N_7369,N_7096,N_7160);
nand U7370 (N_7370,N_7129,N_7113);
xnor U7371 (N_7371,N_7021,N_7175);
nand U7372 (N_7372,N_6962,N_6839);
xnor U7373 (N_7373,N_7135,N_7155);
nor U7374 (N_7374,N_7092,N_7023);
nand U7375 (N_7375,N_6960,N_7104);
and U7376 (N_7376,N_6986,N_7013);
and U7377 (N_7377,N_7164,N_7047);
or U7378 (N_7378,N_6911,N_7060);
or U7379 (N_7379,N_7076,N_7172);
nand U7380 (N_7380,N_7190,N_7105);
nor U7381 (N_7381,N_7132,N_7042);
nor U7382 (N_7382,N_6835,N_6953);
xnor U7383 (N_7383,N_6810,N_7031);
xor U7384 (N_7384,N_6851,N_7065);
xnor U7385 (N_7385,N_6928,N_7176);
or U7386 (N_7386,N_7148,N_7171);
or U7387 (N_7387,N_6941,N_7085);
nor U7388 (N_7388,N_6997,N_7022);
or U7389 (N_7389,N_7110,N_7068);
nor U7390 (N_7390,N_6973,N_7090);
and U7391 (N_7391,N_6847,N_7145);
nand U7392 (N_7392,N_7016,N_7049);
or U7393 (N_7393,N_7198,N_7034);
or U7394 (N_7394,N_7142,N_6896);
xor U7395 (N_7395,N_6818,N_6933);
nor U7396 (N_7396,N_6976,N_7134);
nand U7397 (N_7397,N_6922,N_6932);
nor U7398 (N_7398,N_6908,N_6963);
xnor U7399 (N_7399,N_6874,N_6985);
or U7400 (N_7400,N_7078,N_6896);
or U7401 (N_7401,N_6931,N_6815);
or U7402 (N_7402,N_7137,N_6834);
xnor U7403 (N_7403,N_7016,N_6999);
nand U7404 (N_7404,N_7105,N_6927);
nor U7405 (N_7405,N_6967,N_6927);
and U7406 (N_7406,N_6802,N_7115);
nand U7407 (N_7407,N_6800,N_6903);
xor U7408 (N_7408,N_6852,N_6929);
and U7409 (N_7409,N_7185,N_7072);
nand U7410 (N_7410,N_6960,N_6937);
xor U7411 (N_7411,N_7027,N_7165);
nand U7412 (N_7412,N_6932,N_7138);
nand U7413 (N_7413,N_6883,N_6901);
and U7414 (N_7414,N_6930,N_6969);
and U7415 (N_7415,N_7083,N_6808);
nand U7416 (N_7416,N_6908,N_6974);
xor U7417 (N_7417,N_6991,N_7172);
nor U7418 (N_7418,N_7095,N_7156);
nor U7419 (N_7419,N_6866,N_7072);
or U7420 (N_7420,N_7184,N_6913);
nand U7421 (N_7421,N_6863,N_6887);
xor U7422 (N_7422,N_7185,N_7167);
and U7423 (N_7423,N_6803,N_7180);
nand U7424 (N_7424,N_7032,N_6878);
or U7425 (N_7425,N_6932,N_6800);
or U7426 (N_7426,N_6916,N_6884);
nor U7427 (N_7427,N_7190,N_6801);
nor U7428 (N_7428,N_6917,N_7060);
or U7429 (N_7429,N_6865,N_7144);
xor U7430 (N_7430,N_6973,N_6974);
nand U7431 (N_7431,N_6901,N_6949);
xnor U7432 (N_7432,N_7141,N_6968);
nor U7433 (N_7433,N_6812,N_7120);
nor U7434 (N_7434,N_6859,N_7004);
or U7435 (N_7435,N_6825,N_6906);
nand U7436 (N_7436,N_7058,N_7094);
xnor U7437 (N_7437,N_6860,N_6846);
nor U7438 (N_7438,N_6887,N_6975);
nand U7439 (N_7439,N_6845,N_7014);
nand U7440 (N_7440,N_7096,N_6914);
nor U7441 (N_7441,N_7184,N_7193);
xnor U7442 (N_7442,N_6995,N_6849);
nand U7443 (N_7443,N_6903,N_7114);
nor U7444 (N_7444,N_6818,N_7179);
or U7445 (N_7445,N_6874,N_6888);
or U7446 (N_7446,N_7167,N_6952);
nand U7447 (N_7447,N_7073,N_7154);
nor U7448 (N_7448,N_6897,N_6975);
xor U7449 (N_7449,N_7036,N_6975);
nor U7450 (N_7450,N_6828,N_6937);
nor U7451 (N_7451,N_7197,N_6978);
or U7452 (N_7452,N_7144,N_6933);
and U7453 (N_7453,N_6867,N_6925);
nor U7454 (N_7454,N_7127,N_7195);
nand U7455 (N_7455,N_6921,N_7056);
nor U7456 (N_7456,N_7188,N_7024);
or U7457 (N_7457,N_6813,N_6926);
xnor U7458 (N_7458,N_7167,N_6962);
nor U7459 (N_7459,N_6891,N_6941);
or U7460 (N_7460,N_7045,N_7153);
xnor U7461 (N_7461,N_7133,N_7135);
nand U7462 (N_7462,N_7095,N_6897);
xor U7463 (N_7463,N_7044,N_6950);
and U7464 (N_7464,N_7195,N_6856);
nand U7465 (N_7465,N_7126,N_6916);
and U7466 (N_7466,N_7039,N_6862);
nor U7467 (N_7467,N_6909,N_6911);
or U7468 (N_7468,N_7198,N_7109);
xor U7469 (N_7469,N_6808,N_7030);
and U7470 (N_7470,N_6909,N_6856);
and U7471 (N_7471,N_7029,N_6850);
or U7472 (N_7472,N_7026,N_6942);
nand U7473 (N_7473,N_6980,N_6859);
nor U7474 (N_7474,N_6933,N_6943);
xor U7475 (N_7475,N_6872,N_6834);
and U7476 (N_7476,N_7087,N_6964);
or U7477 (N_7477,N_7159,N_6806);
nand U7478 (N_7478,N_6827,N_7111);
or U7479 (N_7479,N_7182,N_7002);
xnor U7480 (N_7480,N_6801,N_6996);
or U7481 (N_7481,N_7180,N_7075);
nor U7482 (N_7482,N_7056,N_7073);
and U7483 (N_7483,N_7105,N_6970);
or U7484 (N_7484,N_6805,N_6924);
or U7485 (N_7485,N_7190,N_7099);
nor U7486 (N_7486,N_7192,N_7144);
nand U7487 (N_7487,N_6969,N_6858);
xnor U7488 (N_7488,N_6991,N_6969);
nand U7489 (N_7489,N_7124,N_6878);
nand U7490 (N_7490,N_6927,N_7059);
and U7491 (N_7491,N_7174,N_7038);
nand U7492 (N_7492,N_7037,N_7182);
nor U7493 (N_7493,N_6980,N_6849);
nand U7494 (N_7494,N_7131,N_7077);
xnor U7495 (N_7495,N_7131,N_6929);
nor U7496 (N_7496,N_6833,N_6898);
or U7497 (N_7497,N_6985,N_7173);
or U7498 (N_7498,N_6864,N_7162);
and U7499 (N_7499,N_7112,N_7129);
or U7500 (N_7500,N_6949,N_6913);
nor U7501 (N_7501,N_6995,N_6979);
or U7502 (N_7502,N_7120,N_6879);
nor U7503 (N_7503,N_6851,N_6856);
xnor U7504 (N_7504,N_7082,N_7100);
and U7505 (N_7505,N_6832,N_7021);
nor U7506 (N_7506,N_7056,N_6902);
nand U7507 (N_7507,N_7038,N_6858);
xor U7508 (N_7508,N_6998,N_6853);
or U7509 (N_7509,N_6978,N_6949);
and U7510 (N_7510,N_7153,N_7166);
xnor U7511 (N_7511,N_7194,N_6983);
nor U7512 (N_7512,N_6992,N_6913);
and U7513 (N_7513,N_7162,N_7169);
nand U7514 (N_7514,N_7197,N_6892);
nand U7515 (N_7515,N_7070,N_7057);
and U7516 (N_7516,N_6897,N_7178);
and U7517 (N_7517,N_7190,N_6990);
xnor U7518 (N_7518,N_6976,N_6942);
nor U7519 (N_7519,N_6828,N_6824);
nor U7520 (N_7520,N_7000,N_6955);
nand U7521 (N_7521,N_6930,N_7117);
nor U7522 (N_7522,N_7039,N_7175);
or U7523 (N_7523,N_7056,N_6893);
nand U7524 (N_7524,N_7056,N_6944);
nor U7525 (N_7525,N_6864,N_7033);
xor U7526 (N_7526,N_7128,N_7137);
xnor U7527 (N_7527,N_7062,N_7167);
or U7528 (N_7528,N_6936,N_7159);
xnor U7529 (N_7529,N_6816,N_7015);
xor U7530 (N_7530,N_7092,N_7001);
xnor U7531 (N_7531,N_6912,N_7062);
xor U7532 (N_7532,N_7030,N_7061);
and U7533 (N_7533,N_6881,N_6923);
xnor U7534 (N_7534,N_7188,N_6804);
xnor U7535 (N_7535,N_6966,N_7005);
and U7536 (N_7536,N_7008,N_6951);
nand U7537 (N_7537,N_7090,N_6807);
or U7538 (N_7538,N_6894,N_6947);
nor U7539 (N_7539,N_7180,N_6986);
xnor U7540 (N_7540,N_6900,N_7008);
nand U7541 (N_7541,N_6887,N_6877);
nor U7542 (N_7542,N_6859,N_7102);
nand U7543 (N_7543,N_6999,N_6805);
nor U7544 (N_7544,N_7083,N_7082);
xor U7545 (N_7545,N_7140,N_6954);
and U7546 (N_7546,N_7142,N_7034);
nand U7547 (N_7547,N_7119,N_6975);
and U7548 (N_7548,N_6806,N_7119);
or U7549 (N_7549,N_7197,N_7170);
nor U7550 (N_7550,N_7125,N_7070);
or U7551 (N_7551,N_7098,N_6833);
or U7552 (N_7552,N_6901,N_6928);
or U7553 (N_7553,N_6917,N_6950);
or U7554 (N_7554,N_7046,N_7069);
nor U7555 (N_7555,N_6814,N_6993);
nand U7556 (N_7556,N_6907,N_6934);
nor U7557 (N_7557,N_7136,N_7125);
xnor U7558 (N_7558,N_7115,N_7147);
or U7559 (N_7559,N_6845,N_7032);
and U7560 (N_7560,N_6959,N_7074);
nand U7561 (N_7561,N_7082,N_7108);
and U7562 (N_7562,N_7174,N_6828);
nor U7563 (N_7563,N_6846,N_6831);
nor U7564 (N_7564,N_6993,N_6849);
xnor U7565 (N_7565,N_7148,N_6848);
xnor U7566 (N_7566,N_7094,N_7111);
or U7567 (N_7567,N_6942,N_7195);
nor U7568 (N_7568,N_6856,N_6971);
nor U7569 (N_7569,N_7031,N_6814);
or U7570 (N_7570,N_7096,N_7056);
or U7571 (N_7571,N_7139,N_6985);
nand U7572 (N_7572,N_6989,N_7097);
or U7573 (N_7573,N_6903,N_6812);
xnor U7574 (N_7574,N_7083,N_7038);
nand U7575 (N_7575,N_6963,N_6958);
xor U7576 (N_7576,N_7146,N_6847);
xnor U7577 (N_7577,N_7107,N_7094);
nor U7578 (N_7578,N_7046,N_7056);
and U7579 (N_7579,N_6978,N_7121);
xor U7580 (N_7580,N_7138,N_6859);
nor U7581 (N_7581,N_7112,N_7011);
nand U7582 (N_7582,N_7170,N_6921);
nor U7583 (N_7583,N_7182,N_7110);
and U7584 (N_7584,N_6981,N_7178);
or U7585 (N_7585,N_7033,N_7095);
or U7586 (N_7586,N_7032,N_7002);
nor U7587 (N_7587,N_6937,N_7008);
nand U7588 (N_7588,N_7079,N_6815);
xor U7589 (N_7589,N_7144,N_7028);
and U7590 (N_7590,N_6857,N_6881);
nand U7591 (N_7591,N_7169,N_7060);
and U7592 (N_7592,N_7170,N_7169);
and U7593 (N_7593,N_7160,N_7072);
nand U7594 (N_7594,N_7034,N_6884);
and U7595 (N_7595,N_6809,N_6914);
nand U7596 (N_7596,N_7019,N_6834);
xor U7597 (N_7597,N_6824,N_7053);
or U7598 (N_7598,N_7073,N_7002);
nor U7599 (N_7599,N_6907,N_6891);
nand U7600 (N_7600,N_7235,N_7553);
nor U7601 (N_7601,N_7231,N_7323);
and U7602 (N_7602,N_7367,N_7356);
or U7603 (N_7603,N_7426,N_7513);
nand U7604 (N_7604,N_7423,N_7436);
nand U7605 (N_7605,N_7392,N_7437);
nand U7606 (N_7606,N_7237,N_7422);
nor U7607 (N_7607,N_7307,N_7289);
nand U7608 (N_7608,N_7345,N_7523);
nor U7609 (N_7609,N_7252,N_7308);
or U7610 (N_7610,N_7270,N_7201);
nor U7611 (N_7611,N_7324,N_7229);
or U7612 (N_7612,N_7240,N_7226);
nand U7613 (N_7613,N_7203,N_7512);
and U7614 (N_7614,N_7561,N_7468);
or U7615 (N_7615,N_7511,N_7532);
nand U7616 (N_7616,N_7469,N_7258);
and U7617 (N_7617,N_7293,N_7204);
or U7618 (N_7618,N_7350,N_7221);
or U7619 (N_7619,N_7453,N_7597);
and U7620 (N_7620,N_7537,N_7244);
xor U7621 (N_7621,N_7260,N_7488);
nor U7622 (N_7622,N_7373,N_7554);
and U7623 (N_7623,N_7388,N_7556);
nand U7624 (N_7624,N_7572,N_7533);
or U7625 (N_7625,N_7444,N_7310);
xor U7626 (N_7626,N_7410,N_7216);
and U7627 (N_7627,N_7520,N_7263);
nor U7628 (N_7628,N_7313,N_7588);
nand U7629 (N_7629,N_7344,N_7591);
xor U7630 (N_7630,N_7218,N_7342);
nor U7631 (N_7631,N_7247,N_7215);
xnor U7632 (N_7632,N_7476,N_7220);
nor U7633 (N_7633,N_7578,N_7355);
and U7634 (N_7634,N_7301,N_7517);
or U7635 (N_7635,N_7570,N_7208);
nand U7636 (N_7636,N_7489,N_7278);
and U7637 (N_7637,N_7546,N_7411);
nor U7638 (N_7638,N_7299,N_7227);
xor U7639 (N_7639,N_7306,N_7526);
or U7640 (N_7640,N_7292,N_7239);
and U7641 (N_7641,N_7321,N_7459);
nand U7642 (N_7642,N_7399,N_7507);
nand U7643 (N_7643,N_7274,N_7465);
nor U7644 (N_7644,N_7575,N_7398);
nor U7645 (N_7645,N_7331,N_7395);
and U7646 (N_7646,N_7212,N_7294);
xnor U7647 (N_7647,N_7508,N_7416);
nor U7648 (N_7648,N_7234,N_7431);
nand U7649 (N_7649,N_7418,N_7491);
and U7650 (N_7650,N_7576,N_7349);
or U7651 (N_7651,N_7277,N_7592);
and U7652 (N_7652,N_7412,N_7475);
xor U7653 (N_7653,N_7383,N_7358);
xnor U7654 (N_7654,N_7343,N_7389);
nand U7655 (N_7655,N_7429,N_7400);
nand U7656 (N_7656,N_7364,N_7456);
nor U7657 (N_7657,N_7385,N_7320);
and U7658 (N_7658,N_7518,N_7376);
nor U7659 (N_7659,N_7460,N_7405);
xor U7660 (N_7660,N_7454,N_7473);
or U7661 (N_7661,N_7354,N_7505);
and U7662 (N_7662,N_7413,N_7565);
or U7663 (N_7663,N_7580,N_7497);
xnor U7664 (N_7664,N_7503,N_7315);
or U7665 (N_7665,N_7291,N_7573);
or U7666 (N_7666,N_7363,N_7581);
xnor U7667 (N_7667,N_7433,N_7598);
nor U7668 (N_7668,N_7567,N_7595);
nand U7669 (N_7669,N_7304,N_7485);
nand U7670 (N_7670,N_7443,N_7377);
or U7671 (N_7671,N_7256,N_7357);
and U7672 (N_7672,N_7280,N_7547);
nor U7673 (N_7673,N_7255,N_7519);
nand U7674 (N_7674,N_7434,N_7266);
nand U7675 (N_7675,N_7467,N_7502);
or U7676 (N_7676,N_7368,N_7309);
nor U7677 (N_7677,N_7494,N_7415);
or U7678 (N_7678,N_7326,N_7482);
or U7679 (N_7679,N_7574,N_7387);
or U7680 (N_7680,N_7528,N_7250);
or U7681 (N_7681,N_7259,N_7448);
nor U7682 (N_7682,N_7288,N_7243);
and U7683 (N_7683,N_7550,N_7365);
nand U7684 (N_7684,N_7439,N_7462);
nand U7685 (N_7685,N_7312,N_7285);
nand U7686 (N_7686,N_7539,N_7351);
or U7687 (N_7687,N_7262,N_7427);
and U7688 (N_7688,N_7224,N_7269);
xnor U7689 (N_7689,N_7457,N_7481);
nand U7690 (N_7690,N_7441,N_7340);
xor U7691 (N_7691,N_7295,N_7402);
xnor U7692 (N_7692,N_7557,N_7361);
nand U7693 (N_7693,N_7219,N_7401);
xnor U7694 (N_7694,N_7381,N_7425);
nand U7695 (N_7695,N_7500,N_7586);
nor U7696 (N_7696,N_7571,N_7286);
nor U7697 (N_7697,N_7534,N_7463);
nand U7698 (N_7698,N_7577,N_7330);
or U7699 (N_7699,N_7596,N_7509);
xnor U7700 (N_7700,N_7372,N_7371);
or U7701 (N_7701,N_7551,N_7391);
nor U7702 (N_7702,N_7380,N_7296);
or U7703 (N_7703,N_7562,N_7558);
nand U7704 (N_7704,N_7375,N_7382);
nand U7705 (N_7705,N_7404,N_7353);
nand U7706 (N_7706,N_7272,N_7408);
nand U7707 (N_7707,N_7303,N_7492);
xor U7708 (N_7708,N_7257,N_7442);
or U7709 (N_7709,N_7341,N_7403);
nor U7710 (N_7710,N_7450,N_7348);
nand U7711 (N_7711,N_7446,N_7200);
nor U7712 (N_7712,N_7435,N_7214);
xor U7713 (N_7713,N_7594,N_7287);
xnor U7714 (N_7714,N_7318,N_7245);
xnor U7715 (N_7715,N_7205,N_7420);
nor U7716 (N_7716,N_7322,N_7516);
or U7717 (N_7717,N_7440,N_7522);
and U7718 (N_7718,N_7535,N_7529);
or U7719 (N_7719,N_7267,N_7332);
and U7720 (N_7720,N_7360,N_7569);
xor U7721 (N_7721,N_7386,N_7560);
or U7722 (N_7722,N_7328,N_7228);
nand U7723 (N_7723,N_7384,N_7559);
nand U7724 (N_7724,N_7568,N_7447);
or U7725 (N_7725,N_7406,N_7514);
nand U7726 (N_7726,N_7396,N_7589);
and U7727 (N_7727,N_7527,N_7209);
xnor U7728 (N_7728,N_7236,N_7338);
or U7729 (N_7729,N_7233,N_7282);
xor U7730 (N_7730,N_7499,N_7223);
nor U7731 (N_7731,N_7487,N_7261);
and U7732 (N_7732,N_7207,N_7495);
nor U7733 (N_7733,N_7417,N_7333);
and U7734 (N_7734,N_7300,N_7541);
xor U7735 (N_7735,N_7584,N_7249);
nor U7736 (N_7736,N_7335,N_7311);
nand U7737 (N_7737,N_7248,N_7544);
or U7738 (N_7738,N_7316,N_7297);
and U7739 (N_7739,N_7471,N_7419);
xnor U7740 (N_7740,N_7397,N_7302);
and U7741 (N_7741,N_7232,N_7202);
and U7742 (N_7742,N_7409,N_7524);
nor U7743 (N_7743,N_7347,N_7521);
nand U7744 (N_7744,N_7501,N_7414);
or U7745 (N_7745,N_7472,N_7504);
nand U7746 (N_7746,N_7251,N_7336);
xnor U7747 (N_7747,N_7271,N_7370);
nand U7748 (N_7748,N_7477,N_7536);
nor U7749 (N_7749,N_7362,N_7479);
xnor U7750 (N_7750,N_7531,N_7464);
and U7751 (N_7751,N_7242,N_7254);
or U7752 (N_7752,N_7552,N_7359);
or U7753 (N_7753,N_7268,N_7390);
and U7754 (N_7754,N_7430,N_7298);
and U7755 (N_7755,N_7253,N_7498);
xnor U7756 (N_7756,N_7545,N_7455);
nor U7757 (N_7757,N_7379,N_7238);
or U7758 (N_7758,N_7325,N_7276);
and U7759 (N_7759,N_7407,N_7466);
nor U7760 (N_7760,N_7225,N_7540);
xor U7761 (N_7761,N_7555,N_7421);
nand U7762 (N_7762,N_7337,N_7493);
and U7763 (N_7763,N_7478,N_7566);
nand U7764 (N_7764,N_7525,N_7538);
nand U7765 (N_7765,N_7366,N_7530);
nand U7766 (N_7766,N_7275,N_7583);
or U7767 (N_7767,N_7486,N_7563);
nand U7768 (N_7768,N_7281,N_7549);
or U7769 (N_7769,N_7438,N_7327);
or U7770 (N_7770,N_7374,N_7461);
xnor U7771 (N_7771,N_7394,N_7548);
and U7772 (N_7772,N_7480,N_7585);
or U7773 (N_7773,N_7515,N_7496);
xnor U7774 (N_7774,N_7339,N_7279);
nand U7775 (N_7775,N_7564,N_7470);
and U7776 (N_7776,N_7542,N_7305);
nand U7777 (N_7777,N_7369,N_7329);
nor U7778 (N_7778,N_7428,N_7424);
nor U7779 (N_7779,N_7432,N_7284);
nand U7780 (N_7780,N_7246,N_7314);
nor U7781 (N_7781,N_7599,N_7290);
nor U7782 (N_7782,N_7273,N_7230);
nor U7783 (N_7783,N_7452,N_7317);
or U7784 (N_7784,N_7346,N_7211);
xnor U7785 (N_7785,N_7490,N_7213);
or U7786 (N_7786,N_7483,N_7445);
nor U7787 (N_7787,N_7449,N_7451);
or U7788 (N_7788,N_7283,N_7510);
and U7789 (N_7789,N_7210,N_7458);
and U7790 (N_7790,N_7319,N_7593);
nand U7791 (N_7791,N_7241,N_7264);
nor U7792 (N_7792,N_7582,N_7378);
nand U7793 (N_7793,N_7334,N_7265);
nor U7794 (N_7794,N_7206,N_7393);
or U7795 (N_7795,N_7217,N_7590);
and U7796 (N_7796,N_7587,N_7474);
nor U7797 (N_7797,N_7484,N_7543);
xor U7798 (N_7798,N_7352,N_7222);
nand U7799 (N_7799,N_7506,N_7579);
and U7800 (N_7800,N_7404,N_7200);
and U7801 (N_7801,N_7436,N_7414);
nand U7802 (N_7802,N_7505,N_7214);
nor U7803 (N_7803,N_7441,N_7507);
or U7804 (N_7804,N_7226,N_7382);
nor U7805 (N_7805,N_7524,N_7463);
nor U7806 (N_7806,N_7563,N_7368);
nor U7807 (N_7807,N_7550,N_7372);
xnor U7808 (N_7808,N_7327,N_7550);
or U7809 (N_7809,N_7533,N_7304);
nor U7810 (N_7810,N_7416,N_7361);
xnor U7811 (N_7811,N_7591,N_7373);
or U7812 (N_7812,N_7309,N_7593);
or U7813 (N_7813,N_7235,N_7519);
and U7814 (N_7814,N_7406,N_7569);
or U7815 (N_7815,N_7433,N_7312);
nand U7816 (N_7816,N_7583,N_7435);
xor U7817 (N_7817,N_7503,N_7332);
xor U7818 (N_7818,N_7562,N_7481);
or U7819 (N_7819,N_7375,N_7493);
or U7820 (N_7820,N_7363,N_7541);
xnor U7821 (N_7821,N_7350,N_7535);
or U7822 (N_7822,N_7222,N_7240);
nand U7823 (N_7823,N_7594,N_7357);
nor U7824 (N_7824,N_7513,N_7596);
xor U7825 (N_7825,N_7590,N_7465);
nand U7826 (N_7826,N_7269,N_7417);
nand U7827 (N_7827,N_7283,N_7516);
and U7828 (N_7828,N_7360,N_7236);
and U7829 (N_7829,N_7581,N_7574);
or U7830 (N_7830,N_7419,N_7573);
and U7831 (N_7831,N_7241,N_7360);
and U7832 (N_7832,N_7428,N_7550);
nand U7833 (N_7833,N_7314,N_7300);
and U7834 (N_7834,N_7363,N_7347);
nor U7835 (N_7835,N_7316,N_7299);
nand U7836 (N_7836,N_7205,N_7397);
and U7837 (N_7837,N_7505,N_7523);
xnor U7838 (N_7838,N_7402,N_7292);
xnor U7839 (N_7839,N_7266,N_7345);
nor U7840 (N_7840,N_7250,N_7234);
nor U7841 (N_7841,N_7487,N_7412);
nand U7842 (N_7842,N_7426,N_7333);
nand U7843 (N_7843,N_7599,N_7324);
xor U7844 (N_7844,N_7585,N_7200);
nor U7845 (N_7845,N_7560,N_7385);
nand U7846 (N_7846,N_7416,N_7203);
or U7847 (N_7847,N_7562,N_7280);
or U7848 (N_7848,N_7360,N_7599);
and U7849 (N_7849,N_7262,N_7398);
xor U7850 (N_7850,N_7471,N_7279);
or U7851 (N_7851,N_7356,N_7469);
or U7852 (N_7852,N_7305,N_7586);
or U7853 (N_7853,N_7364,N_7503);
or U7854 (N_7854,N_7401,N_7438);
and U7855 (N_7855,N_7369,N_7485);
xnor U7856 (N_7856,N_7276,N_7547);
xnor U7857 (N_7857,N_7272,N_7258);
nor U7858 (N_7858,N_7580,N_7212);
xnor U7859 (N_7859,N_7219,N_7204);
nor U7860 (N_7860,N_7504,N_7271);
nand U7861 (N_7861,N_7480,N_7305);
and U7862 (N_7862,N_7578,N_7308);
or U7863 (N_7863,N_7382,N_7440);
xnor U7864 (N_7864,N_7391,N_7502);
nand U7865 (N_7865,N_7433,N_7531);
nand U7866 (N_7866,N_7460,N_7215);
nand U7867 (N_7867,N_7396,N_7249);
xnor U7868 (N_7868,N_7401,N_7265);
xnor U7869 (N_7869,N_7253,N_7460);
nor U7870 (N_7870,N_7227,N_7212);
or U7871 (N_7871,N_7511,N_7445);
or U7872 (N_7872,N_7424,N_7577);
nor U7873 (N_7873,N_7424,N_7458);
nor U7874 (N_7874,N_7293,N_7524);
nand U7875 (N_7875,N_7572,N_7389);
nand U7876 (N_7876,N_7313,N_7492);
or U7877 (N_7877,N_7271,N_7528);
nor U7878 (N_7878,N_7466,N_7455);
nand U7879 (N_7879,N_7405,N_7324);
xor U7880 (N_7880,N_7448,N_7353);
nor U7881 (N_7881,N_7258,N_7531);
and U7882 (N_7882,N_7319,N_7254);
nor U7883 (N_7883,N_7388,N_7412);
and U7884 (N_7884,N_7355,N_7544);
xnor U7885 (N_7885,N_7511,N_7381);
xor U7886 (N_7886,N_7561,N_7591);
nor U7887 (N_7887,N_7546,N_7486);
or U7888 (N_7888,N_7571,N_7300);
xor U7889 (N_7889,N_7549,N_7222);
xor U7890 (N_7890,N_7409,N_7276);
xor U7891 (N_7891,N_7520,N_7436);
or U7892 (N_7892,N_7532,N_7450);
or U7893 (N_7893,N_7247,N_7310);
nand U7894 (N_7894,N_7367,N_7236);
or U7895 (N_7895,N_7349,N_7511);
or U7896 (N_7896,N_7344,N_7228);
and U7897 (N_7897,N_7270,N_7324);
nor U7898 (N_7898,N_7541,N_7446);
xor U7899 (N_7899,N_7472,N_7577);
or U7900 (N_7900,N_7597,N_7334);
nor U7901 (N_7901,N_7597,N_7560);
and U7902 (N_7902,N_7370,N_7399);
or U7903 (N_7903,N_7296,N_7522);
or U7904 (N_7904,N_7371,N_7252);
and U7905 (N_7905,N_7296,N_7531);
and U7906 (N_7906,N_7437,N_7427);
nor U7907 (N_7907,N_7510,N_7242);
xnor U7908 (N_7908,N_7583,N_7205);
nor U7909 (N_7909,N_7369,N_7298);
nand U7910 (N_7910,N_7481,N_7243);
xor U7911 (N_7911,N_7417,N_7423);
or U7912 (N_7912,N_7419,N_7578);
nand U7913 (N_7913,N_7586,N_7445);
nor U7914 (N_7914,N_7577,N_7220);
nor U7915 (N_7915,N_7282,N_7401);
nor U7916 (N_7916,N_7332,N_7323);
or U7917 (N_7917,N_7451,N_7377);
or U7918 (N_7918,N_7553,N_7207);
and U7919 (N_7919,N_7302,N_7538);
xnor U7920 (N_7920,N_7453,N_7273);
and U7921 (N_7921,N_7585,N_7370);
or U7922 (N_7922,N_7296,N_7340);
nand U7923 (N_7923,N_7352,N_7457);
nand U7924 (N_7924,N_7412,N_7285);
nand U7925 (N_7925,N_7388,N_7598);
or U7926 (N_7926,N_7267,N_7249);
nor U7927 (N_7927,N_7295,N_7403);
nor U7928 (N_7928,N_7235,N_7272);
nand U7929 (N_7929,N_7334,N_7416);
nand U7930 (N_7930,N_7326,N_7478);
and U7931 (N_7931,N_7528,N_7261);
or U7932 (N_7932,N_7348,N_7431);
or U7933 (N_7933,N_7449,N_7420);
and U7934 (N_7934,N_7328,N_7428);
nand U7935 (N_7935,N_7323,N_7279);
or U7936 (N_7936,N_7551,N_7445);
nor U7937 (N_7937,N_7430,N_7510);
nand U7938 (N_7938,N_7595,N_7570);
xnor U7939 (N_7939,N_7218,N_7221);
nor U7940 (N_7940,N_7460,N_7572);
and U7941 (N_7941,N_7396,N_7564);
xnor U7942 (N_7942,N_7593,N_7388);
and U7943 (N_7943,N_7417,N_7405);
nand U7944 (N_7944,N_7242,N_7441);
xor U7945 (N_7945,N_7501,N_7443);
nand U7946 (N_7946,N_7373,N_7599);
nand U7947 (N_7947,N_7403,N_7549);
and U7948 (N_7948,N_7530,N_7511);
and U7949 (N_7949,N_7232,N_7511);
and U7950 (N_7950,N_7483,N_7560);
xor U7951 (N_7951,N_7410,N_7432);
nor U7952 (N_7952,N_7472,N_7546);
xor U7953 (N_7953,N_7324,N_7377);
nor U7954 (N_7954,N_7567,N_7327);
nor U7955 (N_7955,N_7463,N_7283);
nand U7956 (N_7956,N_7548,N_7472);
and U7957 (N_7957,N_7598,N_7386);
nor U7958 (N_7958,N_7471,N_7336);
xor U7959 (N_7959,N_7210,N_7407);
xor U7960 (N_7960,N_7476,N_7430);
xnor U7961 (N_7961,N_7572,N_7530);
xor U7962 (N_7962,N_7542,N_7407);
nand U7963 (N_7963,N_7327,N_7201);
and U7964 (N_7964,N_7516,N_7511);
nor U7965 (N_7965,N_7210,N_7262);
nor U7966 (N_7966,N_7327,N_7472);
and U7967 (N_7967,N_7509,N_7299);
and U7968 (N_7968,N_7568,N_7369);
xnor U7969 (N_7969,N_7520,N_7356);
or U7970 (N_7970,N_7540,N_7238);
nand U7971 (N_7971,N_7206,N_7418);
xnor U7972 (N_7972,N_7501,N_7449);
nand U7973 (N_7973,N_7390,N_7566);
nor U7974 (N_7974,N_7508,N_7279);
or U7975 (N_7975,N_7444,N_7504);
xor U7976 (N_7976,N_7392,N_7363);
and U7977 (N_7977,N_7517,N_7263);
and U7978 (N_7978,N_7363,N_7368);
or U7979 (N_7979,N_7590,N_7595);
xor U7980 (N_7980,N_7217,N_7277);
nand U7981 (N_7981,N_7245,N_7444);
and U7982 (N_7982,N_7277,N_7361);
xor U7983 (N_7983,N_7211,N_7364);
nand U7984 (N_7984,N_7481,N_7415);
and U7985 (N_7985,N_7252,N_7234);
nor U7986 (N_7986,N_7303,N_7265);
nor U7987 (N_7987,N_7528,N_7512);
and U7988 (N_7988,N_7234,N_7255);
or U7989 (N_7989,N_7417,N_7252);
and U7990 (N_7990,N_7448,N_7485);
nand U7991 (N_7991,N_7329,N_7588);
and U7992 (N_7992,N_7479,N_7518);
or U7993 (N_7993,N_7421,N_7298);
xor U7994 (N_7994,N_7216,N_7445);
nand U7995 (N_7995,N_7532,N_7454);
xor U7996 (N_7996,N_7309,N_7433);
and U7997 (N_7997,N_7257,N_7520);
and U7998 (N_7998,N_7257,N_7212);
xnor U7999 (N_7999,N_7355,N_7472);
and U8000 (N_8000,N_7723,N_7825);
xor U8001 (N_8001,N_7979,N_7679);
nor U8002 (N_8002,N_7711,N_7603);
nand U8003 (N_8003,N_7782,N_7929);
xnor U8004 (N_8004,N_7856,N_7790);
nor U8005 (N_8005,N_7738,N_7671);
nand U8006 (N_8006,N_7718,N_7962);
nand U8007 (N_8007,N_7885,N_7713);
and U8008 (N_8008,N_7997,N_7984);
and U8009 (N_8009,N_7892,N_7708);
nor U8010 (N_8010,N_7608,N_7647);
and U8011 (N_8011,N_7677,N_7755);
or U8012 (N_8012,N_7801,N_7833);
nand U8013 (N_8013,N_7682,N_7897);
or U8014 (N_8014,N_7604,N_7800);
xor U8015 (N_8015,N_7823,N_7687);
or U8016 (N_8016,N_7748,N_7891);
nand U8017 (N_8017,N_7803,N_7638);
nand U8018 (N_8018,N_7784,N_7743);
and U8019 (N_8019,N_7927,N_7868);
nand U8020 (N_8020,N_7781,N_7881);
nor U8021 (N_8021,N_7910,N_7642);
xnor U8022 (N_8022,N_7923,N_7889);
nor U8023 (N_8023,N_7834,N_7786);
nor U8024 (N_8024,N_7996,N_7643);
nand U8025 (N_8025,N_7683,N_7785);
nor U8026 (N_8026,N_7837,N_7886);
nand U8027 (N_8027,N_7623,N_7982);
xnor U8028 (N_8028,N_7920,N_7884);
xnor U8029 (N_8029,N_7731,N_7940);
and U8030 (N_8030,N_7878,N_7795);
and U8031 (N_8031,N_7936,N_7760);
or U8032 (N_8032,N_7694,N_7972);
xor U8033 (N_8033,N_7717,N_7930);
and U8034 (N_8034,N_7690,N_7859);
xnor U8035 (N_8035,N_7955,N_7953);
nor U8036 (N_8036,N_7890,N_7775);
xor U8037 (N_8037,N_7975,N_7816);
xnor U8038 (N_8038,N_7753,N_7880);
or U8039 (N_8039,N_7756,N_7733);
nor U8040 (N_8040,N_7635,N_7978);
xnor U8041 (N_8041,N_7624,N_7814);
nor U8042 (N_8042,N_7895,N_7999);
nor U8043 (N_8043,N_7968,N_7605);
and U8044 (N_8044,N_7698,N_7865);
xor U8045 (N_8045,N_7872,N_7609);
and U8046 (N_8046,N_7970,N_7796);
nand U8047 (N_8047,N_7668,N_7934);
nand U8048 (N_8048,N_7730,N_7870);
or U8049 (N_8049,N_7966,N_7893);
or U8050 (N_8050,N_7692,N_7649);
xor U8051 (N_8051,N_7805,N_7774);
xor U8052 (N_8052,N_7697,N_7854);
nor U8053 (N_8053,N_7792,N_7722);
and U8054 (N_8054,N_7744,N_7862);
nand U8055 (N_8055,N_7621,N_7974);
and U8056 (N_8056,N_7848,N_7704);
xnor U8057 (N_8057,N_7830,N_7611);
nand U8058 (N_8058,N_7648,N_7826);
xor U8059 (N_8059,N_7813,N_7663);
xnor U8060 (N_8060,N_7933,N_7625);
nor U8061 (N_8061,N_7860,N_7684);
and U8062 (N_8062,N_7701,N_7789);
nor U8063 (N_8063,N_7778,N_7678);
nor U8064 (N_8064,N_7850,N_7858);
nand U8065 (N_8065,N_7939,N_7739);
nand U8066 (N_8066,N_7991,N_7742);
nand U8067 (N_8067,N_7685,N_7922);
and U8068 (N_8068,N_7716,N_7772);
nor U8069 (N_8069,N_7729,N_7700);
and U8070 (N_8070,N_7846,N_7644);
or U8071 (N_8071,N_7720,N_7757);
nor U8072 (N_8072,N_7610,N_7981);
and U8073 (N_8073,N_7691,N_7740);
or U8074 (N_8074,N_7659,N_7899);
nor U8075 (N_8075,N_7693,N_7932);
and U8076 (N_8076,N_7942,N_7925);
nor U8077 (N_8077,N_7627,N_7606);
xnor U8078 (N_8078,N_7797,N_7959);
nor U8079 (N_8079,N_7902,N_7900);
nand U8080 (N_8080,N_7873,N_7667);
and U8081 (N_8081,N_7946,N_7791);
or U8082 (N_8082,N_7799,N_7887);
and U8083 (N_8083,N_7958,N_7702);
xnor U8084 (N_8084,N_7749,N_7907);
xnor U8085 (N_8085,N_7909,N_7807);
and U8086 (N_8086,N_7793,N_7646);
nand U8087 (N_8087,N_7613,N_7783);
or U8088 (N_8088,N_7812,N_7787);
nand U8089 (N_8089,N_7954,N_7629);
nor U8090 (N_8090,N_7804,N_7802);
and U8091 (N_8091,N_7737,N_7607);
nand U8092 (N_8092,N_7620,N_7715);
and U8093 (N_8093,N_7827,N_7709);
nand U8094 (N_8094,N_7819,N_7714);
nor U8095 (N_8095,N_7965,N_7998);
nand U8096 (N_8096,N_7948,N_7669);
xnor U8097 (N_8097,N_7969,N_7650);
nand U8098 (N_8098,N_7768,N_7658);
and U8099 (N_8099,N_7822,N_7957);
xnor U8100 (N_8100,N_7634,N_7896);
and U8101 (N_8101,N_7911,N_7645);
nand U8102 (N_8102,N_7831,N_7874);
nand U8103 (N_8103,N_7908,N_7943);
xnor U8104 (N_8104,N_7844,N_7655);
nor U8105 (N_8105,N_7843,N_7780);
nor U8106 (N_8106,N_7689,N_7990);
xnor U8107 (N_8107,N_7765,N_7828);
and U8108 (N_8108,N_7836,N_7817);
xnor U8109 (N_8109,N_7675,N_7994);
and U8110 (N_8110,N_7935,N_7806);
and U8111 (N_8111,N_7602,N_7882);
nor U8112 (N_8112,N_7747,N_7761);
xor U8113 (N_8113,N_7937,N_7905);
xor U8114 (N_8114,N_7986,N_7861);
or U8115 (N_8115,N_7764,N_7852);
or U8116 (N_8116,N_7754,N_7773);
nor U8117 (N_8117,N_7995,N_7724);
and U8118 (N_8118,N_7662,N_7815);
or U8119 (N_8119,N_7988,N_7630);
and U8120 (N_8120,N_7867,N_7980);
xnor U8121 (N_8121,N_7849,N_7601);
nor U8122 (N_8122,N_7695,N_7651);
or U8123 (N_8123,N_7736,N_7766);
xor U8124 (N_8124,N_7652,N_7788);
or U8125 (N_8125,N_7759,N_7866);
nor U8126 (N_8126,N_7632,N_7863);
nor U8127 (N_8127,N_7829,N_7924);
nand U8128 (N_8128,N_7944,N_7672);
xor U8129 (N_8129,N_7973,N_7912);
xnor U8130 (N_8130,N_7762,N_7769);
and U8131 (N_8131,N_7853,N_7931);
nor U8132 (N_8132,N_7732,N_7660);
nor U8133 (N_8133,N_7707,N_7915);
xnor U8134 (N_8134,N_7776,N_7661);
or U8135 (N_8135,N_7735,N_7626);
and U8136 (N_8136,N_7993,N_7810);
nor U8137 (N_8137,N_7741,N_7992);
xnor U8138 (N_8138,N_7696,N_7752);
nor U8139 (N_8139,N_7751,N_7664);
nand U8140 (N_8140,N_7951,N_7898);
or U8141 (N_8141,N_7674,N_7916);
or U8142 (N_8142,N_7839,N_7809);
nand U8143 (N_8143,N_7851,N_7628);
nand U8144 (N_8144,N_7964,N_7808);
xnor U8145 (N_8145,N_7767,N_7894);
and U8146 (N_8146,N_7838,N_7821);
xor U8147 (N_8147,N_7681,N_7727);
nand U8148 (N_8148,N_7938,N_7614);
or U8149 (N_8149,N_7726,N_7619);
nor U8150 (N_8150,N_7639,N_7875);
xor U8151 (N_8151,N_7676,N_7616);
nor U8152 (N_8152,N_7928,N_7631);
and U8153 (N_8153,N_7670,N_7949);
xnor U8154 (N_8154,N_7705,N_7921);
xnor U8155 (N_8155,N_7857,N_7941);
xnor U8156 (N_8156,N_7734,N_7869);
nor U8157 (N_8157,N_7706,N_7721);
nand U8158 (N_8158,N_7798,N_7947);
nand U8159 (N_8159,N_7841,N_7612);
nand U8160 (N_8160,N_7855,N_7967);
xor U8161 (N_8161,N_7703,N_7710);
nand U8162 (N_8162,N_7904,N_7976);
and U8163 (N_8163,N_7901,N_7840);
or U8164 (N_8164,N_7641,N_7985);
nand U8165 (N_8165,N_7615,N_7914);
nand U8166 (N_8166,N_7811,N_7794);
nor U8167 (N_8167,N_7637,N_7725);
xnor U8168 (N_8168,N_7983,N_7926);
nand U8169 (N_8169,N_7820,N_7845);
nor U8170 (N_8170,N_7903,N_7745);
or U8171 (N_8171,N_7871,N_7917);
nand U8172 (N_8172,N_7906,N_7879);
or U8173 (N_8173,N_7758,N_7956);
nor U8174 (N_8174,N_7771,N_7673);
xnor U8175 (N_8175,N_7750,N_7779);
nand U8176 (N_8176,N_7832,N_7666);
xor U8177 (N_8177,N_7763,N_7945);
and U8178 (N_8178,N_7657,N_7622);
or U8179 (N_8179,N_7971,N_7719);
nand U8180 (N_8180,N_7686,N_7699);
and U8181 (N_8181,N_7656,N_7770);
nand U8182 (N_8182,N_7876,N_7877);
nor U8183 (N_8183,N_7746,N_7864);
and U8184 (N_8184,N_7950,N_7977);
or U8185 (N_8185,N_7989,N_7777);
nand U8186 (N_8186,N_7665,N_7963);
nand U8187 (N_8187,N_7688,N_7952);
and U8188 (N_8188,N_7728,N_7918);
nor U8189 (N_8189,N_7618,N_7617);
nor U8190 (N_8190,N_7680,N_7600);
and U8191 (N_8191,N_7883,N_7653);
xnor U8192 (N_8192,N_7913,N_7961);
and U8193 (N_8193,N_7636,N_7633);
or U8194 (N_8194,N_7654,N_7712);
or U8195 (N_8195,N_7824,N_7842);
or U8196 (N_8196,N_7847,N_7835);
xnor U8197 (N_8197,N_7640,N_7987);
xor U8198 (N_8198,N_7818,N_7919);
or U8199 (N_8199,N_7888,N_7960);
or U8200 (N_8200,N_7733,N_7899);
xor U8201 (N_8201,N_7941,N_7890);
and U8202 (N_8202,N_7706,N_7971);
or U8203 (N_8203,N_7892,N_7678);
xnor U8204 (N_8204,N_7753,N_7798);
or U8205 (N_8205,N_7916,N_7601);
and U8206 (N_8206,N_7924,N_7731);
and U8207 (N_8207,N_7629,N_7636);
nand U8208 (N_8208,N_7716,N_7762);
or U8209 (N_8209,N_7705,N_7896);
or U8210 (N_8210,N_7877,N_7850);
xor U8211 (N_8211,N_7768,N_7760);
and U8212 (N_8212,N_7655,N_7704);
xor U8213 (N_8213,N_7614,N_7917);
or U8214 (N_8214,N_7874,N_7655);
and U8215 (N_8215,N_7857,N_7665);
nand U8216 (N_8216,N_7710,N_7713);
nand U8217 (N_8217,N_7830,N_7642);
nor U8218 (N_8218,N_7984,N_7610);
and U8219 (N_8219,N_7807,N_7971);
and U8220 (N_8220,N_7992,N_7936);
nand U8221 (N_8221,N_7946,N_7928);
or U8222 (N_8222,N_7993,N_7923);
and U8223 (N_8223,N_7743,N_7841);
nand U8224 (N_8224,N_7940,N_7995);
nand U8225 (N_8225,N_7775,N_7891);
nor U8226 (N_8226,N_7852,N_7636);
nor U8227 (N_8227,N_7671,N_7604);
or U8228 (N_8228,N_7842,N_7695);
xnor U8229 (N_8229,N_7643,N_7612);
and U8230 (N_8230,N_7832,N_7989);
nor U8231 (N_8231,N_7615,N_7710);
nand U8232 (N_8232,N_7641,N_7674);
or U8233 (N_8233,N_7984,N_7674);
and U8234 (N_8234,N_7618,N_7704);
and U8235 (N_8235,N_7783,N_7911);
xnor U8236 (N_8236,N_7711,N_7982);
nor U8237 (N_8237,N_7982,N_7983);
xor U8238 (N_8238,N_7682,N_7715);
nor U8239 (N_8239,N_7891,N_7872);
nor U8240 (N_8240,N_7923,N_7638);
nand U8241 (N_8241,N_7779,N_7867);
or U8242 (N_8242,N_7789,N_7992);
or U8243 (N_8243,N_7664,N_7726);
and U8244 (N_8244,N_7913,N_7969);
xor U8245 (N_8245,N_7768,N_7820);
nand U8246 (N_8246,N_7832,N_7905);
and U8247 (N_8247,N_7826,N_7807);
or U8248 (N_8248,N_7888,N_7931);
nor U8249 (N_8249,N_7964,N_7882);
nor U8250 (N_8250,N_7664,N_7962);
nand U8251 (N_8251,N_7923,N_7942);
xor U8252 (N_8252,N_7703,N_7812);
nand U8253 (N_8253,N_7870,N_7902);
or U8254 (N_8254,N_7711,N_7696);
xnor U8255 (N_8255,N_7960,N_7697);
xnor U8256 (N_8256,N_7875,N_7788);
or U8257 (N_8257,N_7696,N_7693);
xor U8258 (N_8258,N_7830,N_7750);
or U8259 (N_8259,N_7657,N_7726);
xor U8260 (N_8260,N_7604,N_7935);
nor U8261 (N_8261,N_7681,N_7750);
xnor U8262 (N_8262,N_7868,N_7616);
or U8263 (N_8263,N_7737,N_7945);
or U8264 (N_8264,N_7848,N_7724);
xnor U8265 (N_8265,N_7731,N_7981);
nor U8266 (N_8266,N_7852,N_7724);
xnor U8267 (N_8267,N_7733,N_7770);
nor U8268 (N_8268,N_7665,N_7866);
xnor U8269 (N_8269,N_7998,N_7689);
nand U8270 (N_8270,N_7739,N_7773);
nand U8271 (N_8271,N_7984,N_7926);
xnor U8272 (N_8272,N_7829,N_7950);
and U8273 (N_8273,N_7647,N_7786);
xor U8274 (N_8274,N_7697,N_7722);
nand U8275 (N_8275,N_7861,N_7928);
and U8276 (N_8276,N_7885,N_7819);
and U8277 (N_8277,N_7948,N_7809);
xor U8278 (N_8278,N_7882,N_7952);
nand U8279 (N_8279,N_7972,N_7603);
nor U8280 (N_8280,N_7897,N_7985);
nor U8281 (N_8281,N_7729,N_7908);
xnor U8282 (N_8282,N_7869,N_7601);
xnor U8283 (N_8283,N_7805,N_7995);
or U8284 (N_8284,N_7893,N_7946);
nor U8285 (N_8285,N_7864,N_7664);
or U8286 (N_8286,N_7635,N_7935);
and U8287 (N_8287,N_7613,N_7723);
or U8288 (N_8288,N_7790,N_7845);
nand U8289 (N_8289,N_7680,N_7697);
nor U8290 (N_8290,N_7769,N_7746);
nand U8291 (N_8291,N_7807,N_7952);
xor U8292 (N_8292,N_7641,N_7964);
and U8293 (N_8293,N_7878,N_7614);
nand U8294 (N_8294,N_7928,N_7765);
and U8295 (N_8295,N_7785,N_7703);
and U8296 (N_8296,N_7916,N_7611);
xnor U8297 (N_8297,N_7609,N_7801);
xnor U8298 (N_8298,N_7872,N_7840);
and U8299 (N_8299,N_7705,N_7802);
and U8300 (N_8300,N_7735,N_7877);
nor U8301 (N_8301,N_7633,N_7677);
and U8302 (N_8302,N_7755,N_7659);
nor U8303 (N_8303,N_7724,N_7632);
and U8304 (N_8304,N_7791,N_7783);
nand U8305 (N_8305,N_7921,N_7847);
xor U8306 (N_8306,N_7803,N_7872);
nand U8307 (N_8307,N_7775,N_7736);
nand U8308 (N_8308,N_7987,N_7983);
nor U8309 (N_8309,N_7650,N_7798);
nor U8310 (N_8310,N_7611,N_7863);
nor U8311 (N_8311,N_7973,N_7845);
nand U8312 (N_8312,N_7782,N_7832);
and U8313 (N_8313,N_7817,N_7847);
xnor U8314 (N_8314,N_7887,N_7860);
nand U8315 (N_8315,N_7611,N_7672);
nand U8316 (N_8316,N_7811,N_7656);
and U8317 (N_8317,N_7844,N_7944);
xnor U8318 (N_8318,N_7750,N_7664);
nand U8319 (N_8319,N_7642,N_7624);
or U8320 (N_8320,N_7970,N_7668);
nand U8321 (N_8321,N_7973,N_7873);
and U8322 (N_8322,N_7685,N_7806);
or U8323 (N_8323,N_7728,N_7687);
or U8324 (N_8324,N_7788,N_7773);
or U8325 (N_8325,N_7613,N_7897);
nand U8326 (N_8326,N_7946,N_7710);
and U8327 (N_8327,N_7704,N_7938);
nor U8328 (N_8328,N_7655,N_7678);
xor U8329 (N_8329,N_7666,N_7892);
nor U8330 (N_8330,N_7749,N_7632);
nand U8331 (N_8331,N_7948,N_7621);
and U8332 (N_8332,N_7702,N_7731);
or U8333 (N_8333,N_7685,N_7731);
and U8334 (N_8334,N_7709,N_7803);
or U8335 (N_8335,N_7949,N_7824);
or U8336 (N_8336,N_7918,N_7819);
nand U8337 (N_8337,N_7796,N_7645);
xor U8338 (N_8338,N_7729,N_7850);
and U8339 (N_8339,N_7818,N_7996);
and U8340 (N_8340,N_7877,N_7746);
nor U8341 (N_8341,N_7861,N_7660);
xor U8342 (N_8342,N_7628,N_7629);
xor U8343 (N_8343,N_7848,N_7735);
or U8344 (N_8344,N_7753,N_7736);
or U8345 (N_8345,N_7980,N_7762);
xor U8346 (N_8346,N_7819,N_7894);
nand U8347 (N_8347,N_7711,N_7632);
nand U8348 (N_8348,N_7933,N_7757);
and U8349 (N_8349,N_7809,N_7831);
and U8350 (N_8350,N_7733,N_7939);
and U8351 (N_8351,N_7974,N_7814);
or U8352 (N_8352,N_7855,N_7849);
xor U8353 (N_8353,N_7904,N_7974);
xor U8354 (N_8354,N_7718,N_7751);
nand U8355 (N_8355,N_7742,N_7696);
xor U8356 (N_8356,N_7708,N_7917);
xnor U8357 (N_8357,N_7980,N_7633);
nand U8358 (N_8358,N_7963,N_7605);
or U8359 (N_8359,N_7720,N_7670);
or U8360 (N_8360,N_7747,N_7960);
and U8361 (N_8361,N_7903,N_7832);
or U8362 (N_8362,N_7958,N_7835);
nor U8363 (N_8363,N_7832,N_7766);
and U8364 (N_8364,N_7933,N_7713);
nor U8365 (N_8365,N_7850,N_7648);
xnor U8366 (N_8366,N_7951,N_7985);
xor U8367 (N_8367,N_7653,N_7970);
nand U8368 (N_8368,N_7674,N_7678);
and U8369 (N_8369,N_7949,N_7649);
or U8370 (N_8370,N_7823,N_7868);
nand U8371 (N_8371,N_7628,N_7754);
xor U8372 (N_8372,N_7662,N_7991);
nor U8373 (N_8373,N_7980,N_7833);
xor U8374 (N_8374,N_7608,N_7851);
xnor U8375 (N_8375,N_7803,N_7823);
nor U8376 (N_8376,N_7791,N_7877);
and U8377 (N_8377,N_7621,N_7828);
nor U8378 (N_8378,N_7858,N_7635);
nand U8379 (N_8379,N_7715,N_7651);
xor U8380 (N_8380,N_7866,N_7780);
and U8381 (N_8381,N_7947,N_7883);
or U8382 (N_8382,N_7857,N_7912);
nand U8383 (N_8383,N_7770,N_7650);
nand U8384 (N_8384,N_7680,N_7898);
nor U8385 (N_8385,N_7658,N_7892);
nor U8386 (N_8386,N_7689,N_7825);
xnor U8387 (N_8387,N_7937,N_7995);
or U8388 (N_8388,N_7750,N_7749);
and U8389 (N_8389,N_7624,N_7993);
nor U8390 (N_8390,N_7685,N_7705);
nor U8391 (N_8391,N_7929,N_7826);
nor U8392 (N_8392,N_7895,N_7775);
nand U8393 (N_8393,N_7927,N_7943);
and U8394 (N_8394,N_7775,N_7657);
xnor U8395 (N_8395,N_7692,N_7972);
or U8396 (N_8396,N_7903,N_7862);
nand U8397 (N_8397,N_7767,N_7900);
or U8398 (N_8398,N_7833,N_7848);
nor U8399 (N_8399,N_7667,N_7752);
nor U8400 (N_8400,N_8067,N_8321);
nor U8401 (N_8401,N_8225,N_8149);
and U8402 (N_8402,N_8061,N_8376);
xor U8403 (N_8403,N_8363,N_8381);
or U8404 (N_8404,N_8188,N_8009);
xnor U8405 (N_8405,N_8071,N_8319);
nor U8406 (N_8406,N_8287,N_8174);
and U8407 (N_8407,N_8010,N_8161);
nand U8408 (N_8408,N_8013,N_8093);
xor U8409 (N_8409,N_8041,N_8057);
and U8410 (N_8410,N_8270,N_8063);
or U8411 (N_8411,N_8043,N_8290);
and U8412 (N_8412,N_8104,N_8269);
or U8413 (N_8413,N_8175,N_8348);
and U8414 (N_8414,N_8144,N_8142);
or U8415 (N_8415,N_8011,N_8111);
and U8416 (N_8416,N_8140,N_8261);
or U8417 (N_8417,N_8236,N_8073);
and U8418 (N_8418,N_8017,N_8280);
or U8419 (N_8419,N_8024,N_8090);
or U8420 (N_8420,N_8271,N_8323);
nand U8421 (N_8421,N_8293,N_8092);
nand U8422 (N_8422,N_8326,N_8354);
or U8423 (N_8423,N_8184,N_8247);
or U8424 (N_8424,N_8055,N_8322);
or U8425 (N_8425,N_8251,N_8050);
nand U8426 (N_8426,N_8005,N_8203);
xor U8427 (N_8427,N_8302,N_8023);
and U8428 (N_8428,N_8334,N_8276);
xor U8429 (N_8429,N_8353,N_8197);
xnor U8430 (N_8430,N_8231,N_8177);
nand U8431 (N_8431,N_8008,N_8386);
xor U8432 (N_8432,N_8291,N_8033);
nand U8433 (N_8433,N_8153,N_8282);
nor U8434 (N_8434,N_8172,N_8329);
nand U8435 (N_8435,N_8118,N_8000);
xnor U8436 (N_8436,N_8257,N_8341);
and U8437 (N_8437,N_8245,N_8204);
nor U8438 (N_8438,N_8365,N_8106);
nand U8439 (N_8439,N_8345,N_8044);
nand U8440 (N_8440,N_8312,N_8389);
xnor U8441 (N_8441,N_8186,N_8292);
and U8442 (N_8442,N_8187,N_8195);
nand U8443 (N_8443,N_8058,N_8035);
nand U8444 (N_8444,N_8391,N_8128);
xnor U8445 (N_8445,N_8100,N_8301);
nand U8446 (N_8446,N_8121,N_8125);
and U8447 (N_8447,N_8053,N_8029);
nor U8448 (N_8448,N_8311,N_8099);
xnor U8449 (N_8449,N_8374,N_8238);
nor U8450 (N_8450,N_8155,N_8046);
or U8451 (N_8451,N_8239,N_8180);
nor U8452 (N_8452,N_8392,N_8114);
nand U8453 (N_8453,N_8021,N_8042);
nand U8454 (N_8454,N_8022,N_8262);
nor U8455 (N_8455,N_8372,N_8229);
xor U8456 (N_8456,N_8250,N_8325);
nand U8457 (N_8457,N_8030,N_8356);
nand U8458 (N_8458,N_8308,N_8315);
nor U8459 (N_8459,N_8107,N_8281);
or U8460 (N_8460,N_8095,N_8303);
xnor U8461 (N_8461,N_8160,N_8223);
and U8462 (N_8462,N_8131,N_8216);
xnor U8463 (N_8463,N_8332,N_8387);
or U8464 (N_8464,N_8176,N_8335);
nand U8465 (N_8465,N_8163,N_8336);
nand U8466 (N_8466,N_8215,N_8083);
or U8467 (N_8467,N_8265,N_8220);
or U8468 (N_8468,N_8375,N_8091);
or U8469 (N_8469,N_8169,N_8233);
and U8470 (N_8470,N_8117,N_8285);
nor U8471 (N_8471,N_8306,N_8279);
or U8472 (N_8472,N_8004,N_8337);
nand U8473 (N_8473,N_8112,N_8396);
nor U8474 (N_8474,N_8016,N_8190);
xnor U8475 (N_8475,N_8108,N_8137);
nor U8476 (N_8476,N_8059,N_8113);
or U8477 (N_8477,N_8222,N_8317);
nor U8478 (N_8478,N_8380,N_8212);
nor U8479 (N_8479,N_8088,N_8152);
and U8480 (N_8480,N_8079,N_8066);
nand U8481 (N_8481,N_8116,N_8249);
nor U8482 (N_8482,N_8036,N_8006);
and U8483 (N_8483,N_8272,N_8331);
and U8484 (N_8484,N_8367,N_8087);
nor U8485 (N_8485,N_8089,N_8134);
xor U8486 (N_8486,N_8146,N_8235);
nor U8487 (N_8487,N_8358,N_8051);
and U8488 (N_8488,N_8020,N_8343);
nand U8489 (N_8489,N_8098,N_8018);
or U8490 (N_8490,N_8047,N_8031);
nand U8491 (N_8491,N_8344,N_8397);
nor U8492 (N_8492,N_8234,N_8075);
or U8493 (N_8493,N_8065,N_8274);
nor U8494 (N_8494,N_8286,N_8357);
nand U8495 (N_8495,N_8246,N_8283);
or U8496 (N_8496,N_8192,N_8154);
or U8497 (N_8497,N_8384,N_8119);
nor U8498 (N_8498,N_8122,N_8151);
nor U8499 (N_8499,N_8109,N_8295);
nor U8500 (N_8500,N_8252,N_8148);
nand U8501 (N_8501,N_8191,N_8110);
or U8502 (N_8502,N_8143,N_8012);
xnor U8503 (N_8503,N_8294,N_8064);
xnor U8504 (N_8504,N_8040,N_8309);
xnor U8505 (N_8505,N_8318,N_8078);
xor U8506 (N_8506,N_8390,N_8147);
or U8507 (N_8507,N_8362,N_8349);
nand U8508 (N_8508,N_8277,N_8001);
nand U8509 (N_8509,N_8399,N_8048);
or U8510 (N_8510,N_8364,N_8260);
and U8511 (N_8511,N_8217,N_8305);
and U8512 (N_8512,N_8248,N_8346);
or U8513 (N_8513,N_8178,N_8359);
xor U8514 (N_8514,N_8015,N_8237);
or U8515 (N_8515,N_8141,N_8081);
or U8516 (N_8516,N_8227,N_8200);
or U8517 (N_8517,N_8347,N_8136);
nor U8518 (N_8518,N_8313,N_8157);
and U8519 (N_8519,N_8115,N_8077);
and U8520 (N_8520,N_8056,N_8062);
and U8521 (N_8521,N_8162,N_8342);
and U8522 (N_8522,N_8201,N_8264);
xor U8523 (N_8523,N_8070,N_8219);
or U8524 (N_8524,N_8158,N_8310);
and U8525 (N_8525,N_8126,N_8027);
nor U8526 (N_8526,N_8129,N_8330);
xor U8527 (N_8527,N_8241,N_8164);
and U8528 (N_8528,N_8038,N_8068);
or U8529 (N_8529,N_8382,N_8124);
or U8530 (N_8530,N_8103,N_8284);
and U8531 (N_8531,N_8254,N_8352);
nand U8532 (N_8532,N_8307,N_8300);
or U8533 (N_8533,N_8259,N_8338);
xor U8534 (N_8534,N_8086,N_8393);
nor U8535 (N_8535,N_8255,N_8328);
xnor U8536 (N_8536,N_8173,N_8185);
and U8537 (N_8537,N_8355,N_8373);
or U8538 (N_8538,N_8166,N_8368);
nor U8539 (N_8539,N_8139,N_8214);
and U8540 (N_8540,N_8127,N_8206);
xnor U8541 (N_8541,N_8189,N_8130);
nor U8542 (N_8542,N_8032,N_8224);
nor U8543 (N_8543,N_8179,N_8025);
or U8544 (N_8544,N_8094,N_8327);
xnor U8545 (N_8545,N_8275,N_8298);
nand U8546 (N_8546,N_8105,N_8243);
xor U8547 (N_8547,N_8210,N_8181);
nand U8548 (N_8548,N_8034,N_8072);
xor U8549 (N_8549,N_8314,N_8199);
xor U8550 (N_8550,N_8268,N_8054);
or U8551 (N_8551,N_8003,N_8221);
nor U8552 (N_8552,N_8168,N_8288);
xnor U8553 (N_8553,N_8198,N_8232);
xnor U8554 (N_8554,N_8019,N_8266);
xnor U8555 (N_8555,N_8209,N_8202);
and U8556 (N_8556,N_8135,N_8208);
or U8557 (N_8557,N_8028,N_8371);
or U8558 (N_8558,N_8388,N_8213);
nand U8559 (N_8559,N_8256,N_8273);
nand U8560 (N_8560,N_8069,N_8120);
nor U8561 (N_8561,N_8037,N_8320);
or U8562 (N_8562,N_8205,N_8304);
xnor U8563 (N_8563,N_8049,N_8228);
xnor U8564 (N_8564,N_8039,N_8351);
xnor U8565 (N_8565,N_8211,N_8289);
xor U8566 (N_8566,N_8076,N_8002);
nor U8567 (N_8567,N_8026,N_8183);
xnor U8568 (N_8568,N_8014,N_8132);
xor U8569 (N_8569,N_8194,N_8316);
or U8570 (N_8570,N_8145,N_8096);
or U8571 (N_8571,N_8350,N_8366);
xnor U8572 (N_8572,N_8395,N_8102);
nand U8573 (N_8573,N_8165,N_8226);
nor U8574 (N_8574,N_8060,N_8297);
xnor U8575 (N_8575,N_8253,N_8150);
or U8576 (N_8576,N_8156,N_8193);
nand U8577 (N_8577,N_8080,N_8244);
xnor U8578 (N_8578,N_8171,N_8045);
and U8579 (N_8579,N_8133,N_8394);
xnor U8580 (N_8580,N_8361,N_8085);
nand U8581 (N_8581,N_8267,N_8398);
xnor U8582 (N_8582,N_8123,N_8138);
nor U8583 (N_8583,N_8258,N_8324);
nand U8584 (N_8584,N_8360,N_8370);
or U8585 (N_8585,N_8084,N_8383);
nand U8586 (N_8586,N_8379,N_8097);
xor U8587 (N_8587,N_8182,N_8242);
nand U8588 (N_8588,N_8369,N_8167);
xnor U8589 (N_8589,N_8052,N_8230);
and U8590 (N_8590,N_8207,N_8333);
nor U8591 (N_8591,N_8378,N_8377);
and U8592 (N_8592,N_8101,N_8082);
nand U8593 (N_8593,N_8159,N_8299);
xor U8594 (N_8594,N_8074,N_8339);
and U8595 (N_8595,N_8385,N_8263);
nand U8596 (N_8596,N_8007,N_8340);
xnor U8597 (N_8597,N_8170,N_8196);
or U8598 (N_8598,N_8240,N_8278);
xor U8599 (N_8599,N_8296,N_8218);
xnor U8600 (N_8600,N_8130,N_8243);
or U8601 (N_8601,N_8328,N_8198);
and U8602 (N_8602,N_8392,N_8126);
nor U8603 (N_8603,N_8240,N_8292);
nand U8604 (N_8604,N_8242,N_8065);
or U8605 (N_8605,N_8189,N_8036);
nand U8606 (N_8606,N_8121,N_8259);
or U8607 (N_8607,N_8398,N_8356);
and U8608 (N_8608,N_8105,N_8089);
nor U8609 (N_8609,N_8119,N_8102);
nand U8610 (N_8610,N_8020,N_8388);
nand U8611 (N_8611,N_8131,N_8144);
or U8612 (N_8612,N_8107,N_8398);
or U8613 (N_8613,N_8126,N_8357);
xor U8614 (N_8614,N_8273,N_8149);
nor U8615 (N_8615,N_8346,N_8357);
or U8616 (N_8616,N_8246,N_8126);
nand U8617 (N_8617,N_8125,N_8254);
xnor U8618 (N_8618,N_8164,N_8238);
nand U8619 (N_8619,N_8294,N_8183);
xnor U8620 (N_8620,N_8346,N_8034);
or U8621 (N_8621,N_8102,N_8114);
and U8622 (N_8622,N_8356,N_8246);
or U8623 (N_8623,N_8330,N_8033);
xor U8624 (N_8624,N_8122,N_8002);
and U8625 (N_8625,N_8261,N_8340);
nand U8626 (N_8626,N_8209,N_8005);
xnor U8627 (N_8627,N_8016,N_8039);
nor U8628 (N_8628,N_8059,N_8261);
nor U8629 (N_8629,N_8320,N_8002);
xnor U8630 (N_8630,N_8003,N_8336);
and U8631 (N_8631,N_8254,N_8367);
xor U8632 (N_8632,N_8246,N_8141);
nor U8633 (N_8633,N_8122,N_8294);
xnor U8634 (N_8634,N_8204,N_8241);
nand U8635 (N_8635,N_8076,N_8240);
nor U8636 (N_8636,N_8041,N_8291);
or U8637 (N_8637,N_8321,N_8369);
nand U8638 (N_8638,N_8179,N_8260);
nand U8639 (N_8639,N_8031,N_8035);
xor U8640 (N_8640,N_8314,N_8136);
nand U8641 (N_8641,N_8390,N_8337);
or U8642 (N_8642,N_8087,N_8225);
xor U8643 (N_8643,N_8026,N_8093);
and U8644 (N_8644,N_8107,N_8045);
nor U8645 (N_8645,N_8330,N_8008);
and U8646 (N_8646,N_8001,N_8153);
nand U8647 (N_8647,N_8308,N_8015);
or U8648 (N_8648,N_8088,N_8299);
or U8649 (N_8649,N_8163,N_8355);
xor U8650 (N_8650,N_8376,N_8172);
xnor U8651 (N_8651,N_8200,N_8109);
or U8652 (N_8652,N_8156,N_8206);
nand U8653 (N_8653,N_8355,N_8086);
nand U8654 (N_8654,N_8202,N_8031);
and U8655 (N_8655,N_8244,N_8070);
nand U8656 (N_8656,N_8242,N_8184);
xnor U8657 (N_8657,N_8021,N_8154);
and U8658 (N_8658,N_8050,N_8018);
or U8659 (N_8659,N_8200,N_8385);
or U8660 (N_8660,N_8063,N_8119);
and U8661 (N_8661,N_8309,N_8177);
nand U8662 (N_8662,N_8004,N_8046);
or U8663 (N_8663,N_8095,N_8136);
nor U8664 (N_8664,N_8029,N_8387);
nand U8665 (N_8665,N_8054,N_8345);
nor U8666 (N_8666,N_8218,N_8235);
and U8667 (N_8667,N_8302,N_8278);
xnor U8668 (N_8668,N_8233,N_8383);
xnor U8669 (N_8669,N_8152,N_8008);
or U8670 (N_8670,N_8340,N_8118);
nor U8671 (N_8671,N_8075,N_8289);
and U8672 (N_8672,N_8045,N_8304);
nand U8673 (N_8673,N_8189,N_8239);
or U8674 (N_8674,N_8038,N_8215);
nand U8675 (N_8675,N_8157,N_8335);
nor U8676 (N_8676,N_8387,N_8019);
and U8677 (N_8677,N_8265,N_8062);
and U8678 (N_8678,N_8141,N_8075);
nor U8679 (N_8679,N_8142,N_8213);
nand U8680 (N_8680,N_8278,N_8397);
nor U8681 (N_8681,N_8220,N_8335);
nor U8682 (N_8682,N_8320,N_8142);
and U8683 (N_8683,N_8128,N_8274);
nand U8684 (N_8684,N_8191,N_8100);
or U8685 (N_8685,N_8062,N_8381);
or U8686 (N_8686,N_8227,N_8225);
nand U8687 (N_8687,N_8393,N_8186);
xor U8688 (N_8688,N_8250,N_8148);
nand U8689 (N_8689,N_8061,N_8266);
nor U8690 (N_8690,N_8291,N_8251);
or U8691 (N_8691,N_8230,N_8290);
nor U8692 (N_8692,N_8297,N_8057);
xnor U8693 (N_8693,N_8257,N_8148);
or U8694 (N_8694,N_8304,N_8286);
xnor U8695 (N_8695,N_8184,N_8383);
and U8696 (N_8696,N_8113,N_8279);
or U8697 (N_8697,N_8367,N_8187);
or U8698 (N_8698,N_8071,N_8001);
and U8699 (N_8699,N_8020,N_8306);
or U8700 (N_8700,N_8354,N_8095);
or U8701 (N_8701,N_8355,N_8281);
or U8702 (N_8702,N_8199,N_8041);
nand U8703 (N_8703,N_8064,N_8356);
or U8704 (N_8704,N_8042,N_8160);
nand U8705 (N_8705,N_8344,N_8012);
or U8706 (N_8706,N_8258,N_8204);
or U8707 (N_8707,N_8155,N_8309);
or U8708 (N_8708,N_8033,N_8289);
nand U8709 (N_8709,N_8185,N_8096);
and U8710 (N_8710,N_8292,N_8318);
nand U8711 (N_8711,N_8261,N_8248);
or U8712 (N_8712,N_8353,N_8362);
or U8713 (N_8713,N_8088,N_8034);
nor U8714 (N_8714,N_8115,N_8109);
and U8715 (N_8715,N_8085,N_8388);
and U8716 (N_8716,N_8349,N_8041);
nor U8717 (N_8717,N_8065,N_8032);
xor U8718 (N_8718,N_8280,N_8173);
nand U8719 (N_8719,N_8164,N_8022);
nand U8720 (N_8720,N_8050,N_8358);
xor U8721 (N_8721,N_8350,N_8280);
nor U8722 (N_8722,N_8040,N_8237);
nand U8723 (N_8723,N_8042,N_8207);
nand U8724 (N_8724,N_8122,N_8228);
nand U8725 (N_8725,N_8356,N_8276);
nand U8726 (N_8726,N_8072,N_8143);
and U8727 (N_8727,N_8145,N_8287);
xnor U8728 (N_8728,N_8126,N_8147);
nand U8729 (N_8729,N_8054,N_8075);
and U8730 (N_8730,N_8383,N_8328);
nor U8731 (N_8731,N_8159,N_8084);
or U8732 (N_8732,N_8252,N_8354);
and U8733 (N_8733,N_8331,N_8289);
xnor U8734 (N_8734,N_8355,N_8004);
xnor U8735 (N_8735,N_8254,N_8127);
or U8736 (N_8736,N_8064,N_8082);
xnor U8737 (N_8737,N_8385,N_8151);
nand U8738 (N_8738,N_8277,N_8025);
xnor U8739 (N_8739,N_8280,N_8170);
and U8740 (N_8740,N_8204,N_8067);
nand U8741 (N_8741,N_8313,N_8208);
xnor U8742 (N_8742,N_8175,N_8167);
nand U8743 (N_8743,N_8394,N_8052);
or U8744 (N_8744,N_8397,N_8192);
nand U8745 (N_8745,N_8103,N_8131);
nor U8746 (N_8746,N_8293,N_8333);
xnor U8747 (N_8747,N_8114,N_8246);
nand U8748 (N_8748,N_8241,N_8320);
nand U8749 (N_8749,N_8312,N_8029);
or U8750 (N_8750,N_8399,N_8088);
nand U8751 (N_8751,N_8154,N_8211);
xor U8752 (N_8752,N_8105,N_8391);
nor U8753 (N_8753,N_8260,N_8281);
xor U8754 (N_8754,N_8230,N_8316);
xnor U8755 (N_8755,N_8275,N_8146);
or U8756 (N_8756,N_8369,N_8395);
xnor U8757 (N_8757,N_8017,N_8399);
xnor U8758 (N_8758,N_8192,N_8392);
or U8759 (N_8759,N_8259,N_8064);
xnor U8760 (N_8760,N_8111,N_8066);
xor U8761 (N_8761,N_8064,N_8296);
nor U8762 (N_8762,N_8383,N_8150);
nor U8763 (N_8763,N_8146,N_8032);
nand U8764 (N_8764,N_8139,N_8267);
xnor U8765 (N_8765,N_8259,N_8208);
nor U8766 (N_8766,N_8381,N_8007);
and U8767 (N_8767,N_8230,N_8332);
nand U8768 (N_8768,N_8101,N_8221);
nand U8769 (N_8769,N_8233,N_8314);
nor U8770 (N_8770,N_8398,N_8330);
and U8771 (N_8771,N_8329,N_8021);
xor U8772 (N_8772,N_8378,N_8180);
or U8773 (N_8773,N_8180,N_8131);
nor U8774 (N_8774,N_8142,N_8315);
and U8775 (N_8775,N_8207,N_8347);
and U8776 (N_8776,N_8071,N_8064);
and U8777 (N_8777,N_8178,N_8015);
nand U8778 (N_8778,N_8274,N_8148);
nor U8779 (N_8779,N_8144,N_8355);
nor U8780 (N_8780,N_8196,N_8006);
nand U8781 (N_8781,N_8026,N_8166);
nor U8782 (N_8782,N_8376,N_8385);
xnor U8783 (N_8783,N_8333,N_8098);
and U8784 (N_8784,N_8107,N_8289);
nor U8785 (N_8785,N_8102,N_8223);
nand U8786 (N_8786,N_8313,N_8330);
xnor U8787 (N_8787,N_8015,N_8239);
or U8788 (N_8788,N_8133,N_8228);
and U8789 (N_8789,N_8077,N_8107);
and U8790 (N_8790,N_8111,N_8378);
nor U8791 (N_8791,N_8139,N_8268);
or U8792 (N_8792,N_8148,N_8251);
nor U8793 (N_8793,N_8275,N_8292);
nand U8794 (N_8794,N_8154,N_8151);
and U8795 (N_8795,N_8017,N_8310);
or U8796 (N_8796,N_8395,N_8292);
nor U8797 (N_8797,N_8211,N_8261);
and U8798 (N_8798,N_8071,N_8087);
nor U8799 (N_8799,N_8257,N_8003);
nand U8800 (N_8800,N_8784,N_8545);
nand U8801 (N_8801,N_8793,N_8505);
and U8802 (N_8802,N_8508,N_8564);
and U8803 (N_8803,N_8570,N_8483);
nand U8804 (N_8804,N_8704,N_8752);
xor U8805 (N_8805,N_8642,N_8485);
nand U8806 (N_8806,N_8728,N_8684);
xnor U8807 (N_8807,N_8633,N_8490);
or U8808 (N_8808,N_8546,N_8445);
or U8809 (N_8809,N_8475,N_8763);
xor U8810 (N_8810,N_8566,N_8600);
xor U8811 (N_8811,N_8705,N_8405);
nand U8812 (N_8812,N_8640,N_8427);
nor U8813 (N_8813,N_8783,N_8738);
or U8814 (N_8814,N_8658,N_8430);
and U8815 (N_8815,N_8664,N_8726);
xor U8816 (N_8816,N_8671,N_8487);
and U8817 (N_8817,N_8418,N_8429);
and U8818 (N_8818,N_8711,N_8478);
xnor U8819 (N_8819,N_8779,N_8773);
nor U8820 (N_8820,N_8650,N_8404);
nor U8821 (N_8821,N_8562,N_8513);
and U8822 (N_8822,N_8462,N_8608);
nand U8823 (N_8823,N_8695,N_8788);
or U8824 (N_8824,N_8751,N_8764);
or U8825 (N_8825,N_8749,N_8589);
xor U8826 (N_8826,N_8670,N_8424);
xor U8827 (N_8827,N_8786,N_8727);
and U8828 (N_8828,N_8467,N_8472);
and U8829 (N_8829,N_8481,N_8460);
or U8830 (N_8830,N_8482,N_8737);
nor U8831 (N_8831,N_8681,N_8602);
xor U8832 (N_8832,N_8477,N_8451);
or U8833 (N_8833,N_8782,N_8520);
nand U8834 (N_8834,N_8569,N_8753);
and U8835 (N_8835,N_8645,N_8571);
nor U8836 (N_8836,N_8612,N_8506);
nor U8837 (N_8837,N_8497,N_8624);
and U8838 (N_8838,N_8750,N_8628);
or U8839 (N_8839,N_8593,N_8524);
nand U8840 (N_8840,N_8433,N_8551);
or U8841 (N_8841,N_8626,N_8687);
xnor U8842 (N_8842,N_8614,N_8517);
nor U8843 (N_8843,N_8457,N_8573);
nor U8844 (N_8844,N_8748,N_8643);
and U8845 (N_8845,N_8414,N_8426);
nand U8846 (N_8846,N_8438,N_8597);
nand U8847 (N_8847,N_8617,N_8439);
or U8848 (N_8848,N_8436,N_8759);
or U8849 (N_8849,N_8605,N_8618);
xnor U8850 (N_8850,N_8641,N_8534);
and U8851 (N_8851,N_8676,N_8527);
xnor U8852 (N_8852,N_8668,N_8700);
nor U8853 (N_8853,N_8459,N_8548);
nor U8854 (N_8854,N_8494,N_8544);
and U8855 (N_8855,N_8489,N_8563);
and U8856 (N_8856,N_8715,N_8619);
nand U8857 (N_8857,N_8576,N_8568);
nor U8858 (N_8858,N_8796,N_8507);
and U8859 (N_8859,N_8656,N_8722);
and U8860 (N_8860,N_8549,N_8590);
and U8861 (N_8861,N_8678,N_8630);
or U8862 (N_8862,N_8510,N_8615);
and U8863 (N_8863,N_8691,N_8479);
nor U8864 (N_8864,N_8558,N_8532);
xnor U8865 (N_8865,N_8543,N_8606);
xor U8866 (N_8866,N_8537,N_8428);
or U8867 (N_8867,N_8694,N_8635);
nor U8868 (N_8868,N_8542,N_8533);
nand U8869 (N_8869,N_8657,N_8702);
or U8870 (N_8870,N_8789,N_8639);
or U8871 (N_8871,N_8743,N_8447);
nand U8872 (N_8872,N_8667,N_8683);
xnor U8873 (N_8873,N_8578,N_8651);
or U8874 (N_8874,N_8770,N_8735);
xor U8875 (N_8875,N_8781,N_8415);
and U8876 (N_8876,N_8774,N_8791);
and U8877 (N_8877,N_8446,N_8499);
nor U8878 (N_8878,N_8648,N_8586);
nor U8879 (N_8879,N_8692,N_8461);
nand U8880 (N_8880,N_8583,N_8744);
nor U8881 (N_8881,N_8592,N_8453);
or U8882 (N_8882,N_8588,N_8767);
nor U8883 (N_8883,N_8761,N_8598);
or U8884 (N_8884,N_8634,N_8799);
or U8885 (N_8885,N_8525,N_8638);
and U8886 (N_8886,N_8555,N_8714);
or U8887 (N_8887,N_8603,N_8468);
and U8888 (N_8888,N_8416,N_8740);
nand U8889 (N_8889,N_8442,N_8406);
or U8890 (N_8890,N_8538,N_8529);
or U8891 (N_8891,N_8771,N_8491);
and U8892 (N_8892,N_8777,N_8599);
nand U8893 (N_8893,N_8511,N_8709);
nor U8894 (N_8894,N_8402,N_8629);
and U8895 (N_8895,N_8454,N_8495);
nand U8896 (N_8896,N_8504,N_8584);
nand U8897 (N_8897,N_8607,N_8420);
xnor U8898 (N_8898,N_8673,N_8724);
xnor U8899 (N_8899,N_8775,N_8719);
nor U8900 (N_8900,N_8739,N_8492);
nand U8901 (N_8901,N_8536,N_8655);
or U8902 (N_8902,N_8747,N_8723);
or U8903 (N_8903,N_8622,N_8604);
or U8904 (N_8904,N_8456,N_8732);
or U8905 (N_8905,N_8465,N_8473);
or U8906 (N_8906,N_8672,N_8503);
nor U8907 (N_8907,N_8734,N_8682);
nand U8908 (N_8908,N_8403,N_8745);
or U8909 (N_8909,N_8623,N_8413);
and U8910 (N_8910,N_8528,N_8455);
nor U8911 (N_8911,N_8577,N_8541);
nor U8912 (N_8912,N_8706,N_8725);
nand U8913 (N_8913,N_8526,N_8552);
nand U8914 (N_8914,N_8531,N_8610);
xor U8915 (N_8915,N_8449,N_8409);
xor U8916 (N_8916,N_8649,N_8591);
and U8917 (N_8917,N_8470,N_8557);
or U8918 (N_8918,N_8663,N_8572);
or U8919 (N_8919,N_8729,N_8680);
nand U8920 (N_8920,N_8554,N_8441);
nor U8921 (N_8921,N_8720,N_8654);
or U8922 (N_8922,N_8794,N_8458);
nor U8923 (N_8923,N_8718,N_8757);
and U8924 (N_8924,N_8778,N_8741);
nor U8925 (N_8925,N_8686,N_8580);
nor U8926 (N_8926,N_8419,N_8484);
and U8927 (N_8927,N_8579,N_8636);
and U8928 (N_8928,N_8792,N_8733);
nand U8929 (N_8929,N_8594,N_8707);
or U8930 (N_8930,N_8701,N_8712);
and U8931 (N_8931,N_8766,N_8550);
nand U8932 (N_8932,N_8425,N_8561);
or U8933 (N_8933,N_8708,N_8434);
or U8934 (N_8934,N_8448,N_8790);
or U8935 (N_8935,N_8797,N_8486);
nor U8936 (N_8936,N_8755,N_8408);
and U8937 (N_8937,N_8760,N_8469);
nand U8938 (N_8938,N_8768,N_8518);
and U8939 (N_8939,N_8713,N_8567);
xor U8940 (N_8940,N_8652,N_8547);
or U8941 (N_8941,N_8746,N_8535);
xor U8942 (N_8942,N_8466,N_8412);
xor U8943 (N_8943,N_8587,N_8595);
and U8944 (N_8944,N_8776,N_8498);
nor U8945 (N_8945,N_8496,N_8717);
nand U8946 (N_8946,N_8647,N_8488);
nor U8947 (N_8947,N_8710,N_8696);
and U8948 (N_8948,N_8440,N_8798);
nand U8949 (N_8949,N_8693,N_8515);
xor U8950 (N_8950,N_8674,N_8697);
xor U8951 (N_8951,N_8539,N_8690);
nor U8952 (N_8952,N_8574,N_8450);
and U8953 (N_8953,N_8731,N_8613);
or U8954 (N_8954,N_8616,N_8754);
nor U8955 (N_8955,N_8611,N_8500);
or U8956 (N_8956,N_8677,N_8621);
nor U8957 (N_8957,N_8410,N_8407);
nor U8958 (N_8958,N_8501,N_8769);
or U8959 (N_8959,N_8665,N_8516);
and U8960 (N_8960,N_8540,N_8631);
or U8961 (N_8961,N_8582,N_8756);
nor U8962 (N_8962,N_8530,N_8785);
nand U8963 (N_8963,N_8553,N_8758);
xor U8964 (N_8964,N_8685,N_8575);
xnor U8965 (N_8965,N_8679,N_8772);
nand U8966 (N_8966,N_8581,N_8730);
and U8967 (N_8967,N_8417,N_8646);
nor U8968 (N_8968,N_8666,N_8661);
or U8969 (N_8969,N_8502,N_8795);
and U8970 (N_8970,N_8400,N_8653);
nand U8971 (N_8971,N_8476,N_8689);
nand U8972 (N_8972,N_8556,N_8787);
and U8973 (N_8973,N_8422,N_8444);
nand U8974 (N_8974,N_8716,N_8620);
nand U8975 (N_8975,N_8423,N_8601);
xor U8976 (N_8976,N_8780,N_8662);
nand U8977 (N_8977,N_8762,N_8637);
nand U8978 (N_8978,N_8644,N_8452);
or U8979 (N_8979,N_8464,N_8523);
xnor U8980 (N_8980,N_8659,N_8742);
and U8981 (N_8981,N_8435,N_8698);
nor U8982 (N_8982,N_8565,N_8519);
and U8983 (N_8983,N_8703,N_8401);
nor U8984 (N_8984,N_8432,N_8509);
nor U8985 (N_8985,N_8522,N_8512);
xnor U8986 (N_8986,N_8521,N_8474);
or U8987 (N_8987,N_8632,N_8411);
nand U8988 (N_8988,N_8559,N_8514);
nor U8989 (N_8989,N_8721,N_8480);
or U8990 (N_8990,N_8699,N_8625);
nor U8991 (N_8991,N_8675,N_8437);
or U8992 (N_8992,N_8736,N_8627);
or U8993 (N_8993,N_8471,N_8688);
nor U8994 (N_8994,N_8669,N_8463);
and U8995 (N_8995,N_8660,N_8443);
and U8996 (N_8996,N_8493,N_8560);
nor U8997 (N_8997,N_8596,N_8609);
and U8998 (N_8998,N_8421,N_8585);
or U8999 (N_8999,N_8431,N_8765);
or U9000 (N_9000,N_8492,N_8479);
or U9001 (N_9001,N_8510,N_8515);
and U9002 (N_9002,N_8631,N_8488);
nand U9003 (N_9003,N_8686,N_8556);
and U9004 (N_9004,N_8405,N_8571);
and U9005 (N_9005,N_8611,N_8510);
and U9006 (N_9006,N_8542,N_8635);
or U9007 (N_9007,N_8633,N_8685);
and U9008 (N_9008,N_8459,N_8701);
or U9009 (N_9009,N_8778,N_8668);
nand U9010 (N_9010,N_8517,N_8598);
or U9011 (N_9011,N_8653,N_8495);
nand U9012 (N_9012,N_8656,N_8586);
xor U9013 (N_9013,N_8635,N_8427);
or U9014 (N_9014,N_8587,N_8416);
or U9015 (N_9015,N_8593,N_8484);
or U9016 (N_9016,N_8734,N_8441);
nor U9017 (N_9017,N_8640,N_8406);
nand U9018 (N_9018,N_8772,N_8580);
nor U9019 (N_9019,N_8799,N_8596);
and U9020 (N_9020,N_8549,N_8562);
nor U9021 (N_9021,N_8596,N_8525);
xor U9022 (N_9022,N_8529,N_8462);
or U9023 (N_9023,N_8442,N_8400);
nor U9024 (N_9024,N_8581,N_8639);
nand U9025 (N_9025,N_8690,N_8563);
nor U9026 (N_9026,N_8503,N_8443);
nand U9027 (N_9027,N_8594,N_8752);
or U9028 (N_9028,N_8578,N_8551);
or U9029 (N_9029,N_8664,N_8626);
xor U9030 (N_9030,N_8447,N_8449);
nand U9031 (N_9031,N_8523,N_8652);
and U9032 (N_9032,N_8454,N_8594);
and U9033 (N_9033,N_8713,N_8689);
or U9034 (N_9034,N_8427,N_8532);
nor U9035 (N_9035,N_8530,N_8771);
nand U9036 (N_9036,N_8473,N_8464);
nand U9037 (N_9037,N_8511,N_8680);
and U9038 (N_9038,N_8449,N_8793);
nand U9039 (N_9039,N_8783,N_8768);
nand U9040 (N_9040,N_8662,N_8588);
nand U9041 (N_9041,N_8552,N_8515);
or U9042 (N_9042,N_8416,N_8773);
and U9043 (N_9043,N_8673,N_8646);
nand U9044 (N_9044,N_8514,N_8575);
nand U9045 (N_9045,N_8608,N_8658);
or U9046 (N_9046,N_8630,N_8654);
nand U9047 (N_9047,N_8752,N_8513);
xor U9048 (N_9048,N_8464,N_8658);
or U9049 (N_9049,N_8556,N_8687);
and U9050 (N_9050,N_8434,N_8554);
xnor U9051 (N_9051,N_8411,N_8464);
nor U9052 (N_9052,N_8499,N_8517);
xor U9053 (N_9053,N_8696,N_8749);
nand U9054 (N_9054,N_8480,N_8429);
or U9055 (N_9055,N_8501,N_8763);
nand U9056 (N_9056,N_8769,N_8485);
or U9057 (N_9057,N_8563,N_8700);
nor U9058 (N_9058,N_8686,N_8791);
nand U9059 (N_9059,N_8533,N_8603);
or U9060 (N_9060,N_8757,N_8460);
xor U9061 (N_9061,N_8649,N_8482);
nor U9062 (N_9062,N_8517,N_8762);
xnor U9063 (N_9063,N_8477,N_8547);
nor U9064 (N_9064,N_8568,N_8599);
nand U9065 (N_9065,N_8545,N_8631);
nor U9066 (N_9066,N_8435,N_8723);
nand U9067 (N_9067,N_8790,N_8433);
nor U9068 (N_9068,N_8529,N_8658);
and U9069 (N_9069,N_8414,N_8634);
nand U9070 (N_9070,N_8739,N_8628);
nor U9071 (N_9071,N_8656,N_8457);
nand U9072 (N_9072,N_8622,N_8661);
or U9073 (N_9073,N_8623,N_8456);
xor U9074 (N_9074,N_8611,N_8501);
and U9075 (N_9075,N_8422,N_8509);
or U9076 (N_9076,N_8557,N_8455);
or U9077 (N_9077,N_8517,N_8487);
xor U9078 (N_9078,N_8719,N_8560);
xor U9079 (N_9079,N_8430,N_8779);
or U9080 (N_9080,N_8475,N_8705);
and U9081 (N_9081,N_8583,N_8777);
nand U9082 (N_9082,N_8744,N_8405);
nand U9083 (N_9083,N_8765,N_8495);
and U9084 (N_9084,N_8689,N_8504);
nand U9085 (N_9085,N_8648,N_8798);
xnor U9086 (N_9086,N_8709,N_8646);
nand U9087 (N_9087,N_8441,N_8407);
nor U9088 (N_9088,N_8417,N_8605);
nor U9089 (N_9089,N_8663,N_8712);
or U9090 (N_9090,N_8555,N_8679);
xnor U9091 (N_9091,N_8640,N_8795);
xnor U9092 (N_9092,N_8763,N_8701);
nand U9093 (N_9093,N_8725,N_8491);
nand U9094 (N_9094,N_8748,N_8554);
nor U9095 (N_9095,N_8471,N_8755);
and U9096 (N_9096,N_8715,N_8558);
nand U9097 (N_9097,N_8601,N_8582);
nor U9098 (N_9098,N_8650,N_8660);
or U9099 (N_9099,N_8471,N_8582);
or U9100 (N_9100,N_8540,N_8703);
or U9101 (N_9101,N_8415,N_8647);
nor U9102 (N_9102,N_8736,N_8596);
nand U9103 (N_9103,N_8673,N_8526);
nand U9104 (N_9104,N_8505,N_8568);
and U9105 (N_9105,N_8577,N_8728);
or U9106 (N_9106,N_8532,N_8440);
or U9107 (N_9107,N_8750,N_8660);
nand U9108 (N_9108,N_8406,N_8441);
nor U9109 (N_9109,N_8665,N_8428);
xor U9110 (N_9110,N_8771,N_8549);
and U9111 (N_9111,N_8637,N_8766);
nor U9112 (N_9112,N_8475,N_8568);
and U9113 (N_9113,N_8450,N_8783);
nand U9114 (N_9114,N_8747,N_8608);
nor U9115 (N_9115,N_8595,N_8410);
or U9116 (N_9116,N_8475,N_8700);
or U9117 (N_9117,N_8493,N_8733);
nand U9118 (N_9118,N_8729,N_8434);
nor U9119 (N_9119,N_8743,N_8537);
or U9120 (N_9120,N_8768,N_8628);
nor U9121 (N_9121,N_8796,N_8442);
and U9122 (N_9122,N_8410,N_8699);
and U9123 (N_9123,N_8447,N_8719);
or U9124 (N_9124,N_8494,N_8436);
nor U9125 (N_9125,N_8440,N_8484);
and U9126 (N_9126,N_8623,N_8494);
nor U9127 (N_9127,N_8728,N_8759);
nor U9128 (N_9128,N_8788,N_8457);
or U9129 (N_9129,N_8453,N_8438);
xor U9130 (N_9130,N_8498,N_8771);
and U9131 (N_9131,N_8675,N_8738);
and U9132 (N_9132,N_8681,N_8563);
xor U9133 (N_9133,N_8762,N_8736);
nand U9134 (N_9134,N_8497,N_8499);
nand U9135 (N_9135,N_8701,N_8455);
and U9136 (N_9136,N_8799,N_8493);
and U9137 (N_9137,N_8681,N_8453);
nor U9138 (N_9138,N_8484,N_8687);
nor U9139 (N_9139,N_8702,N_8516);
nor U9140 (N_9140,N_8463,N_8622);
and U9141 (N_9141,N_8492,N_8596);
or U9142 (N_9142,N_8442,N_8485);
nand U9143 (N_9143,N_8782,N_8595);
nand U9144 (N_9144,N_8411,N_8633);
xnor U9145 (N_9145,N_8514,N_8508);
and U9146 (N_9146,N_8513,N_8568);
and U9147 (N_9147,N_8556,N_8683);
xor U9148 (N_9148,N_8608,N_8414);
nand U9149 (N_9149,N_8637,N_8543);
nor U9150 (N_9150,N_8477,N_8499);
xor U9151 (N_9151,N_8766,N_8765);
nor U9152 (N_9152,N_8401,N_8719);
and U9153 (N_9153,N_8481,N_8579);
xnor U9154 (N_9154,N_8673,N_8550);
nor U9155 (N_9155,N_8448,N_8689);
or U9156 (N_9156,N_8452,N_8556);
nor U9157 (N_9157,N_8495,N_8516);
and U9158 (N_9158,N_8426,N_8588);
nand U9159 (N_9159,N_8769,N_8570);
and U9160 (N_9160,N_8700,N_8594);
or U9161 (N_9161,N_8435,N_8566);
or U9162 (N_9162,N_8407,N_8769);
xnor U9163 (N_9163,N_8648,N_8776);
or U9164 (N_9164,N_8761,N_8586);
xor U9165 (N_9165,N_8411,N_8528);
nand U9166 (N_9166,N_8735,N_8797);
nand U9167 (N_9167,N_8400,N_8628);
nor U9168 (N_9168,N_8680,N_8446);
xnor U9169 (N_9169,N_8658,N_8445);
nor U9170 (N_9170,N_8736,N_8639);
xnor U9171 (N_9171,N_8602,N_8726);
and U9172 (N_9172,N_8545,N_8638);
nand U9173 (N_9173,N_8677,N_8524);
or U9174 (N_9174,N_8655,N_8604);
nand U9175 (N_9175,N_8581,N_8791);
nor U9176 (N_9176,N_8433,N_8454);
nand U9177 (N_9177,N_8493,N_8588);
nor U9178 (N_9178,N_8426,N_8471);
nor U9179 (N_9179,N_8664,N_8501);
and U9180 (N_9180,N_8546,N_8527);
xor U9181 (N_9181,N_8536,N_8525);
nor U9182 (N_9182,N_8603,N_8705);
xnor U9183 (N_9183,N_8442,N_8454);
nor U9184 (N_9184,N_8558,N_8466);
nor U9185 (N_9185,N_8472,N_8590);
xnor U9186 (N_9186,N_8774,N_8581);
xor U9187 (N_9187,N_8625,N_8601);
nand U9188 (N_9188,N_8588,N_8419);
nand U9189 (N_9189,N_8420,N_8586);
or U9190 (N_9190,N_8466,N_8779);
or U9191 (N_9191,N_8521,N_8577);
or U9192 (N_9192,N_8623,N_8694);
and U9193 (N_9193,N_8690,N_8501);
nand U9194 (N_9194,N_8603,N_8546);
nand U9195 (N_9195,N_8553,N_8757);
nand U9196 (N_9196,N_8453,N_8477);
and U9197 (N_9197,N_8426,N_8571);
nand U9198 (N_9198,N_8459,N_8741);
nor U9199 (N_9199,N_8441,N_8540);
or U9200 (N_9200,N_9177,N_9150);
nand U9201 (N_9201,N_9033,N_9062);
or U9202 (N_9202,N_9197,N_8880);
and U9203 (N_9203,N_9103,N_8839);
xor U9204 (N_9204,N_9098,N_9143);
xor U9205 (N_9205,N_9072,N_9097);
nand U9206 (N_9206,N_9076,N_9090);
nand U9207 (N_9207,N_9000,N_9096);
nor U9208 (N_9208,N_9095,N_8887);
or U9209 (N_9209,N_8970,N_8933);
nor U9210 (N_9210,N_9131,N_9193);
xnor U9211 (N_9211,N_8892,N_8945);
or U9212 (N_9212,N_8873,N_9044);
nor U9213 (N_9213,N_8999,N_8949);
or U9214 (N_9214,N_9048,N_8846);
nor U9215 (N_9215,N_9114,N_8937);
and U9216 (N_9216,N_8849,N_8996);
and U9217 (N_9217,N_9156,N_8883);
or U9218 (N_9218,N_8906,N_8944);
nand U9219 (N_9219,N_9065,N_8909);
nand U9220 (N_9220,N_8868,N_8802);
xor U9221 (N_9221,N_8997,N_8967);
nand U9222 (N_9222,N_8983,N_8953);
and U9223 (N_9223,N_9021,N_9127);
xnor U9224 (N_9224,N_8852,N_9013);
nor U9225 (N_9225,N_8926,N_9027);
and U9226 (N_9226,N_8801,N_8828);
xor U9227 (N_9227,N_8990,N_9088);
xor U9228 (N_9228,N_8918,N_8901);
xnor U9229 (N_9229,N_8946,N_9029);
or U9230 (N_9230,N_8982,N_9020);
or U9231 (N_9231,N_9007,N_9118);
xnor U9232 (N_9232,N_9025,N_9023);
or U9233 (N_9233,N_9064,N_9190);
xnor U9234 (N_9234,N_9077,N_9172);
nand U9235 (N_9235,N_8914,N_9037);
nand U9236 (N_9236,N_9099,N_9028);
nand U9237 (N_9237,N_9043,N_9012);
nand U9238 (N_9238,N_9063,N_9122);
and U9239 (N_9239,N_8837,N_8896);
nor U9240 (N_9240,N_9060,N_9085);
nor U9241 (N_9241,N_9059,N_8863);
xnor U9242 (N_9242,N_9163,N_9100);
xnor U9243 (N_9243,N_9074,N_9191);
nand U9244 (N_9244,N_8934,N_9093);
nor U9245 (N_9245,N_8987,N_8959);
xor U9246 (N_9246,N_8838,N_9052);
xnor U9247 (N_9247,N_8939,N_9015);
or U9248 (N_9248,N_8958,N_8800);
nor U9249 (N_9249,N_9148,N_9089);
or U9250 (N_9250,N_8927,N_8935);
xnor U9251 (N_9251,N_9011,N_9022);
nor U9252 (N_9252,N_8919,N_8973);
nor U9253 (N_9253,N_9109,N_8834);
xnor U9254 (N_9254,N_8832,N_9178);
and U9255 (N_9255,N_9115,N_8859);
xnor U9256 (N_9256,N_9070,N_9182);
nand U9257 (N_9257,N_9174,N_8836);
nand U9258 (N_9258,N_8893,N_8889);
and U9259 (N_9259,N_8948,N_8879);
nand U9260 (N_9260,N_8855,N_8972);
nand U9261 (N_9261,N_8910,N_9054);
xor U9262 (N_9262,N_9030,N_9144);
nand U9263 (N_9263,N_8871,N_8822);
nor U9264 (N_9264,N_9016,N_8843);
and U9265 (N_9265,N_9073,N_8963);
and U9266 (N_9266,N_9196,N_9050);
xor U9267 (N_9267,N_8804,N_9009);
xor U9268 (N_9268,N_9106,N_8856);
and U9269 (N_9269,N_9075,N_8833);
nor U9270 (N_9270,N_8830,N_9175);
or U9271 (N_9271,N_9056,N_8888);
nor U9272 (N_9272,N_9111,N_9080);
nor U9273 (N_9273,N_9117,N_8897);
nand U9274 (N_9274,N_9035,N_8936);
or U9275 (N_9275,N_8842,N_9102);
and U9276 (N_9276,N_8810,N_9181);
or U9277 (N_9277,N_9199,N_8930);
nand U9278 (N_9278,N_9173,N_9040);
nor U9279 (N_9279,N_9116,N_9008);
xor U9280 (N_9280,N_8803,N_9188);
and U9281 (N_9281,N_8924,N_8984);
xnor U9282 (N_9282,N_9042,N_9142);
or U9283 (N_9283,N_9051,N_8976);
and U9284 (N_9284,N_9176,N_9105);
and U9285 (N_9285,N_8890,N_9170);
or U9286 (N_9286,N_9120,N_8813);
or U9287 (N_9287,N_8965,N_9066);
or U9288 (N_9288,N_9146,N_8957);
nor U9289 (N_9289,N_8925,N_9198);
and U9290 (N_9290,N_9183,N_8917);
xnor U9291 (N_9291,N_8942,N_9165);
nand U9292 (N_9292,N_9087,N_8805);
nand U9293 (N_9293,N_8826,N_8898);
or U9294 (N_9294,N_9112,N_8807);
and U9295 (N_9295,N_9002,N_8903);
nand U9296 (N_9296,N_9123,N_9081);
and U9297 (N_9297,N_8818,N_9057);
nor U9298 (N_9298,N_8913,N_8835);
nor U9299 (N_9299,N_9083,N_8850);
nor U9300 (N_9300,N_9166,N_8819);
or U9301 (N_9301,N_9157,N_8829);
xnor U9302 (N_9302,N_9094,N_8941);
xor U9303 (N_9303,N_8827,N_8840);
or U9304 (N_9304,N_8831,N_9079);
nand U9305 (N_9305,N_8845,N_8865);
or U9306 (N_9306,N_8824,N_9107);
nand U9307 (N_9307,N_8841,N_9152);
nand U9308 (N_9308,N_9069,N_8900);
nor U9309 (N_9309,N_9145,N_9137);
nand U9310 (N_9310,N_8811,N_8820);
or U9311 (N_9311,N_9140,N_9017);
nand U9312 (N_9312,N_9187,N_8932);
and U9313 (N_9313,N_8916,N_8886);
xnor U9314 (N_9314,N_8920,N_8931);
nor U9315 (N_9315,N_8995,N_9110);
nand U9316 (N_9316,N_9168,N_9132);
or U9317 (N_9317,N_9001,N_9014);
nand U9318 (N_9318,N_8978,N_8955);
and U9319 (N_9319,N_9134,N_8816);
and U9320 (N_9320,N_9135,N_8851);
xor U9321 (N_9321,N_9159,N_9186);
and U9322 (N_9322,N_8991,N_9055);
xor U9323 (N_9323,N_9113,N_9041);
xor U9324 (N_9324,N_8848,N_9129);
and U9325 (N_9325,N_8823,N_9092);
nor U9326 (N_9326,N_8861,N_8940);
xnor U9327 (N_9327,N_8992,N_8882);
or U9328 (N_9328,N_9068,N_9101);
and U9329 (N_9329,N_9034,N_9124);
nor U9330 (N_9330,N_9046,N_9091);
and U9331 (N_9331,N_8809,N_9179);
nand U9332 (N_9332,N_8956,N_8902);
xor U9333 (N_9333,N_9160,N_8974);
xor U9334 (N_9334,N_9045,N_8962);
and U9335 (N_9335,N_8971,N_9005);
xnor U9336 (N_9336,N_9194,N_8952);
nor U9337 (N_9337,N_8938,N_9180);
xor U9338 (N_9338,N_8885,N_9167);
nand U9339 (N_9339,N_8894,N_9171);
nor U9340 (N_9340,N_8969,N_9154);
and U9341 (N_9341,N_8814,N_8876);
or U9342 (N_9342,N_9031,N_8985);
nand U9343 (N_9343,N_9026,N_9153);
nand U9344 (N_9344,N_8872,N_8928);
and U9345 (N_9345,N_9047,N_9082);
or U9346 (N_9346,N_8881,N_8923);
or U9347 (N_9347,N_9084,N_8993);
nor U9348 (N_9348,N_9130,N_9058);
nand U9349 (N_9349,N_9024,N_8961);
or U9350 (N_9350,N_9006,N_8922);
nor U9351 (N_9351,N_9139,N_8904);
nor U9352 (N_9352,N_8968,N_9038);
xor U9353 (N_9353,N_8825,N_8943);
or U9354 (N_9354,N_9036,N_9067);
or U9355 (N_9355,N_9125,N_9162);
xnor U9356 (N_9356,N_8899,N_8874);
or U9357 (N_9357,N_9189,N_8988);
nor U9358 (N_9358,N_8921,N_8821);
and U9359 (N_9359,N_9003,N_8884);
nor U9360 (N_9360,N_9121,N_8905);
xnor U9361 (N_9361,N_9104,N_9108);
and U9362 (N_9362,N_9149,N_9078);
and U9363 (N_9363,N_8989,N_8812);
xor U9364 (N_9364,N_9184,N_8954);
xor U9365 (N_9365,N_9147,N_9010);
xor U9366 (N_9366,N_8853,N_9086);
and U9367 (N_9367,N_9141,N_9195);
xor U9368 (N_9368,N_9161,N_8977);
or U9369 (N_9369,N_8911,N_9119);
nand U9370 (N_9370,N_8869,N_8907);
or U9371 (N_9371,N_8980,N_8947);
and U9372 (N_9372,N_8857,N_8870);
nand U9373 (N_9373,N_8815,N_9049);
xnor U9374 (N_9374,N_8994,N_8979);
or U9375 (N_9375,N_9053,N_8986);
or U9376 (N_9376,N_9155,N_8806);
nor U9377 (N_9377,N_8866,N_8877);
xor U9378 (N_9378,N_8864,N_9061);
and U9379 (N_9379,N_8867,N_8878);
xnor U9380 (N_9380,N_9039,N_9018);
or U9381 (N_9381,N_8915,N_9032);
or U9382 (N_9382,N_8981,N_8891);
or U9383 (N_9383,N_9071,N_8858);
nor U9384 (N_9384,N_8808,N_9004);
or U9385 (N_9385,N_9136,N_8862);
nor U9386 (N_9386,N_8847,N_8960);
xor U9387 (N_9387,N_8860,N_9151);
xor U9388 (N_9388,N_8908,N_9169);
and U9389 (N_9389,N_8844,N_9185);
xnor U9390 (N_9390,N_8875,N_8975);
nor U9391 (N_9391,N_9164,N_9192);
nor U9392 (N_9392,N_8817,N_8951);
and U9393 (N_9393,N_8929,N_9019);
nand U9394 (N_9394,N_8895,N_9158);
nand U9395 (N_9395,N_8950,N_8998);
or U9396 (N_9396,N_8966,N_8854);
and U9397 (N_9397,N_9138,N_8964);
or U9398 (N_9398,N_8912,N_9128);
nand U9399 (N_9399,N_9126,N_9133);
or U9400 (N_9400,N_8995,N_9132);
nor U9401 (N_9401,N_8908,N_8939);
nor U9402 (N_9402,N_8822,N_9161);
and U9403 (N_9403,N_9012,N_9055);
xnor U9404 (N_9404,N_9072,N_9030);
nor U9405 (N_9405,N_9093,N_9054);
nand U9406 (N_9406,N_9121,N_9124);
nand U9407 (N_9407,N_9134,N_8959);
nand U9408 (N_9408,N_9025,N_9154);
nand U9409 (N_9409,N_8925,N_9079);
xnor U9410 (N_9410,N_9135,N_8902);
and U9411 (N_9411,N_9148,N_9011);
or U9412 (N_9412,N_8957,N_8951);
nor U9413 (N_9413,N_8942,N_8837);
or U9414 (N_9414,N_9013,N_9090);
nor U9415 (N_9415,N_9148,N_8845);
or U9416 (N_9416,N_9077,N_8948);
xor U9417 (N_9417,N_9047,N_9136);
xor U9418 (N_9418,N_9075,N_8952);
nand U9419 (N_9419,N_9123,N_9019);
nand U9420 (N_9420,N_8889,N_9072);
xor U9421 (N_9421,N_9114,N_8980);
and U9422 (N_9422,N_8943,N_9016);
xor U9423 (N_9423,N_8911,N_8832);
and U9424 (N_9424,N_9121,N_9183);
or U9425 (N_9425,N_8962,N_9074);
or U9426 (N_9426,N_8903,N_8998);
nor U9427 (N_9427,N_8839,N_9105);
and U9428 (N_9428,N_9139,N_9170);
and U9429 (N_9429,N_8896,N_8853);
nor U9430 (N_9430,N_9005,N_9167);
or U9431 (N_9431,N_8846,N_8845);
or U9432 (N_9432,N_8818,N_8977);
nor U9433 (N_9433,N_9055,N_9007);
nor U9434 (N_9434,N_9092,N_8928);
or U9435 (N_9435,N_9019,N_8958);
or U9436 (N_9436,N_8937,N_8873);
nor U9437 (N_9437,N_8970,N_8901);
or U9438 (N_9438,N_8918,N_8988);
and U9439 (N_9439,N_9033,N_9100);
nor U9440 (N_9440,N_8894,N_9119);
or U9441 (N_9441,N_9042,N_9091);
and U9442 (N_9442,N_9182,N_9184);
xor U9443 (N_9443,N_8900,N_8880);
or U9444 (N_9444,N_9158,N_9075);
or U9445 (N_9445,N_9033,N_9093);
nand U9446 (N_9446,N_9062,N_8880);
xnor U9447 (N_9447,N_9171,N_9072);
and U9448 (N_9448,N_9163,N_8806);
or U9449 (N_9449,N_8888,N_8925);
or U9450 (N_9450,N_8844,N_8963);
nor U9451 (N_9451,N_8887,N_9154);
nand U9452 (N_9452,N_9080,N_8809);
nor U9453 (N_9453,N_8938,N_9194);
and U9454 (N_9454,N_8887,N_8922);
or U9455 (N_9455,N_8811,N_8821);
nand U9456 (N_9456,N_8948,N_8908);
xor U9457 (N_9457,N_8932,N_9093);
and U9458 (N_9458,N_9110,N_8842);
and U9459 (N_9459,N_9044,N_9013);
xor U9460 (N_9460,N_8972,N_8954);
nand U9461 (N_9461,N_8945,N_8801);
and U9462 (N_9462,N_9178,N_9147);
nand U9463 (N_9463,N_8986,N_9126);
nor U9464 (N_9464,N_8860,N_8898);
nand U9465 (N_9465,N_8862,N_9140);
nor U9466 (N_9466,N_9151,N_8845);
or U9467 (N_9467,N_9117,N_8895);
nor U9468 (N_9468,N_9135,N_8974);
and U9469 (N_9469,N_8844,N_9116);
nor U9470 (N_9470,N_9069,N_8995);
xnor U9471 (N_9471,N_8995,N_8880);
nand U9472 (N_9472,N_8904,N_9104);
nor U9473 (N_9473,N_8890,N_9140);
and U9474 (N_9474,N_9044,N_8915);
nand U9475 (N_9475,N_9094,N_8919);
xnor U9476 (N_9476,N_8882,N_8888);
and U9477 (N_9477,N_8802,N_8841);
xor U9478 (N_9478,N_9007,N_9020);
nand U9479 (N_9479,N_9192,N_8809);
nand U9480 (N_9480,N_9115,N_9148);
nor U9481 (N_9481,N_9140,N_9168);
and U9482 (N_9482,N_9070,N_8884);
xnor U9483 (N_9483,N_9109,N_9172);
xnor U9484 (N_9484,N_9021,N_8966);
or U9485 (N_9485,N_9137,N_8920);
or U9486 (N_9486,N_8831,N_8922);
and U9487 (N_9487,N_8915,N_9074);
nand U9488 (N_9488,N_9052,N_9025);
nor U9489 (N_9489,N_8852,N_9046);
or U9490 (N_9490,N_9188,N_9130);
or U9491 (N_9491,N_8957,N_8983);
xnor U9492 (N_9492,N_9181,N_9055);
xor U9493 (N_9493,N_8975,N_8928);
nor U9494 (N_9494,N_9022,N_9046);
and U9495 (N_9495,N_9112,N_9184);
nand U9496 (N_9496,N_9091,N_9116);
nand U9497 (N_9497,N_9145,N_9031);
and U9498 (N_9498,N_8898,N_8964);
xnor U9499 (N_9499,N_9096,N_8921);
nand U9500 (N_9500,N_8832,N_8955);
and U9501 (N_9501,N_9067,N_9161);
nand U9502 (N_9502,N_8970,N_8957);
or U9503 (N_9503,N_8843,N_8998);
nor U9504 (N_9504,N_8914,N_9112);
xnor U9505 (N_9505,N_9091,N_8901);
or U9506 (N_9506,N_8938,N_8962);
or U9507 (N_9507,N_9179,N_8821);
nor U9508 (N_9508,N_8937,N_8879);
nor U9509 (N_9509,N_9033,N_9087);
or U9510 (N_9510,N_8949,N_8811);
and U9511 (N_9511,N_9098,N_8994);
nand U9512 (N_9512,N_9009,N_8847);
nand U9513 (N_9513,N_8850,N_8954);
or U9514 (N_9514,N_9015,N_9135);
nand U9515 (N_9515,N_9038,N_9116);
xnor U9516 (N_9516,N_9055,N_8825);
xnor U9517 (N_9517,N_9000,N_8876);
or U9518 (N_9518,N_8925,N_8979);
or U9519 (N_9519,N_8912,N_9114);
and U9520 (N_9520,N_9156,N_9033);
xor U9521 (N_9521,N_8811,N_8946);
xor U9522 (N_9522,N_9119,N_8970);
and U9523 (N_9523,N_8894,N_9086);
nor U9524 (N_9524,N_8869,N_9058);
and U9525 (N_9525,N_8839,N_9122);
xor U9526 (N_9526,N_8964,N_9150);
nand U9527 (N_9527,N_9091,N_8937);
and U9528 (N_9528,N_8864,N_8836);
xnor U9529 (N_9529,N_8860,N_9074);
or U9530 (N_9530,N_9114,N_8838);
or U9531 (N_9531,N_9186,N_9060);
nor U9532 (N_9532,N_9083,N_8933);
xnor U9533 (N_9533,N_8847,N_8976);
xor U9534 (N_9534,N_9051,N_8887);
or U9535 (N_9535,N_8909,N_9119);
and U9536 (N_9536,N_8965,N_8814);
or U9537 (N_9537,N_9069,N_8933);
nor U9538 (N_9538,N_9072,N_8861);
xor U9539 (N_9539,N_9128,N_9183);
xor U9540 (N_9540,N_8997,N_9094);
or U9541 (N_9541,N_8942,N_8883);
and U9542 (N_9542,N_9145,N_9013);
nor U9543 (N_9543,N_9017,N_8848);
and U9544 (N_9544,N_9073,N_9015);
xnor U9545 (N_9545,N_9127,N_8884);
or U9546 (N_9546,N_8974,N_8915);
nand U9547 (N_9547,N_8843,N_8951);
nand U9548 (N_9548,N_9099,N_8917);
and U9549 (N_9549,N_8906,N_9169);
or U9550 (N_9550,N_8978,N_9193);
and U9551 (N_9551,N_9133,N_9000);
nor U9552 (N_9552,N_9070,N_9165);
nor U9553 (N_9553,N_8830,N_8841);
nor U9554 (N_9554,N_8946,N_8846);
xor U9555 (N_9555,N_9194,N_9031);
and U9556 (N_9556,N_8923,N_9108);
nand U9557 (N_9557,N_9018,N_8948);
nor U9558 (N_9558,N_9137,N_9073);
xnor U9559 (N_9559,N_9004,N_9141);
xnor U9560 (N_9560,N_9020,N_9112);
nand U9561 (N_9561,N_8948,N_9127);
xnor U9562 (N_9562,N_9139,N_9105);
nand U9563 (N_9563,N_8987,N_9195);
xor U9564 (N_9564,N_9041,N_9076);
xor U9565 (N_9565,N_9055,N_8980);
nor U9566 (N_9566,N_9070,N_9113);
nor U9567 (N_9567,N_9011,N_9166);
nor U9568 (N_9568,N_8925,N_8902);
or U9569 (N_9569,N_8960,N_9009);
xnor U9570 (N_9570,N_8801,N_8842);
or U9571 (N_9571,N_9189,N_9056);
nand U9572 (N_9572,N_8897,N_8965);
or U9573 (N_9573,N_8825,N_8865);
nand U9574 (N_9574,N_8861,N_9094);
and U9575 (N_9575,N_9061,N_8832);
or U9576 (N_9576,N_8867,N_8951);
and U9577 (N_9577,N_8822,N_9175);
and U9578 (N_9578,N_9031,N_8948);
nand U9579 (N_9579,N_8913,N_9057);
xor U9580 (N_9580,N_9136,N_9135);
or U9581 (N_9581,N_9182,N_9136);
xor U9582 (N_9582,N_8923,N_9069);
or U9583 (N_9583,N_9099,N_9092);
nor U9584 (N_9584,N_8919,N_8924);
or U9585 (N_9585,N_9061,N_9122);
nand U9586 (N_9586,N_9091,N_8932);
nor U9587 (N_9587,N_9074,N_9024);
nand U9588 (N_9588,N_8841,N_8816);
xnor U9589 (N_9589,N_8863,N_9124);
nand U9590 (N_9590,N_9065,N_8811);
and U9591 (N_9591,N_9021,N_9091);
nor U9592 (N_9592,N_8849,N_8932);
nor U9593 (N_9593,N_8868,N_8881);
or U9594 (N_9594,N_8882,N_8844);
or U9595 (N_9595,N_8892,N_9126);
xor U9596 (N_9596,N_8967,N_9029);
xor U9597 (N_9597,N_9177,N_9167);
and U9598 (N_9598,N_8846,N_9084);
nor U9599 (N_9599,N_8991,N_9112);
nor U9600 (N_9600,N_9327,N_9389);
nand U9601 (N_9601,N_9200,N_9438);
or U9602 (N_9602,N_9233,N_9317);
or U9603 (N_9603,N_9297,N_9406);
nor U9604 (N_9604,N_9331,N_9275);
nor U9605 (N_9605,N_9516,N_9299);
nor U9606 (N_9606,N_9420,N_9397);
nor U9607 (N_9607,N_9258,N_9321);
xnor U9608 (N_9608,N_9418,N_9525);
nand U9609 (N_9609,N_9293,N_9505);
nor U9610 (N_9610,N_9421,N_9497);
or U9611 (N_9611,N_9555,N_9213);
nand U9612 (N_9612,N_9435,N_9534);
nand U9613 (N_9613,N_9387,N_9352);
nand U9614 (N_9614,N_9262,N_9247);
xnor U9615 (N_9615,N_9443,N_9318);
nor U9616 (N_9616,N_9308,N_9373);
nor U9617 (N_9617,N_9260,N_9557);
xnor U9618 (N_9618,N_9395,N_9562);
xor U9619 (N_9619,N_9205,N_9245);
nor U9620 (N_9620,N_9261,N_9411);
xor U9621 (N_9621,N_9429,N_9502);
nor U9622 (N_9622,N_9504,N_9246);
nor U9623 (N_9623,N_9463,N_9253);
xnor U9624 (N_9624,N_9495,N_9540);
xnor U9625 (N_9625,N_9343,N_9573);
and U9626 (N_9626,N_9524,N_9460);
nand U9627 (N_9627,N_9536,N_9442);
nor U9628 (N_9628,N_9339,N_9263);
xor U9629 (N_9629,N_9423,N_9314);
or U9630 (N_9630,N_9288,N_9486);
nand U9631 (N_9631,N_9431,N_9590);
and U9632 (N_9632,N_9474,N_9307);
xnor U9633 (N_9633,N_9273,N_9394);
nor U9634 (N_9634,N_9466,N_9264);
nand U9635 (N_9635,N_9207,N_9357);
nand U9636 (N_9636,N_9224,N_9329);
nor U9637 (N_9637,N_9455,N_9342);
nor U9638 (N_9638,N_9333,N_9465);
xnor U9639 (N_9639,N_9527,N_9271);
nand U9640 (N_9640,N_9336,N_9252);
or U9641 (N_9641,N_9391,N_9596);
or U9642 (N_9642,N_9518,N_9226);
xor U9643 (N_9643,N_9499,N_9599);
or U9644 (N_9644,N_9239,N_9454);
or U9645 (N_9645,N_9383,N_9316);
and U9646 (N_9646,N_9520,N_9552);
or U9647 (N_9647,N_9202,N_9217);
nor U9648 (N_9648,N_9407,N_9348);
and U9649 (N_9649,N_9284,N_9367);
nand U9650 (N_9650,N_9218,N_9522);
and U9651 (N_9651,N_9294,N_9481);
xor U9652 (N_9652,N_9501,N_9434);
nor U9653 (N_9653,N_9227,N_9400);
xor U9654 (N_9654,N_9507,N_9556);
nand U9655 (N_9655,N_9409,N_9313);
or U9656 (N_9656,N_9249,N_9380);
nor U9657 (N_9657,N_9496,N_9519);
nor U9658 (N_9658,N_9512,N_9240);
nand U9659 (N_9659,N_9542,N_9430);
nand U9660 (N_9660,N_9379,N_9475);
and U9661 (N_9661,N_9493,N_9593);
nand U9662 (N_9662,N_9489,N_9576);
nor U9663 (N_9663,N_9347,N_9267);
and U9664 (N_9664,N_9396,N_9377);
xnor U9665 (N_9665,N_9410,N_9513);
nor U9666 (N_9666,N_9248,N_9359);
xnor U9667 (N_9667,N_9285,N_9509);
and U9668 (N_9668,N_9500,N_9353);
or U9669 (N_9669,N_9565,N_9281);
or U9670 (N_9670,N_9483,N_9488);
nor U9671 (N_9671,N_9553,N_9456);
or U9672 (N_9672,N_9584,N_9444);
xnor U9673 (N_9673,N_9328,N_9365);
xnor U9674 (N_9674,N_9278,N_9424);
xnor U9675 (N_9675,N_9287,N_9309);
xnor U9676 (N_9676,N_9378,N_9458);
nor U9677 (N_9677,N_9485,N_9219);
xnor U9678 (N_9678,N_9335,N_9417);
nand U9679 (N_9679,N_9363,N_9371);
nand U9680 (N_9680,N_9511,N_9404);
and U9681 (N_9681,N_9586,N_9223);
nand U9682 (N_9682,N_9432,N_9243);
xor U9683 (N_9683,N_9256,N_9238);
and U9684 (N_9684,N_9571,N_9598);
xnor U9685 (N_9685,N_9514,N_9543);
xor U9686 (N_9686,N_9490,N_9368);
and U9687 (N_9687,N_9208,N_9366);
xor U9688 (N_9688,N_9515,N_9215);
or U9689 (N_9689,N_9484,N_9228);
xor U9690 (N_9690,N_9459,N_9526);
or U9691 (N_9691,N_9324,N_9374);
xor U9692 (N_9692,N_9203,N_9286);
nor U9693 (N_9693,N_9230,N_9265);
and U9694 (N_9694,N_9473,N_9289);
xor U9695 (N_9695,N_9523,N_9535);
nor U9696 (N_9696,N_9222,N_9541);
nor U9697 (N_9697,N_9320,N_9221);
and U9698 (N_9698,N_9510,N_9436);
xnor U9699 (N_9699,N_9419,N_9425);
and U9700 (N_9700,N_9388,N_9594);
xor U9701 (N_9701,N_9449,N_9390);
and U9702 (N_9702,N_9346,N_9538);
nor U9703 (N_9703,N_9296,N_9482);
and U9704 (N_9704,N_9386,N_9440);
nand U9705 (N_9705,N_9457,N_9376);
nor U9706 (N_9706,N_9530,N_9533);
nor U9707 (N_9707,N_9426,N_9547);
and U9708 (N_9708,N_9298,N_9494);
xnor U9709 (N_9709,N_9393,N_9305);
xnor U9710 (N_9710,N_9259,N_9544);
and U9711 (N_9711,N_9401,N_9597);
and U9712 (N_9712,N_9295,N_9487);
xnor U9713 (N_9713,N_9274,N_9550);
and U9714 (N_9714,N_9572,N_9212);
and U9715 (N_9715,N_9453,N_9560);
or U9716 (N_9716,N_9577,N_9399);
nor U9717 (N_9717,N_9311,N_9301);
nand U9718 (N_9718,N_9372,N_9369);
nor U9719 (N_9719,N_9559,N_9338);
nor U9720 (N_9720,N_9300,N_9537);
nor U9721 (N_9721,N_9508,N_9323);
nor U9722 (N_9722,N_9350,N_9469);
and U9723 (N_9723,N_9567,N_9528);
and U9724 (N_9724,N_9546,N_9472);
nand U9725 (N_9725,N_9351,N_9209);
nor U9726 (N_9726,N_9279,N_9362);
or U9727 (N_9727,N_9204,N_9461);
nor U9728 (N_9728,N_9276,N_9232);
and U9729 (N_9729,N_9201,N_9551);
xnor U9730 (N_9730,N_9579,N_9478);
nand U9731 (N_9731,N_9250,N_9451);
and U9732 (N_9732,N_9445,N_9452);
nor U9733 (N_9733,N_9415,N_9414);
or U9734 (N_9734,N_9548,N_9334);
and U9735 (N_9735,N_9422,N_9545);
and U9736 (N_9736,N_9364,N_9392);
and U9737 (N_9737,N_9467,N_9290);
and U9738 (N_9738,N_9582,N_9437);
nor U9739 (N_9739,N_9585,N_9566);
nor U9740 (N_9740,N_9234,N_9277);
nor U9741 (N_9741,N_9303,N_9464);
nand U9742 (N_9742,N_9428,N_9358);
nand U9743 (N_9743,N_9570,N_9257);
or U9744 (N_9744,N_9448,N_9231);
or U9745 (N_9745,N_9283,N_9402);
and U9746 (N_9746,N_9381,N_9255);
and U9747 (N_9747,N_9587,N_9242);
nand U9748 (N_9748,N_9398,N_9237);
or U9749 (N_9749,N_9589,N_9244);
or U9750 (N_9750,N_9446,N_9355);
nor U9751 (N_9751,N_9549,N_9354);
nor U9752 (N_9752,N_9591,N_9531);
or U9753 (N_9753,N_9498,N_9345);
and U9754 (N_9754,N_9340,N_9225);
nand U9755 (N_9755,N_9349,N_9561);
xor U9756 (N_9756,N_9292,N_9385);
nor U9757 (N_9757,N_9408,N_9574);
or U9758 (N_9758,N_9506,N_9581);
and U9759 (N_9759,N_9583,N_9580);
nor U9760 (N_9760,N_9370,N_9360);
and U9761 (N_9761,N_9206,N_9439);
nand U9762 (N_9762,N_9412,N_9241);
and U9763 (N_9763,N_9269,N_9468);
nand U9764 (N_9764,N_9592,N_9539);
or U9765 (N_9765,N_9306,N_9427);
and U9766 (N_9766,N_9517,N_9235);
and U9767 (N_9767,N_9310,N_9416);
nand U9768 (N_9768,N_9554,N_9384);
xor U9769 (N_9769,N_9280,N_9270);
nand U9770 (N_9770,N_9229,N_9214);
or U9771 (N_9771,N_9413,N_9341);
nand U9772 (N_9772,N_9326,N_9563);
or U9773 (N_9773,N_9337,N_9216);
nor U9774 (N_9774,N_9450,N_9532);
or U9775 (N_9775,N_9382,N_9491);
nor U9776 (N_9776,N_9330,N_9361);
nor U9777 (N_9777,N_9476,N_9325);
nand U9778 (N_9778,N_9220,N_9266);
and U9779 (N_9779,N_9211,N_9480);
nor U9780 (N_9780,N_9254,N_9569);
or U9781 (N_9781,N_9304,N_9272);
nand U9782 (N_9782,N_9568,N_9471);
nand U9783 (N_9783,N_9470,N_9503);
or U9784 (N_9784,N_9319,N_9433);
nor U9785 (N_9785,N_9575,N_9462);
nor U9786 (N_9786,N_9315,N_9344);
and U9787 (N_9787,N_9441,N_9595);
and U9788 (N_9788,N_9332,N_9268);
xor U9789 (N_9789,N_9236,N_9375);
xor U9790 (N_9790,N_9447,N_9492);
nor U9791 (N_9791,N_9558,N_9578);
and U9792 (N_9792,N_9291,N_9403);
and U9793 (N_9793,N_9251,N_9477);
xor U9794 (N_9794,N_9405,N_9312);
and U9795 (N_9795,N_9529,N_9356);
nand U9796 (N_9796,N_9588,N_9302);
and U9797 (N_9797,N_9564,N_9210);
xnor U9798 (N_9798,N_9521,N_9322);
and U9799 (N_9799,N_9479,N_9282);
nor U9800 (N_9800,N_9390,N_9260);
xnor U9801 (N_9801,N_9365,N_9301);
nor U9802 (N_9802,N_9375,N_9578);
and U9803 (N_9803,N_9426,N_9385);
or U9804 (N_9804,N_9383,N_9465);
and U9805 (N_9805,N_9368,N_9591);
xnor U9806 (N_9806,N_9278,N_9235);
nand U9807 (N_9807,N_9488,N_9262);
nor U9808 (N_9808,N_9368,N_9373);
and U9809 (N_9809,N_9338,N_9372);
and U9810 (N_9810,N_9207,N_9406);
nor U9811 (N_9811,N_9502,N_9202);
nand U9812 (N_9812,N_9348,N_9309);
nor U9813 (N_9813,N_9513,N_9474);
and U9814 (N_9814,N_9581,N_9434);
and U9815 (N_9815,N_9380,N_9343);
nor U9816 (N_9816,N_9584,N_9352);
nand U9817 (N_9817,N_9419,N_9550);
or U9818 (N_9818,N_9389,N_9230);
or U9819 (N_9819,N_9202,N_9519);
nand U9820 (N_9820,N_9364,N_9344);
xnor U9821 (N_9821,N_9305,N_9403);
or U9822 (N_9822,N_9405,N_9495);
nand U9823 (N_9823,N_9227,N_9472);
and U9824 (N_9824,N_9393,N_9205);
and U9825 (N_9825,N_9505,N_9570);
or U9826 (N_9826,N_9461,N_9222);
or U9827 (N_9827,N_9507,N_9324);
nand U9828 (N_9828,N_9427,N_9487);
xor U9829 (N_9829,N_9272,N_9494);
xor U9830 (N_9830,N_9524,N_9420);
and U9831 (N_9831,N_9501,N_9353);
nor U9832 (N_9832,N_9253,N_9590);
nand U9833 (N_9833,N_9517,N_9251);
and U9834 (N_9834,N_9351,N_9520);
or U9835 (N_9835,N_9517,N_9322);
nor U9836 (N_9836,N_9492,N_9230);
nor U9837 (N_9837,N_9522,N_9436);
nor U9838 (N_9838,N_9519,N_9410);
and U9839 (N_9839,N_9323,N_9394);
xnor U9840 (N_9840,N_9490,N_9262);
and U9841 (N_9841,N_9271,N_9374);
nand U9842 (N_9842,N_9520,N_9228);
nand U9843 (N_9843,N_9366,N_9454);
and U9844 (N_9844,N_9584,N_9275);
nor U9845 (N_9845,N_9520,N_9484);
and U9846 (N_9846,N_9486,N_9461);
nand U9847 (N_9847,N_9255,N_9327);
or U9848 (N_9848,N_9548,N_9410);
xor U9849 (N_9849,N_9367,N_9200);
or U9850 (N_9850,N_9595,N_9264);
nand U9851 (N_9851,N_9390,N_9494);
xor U9852 (N_9852,N_9498,N_9547);
nand U9853 (N_9853,N_9409,N_9495);
and U9854 (N_9854,N_9291,N_9256);
nor U9855 (N_9855,N_9388,N_9507);
nand U9856 (N_9856,N_9384,N_9340);
nor U9857 (N_9857,N_9510,N_9514);
nand U9858 (N_9858,N_9494,N_9457);
or U9859 (N_9859,N_9339,N_9405);
or U9860 (N_9860,N_9591,N_9382);
or U9861 (N_9861,N_9331,N_9532);
nor U9862 (N_9862,N_9540,N_9411);
nor U9863 (N_9863,N_9598,N_9461);
and U9864 (N_9864,N_9439,N_9549);
nand U9865 (N_9865,N_9517,N_9334);
or U9866 (N_9866,N_9462,N_9401);
or U9867 (N_9867,N_9294,N_9404);
nand U9868 (N_9868,N_9384,N_9363);
and U9869 (N_9869,N_9591,N_9309);
nor U9870 (N_9870,N_9306,N_9495);
nand U9871 (N_9871,N_9536,N_9559);
or U9872 (N_9872,N_9212,N_9421);
nand U9873 (N_9873,N_9563,N_9262);
and U9874 (N_9874,N_9265,N_9450);
nor U9875 (N_9875,N_9226,N_9544);
nor U9876 (N_9876,N_9389,N_9329);
or U9877 (N_9877,N_9520,N_9451);
or U9878 (N_9878,N_9591,N_9575);
xnor U9879 (N_9879,N_9269,N_9228);
xor U9880 (N_9880,N_9455,N_9296);
nand U9881 (N_9881,N_9543,N_9427);
xnor U9882 (N_9882,N_9396,N_9534);
or U9883 (N_9883,N_9364,N_9361);
and U9884 (N_9884,N_9487,N_9423);
or U9885 (N_9885,N_9200,N_9461);
nand U9886 (N_9886,N_9458,N_9583);
nand U9887 (N_9887,N_9349,N_9237);
or U9888 (N_9888,N_9248,N_9356);
and U9889 (N_9889,N_9219,N_9332);
xor U9890 (N_9890,N_9484,N_9580);
or U9891 (N_9891,N_9544,N_9242);
xnor U9892 (N_9892,N_9449,N_9393);
xnor U9893 (N_9893,N_9468,N_9351);
xor U9894 (N_9894,N_9205,N_9550);
nor U9895 (N_9895,N_9208,N_9364);
xor U9896 (N_9896,N_9472,N_9392);
xor U9897 (N_9897,N_9533,N_9226);
nand U9898 (N_9898,N_9217,N_9362);
nor U9899 (N_9899,N_9502,N_9330);
nand U9900 (N_9900,N_9435,N_9249);
or U9901 (N_9901,N_9462,N_9204);
and U9902 (N_9902,N_9462,N_9456);
or U9903 (N_9903,N_9425,N_9253);
nand U9904 (N_9904,N_9262,N_9224);
and U9905 (N_9905,N_9400,N_9247);
nand U9906 (N_9906,N_9342,N_9309);
and U9907 (N_9907,N_9572,N_9426);
xor U9908 (N_9908,N_9440,N_9282);
and U9909 (N_9909,N_9315,N_9386);
nand U9910 (N_9910,N_9262,N_9433);
xnor U9911 (N_9911,N_9543,N_9585);
nor U9912 (N_9912,N_9461,N_9298);
and U9913 (N_9913,N_9440,N_9352);
and U9914 (N_9914,N_9598,N_9527);
and U9915 (N_9915,N_9220,N_9556);
and U9916 (N_9916,N_9595,N_9297);
nand U9917 (N_9917,N_9577,N_9370);
and U9918 (N_9918,N_9491,N_9214);
or U9919 (N_9919,N_9307,N_9523);
nor U9920 (N_9920,N_9460,N_9361);
and U9921 (N_9921,N_9406,N_9427);
xor U9922 (N_9922,N_9402,N_9487);
or U9923 (N_9923,N_9572,N_9542);
nand U9924 (N_9924,N_9533,N_9333);
nor U9925 (N_9925,N_9566,N_9248);
or U9926 (N_9926,N_9519,N_9398);
nor U9927 (N_9927,N_9588,N_9547);
xnor U9928 (N_9928,N_9257,N_9391);
and U9929 (N_9929,N_9436,N_9209);
xor U9930 (N_9930,N_9398,N_9324);
and U9931 (N_9931,N_9504,N_9386);
or U9932 (N_9932,N_9461,N_9403);
xnor U9933 (N_9933,N_9372,N_9342);
xnor U9934 (N_9934,N_9531,N_9241);
xnor U9935 (N_9935,N_9576,N_9598);
and U9936 (N_9936,N_9234,N_9555);
or U9937 (N_9937,N_9575,N_9502);
xor U9938 (N_9938,N_9595,N_9340);
nand U9939 (N_9939,N_9592,N_9233);
nand U9940 (N_9940,N_9419,N_9276);
xor U9941 (N_9941,N_9303,N_9347);
nor U9942 (N_9942,N_9444,N_9277);
xnor U9943 (N_9943,N_9506,N_9554);
xnor U9944 (N_9944,N_9347,N_9481);
or U9945 (N_9945,N_9332,N_9391);
nor U9946 (N_9946,N_9416,N_9235);
or U9947 (N_9947,N_9465,N_9459);
and U9948 (N_9948,N_9501,N_9211);
xor U9949 (N_9949,N_9432,N_9486);
and U9950 (N_9950,N_9583,N_9363);
nor U9951 (N_9951,N_9264,N_9523);
or U9952 (N_9952,N_9297,N_9563);
nor U9953 (N_9953,N_9375,N_9510);
xor U9954 (N_9954,N_9338,N_9364);
nor U9955 (N_9955,N_9586,N_9576);
nor U9956 (N_9956,N_9330,N_9373);
and U9957 (N_9957,N_9580,N_9259);
xor U9958 (N_9958,N_9337,N_9332);
nor U9959 (N_9959,N_9465,N_9494);
and U9960 (N_9960,N_9493,N_9217);
or U9961 (N_9961,N_9253,N_9592);
nand U9962 (N_9962,N_9464,N_9429);
nor U9963 (N_9963,N_9592,N_9417);
and U9964 (N_9964,N_9571,N_9355);
or U9965 (N_9965,N_9393,N_9485);
nand U9966 (N_9966,N_9572,N_9514);
or U9967 (N_9967,N_9360,N_9592);
nand U9968 (N_9968,N_9487,N_9412);
nand U9969 (N_9969,N_9535,N_9507);
xnor U9970 (N_9970,N_9416,N_9342);
nor U9971 (N_9971,N_9435,N_9529);
and U9972 (N_9972,N_9351,N_9389);
and U9973 (N_9973,N_9447,N_9499);
xnor U9974 (N_9974,N_9211,N_9503);
nor U9975 (N_9975,N_9352,N_9312);
nand U9976 (N_9976,N_9412,N_9471);
or U9977 (N_9977,N_9442,N_9244);
or U9978 (N_9978,N_9419,N_9387);
xor U9979 (N_9979,N_9551,N_9593);
or U9980 (N_9980,N_9268,N_9524);
nor U9981 (N_9981,N_9400,N_9328);
nand U9982 (N_9982,N_9268,N_9365);
or U9983 (N_9983,N_9499,N_9531);
nand U9984 (N_9984,N_9481,N_9258);
nor U9985 (N_9985,N_9483,N_9576);
and U9986 (N_9986,N_9430,N_9544);
and U9987 (N_9987,N_9293,N_9542);
xor U9988 (N_9988,N_9317,N_9383);
nor U9989 (N_9989,N_9394,N_9388);
nor U9990 (N_9990,N_9200,N_9550);
nor U9991 (N_9991,N_9569,N_9387);
or U9992 (N_9992,N_9305,N_9427);
and U9993 (N_9993,N_9443,N_9580);
xnor U9994 (N_9994,N_9554,N_9456);
xnor U9995 (N_9995,N_9228,N_9398);
xnor U9996 (N_9996,N_9257,N_9521);
nor U9997 (N_9997,N_9423,N_9287);
nand U9998 (N_9998,N_9441,N_9213);
nand U9999 (N_9999,N_9509,N_9329);
xor U10000 (N_10000,N_9758,N_9749);
nor U10001 (N_10001,N_9848,N_9654);
nand U10002 (N_10002,N_9771,N_9665);
xnor U10003 (N_10003,N_9985,N_9686);
or U10004 (N_10004,N_9897,N_9876);
nand U10005 (N_10005,N_9925,N_9698);
or U10006 (N_10006,N_9933,N_9934);
and U10007 (N_10007,N_9618,N_9647);
xnor U10008 (N_10008,N_9886,N_9947);
nand U10009 (N_10009,N_9645,N_9676);
nor U10010 (N_10010,N_9820,N_9995);
nor U10011 (N_10011,N_9940,N_9778);
nand U10012 (N_10012,N_9720,N_9938);
or U10013 (N_10013,N_9612,N_9866);
xnor U10014 (N_10014,N_9751,N_9785);
and U10015 (N_10015,N_9679,N_9917);
nand U10016 (N_10016,N_9816,N_9712);
or U10017 (N_10017,N_9601,N_9685);
nor U10018 (N_10018,N_9950,N_9682);
xor U10019 (N_10019,N_9613,N_9863);
nor U10020 (N_10020,N_9971,N_9770);
xnor U10021 (N_10021,N_9703,N_9630);
xor U10022 (N_10022,N_9641,N_9834);
nand U10023 (N_10023,N_9677,N_9903);
or U10024 (N_10024,N_9623,N_9632);
and U10025 (N_10025,N_9757,N_9881);
or U10026 (N_10026,N_9901,N_9766);
or U10027 (N_10027,N_9631,N_9616);
xnor U10028 (N_10028,N_9617,N_9857);
or U10029 (N_10029,N_9775,N_9872);
nor U10030 (N_10030,N_9747,N_9941);
and U10031 (N_10031,N_9772,N_9896);
and U10032 (N_10032,N_9909,N_9852);
nor U10033 (N_10033,N_9721,N_9691);
nor U10034 (N_10034,N_9935,N_9688);
and U10035 (N_10035,N_9851,N_9642);
nand U10036 (N_10036,N_9847,N_9798);
or U10037 (N_10037,N_9828,N_9756);
nand U10038 (N_10038,N_9680,N_9754);
and U10039 (N_10039,N_9837,N_9692);
and U10040 (N_10040,N_9982,N_9821);
or U10041 (N_10041,N_9957,N_9892);
and U10042 (N_10042,N_9920,N_9690);
and U10043 (N_10043,N_9929,N_9968);
and U10044 (N_10044,N_9697,N_9998);
nor U10045 (N_10045,N_9625,N_9651);
and U10046 (N_10046,N_9843,N_9604);
and U10047 (N_10047,N_9669,N_9639);
or U10048 (N_10048,N_9660,N_9709);
nor U10049 (N_10049,N_9890,N_9621);
nand U10050 (N_10050,N_9726,N_9769);
or U10051 (N_10051,N_9974,N_9823);
nor U10052 (N_10052,N_9888,N_9755);
or U10053 (N_10053,N_9659,N_9803);
or U10054 (N_10054,N_9839,N_9975);
nand U10055 (N_10055,N_9708,N_9656);
nor U10056 (N_10056,N_9603,N_9814);
nand U10057 (N_10057,N_9646,N_9740);
and U10058 (N_10058,N_9790,N_9629);
or U10059 (N_10059,N_9889,N_9965);
xor U10060 (N_10060,N_9996,N_9614);
xor U10061 (N_10061,N_9915,N_9681);
xnor U10062 (N_10062,N_9817,N_9627);
nor U10063 (N_10063,N_9945,N_9786);
xor U10064 (N_10064,N_9990,N_9832);
or U10065 (N_10065,N_9838,N_9979);
and U10066 (N_10066,N_9622,N_9811);
nand U10067 (N_10067,N_9602,N_9663);
nand U10068 (N_10068,N_9806,N_9735);
xnor U10069 (N_10069,N_9921,N_9760);
nand U10070 (N_10070,N_9946,N_9846);
or U10071 (N_10071,N_9804,N_9661);
xnor U10072 (N_10072,N_9894,N_9900);
nor U10073 (N_10073,N_9650,N_9672);
nor U10074 (N_10074,N_9689,N_9865);
xor U10075 (N_10075,N_9694,N_9992);
nor U10076 (N_10076,N_9981,N_9952);
nand U10077 (N_10077,N_9737,N_9919);
xor U10078 (N_10078,N_9791,N_9729);
or U10079 (N_10079,N_9908,N_9849);
xor U10080 (N_10080,N_9643,N_9706);
nor U10081 (N_10081,N_9931,N_9833);
and U10082 (N_10082,N_9809,N_9731);
or U10083 (N_10083,N_9668,N_9687);
nor U10084 (N_10084,N_9969,N_9793);
and U10085 (N_10085,N_9910,N_9750);
xor U10086 (N_10086,N_9902,N_9762);
or U10087 (N_10087,N_9943,N_9767);
nand U10088 (N_10088,N_9875,N_9815);
or U10089 (N_10089,N_9928,N_9836);
nor U10090 (N_10090,N_9855,N_9776);
or U10091 (N_10091,N_9714,N_9858);
or U10092 (N_10092,N_9695,N_9882);
and U10093 (N_10093,N_9862,N_9779);
xor U10094 (N_10094,N_9609,N_9683);
or U10095 (N_10095,N_9906,N_9784);
and U10096 (N_10096,N_9606,N_9781);
xnor U10097 (N_10097,N_9655,N_9861);
nand U10098 (N_10098,N_9805,N_9727);
nor U10099 (N_10099,N_9693,N_9710);
nor U10100 (N_10100,N_9701,N_9746);
or U10101 (N_10101,N_9895,N_9819);
and U10102 (N_10102,N_9905,N_9640);
and U10103 (N_10103,N_9853,N_9700);
nor U10104 (N_10104,N_9923,N_9671);
and U10105 (N_10105,N_9624,N_9759);
nand U10106 (N_10106,N_9966,N_9868);
nor U10107 (N_10107,N_9796,N_9728);
xnor U10108 (N_10108,N_9818,N_9885);
xor U10109 (N_10109,N_9788,N_9842);
and U10110 (N_10110,N_9761,N_9667);
and U10111 (N_10111,N_9801,N_9636);
xor U10112 (N_10112,N_9730,N_9964);
and U10113 (N_10113,N_9673,N_9955);
nor U10114 (N_10114,N_9711,N_9999);
and U10115 (N_10115,N_9891,N_9829);
or U10116 (N_10116,N_9717,N_9652);
and U10117 (N_10117,N_9987,N_9954);
or U10118 (N_10118,N_9826,N_9963);
nand U10119 (N_10119,N_9744,N_9962);
and U10120 (N_10120,N_9867,N_9926);
xor U10121 (N_10121,N_9997,N_9768);
nor U10122 (N_10122,N_9970,N_9653);
or U10123 (N_10123,N_9907,N_9880);
or U10124 (N_10124,N_9958,N_9859);
and U10125 (N_10125,N_9951,N_9878);
nor U10126 (N_10126,N_9600,N_9854);
nand U10127 (N_10127,N_9719,N_9989);
or U10128 (N_10128,N_9684,N_9723);
and U10129 (N_10129,N_9718,N_9738);
or U10130 (N_10130,N_9637,N_9893);
xnor U10131 (N_10131,N_9911,N_9845);
or U10132 (N_10132,N_9739,N_9939);
or U10133 (N_10133,N_9936,N_9733);
nand U10134 (N_10134,N_9812,N_9944);
and U10135 (N_10135,N_9961,N_9635);
nand U10136 (N_10136,N_9850,N_9972);
xor U10137 (N_10137,N_9658,N_9741);
nor U10138 (N_10138,N_9831,N_9914);
xor U10139 (N_10139,N_9869,N_9634);
or U10140 (N_10140,N_9977,N_9777);
or U10141 (N_10141,N_9976,N_9633);
nand U10142 (N_10142,N_9887,N_9649);
nor U10143 (N_10143,N_9664,N_9874);
xor U10144 (N_10144,N_9657,N_9813);
or U10145 (N_10145,N_9991,N_9644);
or U10146 (N_10146,N_9620,N_9674);
nor U10147 (N_10147,N_9835,N_9864);
nor U10148 (N_10148,N_9988,N_9799);
and U10149 (N_10149,N_9898,N_9752);
nand U10150 (N_10150,N_9716,N_9994);
nand U10151 (N_10151,N_9678,N_9619);
nand U10152 (N_10152,N_9841,N_9794);
and U10153 (N_10153,N_9763,N_9871);
xor U10154 (N_10154,N_9774,N_9980);
or U10155 (N_10155,N_9610,N_9715);
xnor U10156 (N_10156,N_9879,N_9748);
nand U10157 (N_10157,N_9722,N_9840);
xor U10158 (N_10158,N_9916,N_9912);
nand U10159 (N_10159,N_9802,N_9960);
xor U10160 (N_10160,N_9883,N_9666);
and U10161 (N_10161,N_9899,N_9795);
or U10162 (N_10162,N_9808,N_9745);
nand U10163 (N_10163,N_9725,N_9993);
xnor U10164 (N_10164,N_9662,N_9918);
or U10165 (N_10165,N_9670,N_9932);
and U10166 (N_10166,N_9825,N_9611);
xnor U10167 (N_10167,N_9705,N_9856);
xnor U10168 (N_10168,N_9827,N_9956);
or U10169 (N_10169,N_9713,N_9922);
xor U10170 (N_10170,N_9904,N_9967);
or U10171 (N_10171,N_9764,N_9927);
nor U10172 (N_10172,N_9884,N_9734);
nor U10173 (N_10173,N_9983,N_9628);
nand U10174 (N_10174,N_9949,N_9780);
nor U10175 (N_10175,N_9984,N_9810);
and U10176 (N_10176,N_9844,N_9870);
nor U10177 (N_10177,N_9732,N_9787);
nor U10178 (N_10178,N_9959,N_9789);
xnor U10179 (N_10179,N_9800,N_9792);
nand U10180 (N_10180,N_9913,N_9830);
nor U10181 (N_10181,N_9702,N_9675);
xnor U10182 (N_10182,N_9953,N_9807);
xnor U10183 (N_10183,N_9773,N_9948);
nand U10184 (N_10184,N_9607,N_9782);
or U10185 (N_10185,N_9930,N_9605);
nand U10186 (N_10186,N_9724,N_9942);
nand U10187 (N_10187,N_9824,N_9797);
or U10188 (N_10188,N_9626,N_9742);
and U10189 (N_10189,N_9765,N_9783);
or U10190 (N_10190,N_9743,N_9699);
xnor U10191 (N_10191,N_9638,N_9924);
nand U10192 (N_10192,N_9707,N_9736);
nor U10193 (N_10193,N_9615,N_9978);
nor U10194 (N_10194,N_9986,N_9822);
and U10195 (N_10195,N_9648,N_9860);
nor U10196 (N_10196,N_9973,N_9753);
nand U10197 (N_10197,N_9877,N_9937);
nor U10198 (N_10198,N_9696,N_9873);
or U10199 (N_10199,N_9704,N_9608);
or U10200 (N_10200,N_9622,N_9831);
xor U10201 (N_10201,N_9711,N_9604);
or U10202 (N_10202,N_9719,N_9795);
and U10203 (N_10203,N_9942,N_9800);
and U10204 (N_10204,N_9893,N_9796);
xor U10205 (N_10205,N_9833,N_9614);
nand U10206 (N_10206,N_9767,N_9964);
and U10207 (N_10207,N_9617,N_9842);
nor U10208 (N_10208,N_9745,N_9769);
or U10209 (N_10209,N_9602,N_9919);
and U10210 (N_10210,N_9788,N_9694);
nor U10211 (N_10211,N_9740,N_9704);
or U10212 (N_10212,N_9832,N_9945);
nand U10213 (N_10213,N_9938,N_9658);
xnor U10214 (N_10214,N_9842,N_9894);
nand U10215 (N_10215,N_9913,N_9824);
and U10216 (N_10216,N_9801,N_9774);
nand U10217 (N_10217,N_9729,N_9929);
xor U10218 (N_10218,N_9679,N_9716);
or U10219 (N_10219,N_9605,N_9789);
or U10220 (N_10220,N_9933,N_9889);
and U10221 (N_10221,N_9771,N_9704);
or U10222 (N_10222,N_9751,N_9965);
nor U10223 (N_10223,N_9783,N_9854);
and U10224 (N_10224,N_9917,N_9992);
nand U10225 (N_10225,N_9909,N_9605);
xnor U10226 (N_10226,N_9737,N_9645);
nand U10227 (N_10227,N_9631,N_9800);
nand U10228 (N_10228,N_9886,N_9985);
or U10229 (N_10229,N_9915,N_9673);
and U10230 (N_10230,N_9911,N_9721);
and U10231 (N_10231,N_9791,N_9966);
nand U10232 (N_10232,N_9621,N_9887);
nand U10233 (N_10233,N_9643,N_9662);
and U10234 (N_10234,N_9803,N_9887);
xnor U10235 (N_10235,N_9618,N_9792);
nand U10236 (N_10236,N_9847,N_9691);
xor U10237 (N_10237,N_9864,N_9691);
and U10238 (N_10238,N_9801,N_9833);
xnor U10239 (N_10239,N_9792,N_9645);
nand U10240 (N_10240,N_9637,N_9785);
nor U10241 (N_10241,N_9617,N_9608);
or U10242 (N_10242,N_9887,N_9787);
xnor U10243 (N_10243,N_9641,N_9653);
xnor U10244 (N_10244,N_9934,N_9831);
and U10245 (N_10245,N_9806,N_9817);
nor U10246 (N_10246,N_9815,N_9694);
or U10247 (N_10247,N_9790,N_9897);
and U10248 (N_10248,N_9803,N_9660);
xnor U10249 (N_10249,N_9619,N_9673);
or U10250 (N_10250,N_9813,N_9871);
nand U10251 (N_10251,N_9777,N_9944);
nor U10252 (N_10252,N_9641,N_9628);
nor U10253 (N_10253,N_9895,N_9684);
and U10254 (N_10254,N_9643,N_9631);
nor U10255 (N_10255,N_9902,N_9874);
nand U10256 (N_10256,N_9809,N_9928);
and U10257 (N_10257,N_9948,N_9970);
and U10258 (N_10258,N_9704,N_9861);
nor U10259 (N_10259,N_9788,N_9750);
xnor U10260 (N_10260,N_9607,N_9818);
nand U10261 (N_10261,N_9762,N_9751);
or U10262 (N_10262,N_9898,N_9803);
nor U10263 (N_10263,N_9873,N_9712);
or U10264 (N_10264,N_9834,N_9625);
nand U10265 (N_10265,N_9744,N_9632);
nor U10266 (N_10266,N_9692,N_9882);
nand U10267 (N_10267,N_9636,N_9893);
nor U10268 (N_10268,N_9765,N_9841);
nand U10269 (N_10269,N_9840,N_9976);
nor U10270 (N_10270,N_9772,N_9828);
nand U10271 (N_10271,N_9855,N_9791);
xor U10272 (N_10272,N_9733,N_9742);
or U10273 (N_10273,N_9987,N_9614);
nand U10274 (N_10274,N_9663,N_9893);
and U10275 (N_10275,N_9947,N_9789);
xnor U10276 (N_10276,N_9782,N_9698);
xor U10277 (N_10277,N_9803,N_9877);
nor U10278 (N_10278,N_9944,N_9875);
and U10279 (N_10279,N_9893,N_9720);
nand U10280 (N_10280,N_9995,N_9880);
or U10281 (N_10281,N_9611,N_9878);
and U10282 (N_10282,N_9654,N_9635);
nor U10283 (N_10283,N_9967,N_9733);
nand U10284 (N_10284,N_9620,N_9896);
xor U10285 (N_10285,N_9715,N_9871);
nand U10286 (N_10286,N_9967,N_9870);
or U10287 (N_10287,N_9646,N_9601);
nand U10288 (N_10288,N_9679,N_9722);
nor U10289 (N_10289,N_9908,N_9675);
nor U10290 (N_10290,N_9612,N_9706);
or U10291 (N_10291,N_9731,N_9912);
nand U10292 (N_10292,N_9889,N_9630);
or U10293 (N_10293,N_9769,N_9683);
or U10294 (N_10294,N_9995,N_9666);
xor U10295 (N_10295,N_9812,N_9892);
xnor U10296 (N_10296,N_9938,N_9782);
xor U10297 (N_10297,N_9739,N_9865);
and U10298 (N_10298,N_9623,N_9943);
xnor U10299 (N_10299,N_9778,N_9909);
nor U10300 (N_10300,N_9895,N_9954);
or U10301 (N_10301,N_9736,N_9888);
nand U10302 (N_10302,N_9640,N_9626);
and U10303 (N_10303,N_9666,N_9917);
xnor U10304 (N_10304,N_9767,N_9966);
xor U10305 (N_10305,N_9695,N_9666);
and U10306 (N_10306,N_9735,N_9867);
and U10307 (N_10307,N_9997,N_9949);
nor U10308 (N_10308,N_9715,N_9970);
or U10309 (N_10309,N_9895,N_9992);
nand U10310 (N_10310,N_9944,N_9986);
or U10311 (N_10311,N_9818,N_9811);
and U10312 (N_10312,N_9956,N_9614);
nor U10313 (N_10313,N_9787,N_9912);
and U10314 (N_10314,N_9831,N_9997);
nor U10315 (N_10315,N_9775,N_9747);
nor U10316 (N_10316,N_9758,N_9851);
xor U10317 (N_10317,N_9718,N_9918);
and U10318 (N_10318,N_9773,N_9945);
xor U10319 (N_10319,N_9954,N_9781);
and U10320 (N_10320,N_9735,N_9951);
or U10321 (N_10321,N_9939,N_9838);
nor U10322 (N_10322,N_9763,N_9794);
nor U10323 (N_10323,N_9619,N_9775);
nor U10324 (N_10324,N_9724,N_9993);
and U10325 (N_10325,N_9736,N_9843);
nand U10326 (N_10326,N_9898,N_9727);
xor U10327 (N_10327,N_9998,N_9765);
nand U10328 (N_10328,N_9732,N_9819);
xor U10329 (N_10329,N_9836,N_9612);
and U10330 (N_10330,N_9703,N_9738);
and U10331 (N_10331,N_9650,N_9715);
xor U10332 (N_10332,N_9826,N_9662);
nand U10333 (N_10333,N_9942,N_9927);
or U10334 (N_10334,N_9912,N_9822);
xor U10335 (N_10335,N_9836,N_9973);
nor U10336 (N_10336,N_9747,N_9791);
nand U10337 (N_10337,N_9752,N_9934);
nand U10338 (N_10338,N_9767,N_9917);
nor U10339 (N_10339,N_9752,N_9725);
and U10340 (N_10340,N_9671,N_9850);
or U10341 (N_10341,N_9748,N_9769);
and U10342 (N_10342,N_9869,N_9695);
nor U10343 (N_10343,N_9962,N_9781);
xor U10344 (N_10344,N_9612,N_9899);
or U10345 (N_10345,N_9878,N_9749);
nand U10346 (N_10346,N_9843,N_9688);
or U10347 (N_10347,N_9790,N_9760);
or U10348 (N_10348,N_9871,N_9669);
nor U10349 (N_10349,N_9903,N_9852);
and U10350 (N_10350,N_9966,N_9996);
xor U10351 (N_10351,N_9790,N_9781);
and U10352 (N_10352,N_9816,N_9961);
nor U10353 (N_10353,N_9704,N_9828);
nand U10354 (N_10354,N_9909,N_9952);
nand U10355 (N_10355,N_9887,N_9725);
nor U10356 (N_10356,N_9779,N_9948);
nor U10357 (N_10357,N_9718,N_9651);
nand U10358 (N_10358,N_9766,N_9974);
and U10359 (N_10359,N_9693,N_9677);
nor U10360 (N_10360,N_9612,N_9676);
or U10361 (N_10361,N_9631,N_9922);
and U10362 (N_10362,N_9707,N_9765);
or U10363 (N_10363,N_9693,N_9616);
nand U10364 (N_10364,N_9632,N_9912);
or U10365 (N_10365,N_9735,N_9944);
or U10366 (N_10366,N_9665,N_9941);
nand U10367 (N_10367,N_9723,N_9898);
xor U10368 (N_10368,N_9618,N_9622);
nand U10369 (N_10369,N_9836,N_9695);
or U10370 (N_10370,N_9887,N_9702);
and U10371 (N_10371,N_9632,N_9671);
or U10372 (N_10372,N_9657,N_9925);
xor U10373 (N_10373,N_9724,N_9636);
nand U10374 (N_10374,N_9749,N_9921);
xor U10375 (N_10375,N_9884,N_9602);
nand U10376 (N_10376,N_9825,N_9954);
nor U10377 (N_10377,N_9861,N_9972);
nand U10378 (N_10378,N_9981,N_9943);
nor U10379 (N_10379,N_9768,N_9818);
nand U10380 (N_10380,N_9933,N_9827);
and U10381 (N_10381,N_9894,N_9662);
nor U10382 (N_10382,N_9664,N_9896);
xnor U10383 (N_10383,N_9789,N_9934);
nor U10384 (N_10384,N_9971,N_9974);
xnor U10385 (N_10385,N_9686,N_9771);
or U10386 (N_10386,N_9943,N_9923);
nor U10387 (N_10387,N_9778,N_9782);
or U10388 (N_10388,N_9879,N_9972);
nor U10389 (N_10389,N_9627,N_9844);
nand U10390 (N_10390,N_9630,N_9914);
and U10391 (N_10391,N_9834,N_9793);
nand U10392 (N_10392,N_9846,N_9934);
nand U10393 (N_10393,N_9664,N_9826);
nand U10394 (N_10394,N_9786,N_9627);
xnor U10395 (N_10395,N_9914,N_9767);
or U10396 (N_10396,N_9855,N_9963);
xor U10397 (N_10397,N_9758,N_9802);
nand U10398 (N_10398,N_9660,N_9846);
xnor U10399 (N_10399,N_9928,N_9761);
or U10400 (N_10400,N_10387,N_10389);
and U10401 (N_10401,N_10314,N_10143);
or U10402 (N_10402,N_10119,N_10173);
xnor U10403 (N_10403,N_10328,N_10368);
xnor U10404 (N_10404,N_10215,N_10019);
and U10405 (N_10405,N_10185,N_10379);
nand U10406 (N_10406,N_10058,N_10226);
nor U10407 (N_10407,N_10008,N_10045);
nor U10408 (N_10408,N_10041,N_10179);
and U10409 (N_10409,N_10010,N_10157);
and U10410 (N_10410,N_10347,N_10337);
nor U10411 (N_10411,N_10395,N_10114);
nand U10412 (N_10412,N_10305,N_10331);
nor U10413 (N_10413,N_10014,N_10021);
or U10414 (N_10414,N_10348,N_10269);
xnor U10415 (N_10415,N_10077,N_10040);
xnor U10416 (N_10416,N_10270,N_10346);
nand U10417 (N_10417,N_10281,N_10022);
and U10418 (N_10418,N_10304,N_10246);
and U10419 (N_10419,N_10384,N_10311);
or U10420 (N_10420,N_10219,N_10250);
xor U10421 (N_10421,N_10072,N_10096);
and U10422 (N_10422,N_10027,N_10018);
and U10423 (N_10423,N_10135,N_10159);
nand U10424 (N_10424,N_10391,N_10030);
xor U10425 (N_10425,N_10193,N_10071);
or U10426 (N_10426,N_10213,N_10171);
nand U10427 (N_10427,N_10017,N_10189);
xor U10428 (N_10428,N_10342,N_10098);
xnor U10429 (N_10429,N_10266,N_10028);
nor U10430 (N_10430,N_10383,N_10218);
xnor U10431 (N_10431,N_10181,N_10282);
and U10432 (N_10432,N_10099,N_10013);
xor U10433 (N_10433,N_10276,N_10394);
and U10434 (N_10434,N_10116,N_10286);
xnor U10435 (N_10435,N_10052,N_10024);
or U10436 (N_10436,N_10169,N_10122);
and U10437 (N_10437,N_10367,N_10111);
or U10438 (N_10438,N_10128,N_10020);
xor U10439 (N_10439,N_10065,N_10117);
nor U10440 (N_10440,N_10262,N_10325);
nand U10441 (N_10441,N_10032,N_10036);
or U10442 (N_10442,N_10103,N_10156);
or U10443 (N_10443,N_10088,N_10344);
and U10444 (N_10444,N_10033,N_10338);
nand U10445 (N_10445,N_10035,N_10170);
nor U10446 (N_10446,N_10000,N_10222);
xor U10447 (N_10447,N_10086,N_10306);
xnor U10448 (N_10448,N_10341,N_10320);
xor U10449 (N_10449,N_10399,N_10158);
or U10450 (N_10450,N_10199,N_10129);
and U10451 (N_10451,N_10073,N_10139);
xor U10452 (N_10452,N_10288,N_10313);
or U10453 (N_10453,N_10386,N_10121);
xnor U10454 (N_10454,N_10333,N_10370);
xor U10455 (N_10455,N_10049,N_10059);
and U10456 (N_10456,N_10090,N_10223);
nand U10457 (N_10457,N_10107,N_10130);
or U10458 (N_10458,N_10249,N_10228);
xnor U10459 (N_10459,N_10003,N_10234);
or U10460 (N_10460,N_10208,N_10132);
nor U10461 (N_10461,N_10070,N_10016);
or U10462 (N_10462,N_10258,N_10075);
xor U10463 (N_10463,N_10210,N_10082);
nand U10464 (N_10464,N_10069,N_10330);
xor U10465 (N_10465,N_10365,N_10211);
or U10466 (N_10466,N_10050,N_10067);
nor U10467 (N_10467,N_10293,N_10329);
or U10468 (N_10468,N_10340,N_10349);
or U10469 (N_10469,N_10160,N_10186);
and U10470 (N_10470,N_10155,N_10093);
and U10471 (N_10471,N_10255,N_10353);
xnor U10472 (N_10472,N_10298,N_10251);
or U10473 (N_10473,N_10264,N_10112);
nor U10474 (N_10474,N_10303,N_10083);
xnor U10475 (N_10475,N_10241,N_10007);
nand U10476 (N_10476,N_10163,N_10140);
or U10477 (N_10477,N_10108,N_10308);
and U10478 (N_10478,N_10361,N_10363);
or U10479 (N_10479,N_10369,N_10057);
nor U10480 (N_10480,N_10009,N_10180);
nand U10481 (N_10481,N_10081,N_10265);
or U10482 (N_10482,N_10292,N_10191);
xor U10483 (N_10483,N_10201,N_10378);
nor U10484 (N_10484,N_10060,N_10172);
nor U10485 (N_10485,N_10048,N_10183);
and U10486 (N_10486,N_10319,N_10147);
and U10487 (N_10487,N_10321,N_10287);
nand U10488 (N_10488,N_10166,N_10253);
nand U10489 (N_10489,N_10196,N_10327);
nor U10490 (N_10490,N_10230,N_10091);
or U10491 (N_10491,N_10373,N_10259);
nor U10492 (N_10492,N_10376,N_10203);
nor U10493 (N_10493,N_10026,N_10153);
or U10494 (N_10494,N_10056,N_10012);
nor U10495 (N_10495,N_10097,N_10233);
nor U10496 (N_10496,N_10221,N_10295);
xnor U10497 (N_10497,N_10209,N_10307);
or U10498 (N_10498,N_10377,N_10204);
nand U10499 (N_10499,N_10289,N_10053);
nor U10500 (N_10500,N_10388,N_10029);
and U10501 (N_10501,N_10165,N_10302);
and U10502 (N_10502,N_10089,N_10174);
xor U10503 (N_10503,N_10312,N_10225);
nor U10504 (N_10504,N_10146,N_10192);
nor U10505 (N_10505,N_10214,N_10125);
nand U10506 (N_10506,N_10274,N_10359);
or U10507 (N_10507,N_10212,N_10152);
and U10508 (N_10508,N_10120,N_10161);
and U10509 (N_10509,N_10002,N_10291);
or U10510 (N_10510,N_10127,N_10110);
or U10511 (N_10511,N_10323,N_10277);
nand U10512 (N_10512,N_10334,N_10038);
or U10513 (N_10513,N_10194,N_10123);
nand U10514 (N_10514,N_10094,N_10364);
xor U10515 (N_10515,N_10271,N_10336);
nor U10516 (N_10516,N_10006,N_10015);
xnor U10517 (N_10517,N_10380,N_10102);
and U10518 (N_10518,N_10118,N_10175);
nand U10519 (N_10519,N_10182,N_10248);
xor U10520 (N_10520,N_10243,N_10326);
nand U10521 (N_10521,N_10285,N_10142);
or U10522 (N_10522,N_10252,N_10245);
xnor U10523 (N_10523,N_10247,N_10109);
and U10524 (N_10524,N_10309,N_10134);
nand U10525 (N_10525,N_10374,N_10355);
nor U10526 (N_10526,N_10339,N_10239);
nor U10527 (N_10527,N_10263,N_10074);
and U10528 (N_10528,N_10138,N_10238);
and U10529 (N_10529,N_10188,N_10100);
or U10530 (N_10530,N_10352,N_10345);
and U10531 (N_10531,N_10316,N_10362);
or U10532 (N_10532,N_10106,N_10197);
xnor U10533 (N_10533,N_10240,N_10358);
and U10534 (N_10534,N_10244,N_10260);
or U10535 (N_10535,N_10136,N_10063);
nand U10536 (N_10536,N_10393,N_10350);
xor U10537 (N_10537,N_10084,N_10392);
nand U10538 (N_10538,N_10220,N_10356);
nand U10539 (N_10539,N_10137,N_10039);
and U10540 (N_10540,N_10124,N_10055);
nor U10541 (N_10541,N_10318,N_10062);
or U10542 (N_10542,N_10216,N_10343);
nor U10543 (N_10543,N_10275,N_10317);
xnor U10544 (N_10544,N_10200,N_10149);
nand U10545 (N_10545,N_10390,N_10080);
nand U10546 (N_10546,N_10202,N_10284);
nor U10547 (N_10547,N_10396,N_10372);
or U10548 (N_10548,N_10351,N_10354);
nor U10549 (N_10549,N_10066,N_10131);
xor U10550 (N_10550,N_10092,N_10294);
and U10551 (N_10551,N_10267,N_10068);
nand U10552 (N_10552,N_10104,N_10280);
xor U10553 (N_10553,N_10296,N_10207);
or U10554 (N_10554,N_10315,N_10261);
nand U10555 (N_10555,N_10300,N_10257);
and U10556 (N_10556,N_10278,N_10037);
nor U10557 (N_10557,N_10076,N_10005);
and U10558 (N_10558,N_10047,N_10232);
nand U10559 (N_10559,N_10256,N_10375);
or U10560 (N_10560,N_10187,N_10031);
and U10561 (N_10561,N_10335,N_10385);
and U10562 (N_10562,N_10004,N_10397);
xor U10563 (N_10563,N_10095,N_10101);
or U10564 (N_10564,N_10087,N_10001);
xnor U10565 (N_10565,N_10279,N_10217);
nor U10566 (N_10566,N_10398,N_10078);
nand U10567 (N_10567,N_10151,N_10023);
nor U10568 (N_10568,N_10310,N_10236);
and U10569 (N_10569,N_10042,N_10268);
and U10570 (N_10570,N_10043,N_10357);
xor U10571 (N_10571,N_10366,N_10150);
nand U10572 (N_10572,N_10167,N_10079);
nor U10573 (N_10573,N_10242,N_10061);
nor U10574 (N_10574,N_10113,N_10148);
nor U10575 (N_10575,N_10184,N_10141);
xor U10576 (N_10576,N_10332,N_10235);
nand U10577 (N_10577,N_10283,N_10085);
nand U10578 (N_10578,N_10381,N_10195);
xor U10579 (N_10579,N_10205,N_10322);
and U10580 (N_10580,N_10206,N_10299);
or U10581 (N_10581,N_10273,N_10168);
nor U10582 (N_10582,N_10178,N_10164);
nand U10583 (N_10583,N_10198,N_10231);
xnor U10584 (N_10584,N_10144,N_10224);
nor U10585 (N_10585,N_10301,N_10105);
or U10586 (N_10586,N_10237,N_10051);
nor U10587 (N_10587,N_10290,N_10177);
nor U10588 (N_10588,N_10025,N_10227);
nand U10589 (N_10589,N_10044,N_10126);
xor U10590 (N_10590,N_10145,N_10272);
nand U10591 (N_10591,N_10324,N_10064);
xor U10592 (N_10592,N_10254,N_10133);
nand U10593 (N_10593,N_10360,N_10034);
nor U10594 (N_10594,N_10054,N_10011);
or U10595 (N_10595,N_10176,N_10115);
or U10596 (N_10596,N_10382,N_10297);
nand U10597 (N_10597,N_10190,N_10229);
and U10598 (N_10598,N_10046,N_10371);
and U10599 (N_10599,N_10162,N_10154);
nand U10600 (N_10600,N_10072,N_10297);
nand U10601 (N_10601,N_10336,N_10115);
nor U10602 (N_10602,N_10292,N_10313);
nor U10603 (N_10603,N_10307,N_10095);
and U10604 (N_10604,N_10287,N_10208);
or U10605 (N_10605,N_10261,N_10349);
xor U10606 (N_10606,N_10003,N_10292);
nand U10607 (N_10607,N_10254,N_10087);
and U10608 (N_10608,N_10056,N_10214);
or U10609 (N_10609,N_10099,N_10126);
nor U10610 (N_10610,N_10096,N_10059);
nand U10611 (N_10611,N_10289,N_10131);
nand U10612 (N_10612,N_10377,N_10326);
nor U10613 (N_10613,N_10393,N_10111);
nand U10614 (N_10614,N_10280,N_10355);
xnor U10615 (N_10615,N_10242,N_10197);
or U10616 (N_10616,N_10228,N_10279);
and U10617 (N_10617,N_10003,N_10304);
or U10618 (N_10618,N_10153,N_10132);
xor U10619 (N_10619,N_10253,N_10190);
and U10620 (N_10620,N_10251,N_10329);
or U10621 (N_10621,N_10357,N_10116);
nor U10622 (N_10622,N_10144,N_10223);
nand U10623 (N_10623,N_10082,N_10112);
xor U10624 (N_10624,N_10338,N_10176);
nand U10625 (N_10625,N_10033,N_10382);
nand U10626 (N_10626,N_10184,N_10230);
nor U10627 (N_10627,N_10203,N_10386);
and U10628 (N_10628,N_10224,N_10092);
and U10629 (N_10629,N_10071,N_10333);
and U10630 (N_10630,N_10071,N_10056);
xor U10631 (N_10631,N_10096,N_10142);
or U10632 (N_10632,N_10261,N_10353);
xor U10633 (N_10633,N_10396,N_10370);
nor U10634 (N_10634,N_10295,N_10175);
nor U10635 (N_10635,N_10308,N_10114);
nor U10636 (N_10636,N_10231,N_10146);
nand U10637 (N_10637,N_10276,N_10348);
and U10638 (N_10638,N_10364,N_10227);
or U10639 (N_10639,N_10139,N_10226);
nor U10640 (N_10640,N_10262,N_10289);
and U10641 (N_10641,N_10269,N_10367);
xor U10642 (N_10642,N_10003,N_10379);
and U10643 (N_10643,N_10198,N_10237);
nand U10644 (N_10644,N_10043,N_10308);
xnor U10645 (N_10645,N_10267,N_10285);
xor U10646 (N_10646,N_10248,N_10313);
and U10647 (N_10647,N_10141,N_10385);
xnor U10648 (N_10648,N_10280,N_10188);
xor U10649 (N_10649,N_10287,N_10141);
nor U10650 (N_10650,N_10132,N_10385);
and U10651 (N_10651,N_10089,N_10056);
and U10652 (N_10652,N_10089,N_10369);
xor U10653 (N_10653,N_10003,N_10165);
and U10654 (N_10654,N_10089,N_10156);
xor U10655 (N_10655,N_10013,N_10252);
xnor U10656 (N_10656,N_10200,N_10122);
nor U10657 (N_10657,N_10127,N_10073);
and U10658 (N_10658,N_10041,N_10127);
nand U10659 (N_10659,N_10365,N_10023);
nand U10660 (N_10660,N_10240,N_10040);
or U10661 (N_10661,N_10084,N_10133);
nor U10662 (N_10662,N_10168,N_10217);
nand U10663 (N_10663,N_10065,N_10241);
xor U10664 (N_10664,N_10144,N_10184);
xnor U10665 (N_10665,N_10111,N_10116);
or U10666 (N_10666,N_10034,N_10251);
xnor U10667 (N_10667,N_10010,N_10370);
xor U10668 (N_10668,N_10148,N_10216);
xor U10669 (N_10669,N_10326,N_10299);
or U10670 (N_10670,N_10141,N_10064);
xor U10671 (N_10671,N_10084,N_10016);
nand U10672 (N_10672,N_10301,N_10099);
xnor U10673 (N_10673,N_10103,N_10199);
nand U10674 (N_10674,N_10083,N_10299);
nand U10675 (N_10675,N_10071,N_10057);
or U10676 (N_10676,N_10103,N_10286);
and U10677 (N_10677,N_10087,N_10082);
nand U10678 (N_10678,N_10390,N_10332);
xnor U10679 (N_10679,N_10164,N_10050);
xnor U10680 (N_10680,N_10251,N_10053);
xnor U10681 (N_10681,N_10063,N_10299);
nand U10682 (N_10682,N_10122,N_10141);
or U10683 (N_10683,N_10130,N_10064);
or U10684 (N_10684,N_10338,N_10145);
xor U10685 (N_10685,N_10196,N_10027);
xnor U10686 (N_10686,N_10148,N_10256);
nand U10687 (N_10687,N_10004,N_10113);
xor U10688 (N_10688,N_10052,N_10147);
nor U10689 (N_10689,N_10224,N_10394);
nor U10690 (N_10690,N_10164,N_10373);
xor U10691 (N_10691,N_10236,N_10111);
or U10692 (N_10692,N_10070,N_10379);
or U10693 (N_10693,N_10296,N_10274);
xor U10694 (N_10694,N_10002,N_10302);
xnor U10695 (N_10695,N_10243,N_10382);
xnor U10696 (N_10696,N_10194,N_10095);
and U10697 (N_10697,N_10321,N_10173);
nand U10698 (N_10698,N_10249,N_10395);
and U10699 (N_10699,N_10127,N_10337);
nor U10700 (N_10700,N_10249,N_10274);
or U10701 (N_10701,N_10192,N_10026);
nand U10702 (N_10702,N_10087,N_10013);
nor U10703 (N_10703,N_10273,N_10235);
and U10704 (N_10704,N_10177,N_10200);
nor U10705 (N_10705,N_10037,N_10157);
or U10706 (N_10706,N_10360,N_10293);
nor U10707 (N_10707,N_10236,N_10102);
xor U10708 (N_10708,N_10344,N_10043);
or U10709 (N_10709,N_10004,N_10382);
and U10710 (N_10710,N_10190,N_10181);
and U10711 (N_10711,N_10340,N_10363);
nor U10712 (N_10712,N_10153,N_10040);
nor U10713 (N_10713,N_10075,N_10303);
xor U10714 (N_10714,N_10232,N_10174);
nor U10715 (N_10715,N_10295,N_10218);
nand U10716 (N_10716,N_10065,N_10293);
or U10717 (N_10717,N_10281,N_10169);
and U10718 (N_10718,N_10232,N_10085);
xnor U10719 (N_10719,N_10304,N_10390);
and U10720 (N_10720,N_10395,N_10362);
nand U10721 (N_10721,N_10291,N_10263);
and U10722 (N_10722,N_10072,N_10057);
and U10723 (N_10723,N_10138,N_10320);
xnor U10724 (N_10724,N_10127,N_10263);
nor U10725 (N_10725,N_10203,N_10249);
nand U10726 (N_10726,N_10109,N_10285);
nor U10727 (N_10727,N_10263,N_10174);
xnor U10728 (N_10728,N_10157,N_10227);
xnor U10729 (N_10729,N_10149,N_10276);
and U10730 (N_10730,N_10143,N_10253);
nand U10731 (N_10731,N_10195,N_10004);
nand U10732 (N_10732,N_10349,N_10279);
and U10733 (N_10733,N_10029,N_10156);
and U10734 (N_10734,N_10293,N_10055);
nand U10735 (N_10735,N_10326,N_10269);
xnor U10736 (N_10736,N_10389,N_10211);
or U10737 (N_10737,N_10332,N_10383);
nor U10738 (N_10738,N_10377,N_10322);
xor U10739 (N_10739,N_10103,N_10139);
nand U10740 (N_10740,N_10081,N_10169);
or U10741 (N_10741,N_10091,N_10227);
and U10742 (N_10742,N_10229,N_10154);
or U10743 (N_10743,N_10167,N_10025);
and U10744 (N_10744,N_10251,N_10385);
nor U10745 (N_10745,N_10273,N_10213);
nor U10746 (N_10746,N_10079,N_10383);
and U10747 (N_10747,N_10321,N_10297);
nand U10748 (N_10748,N_10249,N_10129);
nor U10749 (N_10749,N_10306,N_10303);
nand U10750 (N_10750,N_10069,N_10257);
nor U10751 (N_10751,N_10190,N_10386);
nand U10752 (N_10752,N_10093,N_10080);
xor U10753 (N_10753,N_10392,N_10202);
nor U10754 (N_10754,N_10290,N_10337);
nor U10755 (N_10755,N_10121,N_10147);
nand U10756 (N_10756,N_10029,N_10196);
and U10757 (N_10757,N_10270,N_10309);
xor U10758 (N_10758,N_10112,N_10231);
or U10759 (N_10759,N_10378,N_10112);
nand U10760 (N_10760,N_10076,N_10150);
nor U10761 (N_10761,N_10362,N_10104);
nor U10762 (N_10762,N_10360,N_10180);
nand U10763 (N_10763,N_10330,N_10201);
xnor U10764 (N_10764,N_10033,N_10397);
nor U10765 (N_10765,N_10032,N_10087);
xnor U10766 (N_10766,N_10027,N_10262);
or U10767 (N_10767,N_10285,N_10209);
xnor U10768 (N_10768,N_10032,N_10149);
or U10769 (N_10769,N_10102,N_10254);
nor U10770 (N_10770,N_10270,N_10140);
xnor U10771 (N_10771,N_10170,N_10173);
and U10772 (N_10772,N_10262,N_10183);
nor U10773 (N_10773,N_10343,N_10099);
or U10774 (N_10774,N_10340,N_10063);
xor U10775 (N_10775,N_10206,N_10281);
and U10776 (N_10776,N_10029,N_10111);
nand U10777 (N_10777,N_10201,N_10179);
and U10778 (N_10778,N_10142,N_10034);
nand U10779 (N_10779,N_10127,N_10360);
nor U10780 (N_10780,N_10112,N_10312);
nor U10781 (N_10781,N_10231,N_10085);
or U10782 (N_10782,N_10018,N_10212);
nor U10783 (N_10783,N_10137,N_10204);
xor U10784 (N_10784,N_10076,N_10007);
nor U10785 (N_10785,N_10082,N_10211);
or U10786 (N_10786,N_10054,N_10042);
or U10787 (N_10787,N_10134,N_10149);
nand U10788 (N_10788,N_10070,N_10081);
nand U10789 (N_10789,N_10164,N_10313);
and U10790 (N_10790,N_10365,N_10100);
or U10791 (N_10791,N_10153,N_10388);
nand U10792 (N_10792,N_10327,N_10290);
nand U10793 (N_10793,N_10325,N_10300);
and U10794 (N_10794,N_10098,N_10075);
xor U10795 (N_10795,N_10248,N_10354);
and U10796 (N_10796,N_10346,N_10041);
xor U10797 (N_10797,N_10359,N_10084);
or U10798 (N_10798,N_10174,N_10344);
nand U10799 (N_10799,N_10389,N_10150);
nor U10800 (N_10800,N_10530,N_10403);
or U10801 (N_10801,N_10686,N_10755);
nor U10802 (N_10802,N_10516,N_10771);
nor U10803 (N_10803,N_10684,N_10749);
and U10804 (N_10804,N_10654,N_10578);
nand U10805 (N_10805,N_10583,N_10780);
xor U10806 (N_10806,N_10490,N_10413);
nor U10807 (N_10807,N_10541,N_10676);
nor U10808 (N_10808,N_10742,N_10434);
nand U10809 (N_10809,N_10406,N_10540);
and U10810 (N_10810,N_10694,N_10493);
nand U10811 (N_10811,N_10552,N_10639);
and U10812 (N_10812,N_10501,N_10419);
xnor U10813 (N_10813,N_10785,N_10566);
nor U10814 (N_10814,N_10622,N_10751);
or U10815 (N_10815,N_10740,N_10645);
and U10816 (N_10816,N_10758,N_10586);
nand U10817 (N_10817,N_10709,N_10573);
xnor U10818 (N_10818,N_10750,N_10519);
nor U10819 (N_10819,N_10648,N_10559);
or U10820 (N_10820,N_10675,N_10706);
and U10821 (N_10821,N_10420,N_10596);
nand U10822 (N_10822,N_10599,N_10729);
nor U10823 (N_10823,N_10439,N_10617);
nand U10824 (N_10824,N_10746,N_10428);
or U10825 (N_10825,N_10691,N_10455);
nor U10826 (N_10826,N_10470,N_10415);
nand U10827 (N_10827,N_10792,N_10688);
and U10828 (N_10828,N_10651,N_10492);
nand U10829 (N_10829,N_10575,N_10494);
xnor U10830 (N_10830,N_10579,N_10795);
nor U10831 (N_10831,N_10695,N_10507);
or U10832 (N_10832,N_10734,N_10679);
or U10833 (N_10833,N_10550,N_10497);
or U10834 (N_10834,N_10644,N_10765);
and U10835 (N_10835,N_10607,N_10449);
or U10836 (N_10836,N_10621,N_10754);
and U10837 (N_10837,N_10782,N_10433);
and U10838 (N_10838,N_10739,N_10557);
xnor U10839 (N_10839,N_10593,N_10549);
nand U10840 (N_10840,N_10441,N_10712);
or U10841 (N_10841,N_10636,N_10738);
or U10842 (N_10842,N_10603,N_10756);
nor U10843 (N_10843,N_10558,N_10569);
and U10844 (N_10844,N_10757,N_10421);
nor U10845 (N_10845,N_10789,N_10635);
nor U10846 (N_10846,N_10656,N_10685);
or U10847 (N_10847,N_10791,N_10658);
and U10848 (N_10848,N_10741,N_10626);
nor U10849 (N_10849,N_10776,N_10580);
nor U10850 (N_10850,N_10669,N_10662);
nor U10851 (N_10851,N_10605,N_10521);
nor U10852 (N_10852,N_10660,N_10401);
nand U10853 (N_10853,N_10400,N_10611);
xnor U10854 (N_10854,N_10546,N_10799);
and U10855 (N_10855,N_10444,N_10663);
nor U10856 (N_10856,N_10479,N_10736);
or U10857 (N_10857,N_10601,N_10481);
nand U10858 (N_10858,N_10752,N_10404);
and U10859 (N_10859,N_10504,N_10784);
nand U10860 (N_10860,N_10667,N_10445);
nand U10861 (N_10861,N_10589,N_10430);
nor U10862 (N_10862,N_10683,N_10721);
or U10863 (N_10863,N_10598,N_10618);
xor U10864 (N_10864,N_10506,N_10567);
and U10865 (N_10865,N_10597,N_10769);
and U10866 (N_10866,N_10787,N_10630);
nor U10867 (N_10867,N_10475,N_10527);
and U10868 (N_10868,N_10582,N_10454);
xnor U10869 (N_10869,N_10747,N_10581);
xor U10870 (N_10870,N_10446,N_10513);
nor U10871 (N_10871,N_10543,N_10783);
xnor U10872 (N_10872,N_10466,N_10606);
and U10873 (N_10873,N_10531,N_10779);
and U10874 (N_10874,N_10687,N_10767);
or U10875 (N_10875,N_10710,N_10609);
nor U10876 (N_10876,N_10517,N_10778);
nand U10877 (N_10877,N_10637,N_10487);
nor U10878 (N_10878,N_10650,N_10604);
nand U10879 (N_10879,N_10777,N_10483);
and U10880 (N_10880,N_10774,N_10463);
xor U10881 (N_10881,N_10499,N_10722);
nor U10882 (N_10882,N_10514,N_10797);
or U10883 (N_10883,N_10717,N_10563);
nor U10884 (N_10884,N_10476,N_10733);
nor U10885 (N_10885,N_10763,N_10544);
nand U10886 (N_10886,N_10759,N_10697);
and U10887 (N_10887,N_10732,N_10555);
xor U10888 (N_10888,N_10459,N_10786);
nand U10889 (N_10889,N_10461,N_10526);
xor U10890 (N_10890,N_10737,N_10659);
xnor U10891 (N_10891,N_10704,N_10608);
nor U10892 (N_10892,N_10690,N_10432);
or U10893 (N_10893,N_10408,N_10595);
nand U10894 (N_10894,N_10615,N_10653);
nand U10895 (N_10895,N_10716,N_10447);
nor U10896 (N_10896,N_10701,N_10594);
nor U10897 (N_10897,N_10692,N_10437);
nand U10898 (N_10898,N_10587,N_10562);
nand U10899 (N_10899,N_10511,N_10713);
or U10900 (N_10900,N_10484,N_10533);
nand U10901 (N_10901,N_10711,N_10515);
or U10902 (N_10902,N_10631,N_10418);
nand U10903 (N_10903,N_10423,N_10471);
nand U10904 (N_10904,N_10643,N_10467);
xnor U10905 (N_10905,N_10551,N_10409);
xnor U10906 (N_10906,N_10477,N_10681);
nand U10907 (N_10907,N_10538,N_10560);
xnor U10908 (N_10908,N_10762,N_10529);
xor U10909 (N_10909,N_10480,N_10632);
and U10910 (N_10910,N_10495,N_10796);
and U10911 (N_10911,N_10612,N_10468);
nand U10912 (N_10912,N_10705,N_10748);
xor U10913 (N_10913,N_10781,N_10646);
xnor U10914 (N_10914,N_10440,N_10642);
xnor U10915 (N_10915,N_10728,N_10661);
nand U10916 (N_10916,N_10590,N_10509);
nor U10917 (N_10917,N_10491,N_10700);
nor U10918 (N_10918,N_10414,N_10613);
and U10919 (N_10919,N_10458,N_10510);
and U10920 (N_10920,N_10496,N_10435);
and U10921 (N_10921,N_10405,N_10652);
xnor U10922 (N_10922,N_10469,N_10693);
and U10923 (N_10923,N_10453,N_10528);
xnor U10924 (N_10924,N_10680,N_10638);
and U10925 (N_10925,N_10610,N_10503);
and U10926 (N_10926,N_10462,N_10518);
xor U10927 (N_10927,N_10649,N_10625);
or U10928 (N_10928,N_10720,N_10422);
or U10929 (N_10929,N_10678,N_10426);
or U10930 (N_10930,N_10772,N_10773);
nor U10931 (N_10931,N_10554,N_10523);
nand U10932 (N_10932,N_10502,N_10410);
nand U10933 (N_10933,N_10666,N_10794);
nand U10934 (N_10934,N_10505,N_10485);
nand U10935 (N_10935,N_10629,N_10412);
xor U10936 (N_10936,N_10760,N_10539);
nor U10937 (N_10937,N_10627,N_10745);
xor U10938 (N_10938,N_10744,N_10585);
xnor U10939 (N_10939,N_10714,N_10620);
xnor U10940 (N_10940,N_10535,N_10464);
or U10941 (N_10941,N_10465,N_10548);
and U10942 (N_10942,N_10565,N_10614);
nand U10943 (N_10943,N_10570,N_10634);
nand U10944 (N_10944,N_10640,N_10724);
xor U10945 (N_10945,N_10766,N_10790);
nand U10946 (N_10946,N_10624,N_10670);
nand U10947 (N_10947,N_10473,N_10671);
xnor U10948 (N_10948,N_10715,N_10698);
nand U10949 (N_10949,N_10668,N_10703);
xor U10950 (N_10950,N_10488,N_10577);
nor U10951 (N_10951,N_10619,N_10677);
nand U10952 (N_10952,N_10768,N_10508);
nor U10953 (N_10953,N_10574,N_10628);
xor U10954 (N_10954,N_10478,N_10672);
nand U10955 (N_10955,N_10568,N_10664);
nor U10956 (N_10956,N_10775,N_10584);
nor U10957 (N_10957,N_10682,N_10556);
and U10958 (N_10958,N_10743,N_10592);
and U10959 (N_10959,N_10793,N_10512);
xnor U10960 (N_10960,N_10719,N_10770);
and U10961 (N_10961,N_10647,N_10731);
nor U10962 (N_10962,N_10457,N_10498);
and U10963 (N_10963,N_10436,N_10602);
xnor U10964 (N_10964,N_10798,N_10616);
nor U10965 (N_10965,N_10633,N_10673);
nand U10966 (N_10966,N_10536,N_10431);
and U10967 (N_10967,N_10486,N_10542);
nor U10968 (N_10968,N_10520,N_10708);
or U10969 (N_10969,N_10761,N_10451);
or U10970 (N_10970,N_10411,N_10730);
nor U10971 (N_10971,N_10623,N_10525);
and U10972 (N_10972,N_10726,N_10532);
or U10973 (N_10973,N_10452,N_10689);
or U10974 (N_10974,N_10553,N_10753);
xor U10975 (N_10975,N_10460,N_10788);
nor U10976 (N_10976,N_10545,N_10657);
nor U10977 (N_10977,N_10424,N_10564);
nand U10978 (N_10978,N_10735,N_10425);
or U10979 (N_10979,N_10764,N_10699);
nor U10980 (N_10980,N_10522,N_10534);
and U10981 (N_10981,N_10727,N_10438);
or U10982 (N_10982,N_10427,N_10500);
or U10983 (N_10983,N_10407,N_10600);
nor U10984 (N_10984,N_10416,N_10588);
xnor U10985 (N_10985,N_10696,N_10472);
xnor U10986 (N_10986,N_10707,N_10723);
nand U10987 (N_10987,N_10641,N_10655);
and U10988 (N_10988,N_10450,N_10547);
xor U10989 (N_10989,N_10474,N_10537);
or U10990 (N_10990,N_10571,N_10576);
nor U10991 (N_10991,N_10482,N_10665);
and U10992 (N_10992,N_10702,N_10448);
or U10993 (N_10993,N_10725,N_10489);
and U10994 (N_10994,N_10718,N_10456);
nor U10995 (N_10995,N_10443,N_10572);
and U10996 (N_10996,N_10417,N_10429);
xnor U10997 (N_10997,N_10402,N_10561);
nand U10998 (N_10998,N_10524,N_10591);
xor U10999 (N_10999,N_10674,N_10442);
or U11000 (N_11000,N_10730,N_10557);
or U11001 (N_11001,N_10542,N_10402);
xor U11002 (N_11002,N_10476,N_10603);
nor U11003 (N_11003,N_10756,N_10612);
and U11004 (N_11004,N_10632,N_10457);
or U11005 (N_11005,N_10483,N_10669);
and U11006 (N_11006,N_10716,N_10560);
and U11007 (N_11007,N_10615,N_10575);
or U11008 (N_11008,N_10770,N_10607);
xor U11009 (N_11009,N_10681,N_10713);
nor U11010 (N_11010,N_10442,N_10692);
and U11011 (N_11011,N_10732,N_10620);
and U11012 (N_11012,N_10776,N_10692);
and U11013 (N_11013,N_10455,N_10754);
xor U11014 (N_11014,N_10554,N_10786);
and U11015 (N_11015,N_10776,N_10731);
and U11016 (N_11016,N_10424,N_10701);
or U11017 (N_11017,N_10574,N_10411);
or U11018 (N_11018,N_10541,N_10559);
nand U11019 (N_11019,N_10740,N_10793);
nor U11020 (N_11020,N_10456,N_10469);
or U11021 (N_11021,N_10464,N_10551);
and U11022 (N_11022,N_10561,N_10668);
or U11023 (N_11023,N_10779,N_10694);
or U11024 (N_11024,N_10697,N_10724);
nor U11025 (N_11025,N_10651,N_10678);
nand U11026 (N_11026,N_10471,N_10634);
xnor U11027 (N_11027,N_10537,N_10512);
and U11028 (N_11028,N_10413,N_10654);
nand U11029 (N_11029,N_10447,N_10645);
xnor U11030 (N_11030,N_10542,N_10458);
or U11031 (N_11031,N_10791,N_10476);
or U11032 (N_11032,N_10555,N_10479);
xnor U11033 (N_11033,N_10402,N_10481);
xnor U11034 (N_11034,N_10529,N_10629);
or U11035 (N_11035,N_10557,N_10795);
or U11036 (N_11036,N_10716,N_10698);
nand U11037 (N_11037,N_10672,N_10565);
and U11038 (N_11038,N_10538,N_10412);
xor U11039 (N_11039,N_10479,N_10773);
nand U11040 (N_11040,N_10779,N_10614);
nand U11041 (N_11041,N_10448,N_10507);
and U11042 (N_11042,N_10688,N_10672);
and U11043 (N_11043,N_10490,N_10469);
nand U11044 (N_11044,N_10569,N_10753);
xor U11045 (N_11045,N_10730,N_10570);
or U11046 (N_11046,N_10520,N_10789);
or U11047 (N_11047,N_10490,N_10517);
and U11048 (N_11048,N_10779,N_10778);
or U11049 (N_11049,N_10791,N_10768);
and U11050 (N_11050,N_10407,N_10500);
or U11051 (N_11051,N_10509,N_10750);
nor U11052 (N_11052,N_10455,N_10782);
nor U11053 (N_11053,N_10472,N_10566);
nor U11054 (N_11054,N_10677,N_10725);
or U11055 (N_11055,N_10609,N_10452);
nand U11056 (N_11056,N_10543,N_10682);
nand U11057 (N_11057,N_10753,N_10730);
nand U11058 (N_11058,N_10439,N_10480);
nand U11059 (N_11059,N_10630,N_10480);
nor U11060 (N_11060,N_10577,N_10464);
nor U11061 (N_11061,N_10551,N_10615);
nor U11062 (N_11062,N_10569,N_10625);
xor U11063 (N_11063,N_10629,N_10626);
nand U11064 (N_11064,N_10651,N_10623);
or U11065 (N_11065,N_10543,N_10725);
nor U11066 (N_11066,N_10541,N_10693);
xnor U11067 (N_11067,N_10722,N_10582);
nand U11068 (N_11068,N_10553,N_10489);
and U11069 (N_11069,N_10608,N_10410);
nor U11070 (N_11070,N_10512,N_10626);
nor U11071 (N_11071,N_10591,N_10716);
nor U11072 (N_11072,N_10717,N_10686);
xnor U11073 (N_11073,N_10777,N_10789);
or U11074 (N_11074,N_10408,N_10565);
xor U11075 (N_11075,N_10434,N_10510);
and U11076 (N_11076,N_10665,N_10731);
nor U11077 (N_11077,N_10736,N_10585);
and U11078 (N_11078,N_10643,N_10613);
nand U11079 (N_11079,N_10500,N_10620);
and U11080 (N_11080,N_10606,N_10654);
xor U11081 (N_11081,N_10721,N_10626);
nand U11082 (N_11082,N_10608,N_10742);
and U11083 (N_11083,N_10692,N_10581);
and U11084 (N_11084,N_10523,N_10689);
and U11085 (N_11085,N_10607,N_10645);
nand U11086 (N_11086,N_10443,N_10665);
nand U11087 (N_11087,N_10457,N_10563);
xnor U11088 (N_11088,N_10502,N_10707);
or U11089 (N_11089,N_10766,N_10557);
and U11090 (N_11090,N_10549,N_10567);
or U11091 (N_11091,N_10478,N_10557);
or U11092 (N_11092,N_10579,N_10613);
or U11093 (N_11093,N_10456,N_10437);
or U11094 (N_11094,N_10433,N_10783);
xor U11095 (N_11095,N_10600,N_10408);
nor U11096 (N_11096,N_10595,N_10651);
nor U11097 (N_11097,N_10672,N_10475);
xnor U11098 (N_11098,N_10677,N_10457);
xnor U11099 (N_11099,N_10496,N_10603);
nor U11100 (N_11100,N_10542,N_10578);
and U11101 (N_11101,N_10742,N_10761);
and U11102 (N_11102,N_10765,N_10491);
or U11103 (N_11103,N_10400,N_10696);
nand U11104 (N_11104,N_10455,N_10612);
xnor U11105 (N_11105,N_10786,N_10667);
nand U11106 (N_11106,N_10650,N_10660);
nor U11107 (N_11107,N_10488,N_10570);
xnor U11108 (N_11108,N_10434,N_10450);
and U11109 (N_11109,N_10581,N_10525);
and U11110 (N_11110,N_10795,N_10479);
xnor U11111 (N_11111,N_10410,N_10518);
or U11112 (N_11112,N_10553,N_10458);
nand U11113 (N_11113,N_10454,N_10779);
xnor U11114 (N_11114,N_10790,N_10425);
or U11115 (N_11115,N_10795,N_10566);
or U11116 (N_11116,N_10458,N_10476);
and U11117 (N_11117,N_10700,N_10652);
or U11118 (N_11118,N_10436,N_10567);
nor U11119 (N_11119,N_10402,N_10744);
and U11120 (N_11120,N_10683,N_10606);
xor U11121 (N_11121,N_10503,N_10744);
nor U11122 (N_11122,N_10741,N_10716);
nor U11123 (N_11123,N_10604,N_10408);
and U11124 (N_11124,N_10716,N_10616);
or U11125 (N_11125,N_10458,N_10726);
or U11126 (N_11126,N_10503,N_10690);
xnor U11127 (N_11127,N_10572,N_10552);
nand U11128 (N_11128,N_10585,N_10590);
xnor U11129 (N_11129,N_10793,N_10714);
nand U11130 (N_11130,N_10508,N_10558);
nand U11131 (N_11131,N_10688,N_10429);
nand U11132 (N_11132,N_10740,N_10613);
nor U11133 (N_11133,N_10569,N_10643);
xor U11134 (N_11134,N_10678,N_10793);
nand U11135 (N_11135,N_10687,N_10556);
nand U11136 (N_11136,N_10490,N_10793);
nor U11137 (N_11137,N_10525,N_10422);
or U11138 (N_11138,N_10464,N_10701);
and U11139 (N_11139,N_10611,N_10578);
and U11140 (N_11140,N_10451,N_10731);
nand U11141 (N_11141,N_10777,N_10517);
nand U11142 (N_11142,N_10559,N_10790);
nor U11143 (N_11143,N_10408,N_10550);
nor U11144 (N_11144,N_10556,N_10431);
nor U11145 (N_11145,N_10697,N_10725);
nand U11146 (N_11146,N_10558,N_10655);
nand U11147 (N_11147,N_10604,N_10438);
xor U11148 (N_11148,N_10737,N_10446);
or U11149 (N_11149,N_10520,N_10436);
and U11150 (N_11150,N_10787,N_10432);
nor U11151 (N_11151,N_10733,N_10575);
and U11152 (N_11152,N_10667,N_10405);
nand U11153 (N_11153,N_10433,N_10718);
or U11154 (N_11154,N_10763,N_10743);
or U11155 (N_11155,N_10667,N_10640);
xnor U11156 (N_11156,N_10781,N_10619);
nor U11157 (N_11157,N_10685,N_10448);
or U11158 (N_11158,N_10528,N_10766);
xor U11159 (N_11159,N_10633,N_10571);
and U11160 (N_11160,N_10662,N_10729);
nor U11161 (N_11161,N_10784,N_10623);
and U11162 (N_11162,N_10524,N_10459);
or U11163 (N_11163,N_10685,N_10695);
nand U11164 (N_11164,N_10717,N_10627);
nor U11165 (N_11165,N_10742,N_10479);
and U11166 (N_11166,N_10587,N_10712);
or U11167 (N_11167,N_10575,N_10764);
xnor U11168 (N_11168,N_10509,N_10715);
xnor U11169 (N_11169,N_10797,N_10593);
nand U11170 (N_11170,N_10469,N_10781);
or U11171 (N_11171,N_10467,N_10656);
xor U11172 (N_11172,N_10587,N_10711);
xor U11173 (N_11173,N_10472,N_10482);
nand U11174 (N_11174,N_10625,N_10709);
or U11175 (N_11175,N_10577,N_10555);
or U11176 (N_11176,N_10410,N_10789);
and U11177 (N_11177,N_10731,N_10703);
xor U11178 (N_11178,N_10479,N_10551);
xnor U11179 (N_11179,N_10575,N_10753);
or U11180 (N_11180,N_10527,N_10638);
nand U11181 (N_11181,N_10589,N_10422);
nand U11182 (N_11182,N_10632,N_10464);
or U11183 (N_11183,N_10643,N_10671);
xor U11184 (N_11184,N_10674,N_10454);
nand U11185 (N_11185,N_10733,N_10405);
nand U11186 (N_11186,N_10468,N_10674);
nand U11187 (N_11187,N_10553,N_10554);
xor U11188 (N_11188,N_10606,N_10646);
nor U11189 (N_11189,N_10677,N_10451);
and U11190 (N_11190,N_10456,N_10790);
xor U11191 (N_11191,N_10561,N_10522);
nor U11192 (N_11192,N_10741,N_10737);
and U11193 (N_11193,N_10453,N_10564);
nor U11194 (N_11194,N_10556,N_10442);
nand U11195 (N_11195,N_10445,N_10696);
and U11196 (N_11196,N_10505,N_10439);
or U11197 (N_11197,N_10466,N_10541);
nand U11198 (N_11198,N_10549,N_10471);
or U11199 (N_11199,N_10400,N_10541);
or U11200 (N_11200,N_10837,N_10985);
nor U11201 (N_11201,N_10884,N_10857);
or U11202 (N_11202,N_10965,N_11067);
and U11203 (N_11203,N_10982,N_11167);
nand U11204 (N_11204,N_11106,N_11081);
nor U11205 (N_11205,N_10858,N_11163);
and U11206 (N_11206,N_11033,N_10961);
nor U11207 (N_11207,N_10991,N_10841);
or U11208 (N_11208,N_11117,N_11122);
or U11209 (N_11209,N_11056,N_11003);
or U11210 (N_11210,N_11107,N_11159);
nand U11211 (N_11211,N_11176,N_10959);
or U11212 (N_11212,N_10828,N_10878);
or U11213 (N_11213,N_11145,N_11057);
or U11214 (N_11214,N_11080,N_11127);
and U11215 (N_11215,N_11153,N_10865);
nor U11216 (N_11216,N_11155,N_10815);
and U11217 (N_11217,N_11087,N_11051);
nand U11218 (N_11218,N_10939,N_10847);
nor U11219 (N_11219,N_10926,N_11169);
and U11220 (N_11220,N_11017,N_10854);
and U11221 (N_11221,N_11074,N_10936);
nor U11222 (N_11222,N_10973,N_10941);
and U11223 (N_11223,N_11068,N_10819);
or U11224 (N_11224,N_11054,N_11035);
and U11225 (N_11225,N_11177,N_11013);
xnor U11226 (N_11226,N_11042,N_10824);
nor U11227 (N_11227,N_10832,N_10812);
or U11228 (N_11228,N_10954,N_11034);
and U11229 (N_11229,N_10881,N_11114);
nor U11230 (N_11230,N_10803,N_11036);
or U11231 (N_11231,N_10953,N_10901);
nor U11232 (N_11232,N_11046,N_10975);
and U11233 (N_11233,N_11148,N_11133);
xnor U11234 (N_11234,N_10964,N_11020);
and U11235 (N_11235,N_10810,N_10919);
nand U11236 (N_11236,N_11016,N_11093);
nand U11237 (N_11237,N_11089,N_11031);
nand U11238 (N_11238,N_10915,N_10940);
nand U11239 (N_11239,N_10852,N_10823);
nor U11240 (N_11240,N_10826,N_11053);
nand U11241 (N_11241,N_10846,N_11158);
nor U11242 (N_11242,N_10821,N_11124);
and U11243 (N_11243,N_10989,N_11041);
or U11244 (N_11244,N_11043,N_10978);
xor U11245 (N_11245,N_10877,N_10909);
nand U11246 (N_11246,N_11160,N_10920);
or U11247 (N_11247,N_11129,N_11109);
xor U11248 (N_11248,N_11065,N_11029);
xor U11249 (N_11249,N_10995,N_11125);
and U11250 (N_11250,N_11086,N_10814);
or U11251 (N_11251,N_11126,N_10931);
nor U11252 (N_11252,N_10840,N_10938);
nor U11253 (N_11253,N_10908,N_10893);
nor U11254 (N_11254,N_10952,N_10983);
nand U11255 (N_11255,N_11078,N_10808);
nand U11256 (N_11256,N_10862,N_11099);
nand U11257 (N_11257,N_10816,N_10971);
and U11258 (N_11258,N_11181,N_11165);
or U11259 (N_11259,N_10904,N_10876);
nand U11260 (N_11260,N_11130,N_11192);
and U11261 (N_11261,N_10911,N_11026);
nor U11262 (N_11262,N_11194,N_11154);
nand U11263 (N_11263,N_11037,N_10831);
nand U11264 (N_11264,N_10935,N_10805);
nand U11265 (N_11265,N_11195,N_10871);
or U11266 (N_11266,N_10958,N_10890);
and U11267 (N_11267,N_11073,N_11149);
nor U11268 (N_11268,N_10905,N_10998);
nor U11269 (N_11269,N_11140,N_10800);
xor U11270 (N_11270,N_10801,N_10850);
xor U11271 (N_11271,N_11151,N_10848);
nor U11272 (N_11272,N_10955,N_11115);
or U11273 (N_11273,N_11123,N_10844);
nor U11274 (N_11274,N_10833,N_10923);
xor U11275 (N_11275,N_11139,N_10963);
and U11276 (N_11276,N_10868,N_11076);
xor U11277 (N_11277,N_11146,N_10818);
or U11278 (N_11278,N_11103,N_10887);
xnor U11279 (N_11279,N_11193,N_11105);
nand U11280 (N_11280,N_10933,N_11072);
nor U11281 (N_11281,N_10980,N_10987);
or U11282 (N_11282,N_11100,N_11136);
or U11283 (N_11283,N_10928,N_10891);
or U11284 (N_11284,N_10875,N_10898);
or U11285 (N_11285,N_10918,N_10853);
and U11286 (N_11286,N_11083,N_10999);
or U11287 (N_11287,N_11059,N_10910);
nor U11288 (N_11288,N_10830,N_11023);
or U11289 (N_11289,N_11096,N_10834);
or U11290 (N_11290,N_11113,N_10897);
and U11291 (N_11291,N_11164,N_10925);
or U11292 (N_11292,N_10932,N_10924);
nor U11293 (N_11293,N_11022,N_11183);
nor U11294 (N_11294,N_10946,N_11061);
nand U11295 (N_11295,N_10900,N_11079);
xor U11296 (N_11296,N_10855,N_11062);
or U11297 (N_11297,N_11199,N_11075);
xnor U11298 (N_11298,N_11110,N_11173);
and U11299 (N_11299,N_11048,N_10966);
or U11300 (N_11300,N_10916,N_10951);
xnor U11301 (N_11301,N_11085,N_11161);
or U11302 (N_11302,N_11063,N_11121);
nor U11303 (N_11303,N_11050,N_11077);
nand U11304 (N_11304,N_10996,N_10930);
and U11305 (N_11305,N_11040,N_10907);
nor U11306 (N_11306,N_10820,N_11104);
and U11307 (N_11307,N_11197,N_10992);
nor U11308 (N_11308,N_10943,N_10839);
and U11309 (N_11309,N_11002,N_10825);
or U11310 (N_11310,N_10969,N_11196);
nand U11311 (N_11311,N_10949,N_11116);
nand U11312 (N_11312,N_10896,N_10867);
or U11313 (N_11313,N_11012,N_11144);
nor U11314 (N_11314,N_11018,N_10906);
or U11315 (N_11315,N_10836,N_10804);
xnor U11316 (N_11316,N_10937,N_11052);
nor U11317 (N_11317,N_11198,N_11188);
and U11318 (N_11318,N_10993,N_10988);
xnor U11319 (N_11319,N_11157,N_11191);
nor U11320 (N_11320,N_11028,N_10956);
or U11321 (N_11321,N_11070,N_11166);
and U11322 (N_11322,N_11189,N_11011);
or U11323 (N_11323,N_10986,N_11019);
xnor U11324 (N_11324,N_11128,N_11112);
or U11325 (N_11325,N_11141,N_10972);
and U11326 (N_11326,N_11094,N_10838);
nor U11327 (N_11327,N_11185,N_11135);
or U11328 (N_11328,N_10912,N_10843);
nor U11329 (N_11329,N_10914,N_11049);
and U11330 (N_11330,N_10869,N_10809);
or U11331 (N_11331,N_11171,N_11071);
and U11332 (N_11332,N_11172,N_10957);
xor U11333 (N_11333,N_10886,N_10960);
nand U11334 (N_11334,N_11152,N_10894);
and U11335 (N_11335,N_11039,N_10970);
or U11336 (N_11336,N_10817,N_11060);
and U11337 (N_11337,N_11147,N_11025);
or U11338 (N_11338,N_10913,N_10922);
xor U11339 (N_11339,N_11004,N_10849);
or U11340 (N_11340,N_11027,N_11001);
nor U11341 (N_11341,N_10866,N_11007);
and U11342 (N_11342,N_10944,N_10942);
and U11343 (N_11343,N_10827,N_10927);
xor U11344 (N_11344,N_10945,N_11184);
or U11345 (N_11345,N_11024,N_11180);
nor U11346 (N_11346,N_11182,N_11131);
and U11347 (N_11347,N_10845,N_10962);
nor U11348 (N_11348,N_11187,N_11111);
and U11349 (N_11349,N_10811,N_11101);
and U11350 (N_11350,N_11038,N_11097);
nand U11351 (N_11351,N_11179,N_10967);
xor U11352 (N_11352,N_11102,N_10921);
and U11353 (N_11353,N_10829,N_11143);
nand U11354 (N_11354,N_10822,N_11091);
xor U11355 (N_11355,N_10874,N_10813);
xor U11356 (N_11356,N_11009,N_10883);
or U11357 (N_11357,N_11134,N_10947);
nand U11358 (N_11358,N_10948,N_10864);
or U11359 (N_11359,N_11030,N_10842);
or U11360 (N_11360,N_10968,N_10990);
or U11361 (N_11361,N_10892,N_10981);
xnor U11362 (N_11362,N_10863,N_11000);
nand U11363 (N_11363,N_10835,N_10859);
nor U11364 (N_11364,N_11132,N_11015);
nand U11365 (N_11365,N_11098,N_10882);
or U11366 (N_11366,N_11137,N_10872);
nor U11367 (N_11367,N_11170,N_11014);
xnor U11368 (N_11368,N_10861,N_11108);
nor U11369 (N_11369,N_10950,N_11088);
and U11370 (N_11370,N_10851,N_11186);
xor U11371 (N_11371,N_10929,N_10902);
xor U11372 (N_11372,N_10856,N_10873);
or U11373 (N_11373,N_10934,N_11178);
nand U11374 (N_11374,N_10997,N_10880);
xnor U11375 (N_11375,N_11162,N_10885);
and U11376 (N_11376,N_11092,N_10979);
and U11377 (N_11377,N_10860,N_11156);
or U11378 (N_11378,N_11190,N_11095);
xor U11379 (N_11379,N_10976,N_11010);
nor U11380 (N_11380,N_10807,N_11069);
nor U11381 (N_11381,N_11066,N_11175);
xor U11382 (N_11382,N_11142,N_11090);
and U11383 (N_11383,N_11150,N_11138);
xor U11384 (N_11384,N_11045,N_11082);
and U11385 (N_11385,N_10889,N_10899);
or U11386 (N_11386,N_11174,N_11120);
xnor U11387 (N_11387,N_11005,N_11058);
xor U11388 (N_11388,N_10994,N_11118);
nor U11389 (N_11389,N_11021,N_10895);
nor U11390 (N_11390,N_11119,N_11064);
xnor U11391 (N_11391,N_10974,N_10917);
or U11392 (N_11392,N_10806,N_11032);
or U11393 (N_11393,N_11055,N_11047);
and U11394 (N_11394,N_11168,N_11044);
xnor U11395 (N_11395,N_10977,N_11008);
nand U11396 (N_11396,N_10870,N_10802);
xor U11397 (N_11397,N_11006,N_10984);
xnor U11398 (N_11398,N_10903,N_10888);
nand U11399 (N_11399,N_11084,N_10879);
xor U11400 (N_11400,N_11130,N_11126);
nand U11401 (N_11401,N_10980,N_11108);
or U11402 (N_11402,N_11064,N_11081);
nor U11403 (N_11403,N_10801,N_11155);
nor U11404 (N_11404,N_10886,N_10883);
or U11405 (N_11405,N_10947,N_10836);
nor U11406 (N_11406,N_10888,N_10964);
nor U11407 (N_11407,N_11157,N_10942);
and U11408 (N_11408,N_10956,N_11165);
or U11409 (N_11409,N_10989,N_11005);
nor U11410 (N_11410,N_10961,N_11031);
and U11411 (N_11411,N_10960,N_10972);
xor U11412 (N_11412,N_10827,N_11042);
xor U11413 (N_11413,N_10931,N_10838);
nand U11414 (N_11414,N_11093,N_10952);
or U11415 (N_11415,N_11057,N_11154);
or U11416 (N_11416,N_11072,N_11032);
nand U11417 (N_11417,N_11127,N_11132);
xnor U11418 (N_11418,N_10812,N_11068);
or U11419 (N_11419,N_11188,N_11011);
and U11420 (N_11420,N_11028,N_10980);
xor U11421 (N_11421,N_10941,N_11099);
and U11422 (N_11422,N_10841,N_11148);
and U11423 (N_11423,N_10969,N_11074);
nor U11424 (N_11424,N_11034,N_11040);
nor U11425 (N_11425,N_11078,N_10836);
nand U11426 (N_11426,N_10977,N_11034);
or U11427 (N_11427,N_11023,N_11008);
xnor U11428 (N_11428,N_10831,N_10921);
or U11429 (N_11429,N_11126,N_10983);
or U11430 (N_11430,N_11191,N_11113);
and U11431 (N_11431,N_11017,N_11150);
nand U11432 (N_11432,N_11000,N_11056);
xnor U11433 (N_11433,N_10827,N_11128);
or U11434 (N_11434,N_10898,N_10940);
nand U11435 (N_11435,N_10911,N_10949);
xor U11436 (N_11436,N_11129,N_11089);
xnor U11437 (N_11437,N_10806,N_11111);
nand U11438 (N_11438,N_10979,N_10821);
xnor U11439 (N_11439,N_10962,N_11099);
and U11440 (N_11440,N_10846,N_10827);
or U11441 (N_11441,N_11195,N_10808);
nand U11442 (N_11442,N_10834,N_10961);
and U11443 (N_11443,N_11125,N_10966);
xor U11444 (N_11444,N_10836,N_10876);
xor U11445 (N_11445,N_11138,N_11168);
xor U11446 (N_11446,N_10893,N_11086);
nand U11447 (N_11447,N_11099,N_10900);
xor U11448 (N_11448,N_11168,N_10826);
nand U11449 (N_11449,N_10952,N_11019);
xor U11450 (N_11450,N_11045,N_11188);
nand U11451 (N_11451,N_11076,N_10991);
nor U11452 (N_11452,N_11046,N_11009);
nor U11453 (N_11453,N_11197,N_10820);
nand U11454 (N_11454,N_11073,N_10838);
nor U11455 (N_11455,N_11161,N_11191);
nor U11456 (N_11456,N_10901,N_11127);
nor U11457 (N_11457,N_11026,N_11127);
or U11458 (N_11458,N_11105,N_10826);
nand U11459 (N_11459,N_11192,N_11165);
nand U11460 (N_11460,N_10893,N_10839);
nand U11461 (N_11461,N_10819,N_10890);
xor U11462 (N_11462,N_11103,N_10907);
or U11463 (N_11463,N_11190,N_10865);
and U11464 (N_11464,N_11079,N_11172);
nand U11465 (N_11465,N_10830,N_10925);
or U11466 (N_11466,N_10931,N_11009);
nor U11467 (N_11467,N_11003,N_11113);
nor U11468 (N_11468,N_10959,N_10956);
or U11469 (N_11469,N_10866,N_11183);
or U11470 (N_11470,N_10970,N_11176);
nand U11471 (N_11471,N_11191,N_10939);
and U11472 (N_11472,N_11113,N_10824);
or U11473 (N_11473,N_11157,N_11106);
or U11474 (N_11474,N_11007,N_11033);
nand U11475 (N_11475,N_11190,N_11129);
and U11476 (N_11476,N_11102,N_11045);
nor U11477 (N_11477,N_11054,N_11034);
or U11478 (N_11478,N_11128,N_11089);
and U11479 (N_11479,N_11161,N_11013);
nor U11480 (N_11480,N_10964,N_11130);
xor U11481 (N_11481,N_10920,N_11179);
and U11482 (N_11482,N_10979,N_11133);
nand U11483 (N_11483,N_11015,N_10937);
nand U11484 (N_11484,N_10817,N_10940);
xor U11485 (N_11485,N_11116,N_10833);
and U11486 (N_11486,N_10932,N_11059);
nor U11487 (N_11487,N_11192,N_10882);
nand U11488 (N_11488,N_10945,N_11100);
and U11489 (N_11489,N_11029,N_11127);
or U11490 (N_11490,N_11006,N_11174);
and U11491 (N_11491,N_10834,N_10872);
or U11492 (N_11492,N_11118,N_11155);
xnor U11493 (N_11493,N_11006,N_11176);
nand U11494 (N_11494,N_11107,N_11028);
and U11495 (N_11495,N_10949,N_11073);
or U11496 (N_11496,N_11141,N_10942);
nand U11497 (N_11497,N_11104,N_10800);
nor U11498 (N_11498,N_10977,N_11018);
nand U11499 (N_11499,N_10935,N_10820);
nor U11500 (N_11500,N_11057,N_10893);
and U11501 (N_11501,N_10943,N_10907);
nand U11502 (N_11502,N_10962,N_10831);
and U11503 (N_11503,N_10871,N_11147);
xnor U11504 (N_11504,N_10824,N_10855);
nand U11505 (N_11505,N_11026,N_10957);
xor U11506 (N_11506,N_10908,N_11002);
xor U11507 (N_11507,N_11175,N_11061);
or U11508 (N_11508,N_11178,N_10930);
and U11509 (N_11509,N_10989,N_11037);
and U11510 (N_11510,N_10831,N_10918);
and U11511 (N_11511,N_10981,N_10959);
nor U11512 (N_11512,N_11045,N_11120);
nand U11513 (N_11513,N_10823,N_11123);
nor U11514 (N_11514,N_10972,N_11079);
xor U11515 (N_11515,N_10881,N_11016);
nor U11516 (N_11516,N_11155,N_11022);
or U11517 (N_11517,N_10834,N_10816);
xor U11518 (N_11518,N_10815,N_11128);
nand U11519 (N_11519,N_10878,N_10868);
nor U11520 (N_11520,N_11049,N_11019);
and U11521 (N_11521,N_10957,N_10976);
or U11522 (N_11522,N_10993,N_11028);
nand U11523 (N_11523,N_10974,N_10927);
xnor U11524 (N_11524,N_10898,N_10801);
nand U11525 (N_11525,N_10869,N_10940);
nor U11526 (N_11526,N_10820,N_11003);
or U11527 (N_11527,N_11155,N_10962);
nor U11528 (N_11528,N_10833,N_10828);
xnor U11529 (N_11529,N_11057,N_11164);
nand U11530 (N_11530,N_11023,N_11152);
nor U11531 (N_11531,N_10862,N_10808);
nor U11532 (N_11532,N_11148,N_10849);
nor U11533 (N_11533,N_11011,N_11104);
and U11534 (N_11534,N_10995,N_10882);
xor U11535 (N_11535,N_11178,N_11095);
and U11536 (N_11536,N_10814,N_10980);
and U11537 (N_11537,N_10809,N_11115);
nand U11538 (N_11538,N_11034,N_10869);
and U11539 (N_11539,N_11164,N_10872);
or U11540 (N_11540,N_10807,N_11172);
nand U11541 (N_11541,N_11080,N_11032);
or U11542 (N_11542,N_11057,N_11152);
nand U11543 (N_11543,N_11128,N_11010);
or U11544 (N_11544,N_11013,N_10989);
and U11545 (N_11545,N_10805,N_10804);
nand U11546 (N_11546,N_10875,N_11002);
nand U11547 (N_11547,N_10913,N_10804);
xnor U11548 (N_11548,N_10965,N_11157);
xnor U11549 (N_11549,N_11096,N_10816);
nor U11550 (N_11550,N_11110,N_10959);
nor U11551 (N_11551,N_10977,N_11182);
or U11552 (N_11552,N_10960,N_11075);
nor U11553 (N_11553,N_10988,N_11123);
and U11554 (N_11554,N_10882,N_10833);
xnor U11555 (N_11555,N_11106,N_10873);
nor U11556 (N_11556,N_10993,N_11175);
and U11557 (N_11557,N_11120,N_10931);
nor U11558 (N_11558,N_10818,N_10941);
nor U11559 (N_11559,N_10867,N_10923);
xor U11560 (N_11560,N_11017,N_10822);
and U11561 (N_11561,N_11185,N_11016);
and U11562 (N_11562,N_10909,N_11085);
and U11563 (N_11563,N_11168,N_10888);
nand U11564 (N_11564,N_11077,N_10969);
and U11565 (N_11565,N_10857,N_10987);
nand U11566 (N_11566,N_10962,N_10975);
nor U11567 (N_11567,N_11143,N_11114);
or U11568 (N_11568,N_11078,N_11010);
xor U11569 (N_11569,N_11025,N_11156);
nand U11570 (N_11570,N_11142,N_11091);
and U11571 (N_11571,N_11079,N_11088);
nor U11572 (N_11572,N_10865,N_10816);
and U11573 (N_11573,N_11121,N_10865);
nor U11574 (N_11574,N_11148,N_11177);
xor U11575 (N_11575,N_10918,N_10934);
and U11576 (N_11576,N_11180,N_11151);
and U11577 (N_11577,N_11133,N_11092);
xnor U11578 (N_11578,N_10866,N_10951);
nand U11579 (N_11579,N_10822,N_11047);
or U11580 (N_11580,N_11181,N_11170);
and U11581 (N_11581,N_10914,N_11108);
and U11582 (N_11582,N_11017,N_11056);
nor U11583 (N_11583,N_10823,N_11112);
nor U11584 (N_11584,N_10854,N_11092);
nor U11585 (N_11585,N_10846,N_10891);
nand U11586 (N_11586,N_10836,N_11009);
or U11587 (N_11587,N_10855,N_11119);
xnor U11588 (N_11588,N_10910,N_11193);
nor U11589 (N_11589,N_10927,N_11107);
and U11590 (N_11590,N_10830,N_10988);
or U11591 (N_11591,N_11000,N_11119);
and U11592 (N_11592,N_11188,N_10884);
nand U11593 (N_11593,N_10803,N_11122);
nand U11594 (N_11594,N_11028,N_11073);
and U11595 (N_11595,N_10866,N_10860);
nand U11596 (N_11596,N_10846,N_11034);
nor U11597 (N_11597,N_10938,N_11134);
xor U11598 (N_11598,N_11026,N_11038);
nor U11599 (N_11599,N_11178,N_10863);
nand U11600 (N_11600,N_11296,N_11205);
and U11601 (N_11601,N_11569,N_11251);
and U11602 (N_11602,N_11259,N_11281);
nand U11603 (N_11603,N_11518,N_11439);
nor U11604 (N_11604,N_11466,N_11527);
or U11605 (N_11605,N_11303,N_11595);
nand U11606 (N_11606,N_11278,N_11414);
or U11607 (N_11607,N_11272,N_11548);
and U11608 (N_11608,N_11556,N_11574);
or U11609 (N_11609,N_11509,N_11394);
and U11610 (N_11610,N_11552,N_11382);
nor U11611 (N_11611,N_11521,N_11242);
nor U11612 (N_11612,N_11430,N_11557);
and U11613 (N_11613,N_11338,N_11500);
or U11614 (N_11614,N_11555,N_11495);
and U11615 (N_11615,N_11597,N_11508);
and U11616 (N_11616,N_11565,N_11250);
xnor U11617 (N_11617,N_11260,N_11219);
nor U11618 (N_11618,N_11547,N_11586);
or U11619 (N_11619,N_11315,N_11328);
nor U11620 (N_11620,N_11368,N_11332);
nand U11621 (N_11621,N_11443,N_11375);
or U11622 (N_11622,N_11519,N_11531);
xor U11623 (N_11623,N_11475,N_11481);
nand U11624 (N_11624,N_11476,N_11346);
xnor U11625 (N_11625,N_11232,N_11596);
nor U11626 (N_11626,N_11397,N_11458);
or U11627 (N_11627,N_11350,N_11451);
and U11628 (N_11628,N_11222,N_11316);
or U11629 (N_11629,N_11284,N_11321);
xnor U11630 (N_11630,N_11352,N_11313);
xor U11631 (N_11631,N_11302,N_11479);
xnor U11632 (N_11632,N_11325,N_11246);
nor U11633 (N_11633,N_11317,N_11238);
or U11634 (N_11634,N_11429,N_11487);
nor U11635 (N_11635,N_11357,N_11459);
nor U11636 (N_11636,N_11228,N_11378);
nor U11637 (N_11637,N_11270,N_11499);
and U11638 (N_11638,N_11482,N_11204);
and U11639 (N_11639,N_11422,N_11209);
xnor U11640 (N_11640,N_11478,N_11288);
or U11641 (N_11641,N_11431,N_11513);
xnor U11642 (N_11642,N_11269,N_11493);
xnor U11643 (N_11643,N_11541,N_11572);
nor U11644 (N_11644,N_11584,N_11588);
xor U11645 (N_11645,N_11523,N_11449);
nor U11646 (N_11646,N_11336,N_11593);
or U11647 (N_11647,N_11585,N_11471);
xnor U11648 (N_11648,N_11410,N_11225);
nor U11649 (N_11649,N_11477,N_11327);
nand U11650 (N_11650,N_11544,N_11575);
or U11651 (N_11651,N_11501,N_11448);
nand U11652 (N_11652,N_11267,N_11516);
xor U11653 (N_11653,N_11230,N_11582);
and U11654 (N_11654,N_11229,N_11530);
xor U11655 (N_11655,N_11420,N_11245);
nand U11656 (N_11656,N_11413,N_11559);
or U11657 (N_11657,N_11247,N_11221);
nand U11658 (N_11658,N_11533,N_11571);
nor U11659 (N_11659,N_11208,N_11224);
xnor U11660 (N_11660,N_11432,N_11291);
nand U11661 (N_11661,N_11517,N_11457);
xnor U11662 (N_11662,N_11416,N_11223);
or U11663 (N_11663,N_11570,N_11212);
nand U11664 (N_11664,N_11507,N_11384);
nor U11665 (N_11665,N_11203,N_11268);
nand U11666 (N_11666,N_11265,N_11337);
nand U11667 (N_11667,N_11253,N_11442);
and U11668 (N_11668,N_11347,N_11386);
and U11669 (N_11669,N_11436,N_11496);
or U11670 (N_11670,N_11463,N_11262);
nor U11671 (N_11671,N_11578,N_11470);
nor U11672 (N_11672,N_11445,N_11280);
xnor U11673 (N_11673,N_11399,N_11240);
and U11674 (N_11674,N_11279,N_11558);
xnor U11675 (N_11675,N_11423,N_11522);
xor U11676 (N_11676,N_11535,N_11402);
or U11677 (N_11677,N_11294,N_11322);
nor U11678 (N_11678,N_11453,N_11235);
nor U11679 (N_11679,N_11485,N_11591);
xor U11680 (N_11680,N_11371,N_11292);
nor U11681 (N_11681,N_11381,N_11231);
or U11682 (N_11682,N_11392,N_11307);
nand U11683 (N_11683,N_11455,N_11213);
nor U11684 (N_11684,N_11543,N_11217);
and U11685 (N_11685,N_11526,N_11576);
and U11686 (N_11686,N_11363,N_11456);
xnor U11687 (N_11687,N_11318,N_11335);
nand U11688 (N_11688,N_11549,N_11324);
nand U11689 (N_11689,N_11540,N_11323);
xnor U11690 (N_11690,N_11202,N_11227);
nand U11691 (N_11691,N_11465,N_11274);
nor U11692 (N_11692,N_11305,N_11329);
xnor U11693 (N_11693,N_11297,N_11215);
nand U11694 (N_11694,N_11362,N_11320);
or U11695 (N_11695,N_11464,N_11511);
or U11696 (N_11696,N_11408,N_11514);
xor U11697 (N_11697,N_11441,N_11360);
nor U11698 (N_11698,N_11539,N_11405);
nand U11699 (N_11699,N_11427,N_11390);
xor U11700 (N_11700,N_11568,N_11248);
nand U11701 (N_11701,N_11277,N_11306);
xnor U11702 (N_11702,N_11314,N_11377);
xor U11703 (N_11703,N_11473,N_11218);
xnor U11704 (N_11704,N_11435,N_11234);
nor U11705 (N_11705,N_11271,N_11403);
xor U11706 (N_11706,N_11319,N_11486);
xnor U11707 (N_11707,N_11404,N_11415);
nand U11708 (N_11708,N_11469,N_11354);
or U11709 (N_11709,N_11450,N_11480);
and U11710 (N_11710,N_11446,N_11400);
xor U11711 (N_11711,N_11560,N_11254);
nand U11712 (N_11712,N_11233,N_11348);
nor U11713 (N_11713,N_11241,N_11287);
nor U11714 (N_11714,N_11359,N_11428);
and U11715 (N_11715,N_11351,N_11290);
and U11716 (N_11716,N_11411,N_11433);
nand U11717 (N_11717,N_11452,N_11379);
or U11718 (N_11718,N_11258,N_11344);
and U11719 (N_11719,N_11525,N_11580);
xor U11720 (N_11720,N_11528,N_11583);
nor U11721 (N_11721,N_11372,N_11373);
nand U11722 (N_11722,N_11255,N_11524);
xor U11723 (N_11723,N_11538,N_11587);
or U11724 (N_11724,N_11356,N_11299);
and U11725 (N_11725,N_11564,N_11401);
nand U11726 (N_11726,N_11562,N_11304);
nand U11727 (N_11727,N_11505,N_11542);
xor U11728 (N_11728,N_11236,N_11343);
nand U11729 (N_11729,N_11506,N_11283);
xor U11730 (N_11730,N_11207,N_11590);
nand U11731 (N_11731,N_11437,N_11285);
and U11732 (N_11732,N_11494,N_11554);
or U11733 (N_11733,N_11257,N_11594);
or U11734 (N_11734,N_11491,N_11358);
and U11735 (N_11735,N_11200,N_11388);
and U11736 (N_11736,N_11504,N_11550);
xor U11737 (N_11737,N_11497,N_11282);
xnor U11738 (N_11738,N_11308,N_11383);
or U11739 (N_11739,N_11276,N_11598);
or U11740 (N_11740,N_11563,N_11421);
and U11741 (N_11741,N_11395,N_11330);
nand U11742 (N_11742,N_11488,N_11252);
nor U11743 (N_11743,N_11561,N_11370);
nor U11744 (N_11744,N_11345,N_11364);
xor U11745 (N_11745,N_11300,N_11532);
xor U11746 (N_11746,N_11366,N_11461);
nand U11747 (N_11747,N_11226,N_11365);
xor U11748 (N_11748,N_11220,N_11310);
nor U11749 (N_11749,N_11483,N_11418);
nand U11750 (N_11750,N_11447,N_11599);
nand U11751 (N_11751,N_11367,N_11264);
or U11752 (N_11752,N_11326,N_11341);
xnor U11753 (N_11753,N_11492,N_11396);
xor U11754 (N_11754,N_11520,N_11334);
xnor U11755 (N_11755,N_11286,N_11536);
nor U11756 (N_11756,N_11424,N_11349);
nor U11757 (N_11757,N_11331,N_11407);
xnor U11758 (N_11758,N_11275,N_11211);
and U11759 (N_11759,N_11376,N_11293);
nor U11760 (N_11760,N_11398,N_11273);
nor U11761 (N_11761,N_11534,N_11342);
and U11762 (N_11762,N_11412,N_11256);
nor U11763 (N_11763,N_11425,N_11460);
xnor U11764 (N_11764,N_11261,N_11545);
nor U11765 (N_11765,N_11369,N_11489);
and U11766 (N_11766,N_11417,N_11566);
nand U11767 (N_11767,N_11440,N_11361);
xor U11768 (N_11768,N_11573,N_11406);
or U11769 (N_11769,N_11537,N_11340);
and U11770 (N_11770,N_11263,N_11515);
and U11771 (N_11771,N_11385,N_11214);
or U11772 (N_11772,N_11553,N_11462);
nand U11773 (N_11773,N_11266,N_11589);
nor U11774 (N_11774,N_11510,N_11311);
xor U11775 (N_11775,N_11309,N_11298);
nor U11776 (N_11776,N_11577,N_11454);
xnor U11777 (N_11777,N_11474,N_11592);
nand U11778 (N_11778,N_11216,N_11312);
and U11779 (N_11779,N_11374,N_11444);
xnor U11780 (N_11780,N_11484,N_11355);
nand U11781 (N_11781,N_11426,N_11468);
and U11782 (N_11782,N_11502,N_11301);
xnor U11783 (N_11783,N_11581,N_11579);
and U11784 (N_11784,N_11546,N_11389);
nand U11785 (N_11785,N_11498,N_11339);
nand U11786 (N_11786,N_11295,N_11393);
xnor U11787 (N_11787,N_11434,N_11237);
or U11788 (N_11788,N_11512,N_11249);
or U11789 (N_11789,N_11353,N_11210);
xnor U11790 (N_11790,N_11472,N_11289);
xnor U11791 (N_11791,N_11551,N_11438);
and U11792 (N_11792,N_11391,N_11387);
nand U11793 (N_11793,N_11333,N_11409);
nand U11794 (N_11794,N_11244,N_11490);
or U11795 (N_11795,N_11503,N_11467);
or U11796 (N_11796,N_11201,N_11567);
nor U11797 (N_11797,N_11419,N_11206);
xnor U11798 (N_11798,N_11529,N_11380);
xnor U11799 (N_11799,N_11239,N_11243);
or U11800 (N_11800,N_11417,N_11276);
and U11801 (N_11801,N_11396,N_11504);
xor U11802 (N_11802,N_11518,N_11376);
nand U11803 (N_11803,N_11421,N_11417);
nand U11804 (N_11804,N_11537,N_11335);
or U11805 (N_11805,N_11505,N_11562);
or U11806 (N_11806,N_11355,N_11345);
or U11807 (N_11807,N_11577,N_11412);
and U11808 (N_11808,N_11588,N_11339);
xnor U11809 (N_11809,N_11371,N_11362);
and U11810 (N_11810,N_11336,N_11298);
nand U11811 (N_11811,N_11457,N_11503);
nor U11812 (N_11812,N_11364,N_11597);
and U11813 (N_11813,N_11286,N_11470);
nand U11814 (N_11814,N_11422,N_11227);
nand U11815 (N_11815,N_11563,N_11290);
nand U11816 (N_11816,N_11495,N_11206);
or U11817 (N_11817,N_11286,N_11531);
nand U11818 (N_11818,N_11245,N_11432);
nor U11819 (N_11819,N_11358,N_11457);
nor U11820 (N_11820,N_11563,N_11533);
xor U11821 (N_11821,N_11516,N_11491);
nand U11822 (N_11822,N_11208,N_11386);
nor U11823 (N_11823,N_11431,N_11596);
xor U11824 (N_11824,N_11446,N_11334);
nor U11825 (N_11825,N_11358,N_11587);
or U11826 (N_11826,N_11398,N_11468);
nand U11827 (N_11827,N_11237,N_11568);
or U11828 (N_11828,N_11244,N_11342);
nor U11829 (N_11829,N_11412,N_11499);
nor U11830 (N_11830,N_11404,N_11551);
nor U11831 (N_11831,N_11381,N_11239);
nor U11832 (N_11832,N_11350,N_11414);
nor U11833 (N_11833,N_11221,N_11278);
xnor U11834 (N_11834,N_11549,N_11516);
nand U11835 (N_11835,N_11304,N_11345);
and U11836 (N_11836,N_11380,N_11532);
nor U11837 (N_11837,N_11553,N_11276);
xnor U11838 (N_11838,N_11477,N_11394);
xor U11839 (N_11839,N_11401,N_11413);
and U11840 (N_11840,N_11383,N_11232);
nand U11841 (N_11841,N_11561,N_11309);
xnor U11842 (N_11842,N_11575,N_11540);
nand U11843 (N_11843,N_11493,N_11404);
nor U11844 (N_11844,N_11263,N_11507);
nand U11845 (N_11845,N_11411,N_11473);
nand U11846 (N_11846,N_11353,N_11342);
nand U11847 (N_11847,N_11523,N_11325);
nor U11848 (N_11848,N_11562,N_11514);
or U11849 (N_11849,N_11390,N_11490);
nor U11850 (N_11850,N_11489,N_11375);
xor U11851 (N_11851,N_11584,N_11405);
or U11852 (N_11852,N_11545,N_11305);
nor U11853 (N_11853,N_11495,N_11235);
xnor U11854 (N_11854,N_11287,N_11567);
nand U11855 (N_11855,N_11324,N_11214);
xor U11856 (N_11856,N_11301,N_11476);
nand U11857 (N_11857,N_11309,N_11435);
or U11858 (N_11858,N_11247,N_11375);
or U11859 (N_11859,N_11539,N_11301);
xnor U11860 (N_11860,N_11349,N_11499);
nand U11861 (N_11861,N_11409,N_11536);
xor U11862 (N_11862,N_11398,N_11452);
nor U11863 (N_11863,N_11366,N_11486);
xnor U11864 (N_11864,N_11384,N_11291);
nand U11865 (N_11865,N_11472,N_11257);
and U11866 (N_11866,N_11478,N_11261);
xor U11867 (N_11867,N_11443,N_11263);
or U11868 (N_11868,N_11286,N_11412);
or U11869 (N_11869,N_11416,N_11554);
or U11870 (N_11870,N_11423,N_11374);
xor U11871 (N_11871,N_11414,N_11462);
nor U11872 (N_11872,N_11425,N_11379);
or U11873 (N_11873,N_11542,N_11256);
xnor U11874 (N_11874,N_11255,N_11458);
and U11875 (N_11875,N_11405,N_11265);
nand U11876 (N_11876,N_11524,N_11519);
nand U11877 (N_11877,N_11551,N_11498);
or U11878 (N_11878,N_11506,N_11370);
or U11879 (N_11879,N_11477,N_11246);
or U11880 (N_11880,N_11441,N_11299);
nor U11881 (N_11881,N_11253,N_11399);
nand U11882 (N_11882,N_11400,N_11405);
or U11883 (N_11883,N_11303,N_11373);
or U11884 (N_11884,N_11269,N_11258);
nand U11885 (N_11885,N_11400,N_11302);
and U11886 (N_11886,N_11561,N_11388);
or U11887 (N_11887,N_11497,N_11217);
nor U11888 (N_11888,N_11322,N_11266);
and U11889 (N_11889,N_11539,N_11409);
and U11890 (N_11890,N_11306,N_11543);
nand U11891 (N_11891,N_11214,N_11465);
nand U11892 (N_11892,N_11532,N_11363);
nand U11893 (N_11893,N_11277,N_11430);
nand U11894 (N_11894,N_11302,N_11266);
or U11895 (N_11895,N_11501,N_11388);
or U11896 (N_11896,N_11367,N_11429);
or U11897 (N_11897,N_11545,N_11291);
xnor U11898 (N_11898,N_11575,N_11409);
xor U11899 (N_11899,N_11201,N_11399);
nor U11900 (N_11900,N_11436,N_11507);
and U11901 (N_11901,N_11460,N_11494);
or U11902 (N_11902,N_11222,N_11265);
and U11903 (N_11903,N_11531,N_11374);
nor U11904 (N_11904,N_11273,N_11380);
xnor U11905 (N_11905,N_11383,N_11587);
xnor U11906 (N_11906,N_11496,N_11452);
or U11907 (N_11907,N_11502,N_11517);
nor U11908 (N_11908,N_11392,N_11513);
or U11909 (N_11909,N_11314,N_11349);
or U11910 (N_11910,N_11561,N_11482);
xnor U11911 (N_11911,N_11547,N_11456);
or U11912 (N_11912,N_11306,N_11400);
xor U11913 (N_11913,N_11298,N_11519);
or U11914 (N_11914,N_11519,N_11476);
nor U11915 (N_11915,N_11416,N_11285);
nand U11916 (N_11916,N_11505,N_11208);
nor U11917 (N_11917,N_11382,N_11275);
nand U11918 (N_11918,N_11518,N_11247);
xnor U11919 (N_11919,N_11412,N_11454);
nand U11920 (N_11920,N_11246,N_11304);
nor U11921 (N_11921,N_11338,N_11474);
nand U11922 (N_11922,N_11440,N_11481);
nand U11923 (N_11923,N_11483,N_11394);
xor U11924 (N_11924,N_11394,N_11424);
xor U11925 (N_11925,N_11292,N_11551);
nand U11926 (N_11926,N_11566,N_11590);
and U11927 (N_11927,N_11262,N_11295);
or U11928 (N_11928,N_11342,N_11344);
nand U11929 (N_11929,N_11301,N_11451);
nor U11930 (N_11930,N_11201,N_11503);
or U11931 (N_11931,N_11348,N_11312);
nand U11932 (N_11932,N_11317,N_11307);
or U11933 (N_11933,N_11386,N_11324);
nor U11934 (N_11934,N_11358,N_11438);
or U11935 (N_11935,N_11531,N_11278);
xnor U11936 (N_11936,N_11346,N_11353);
and U11937 (N_11937,N_11428,N_11588);
and U11938 (N_11938,N_11383,N_11577);
or U11939 (N_11939,N_11371,N_11328);
or U11940 (N_11940,N_11304,N_11269);
nand U11941 (N_11941,N_11379,N_11268);
or U11942 (N_11942,N_11309,N_11248);
nand U11943 (N_11943,N_11292,N_11293);
nand U11944 (N_11944,N_11391,N_11233);
nand U11945 (N_11945,N_11266,N_11258);
xnor U11946 (N_11946,N_11281,N_11499);
xnor U11947 (N_11947,N_11361,N_11597);
or U11948 (N_11948,N_11300,N_11269);
nor U11949 (N_11949,N_11385,N_11546);
and U11950 (N_11950,N_11484,N_11528);
xnor U11951 (N_11951,N_11315,N_11216);
nand U11952 (N_11952,N_11470,N_11428);
nand U11953 (N_11953,N_11291,N_11386);
nor U11954 (N_11954,N_11503,N_11360);
nor U11955 (N_11955,N_11390,N_11461);
nor U11956 (N_11956,N_11339,N_11561);
nor U11957 (N_11957,N_11427,N_11252);
xor U11958 (N_11958,N_11331,N_11516);
xor U11959 (N_11959,N_11487,N_11542);
xor U11960 (N_11960,N_11504,N_11224);
or U11961 (N_11961,N_11493,N_11337);
or U11962 (N_11962,N_11239,N_11465);
xnor U11963 (N_11963,N_11317,N_11327);
xor U11964 (N_11964,N_11311,N_11240);
nand U11965 (N_11965,N_11495,N_11532);
and U11966 (N_11966,N_11372,N_11396);
xor U11967 (N_11967,N_11535,N_11218);
or U11968 (N_11968,N_11255,N_11535);
xor U11969 (N_11969,N_11366,N_11598);
nand U11970 (N_11970,N_11515,N_11368);
nand U11971 (N_11971,N_11401,N_11562);
nand U11972 (N_11972,N_11526,N_11451);
or U11973 (N_11973,N_11293,N_11486);
and U11974 (N_11974,N_11352,N_11505);
nand U11975 (N_11975,N_11299,N_11329);
xor U11976 (N_11976,N_11479,N_11360);
xnor U11977 (N_11977,N_11242,N_11252);
nor U11978 (N_11978,N_11248,N_11461);
or U11979 (N_11979,N_11254,N_11503);
xnor U11980 (N_11980,N_11475,N_11435);
nor U11981 (N_11981,N_11493,N_11435);
nand U11982 (N_11982,N_11436,N_11537);
and U11983 (N_11983,N_11589,N_11556);
or U11984 (N_11984,N_11392,N_11364);
nand U11985 (N_11985,N_11589,N_11483);
xor U11986 (N_11986,N_11408,N_11530);
or U11987 (N_11987,N_11575,N_11437);
and U11988 (N_11988,N_11570,N_11363);
nand U11989 (N_11989,N_11448,N_11434);
nor U11990 (N_11990,N_11465,N_11225);
nor U11991 (N_11991,N_11285,N_11504);
nand U11992 (N_11992,N_11208,N_11560);
xor U11993 (N_11993,N_11547,N_11397);
or U11994 (N_11994,N_11397,N_11267);
xnor U11995 (N_11995,N_11550,N_11529);
xor U11996 (N_11996,N_11444,N_11237);
or U11997 (N_11997,N_11388,N_11457);
or U11998 (N_11998,N_11552,N_11457);
nand U11999 (N_11999,N_11413,N_11526);
nor U12000 (N_12000,N_11896,N_11678);
or U12001 (N_12001,N_11979,N_11984);
nor U12002 (N_12002,N_11692,N_11838);
nor U12003 (N_12003,N_11869,N_11889);
nor U12004 (N_12004,N_11879,N_11609);
xor U12005 (N_12005,N_11722,N_11835);
nor U12006 (N_12006,N_11618,N_11898);
nand U12007 (N_12007,N_11754,N_11736);
and U12008 (N_12008,N_11657,N_11630);
xor U12009 (N_12009,N_11848,N_11825);
xor U12010 (N_12010,N_11847,N_11788);
nor U12011 (N_12011,N_11923,N_11855);
nand U12012 (N_12012,N_11769,N_11715);
xnor U12013 (N_12013,N_11802,N_11860);
xor U12014 (N_12014,N_11940,N_11866);
xnor U12015 (N_12015,N_11737,N_11850);
xnor U12016 (N_12016,N_11702,N_11627);
nor U12017 (N_12017,N_11809,N_11871);
or U12018 (N_12018,N_11805,N_11713);
nor U12019 (N_12019,N_11995,N_11697);
xnor U12020 (N_12020,N_11915,N_11768);
or U12021 (N_12021,N_11732,N_11971);
and U12022 (N_12022,N_11683,N_11632);
and U12023 (N_12023,N_11767,N_11990);
nand U12024 (N_12024,N_11677,N_11749);
xor U12025 (N_12025,N_11910,N_11635);
nand U12026 (N_12026,N_11956,N_11913);
nor U12027 (N_12027,N_11942,N_11954);
and U12028 (N_12028,N_11718,N_11777);
or U12029 (N_12029,N_11804,N_11872);
or U12030 (N_12030,N_11852,N_11779);
nor U12031 (N_12031,N_11798,N_11792);
or U12032 (N_12032,N_11636,N_11953);
nand U12033 (N_12033,N_11861,N_11967);
xor U12034 (N_12034,N_11960,N_11880);
xnor U12035 (N_12035,N_11631,N_11884);
nor U12036 (N_12036,N_11753,N_11959);
or U12037 (N_12037,N_11729,N_11914);
or U12038 (N_12038,N_11989,N_11890);
and U12039 (N_12039,N_11602,N_11626);
or U12040 (N_12040,N_11703,N_11646);
and U12041 (N_12041,N_11909,N_11751);
or U12042 (N_12042,N_11625,N_11854);
nor U12043 (N_12043,N_11998,N_11795);
and U12044 (N_12044,N_11694,N_11710);
or U12045 (N_12045,N_11965,N_11653);
nor U12046 (N_12046,N_11658,N_11641);
and U12047 (N_12047,N_11778,N_11799);
and U12048 (N_12048,N_11770,N_11665);
and U12049 (N_12049,N_11862,N_11681);
nor U12050 (N_12050,N_11743,N_11711);
and U12051 (N_12051,N_11654,N_11992);
or U12052 (N_12052,N_11708,N_11873);
xnor U12053 (N_12053,N_11687,N_11925);
xnor U12054 (N_12054,N_11933,N_11941);
xnor U12055 (N_12055,N_11733,N_11976);
xor U12056 (N_12056,N_11858,N_11801);
or U12057 (N_12057,N_11755,N_11741);
nor U12058 (N_12058,N_11904,N_11642);
and U12059 (N_12059,N_11859,N_11846);
xor U12060 (N_12060,N_11975,N_11922);
xnor U12061 (N_12061,N_11887,N_11908);
xnor U12062 (N_12062,N_11693,N_11810);
xor U12063 (N_12063,N_11747,N_11652);
and U12064 (N_12064,N_11669,N_11765);
nor U12065 (N_12065,N_11757,N_11981);
or U12066 (N_12066,N_11885,N_11853);
and U12067 (N_12067,N_11695,N_11672);
xor U12068 (N_12068,N_11845,N_11704);
nand U12069 (N_12069,N_11948,N_11706);
and U12070 (N_12070,N_11790,N_11803);
or U12071 (N_12071,N_11963,N_11993);
xnor U12072 (N_12072,N_11621,N_11728);
nand U12073 (N_12073,N_11856,N_11814);
xor U12074 (N_12074,N_11837,N_11726);
nand U12075 (N_12075,N_11813,N_11603);
nor U12076 (N_12076,N_11902,N_11829);
nor U12077 (N_12077,N_11916,N_11800);
nor U12078 (N_12078,N_11828,N_11707);
nor U12079 (N_12079,N_11774,N_11867);
or U12080 (N_12080,N_11870,N_11951);
and U12081 (N_12081,N_11673,N_11667);
and U12082 (N_12082,N_11688,N_11727);
and U12083 (N_12083,N_11857,N_11629);
nand U12084 (N_12084,N_11615,N_11750);
nor U12085 (N_12085,N_11843,N_11842);
nand U12086 (N_12086,N_11931,N_11983);
and U12087 (N_12087,N_11991,N_11988);
and U12088 (N_12088,N_11608,N_11651);
nor U12089 (N_12089,N_11700,N_11886);
nand U12090 (N_12090,N_11781,N_11827);
xor U12091 (N_12091,N_11738,N_11771);
nand U12092 (N_12092,N_11675,N_11806);
or U12093 (N_12093,N_11935,N_11607);
or U12094 (N_12094,N_11999,N_11878);
xnor U12095 (N_12095,N_11811,N_11920);
or U12096 (N_12096,N_11944,N_11637);
or U12097 (N_12097,N_11823,N_11901);
nand U12098 (N_12098,N_11624,N_11900);
nor U12099 (N_12099,N_11875,N_11662);
or U12100 (N_12100,N_11968,N_11907);
and U12101 (N_12101,N_11773,N_11994);
xor U12102 (N_12102,N_11696,N_11936);
and U12103 (N_12103,N_11744,N_11705);
and U12104 (N_12104,N_11740,N_11943);
nand U12105 (N_12105,N_11912,N_11776);
or U12106 (N_12106,N_11945,N_11611);
nor U12107 (N_12107,N_11946,N_11821);
nand U12108 (N_12108,N_11671,N_11689);
nand U12109 (N_12109,N_11698,N_11863);
or U12110 (N_12110,N_11721,N_11610);
nand U12111 (N_12111,N_11832,N_11834);
or U12112 (N_12112,N_11785,N_11731);
nor U12113 (N_12113,N_11883,N_11679);
and U12114 (N_12114,N_11868,N_11633);
nand U12115 (N_12115,N_11882,N_11762);
xor U12116 (N_12116,N_11605,N_11796);
nor U12117 (N_12117,N_11760,N_11623);
nor U12118 (N_12118,N_11962,N_11905);
nor U12119 (N_12119,N_11972,N_11808);
nor U12120 (N_12120,N_11978,N_11840);
xor U12121 (N_12121,N_11685,N_11864);
nand U12122 (N_12122,N_11682,N_11691);
or U12123 (N_12123,N_11830,N_11877);
nand U12124 (N_12124,N_11717,N_11622);
nor U12125 (N_12125,N_11930,N_11874);
nor U12126 (N_12126,N_11664,N_11929);
or U12127 (N_12127,N_11600,N_11670);
or U12128 (N_12128,N_11911,N_11894);
nand U12129 (N_12129,N_11977,N_11906);
and U12130 (N_12130,N_11876,N_11899);
or U12131 (N_12131,N_11612,N_11759);
or U12132 (N_12132,N_11649,N_11820);
nor U12133 (N_12133,N_11724,N_11746);
nand U12134 (N_12134,N_11921,N_11684);
xor U12135 (N_12135,N_11739,N_11614);
nand U12136 (N_12136,N_11761,N_11938);
nor U12137 (N_12137,N_11985,N_11644);
xor U12138 (N_12138,N_11734,N_11676);
nand U12139 (N_12139,N_11789,N_11783);
nor U12140 (N_12140,N_11613,N_11974);
or U12141 (N_12141,N_11819,N_11639);
xnor U12142 (N_12142,N_11888,N_11780);
nor U12143 (N_12143,N_11797,N_11714);
nor U12144 (N_12144,N_11952,N_11833);
or U12145 (N_12145,N_11961,N_11817);
or U12146 (N_12146,N_11643,N_11659);
or U12147 (N_12147,N_11604,N_11616);
nor U12148 (N_12148,N_11656,N_11824);
nand U12149 (N_12149,N_11674,N_11947);
nand U12150 (N_12150,N_11836,N_11786);
xnor U12151 (N_12151,N_11892,N_11663);
xnor U12152 (N_12152,N_11865,N_11903);
and U12153 (N_12153,N_11895,N_11793);
xor U12154 (N_12154,N_11668,N_11709);
and U12155 (N_12155,N_11969,N_11849);
nand U12156 (N_12156,N_11686,N_11617);
xor U12157 (N_12157,N_11917,N_11660);
xor U12158 (N_12158,N_11807,N_11628);
nand U12159 (N_12159,N_11716,N_11742);
or U12160 (N_12160,N_11996,N_11766);
or U12161 (N_12161,N_11949,N_11794);
or U12162 (N_12162,N_11937,N_11745);
xnor U12163 (N_12163,N_11723,N_11939);
or U12164 (N_12164,N_11634,N_11973);
xor U12165 (N_12165,N_11841,N_11666);
xnor U12166 (N_12166,N_11791,N_11712);
or U12167 (N_12167,N_11606,N_11918);
and U12168 (N_12168,N_11897,N_11881);
nor U12169 (N_12169,N_11851,N_11987);
xnor U12170 (N_12170,N_11764,N_11720);
xnor U12171 (N_12171,N_11645,N_11950);
nand U12172 (N_12172,N_11680,N_11756);
nor U12173 (N_12173,N_11752,N_11839);
xor U12174 (N_12174,N_11730,N_11844);
xor U12175 (N_12175,N_11640,N_11775);
and U12176 (N_12176,N_11772,N_11701);
xnor U12177 (N_12177,N_11919,N_11815);
or U12178 (N_12178,N_11650,N_11661);
and U12179 (N_12179,N_11826,N_11699);
and U12180 (N_12180,N_11648,N_11822);
and U12181 (N_12181,N_11818,N_11831);
nor U12182 (N_12182,N_11782,N_11927);
and U12183 (N_12183,N_11964,N_11784);
or U12184 (N_12184,N_11924,N_11955);
xnor U12185 (N_12185,N_11966,N_11982);
and U12186 (N_12186,N_11620,N_11997);
and U12187 (N_12187,N_11763,N_11928);
and U12188 (N_12188,N_11980,N_11958);
or U12189 (N_12189,N_11758,N_11725);
or U12190 (N_12190,N_11619,N_11812);
and U12191 (N_12191,N_11787,N_11893);
or U12192 (N_12192,N_11638,N_11735);
xor U12193 (N_12193,N_11932,N_11748);
xnor U12194 (N_12194,N_11926,N_11647);
xor U12195 (N_12195,N_11690,N_11957);
nor U12196 (N_12196,N_11986,N_11601);
nand U12197 (N_12197,N_11719,N_11934);
nand U12198 (N_12198,N_11655,N_11970);
and U12199 (N_12199,N_11891,N_11816);
nor U12200 (N_12200,N_11870,N_11610);
or U12201 (N_12201,N_11651,N_11773);
xnor U12202 (N_12202,N_11992,N_11813);
and U12203 (N_12203,N_11826,N_11773);
nand U12204 (N_12204,N_11626,N_11621);
nand U12205 (N_12205,N_11732,N_11887);
or U12206 (N_12206,N_11893,N_11974);
or U12207 (N_12207,N_11748,N_11838);
and U12208 (N_12208,N_11809,N_11718);
nor U12209 (N_12209,N_11929,N_11645);
and U12210 (N_12210,N_11978,N_11927);
nand U12211 (N_12211,N_11904,N_11620);
nor U12212 (N_12212,N_11758,N_11855);
or U12213 (N_12213,N_11604,N_11738);
nand U12214 (N_12214,N_11926,N_11600);
xnor U12215 (N_12215,N_11807,N_11831);
and U12216 (N_12216,N_11869,N_11834);
xor U12217 (N_12217,N_11821,N_11833);
and U12218 (N_12218,N_11991,N_11775);
or U12219 (N_12219,N_11718,N_11738);
and U12220 (N_12220,N_11964,N_11826);
or U12221 (N_12221,N_11739,N_11695);
nor U12222 (N_12222,N_11877,N_11887);
and U12223 (N_12223,N_11901,N_11789);
nand U12224 (N_12224,N_11679,N_11761);
and U12225 (N_12225,N_11838,N_11717);
nand U12226 (N_12226,N_11774,N_11668);
xor U12227 (N_12227,N_11791,N_11604);
and U12228 (N_12228,N_11722,N_11633);
xnor U12229 (N_12229,N_11637,N_11922);
xnor U12230 (N_12230,N_11888,N_11621);
or U12231 (N_12231,N_11721,N_11704);
nor U12232 (N_12232,N_11887,N_11657);
xor U12233 (N_12233,N_11922,N_11960);
nand U12234 (N_12234,N_11958,N_11749);
or U12235 (N_12235,N_11692,N_11933);
nor U12236 (N_12236,N_11937,N_11696);
or U12237 (N_12237,N_11678,N_11851);
xor U12238 (N_12238,N_11738,N_11808);
or U12239 (N_12239,N_11949,N_11685);
nor U12240 (N_12240,N_11783,N_11812);
nand U12241 (N_12241,N_11896,N_11843);
nor U12242 (N_12242,N_11800,N_11945);
nand U12243 (N_12243,N_11886,N_11769);
xnor U12244 (N_12244,N_11671,N_11730);
and U12245 (N_12245,N_11754,N_11946);
xnor U12246 (N_12246,N_11852,N_11946);
and U12247 (N_12247,N_11889,N_11640);
nand U12248 (N_12248,N_11666,N_11736);
xnor U12249 (N_12249,N_11720,N_11627);
nor U12250 (N_12250,N_11622,N_11791);
and U12251 (N_12251,N_11854,N_11606);
and U12252 (N_12252,N_11757,N_11932);
xnor U12253 (N_12253,N_11910,N_11936);
nor U12254 (N_12254,N_11896,N_11851);
xor U12255 (N_12255,N_11898,N_11952);
and U12256 (N_12256,N_11670,N_11870);
or U12257 (N_12257,N_11994,N_11687);
and U12258 (N_12258,N_11725,N_11908);
xnor U12259 (N_12259,N_11874,N_11950);
nor U12260 (N_12260,N_11899,N_11670);
nor U12261 (N_12261,N_11608,N_11994);
nand U12262 (N_12262,N_11860,N_11988);
or U12263 (N_12263,N_11794,N_11854);
or U12264 (N_12264,N_11806,N_11875);
xnor U12265 (N_12265,N_11735,N_11991);
and U12266 (N_12266,N_11928,N_11786);
nand U12267 (N_12267,N_11602,N_11907);
nor U12268 (N_12268,N_11806,N_11694);
or U12269 (N_12269,N_11815,N_11921);
nor U12270 (N_12270,N_11999,N_11936);
xnor U12271 (N_12271,N_11689,N_11997);
xor U12272 (N_12272,N_11792,N_11840);
nor U12273 (N_12273,N_11762,N_11731);
xnor U12274 (N_12274,N_11762,N_11899);
nor U12275 (N_12275,N_11688,N_11626);
or U12276 (N_12276,N_11918,N_11950);
nor U12277 (N_12277,N_11791,N_11935);
nand U12278 (N_12278,N_11878,N_11823);
and U12279 (N_12279,N_11790,N_11702);
nor U12280 (N_12280,N_11775,N_11607);
or U12281 (N_12281,N_11984,N_11778);
and U12282 (N_12282,N_11908,N_11931);
nand U12283 (N_12283,N_11817,N_11752);
nor U12284 (N_12284,N_11870,N_11641);
nand U12285 (N_12285,N_11624,N_11819);
or U12286 (N_12286,N_11626,N_11972);
or U12287 (N_12287,N_11656,N_11682);
nor U12288 (N_12288,N_11887,N_11935);
nand U12289 (N_12289,N_11700,N_11653);
or U12290 (N_12290,N_11757,N_11899);
nor U12291 (N_12291,N_11787,N_11762);
and U12292 (N_12292,N_11802,N_11759);
nand U12293 (N_12293,N_11634,N_11710);
nor U12294 (N_12294,N_11906,N_11746);
xor U12295 (N_12295,N_11857,N_11740);
nor U12296 (N_12296,N_11961,N_11988);
xor U12297 (N_12297,N_11910,N_11841);
nand U12298 (N_12298,N_11760,N_11745);
nor U12299 (N_12299,N_11750,N_11721);
xnor U12300 (N_12300,N_11746,N_11715);
and U12301 (N_12301,N_11714,N_11910);
nor U12302 (N_12302,N_11930,N_11640);
and U12303 (N_12303,N_11687,N_11785);
xor U12304 (N_12304,N_11600,N_11708);
nand U12305 (N_12305,N_11883,N_11843);
or U12306 (N_12306,N_11651,N_11960);
nor U12307 (N_12307,N_11671,N_11790);
or U12308 (N_12308,N_11933,N_11780);
and U12309 (N_12309,N_11945,N_11711);
nor U12310 (N_12310,N_11653,N_11620);
nand U12311 (N_12311,N_11963,N_11736);
or U12312 (N_12312,N_11883,N_11869);
and U12313 (N_12313,N_11988,N_11809);
and U12314 (N_12314,N_11740,N_11702);
nand U12315 (N_12315,N_11782,N_11796);
xor U12316 (N_12316,N_11852,N_11703);
nand U12317 (N_12317,N_11735,N_11747);
nor U12318 (N_12318,N_11841,N_11832);
xnor U12319 (N_12319,N_11974,N_11647);
and U12320 (N_12320,N_11825,N_11768);
nor U12321 (N_12321,N_11713,N_11878);
nand U12322 (N_12322,N_11821,N_11868);
and U12323 (N_12323,N_11769,N_11971);
nor U12324 (N_12324,N_11660,N_11843);
and U12325 (N_12325,N_11766,N_11831);
nand U12326 (N_12326,N_11782,N_11628);
and U12327 (N_12327,N_11840,N_11899);
and U12328 (N_12328,N_11690,N_11737);
xnor U12329 (N_12329,N_11627,N_11807);
xor U12330 (N_12330,N_11981,N_11678);
or U12331 (N_12331,N_11812,N_11793);
xor U12332 (N_12332,N_11773,N_11766);
nor U12333 (N_12333,N_11604,N_11965);
nor U12334 (N_12334,N_11773,N_11751);
and U12335 (N_12335,N_11651,N_11769);
xnor U12336 (N_12336,N_11605,N_11917);
and U12337 (N_12337,N_11693,N_11646);
nor U12338 (N_12338,N_11650,N_11920);
xnor U12339 (N_12339,N_11855,N_11682);
and U12340 (N_12340,N_11944,N_11974);
xor U12341 (N_12341,N_11988,N_11613);
nand U12342 (N_12342,N_11894,N_11740);
nand U12343 (N_12343,N_11714,N_11758);
and U12344 (N_12344,N_11817,N_11718);
nor U12345 (N_12345,N_11708,N_11855);
and U12346 (N_12346,N_11703,N_11791);
nor U12347 (N_12347,N_11762,N_11604);
and U12348 (N_12348,N_11784,N_11781);
nor U12349 (N_12349,N_11714,N_11738);
nand U12350 (N_12350,N_11631,N_11974);
nand U12351 (N_12351,N_11683,N_11823);
nor U12352 (N_12352,N_11669,N_11747);
and U12353 (N_12353,N_11939,N_11669);
nand U12354 (N_12354,N_11733,N_11978);
or U12355 (N_12355,N_11897,N_11947);
nand U12356 (N_12356,N_11826,N_11731);
and U12357 (N_12357,N_11884,N_11688);
or U12358 (N_12358,N_11818,N_11982);
nand U12359 (N_12359,N_11644,N_11701);
nand U12360 (N_12360,N_11785,N_11606);
nor U12361 (N_12361,N_11978,N_11775);
nor U12362 (N_12362,N_11602,N_11994);
and U12363 (N_12363,N_11713,N_11644);
nand U12364 (N_12364,N_11760,N_11990);
and U12365 (N_12365,N_11975,N_11796);
nand U12366 (N_12366,N_11938,N_11828);
xnor U12367 (N_12367,N_11606,N_11966);
xnor U12368 (N_12368,N_11644,N_11786);
xnor U12369 (N_12369,N_11988,N_11635);
nor U12370 (N_12370,N_11714,N_11759);
xnor U12371 (N_12371,N_11964,N_11951);
nor U12372 (N_12372,N_11671,N_11743);
xnor U12373 (N_12373,N_11880,N_11714);
and U12374 (N_12374,N_11902,N_11647);
nor U12375 (N_12375,N_11938,N_11630);
nor U12376 (N_12376,N_11795,N_11636);
xnor U12377 (N_12377,N_11602,N_11764);
nor U12378 (N_12378,N_11953,N_11729);
or U12379 (N_12379,N_11832,N_11623);
nand U12380 (N_12380,N_11971,N_11863);
and U12381 (N_12381,N_11678,N_11625);
nand U12382 (N_12382,N_11926,N_11853);
nand U12383 (N_12383,N_11907,N_11710);
or U12384 (N_12384,N_11957,N_11857);
or U12385 (N_12385,N_11634,N_11693);
or U12386 (N_12386,N_11855,N_11893);
or U12387 (N_12387,N_11761,N_11936);
xnor U12388 (N_12388,N_11672,N_11637);
and U12389 (N_12389,N_11718,N_11887);
or U12390 (N_12390,N_11710,N_11787);
nand U12391 (N_12391,N_11927,N_11945);
and U12392 (N_12392,N_11816,N_11926);
nor U12393 (N_12393,N_11998,N_11843);
xnor U12394 (N_12394,N_11907,N_11813);
or U12395 (N_12395,N_11875,N_11970);
nand U12396 (N_12396,N_11812,N_11833);
xnor U12397 (N_12397,N_11638,N_11675);
xor U12398 (N_12398,N_11934,N_11613);
nor U12399 (N_12399,N_11700,N_11800);
xor U12400 (N_12400,N_12343,N_12064);
nor U12401 (N_12401,N_12154,N_12376);
or U12402 (N_12402,N_12012,N_12128);
nor U12403 (N_12403,N_12312,N_12230);
nor U12404 (N_12404,N_12037,N_12075);
nor U12405 (N_12405,N_12236,N_12097);
nor U12406 (N_12406,N_12076,N_12023);
and U12407 (N_12407,N_12375,N_12111);
and U12408 (N_12408,N_12275,N_12098);
nor U12409 (N_12409,N_12115,N_12301);
and U12410 (N_12410,N_12252,N_12271);
nor U12411 (N_12411,N_12381,N_12223);
xnor U12412 (N_12412,N_12318,N_12150);
nor U12413 (N_12413,N_12380,N_12132);
xor U12414 (N_12414,N_12277,N_12212);
nand U12415 (N_12415,N_12279,N_12069);
xnor U12416 (N_12416,N_12329,N_12260);
nand U12417 (N_12417,N_12029,N_12296);
or U12418 (N_12418,N_12203,N_12281);
or U12419 (N_12419,N_12269,N_12227);
nor U12420 (N_12420,N_12049,N_12100);
nor U12421 (N_12421,N_12226,N_12328);
nor U12422 (N_12422,N_12040,N_12104);
nand U12423 (N_12423,N_12189,N_12015);
and U12424 (N_12424,N_12047,N_12387);
xnor U12425 (N_12425,N_12370,N_12042);
or U12426 (N_12426,N_12221,N_12332);
or U12427 (N_12427,N_12021,N_12011);
and U12428 (N_12428,N_12385,N_12176);
or U12429 (N_12429,N_12129,N_12025);
nor U12430 (N_12430,N_12167,N_12398);
nor U12431 (N_12431,N_12180,N_12106);
and U12432 (N_12432,N_12182,N_12399);
nand U12433 (N_12433,N_12295,N_12079);
and U12434 (N_12434,N_12063,N_12033);
and U12435 (N_12435,N_12346,N_12026);
nor U12436 (N_12436,N_12308,N_12233);
nand U12437 (N_12437,N_12157,N_12204);
xor U12438 (N_12438,N_12373,N_12061);
or U12439 (N_12439,N_12067,N_12323);
nor U12440 (N_12440,N_12282,N_12263);
and U12441 (N_12441,N_12344,N_12261);
nor U12442 (N_12442,N_12144,N_12175);
and U12443 (N_12443,N_12056,N_12302);
and U12444 (N_12444,N_12248,N_12156);
xnor U12445 (N_12445,N_12300,N_12166);
nand U12446 (N_12446,N_12149,N_12058);
or U12447 (N_12447,N_12306,N_12137);
nor U12448 (N_12448,N_12081,N_12022);
or U12449 (N_12449,N_12065,N_12148);
nor U12450 (N_12450,N_12276,N_12341);
nand U12451 (N_12451,N_12340,N_12134);
nand U12452 (N_12452,N_12059,N_12225);
nor U12453 (N_12453,N_12146,N_12270);
and U12454 (N_12454,N_12000,N_12354);
and U12455 (N_12455,N_12294,N_12024);
and U12456 (N_12456,N_12374,N_12108);
and U12457 (N_12457,N_12322,N_12359);
and U12458 (N_12458,N_12384,N_12034);
xor U12459 (N_12459,N_12351,N_12158);
and U12460 (N_12460,N_12288,N_12237);
nand U12461 (N_12461,N_12155,N_12043);
and U12462 (N_12462,N_12193,N_12125);
nand U12463 (N_12463,N_12215,N_12297);
xnor U12464 (N_12464,N_12319,N_12256);
nand U12465 (N_12465,N_12348,N_12030);
and U12466 (N_12466,N_12358,N_12194);
xor U12467 (N_12467,N_12084,N_12031);
and U12468 (N_12468,N_12317,N_12283);
nor U12469 (N_12469,N_12257,N_12095);
xor U12470 (N_12470,N_12377,N_12016);
or U12471 (N_12471,N_12138,N_12246);
xor U12472 (N_12472,N_12367,N_12052);
nor U12473 (N_12473,N_12174,N_12334);
nand U12474 (N_12474,N_12267,N_12038);
or U12475 (N_12475,N_12143,N_12378);
or U12476 (N_12476,N_12159,N_12187);
xor U12477 (N_12477,N_12124,N_12107);
nor U12478 (N_12478,N_12085,N_12179);
xnor U12479 (N_12479,N_12003,N_12220);
or U12480 (N_12480,N_12044,N_12219);
xor U12481 (N_12481,N_12369,N_12208);
nand U12482 (N_12482,N_12382,N_12390);
or U12483 (N_12483,N_12083,N_12185);
nand U12484 (N_12484,N_12305,N_12372);
xnor U12485 (N_12485,N_12020,N_12036);
nor U12486 (N_12486,N_12259,N_12073);
xor U12487 (N_12487,N_12184,N_12045);
nor U12488 (N_12488,N_12333,N_12360);
nand U12489 (N_12489,N_12014,N_12264);
xnor U12490 (N_12490,N_12074,N_12243);
xnor U12491 (N_12491,N_12119,N_12126);
nor U12492 (N_12492,N_12162,N_12395);
xor U12493 (N_12493,N_12213,N_12165);
and U12494 (N_12494,N_12035,N_12130);
xor U12495 (N_12495,N_12013,N_12392);
xnor U12496 (N_12496,N_12335,N_12254);
and U12497 (N_12497,N_12196,N_12088);
and U12498 (N_12498,N_12345,N_12090);
nand U12499 (N_12499,N_12087,N_12389);
or U12500 (N_12500,N_12153,N_12338);
xnor U12501 (N_12501,N_12394,N_12068);
nor U12502 (N_12502,N_12094,N_12242);
or U12503 (N_12503,N_12214,N_12139);
xnor U12504 (N_12504,N_12018,N_12353);
or U12505 (N_12505,N_12347,N_12071);
xnor U12506 (N_12506,N_12195,N_12352);
or U12507 (N_12507,N_12114,N_12320);
or U12508 (N_12508,N_12077,N_12057);
xnor U12509 (N_12509,N_12274,N_12238);
nor U12510 (N_12510,N_12321,N_12009);
xor U12511 (N_12511,N_12122,N_12231);
xnor U12512 (N_12512,N_12298,N_12164);
and U12513 (N_12513,N_12062,N_12188);
or U12514 (N_12514,N_12161,N_12050);
or U12515 (N_12515,N_12356,N_12170);
or U12516 (N_12516,N_12112,N_12209);
nor U12517 (N_12517,N_12070,N_12330);
and U12518 (N_12518,N_12113,N_12082);
and U12519 (N_12519,N_12105,N_12310);
xor U12520 (N_12520,N_12039,N_12152);
xor U12521 (N_12521,N_12285,N_12198);
nand U12522 (N_12522,N_12292,N_12217);
nand U12523 (N_12523,N_12262,N_12383);
nor U12524 (N_12524,N_12120,N_12041);
or U12525 (N_12525,N_12032,N_12171);
and U12526 (N_12526,N_12265,N_12110);
or U12527 (N_12527,N_12191,N_12304);
and U12528 (N_12528,N_12218,N_12313);
or U12529 (N_12529,N_12240,N_12361);
nor U12530 (N_12530,N_12116,N_12258);
nand U12531 (N_12531,N_12235,N_12140);
nor U12532 (N_12532,N_12117,N_12314);
and U12533 (N_12533,N_12109,N_12363);
xor U12534 (N_12534,N_12350,N_12123);
xnor U12535 (N_12535,N_12244,N_12255);
and U12536 (N_12536,N_12190,N_12206);
or U12537 (N_12537,N_12250,N_12053);
nand U12538 (N_12538,N_12096,N_12299);
nor U12539 (N_12539,N_12241,N_12247);
nand U12540 (N_12540,N_12202,N_12183);
or U12541 (N_12541,N_12207,N_12201);
xnor U12542 (N_12542,N_12397,N_12197);
or U12543 (N_12543,N_12232,N_12093);
nand U12544 (N_12544,N_12089,N_12200);
and U12545 (N_12545,N_12365,N_12133);
or U12546 (N_12546,N_12181,N_12142);
nand U12547 (N_12547,N_12136,N_12172);
xor U12548 (N_12548,N_12234,N_12001);
nand U12549 (N_12549,N_12249,N_12268);
and U12550 (N_12550,N_12121,N_12051);
xnor U12551 (N_12551,N_12251,N_12135);
nor U12552 (N_12552,N_12222,N_12278);
nand U12553 (N_12553,N_12366,N_12357);
and U12554 (N_12554,N_12386,N_12266);
nor U12555 (N_12555,N_12391,N_12055);
and U12556 (N_12556,N_12008,N_12091);
nand U12557 (N_12557,N_12368,N_12028);
nand U12558 (N_12558,N_12066,N_12192);
nor U12559 (N_12559,N_12211,N_12339);
nand U12560 (N_12560,N_12362,N_12364);
xnor U12561 (N_12561,N_12291,N_12131);
nor U12562 (N_12562,N_12303,N_12379);
nand U12563 (N_12563,N_12017,N_12006);
nand U12564 (N_12564,N_12177,N_12010);
nor U12565 (N_12565,N_12309,N_12349);
and U12566 (N_12566,N_12127,N_12393);
and U12567 (N_12567,N_12293,N_12102);
nand U12568 (N_12568,N_12054,N_12160);
and U12569 (N_12569,N_12046,N_12169);
or U12570 (N_12570,N_12173,N_12229);
or U12571 (N_12571,N_12078,N_12287);
and U12572 (N_12572,N_12342,N_12163);
and U12573 (N_12573,N_12326,N_12336);
and U12574 (N_12574,N_12103,N_12086);
xor U12575 (N_12575,N_12004,N_12331);
or U12576 (N_12576,N_12141,N_12228);
xor U12577 (N_12577,N_12019,N_12396);
xor U12578 (N_12578,N_12290,N_12325);
or U12579 (N_12579,N_12224,N_12007);
nor U12580 (N_12580,N_12118,N_12186);
or U12581 (N_12581,N_12027,N_12253);
and U12582 (N_12582,N_12337,N_12151);
or U12583 (N_12583,N_12092,N_12280);
nor U12584 (N_12584,N_12245,N_12272);
or U12585 (N_12585,N_12289,N_12199);
or U12586 (N_12586,N_12239,N_12048);
xnor U12587 (N_12587,N_12327,N_12371);
nor U12588 (N_12588,N_12388,N_12284);
nand U12589 (N_12589,N_12080,N_12315);
xnor U12590 (N_12590,N_12216,N_12101);
nand U12591 (N_12591,N_12147,N_12311);
or U12592 (N_12592,N_12205,N_12286);
nor U12593 (N_12593,N_12002,N_12307);
nand U12594 (N_12594,N_12145,N_12210);
xor U12595 (N_12595,N_12168,N_12060);
nand U12596 (N_12596,N_12316,N_12178);
nor U12597 (N_12597,N_12005,N_12324);
xor U12598 (N_12598,N_12355,N_12273);
and U12599 (N_12599,N_12072,N_12099);
and U12600 (N_12600,N_12399,N_12160);
and U12601 (N_12601,N_12163,N_12325);
xor U12602 (N_12602,N_12078,N_12238);
nand U12603 (N_12603,N_12383,N_12247);
nor U12604 (N_12604,N_12102,N_12302);
xnor U12605 (N_12605,N_12230,N_12321);
nor U12606 (N_12606,N_12048,N_12281);
or U12607 (N_12607,N_12324,N_12183);
or U12608 (N_12608,N_12335,N_12215);
and U12609 (N_12609,N_12273,N_12217);
xnor U12610 (N_12610,N_12353,N_12186);
xor U12611 (N_12611,N_12074,N_12294);
nor U12612 (N_12612,N_12386,N_12103);
xor U12613 (N_12613,N_12217,N_12102);
nand U12614 (N_12614,N_12361,N_12148);
nor U12615 (N_12615,N_12206,N_12148);
nor U12616 (N_12616,N_12166,N_12126);
nor U12617 (N_12617,N_12089,N_12026);
xnor U12618 (N_12618,N_12025,N_12285);
nor U12619 (N_12619,N_12108,N_12136);
nand U12620 (N_12620,N_12079,N_12147);
nor U12621 (N_12621,N_12065,N_12309);
xnor U12622 (N_12622,N_12343,N_12053);
nand U12623 (N_12623,N_12356,N_12394);
or U12624 (N_12624,N_12154,N_12198);
nand U12625 (N_12625,N_12134,N_12067);
nand U12626 (N_12626,N_12139,N_12259);
or U12627 (N_12627,N_12100,N_12106);
xor U12628 (N_12628,N_12234,N_12322);
and U12629 (N_12629,N_12234,N_12054);
and U12630 (N_12630,N_12297,N_12090);
and U12631 (N_12631,N_12081,N_12395);
or U12632 (N_12632,N_12014,N_12227);
nor U12633 (N_12633,N_12044,N_12174);
or U12634 (N_12634,N_12256,N_12267);
nor U12635 (N_12635,N_12031,N_12317);
nand U12636 (N_12636,N_12064,N_12394);
nand U12637 (N_12637,N_12266,N_12040);
or U12638 (N_12638,N_12302,N_12394);
or U12639 (N_12639,N_12142,N_12310);
or U12640 (N_12640,N_12077,N_12299);
xor U12641 (N_12641,N_12142,N_12159);
xor U12642 (N_12642,N_12385,N_12302);
and U12643 (N_12643,N_12106,N_12316);
nor U12644 (N_12644,N_12128,N_12311);
nand U12645 (N_12645,N_12313,N_12104);
xnor U12646 (N_12646,N_12357,N_12241);
nand U12647 (N_12647,N_12042,N_12098);
or U12648 (N_12648,N_12351,N_12305);
and U12649 (N_12649,N_12031,N_12014);
nor U12650 (N_12650,N_12119,N_12204);
xor U12651 (N_12651,N_12341,N_12051);
or U12652 (N_12652,N_12264,N_12100);
nor U12653 (N_12653,N_12261,N_12063);
nor U12654 (N_12654,N_12136,N_12013);
nor U12655 (N_12655,N_12045,N_12073);
and U12656 (N_12656,N_12280,N_12150);
xnor U12657 (N_12657,N_12048,N_12035);
nor U12658 (N_12658,N_12227,N_12394);
or U12659 (N_12659,N_12079,N_12190);
xnor U12660 (N_12660,N_12368,N_12251);
nand U12661 (N_12661,N_12061,N_12301);
and U12662 (N_12662,N_12226,N_12278);
and U12663 (N_12663,N_12386,N_12153);
xor U12664 (N_12664,N_12366,N_12348);
or U12665 (N_12665,N_12384,N_12076);
or U12666 (N_12666,N_12339,N_12212);
or U12667 (N_12667,N_12392,N_12025);
nand U12668 (N_12668,N_12124,N_12239);
nand U12669 (N_12669,N_12025,N_12028);
xnor U12670 (N_12670,N_12337,N_12130);
and U12671 (N_12671,N_12064,N_12348);
nand U12672 (N_12672,N_12035,N_12388);
nand U12673 (N_12673,N_12294,N_12071);
and U12674 (N_12674,N_12074,N_12316);
xnor U12675 (N_12675,N_12067,N_12335);
nand U12676 (N_12676,N_12138,N_12133);
xnor U12677 (N_12677,N_12053,N_12365);
nand U12678 (N_12678,N_12131,N_12290);
nand U12679 (N_12679,N_12004,N_12001);
and U12680 (N_12680,N_12182,N_12097);
and U12681 (N_12681,N_12371,N_12281);
or U12682 (N_12682,N_12068,N_12193);
xnor U12683 (N_12683,N_12000,N_12298);
and U12684 (N_12684,N_12231,N_12024);
and U12685 (N_12685,N_12048,N_12054);
xor U12686 (N_12686,N_12248,N_12119);
nor U12687 (N_12687,N_12278,N_12036);
nor U12688 (N_12688,N_12004,N_12204);
and U12689 (N_12689,N_12260,N_12120);
or U12690 (N_12690,N_12158,N_12223);
xor U12691 (N_12691,N_12224,N_12281);
nand U12692 (N_12692,N_12288,N_12303);
nor U12693 (N_12693,N_12265,N_12093);
nand U12694 (N_12694,N_12116,N_12340);
nor U12695 (N_12695,N_12225,N_12302);
xor U12696 (N_12696,N_12210,N_12391);
nand U12697 (N_12697,N_12337,N_12395);
nand U12698 (N_12698,N_12307,N_12286);
or U12699 (N_12699,N_12332,N_12048);
and U12700 (N_12700,N_12239,N_12171);
and U12701 (N_12701,N_12054,N_12386);
or U12702 (N_12702,N_12026,N_12158);
nand U12703 (N_12703,N_12155,N_12089);
nand U12704 (N_12704,N_12315,N_12319);
and U12705 (N_12705,N_12328,N_12239);
nor U12706 (N_12706,N_12054,N_12280);
or U12707 (N_12707,N_12076,N_12303);
xnor U12708 (N_12708,N_12376,N_12153);
xor U12709 (N_12709,N_12173,N_12356);
and U12710 (N_12710,N_12332,N_12397);
nand U12711 (N_12711,N_12062,N_12000);
nor U12712 (N_12712,N_12005,N_12052);
xor U12713 (N_12713,N_12255,N_12256);
and U12714 (N_12714,N_12165,N_12103);
nor U12715 (N_12715,N_12034,N_12237);
nor U12716 (N_12716,N_12074,N_12335);
nand U12717 (N_12717,N_12277,N_12116);
nand U12718 (N_12718,N_12010,N_12311);
and U12719 (N_12719,N_12349,N_12335);
and U12720 (N_12720,N_12203,N_12300);
and U12721 (N_12721,N_12384,N_12303);
and U12722 (N_12722,N_12281,N_12227);
nand U12723 (N_12723,N_12189,N_12183);
nand U12724 (N_12724,N_12150,N_12338);
or U12725 (N_12725,N_12328,N_12334);
nand U12726 (N_12726,N_12305,N_12397);
or U12727 (N_12727,N_12054,N_12022);
nor U12728 (N_12728,N_12301,N_12290);
nand U12729 (N_12729,N_12188,N_12298);
xor U12730 (N_12730,N_12166,N_12135);
and U12731 (N_12731,N_12285,N_12288);
or U12732 (N_12732,N_12088,N_12278);
nor U12733 (N_12733,N_12035,N_12141);
or U12734 (N_12734,N_12291,N_12027);
nand U12735 (N_12735,N_12083,N_12029);
nand U12736 (N_12736,N_12336,N_12188);
xor U12737 (N_12737,N_12109,N_12287);
or U12738 (N_12738,N_12038,N_12323);
nor U12739 (N_12739,N_12252,N_12170);
nand U12740 (N_12740,N_12009,N_12212);
xnor U12741 (N_12741,N_12283,N_12173);
and U12742 (N_12742,N_12330,N_12028);
and U12743 (N_12743,N_12206,N_12033);
xor U12744 (N_12744,N_12360,N_12181);
nand U12745 (N_12745,N_12118,N_12165);
and U12746 (N_12746,N_12252,N_12206);
and U12747 (N_12747,N_12340,N_12150);
or U12748 (N_12748,N_12348,N_12379);
nor U12749 (N_12749,N_12324,N_12343);
and U12750 (N_12750,N_12120,N_12122);
xnor U12751 (N_12751,N_12289,N_12334);
xnor U12752 (N_12752,N_12169,N_12384);
xnor U12753 (N_12753,N_12170,N_12245);
xor U12754 (N_12754,N_12242,N_12037);
xnor U12755 (N_12755,N_12321,N_12208);
or U12756 (N_12756,N_12174,N_12261);
xnor U12757 (N_12757,N_12334,N_12038);
nor U12758 (N_12758,N_12268,N_12348);
or U12759 (N_12759,N_12034,N_12349);
or U12760 (N_12760,N_12125,N_12181);
or U12761 (N_12761,N_12205,N_12272);
nor U12762 (N_12762,N_12381,N_12301);
nor U12763 (N_12763,N_12305,N_12123);
nand U12764 (N_12764,N_12296,N_12044);
xnor U12765 (N_12765,N_12146,N_12368);
xnor U12766 (N_12766,N_12380,N_12009);
or U12767 (N_12767,N_12273,N_12174);
xnor U12768 (N_12768,N_12354,N_12304);
or U12769 (N_12769,N_12052,N_12066);
nand U12770 (N_12770,N_12100,N_12179);
and U12771 (N_12771,N_12256,N_12026);
or U12772 (N_12772,N_12213,N_12072);
or U12773 (N_12773,N_12142,N_12195);
or U12774 (N_12774,N_12033,N_12181);
or U12775 (N_12775,N_12115,N_12195);
xor U12776 (N_12776,N_12160,N_12180);
xor U12777 (N_12777,N_12038,N_12352);
or U12778 (N_12778,N_12331,N_12231);
xnor U12779 (N_12779,N_12389,N_12252);
or U12780 (N_12780,N_12249,N_12257);
nor U12781 (N_12781,N_12163,N_12226);
nor U12782 (N_12782,N_12356,N_12004);
nor U12783 (N_12783,N_12348,N_12062);
and U12784 (N_12784,N_12100,N_12363);
or U12785 (N_12785,N_12370,N_12171);
nor U12786 (N_12786,N_12162,N_12008);
or U12787 (N_12787,N_12318,N_12223);
nand U12788 (N_12788,N_12388,N_12022);
nor U12789 (N_12789,N_12096,N_12155);
xor U12790 (N_12790,N_12282,N_12193);
or U12791 (N_12791,N_12161,N_12358);
nand U12792 (N_12792,N_12134,N_12288);
and U12793 (N_12793,N_12069,N_12113);
xor U12794 (N_12794,N_12218,N_12311);
or U12795 (N_12795,N_12353,N_12012);
and U12796 (N_12796,N_12051,N_12142);
or U12797 (N_12797,N_12095,N_12139);
nand U12798 (N_12798,N_12038,N_12283);
xnor U12799 (N_12799,N_12097,N_12053);
nor U12800 (N_12800,N_12717,N_12478);
nor U12801 (N_12801,N_12568,N_12546);
or U12802 (N_12802,N_12796,N_12547);
xor U12803 (N_12803,N_12778,N_12714);
and U12804 (N_12804,N_12465,N_12735);
nand U12805 (N_12805,N_12740,N_12578);
and U12806 (N_12806,N_12403,N_12701);
nand U12807 (N_12807,N_12769,N_12425);
xnor U12808 (N_12808,N_12510,N_12473);
xor U12809 (N_12809,N_12766,N_12628);
nor U12810 (N_12810,N_12548,N_12502);
and U12811 (N_12811,N_12542,N_12794);
and U12812 (N_12812,N_12655,N_12692);
xnor U12813 (N_12813,N_12448,N_12762);
or U12814 (N_12814,N_12688,N_12720);
nor U12815 (N_12815,N_12697,N_12506);
xnor U12816 (N_12816,N_12537,N_12683);
xor U12817 (N_12817,N_12677,N_12700);
xor U12818 (N_12818,N_12518,N_12445);
and U12819 (N_12819,N_12786,N_12704);
nor U12820 (N_12820,N_12507,N_12638);
nand U12821 (N_12821,N_12596,N_12637);
xor U12822 (N_12822,N_12587,N_12772);
or U12823 (N_12823,N_12513,N_12577);
nand U12824 (N_12824,N_12758,N_12503);
or U12825 (N_12825,N_12671,N_12779);
or U12826 (N_12826,N_12439,N_12645);
nand U12827 (N_12827,N_12440,N_12583);
and U12828 (N_12828,N_12595,N_12526);
or U12829 (N_12829,N_12742,N_12715);
xnor U12830 (N_12830,N_12410,N_12543);
or U12831 (N_12831,N_12711,N_12636);
nand U12832 (N_12832,N_12625,N_12746);
and U12833 (N_12833,N_12680,N_12748);
xor U12834 (N_12834,N_12593,N_12451);
xnor U12835 (N_12835,N_12405,N_12505);
nand U12836 (N_12836,N_12571,N_12592);
nand U12837 (N_12837,N_12570,N_12629);
xnor U12838 (N_12838,N_12653,N_12633);
nor U12839 (N_12839,N_12659,N_12552);
nor U12840 (N_12840,N_12749,N_12544);
and U12841 (N_12841,N_12418,N_12420);
nand U12842 (N_12842,N_12444,N_12512);
nor U12843 (N_12843,N_12624,N_12459);
or U12844 (N_12844,N_12608,N_12569);
nand U12845 (N_12845,N_12446,N_12453);
and U12846 (N_12846,N_12771,N_12631);
or U12847 (N_12847,N_12400,N_12793);
nand U12848 (N_12848,N_12763,N_12666);
xnor U12849 (N_12849,N_12588,N_12450);
nand U12850 (N_12850,N_12558,N_12675);
nand U12851 (N_12851,N_12780,N_12469);
or U12852 (N_12852,N_12611,N_12422);
nand U12853 (N_12853,N_12651,N_12407);
xor U12854 (N_12854,N_12457,N_12464);
xor U12855 (N_12855,N_12643,N_12534);
or U12856 (N_12856,N_12718,N_12733);
nand U12857 (N_12857,N_12663,N_12723);
and U12858 (N_12858,N_12460,N_12566);
nand U12859 (N_12859,N_12560,N_12454);
or U12860 (N_12860,N_12756,N_12712);
and U12861 (N_12861,N_12589,N_12797);
nand U12862 (N_12862,N_12564,N_12644);
xnor U12863 (N_12863,N_12549,N_12461);
nand U12864 (N_12864,N_12412,N_12795);
or U12865 (N_12865,N_12606,N_12646);
and U12866 (N_12866,N_12437,N_12759);
xnor U12867 (N_12867,N_12743,N_12480);
and U12868 (N_12868,N_12575,N_12408);
nor U12869 (N_12869,N_12556,N_12703);
or U12870 (N_12870,N_12545,N_12533);
xnor U12871 (N_12871,N_12495,N_12431);
or U12872 (N_12872,N_12672,N_12550);
and U12873 (N_12873,N_12661,N_12551);
and U12874 (N_12874,N_12471,N_12541);
nand U12875 (N_12875,N_12498,N_12630);
and U12876 (N_12876,N_12785,N_12515);
or U12877 (N_12877,N_12652,N_12486);
xnor U12878 (N_12878,N_12438,N_12623);
and U12879 (N_12879,N_12790,N_12657);
or U12880 (N_12880,N_12530,N_12484);
or U12881 (N_12881,N_12674,N_12741);
xnor U12882 (N_12882,N_12591,N_12788);
nor U12883 (N_12883,N_12435,N_12580);
nand U12884 (N_12884,N_12719,N_12601);
and U12885 (N_12885,N_12521,N_12658);
or U12886 (N_12886,N_12693,N_12501);
nor U12887 (N_12887,N_12477,N_12737);
and U12888 (N_12888,N_12557,N_12713);
nand U12889 (N_12889,N_12555,N_12690);
nand U12890 (N_12890,N_12782,N_12561);
xnor U12891 (N_12891,N_12667,N_12662);
and U12892 (N_12892,N_12567,N_12724);
and U12893 (N_12893,N_12668,N_12642);
and U12894 (N_12894,N_12509,N_12791);
or U12895 (N_12895,N_12789,N_12590);
and U12896 (N_12896,N_12770,N_12524);
xor U12897 (N_12897,N_12582,N_12679);
nand U12898 (N_12898,N_12572,N_12436);
and U12899 (N_12899,N_12665,N_12494);
or U12900 (N_12900,N_12585,N_12433);
and U12901 (N_12901,N_12520,N_12691);
nand U12902 (N_12902,N_12532,N_12670);
nand U12903 (N_12903,N_12783,N_12508);
nand U12904 (N_12904,N_12784,N_12415);
xnor U12905 (N_12905,N_12777,N_12621);
nor U12906 (N_12906,N_12517,N_12626);
and U12907 (N_12907,N_12710,N_12490);
nor U12908 (N_12908,N_12727,N_12765);
nor U12909 (N_12909,N_12615,N_12491);
xor U12910 (N_12910,N_12401,N_12726);
and U12911 (N_12911,N_12604,N_12755);
xnor U12912 (N_12912,N_12522,N_12619);
or U12913 (N_12913,N_12443,N_12773);
nor U12914 (N_12914,N_12747,N_12722);
and U12915 (N_12915,N_12634,N_12540);
nor U12916 (N_12916,N_12760,N_12479);
nor U12917 (N_12917,N_12599,N_12620);
and U12918 (N_12918,N_12493,N_12482);
nor U12919 (N_12919,N_12409,N_12768);
nand U12920 (N_12920,N_12622,N_12475);
nand U12921 (N_12921,N_12514,N_12685);
and U12922 (N_12922,N_12707,N_12417);
nand U12923 (N_12923,N_12496,N_12776);
or U12924 (N_12924,N_12456,N_12617);
or U12925 (N_12925,N_12528,N_12488);
nand U12926 (N_12926,N_12654,N_12468);
nor U12927 (N_12927,N_12535,N_12581);
xnor U12928 (N_12928,N_12676,N_12799);
or U12929 (N_12929,N_12467,N_12753);
or U12930 (N_12930,N_12492,N_12739);
nand U12931 (N_12931,N_12481,N_12734);
nand U12932 (N_12932,N_12648,N_12519);
or U12933 (N_12933,N_12413,N_12664);
and U12934 (N_12934,N_12761,N_12728);
and U12935 (N_12935,N_12442,N_12466);
or U12936 (N_12936,N_12736,N_12757);
nor U12937 (N_12937,N_12787,N_12529);
or U12938 (N_12938,N_12750,N_12455);
and U12939 (N_12939,N_12428,N_12774);
nand U12940 (N_12940,N_12602,N_12419);
and U12941 (N_12941,N_12536,N_12525);
and U12942 (N_12942,N_12798,N_12612);
and U12943 (N_12943,N_12603,N_12434);
or U12944 (N_12944,N_12694,N_12605);
nor U12945 (N_12945,N_12708,N_12754);
and U12946 (N_12946,N_12476,N_12553);
nor U12947 (N_12947,N_12452,N_12686);
or U12948 (N_12948,N_12424,N_12538);
nor U12949 (N_12949,N_12689,N_12632);
nand U12950 (N_12950,N_12745,N_12576);
or U12951 (N_12951,N_12660,N_12504);
nand U12952 (N_12952,N_12427,N_12565);
xor U12953 (N_12953,N_12695,N_12579);
nand U12954 (N_12954,N_12573,N_12554);
and U12955 (N_12955,N_12709,N_12406);
and U12956 (N_12956,N_12649,N_12411);
or U12957 (N_12957,N_12489,N_12681);
nand U12958 (N_12958,N_12559,N_12721);
xnor U12959 (N_12959,N_12656,N_12775);
and U12960 (N_12960,N_12430,N_12716);
nand U12961 (N_12961,N_12627,N_12635);
xor U12962 (N_12962,N_12449,N_12730);
and U12963 (N_12963,N_12426,N_12421);
nor U12964 (N_12964,N_12767,N_12563);
nand U12965 (N_12965,N_12499,N_12462);
and U12966 (N_12966,N_12527,N_12640);
and U12967 (N_12967,N_12669,N_12600);
xor U12968 (N_12968,N_12539,N_12609);
nor U12969 (N_12969,N_12447,N_12497);
or U12970 (N_12970,N_12607,N_12511);
nand U12971 (N_12971,N_12682,N_12610);
nand U12972 (N_12972,N_12641,N_12729);
and U12973 (N_12973,N_12402,N_12485);
nor U12974 (N_12974,N_12441,N_12706);
xnor U12975 (N_12975,N_12594,N_12687);
nand U12976 (N_12976,N_12423,N_12616);
nor U12977 (N_12977,N_12562,N_12751);
and U12978 (N_12978,N_12792,N_12500);
xnor U12979 (N_12979,N_12699,N_12574);
and U12980 (N_12980,N_12598,N_12764);
and U12981 (N_12981,N_12470,N_12732);
nand U12982 (N_12982,N_12584,N_12458);
xor U12983 (N_12983,N_12516,N_12487);
or U12984 (N_12984,N_12472,N_12725);
nand U12985 (N_12985,N_12586,N_12738);
or U12986 (N_12986,N_12702,N_12696);
nor U12987 (N_12987,N_12614,N_12429);
nand U12988 (N_12988,N_12781,N_12432);
nor U12989 (N_12989,N_12744,N_12416);
xnor U12990 (N_12990,N_12731,N_12414);
nor U12991 (N_12991,N_12673,N_12705);
xnor U12992 (N_12992,N_12678,N_12639);
and U12993 (N_12993,N_12647,N_12597);
nor U12994 (N_12994,N_12531,N_12650);
and U12995 (N_12995,N_12463,N_12613);
nand U12996 (N_12996,N_12483,N_12618);
nor U12997 (N_12997,N_12523,N_12404);
xnor U12998 (N_12998,N_12698,N_12684);
nor U12999 (N_12999,N_12474,N_12752);
xor U13000 (N_13000,N_12507,N_12473);
nor U13001 (N_13001,N_12639,N_12572);
or U13002 (N_13002,N_12405,N_12765);
and U13003 (N_13003,N_12551,N_12738);
nand U13004 (N_13004,N_12575,N_12506);
or U13005 (N_13005,N_12574,N_12596);
and U13006 (N_13006,N_12788,N_12535);
or U13007 (N_13007,N_12566,N_12478);
nor U13008 (N_13008,N_12767,N_12766);
or U13009 (N_13009,N_12540,N_12715);
nand U13010 (N_13010,N_12686,N_12671);
nand U13011 (N_13011,N_12476,N_12767);
nand U13012 (N_13012,N_12677,N_12713);
and U13013 (N_13013,N_12408,N_12620);
nand U13014 (N_13014,N_12540,N_12640);
or U13015 (N_13015,N_12776,N_12507);
nor U13016 (N_13016,N_12544,N_12425);
xnor U13017 (N_13017,N_12447,N_12519);
nand U13018 (N_13018,N_12402,N_12798);
nor U13019 (N_13019,N_12450,N_12665);
nand U13020 (N_13020,N_12588,N_12755);
and U13021 (N_13021,N_12490,N_12438);
xnor U13022 (N_13022,N_12526,N_12705);
and U13023 (N_13023,N_12747,N_12712);
nand U13024 (N_13024,N_12418,N_12477);
xor U13025 (N_13025,N_12470,N_12653);
and U13026 (N_13026,N_12423,N_12654);
or U13027 (N_13027,N_12617,N_12503);
and U13028 (N_13028,N_12766,N_12454);
nor U13029 (N_13029,N_12535,N_12612);
nor U13030 (N_13030,N_12580,N_12613);
and U13031 (N_13031,N_12461,N_12605);
nor U13032 (N_13032,N_12486,N_12602);
or U13033 (N_13033,N_12785,N_12685);
and U13034 (N_13034,N_12429,N_12688);
xor U13035 (N_13035,N_12719,N_12797);
and U13036 (N_13036,N_12776,N_12760);
or U13037 (N_13037,N_12741,N_12506);
nor U13038 (N_13038,N_12421,N_12516);
xnor U13039 (N_13039,N_12776,N_12616);
nand U13040 (N_13040,N_12486,N_12785);
xor U13041 (N_13041,N_12777,N_12467);
or U13042 (N_13042,N_12437,N_12499);
nand U13043 (N_13043,N_12587,N_12668);
nand U13044 (N_13044,N_12610,N_12757);
xnor U13045 (N_13045,N_12571,N_12581);
xnor U13046 (N_13046,N_12502,N_12421);
or U13047 (N_13047,N_12432,N_12641);
and U13048 (N_13048,N_12528,N_12415);
nor U13049 (N_13049,N_12403,N_12577);
xor U13050 (N_13050,N_12667,N_12441);
or U13051 (N_13051,N_12403,N_12418);
xnor U13052 (N_13052,N_12677,N_12705);
or U13053 (N_13053,N_12476,N_12558);
xnor U13054 (N_13054,N_12758,N_12782);
nand U13055 (N_13055,N_12581,N_12454);
xor U13056 (N_13056,N_12415,N_12711);
nand U13057 (N_13057,N_12628,N_12494);
nand U13058 (N_13058,N_12540,N_12793);
or U13059 (N_13059,N_12551,N_12714);
or U13060 (N_13060,N_12635,N_12746);
nor U13061 (N_13061,N_12624,N_12520);
nand U13062 (N_13062,N_12685,N_12766);
or U13063 (N_13063,N_12567,N_12421);
and U13064 (N_13064,N_12481,N_12533);
or U13065 (N_13065,N_12752,N_12740);
nand U13066 (N_13066,N_12712,N_12779);
nand U13067 (N_13067,N_12479,N_12775);
or U13068 (N_13068,N_12737,N_12460);
and U13069 (N_13069,N_12780,N_12658);
and U13070 (N_13070,N_12508,N_12547);
nand U13071 (N_13071,N_12588,N_12638);
nor U13072 (N_13072,N_12419,N_12675);
and U13073 (N_13073,N_12493,N_12489);
or U13074 (N_13074,N_12590,N_12464);
xnor U13075 (N_13075,N_12725,N_12431);
nand U13076 (N_13076,N_12470,N_12589);
and U13077 (N_13077,N_12483,N_12614);
and U13078 (N_13078,N_12732,N_12401);
nor U13079 (N_13079,N_12764,N_12757);
and U13080 (N_13080,N_12682,N_12608);
or U13081 (N_13081,N_12423,N_12434);
nand U13082 (N_13082,N_12509,N_12433);
nor U13083 (N_13083,N_12478,N_12594);
xnor U13084 (N_13084,N_12714,N_12438);
nand U13085 (N_13085,N_12556,N_12715);
nand U13086 (N_13086,N_12720,N_12484);
nor U13087 (N_13087,N_12491,N_12531);
and U13088 (N_13088,N_12566,N_12570);
xnor U13089 (N_13089,N_12631,N_12405);
xor U13090 (N_13090,N_12488,N_12435);
xor U13091 (N_13091,N_12538,N_12784);
xor U13092 (N_13092,N_12512,N_12695);
nand U13093 (N_13093,N_12543,N_12777);
or U13094 (N_13094,N_12636,N_12752);
and U13095 (N_13095,N_12572,N_12746);
nand U13096 (N_13096,N_12519,N_12643);
and U13097 (N_13097,N_12755,N_12444);
nor U13098 (N_13098,N_12600,N_12687);
and U13099 (N_13099,N_12677,N_12739);
nor U13100 (N_13100,N_12793,N_12476);
or U13101 (N_13101,N_12467,N_12785);
xnor U13102 (N_13102,N_12535,N_12532);
nand U13103 (N_13103,N_12754,N_12441);
xnor U13104 (N_13104,N_12753,N_12584);
and U13105 (N_13105,N_12508,N_12777);
nor U13106 (N_13106,N_12633,N_12494);
nor U13107 (N_13107,N_12465,N_12497);
nor U13108 (N_13108,N_12426,N_12719);
or U13109 (N_13109,N_12422,N_12616);
and U13110 (N_13110,N_12474,N_12473);
xor U13111 (N_13111,N_12640,N_12632);
or U13112 (N_13112,N_12539,N_12579);
xor U13113 (N_13113,N_12682,N_12607);
xnor U13114 (N_13114,N_12456,N_12532);
nand U13115 (N_13115,N_12644,N_12400);
nand U13116 (N_13116,N_12661,N_12427);
and U13117 (N_13117,N_12573,N_12799);
and U13118 (N_13118,N_12512,N_12671);
nand U13119 (N_13119,N_12772,N_12749);
and U13120 (N_13120,N_12436,N_12603);
nor U13121 (N_13121,N_12788,N_12554);
nand U13122 (N_13122,N_12740,N_12566);
or U13123 (N_13123,N_12639,N_12603);
xor U13124 (N_13124,N_12635,N_12789);
xnor U13125 (N_13125,N_12490,N_12759);
nor U13126 (N_13126,N_12766,N_12470);
nor U13127 (N_13127,N_12506,N_12618);
xnor U13128 (N_13128,N_12534,N_12786);
xor U13129 (N_13129,N_12610,N_12678);
nand U13130 (N_13130,N_12552,N_12437);
nor U13131 (N_13131,N_12495,N_12536);
nand U13132 (N_13132,N_12749,N_12709);
nor U13133 (N_13133,N_12484,N_12687);
nor U13134 (N_13134,N_12760,N_12651);
nor U13135 (N_13135,N_12627,N_12499);
and U13136 (N_13136,N_12678,N_12485);
or U13137 (N_13137,N_12757,N_12754);
nor U13138 (N_13138,N_12488,N_12534);
or U13139 (N_13139,N_12671,N_12792);
nor U13140 (N_13140,N_12584,N_12445);
xnor U13141 (N_13141,N_12690,N_12715);
and U13142 (N_13142,N_12738,N_12423);
nand U13143 (N_13143,N_12575,N_12503);
nor U13144 (N_13144,N_12636,N_12784);
nor U13145 (N_13145,N_12501,N_12660);
or U13146 (N_13146,N_12623,N_12463);
or U13147 (N_13147,N_12657,N_12514);
xnor U13148 (N_13148,N_12668,N_12446);
nand U13149 (N_13149,N_12741,N_12726);
and U13150 (N_13150,N_12416,N_12763);
or U13151 (N_13151,N_12577,N_12706);
nor U13152 (N_13152,N_12505,N_12755);
and U13153 (N_13153,N_12611,N_12769);
and U13154 (N_13154,N_12658,N_12727);
nor U13155 (N_13155,N_12520,N_12477);
or U13156 (N_13156,N_12531,N_12749);
and U13157 (N_13157,N_12678,N_12747);
xor U13158 (N_13158,N_12490,N_12631);
and U13159 (N_13159,N_12504,N_12667);
xnor U13160 (N_13160,N_12505,N_12442);
xor U13161 (N_13161,N_12707,N_12621);
and U13162 (N_13162,N_12636,N_12430);
and U13163 (N_13163,N_12558,N_12680);
nand U13164 (N_13164,N_12789,N_12494);
nand U13165 (N_13165,N_12742,N_12489);
nor U13166 (N_13166,N_12747,N_12775);
xnor U13167 (N_13167,N_12769,N_12448);
or U13168 (N_13168,N_12469,N_12671);
xnor U13169 (N_13169,N_12438,N_12738);
nand U13170 (N_13170,N_12714,N_12474);
and U13171 (N_13171,N_12452,N_12735);
nand U13172 (N_13172,N_12462,N_12524);
nor U13173 (N_13173,N_12434,N_12508);
xnor U13174 (N_13174,N_12434,N_12504);
nor U13175 (N_13175,N_12670,N_12561);
or U13176 (N_13176,N_12518,N_12709);
nand U13177 (N_13177,N_12458,N_12493);
and U13178 (N_13178,N_12514,N_12643);
nor U13179 (N_13179,N_12415,N_12531);
and U13180 (N_13180,N_12655,N_12773);
nor U13181 (N_13181,N_12761,N_12529);
or U13182 (N_13182,N_12464,N_12553);
and U13183 (N_13183,N_12795,N_12775);
nand U13184 (N_13184,N_12638,N_12586);
or U13185 (N_13185,N_12584,N_12621);
or U13186 (N_13186,N_12767,N_12575);
and U13187 (N_13187,N_12538,N_12676);
nand U13188 (N_13188,N_12623,N_12736);
nor U13189 (N_13189,N_12675,N_12784);
nor U13190 (N_13190,N_12544,N_12434);
or U13191 (N_13191,N_12607,N_12681);
and U13192 (N_13192,N_12453,N_12763);
or U13193 (N_13193,N_12736,N_12553);
nand U13194 (N_13194,N_12725,N_12628);
nand U13195 (N_13195,N_12750,N_12679);
nand U13196 (N_13196,N_12610,N_12724);
and U13197 (N_13197,N_12621,N_12556);
and U13198 (N_13198,N_12566,N_12769);
and U13199 (N_13199,N_12567,N_12409);
and U13200 (N_13200,N_12962,N_13024);
nor U13201 (N_13201,N_13062,N_12911);
or U13202 (N_13202,N_13102,N_13058);
or U13203 (N_13203,N_13159,N_13185);
nor U13204 (N_13204,N_12864,N_12814);
xnor U13205 (N_13205,N_12832,N_12822);
or U13206 (N_13206,N_12921,N_13028);
or U13207 (N_13207,N_13035,N_12840);
xnor U13208 (N_13208,N_13195,N_13050);
and U13209 (N_13209,N_12802,N_12837);
nor U13210 (N_13210,N_12983,N_13044);
nand U13211 (N_13211,N_13116,N_13042);
xnor U13212 (N_13212,N_12823,N_13096);
xor U13213 (N_13213,N_13049,N_13070);
xor U13214 (N_13214,N_12855,N_12844);
nand U13215 (N_13215,N_12945,N_12841);
nor U13216 (N_13216,N_12949,N_13183);
or U13217 (N_13217,N_12904,N_12984);
or U13218 (N_13218,N_13182,N_13043);
and U13219 (N_13219,N_12878,N_13147);
nand U13220 (N_13220,N_12815,N_12957);
and U13221 (N_13221,N_12849,N_12929);
xnor U13222 (N_13222,N_13064,N_13073);
or U13223 (N_13223,N_13138,N_12835);
xnor U13224 (N_13224,N_12915,N_13016);
nand U13225 (N_13225,N_12946,N_12803);
and U13226 (N_13226,N_12991,N_12971);
nor U13227 (N_13227,N_13004,N_12977);
and U13228 (N_13228,N_12843,N_13023);
xnor U13229 (N_13229,N_12948,N_12910);
xnor U13230 (N_13230,N_12887,N_12830);
nand U13231 (N_13231,N_13128,N_13082);
or U13232 (N_13232,N_12892,N_12933);
nand U13233 (N_13233,N_12839,N_13099);
xnor U13234 (N_13234,N_12992,N_12975);
nand U13235 (N_13235,N_12817,N_13157);
nand U13236 (N_13236,N_12859,N_12987);
or U13237 (N_13237,N_12931,N_12965);
nor U13238 (N_13238,N_13119,N_13075);
nor U13239 (N_13239,N_12934,N_12954);
or U13240 (N_13240,N_13091,N_13100);
or U13241 (N_13241,N_13153,N_13010);
and U13242 (N_13242,N_12842,N_13041);
nand U13243 (N_13243,N_12979,N_13008);
nand U13244 (N_13244,N_13162,N_12923);
and U13245 (N_13245,N_12937,N_12994);
nand U13246 (N_13246,N_13191,N_13065);
xnor U13247 (N_13247,N_13142,N_13045);
and U13248 (N_13248,N_13000,N_13127);
xnor U13249 (N_13249,N_13144,N_13137);
nand U13250 (N_13250,N_13103,N_12893);
or U13251 (N_13251,N_13177,N_13090);
or U13252 (N_13252,N_12908,N_13145);
or U13253 (N_13253,N_12953,N_12821);
nand U13254 (N_13254,N_13033,N_12881);
or U13255 (N_13255,N_13110,N_12877);
nor U13256 (N_13256,N_12860,N_13029);
xor U13257 (N_13257,N_13052,N_12996);
xor U13258 (N_13258,N_13188,N_12826);
nor U13259 (N_13259,N_13037,N_12919);
nand U13260 (N_13260,N_13131,N_12970);
nand U13261 (N_13261,N_13186,N_12820);
or U13262 (N_13262,N_12875,N_13164);
xor U13263 (N_13263,N_13166,N_13022);
and U13264 (N_13264,N_13151,N_12952);
or U13265 (N_13265,N_12813,N_13093);
and U13266 (N_13266,N_12905,N_13150);
or U13267 (N_13267,N_13122,N_13072);
and U13268 (N_13268,N_13101,N_13179);
nor U13269 (N_13269,N_12907,N_13086);
and U13270 (N_13270,N_13002,N_12891);
xnor U13271 (N_13271,N_13154,N_13094);
and U13272 (N_13272,N_13059,N_13158);
xnor U13273 (N_13273,N_13114,N_13098);
or U13274 (N_13274,N_13143,N_13141);
xor U13275 (N_13275,N_12944,N_12871);
or U13276 (N_13276,N_13178,N_12872);
or U13277 (N_13277,N_12914,N_13057);
xnor U13278 (N_13278,N_12967,N_13140);
nor U13279 (N_13279,N_13174,N_12913);
or U13280 (N_13280,N_13014,N_12870);
nand U13281 (N_13281,N_12938,N_13197);
and U13282 (N_13282,N_12828,N_12988);
xnor U13283 (N_13283,N_13148,N_12998);
nand U13284 (N_13284,N_13112,N_12909);
nand U13285 (N_13285,N_13163,N_13189);
nand U13286 (N_13286,N_12856,N_12883);
and U13287 (N_13287,N_12951,N_12978);
or U13288 (N_13288,N_12972,N_13034);
nand U13289 (N_13289,N_13048,N_12867);
and U13290 (N_13290,N_13001,N_13085);
nand U13291 (N_13291,N_13165,N_13107);
nor U13292 (N_13292,N_12825,N_12894);
and U13293 (N_13293,N_12916,N_13026);
nor U13294 (N_13294,N_12993,N_13095);
xnor U13295 (N_13295,N_13192,N_12981);
nor U13296 (N_13296,N_13190,N_12806);
xnor U13297 (N_13297,N_13184,N_13152);
nand U13298 (N_13298,N_12906,N_12804);
nand U13299 (N_13299,N_13079,N_12846);
nor U13300 (N_13300,N_12874,N_12897);
nand U13301 (N_13301,N_12941,N_12833);
nor U13302 (N_13302,N_12973,N_12819);
or U13303 (N_13303,N_13092,N_13125);
nand U13304 (N_13304,N_12927,N_12964);
xnor U13305 (N_13305,N_13194,N_13134);
and U13306 (N_13306,N_13061,N_13007);
xnor U13307 (N_13307,N_13129,N_12958);
and U13308 (N_13308,N_13169,N_13139);
xor U13309 (N_13309,N_12903,N_12918);
nor U13310 (N_13310,N_12924,N_12940);
or U13311 (N_13311,N_12876,N_12880);
nor U13312 (N_13312,N_13066,N_12807);
nor U13313 (N_13313,N_12836,N_12898);
nand U13314 (N_13314,N_12800,N_13080);
and U13315 (N_13315,N_13135,N_12812);
and U13316 (N_13316,N_12805,N_13077);
and U13317 (N_13317,N_12926,N_13132);
and U13318 (N_13318,N_12816,N_13051);
nor U13319 (N_13319,N_13104,N_12861);
nor U13320 (N_13320,N_13060,N_13088);
xor U13321 (N_13321,N_13167,N_13017);
nand U13322 (N_13322,N_13047,N_13133);
nor U13323 (N_13323,N_12869,N_13046);
xor U13324 (N_13324,N_12935,N_12968);
and U13325 (N_13325,N_13021,N_12969);
nor U13326 (N_13326,N_12884,N_12801);
nor U13327 (N_13327,N_12922,N_12809);
or U13328 (N_13328,N_13121,N_13180);
and U13329 (N_13329,N_13020,N_13068);
nor U13330 (N_13330,N_13123,N_12834);
nand U13331 (N_13331,N_12990,N_13146);
nand U13332 (N_13332,N_12902,N_13032);
nor U13333 (N_13333,N_13013,N_12857);
nand U13334 (N_13334,N_13170,N_13196);
nand U13335 (N_13335,N_13175,N_12966);
nor U13336 (N_13336,N_12879,N_13011);
or U13337 (N_13337,N_13069,N_13130);
or U13338 (N_13338,N_12930,N_13009);
nand U13339 (N_13339,N_13063,N_12885);
nor U13340 (N_13340,N_12999,N_13089);
nor U13341 (N_13341,N_12963,N_13173);
and U13342 (N_13342,N_12827,N_12852);
xor U13343 (N_13343,N_12989,N_12811);
xor U13344 (N_13344,N_13108,N_13040);
and U13345 (N_13345,N_13081,N_12895);
nand U13346 (N_13346,N_13067,N_13161);
nor U13347 (N_13347,N_12882,N_13055);
nor U13348 (N_13348,N_13076,N_12955);
or U13349 (N_13349,N_13083,N_12808);
nand U13350 (N_13350,N_12818,N_13160);
or U13351 (N_13351,N_13198,N_13181);
or U13352 (N_13352,N_13199,N_12942);
or U13353 (N_13353,N_13120,N_13176);
xnor U13354 (N_13354,N_12863,N_12824);
nand U13355 (N_13355,N_13136,N_12986);
nand U13356 (N_13356,N_13106,N_13087);
or U13357 (N_13357,N_12980,N_12847);
or U13358 (N_13358,N_13097,N_13018);
nand U13359 (N_13359,N_12810,N_12932);
and U13360 (N_13360,N_13031,N_13019);
xnor U13361 (N_13361,N_13027,N_12982);
xnor U13362 (N_13362,N_13156,N_12939);
or U13363 (N_13363,N_13030,N_12959);
or U13364 (N_13364,N_13071,N_12831);
xnor U13365 (N_13365,N_12976,N_12960);
nand U13366 (N_13366,N_12853,N_12865);
nor U13367 (N_13367,N_12943,N_12889);
or U13368 (N_13368,N_13056,N_12886);
nor U13369 (N_13369,N_13039,N_12888);
or U13370 (N_13370,N_12985,N_12866);
and U13371 (N_13371,N_12928,N_13078);
and U13372 (N_13372,N_13038,N_13025);
or U13373 (N_13373,N_12890,N_13171);
nand U13374 (N_13374,N_13054,N_12995);
or U13375 (N_13375,N_12900,N_12845);
nor U13376 (N_13376,N_12961,N_13005);
and U13377 (N_13377,N_12850,N_13118);
xnor U13378 (N_13378,N_13074,N_13149);
and U13379 (N_13379,N_12854,N_12974);
nor U13380 (N_13380,N_12899,N_12947);
nand U13381 (N_13381,N_12862,N_13172);
xor U13382 (N_13382,N_13168,N_13113);
and U13383 (N_13383,N_12848,N_12997);
nand U13384 (N_13384,N_13084,N_13053);
xor U13385 (N_13385,N_13126,N_12917);
nor U13386 (N_13386,N_13117,N_12838);
xor U13387 (N_13387,N_12925,N_13111);
xor U13388 (N_13388,N_12956,N_13187);
or U13389 (N_13389,N_13006,N_12868);
nand U13390 (N_13390,N_13012,N_13036);
nand U13391 (N_13391,N_13015,N_13155);
nand U13392 (N_13392,N_13115,N_13109);
xor U13393 (N_13393,N_12858,N_12950);
or U13394 (N_13394,N_12851,N_12936);
or U13395 (N_13395,N_12901,N_12829);
xor U13396 (N_13396,N_12920,N_13003);
and U13397 (N_13397,N_12912,N_12896);
nand U13398 (N_13398,N_13105,N_12873);
nand U13399 (N_13399,N_13124,N_13193);
and U13400 (N_13400,N_13105,N_12983);
nor U13401 (N_13401,N_12981,N_12826);
nand U13402 (N_13402,N_13187,N_13021);
nand U13403 (N_13403,N_13042,N_12883);
xor U13404 (N_13404,N_12955,N_12951);
nand U13405 (N_13405,N_12884,N_13018);
or U13406 (N_13406,N_12993,N_12902);
or U13407 (N_13407,N_12980,N_13157);
nand U13408 (N_13408,N_13030,N_12956);
or U13409 (N_13409,N_13093,N_12882);
nor U13410 (N_13410,N_12888,N_12983);
and U13411 (N_13411,N_13146,N_12814);
xor U13412 (N_13412,N_12833,N_12800);
xnor U13413 (N_13413,N_13050,N_13005);
xor U13414 (N_13414,N_12909,N_13069);
and U13415 (N_13415,N_13128,N_13086);
or U13416 (N_13416,N_13101,N_12811);
nor U13417 (N_13417,N_13093,N_12836);
nand U13418 (N_13418,N_13150,N_13026);
or U13419 (N_13419,N_12967,N_13160);
nand U13420 (N_13420,N_13044,N_12810);
nand U13421 (N_13421,N_13119,N_12825);
and U13422 (N_13422,N_12876,N_13183);
or U13423 (N_13423,N_12839,N_12849);
or U13424 (N_13424,N_12816,N_13063);
and U13425 (N_13425,N_13079,N_13173);
or U13426 (N_13426,N_13130,N_13128);
and U13427 (N_13427,N_12829,N_13123);
and U13428 (N_13428,N_13018,N_13091);
xor U13429 (N_13429,N_13146,N_13062);
nand U13430 (N_13430,N_12989,N_12940);
xor U13431 (N_13431,N_12826,N_12877);
nand U13432 (N_13432,N_12886,N_13033);
or U13433 (N_13433,N_12956,N_13166);
nand U13434 (N_13434,N_13168,N_13040);
xnor U13435 (N_13435,N_13025,N_12814);
xor U13436 (N_13436,N_13136,N_13098);
and U13437 (N_13437,N_13060,N_13164);
or U13438 (N_13438,N_12800,N_13064);
xnor U13439 (N_13439,N_13027,N_13190);
and U13440 (N_13440,N_12932,N_12961);
or U13441 (N_13441,N_13192,N_13044);
nand U13442 (N_13442,N_12895,N_12817);
or U13443 (N_13443,N_13180,N_13066);
or U13444 (N_13444,N_13141,N_12850);
xnor U13445 (N_13445,N_13161,N_12830);
and U13446 (N_13446,N_13031,N_13000);
nand U13447 (N_13447,N_13056,N_13112);
and U13448 (N_13448,N_13042,N_12969);
nand U13449 (N_13449,N_13075,N_13032);
or U13450 (N_13450,N_12805,N_12902);
nor U13451 (N_13451,N_12896,N_12882);
xor U13452 (N_13452,N_12851,N_13140);
xnor U13453 (N_13453,N_13165,N_13108);
or U13454 (N_13454,N_13017,N_13094);
and U13455 (N_13455,N_12975,N_13087);
nor U13456 (N_13456,N_12977,N_12838);
nor U13457 (N_13457,N_12926,N_12956);
nand U13458 (N_13458,N_13090,N_12847);
or U13459 (N_13459,N_12995,N_13066);
xor U13460 (N_13460,N_12929,N_13039);
and U13461 (N_13461,N_12874,N_13166);
nor U13462 (N_13462,N_12991,N_13126);
and U13463 (N_13463,N_13072,N_12881);
or U13464 (N_13464,N_13131,N_13003);
nor U13465 (N_13465,N_12910,N_13148);
xor U13466 (N_13466,N_13191,N_13171);
or U13467 (N_13467,N_13163,N_13030);
nand U13468 (N_13468,N_12989,N_12897);
and U13469 (N_13469,N_12884,N_13158);
nand U13470 (N_13470,N_13000,N_13078);
nor U13471 (N_13471,N_12961,N_12805);
and U13472 (N_13472,N_13063,N_13144);
nor U13473 (N_13473,N_12832,N_12859);
or U13474 (N_13474,N_13178,N_13132);
and U13475 (N_13475,N_13055,N_12997);
xor U13476 (N_13476,N_12997,N_12836);
nand U13477 (N_13477,N_13089,N_13051);
nor U13478 (N_13478,N_12989,N_13136);
or U13479 (N_13479,N_13064,N_12969);
or U13480 (N_13480,N_13049,N_13147);
xor U13481 (N_13481,N_12936,N_12878);
xnor U13482 (N_13482,N_13120,N_12943);
and U13483 (N_13483,N_13041,N_12937);
nand U13484 (N_13484,N_13144,N_12873);
nand U13485 (N_13485,N_13066,N_12873);
nor U13486 (N_13486,N_12905,N_13115);
nand U13487 (N_13487,N_12854,N_13153);
and U13488 (N_13488,N_13123,N_12867);
or U13489 (N_13489,N_12874,N_13011);
or U13490 (N_13490,N_13177,N_12990);
xnor U13491 (N_13491,N_12895,N_13057);
nor U13492 (N_13492,N_12967,N_12860);
xor U13493 (N_13493,N_12962,N_13137);
nand U13494 (N_13494,N_12828,N_12982);
nor U13495 (N_13495,N_12986,N_13057);
nor U13496 (N_13496,N_12933,N_12849);
nand U13497 (N_13497,N_13063,N_13012);
or U13498 (N_13498,N_12959,N_13143);
or U13499 (N_13499,N_12823,N_13047);
or U13500 (N_13500,N_12871,N_13094);
or U13501 (N_13501,N_12847,N_12875);
and U13502 (N_13502,N_13053,N_12991);
nor U13503 (N_13503,N_12922,N_12986);
nand U13504 (N_13504,N_13145,N_12859);
and U13505 (N_13505,N_13121,N_12975);
and U13506 (N_13506,N_12817,N_12873);
xor U13507 (N_13507,N_13111,N_12990);
or U13508 (N_13508,N_12807,N_12938);
nor U13509 (N_13509,N_12840,N_12936);
or U13510 (N_13510,N_13062,N_12895);
nand U13511 (N_13511,N_12954,N_12841);
and U13512 (N_13512,N_12875,N_13119);
nand U13513 (N_13513,N_12972,N_12954);
nand U13514 (N_13514,N_12866,N_12897);
and U13515 (N_13515,N_12884,N_12975);
nand U13516 (N_13516,N_13059,N_13195);
nand U13517 (N_13517,N_13166,N_13079);
and U13518 (N_13518,N_13193,N_13050);
or U13519 (N_13519,N_13001,N_13151);
and U13520 (N_13520,N_13171,N_12968);
or U13521 (N_13521,N_12970,N_12943);
and U13522 (N_13522,N_13047,N_13044);
nand U13523 (N_13523,N_13123,N_13102);
nor U13524 (N_13524,N_13034,N_12800);
nor U13525 (N_13525,N_12979,N_13096);
nand U13526 (N_13526,N_13107,N_12873);
and U13527 (N_13527,N_13015,N_13181);
nor U13528 (N_13528,N_12804,N_13089);
and U13529 (N_13529,N_12912,N_13044);
nor U13530 (N_13530,N_12940,N_13002);
nor U13531 (N_13531,N_13170,N_13043);
or U13532 (N_13532,N_13006,N_13163);
xor U13533 (N_13533,N_12904,N_13085);
nand U13534 (N_13534,N_13130,N_13092);
nor U13535 (N_13535,N_13184,N_13191);
nor U13536 (N_13536,N_13073,N_12829);
xnor U13537 (N_13537,N_13064,N_12915);
or U13538 (N_13538,N_13114,N_13164);
and U13539 (N_13539,N_13084,N_13107);
nand U13540 (N_13540,N_13015,N_13032);
or U13541 (N_13541,N_13041,N_13162);
and U13542 (N_13542,N_12803,N_13015);
and U13543 (N_13543,N_13086,N_13148);
and U13544 (N_13544,N_13115,N_12910);
nand U13545 (N_13545,N_12855,N_12907);
xor U13546 (N_13546,N_13175,N_12830);
xor U13547 (N_13547,N_12845,N_12966);
nor U13548 (N_13548,N_12811,N_13016);
and U13549 (N_13549,N_12829,N_13142);
xnor U13550 (N_13550,N_13105,N_12890);
or U13551 (N_13551,N_12933,N_12852);
nor U13552 (N_13552,N_13090,N_12843);
nand U13553 (N_13553,N_13103,N_13067);
nand U13554 (N_13554,N_13000,N_12891);
and U13555 (N_13555,N_12893,N_13050);
xnor U13556 (N_13556,N_12863,N_12857);
or U13557 (N_13557,N_12868,N_13023);
xor U13558 (N_13558,N_12988,N_13039);
nand U13559 (N_13559,N_12855,N_13089);
nor U13560 (N_13560,N_12932,N_13136);
nor U13561 (N_13561,N_12946,N_13178);
or U13562 (N_13562,N_12936,N_13006);
nor U13563 (N_13563,N_13027,N_12921);
and U13564 (N_13564,N_12841,N_13027);
nand U13565 (N_13565,N_12948,N_12957);
nand U13566 (N_13566,N_12886,N_12847);
xnor U13567 (N_13567,N_12960,N_12977);
or U13568 (N_13568,N_12890,N_12847);
nand U13569 (N_13569,N_12923,N_13098);
and U13570 (N_13570,N_13079,N_12958);
nand U13571 (N_13571,N_13173,N_13144);
nand U13572 (N_13572,N_13067,N_12924);
nor U13573 (N_13573,N_12989,N_13004);
or U13574 (N_13574,N_12835,N_13148);
nand U13575 (N_13575,N_12940,N_12872);
nor U13576 (N_13576,N_13077,N_12963);
or U13577 (N_13577,N_12931,N_13026);
nand U13578 (N_13578,N_12884,N_12907);
xnor U13579 (N_13579,N_12989,N_13152);
xnor U13580 (N_13580,N_13125,N_12815);
nor U13581 (N_13581,N_12985,N_12838);
xnor U13582 (N_13582,N_13044,N_12903);
nand U13583 (N_13583,N_13061,N_13111);
xnor U13584 (N_13584,N_13134,N_12878);
nand U13585 (N_13585,N_13045,N_12889);
or U13586 (N_13586,N_12872,N_13072);
nand U13587 (N_13587,N_12971,N_13118);
nand U13588 (N_13588,N_12917,N_13133);
or U13589 (N_13589,N_13014,N_12961);
and U13590 (N_13590,N_12843,N_13022);
nor U13591 (N_13591,N_13136,N_12862);
or U13592 (N_13592,N_13183,N_13137);
xnor U13593 (N_13593,N_13000,N_13009);
or U13594 (N_13594,N_13014,N_13067);
and U13595 (N_13595,N_12912,N_13198);
xor U13596 (N_13596,N_13103,N_12804);
and U13597 (N_13597,N_13023,N_13018);
and U13598 (N_13598,N_13173,N_13086);
xnor U13599 (N_13599,N_13044,N_12899);
or U13600 (N_13600,N_13407,N_13322);
nand U13601 (N_13601,N_13425,N_13561);
nand U13602 (N_13602,N_13507,N_13538);
xnor U13603 (N_13603,N_13473,N_13261);
nand U13604 (N_13604,N_13483,N_13280);
or U13605 (N_13605,N_13239,N_13206);
nor U13606 (N_13606,N_13581,N_13568);
xor U13607 (N_13607,N_13565,N_13479);
xor U13608 (N_13608,N_13505,N_13447);
nand U13609 (N_13609,N_13377,N_13274);
nand U13610 (N_13610,N_13435,N_13563);
nand U13611 (N_13611,N_13521,N_13552);
nor U13612 (N_13612,N_13354,N_13331);
and U13613 (N_13613,N_13550,N_13247);
nor U13614 (N_13614,N_13311,N_13293);
or U13615 (N_13615,N_13528,N_13269);
and U13616 (N_13616,N_13590,N_13352);
nand U13617 (N_13617,N_13591,N_13275);
and U13618 (N_13618,N_13276,N_13418);
or U13619 (N_13619,N_13502,N_13262);
nand U13620 (N_13620,N_13555,N_13258);
or U13621 (N_13621,N_13281,N_13303);
or U13622 (N_13622,N_13388,N_13395);
xor U13623 (N_13623,N_13490,N_13214);
nand U13624 (N_13624,N_13298,N_13254);
and U13625 (N_13625,N_13353,N_13569);
nor U13626 (N_13626,N_13558,N_13582);
nor U13627 (N_13627,N_13288,N_13336);
nor U13628 (N_13628,N_13575,N_13365);
and U13629 (N_13629,N_13235,N_13406);
xor U13630 (N_13630,N_13431,N_13291);
nand U13631 (N_13631,N_13452,N_13273);
nor U13632 (N_13632,N_13233,N_13500);
and U13633 (N_13633,N_13376,N_13351);
nor U13634 (N_13634,N_13559,N_13396);
and U13635 (N_13635,N_13543,N_13468);
and U13636 (N_13636,N_13339,N_13344);
xor U13637 (N_13637,N_13211,N_13284);
nor U13638 (N_13638,N_13330,N_13263);
xor U13639 (N_13639,N_13494,N_13266);
or U13640 (N_13640,N_13402,N_13333);
nor U13641 (N_13641,N_13485,N_13207);
nor U13642 (N_13642,N_13245,N_13203);
nor U13643 (N_13643,N_13212,N_13440);
xnor U13644 (N_13644,N_13516,N_13533);
nand U13645 (N_13645,N_13222,N_13551);
xnor U13646 (N_13646,N_13537,N_13314);
nand U13647 (N_13647,N_13340,N_13299);
and U13648 (N_13648,N_13360,N_13429);
nor U13649 (N_13649,N_13520,N_13259);
nand U13650 (N_13650,N_13545,N_13373);
nand U13651 (N_13651,N_13236,N_13470);
xnor U13652 (N_13652,N_13327,N_13315);
and U13653 (N_13653,N_13271,N_13387);
nand U13654 (N_13654,N_13290,N_13515);
nor U13655 (N_13655,N_13454,N_13240);
nor U13656 (N_13656,N_13488,N_13564);
or U13657 (N_13657,N_13328,N_13567);
and U13658 (N_13658,N_13560,N_13292);
xnor U13659 (N_13659,N_13209,N_13216);
nand U13660 (N_13660,N_13383,N_13295);
nor U13661 (N_13661,N_13498,N_13566);
xnor U13662 (N_13662,N_13369,N_13389);
or U13663 (N_13663,N_13326,N_13242);
and U13664 (N_13664,N_13296,N_13519);
or U13665 (N_13665,N_13524,N_13324);
or U13666 (N_13666,N_13231,N_13532);
nor U13667 (N_13667,N_13474,N_13596);
nand U13668 (N_13668,N_13514,N_13448);
nor U13669 (N_13669,N_13576,N_13244);
and U13670 (N_13670,N_13487,N_13204);
xnor U13671 (N_13671,N_13257,N_13285);
or U13672 (N_13672,N_13599,N_13363);
or U13673 (N_13673,N_13584,N_13335);
and U13674 (N_13674,N_13219,N_13531);
xnor U13675 (N_13675,N_13462,N_13409);
and U13676 (N_13676,N_13393,N_13323);
xor U13677 (N_13677,N_13509,N_13345);
nand U13678 (N_13678,N_13422,N_13405);
or U13679 (N_13679,N_13415,N_13234);
nand U13680 (N_13680,N_13264,N_13268);
xnor U13681 (N_13681,N_13398,N_13399);
and U13682 (N_13682,N_13530,N_13278);
or U13683 (N_13683,N_13541,N_13302);
nor U13684 (N_13684,N_13392,N_13546);
xor U13685 (N_13685,N_13381,N_13442);
or U13686 (N_13686,N_13391,N_13217);
xor U13687 (N_13687,N_13362,N_13346);
and U13688 (N_13688,N_13410,N_13441);
and U13689 (N_13689,N_13578,N_13492);
nor U13690 (N_13690,N_13553,N_13421);
or U13691 (N_13691,N_13301,N_13224);
and U13692 (N_13692,N_13501,N_13310);
nor U13693 (N_13693,N_13526,N_13510);
nor U13694 (N_13694,N_13549,N_13400);
nand U13695 (N_13695,N_13478,N_13408);
or U13696 (N_13696,N_13243,N_13556);
or U13697 (N_13697,N_13256,N_13282);
or U13698 (N_13698,N_13597,N_13270);
xor U13699 (N_13699,N_13542,N_13300);
and U13700 (N_13700,N_13205,N_13202);
xnor U13701 (N_13701,N_13332,N_13229);
nor U13702 (N_13702,N_13428,N_13417);
and U13703 (N_13703,N_13249,N_13252);
and U13704 (N_13704,N_13313,N_13367);
xor U13705 (N_13705,N_13529,N_13347);
nand U13706 (N_13706,N_13572,N_13312);
and U13707 (N_13707,N_13227,N_13592);
nor U13708 (N_13708,N_13366,N_13380);
or U13709 (N_13709,N_13469,N_13342);
xor U13710 (N_13710,N_13465,N_13201);
xor U13711 (N_13711,N_13386,N_13309);
or U13712 (N_13712,N_13458,N_13426);
xnor U13713 (N_13713,N_13489,N_13588);
nand U13714 (N_13714,N_13503,N_13277);
and U13715 (N_13715,N_13359,N_13595);
nor U13716 (N_13716,N_13539,N_13329);
and U13717 (N_13717,N_13449,N_13464);
nand U13718 (N_13718,N_13397,N_13210);
and U13719 (N_13719,N_13238,N_13385);
nor U13720 (N_13720,N_13356,N_13368);
nand U13721 (N_13721,N_13272,N_13294);
and U13722 (N_13722,N_13598,N_13308);
and U13723 (N_13723,N_13466,N_13304);
and U13724 (N_13724,N_13414,N_13562);
or U13725 (N_13725,N_13225,N_13355);
xnor U13726 (N_13726,N_13265,N_13477);
or U13727 (N_13727,N_13427,N_13350);
and U13728 (N_13728,N_13484,N_13499);
nand U13729 (N_13729,N_13475,N_13547);
xor U13730 (N_13730,N_13585,N_13544);
and U13731 (N_13731,N_13594,N_13432);
nor U13732 (N_13732,N_13446,N_13453);
xor U13733 (N_13733,N_13525,N_13450);
and U13734 (N_13734,N_13237,N_13341);
or U13735 (N_13735,N_13416,N_13384);
and U13736 (N_13736,N_13451,N_13434);
xor U13737 (N_13737,N_13493,N_13444);
and U13738 (N_13738,N_13583,N_13320);
nand U13739 (N_13739,N_13511,N_13480);
xor U13740 (N_13740,N_13589,N_13349);
xor U13741 (N_13741,N_13289,N_13213);
or U13742 (N_13742,N_13218,N_13587);
nand U13743 (N_13743,N_13443,N_13403);
and U13744 (N_13744,N_13506,N_13548);
or U13745 (N_13745,N_13423,N_13445);
nand U13746 (N_13746,N_13456,N_13574);
nor U13747 (N_13747,N_13325,N_13250);
nand U13748 (N_13748,N_13573,N_13287);
or U13749 (N_13749,N_13371,N_13241);
nand U13750 (N_13750,N_13557,N_13580);
and U13751 (N_13751,N_13246,N_13253);
nor U13752 (N_13752,N_13482,N_13316);
nor U13753 (N_13753,N_13455,N_13372);
nand U13754 (N_13754,N_13404,N_13215);
nand U13755 (N_13755,N_13226,N_13438);
nand U13756 (N_13756,N_13279,N_13518);
and U13757 (N_13757,N_13471,N_13413);
nor U13758 (N_13758,N_13463,N_13394);
nand U13759 (N_13759,N_13481,N_13297);
nor U13760 (N_13760,N_13579,N_13461);
xnor U13761 (N_13761,N_13439,N_13267);
xnor U13762 (N_13762,N_13255,N_13221);
or U13763 (N_13763,N_13593,N_13251);
nand U13764 (N_13764,N_13348,N_13419);
or U13765 (N_13765,N_13437,N_13486);
nand U13766 (N_13766,N_13390,N_13554);
and U13767 (N_13767,N_13586,N_13220);
nand U13768 (N_13768,N_13200,N_13307);
xnor U13769 (N_13769,N_13523,N_13286);
xor U13770 (N_13770,N_13305,N_13319);
xor U13771 (N_13771,N_13459,N_13321);
xnor U13772 (N_13772,N_13527,N_13374);
nor U13773 (N_13773,N_13248,N_13412);
and U13774 (N_13774,N_13338,N_13508);
xnor U13775 (N_13775,N_13378,N_13424);
and U13776 (N_13776,N_13513,N_13306);
and U13777 (N_13777,N_13472,N_13512);
and U13778 (N_13778,N_13357,N_13534);
or U13779 (N_13779,N_13467,N_13379);
or U13780 (N_13780,N_13497,N_13577);
or U13781 (N_13781,N_13318,N_13223);
and U13782 (N_13782,N_13334,N_13536);
and U13783 (N_13783,N_13230,N_13495);
nor U13784 (N_13784,N_13430,N_13491);
xnor U13785 (N_13785,N_13260,N_13436);
or U13786 (N_13786,N_13522,N_13401);
or U13787 (N_13787,N_13433,N_13540);
xnor U13788 (N_13788,N_13535,N_13496);
nor U13789 (N_13789,N_13382,N_13358);
xnor U13790 (N_13790,N_13571,N_13228);
nor U13791 (N_13791,N_13232,N_13375);
and U13792 (N_13792,N_13457,N_13476);
or U13793 (N_13793,N_13370,N_13283);
xnor U13794 (N_13794,N_13570,N_13364);
nor U13795 (N_13795,N_13504,N_13460);
nor U13796 (N_13796,N_13517,N_13317);
and U13797 (N_13797,N_13420,N_13411);
and U13798 (N_13798,N_13208,N_13361);
xnor U13799 (N_13799,N_13343,N_13337);
and U13800 (N_13800,N_13558,N_13480);
xor U13801 (N_13801,N_13361,N_13551);
nor U13802 (N_13802,N_13582,N_13544);
or U13803 (N_13803,N_13401,N_13499);
xor U13804 (N_13804,N_13543,N_13463);
and U13805 (N_13805,N_13288,N_13425);
or U13806 (N_13806,N_13416,N_13483);
xor U13807 (N_13807,N_13291,N_13311);
nand U13808 (N_13808,N_13388,N_13483);
nand U13809 (N_13809,N_13251,N_13499);
xnor U13810 (N_13810,N_13308,N_13411);
nand U13811 (N_13811,N_13363,N_13231);
nand U13812 (N_13812,N_13410,N_13453);
nor U13813 (N_13813,N_13272,N_13461);
and U13814 (N_13814,N_13222,N_13554);
nand U13815 (N_13815,N_13438,N_13462);
and U13816 (N_13816,N_13471,N_13254);
nand U13817 (N_13817,N_13248,N_13425);
nor U13818 (N_13818,N_13443,N_13322);
nand U13819 (N_13819,N_13227,N_13268);
or U13820 (N_13820,N_13379,N_13268);
and U13821 (N_13821,N_13313,N_13265);
nor U13822 (N_13822,N_13354,N_13244);
nand U13823 (N_13823,N_13231,N_13514);
nand U13824 (N_13824,N_13519,N_13596);
xor U13825 (N_13825,N_13480,N_13451);
nand U13826 (N_13826,N_13576,N_13510);
xor U13827 (N_13827,N_13572,N_13269);
nand U13828 (N_13828,N_13474,N_13494);
nand U13829 (N_13829,N_13541,N_13398);
and U13830 (N_13830,N_13513,N_13260);
and U13831 (N_13831,N_13593,N_13369);
and U13832 (N_13832,N_13235,N_13444);
nor U13833 (N_13833,N_13282,N_13489);
nor U13834 (N_13834,N_13509,N_13362);
nand U13835 (N_13835,N_13270,N_13423);
or U13836 (N_13836,N_13518,N_13261);
xor U13837 (N_13837,N_13550,N_13589);
nand U13838 (N_13838,N_13202,N_13317);
nor U13839 (N_13839,N_13237,N_13313);
and U13840 (N_13840,N_13329,N_13268);
and U13841 (N_13841,N_13493,N_13418);
nor U13842 (N_13842,N_13310,N_13508);
xor U13843 (N_13843,N_13223,N_13353);
xor U13844 (N_13844,N_13268,N_13525);
nand U13845 (N_13845,N_13328,N_13389);
or U13846 (N_13846,N_13213,N_13481);
or U13847 (N_13847,N_13532,N_13465);
nor U13848 (N_13848,N_13578,N_13371);
or U13849 (N_13849,N_13558,N_13342);
nand U13850 (N_13850,N_13239,N_13448);
xor U13851 (N_13851,N_13349,N_13297);
or U13852 (N_13852,N_13357,N_13220);
xor U13853 (N_13853,N_13216,N_13480);
nand U13854 (N_13854,N_13390,N_13312);
and U13855 (N_13855,N_13323,N_13593);
nor U13856 (N_13856,N_13307,N_13525);
nand U13857 (N_13857,N_13218,N_13364);
nand U13858 (N_13858,N_13591,N_13274);
or U13859 (N_13859,N_13321,N_13305);
nand U13860 (N_13860,N_13392,N_13252);
or U13861 (N_13861,N_13560,N_13466);
nor U13862 (N_13862,N_13280,N_13434);
nand U13863 (N_13863,N_13407,N_13593);
xnor U13864 (N_13864,N_13527,N_13483);
nand U13865 (N_13865,N_13268,N_13327);
nand U13866 (N_13866,N_13313,N_13317);
nor U13867 (N_13867,N_13535,N_13391);
or U13868 (N_13868,N_13306,N_13353);
xnor U13869 (N_13869,N_13518,N_13253);
nor U13870 (N_13870,N_13505,N_13317);
nand U13871 (N_13871,N_13332,N_13266);
xnor U13872 (N_13872,N_13343,N_13552);
or U13873 (N_13873,N_13383,N_13227);
nand U13874 (N_13874,N_13511,N_13443);
nand U13875 (N_13875,N_13274,N_13487);
xor U13876 (N_13876,N_13524,N_13558);
nand U13877 (N_13877,N_13551,N_13490);
nand U13878 (N_13878,N_13314,N_13576);
nand U13879 (N_13879,N_13257,N_13325);
or U13880 (N_13880,N_13579,N_13450);
and U13881 (N_13881,N_13287,N_13452);
and U13882 (N_13882,N_13368,N_13461);
and U13883 (N_13883,N_13307,N_13597);
and U13884 (N_13884,N_13226,N_13464);
nor U13885 (N_13885,N_13521,N_13250);
nand U13886 (N_13886,N_13405,N_13336);
xor U13887 (N_13887,N_13236,N_13248);
and U13888 (N_13888,N_13508,N_13577);
xor U13889 (N_13889,N_13244,N_13516);
or U13890 (N_13890,N_13553,N_13351);
or U13891 (N_13891,N_13267,N_13527);
or U13892 (N_13892,N_13417,N_13392);
or U13893 (N_13893,N_13353,N_13231);
or U13894 (N_13894,N_13448,N_13506);
or U13895 (N_13895,N_13381,N_13382);
xor U13896 (N_13896,N_13518,N_13242);
and U13897 (N_13897,N_13383,N_13422);
and U13898 (N_13898,N_13522,N_13524);
nand U13899 (N_13899,N_13319,N_13476);
xnor U13900 (N_13900,N_13363,N_13451);
nor U13901 (N_13901,N_13574,N_13245);
and U13902 (N_13902,N_13297,N_13425);
nand U13903 (N_13903,N_13482,N_13497);
nor U13904 (N_13904,N_13233,N_13205);
xnor U13905 (N_13905,N_13479,N_13380);
nand U13906 (N_13906,N_13290,N_13350);
or U13907 (N_13907,N_13440,N_13552);
xnor U13908 (N_13908,N_13533,N_13359);
nand U13909 (N_13909,N_13202,N_13367);
xor U13910 (N_13910,N_13343,N_13400);
or U13911 (N_13911,N_13563,N_13588);
xor U13912 (N_13912,N_13260,N_13206);
or U13913 (N_13913,N_13290,N_13388);
or U13914 (N_13914,N_13374,N_13239);
or U13915 (N_13915,N_13251,N_13354);
nor U13916 (N_13916,N_13479,N_13428);
nor U13917 (N_13917,N_13223,N_13316);
nand U13918 (N_13918,N_13240,N_13286);
and U13919 (N_13919,N_13317,N_13518);
or U13920 (N_13920,N_13579,N_13377);
or U13921 (N_13921,N_13384,N_13514);
nor U13922 (N_13922,N_13408,N_13242);
xor U13923 (N_13923,N_13510,N_13450);
and U13924 (N_13924,N_13265,N_13577);
xnor U13925 (N_13925,N_13246,N_13584);
or U13926 (N_13926,N_13350,N_13280);
or U13927 (N_13927,N_13560,N_13455);
or U13928 (N_13928,N_13335,N_13473);
nand U13929 (N_13929,N_13472,N_13295);
xor U13930 (N_13930,N_13548,N_13231);
xnor U13931 (N_13931,N_13518,N_13423);
or U13932 (N_13932,N_13409,N_13229);
nor U13933 (N_13933,N_13344,N_13209);
and U13934 (N_13934,N_13421,N_13499);
nor U13935 (N_13935,N_13325,N_13573);
nor U13936 (N_13936,N_13477,N_13208);
or U13937 (N_13937,N_13211,N_13374);
xnor U13938 (N_13938,N_13559,N_13402);
xnor U13939 (N_13939,N_13360,N_13384);
and U13940 (N_13940,N_13457,N_13470);
xnor U13941 (N_13941,N_13290,N_13300);
nand U13942 (N_13942,N_13324,N_13517);
and U13943 (N_13943,N_13598,N_13572);
nor U13944 (N_13944,N_13306,N_13229);
xnor U13945 (N_13945,N_13200,N_13587);
nor U13946 (N_13946,N_13477,N_13362);
nor U13947 (N_13947,N_13477,N_13465);
nand U13948 (N_13948,N_13508,N_13230);
nand U13949 (N_13949,N_13415,N_13342);
nor U13950 (N_13950,N_13474,N_13503);
nand U13951 (N_13951,N_13432,N_13333);
nand U13952 (N_13952,N_13323,N_13534);
xor U13953 (N_13953,N_13290,N_13309);
xnor U13954 (N_13954,N_13543,N_13488);
and U13955 (N_13955,N_13407,N_13513);
nand U13956 (N_13956,N_13535,N_13325);
nand U13957 (N_13957,N_13367,N_13292);
and U13958 (N_13958,N_13378,N_13369);
and U13959 (N_13959,N_13526,N_13384);
nand U13960 (N_13960,N_13395,N_13389);
or U13961 (N_13961,N_13488,N_13429);
nand U13962 (N_13962,N_13434,N_13450);
and U13963 (N_13963,N_13595,N_13213);
nand U13964 (N_13964,N_13409,N_13248);
xnor U13965 (N_13965,N_13281,N_13504);
or U13966 (N_13966,N_13245,N_13347);
nor U13967 (N_13967,N_13451,N_13331);
nor U13968 (N_13968,N_13249,N_13334);
xnor U13969 (N_13969,N_13478,N_13436);
nor U13970 (N_13970,N_13509,N_13598);
nand U13971 (N_13971,N_13500,N_13473);
and U13972 (N_13972,N_13569,N_13248);
or U13973 (N_13973,N_13215,N_13325);
xnor U13974 (N_13974,N_13256,N_13343);
nand U13975 (N_13975,N_13287,N_13588);
nand U13976 (N_13976,N_13322,N_13363);
or U13977 (N_13977,N_13310,N_13381);
and U13978 (N_13978,N_13599,N_13373);
and U13979 (N_13979,N_13430,N_13530);
nand U13980 (N_13980,N_13335,N_13431);
nand U13981 (N_13981,N_13489,N_13331);
and U13982 (N_13982,N_13356,N_13570);
or U13983 (N_13983,N_13475,N_13267);
xor U13984 (N_13984,N_13330,N_13200);
nand U13985 (N_13985,N_13399,N_13251);
nor U13986 (N_13986,N_13266,N_13246);
or U13987 (N_13987,N_13551,N_13330);
nand U13988 (N_13988,N_13426,N_13241);
and U13989 (N_13989,N_13239,N_13407);
nor U13990 (N_13990,N_13506,N_13556);
or U13991 (N_13991,N_13476,N_13396);
nand U13992 (N_13992,N_13588,N_13273);
nand U13993 (N_13993,N_13529,N_13482);
nor U13994 (N_13994,N_13398,N_13345);
or U13995 (N_13995,N_13356,N_13556);
nand U13996 (N_13996,N_13258,N_13245);
and U13997 (N_13997,N_13213,N_13575);
nor U13998 (N_13998,N_13294,N_13596);
xor U13999 (N_13999,N_13358,N_13329);
xnor U14000 (N_14000,N_13836,N_13875);
xor U14001 (N_14001,N_13724,N_13742);
nand U14002 (N_14002,N_13757,N_13796);
and U14003 (N_14003,N_13827,N_13865);
nor U14004 (N_14004,N_13993,N_13922);
xnor U14005 (N_14005,N_13741,N_13876);
nor U14006 (N_14006,N_13643,N_13846);
nand U14007 (N_14007,N_13961,N_13659);
xor U14008 (N_14008,N_13889,N_13957);
or U14009 (N_14009,N_13866,N_13853);
or U14010 (N_14010,N_13821,N_13691);
xnor U14011 (N_14011,N_13744,N_13705);
and U14012 (N_14012,N_13621,N_13829);
and U14013 (N_14013,N_13727,N_13650);
or U14014 (N_14014,N_13847,N_13785);
or U14015 (N_14015,N_13946,N_13607);
xnor U14016 (N_14016,N_13902,N_13817);
nor U14017 (N_14017,N_13604,N_13699);
nor U14018 (N_14018,N_13629,N_13769);
or U14019 (N_14019,N_13845,N_13759);
xor U14020 (N_14020,N_13996,N_13802);
nand U14021 (N_14021,N_13767,N_13894);
nand U14022 (N_14022,N_13735,N_13789);
nand U14023 (N_14023,N_13893,N_13753);
or U14024 (N_14024,N_13861,N_13891);
xnor U14025 (N_14025,N_13901,N_13873);
nand U14026 (N_14026,N_13954,N_13608);
nor U14027 (N_14027,N_13858,N_13755);
or U14028 (N_14028,N_13684,N_13663);
and U14029 (N_14029,N_13927,N_13968);
xor U14030 (N_14030,N_13812,N_13952);
or U14031 (N_14031,N_13740,N_13716);
and U14032 (N_14032,N_13850,N_13959);
and U14033 (N_14033,N_13841,N_13973);
nor U14034 (N_14034,N_13636,N_13931);
and U14035 (N_14035,N_13985,N_13635);
nand U14036 (N_14036,N_13881,N_13696);
or U14037 (N_14037,N_13765,N_13761);
nor U14038 (N_14038,N_13774,N_13868);
nor U14039 (N_14039,N_13899,N_13647);
nor U14040 (N_14040,N_13786,N_13864);
and U14041 (N_14041,N_13654,N_13657);
or U14042 (N_14042,N_13667,N_13860);
xnor U14043 (N_14043,N_13736,N_13780);
or U14044 (N_14044,N_13794,N_13668);
nor U14045 (N_14045,N_13665,N_13932);
nor U14046 (N_14046,N_13750,N_13711);
nand U14047 (N_14047,N_13944,N_13805);
and U14048 (N_14048,N_13690,N_13921);
and U14049 (N_14049,N_13801,N_13658);
and U14050 (N_14050,N_13601,N_13809);
or U14051 (N_14051,N_13938,N_13910);
or U14052 (N_14052,N_13631,N_13987);
nand U14053 (N_14053,N_13628,N_13625);
xor U14054 (N_14054,N_13939,N_13630);
xor U14055 (N_14055,N_13862,N_13773);
nor U14056 (N_14056,N_13984,N_13649);
nor U14057 (N_14057,N_13883,N_13977);
nor U14058 (N_14058,N_13639,N_13733);
nand U14059 (N_14059,N_13723,N_13760);
xor U14060 (N_14060,N_13701,N_13686);
nand U14061 (N_14061,N_13803,N_13721);
or U14062 (N_14062,N_13816,N_13634);
xor U14063 (N_14063,N_13675,N_13791);
and U14064 (N_14064,N_13758,N_13937);
nand U14065 (N_14065,N_13855,N_13974);
nor U14066 (N_14066,N_13678,N_13818);
xor U14067 (N_14067,N_13605,N_13839);
nand U14068 (N_14068,N_13978,N_13895);
and U14069 (N_14069,N_13660,N_13790);
nor U14070 (N_14070,N_13702,N_13618);
nand U14071 (N_14071,N_13935,N_13926);
xor U14072 (N_14072,N_13900,N_13924);
nand U14073 (N_14073,N_13971,N_13824);
xor U14074 (N_14074,N_13698,N_13929);
xnor U14075 (N_14075,N_13911,N_13933);
nand U14076 (N_14076,N_13754,N_13612);
nor U14077 (N_14077,N_13898,N_13897);
and U14078 (N_14078,N_13693,N_13857);
xnor U14079 (N_14079,N_13848,N_13787);
nand U14080 (N_14080,N_13700,N_13999);
xor U14081 (N_14081,N_13854,N_13990);
nor U14082 (N_14082,N_13718,N_13732);
xnor U14083 (N_14083,N_13603,N_13651);
or U14084 (N_14084,N_13619,N_13804);
xnor U14085 (N_14085,N_13878,N_13709);
nor U14086 (N_14086,N_13772,N_13731);
xnor U14087 (N_14087,N_13956,N_13793);
xnor U14088 (N_14088,N_13997,N_13670);
or U14089 (N_14089,N_13947,N_13975);
xor U14090 (N_14090,N_13638,N_13783);
nor U14091 (N_14091,N_13674,N_13842);
xor U14092 (N_14092,N_13917,N_13979);
nor U14093 (N_14093,N_13882,N_13676);
nor U14094 (N_14094,N_13697,N_13799);
and U14095 (N_14095,N_13943,N_13913);
xor U14096 (N_14096,N_13720,N_13749);
and U14097 (N_14097,N_13710,N_13872);
xnor U14098 (N_14098,N_13967,N_13677);
and U14099 (N_14099,N_13989,N_13641);
and U14100 (N_14100,N_13907,N_13906);
nor U14101 (N_14101,N_13779,N_13714);
and U14102 (N_14102,N_13622,N_13934);
nor U14103 (N_14103,N_13832,N_13752);
or U14104 (N_14104,N_13653,N_13645);
nor U14105 (N_14105,N_13879,N_13813);
or U14106 (N_14106,N_13940,N_13828);
and U14107 (N_14107,N_13852,N_13915);
xnor U14108 (N_14108,N_13781,N_13689);
and U14109 (N_14109,N_13726,N_13942);
or U14110 (N_14110,N_13916,N_13912);
or U14111 (N_14111,N_13719,N_13806);
and U14112 (N_14112,N_13950,N_13775);
nor U14113 (N_14113,N_13771,N_13725);
nor U14114 (N_14114,N_13648,N_13664);
and U14115 (N_14115,N_13666,N_13729);
and U14116 (N_14116,N_13966,N_13888);
nand U14117 (N_14117,N_13712,N_13609);
and U14118 (N_14118,N_13751,N_13885);
or U14119 (N_14119,N_13962,N_13994);
and U14120 (N_14120,N_13682,N_13834);
or U14121 (N_14121,N_13615,N_13970);
xnor U14122 (N_14122,N_13953,N_13814);
xor U14123 (N_14123,N_13798,N_13851);
nor U14124 (N_14124,N_13976,N_13863);
or U14125 (N_14125,N_13919,N_13884);
or U14126 (N_14126,N_13811,N_13825);
nor U14127 (N_14127,N_13903,N_13887);
nand U14128 (N_14128,N_13715,N_13672);
nand U14129 (N_14129,N_13688,N_13958);
or U14130 (N_14130,N_13788,N_13837);
xnor U14131 (N_14131,N_13764,N_13965);
xor U14132 (N_14132,N_13964,N_13998);
and U14133 (N_14133,N_13920,N_13610);
xnor U14134 (N_14134,N_13632,N_13704);
nor U14135 (N_14135,N_13745,N_13614);
nor U14136 (N_14136,N_13844,N_13706);
xnor U14137 (N_14137,N_13835,N_13722);
and U14138 (N_14138,N_13683,N_13792);
nor U14139 (N_14139,N_13661,N_13830);
or U14140 (N_14140,N_13877,N_13948);
xnor U14141 (N_14141,N_13856,N_13826);
or U14142 (N_14142,N_13743,N_13928);
or U14143 (N_14143,N_13695,N_13646);
xor U14144 (N_14144,N_13949,N_13748);
nand U14145 (N_14145,N_13822,N_13728);
nor U14146 (N_14146,N_13738,N_13692);
nand U14147 (N_14147,N_13681,N_13685);
nor U14148 (N_14148,N_13747,N_13810);
nor U14149 (N_14149,N_13746,N_13995);
nand U14150 (N_14150,N_13980,N_13880);
nor U14151 (N_14151,N_13800,N_13823);
or U14152 (N_14152,N_13623,N_13662);
and U14153 (N_14153,N_13784,N_13673);
or U14154 (N_14154,N_13963,N_13627);
nand U14155 (N_14155,N_13960,N_13730);
or U14156 (N_14156,N_13782,N_13819);
nand U14157 (N_14157,N_13909,N_13611);
xor U14158 (N_14158,N_13869,N_13708);
and U14159 (N_14159,N_13951,N_13671);
and U14160 (N_14160,N_13763,N_13840);
nor U14161 (N_14161,N_13988,N_13905);
xor U14162 (N_14162,N_13886,N_13624);
xor U14163 (N_14163,N_13707,N_13797);
nand U14164 (N_14164,N_13870,N_13602);
and U14165 (N_14165,N_13778,N_13859);
xor U14166 (N_14166,N_13713,N_13871);
xnor U14167 (N_14167,N_13892,N_13896);
nor U14168 (N_14168,N_13890,N_13756);
or U14169 (N_14169,N_13982,N_13992);
xor U14170 (N_14170,N_13640,N_13637);
or U14171 (N_14171,N_13777,N_13680);
and U14172 (N_14172,N_13655,N_13981);
nor U14173 (N_14173,N_13633,N_13669);
and U14174 (N_14174,N_13936,N_13955);
and U14175 (N_14175,N_13904,N_13613);
nand U14176 (N_14176,N_13795,N_13867);
nor U14177 (N_14177,N_13991,N_13644);
xor U14178 (N_14178,N_13983,N_13734);
or U14179 (N_14179,N_13831,N_13606);
nor U14180 (N_14180,N_13737,N_13656);
and U14181 (N_14181,N_13808,N_13843);
nor U14182 (N_14182,N_13923,N_13617);
nand U14183 (N_14183,N_13600,N_13838);
xnor U14184 (N_14184,N_13815,N_13620);
nor U14185 (N_14185,N_13941,N_13930);
xnor U14186 (N_14186,N_13717,N_13986);
xnor U14187 (N_14187,N_13945,N_13914);
nor U14188 (N_14188,N_13972,N_13770);
or U14189 (N_14189,N_13908,N_13626);
nand U14190 (N_14190,N_13703,N_13679);
or U14191 (N_14191,N_13874,N_13776);
xnor U14192 (N_14192,N_13642,N_13969);
nand U14193 (N_14193,N_13925,N_13849);
nand U14194 (N_14194,N_13833,N_13762);
xor U14195 (N_14195,N_13652,N_13807);
xor U14196 (N_14196,N_13918,N_13820);
nand U14197 (N_14197,N_13616,N_13768);
nor U14198 (N_14198,N_13739,N_13694);
nor U14199 (N_14199,N_13766,N_13687);
and U14200 (N_14200,N_13811,N_13772);
xor U14201 (N_14201,N_13986,N_13802);
nor U14202 (N_14202,N_13963,N_13907);
xnor U14203 (N_14203,N_13823,N_13910);
and U14204 (N_14204,N_13843,N_13889);
or U14205 (N_14205,N_13603,N_13983);
nand U14206 (N_14206,N_13798,N_13626);
xnor U14207 (N_14207,N_13695,N_13836);
nor U14208 (N_14208,N_13974,N_13822);
and U14209 (N_14209,N_13998,N_13706);
or U14210 (N_14210,N_13998,N_13968);
nand U14211 (N_14211,N_13807,N_13680);
nor U14212 (N_14212,N_13754,N_13616);
and U14213 (N_14213,N_13700,N_13974);
nor U14214 (N_14214,N_13775,N_13899);
or U14215 (N_14215,N_13911,N_13878);
or U14216 (N_14216,N_13603,N_13893);
nor U14217 (N_14217,N_13956,N_13872);
nor U14218 (N_14218,N_13832,N_13864);
nor U14219 (N_14219,N_13635,N_13945);
xnor U14220 (N_14220,N_13681,N_13844);
xnor U14221 (N_14221,N_13821,N_13733);
xnor U14222 (N_14222,N_13907,N_13926);
and U14223 (N_14223,N_13974,N_13804);
nand U14224 (N_14224,N_13741,N_13695);
nand U14225 (N_14225,N_13911,N_13674);
xor U14226 (N_14226,N_13666,N_13748);
nand U14227 (N_14227,N_13720,N_13787);
nand U14228 (N_14228,N_13709,N_13615);
or U14229 (N_14229,N_13882,N_13942);
nand U14230 (N_14230,N_13794,N_13843);
and U14231 (N_14231,N_13614,N_13786);
or U14232 (N_14232,N_13904,N_13910);
nand U14233 (N_14233,N_13625,N_13668);
or U14234 (N_14234,N_13607,N_13684);
nand U14235 (N_14235,N_13637,N_13804);
and U14236 (N_14236,N_13807,N_13933);
nand U14237 (N_14237,N_13694,N_13905);
nor U14238 (N_14238,N_13885,N_13977);
xor U14239 (N_14239,N_13609,N_13659);
or U14240 (N_14240,N_13638,N_13634);
xnor U14241 (N_14241,N_13759,N_13795);
nor U14242 (N_14242,N_13928,N_13979);
and U14243 (N_14243,N_13842,N_13688);
xor U14244 (N_14244,N_13990,N_13634);
nand U14245 (N_14245,N_13688,N_13754);
xnor U14246 (N_14246,N_13697,N_13660);
or U14247 (N_14247,N_13870,N_13960);
xor U14248 (N_14248,N_13955,N_13792);
nor U14249 (N_14249,N_13860,N_13916);
and U14250 (N_14250,N_13751,N_13877);
or U14251 (N_14251,N_13932,N_13662);
or U14252 (N_14252,N_13973,N_13793);
nor U14253 (N_14253,N_13749,N_13671);
xor U14254 (N_14254,N_13771,N_13755);
and U14255 (N_14255,N_13799,N_13990);
nand U14256 (N_14256,N_13972,N_13916);
or U14257 (N_14257,N_13625,N_13790);
or U14258 (N_14258,N_13743,N_13757);
or U14259 (N_14259,N_13682,N_13615);
or U14260 (N_14260,N_13743,N_13813);
or U14261 (N_14261,N_13988,N_13718);
and U14262 (N_14262,N_13887,N_13763);
or U14263 (N_14263,N_13977,N_13621);
or U14264 (N_14264,N_13757,N_13861);
nand U14265 (N_14265,N_13814,N_13952);
nor U14266 (N_14266,N_13710,N_13772);
xnor U14267 (N_14267,N_13607,N_13942);
and U14268 (N_14268,N_13682,N_13813);
nor U14269 (N_14269,N_13745,N_13874);
nor U14270 (N_14270,N_13844,N_13867);
nand U14271 (N_14271,N_13766,N_13991);
and U14272 (N_14272,N_13729,N_13807);
nor U14273 (N_14273,N_13738,N_13778);
and U14274 (N_14274,N_13780,N_13904);
xnor U14275 (N_14275,N_13912,N_13958);
xor U14276 (N_14276,N_13984,N_13664);
nand U14277 (N_14277,N_13747,N_13894);
xor U14278 (N_14278,N_13747,N_13778);
xor U14279 (N_14279,N_13658,N_13675);
nor U14280 (N_14280,N_13825,N_13928);
and U14281 (N_14281,N_13899,N_13955);
or U14282 (N_14282,N_13675,N_13861);
nand U14283 (N_14283,N_13816,N_13670);
and U14284 (N_14284,N_13786,N_13871);
nand U14285 (N_14285,N_13677,N_13958);
nand U14286 (N_14286,N_13862,N_13822);
or U14287 (N_14287,N_13782,N_13813);
and U14288 (N_14288,N_13739,N_13890);
or U14289 (N_14289,N_13842,N_13979);
and U14290 (N_14290,N_13929,N_13662);
nor U14291 (N_14291,N_13817,N_13923);
nor U14292 (N_14292,N_13992,N_13918);
xor U14293 (N_14293,N_13888,N_13734);
and U14294 (N_14294,N_13971,N_13805);
xnor U14295 (N_14295,N_13964,N_13871);
xor U14296 (N_14296,N_13849,N_13748);
xor U14297 (N_14297,N_13999,N_13773);
xnor U14298 (N_14298,N_13911,N_13831);
xnor U14299 (N_14299,N_13957,N_13829);
nor U14300 (N_14300,N_13630,N_13709);
and U14301 (N_14301,N_13804,N_13635);
nand U14302 (N_14302,N_13861,N_13614);
or U14303 (N_14303,N_13648,N_13854);
nor U14304 (N_14304,N_13803,N_13873);
nand U14305 (N_14305,N_13784,N_13982);
or U14306 (N_14306,N_13693,N_13977);
and U14307 (N_14307,N_13709,N_13776);
and U14308 (N_14308,N_13874,N_13987);
xnor U14309 (N_14309,N_13788,N_13630);
nand U14310 (N_14310,N_13839,N_13756);
and U14311 (N_14311,N_13857,N_13844);
nor U14312 (N_14312,N_13826,N_13753);
xnor U14313 (N_14313,N_13676,N_13861);
and U14314 (N_14314,N_13852,N_13917);
xor U14315 (N_14315,N_13683,N_13759);
xor U14316 (N_14316,N_13887,N_13711);
xor U14317 (N_14317,N_13783,N_13601);
nand U14318 (N_14318,N_13635,N_13699);
nor U14319 (N_14319,N_13606,N_13608);
or U14320 (N_14320,N_13936,N_13823);
nand U14321 (N_14321,N_13882,N_13993);
nor U14322 (N_14322,N_13908,N_13845);
nor U14323 (N_14323,N_13847,N_13805);
nor U14324 (N_14324,N_13792,N_13903);
nor U14325 (N_14325,N_13722,N_13635);
or U14326 (N_14326,N_13675,N_13763);
nand U14327 (N_14327,N_13675,N_13670);
nor U14328 (N_14328,N_13661,N_13971);
and U14329 (N_14329,N_13631,N_13801);
xnor U14330 (N_14330,N_13834,N_13664);
nor U14331 (N_14331,N_13849,N_13977);
or U14332 (N_14332,N_13981,N_13735);
and U14333 (N_14333,N_13867,N_13738);
nor U14334 (N_14334,N_13865,N_13861);
xor U14335 (N_14335,N_13896,N_13727);
or U14336 (N_14336,N_13644,N_13946);
nand U14337 (N_14337,N_13927,N_13899);
nand U14338 (N_14338,N_13691,N_13883);
and U14339 (N_14339,N_13776,N_13737);
nand U14340 (N_14340,N_13838,N_13768);
and U14341 (N_14341,N_13927,N_13797);
nor U14342 (N_14342,N_13873,N_13725);
nor U14343 (N_14343,N_13647,N_13732);
nor U14344 (N_14344,N_13729,N_13653);
or U14345 (N_14345,N_13999,N_13779);
nor U14346 (N_14346,N_13754,N_13625);
nand U14347 (N_14347,N_13649,N_13682);
or U14348 (N_14348,N_13912,N_13880);
nand U14349 (N_14349,N_13884,N_13668);
nor U14350 (N_14350,N_13975,N_13611);
and U14351 (N_14351,N_13698,N_13783);
and U14352 (N_14352,N_13769,N_13874);
nand U14353 (N_14353,N_13817,N_13829);
nand U14354 (N_14354,N_13928,N_13706);
xor U14355 (N_14355,N_13846,N_13743);
and U14356 (N_14356,N_13737,N_13821);
and U14357 (N_14357,N_13701,N_13746);
nand U14358 (N_14358,N_13720,N_13818);
nor U14359 (N_14359,N_13807,N_13926);
and U14360 (N_14360,N_13890,N_13627);
and U14361 (N_14361,N_13905,N_13940);
and U14362 (N_14362,N_13614,N_13905);
and U14363 (N_14363,N_13861,N_13828);
nand U14364 (N_14364,N_13883,N_13789);
xor U14365 (N_14365,N_13949,N_13957);
or U14366 (N_14366,N_13640,N_13881);
xnor U14367 (N_14367,N_13639,N_13613);
or U14368 (N_14368,N_13628,N_13612);
nand U14369 (N_14369,N_13774,N_13653);
and U14370 (N_14370,N_13743,N_13784);
or U14371 (N_14371,N_13729,N_13903);
or U14372 (N_14372,N_13849,N_13905);
nor U14373 (N_14373,N_13646,N_13854);
nor U14374 (N_14374,N_13801,N_13686);
xor U14375 (N_14375,N_13824,N_13987);
nor U14376 (N_14376,N_13716,N_13606);
nand U14377 (N_14377,N_13927,N_13919);
nor U14378 (N_14378,N_13973,N_13666);
or U14379 (N_14379,N_13936,N_13644);
nor U14380 (N_14380,N_13702,N_13621);
and U14381 (N_14381,N_13801,N_13920);
xnor U14382 (N_14382,N_13884,N_13804);
nor U14383 (N_14383,N_13892,N_13799);
or U14384 (N_14384,N_13660,N_13691);
xor U14385 (N_14385,N_13858,N_13977);
xor U14386 (N_14386,N_13999,N_13914);
or U14387 (N_14387,N_13882,N_13655);
and U14388 (N_14388,N_13682,N_13965);
xnor U14389 (N_14389,N_13997,N_13729);
and U14390 (N_14390,N_13764,N_13755);
and U14391 (N_14391,N_13692,N_13828);
or U14392 (N_14392,N_13911,N_13741);
nor U14393 (N_14393,N_13809,N_13894);
or U14394 (N_14394,N_13850,N_13970);
or U14395 (N_14395,N_13780,N_13940);
xnor U14396 (N_14396,N_13624,N_13774);
nor U14397 (N_14397,N_13743,N_13978);
or U14398 (N_14398,N_13763,N_13624);
xor U14399 (N_14399,N_13660,N_13783);
nand U14400 (N_14400,N_14266,N_14328);
or U14401 (N_14401,N_14320,N_14073);
xor U14402 (N_14402,N_14097,N_14282);
or U14403 (N_14403,N_14265,N_14160);
or U14404 (N_14404,N_14386,N_14177);
or U14405 (N_14405,N_14192,N_14157);
xor U14406 (N_14406,N_14311,N_14388);
and U14407 (N_14407,N_14348,N_14039);
or U14408 (N_14408,N_14061,N_14349);
xnor U14409 (N_14409,N_14333,N_14297);
nand U14410 (N_14410,N_14295,N_14197);
xor U14411 (N_14411,N_14245,N_14326);
nor U14412 (N_14412,N_14281,N_14151);
nand U14413 (N_14413,N_14307,N_14162);
nor U14414 (N_14414,N_14154,N_14389);
and U14415 (N_14415,N_14150,N_14263);
nand U14416 (N_14416,N_14004,N_14027);
xnor U14417 (N_14417,N_14082,N_14371);
nor U14418 (N_14418,N_14238,N_14274);
or U14419 (N_14419,N_14038,N_14012);
nor U14420 (N_14420,N_14092,N_14342);
nor U14421 (N_14421,N_14272,N_14122);
or U14422 (N_14422,N_14290,N_14198);
xnor U14423 (N_14423,N_14207,N_14341);
xor U14424 (N_14424,N_14277,N_14070);
or U14425 (N_14425,N_14099,N_14362);
and U14426 (N_14426,N_14114,N_14374);
nor U14427 (N_14427,N_14060,N_14105);
nor U14428 (N_14428,N_14120,N_14128);
xnor U14429 (N_14429,N_14392,N_14393);
nand U14430 (N_14430,N_14024,N_14344);
xnor U14431 (N_14431,N_14208,N_14214);
and U14432 (N_14432,N_14190,N_14353);
nand U14433 (N_14433,N_14255,N_14201);
and U14434 (N_14434,N_14074,N_14308);
and U14435 (N_14435,N_14111,N_14226);
and U14436 (N_14436,N_14303,N_14159);
xnor U14437 (N_14437,N_14363,N_14211);
or U14438 (N_14438,N_14279,N_14368);
nor U14439 (N_14439,N_14365,N_14137);
or U14440 (N_14440,N_14072,N_14324);
or U14441 (N_14441,N_14296,N_14172);
nand U14442 (N_14442,N_14025,N_14357);
nand U14443 (N_14443,N_14227,N_14140);
and U14444 (N_14444,N_14254,N_14044);
nand U14445 (N_14445,N_14045,N_14204);
nand U14446 (N_14446,N_14009,N_14314);
or U14447 (N_14447,N_14228,N_14185);
nor U14448 (N_14448,N_14196,N_14136);
or U14449 (N_14449,N_14306,N_14338);
or U14450 (N_14450,N_14123,N_14343);
nand U14451 (N_14451,N_14098,N_14110);
xor U14452 (N_14452,N_14301,N_14148);
or U14453 (N_14453,N_14218,N_14315);
xor U14454 (N_14454,N_14312,N_14260);
xnor U14455 (N_14455,N_14212,N_14232);
xor U14456 (N_14456,N_14119,N_14370);
or U14457 (N_14457,N_14037,N_14210);
or U14458 (N_14458,N_14209,N_14133);
nand U14459 (N_14459,N_14020,N_14135);
nand U14460 (N_14460,N_14294,N_14355);
xnor U14461 (N_14461,N_14068,N_14077);
and U14462 (N_14462,N_14256,N_14216);
and U14463 (N_14463,N_14375,N_14166);
and U14464 (N_14464,N_14002,N_14213);
xor U14465 (N_14465,N_14359,N_14366);
or U14466 (N_14466,N_14367,N_14270);
xnor U14467 (N_14467,N_14138,N_14113);
xnor U14468 (N_14468,N_14052,N_14396);
and U14469 (N_14469,N_14088,N_14143);
nor U14470 (N_14470,N_14101,N_14283);
nor U14471 (N_14471,N_14167,N_14066);
or U14472 (N_14472,N_14153,N_14164);
and U14473 (N_14473,N_14243,N_14183);
nor U14474 (N_14474,N_14313,N_14079);
and U14475 (N_14475,N_14316,N_14321);
nand U14476 (N_14476,N_14076,N_14332);
or U14477 (N_14477,N_14331,N_14284);
nor U14478 (N_14478,N_14309,N_14129);
nor U14479 (N_14479,N_14194,N_14398);
xor U14480 (N_14480,N_14174,N_14013);
nand U14481 (N_14481,N_14125,N_14250);
nor U14482 (N_14482,N_14147,N_14291);
nand U14483 (N_14483,N_14087,N_14195);
nor U14484 (N_14484,N_14188,N_14369);
and U14485 (N_14485,N_14053,N_14121);
nand U14486 (N_14486,N_14117,N_14221);
xnor U14487 (N_14487,N_14134,N_14000);
xor U14488 (N_14488,N_14032,N_14382);
nor U14489 (N_14489,N_14163,N_14030);
xnor U14490 (N_14490,N_14397,N_14050);
or U14491 (N_14491,N_14399,N_14086);
nand U14492 (N_14492,N_14028,N_14305);
nand U14493 (N_14493,N_14327,N_14175);
xnor U14494 (N_14494,N_14288,N_14299);
and U14495 (N_14495,N_14035,N_14139);
xor U14496 (N_14496,N_14394,N_14253);
nand U14497 (N_14497,N_14340,N_14006);
nor U14498 (N_14498,N_14161,N_14026);
nand U14499 (N_14499,N_14247,N_14352);
nand U14500 (N_14500,N_14023,N_14176);
nand U14501 (N_14501,N_14165,N_14078);
and U14502 (N_14502,N_14054,N_14132);
xor U14503 (N_14503,N_14219,N_14081);
or U14504 (N_14504,N_14107,N_14093);
xnor U14505 (N_14505,N_14378,N_14347);
or U14506 (N_14506,N_14285,N_14156);
xor U14507 (N_14507,N_14067,N_14115);
or U14508 (N_14508,N_14267,N_14003);
and U14509 (N_14509,N_14130,N_14178);
and U14510 (N_14510,N_14109,N_14293);
nand U14511 (N_14511,N_14395,N_14036);
nor U14512 (N_14512,N_14155,N_14339);
xor U14513 (N_14513,N_14335,N_14016);
xor U14514 (N_14514,N_14276,N_14055);
or U14515 (N_14515,N_14298,N_14126);
nor U14516 (N_14516,N_14096,N_14206);
nor U14517 (N_14517,N_14231,N_14018);
xor U14518 (N_14518,N_14080,N_14257);
nand U14519 (N_14519,N_14358,N_14259);
nand U14520 (N_14520,N_14318,N_14031);
xnor U14521 (N_14521,N_14381,N_14390);
nand U14522 (N_14522,N_14225,N_14051);
xor U14523 (N_14523,N_14391,N_14350);
nand U14524 (N_14524,N_14236,N_14075);
or U14525 (N_14525,N_14102,N_14233);
xor U14526 (N_14526,N_14095,N_14220);
xnor U14527 (N_14527,N_14149,N_14071);
xor U14528 (N_14528,N_14189,N_14083);
or U14529 (N_14529,N_14187,N_14124);
nor U14530 (N_14530,N_14289,N_14364);
or U14531 (N_14531,N_14021,N_14062);
and U14532 (N_14532,N_14262,N_14323);
xnor U14533 (N_14533,N_14043,N_14380);
nor U14534 (N_14534,N_14215,N_14084);
or U14535 (N_14535,N_14063,N_14317);
nand U14536 (N_14536,N_14372,N_14385);
nor U14537 (N_14537,N_14180,N_14361);
nor U14538 (N_14538,N_14376,N_14251);
nand U14539 (N_14539,N_14104,N_14108);
or U14540 (N_14540,N_14015,N_14235);
nand U14541 (N_14541,N_14239,N_14041);
xor U14542 (N_14542,N_14005,N_14103);
and U14543 (N_14543,N_14040,N_14058);
and U14544 (N_14544,N_14186,N_14152);
xnor U14545 (N_14545,N_14230,N_14203);
xor U14546 (N_14546,N_14089,N_14345);
nor U14547 (N_14547,N_14278,N_14173);
or U14548 (N_14548,N_14240,N_14275);
and U14549 (N_14549,N_14168,N_14094);
nor U14550 (N_14550,N_14034,N_14019);
and U14551 (N_14551,N_14127,N_14319);
nand U14552 (N_14552,N_14202,N_14179);
or U14553 (N_14553,N_14310,N_14205);
xnor U14554 (N_14554,N_14191,N_14141);
xnor U14555 (N_14555,N_14056,N_14325);
nand U14556 (N_14556,N_14100,N_14118);
and U14557 (N_14557,N_14229,N_14384);
or U14558 (N_14558,N_14354,N_14142);
nor U14559 (N_14559,N_14112,N_14046);
nor U14560 (N_14560,N_14171,N_14090);
nand U14561 (N_14561,N_14377,N_14057);
nand U14562 (N_14562,N_14302,N_14047);
and U14563 (N_14563,N_14106,N_14346);
or U14564 (N_14564,N_14329,N_14008);
nor U14565 (N_14565,N_14182,N_14200);
and U14566 (N_14566,N_14387,N_14234);
nand U14567 (N_14567,N_14193,N_14286);
and U14568 (N_14568,N_14199,N_14059);
nand U14569 (N_14569,N_14287,N_14224);
nor U14570 (N_14570,N_14249,N_14258);
and U14571 (N_14571,N_14269,N_14222);
and U14572 (N_14572,N_14170,N_14337);
nor U14573 (N_14573,N_14322,N_14237);
xor U14574 (N_14574,N_14158,N_14007);
nand U14575 (N_14575,N_14069,N_14336);
or U14576 (N_14576,N_14091,N_14252);
or U14577 (N_14577,N_14268,N_14304);
nor U14578 (N_14578,N_14383,N_14292);
xor U14579 (N_14579,N_14181,N_14022);
xor U14580 (N_14580,N_14261,N_14273);
or U14581 (N_14581,N_14351,N_14029);
nor U14582 (N_14582,N_14330,N_14264);
nor U14583 (N_14583,N_14373,N_14010);
xnor U14584 (N_14584,N_14223,N_14379);
xor U14585 (N_14585,N_14242,N_14048);
or U14586 (N_14586,N_14217,N_14049);
nand U14587 (N_14587,N_14001,N_14184);
and U14588 (N_14588,N_14244,N_14085);
xor U14589 (N_14589,N_14017,N_14241);
and U14590 (N_14590,N_14145,N_14356);
nor U14591 (N_14591,N_14144,N_14131);
or U14592 (N_14592,N_14360,N_14248);
xnor U14593 (N_14593,N_14271,N_14246);
or U14594 (N_14594,N_14033,N_14334);
nor U14595 (N_14595,N_14014,N_14280);
nor U14596 (N_14596,N_14116,N_14169);
and U14597 (N_14597,N_14300,N_14065);
xor U14598 (N_14598,N_14011,N_14064);
and U14599 (N_14599,N_14146,N_14042);
nand U14600 (N_14600,N_14320,N_14028);
nand U14601 (N_14601,N_14272,N_14066);
nand U14602 (N_14602,N_14346,N_14242);
and U14603 (N_14603,N_14362,N_14304);
and U14604 (N_14604,N_14264,N_14365);
or U14605 (N_14605,N_14064,N_14217);
nor U14606 (N_14606,N_14203,N_14283);
or U14607 (N_14607,N_14393,N_14253);
nand U14608 (N_14608,N_14382,N_14185);
or U14609 (N_14609,N_14170,N_14058);
nand U14610 (N_14610,N_14234,N_14146);
nand U14611 (N_14611,N_14074,N_14386);
and U14612 (N_14612,N_14333,N_14284);
and U14613 (N_14613,N_14370,N_14254);
xnor U14614 (N_14614,N_14112,N_14255);
xnor U14615 (N_14615,N_14324,N_14303);
and U14616 (N_14616,N_14163,N_14223);
and U14617 (N_14617,N_14295,N_14227);
xnor U14618 (N_14618,N_14222,N_14178);
or U14619 (N_14619,N_14224,N_14355);
xnor U14620 (N_14620,N_14164,N_14188);
xnor U14621 (N_14621,N_14096,N_14280);
xnor U14622 (N_14622,N_14377,N_14153);
xnor U14623 (N_14623,N_14342,N_14114);
nand U14624 (N_14624,N_14114,N_14090);
nand U14625 (N_14625,N_14269,N_14398);
nand U14626 (N_14626,N_14377,N_14265);
nor U14627 (N_14627,N_14130,N_14396);
and U14628 (N_14628,N_14358,N_14238);
or U14629 (N_14629,N_14376,N_14281);
and U14630 (N_14630,N_14079,N_14224);
nor U14631 (N_14631,N_14187,N_14095);
xnor U14632 (N_14632,N_14206,N_14335);
nor U14633 (N_14633,N_14358,N_14332);
xnor U14634 (N_14634,N_14357,N_14230);
and U14635 (N_14635,N_14372,N_14160);
and U14636 (N_14636,N_14342,N_14097);
nand U14637 (N_14637,N_14314,N_14035);
or U14638 (N_14638,N_14003,N_14304);
nand U14639 (N_14639,N_14223,N_14081);
and U14640 (N_14640,N_14043,N_14252);
nor U14641 (N_14641,N_14048,N_14179);
and U14642 (N_14642,N_14335,N_14128);
xor U14643 (N_14643,N_14105,N_14251);
nand U14644 (N_14644,N_14308,N_14351);
nor U14645 (N_14645,N_14268,N_14354);
or U14646 (N_14646,N_14214,N_14376);
xor U14647 (N_14647,N_14260,N_14069);
and U14648 (N_14648,N_14236,N_14055);
xnor U14649 (N_14649,N_14210,N_14272);
nand U14650 (N_14650,N_14340,N_14026);
nor U14651 (N_14651,N_14338,N_14077);
and U14652 (N_14652,N_14027,N_14345);
or U14653 (N_14653,N_14165,N_14221);
or U14654 (N_14654,N_14334,N_14245);
xor U14655 (N_14655,N_14296,N_14331);
and U14656 (N_14656,N_14262,N_14181);
nand U14657 (N_14657,N_14345,N_14341);
or U14658 (N_14658,N_14272,N_14320);
nor U14659 (N_14659,N_14115,N_14332);
and U14660 (N_14660,N_14246,N_14294);
or U14661 (N_14661,N_14205,N_14359);
nand U14662 (N_14662,N_14301,N_14105);
nand U14663 (N_14663,N_14390,N_14255);
and U14664 (N_14664,N_14225,N_14362);
and U14665 (N_14665,N_14132,N_14206);
nand U14666 (N_14666,N_14213,N_14180);
and U14667 (N_14667,N_14318,N_14397);
and U14668 (N_14668,N_14299,N_14103);
or U14669 (N_14669,N_14255,N_14142);
xnor U14670 (N_14670,N_14060,N_14352);
nand U14671 (N_14671,N_14161,N_14247);
nor U14672 (N_14672,N_14230,N_14197);
and U14673 (N_14673,N_14399,N_14298);
nor U14674 (N_14674,N_14158,N_14246);
nand U14675 (N_14675,N_14010,N_14121);
and U14676 (N_14676,N_14127,N_14154);
nor U14677 (N_14677,N_14283,N_14261);
nand U14678 (N_14678,N_14168,N_14230);
nand U14679 (N_14679,N_14102,N_14059);
nor U14680 (N_14680,N_14272,N_14072);
xor U14681 (N_14681,N_14062,N_14248);
xnor U14682 (N_14682,N_14160,N_14163);
nor U14683 (N_14683,N_14335,N_14136);
nand U14684 (N_14684,N_14103,N_14119);
or U14685 (N_14685,N_14232,N_14004);
xor U14686 (N_14686,N_14285,N_14253);
or U14687 (N_14687,N_14393,N_14111);
nor U14688 (N_14688,N_14063,N_14034);
nand U14689 (N_14689,N_14096,N_14311);
and U14690 (N_14690,N_14351,N_14358);
and U14691 (N_14691,N_14205,N_14221);
xor U14692 (N_14692,N_14127,N_14134);
and U14693 (N_14693,N_14028,N_14052);
xnor U14694 (N_14694,N_14278,N_14140);
xnor U14695 (N_14695,N_14254,N_14280);
xnor U14696 (N_14696,N_14229,N_14380);
nor U14697 (N_14697,N_14272,N_14204);
and U14698 (N_14698,N_14234,N_14325);
nand U14699 (N_14699,N_14138,N_14313);
xnor U14700 (N_14700,N_14026,N_14282);
nand U14701 (N_14701,N_14234,N_14128);
nand U14702 (N_14702,N_14323,N_14186);
nand U14703 (N_14703,N_14130,N_14174);
nand U14704 (N_14704,N_14126,N_14346);
nand U14705 (N_14705,N_14250,N_14365);
or U14706 (N_14706,N_14057,N_14189);
or U14707 (N_14707,N_14340,N_14043);
or U14708 (N_14708,N_14191,N_14337);
nor U14709 (N_14709,N_14205,N_14138);
or U14710 (N_14710,N_14276,N_14152);
or U14711 (N_14711,N_14171,N_14054);
xnor U14712 (N_14712,N_14346,N_14214);
or U14713 (N_14713,N_14377,N_14214);
nand U14714 (N_14714,N_14252,N_14021);
or U14715 (N_14715,N_14122,N_14036);
nor U14716 (N_14716,N_14228,N_14247);
and U14717 (N_14717,N_14254,N_14388);
nor U14718 (N_14718,N_14182,N_14298);
or U14719 (N_14719,N_14271,N_14065);
and U14720 (N_14720,N_14221,N_14213);
or U14721 (N_14721,N_14247,N_14128);
and U14722 (N_14722,N_14093,N_14147);
or U14723 (N_14723,N_14283,N_14251);
xnor U14724 (N_14724,N_14151,N_14374);
or U14725 (N_14725,N_14079,N_14022);
xor U14726 (N_14726,N_14004,N_14116);
nor U14727 (N_14727,N_14041,N_14198);
xnor U14728 (N_14728,N_14078,N_14300);
xor U14729 (N_14729,N_14335,N_14028);
xnor U14730 (N_14730,N_14046,N_14379);
nor U14731 (N_14731,N_14037,N_14300);
and U14732 (N_14732,N_14243,N_14293);
or U14733 (N_14733,N_14380,N_14276);
and U14734 (N_14734,N_14238,N_14188);
and U14735 (N_14735,N_14086,N_14013);
nand U14736 (N_14736,N_14350,N_14011);
nand U14737 (N_14737,N_14326,N_14262);
and U14738 (N_14738,N_14035,N_14067);
or U14739 (N_14739,N_14268,N_14235);
and U14740 (N_14740,N_14128,N_14000);
nand U14741 (N_14741,N_14380,N_14144);
or U14742 (N_14742,N_14303,N_14296);
nor U14743 (N_14743,N_14119,N_14286);
xor U14744 (N_14744,N_14138,N_14261);
and U14745 (N_14745,N_14208,N_14203);
or U14746 (N_14746,N_14252,N_14059);
nor U14747 (N_14747,N_14088,N_14272);
and U14748 (N_14748,N_14338,N_14398);
nand U14749 (N_14749,N_14173,N_14098);
or U14750 (N_14750,N_14009,N_14372);
and U14751 (N_14751,N_14368,N_14198);
or U14752 (N_14752,N_14189,N_14046);
nand U14753 (N_14753,N_14332,N_14176);
nand U14754 (N_14754,N_14068,N_14372);
and U14755 (N_14755,N_14164,N_14060);
and U14756 (N_14756,N_14246,N_14175);
and U14757 (N_14757,N_14224,N_14163);
xnor U14758 (N_14758,N_14289,N_14005);
and U14759 (N_14759,N_14331,N_14127);
and U14760 (N_14760,N_14004,N_14073);
xor U14761 (N_14761,N_14344,N_14071);
nor U14762 (N_14762,N_14081,N_14311);
nand U14763 (N_14763,N_14280,N_14179);
nand U14764 (N_14764,N_14120,N_14178);
and U14765 (N_14765,N_14094,N_14187);
or U14766 (N_14766,N_14125,N_14261);
or U14767 (N_14767,N_14319,N_14180);
and U14768 (N_14768,N_14126,N_14063);
or U14769 (N_14769,N_14003,N_14241);
nand U14770 (N_14770,N_14079,N_14024);
or U14771 (N_14771,N_14042,N_14230);
nand U14772 (N_14772,N_14218,N_14280);
and U14773 (N_14773,N_14169,N_14125);
and U14774 (N_14774,N_14312,N_14122);
or U14775 (N_14775,N_14154,N_14148);
or U14776 (N_14776,N_14075,N_14161);
xor U14777 (N_14777,N_14251,N_14134);
nand U14778 (N_14778,N_14293,N_14193);
or U14779 (N_14779,N_14232,N_14078);
nand U14780 (N_14780,N_14324,N_14299);
or U14781 (N_14781,N_14042,N_14267);
xor U14782 (N_14782,N_14393,N_14145);
xnor U14783 (N_14783,N_14035,N_14200);
xor U14784 (N_14784,N_14033,N_14117);
nor U14785 (N_14785,N_14338,N_14281);
xor U14786 (N_14786,N_14387,N_14252);
and U14787 (N_14787,N_14231,N_14131);
nor U14788 (N_14788,N_14256,N_14365);
and U14789 (N_14789,N_14295,N_14018);
or U14790 (N_14790,N_14194,N_14167);
xor U14791 (N_14791,N_14103,N_14394);
or U14792 (N_14792,N_14155,N_14011);
and U14793 (N_14793,N_14019,N_14187);
nor U14794 (N_14794,N_14158,N_14032);
nand U14795 (N_14795,N_14218,N_14393);
xnor U14796 (N_14796,N_14109,N_14356);
or U14797 (N_14797,N_14363,N_14245);
xor U14798 (N_14798,N_14030,N_14021);
nor U14799 (N_14799,N_14373,N_14063);
or U14800 (N_14800,N_14685,N_14448);
xor U14801 (N_14801,N_14626,N_14738);
nand U14802 (N_14802,N_14405,N_14794);
and U14803 (N_14803,N_14759,N_14535);
xnor U14804 (N_14804,N_14744,N_14750);
nor U14805 (N_14805,N_14472,N_14428);
nor U14806 (N_14806,N_14491,N_14436);
nor U14807 (N_14807,N_14758,N_14409);
and U14808 (N_14808,N_14473,N_14585);
nor U14809 (N_14809,N_14665,N_14781);
nand U14810 (N_14810,N_14414,N_14559);
or U14811 (N_14811,N_14568,N_14505);
nand U14812 (N_14812,N_14523,N_14517);
nor U14813 (N_14813,N_14779,N_14466);
xor U14814 (N_14814,N_14459,N_14542);
nor U14815 (N_14815,N_14449,N_14622);
nor U14816 (N_14816,N_14403,N_14538);
xnor U14817 (N_14817,N_14760,N_14445);
and U14818 (N_14818,N_14704,N_14452);
and U14819 (N_14819,N_14765,N_14516);
nor U14820 (N_14820,N_14700,N_14745);
and U14821 (N_14821,N_14601,N_14737);
nand U14822 (N_14822,N_14537,N_14690);
xor U14823 (N_14823,N_14464,N_14769);
nor U14824 (N_14824,N_14788,N_14584);
and U14825 (N_14825,N_14660,N_14504);
nand U14826 (N_14826,N_14512,N_14555);
xnor U14827 (N_14827,N_14733,N_14729);
and U14828 (N_14828,N_14574,N_14708);
and U14829 (N_14829,N_14619,N_14616);
or U14830 (N_14830,N_14688,N_14446);
or U14831 (N_14831,N_14698,N_14582);
and U14832 (N_14832,N_14757,N_14544);
nand U14833 (N_14833,N_14790,N_14402);
nand U14834 (N_14834,N_14599,N_14486);
nor U14835 (N_14835,N_14623,N_14653);
nor U14836 (N_14836,N_14454,N_14628);
xnor U14837 (N_14837,N_14477,N_14658);
or U14838 (N_14838,N_14670,N_14720);
xnor U14839 (N_14839,N_14485,N_14451);
and U14840 (N_14840,N_14596,N_14499);
nand U14841 (N_14841,N_14591,N_14426);
xnor U14842 (N_14842,N_14631,N_14749);
nand U14843 (N_14843,N_14427,N_14641);
or U14844 (N_14844,N_14595,N_14593);
nor U14845 (N_14845,N_14598,N_14527);
nor U14846 (N_14846,N_14672,N_14719);
nor U14847 (N_14847,N_14606,N_14659);
nor U14848 (N_14848,N_14774,N_14488);
nand U14849 (N_14849,N_14566,N_14586);
or U14850 (N_14850,N_14649,N_14524);
and U14851 (N_14851,N_14753,N_14764);
or U14852 (N_14852,N_14681,N_14652);
and U14853 (N_14853,N_14715,N_14514);
nand U14854 (N_14854,N_14554,N_14754);
and U14855 (N_14855,N_14518,N_14430);
and U14856 (N_14856,N_14705,N_14410);
and U14857 (N_14857,N_14456,N_14742);
xnor U14858 (N_14858,N_14493,N_14716);
and U14859 (N_14859,N_14655,N_14689);
nand U14860 (N_14860,N_14510,N_14480);
and U14861 (N_14861,N_14701,N_14686);
xnor U14862 (N_14862,N_14597,N_14792);
and U14863 (N_14863,N_14608,N_14576);
or U14864 (N_14864,N_14588,N_14646);
or U14865 (N_14865,N_14422,N_14661);
or U14866 (N_14866,N_14425,N_14400);
nor U14867 (N_14867,N_14479,N_14650);
nor U14868 (N_14868,N_14693,N_14780);
nor U14869 (N_14869,N_14755,N_14478);
nor U14870 (N_14870,N_14613,N_14432);
nor U14871 (N_14871,N_14547,N_14577);
nor U14872 (N_14872,N_14522,N_14723);
xnor U14873 (N_14873,N_14531,N_14447);
or U14874 (N_14874,N_14590,N_14564);
nand U14875 (N_14875,N_14444,N_14634);
xor U14876 (N_14876,N_14567,N_14640);
or U14877 (N_14877,N_14408,N_14533);
nand U14878 (N_14878,N_14740,N_14416);
nand U14879 (N_14879,N_14691,N_14743);
and U14880 (N_14880,N_14766,N_14415);
nor U14881 (N_14881,N_14607,N_14433);
or U14882 (N_14882,N_14696,N_14471);
and U14883 (N_14883,N_14682,N_14530);
nand U14884 (N_14884,N_14508,N_14437);
and U14885 (N_14885,N_14761,N_14552);
and U14886 (N_14886,N_14594,N_14721);
nor U14887 (N_14887,N_14679,N_14560);
nand U14888 (N_14888,N_14673,N_14789);
nor U14889 (N_14889,N_14773,N_14618);
or U14890 (N_14890,N_14797,N_14741);
or U14891 (N_14891,N_14467,N_14777);
nor U14892 (N_14892,N_14614,N_14419);
nor U14893 (N_14893,N_14482,N_14624);
nand U14894 (N_14894,N_14589,N_14475);
nand U14895 (N_14895,N_14726,N_14648);
and U14896 (N_14896,N_14731,N_14602);
or U14897 (N_14897,N_14639,N_14645);
xor U14898 (N_14898,N_14534,N_14664);
or U14899 (N_14899,N_14787,N_14748);
nor U14900 (N_14900,N_14735,N_14651);
nor U14901 (N_14901,N_14610,N_14439);
or U14902 (N_14902,N_14717,N_14553);
or U14903 (N_14903,N_14751,N_14718);
or U14904 (N_14904,N_14644,N_14462);
nor U14905 (N_14905,N_14418,N_14404);
and U14906 (N_14906,N_14487,N_14540);
and U14907 (N_14907,N_14711,N_14621);
or U14908 (N_14908,N_14775,N_14678);
or U14909 (N_14909,N_14550,N_14662);
nor U14910 (N_14910,N_14793,N_14656);
nor U14911 (N_14911,N_14627,N_14529);
nor U14912 (N_14912,N_14495,N_14615);
or U14913 (N_14913,N_14581,N_14706);
nor U14914 (N_14914,N_14450,N_14580);
nor U14915 (N_14915,N_14677,N_14785);
xnor U14916 (N_14916,N_14521,N_14736);
and U14917 (N_14917,N_14515,N_14481);
or U14918 (N_14918,N_14675,N_14676);
nor U14919 (N_14919,N_14669,N_14710);
nand U14920 (N_14920,N_14603,N_14712);
xor U14921 (N_14921,N_14509,N_14539);
nand U14922 (N_14922,N_14635,N_14578);
and U14923 (N_14923,N_14500,N_14506);
xnor U14924 (N_14924,N_14674,N_14734);
or U14925 (N_14925,N_14440,N_14784);
xor U14926 (N_14926,N_14490,N_14697);
or U14927 (N_14927,N_14747,N_14470);
xor U14928 (N_14928,N_14667,N_14556);
nor U14929 (N_14929,N_14507,N_14489);
nand U14930 (N_14930,N_14474,N_14543);
nand U14931 (N_14931,N_14727,N_14548);
and U14932 (N_14932,N_14722,N_14438);
nand U14933 (N_14933,N_14546,N_14767);
and U14934 (N_14934,N_14483,N_14457);
nor U14935 (N_14935,N_14782,N_14545);
or U14936 (N_14936,N_14768,N_14680);
xnor U14937 (N_14937,N_14569,N_14783);
xnor U14938 (N_14938,N_14604,N_14429);
xnor U14939 (N_14939,N_14776,N_14513);
xnor U14940 (N_14940,N_14746,N_14497);
or U14941 (N_14941,N_14709,N_14630);
and U14942 (N_14942,N_14494,N_14632);
or U14943 (N_14943,N_14638,N_14573);
nand U14944 (N_14944,N_14694,N_14519);
nand U14945 (N_14945,N_14756,N_14687);
xor U14946 (N_14946,N_14695,N_14579);
or U14947 (N_14947,N_14571,N_14778);
or U14948 (N_14948,N_14625,N_14460);
nand U14949 (N_14949,N_14558,N_14707);
or U14950 (N_14950,N_14411,N_14570);
or U14951 (N_14951,N_14423,N_14633);
nand U14952 (N_14952,N_14458,N_14730);
xnor U14953 (N_14953,N_14565,N_14786);
and U14954 (N_14954,N_14572,N_14463);
and U14955 (N_14955,N_14420,N_14770);
xnor U14956 (N_14956,N_14600,N_14434);
nand U14957 (N_14957,N_14703,N_14654);
xor U14958 (N_14958,N_14683,N_14668);
xnor U14959 (N_14959,N_14739,N_14699);
nand U14960 (N_14960,N_14526,N_14771);
nand U14961 (N_14961,N_14637,N_14611);
or U14962 (N_14962,N_14549,N_14443);
or U14963 (N_14963,N_14441,N_14763);
xor U14964 (N_14964,N_14609,N_14413);
nand U14965 (N_14965,N_14476,N_14563);
and U14966 (N_14966,N_14502,N_14692);
nand U14967 (N_14967,N_14498,N_14684);
or U14968 (N_14968,N_14612,N_14732);
xor U14969 (N_14969,N_14551,N_14752);
xor U14970 (N_14970,N_14671,N_14442);
nor U14971 (N_14971,N_14562,N_14605);
xnor U14972 (N_14972,N_14617,N_14762);
or U14973 (N_14973,N_14407,N_14575);
nand U14974 (N_14974,N_14528,N_14666);
xnor U14975 (N_14975,N_14663,N_14647);
or U14976 (N_14976,N_14453,N_14557);
xor U14977 (N_14977,N_14424,N_14468);
and U14978 (N_14978,N_14714,N_14469);
or U14979 (N_14979,N_14401,N_14406);
nor U14980 (N_14980,N_14435,N_14713);
and U14981 (N_14981,N_14412,N_14724);
or U14982 (N_14982,N_14791,N_14702);
nand U14983 (N_14983,N_14511,N_14520);
nor U14984 (N_14984,N_14629,N_14642);
xor U14985 (N_14985,N_14541,N_14799);
xnor U14986 (N_14986,N_14484,N_14461);
or U14987 (N_14987,N_14536,N_14620);
xor U14988 (N_14988,N_14583,N_14525);
or U14989 (N_14989,N_14587,N_14455);
nand U14990 (N_14990,N_14798,N_14795);
or U14991 (N_14991,N_14532,N_14431);
nor U14992 (N_14992,N_14772,N_14421);
xor U14993 (N_14993,N_14636,N_14643);
and U14994 (N_14994,N_14503,N_14725);
nor U14995 (N_14995,N_14728,N_14657);
and U14996 (N_14996,N_14561,N_14796);
nor U14997 (N_14997,N_14496,N_14492);
xor U14998 (N_14998,N_14417,N_14465);
or U14999 (N_14999,N_14501,N_14592);
nand U15000 (N_15000,N_14725,N_14489);
nor U15001 (N_15001,N_14432,N_14472);
nor U15002 (N_15002,N_14527,N_14500);
or U15003 (N_15003,N_14695,N_14559);
and U15004 (N_15004,N_14460,N_14786);
and U15005 (N_15005,N_14690,N_14616);
or U15006 (N_15006,N_14518,N_14613);
nor U15007 (N_15007,N_14744,N_14513);
nand U15008 (N_15008,N_14624,N_14788);
xor U15009 (N_15009,N_14653,N_14597);
nand U15010 (N_15010,N_14763,N_14781);
nand U15011 (N_15011,N_14515,N_14680);
or U15012 (N_15012,N_14536,N_14658);
or U15013 (N_15013,N_14586,N_14474);
or U15014 (N_15014,N_14773,N_14560);
xnor U15015 (N_15015,N_14691,N_14612);
and U15016 (N_15016,N_14576,N_14545);
or U15017 (N_15017,N_14430,N_14720);
xor U15018 (N_15018,N_14436,N_14478);
or U15019 (N_15019,N_14614,N_14608);
nand U15020 (N_15020,N_14672,N_14617);
xor U15021 (N_15021,N_14544,N_14431);
and U15022 (N_15022,N_14661,N_14570);
and U15023 (N_15023,N_14795,N_14731);
and U15024 (N_15024,N_14679,N_14401);
and U15025 (N_15025,N_14445,N_14413);
nor U15026 (N_15026,N_14715,N_14651);
and U15027 (N_15027,N_14473,N_14768);
xnor U15028 (N_15028,N_14643,N_14624);
nand U15029 (N_15029,N_14676,N_14604);
and U15030 (N_15030,N_14641,N_14631);
or U15031 (N_15031,N_14522,N_14524);
and U15032 (N_15032,N_14707,N_14647);
or U15033 (N_15033,N_14549,N_14770);
xnor U15034 (N_15034,N_14413,N_14776);
nor U15035 (N_15035,N_14760,N_14439);
xnor U15036 (N_15036,N_14441,N_14687);
and U15037 (N_15037,N_14772,N_14681);
and U15038 (N_15038,N_14534,N_14743);
and U15039 (N_15039,N_14661,N_14435);
xor U15040 (N_15040,N_14752,N_14404);
nand U15041 (N_15041,N_14665,N_14630);
and U15042 (N_15042,N_14617,N_14596);
nand U15043 (N_15043,N_14582,N_14489);
and U15044 (N_15044,N_14544,N_14405);
nand U15045 (N_15045,N_14611,N_14782);
nand U15046 (N_15046,N_14416,N_14624);
or U15047 (N_15047,N_14454,N_14726);
xor U15048 (N_15048,N_14753,N_14570);
or U15049 (N_15049,N_14692,N_14518);
and U15050 (N_15050,N_14589,N_14722);
or U15051 (N_15051,N_14401,N_14433);
xor U15052 (N_15052,N_14758,N_14630);
or U15053 (N_15053,N_14689,N_14788);
nor U15054 (N_15054,N_14751,N_14679);
xor U15055 (N_15055,N_14636,N_14525);
nor U15056 (N_15056,N_14582,N_14424);
or U15057 (N_15057,N_14532,N_14594);
nor U15058 (N_15058,N_14610,N_14404);
or U15059 (N_15059,N_14771,N_14779);
nand U15060 (N_15060,N_14689,N_14456);
xor U15061 (N_15061,N_14650,N_14754);
nand U15062 (N_15062,N_14438,N_14569);
or U15063 (N_15063,N_14674,N_14458);
nand U15064 (N_15064,N_14446,N_14546);
nor U15065 (N_15065,N_14579,N_14656);
xnor U15066 (N_15066,N_14469,N_14618);
xor U15067 (N_15067,N_14424,N_14612);
and U15068 (N_15068,N_14404,N_14650);
and U15069 (N_15069,N_14428,N_14792);
nand U15070 (N_15070,N_14408,N_14633);
xnor U15071 (N_15071,N_14777,N_14730);
xor U15072 (N_15072,N_14688,N_14790);
and U15073 (N_15073,N_14757,N_14477);
xor U15074 (N_15074,N_14628,N_14737);
or U15075 (N_15075,N_14544,N_14407);
nor U15076 (N_15076,N_14487,N_14550);
or U15077 (N_15077,N_14760,N_14791);
or U15078 (N_15078,N_14585,N_14461);
nand U15079 (N_15079,N_14652,N_14690);
xnor U15080 (N_15080,N_14786,N_14749);
xor U15081 (N_15081,N_14778,N_14400);
and U15082 (N_15082,N_14644,N_14499);
xor U15083 (N_15083,N_14640,N_14756);
or U15084 (N_15084,N_14415,N_14494);
nor U15085 (N_15085,N_14435,N_14574);
or U15086 (N_15086,N_14616,N_14546);
nor U15087 (N_15087,N_14549,N_14785);
nand U15088 (N_15088,N_14607,N_14741);
xnor U15089 (N_15089,N_14434,N_14495);
xor U15090 (N_15090,N_14670,N_14444);
nand U15091 (N_15091,N_14670,N_14497);
or U15092 (N_15092,N_14587,N_14581);
nand U15093 (N_15093,N_14713,N_14474);
and U15094 (N_15094,N_14646,N_14485);
nor U15095 (N_15095,N_14542,N_14700);
xnor U15096 (N_15096,N_14495,N_14596);
and U15097 (N_15097,N_14447,N_14494);
or U15098 (N_15098,N_14761,N_14428);
xor U15099 (N_15099,N_14691,N_14783);
xnor U15100 (N_15100,N_14514,N_14460);
or U15101 (N_15101,N_14765,N_14489);
nand U15102 (N_15102,N_14611,N_14569);
xor U15103 (N_15103,N_14766,N_14745);
or U15104 (N_15104,N_14529,N_14540);
nand U15105 (N_15105,N_14421,N_14488);
and U15106 (N_15106,N_14518,N_14439);
and U15107 (N_15107,N_14643,N_14743);
xnor U15108 (N_15108,N_14462,N_14638);
nor U15109 (N_15109,N_14787,N_14497);
nor U15110 (N_15110,N_14680,N_14766);
nand U15111 (N_15111,N_14728,N_14413);
nor U15112 (N_15112,N_14617,N_14472);
xor U15113 (N_15113,N_14527,N_14495);
or U15114 (N_15114,N_14422,N_14566);
nand U15115 (N_15115,N_14751,N_14724);
nand U15116 (N_15116,N_14711,N_14503);
nor U15117 (N_15117,N_14762,N_14451);
and U15118 (N_15118,N_14530,N_14461);
xnor U15119 (N_15119,N_14762,N_14755);
nand U15120 (N_15120,N_14504,N_14792);
nor U15121 (N_15121,N_14601,N_14612);
and U15122 (N_15122,N_14791,N_14507);
and U15123 (N_15123,N_14519,N_14784);
and U15124 (N_15124,N_14488,N_14593);
and U15125 (N_15125,N_14694,N_14587);
nor U15126 (N_15126,N_14568,N_14564);
nor U15127 (N_15127,N_14480,N_14496);
and U15128 (N_15128,N_14504,N_14614);
nor U15129 (N_15129,N_14776,N_14485);
or U15130 (N_15130,N_14594,N_14461);
xor U15131 (N_15131,N_14779,N_14461);
nor U15132 (N_15132,N_14766,N_14655);
nor U15133 (N_15133,N_14668,N_14718);
or U15134 (N_15134,N_14551,N_14558);
or U15135 (N_15135,N_14624,N_14503);
or U15136 (N_15136,N_14451,N_14606);
and U15137 (N_15137,N_14753,N_14410);
xor U15138 (N_15138,N_14411,N_14796);
nand U15139 (N_15139,N_14730,N_14539);
nand U15140 (N_15140,N_14699,N_14659);
xor U15141 (N_15141,N_14528,N_14789);
nor U15142 (N_15142,N_14477,N_14748);
or U15143 (N_15143,N_14783,N_14469);
xor U15144 (N_15144,N_14549,N_14425);
xnor U15145 (N_15145,N_14421,N_14658);
or U15146 (N_15146,N_14710,N_14707);
or U15147 (N_15147,N_14689,N_14501);
nor U15148 (N_15148,N_14439,N_14647);
or U15149 (N_15149,N_14619,N_14493);
and U15150 (N_15150,N_14573,N_14400);
xnor U15151 (N_15151,N_14764,N_14517);
and U15152 (N_15152,N_14726,N_14664);
xnor U15153 (N_15153,N_14630,N_14607);
and U15154 (N_15154,N_14672,N_14720);
nand U15155 (N_15155,N_14608,N_14644);
nor U15156 (N_15156,N_14636,N_14468);
and U15157 (N_15157,N_14788,N_14529);
nor U15158 (N_15158,N_14652,N_14656);
and U15159 (N_15159,N_14623,N_14446);
nand U15160 (N_15160,N_14710,N_14760);
nand U15161 (N_15161,N_14651,N_14406);
or U15162 (N_15162,N_14758,N_14410);
xnor U15163 (N_15163,N_14451,N_14622);
nand U15164 (N_15164,N_14660,N_14622);
and U15165 (N_15165,N_14764,N_14782);
and U15166 (N_15166,N_14615,N_14608);
nor U15167 (N_15167,N_14605,N_14669);
nand U15168 (N_15168,N_14517,N_14633);
nand U15169 (N_15169,N_14444,N_14739);
nor U15170 (N_15170,N_14478,N_14541);
xnor U15171 (N_15171,N_14605,N_14500);
xnor U15172 (N_15172,N_14620,N_14665);
or U15173 (N_15173,N_14409,N_14642);
nor U15174 (N_15174,N_14428,N_14600);
or U15175 (N_15175,N_14440,N_14653);
or U15176 (N_15176,N_14569,N_14527);
nor U15177 (N_15177,N_14501,N_14696);
xor U15178 (N_15178,N_14461,N_14465);
nand U15179 (N_15179,N_14482,N_14600);
nand U15180 (N_15180,N_14501,N_14768);
and U15181 (N_15181,N_14704,N_14555);
and U15182 (N_15182,N_14558,N_14442);
and U15183 (N_15183,N_14772,N_14409);
and U15184 (N_15184,N_14559,N_14457);
or U15185 (N_15185,N_14765,N_14672);
and U15186 (N_15186,N_14731,N_14509);
or U15187 (N_15187,N_14493,N_14703);
xor U15188 (N_15188,N_14798,N_14562);
and U15189 (N_15189,N_14565,N_14408);
xnor U15190 (N_15190,N_14739,N_14628);
nor U15191 (N_15191,N_14653,N_14532);
xnor U15192 (N_15192,N_14432,N_14485);
nand U15193 (N_15193,N_14462,N_14696);
or U15194 (N_15194,N_14669,N_14760);
nor U15195 (N_15195,N_14465,N_14720);
or U15196 (N_15196,N_14479,N_14561);
nor U15197 (N_15197,N_14492,N_14418);
and U15198 (N_15198,N_14529,N_14618);
nand U15199 (N_15199,N_14547,N_14716);
nor U15200 (N_15200,N_14911,N_15180);
or U15201 (N_15201,N_14804,N_14909);
nand U15202 (N_15202,N_14940,N_14918);
nor U15203 (N_15203,N_15065,N_15111);
nand U15204 (N_15204,N_15027,N_15073);
or U15205 (N_15205,N_15183,N_14974);
nand U15206 (N_15206,N_15179,N_15174);
xor U15207 (N_15207,N_15165,N_14817);
nand U15208 (N_15208,N_14815,N_14941);
xor U15209 (N_15209,N_14982,N_14973);
nor U15210 (N_15210,N_14845,N_14983);
nor U15211 (N_15211,N_14829,N_14824);
xor U15212 (N_15212,N_14871,N_15006);
or U15213 (N_15213,N_14931,N_14981);
and U15214 (N_15214,N_15169,N_15019);
nand U15215 (N_15215,N_15177,N_14843);
nand U15216 (N_15216,N_15157,N_15123);
and U15217 (N_15217,N_14830,N_14886);
nor U15218 (N_15218,N_14863,N_15154);
and U15219 (N_15219,N_15124,N_15029);
nand U15220 (N_15220,N_15064,N_15198);
nand U15221 (N_15221,N_15148,N_15127);
nor U15222 (N_15222,N_14857,N_14809);
nand U15223 (N_15223,N_15066,N_15038);
nand U15224 (N_15224,N_15057,N_15094);
and U15225 (N_15225,N_15014,N_14938);
nor U15226 (N_15226,N_14903,N_15004);
xnor U15227 (N_15227,N_15086,N_15101);
nand U15228 (N_15228,N_15055,N_14884);
nor U15229 (N_15229,N_14963,N_15125);
xnor U15230 (N_15230,N_15001,N_15097);
xor U15231 (N_15231,N_15095,N_15079);
or U15232 (N_15232,N_15056,N_14870);
and U15233 (N_15233,N_15035,N_15092);
and U15234 (N_15234,N_15051,N_15189);
xnor U15235 (N_15235,N_14842,N_14819);
or U15236 (N_15236,N_15159,N_15085);
and U15237 (N_15237,N_15025,N_15196);
or U15238 (N_15238,N_14885,N_15145);
nor U15239 (N_15239,N_15175,N_15090);
nand U15240 (N_15240,N_14822,N_15089);
or U15241 (N_15241,N_15146,N_15068);
nand U15242 (N_15242,N_15100,N_14896);
or U15243 (N_15243,N_14844,N_14979);
or U15244 (N_15244,N_15043,N_15067);
nand U15245 (N_15245,N_14808,N_15144);
or U15246 (N_15246,N_15153,N_14917);
nor U15247 (N_15247,N_14860,N_14943);
xnor U15248 (N_15248,N_14953,N_15039);
and U15249 (N_15249,N_14801,N_14855);
nor U15250 (N_15250,N_14881,N_15131);
and U15251 (N_15251,N_14991,N_14806);
xnor U15252 (N_15252,N_14897,N_15077);
or U15253 (N_15253,N_14948,N_15063);
xnor U15254 (N_15254,N_14840,N_15115);
or U15255 (N_15255,N_14847,N_14805);
and U15256 (N_15256,N_14978,N_15186);
or U15257 (N_15257,N_15072,N_14828);
xnor U15258 (N_15258,N_15158,N_14852);
nor U15259 (N_15259,N_14971,N_15133);
or U15260 (N_15260,N_14803,N_15190);
nor U15261 (N_15261,N_14949,N_14883);
and U15262 (N_15262,N_14825,N_15110);
or U15263 (N_15263,N_15060,N_15135);
xnor U15264 (N_15264,N_15136,N_14950);
and U15265 (N_15265,N_14928,N_15098);
nand U15266 (N_15266,N_15023,N_15058);
nor U15267 (N_15267,N_14891,N_15096);
or U15268 (N_15268,N_15137,N_14932);
xor U15269 (N_15269,N_14868,N_15181);
or U15270 (N_15270,N_14838,N_15160);
nor U15271 (N_15271,N_14814,N_15193);
nand U15272 (N_15272,N_15061,N_14962);
xnor U15273 (N_15273,N_14858,N_15112);
or U15274 (N_15274,N_15173,N_15026);
nand U15275 (N_15275,N_14929,N_14992);
xnor U15276 (N_15276,N_14901,N_15007);
and U15277 (N_15277,N_14837,N_15191);
and U15278 (N_15278,N_15031,N_15088);
nor U15279 (N_15279,N_15016,N_14894);
nand U15280 (N_15280,N_15132,N_15069);
nor U15281 (N_15281,N_14807,N_14997);
nor U15282 (N_15282,N_14960,N_15184);
and U15283 (N_15283,N_14937,N_15104);
or U15284 (N_15284,N_14914,N_15082);
and U15285 (N_15285,N_14827,N_14985);
or U15286 (N_15286,N_14998,N_14867);
nor U15287 (N_15287,N_15120,N_14966);
nor U15288 (N_15288,N_14935,N_14873);
nor U15289 (N_15289,N_15099,N_15114);
and U15290 (N_15290,N_15046,N_14878);
and U15291 (N_15291,N_15113,N_14802);
xnor U15292 (N_15292,N_15167,N_15045);
nor U15293 (N_15293,N_15109,N_15134);
and U15294 (N_15294,N_15117,N_14812);
nor U15295 (N_15295,N_15149,N_15192);
nor U15296 (N_15296,N_14899,N_15147);
xnor U15297 (N_15297,N_15053,N_14965);
xor U15298 (N_15298,N_14924,N_14848);
and U15299 (N_15299,N_15141,N_15034);
and U15300 (N_15300,N_14995,N_15024);
xor U15301 (N_15301,N_15076,N_15152);
nand U15302 (N_15302,N_14993,N_15021);
xor U15303 (N_15303,N_14826,N_14839);
nand U15304 (N_15304,N_14864,N_14926);
or U15305 (N_15305,N_14850,N_14919);
xnor U15306 (N_15306,N_14927,N_14916);
xor U15307 (N_15307,N_14984,N_14930);
or U15308 (N_15308,N_14913,N_15170);
nand U15309 (N_15309,N_14853,N_14975);
nor U15310 (N_15310,N_14972,N_15008);
nor U15311 (N_15311,N_15126,N_14970);
and U15312 (N_15312,N_14862,N_15071);
xnor U15313 (N_15313,N_14936,N_14811);
or U15314 (N_15314,N_14813,N_15017);
xor U15315 (N_15315,N_14831,N_15005);
nand U15316 (N_15316,N_14958,N_15059);
nor U15317 (N_15317,N_14922,N_14951);
or U15318 (N_15318,N_15163,N_15050);
xor U15319 (N_15319,N_15028,N_14920);
and U15320 (N_15320,N_15033,N_15140);
nand U15321 (N_15321,N_14959,N_14989);
nor U15322 (N_15322,N_14942,N_15168);
nor U15323 (N_15323,N_14835,N_15030);
nand U15324 (N_15324,N_15128,N_14818);
or U15325 (N_15325,N_14976,N_15062);
nor U15326 (N_15326,N_14890,N_15102);
nor U15327 (N_15327,N_15000,N_15003);
xnor U15328 (N_15328,N_15182,N_15103);
nand U15329 (N_15329,N_15074,N_14908);
or U15330 (N_15330,N_14882,N_15199);
nand U15331 (N_15331,N_14833,N_15121);
nor U15332 (N_15332,N_14956,N_15078);
or U15333 (N_15333,N_14872,N_14969);
and U15334 (N_15334,N_15195,N_15129);
and U15335 (N_15335,N_14880,N_14987);
and U15336 (N_15336,N_14925,N_15036);
and U15337 (N_15337,N_14820,N_15042);
and U15338 (N_15338,N_15171,N_14980);
nand U15339 (N_15339,N_14877,N_14810);
nand U15340 (N_15340,N_14907,N_15084);
nand U15341 (N_15341,N_15009,N_14921);
nand U15342 (N_15342,N_15047,N_14892);
xnor U15343 (N_15343,N_14898,N_15164);
nand U15344 (N_15344,N_15138,N_14947);
and U15345 (N_15345,N_15178,N_15176);
nor U15346 (N_15346,N_14866,N_15162);
nor U15347 (N_15347,N_14996,N_15093);
and U15348 (N_15348,N_14889,N_14954);
nor U15349 (N_15349,N_15048,N_14952);
xor U15350 (N_15350,N_15156,N_14967);
and U15351 (N_15351,N_14854,N_15037);
and U15352 (N_15352,N_14994,N_14836);
xor U15353 (N_15353,N_14887,N_14939);
or U15354 (N_15354,N_14841,N_14800);
and U15355 (N_15355,N_15049,N_14879);
and U15356 (N_15356,N_14902,N_14816);
and U15357 (N_15357,N_14888,N_14861);
xnor U15358 (N_15358,N_15015,N_14874);
xor U15359 (N_15359,N_14933,N_14968);
nand U15360 (N_15360,N_15012,N_14955);
and U15361 (N_15361,N_14869,N_15166);
or U15362 (N_15362,N_15130,N_15081);
and U15363 (N_15363,N_15022,N_15013);
xor U15364 (N_15364,N_15143,N_15032);
or U15365 (N_15365,N_14904,N_15187);
xor U15366 (N_15366,N_14876,N_14946);
and U15367 (N_15367,N_15052,N_14999);
nor U15368 (N_15368,N_14923,N_14912);
and U15369 (N_15369,N_14900,N_15151);
and U15370 (N_15370,N_15188,N_14893);
nand U15371 (N_15371,N_15106,N_14895);
or U15372 (N_15372,N_14859,N_15194);
and U15373 (N_15373,N_14957,N_14851);
or U15374 (N_15374,N_14945,N_15139);
nor U15375 (N_15375,N_14910,N_14849);
xnor U15376 (N_15376,N_14856,N_15197);
and U15377 (N_15377,N_15161,N_14905);
nand U15378 (N_15378,N_14986,N_14915);
and U15379 (N_15379,N_15010,N_14823);
xnor U15380 (N_15380,N_14990,N_15105);
xnor U15381 (N_15381,N_15080,N_15185);
or U15382 (N_15382,N_15087,N_14977);
nand U15383 (N_15383,N_15041,N_14834);
or U15384 (N_15384,N_15116,N_15091);
nand U15385 (N_15385,N_15108,N_15040);
nor U15386 (N_15386,N_15075,N_14832);
nor U15387 (N_15387,N_15172,N_14906);
xor U15388 (N_15388,N_14875,N_15118);
nor U15389 (N_15389,N_15018,N_15044);
or U15390 (N_15390,N_15150,N_14821);
nor U15391 (N_15391,N_15020,N_14988);
and U15392 (N_15392,N_14964,N_14961);
and U15393 (N_15393,N_15002,N_15070);
or U15394 (N_15394,N_15142,N_15122);
and U15395 (N_15395,N_15083,N_15119);
or U15396 (N_15396,N_14865,N_14934);
and U15397 (N_15397,N_14846,N_14944);
or U15398 (N_15398,N_15054,N_15107);
nor U15399 (N_15399,N_15011,N_15155);
or U15400 (N_15400,N_14881,N_15157);
and U15401 (N_15401,N_14801,N_15091);
nand U15402 (N_15402,N_14956,N_15023);
nand U15403 (N_15403,N_15117,N_14880);
nand U15404 (N_15404,N_15089,N_14876);
and U15405 (N_15405,N_14965,N_14892);
and U15406 (N_15406,N_14950,N_15146);
nor U15407 (N_15407,N_15088,N_15108);
nor U15408 (N_15408,N_15180,N_15100);
or U15409 (N_15409,N_15086,N_15010);
nor U15410 (N_15410,N_14857,N_15004);
nor U15411 (N_15411,N_15142,N_14865);
nor U15412 (N_15412,N_14923,N_14865);
nor U15413 (N_15413,N_14998,N_14918);
or U15414 (N_15414,N_15096,N_14909);
nand U15415 (N_15415,N_15127,N_14845);
nor U15416 (N_15416,N_14901,N_15076);
xnor U15417 (N_15417,N_15138,N_15105);
or U15418 (N_15418,N_15191,N_14971);
or U15419 (N_15419,N_15190,N_15096);
nand U15420 (N_15420,N_14978,N_15060);
and U15421 (N_15421,N_14820,N_14951);
and U15422 (N_15422,N_15147,N_14866);
and U15423 (N_15423,N_14859,N_14953);
or U15424 (N_15424,N_14896,N_14970);
nor U15425 (N_15425,N_14916,N_14885);
nand U15426 (N_15426,N_14960,N_14918);
nor U15427 (N_15427,N_15156,N_14868);
nor U15428 (N_15428,N_14910,N_14962);
and U15429 (N_15429,N_14971,N_14912);
or U15430 (N_15430,N_15094,N_15039);
nor U15431 (N_15431,N_15044,N_15036);
nor U15432 (N_15432,N_15142,N_15061);
nor U15433 (N_15433,N_14966,N_15102);
and U15434 (N_15434,N_14979,N_14994);
or U15435 (N_15435,N_15161,N_15123);
nand U15436 (N_15436,N_15125,N_15044);
or U15437 (N_15437,N_14898,N_15113);
nand U15438 (N_15438,N_15106,N_15120);
and U15439 (N_15439,N_15027,N_15001);
nor U15440 (N_15440,N_14935,N_14844);
xnor U15441 (N_15441,N_14875,N_15040);
xnor U15442 (N_15442,N_15022,N_14965);
nor U15443 (N_15443,N_14973,N_15196);
nand U15444 (N_15444,N_15115,N_14849);
or U15445 (N_15445,N_15037,N_15060);
xnor U15446 (N_15446,N_15193,N_14951);
nor U15447 (N_15447,N_15040,N_14827);
or U15448 (N_15448,N_15187,N_14811);
and U15449 (N_15449,N_14928,N_15126);
xnor U15450 (N_15450,N_15037,N_15021);
nand U15451 (N_15451,N_15036,N_14992);
nand U15452 (N_15452,N_14824,N_14889);
or U15453 (N_15453,N_15074,N_14866);
and U15454 (N_15454,N_14990,N_14958);
and U15455 (N_15455,N_14941,N_15064);
xor U15456 (N_15456,N_15016,N_14907);
and U15457 (N_15457,N_15051,N_14914);
and U15458 (N_15458,N_14816,N_15113);
or U15459 (N_15459,N_14876,N_15060);
nand U15460 (N_15460,N_15029,N_14835);
nor U15461 (N_15461,N_14980,N_14941);
or U15462 (N_15462,N_14859,N_15096);
nor U15463 (N_15463,N_14914,N_15098);
or U15464 (N_15464,N_15184,N_14981);
nand U15465 (N_15465,N_14827,N_14981);
nor U15466 (N_15466,N_15164,N_15121);
nor U15467 (N_15467,N_15048,N_15098);
or U15468 (N_15468,N_14816,N_15121);
nor U15469 (N_15469,N_14801,N_14908);
and U15470 (N_15470,N_15057,N_14818);
and U15471 (N_15471,N_14812,N_15077);
xnor U15472 (N_15472,N_14824,N_14874);
nor U15473 (N_15473,N_14954,N_14985);
xor U15474 (N_15474,N_15075,N_15100);
and U15475 (N_15475,N_15091,N_14996);
xnor U15476 (N_15476,N_15127,N_14971);
nor U15477 (N_15477,N_14981,N_14870);
or U15478 (N_15478,N_14937,N_14909);
xor U15479 (N_15479,N_14891,N_15113);
nand U15480 (N_15480,N_15020,N_15115);
or U15481 (N_15481,N_15036,N_14920);
nor U15482 (N_15482,N_14805,N_14824);
xor U15483 (N_15483,N_15055,N_15094);
and U15484 (N_15484,N_14927,N_14972);
xor U15485 (N_15485,N_15124,N_14858);
nor U15486 (N_15486,N_15140,N_15030);
and U15487 (N_15487,N_15085,N_15100);
nor U15488 (N_15488,N_15106,N_15037);
or U15489 (N_15489,N_14984,N_15043);
or U15490 (N_15490,N_15123,N_14935);
xnor U15491 (N_15491,N_15121,N_15045);
or U15492 (N_15492,N_14928,N_15071);
nor U15493 (N_15493,N_15039,N_15098);
nand U15494 (N_15494,N_14803,N_15018);
nand U15495 (N_15495,N_14962,N_15053);
xnor U15496 (N_15496,N_15168,N_14876);
xnor U15497 (N_15497,N_14916,N_14868);
xor U15498 (N_15498,N_15106,N_14861);
xnor U15499 (N_15499,N_15049,N_15024);
and U15500 (N_15500,N_15022,N_14880);
and U15501 (N_15501,N_15077,N_14953);
or U15502 (N_15502,N_15035,N_15041);
and U15503 (N_15503,N_14842,N_15023);
nand U15504 (N_15504,N_15072,N_14807);
nor U15505 (N_15505,N_14845,N_14935);
xnor U15506 (N_15506,N_15070,N_14886);
xor U15507 (N_15507,N_15129,N_14914);
or U15508 (N_15508,N_14827,N_15095);
and U15509 (N_15509,N_14898,N_15152);
xor U15510 (N_15510,N_14902,N_14881);
or U15511 (N_15511,N_14813,N_15081);
and U15512 (N_15512,N_14851,N_15147);
nand U15513 (N_15513,N_15118,N_15061);
and U15514 (N_15514,N_14970,N_15049);
or U15515 (N_15515,N_15173,N_14901);
xnor U15516 (N_15516,N_14979,N_14901);
and U15517 (N_15517,N_15048,N_14940);
or U15518 (N_15518,N_15147,N_15158);
and U15519 (N_15519,N_14929,N_15131);
and U15520 (N_15520,N_15131,N_14806);
nor U15521 (N_15521,N_14868,N_14955);
or U15522 (N_15522,N_15074,N_14876);
nand U15523 (N_15523,N_14849,N_14975);
and U15524 (N_15524,N_15010,N_15171);
nor U15525 (N_15525,N_15192,N_15031);
nand U15526 (N_15526,N_15101,N_15116);
and U15527 (N_15527,N_15070,N_14924);
xnor U15528 (N_15528,N_14842,N_15107);
xnor U15529 (N_15529,N_15149,N_14894);
xnor U15530 (N_15530,N_15076,N_15050);
nor U15531 (N_15531,N_15110,N_15080);
nor U15532 (N_15532,N_15140,N_14839);
nand U15533 (N_15533,N_14948,N_15057);
xor U15534 (N_15534,N_15003,N_14977);
and U15535 (N_15535,N_14880,N_14816);
or U15536 (N_15536,N_14827,N_14967);
xnor U15537 (N_15537,N_14976,N_15127);
nand U15538 (N_15538,N_14901,N_15088);
xnor U15539 (N_15539,N_15053,N_14859);
and U15540 (N_15540,N_14841,N_15009);
nand U15541 (N_15541,N_15086,N_15025);
xor U15542 (N_15542,N_14938,N_14986);
or U15543 (N_15543,N_14859,N_14825);
nor U15544 (N_15544,N_15063,N_15074);
xnor U15545 (N_15545,N_14890,N_14884);
xor U15546 (N_15546,N_15009,N_15176);
nor U15547 (N_15547,N_14910,N_15087);
xor U15548 (N_15548,N_15176,N_15139);
nor U15549 (N_15549,N_14959,N_14871);
or U15550 (N_15550,N_15061,N_15164);
nor U15551 (N_15551,N_15010,N_15057);
nand U15552 (N_15552,N_14923,N_14854);
xnor U15553 (N_15553,N_14905,N_15123);
nand U15554 (N_15554,N_14896,N_14829);
nand U15555 (N_15555,N_14964,N_15057);
xnor U15556 (N_15556,N_14825,N_14915);
or U15557 (N_15557,N_14947,N_14994);
nand U15558 (N_15558,N_15137,N_15140);
and U15559 (N_15559,N_15188,N_15054);
nor U15560 (N_15560,N_15024,N_15186);
or U15561 (N_15561,N_14916,N_14802);
nor U15562 (N_15562,N_14822,N_15019);
and U15563 (N_15563,N_14947,N_14800);
xor U15564 (N_15564,N_15028,N_15136);
or U15565 (N_15565,N_14835,N_15127);
and U15566 (N_15566,N_14851,N_15055);
and U15567 (N_15567,N_14856,N_15132);
and U15568 (N_15568,N_14840,N_14978);
and U15569 (N_15569,N_14986,N_15173);
or U15570 (N_15570,N_14907,N_14970);
or U15571 (N_15571,N_14935,N_15073);
nand U15572 (N_15572,N_15156,N_15196);
nor U15573 (N_15573,N_15123,N_15146);
and U15574 (N_15574,N_14823,N_15064);
xor U15575 (N_15575,N_14920,N_15076);
or U15576 (N_15576,N_14894,N_14995);
nor U15577 (N_15577,N_14869,N_14914);
and U15578 (N_15578,N_15105,N_14919);
and U15579 (N_15579,N_14892,N_14983);
xnor U15580 (N_15580,N_14852,N_15070);
nor U15581 (N_15581,N_15075,N_14878);
xnor U15582 (N_15582,N_15118,N_15045);
nand U15583 (N_15583,N_15079,N_15110);
nor U15584 (N_15584,N_14914,N_14987);
nor U15585 (N_15585,N_15036,N_15195);
nor U15586 (N_15586,N_14898,N_15006);
xnor U15587 (N_15587,N_15198,N_15110);
nand U15588 (N_15588,N_14863,N_15105);
nor U15589 (N_15589,N_14959,N_14860);
nand U15590 (N_15590,N_14945,N_14973);
nand U15591 (N_15591,N_15031,N_14973);
xnor U15592 (N_15592,N_14831,N_14911);
nand U15593 (N_15593,N_14861,N_15131);
nor U15594 (N_15594,N_14848,N_14887);
and U15595 (N_15595,N_14872,N_15049);
nor U15596 (N_15596,N_14836,N_15162);
xnor U15597 (N_15597,N_15080,N_15170);
or U15598 (N_15598,N_14904,N_14968);
xor U15599 (N_15599,N_14897,N_14808);
nor U15600 (N_15600,N_15588,N_15400);
or U15601 (N_15601,N_15460,N_15562);
nand U15602 (N_15602,N_15315,N_15571);
or U15603 (N_15603,N_15260,N_15323);
nand U15604 (N_15604,N_15381,N_15222);
or U15605 (N_15605,N_15259,N_15499);
nor U15606 (N_15606,N_15268,N_15475);
nand U15607 (N_15607,N_15547,N_15577);
and U15608 (N_15608,N_15466,N_15566);
xor U15609 (N_15609,N_15580,N_15212);
nor U15610 (N_15610,N_15354,N_15204);
nor U15611 (N_15611,N_15350,N_15399);
nand U15612 (N_15612,N_15373,N_15385);
nand U15613 (N_15613,N_15532,N_15286);
xor U15614 (N_15614,N_15255,N_15575);
nand U15615 (N_15615,N_15447,N_15213);
xor U15616 (N_15616,N_15491,N_15342);
nand U15617 (N_15617,N_15244,N_15257);
nand U15618 (N_15618,N_15250,N_15567);
and U15619 (N_15619,N_15390,N_15296);
or U15620 (N_15620,N_15359,N_15589);
or U15621 (N_15621,N_15336,N_15526);
and U15622 (N_15622,N_15308,N_15267);
nor U15623 (N_15623,N_15574,N_15576);
nand U15624 (N_15624,N_15496,N_15481);
xor U15625 (N_15625,N_15539,N_15507);
xnor U15626 (N_15626,N_15572,N_15472);
nand U15627 (N_15627,N_15500,N_15553);
nor U15628 (N_15628,N_15469,N_15289);
or U15629 (N_15629,N_15455,N_15549);
and U15630 (N_15630,N_15263,N_15420);
and U15631 (N_15631,N_15464,N_15211);
and U15632 (N_15632,N_15246,N_15595);
nor U15633 (N_15633,N_15265,N_15438);
nand U15634 (N_15634,N_15531,N_15295);
xor U15635 (N_15635,N_15482,N_15473);
xnor U15636 (N_15636,N_15243,N_15306);
and U15637 (N_15637,N_15486,N_15294);
nand U15638 (N_15638,N_15396,N_15559);
and U15639 (N_15639,N_15565,N_15224);
nor U15640 (N_15640,N_15210,N_15394);
or U15641 (N_15641,N_15517,N_15449);
or U15642 (N_15642,N_15388,N_15584);
nand U15643 (N_15643,N_15330,N_15377);
or U15644 (N_15644,N_15581,N_15280);
xnor U15645 (N_15645,N_15546,N_15261);
nor U15646 (N_15646,N_15374,N_15321);
nor U15647 (N_15647,N_15439,N_15226);
or U15648 (N_15648,N_15483,N_15535);
nand U15649 (N_15649,N_15587,N_15533);
and U15650 (N_15650,N_15470,N_15578);
and U15651 (N_15651,N_15326,N_15441);
or U15652 (N_15652,N_15314,N_15348);
or U15653 (N_15653,N_15242,N_15521);
and U15654 (N_15654,N_15407,N_15415);
nor U15655 (N_15655,N_15510,N_15492);
or U15656 (N_15656,N_15442,N_15513);
or U15657 (N_15657,N_15231,N_15304);
nand U15658 (N_15658,N_15298,N_15346);
and U15659 (N_15659,N_15356,N_15252);
nor U15660 (N_15660,N_15555,N_15471);
xnor U15661 (N_15661,N_15520,N_15506);
nand U15662 (N_15662,N_15456,N_15542);
or U15663 (N_15663,N_15287,N_15347);
nand U15664 (N_15664,N_15364,N_15380);
nand U15665 (N_15665,N_15508,N_15525);
nor U15666 (N_15666,N_15227,N_15239);
nor U15667 (N_15667,N_15215,N_15479);
or U15668 (N_15668,N_15556,N_15230);
or U15669 (N_15669,N_15349,N_15540);
nor U15670 (N_15670,N_15568,N_15478);
xor U15671 (N_15671,N_15233,N_15344);
nor U15672 (N_15672,N_15550,N_15480);
or U15673 (N_15673,N_15220,N_15214);
and U15674 (N_15674,N_15545,N_15262);
and U15675 (N_15675,N_15427,N_15530);
xnor U15676 (N_15676,N_15573,N_15335);
nor U15677 (N_15677,N_15319,N_15487);
or U15678 (N_15678,N_15461,N_15237);
and U15679 (N_15679,N_15276,N_15516);
nor U15680 (N_15680,N_15279,N_15452);
xor U15681 (N_15681,N_15376,N_15217);
and U15682 (N_15682,N_15372,N_15256);
nor U15683 (N_15683,N_15503,N_15501);
xnor U15684 (N_15684,N_15544,N_15241);
nor U15685 (N_15685,N_15218,N_15435);
nand U15686 (N_15686,N_15412,N_15369);
nand U15687 (N_15687,N_15254,N_15292);
nor U15688 (N_15688,N_15311,N_15351);
or U15689 (N_15689,N_15291,N_15317);
xor U15690 (N_15690,N_15225,N_15368);
xnor U15691 (N_15691,N_15277,N_15320);
or U15692 (N_15692,N_15322,N_15375);
xor U15693 (N_15693,N_15303,N_15552);
and U15694 (N_15694,N_15465,N_15301);
and U15695 (N_15695,N_15596,N_15493);
xor U15696 (N_15696,N_15309,N_15383);
xor U15697 (N_15697,N_15305,N_15258);
nor U15698 (N_15698,N_15561,N_15272);
or U15699 (N_15699,N_15490,N_15515);
or U15700 (N_15700,N_15458,N_15467);
and U15701 (N_15701,N_15509,N_15201);
or U15702 (N_15702,N_15504,N_15564);
xor U15703 (N_15703,N_15360,N_15583);
or U15704 (N_15704,N_15457,N_15297);
xnor U15705 (N_15705,N_15398,N_15590);
nor U15706 (N_15706,N_15269,N_15451);
xor U15707 (N_15707,N_15270,N_15430);
nand U15708 (N_15708,N_15426,N_15238);
and U15709 (N_15709,N_15423,N_15382);
and U15710 (N_15710,N_15299,N_15312);
and U15711 (N_15711,N_15236,N_15463);
and U15712 (N_15712,N_15433,N_15599);
nand U15713 (N_15713,N_15207,N_15389);
or U15714 (N_15714,N_15440,N_15477);
nand U15715 (N_15715,N_15489,N_15307);
nor U15716 (N_15716,N_15485,N_15205);
or U15717 (N_15717,N_15448,N_15318);
xnor U15718 (N_15718,N_15411,N_15512);
or U15719 (N_15719,N_15536,N_15444);
or U15720 (N_15720,N_15332,N_15221);
xnor U15721 (N_15721,N_15245,N_15534);
nor U15722 (N_15722,N_15402,N_15325);
xnor U15723 (N_15723,N_15410,N_15216);
nor U15724 (N_15724,N_15484,N_15497);
and U15725 (N_15725,N_15345,N_15251);
nor U15726 (N_15726,N_15288,N_15570);
and U15727 (N_15727,N_15229,N_15431);
nor U15728 (N_15728,N_15502,N_15284);
or U15729 (N_15729,N_15274,N_15392);
nand U15730 (N_15730,N_15537,N_15264);
nor U15731 (N_15731,N_15505,N_15495);
or U15732 (N_15732,N_15313,N_15579);
xnor U15733 (N_15733,N_15408,N_15355);
and U15734 (N_15734,N_15202,N_15476);
nand U15735 (N_15735,N_15582,N_15391);
nor U15736 (N_15736,N_15593,N_15340);
and U15737 (N_15737,N_15428,N_15529);
nand U15738 (N_15738,N_15334,N_15232);
xnor U15739 (N_15739,N_15324,N_15454);
and U15740 (N_15740,N_15271,N_15453);
or U15741 (N_15741,N_15560,N_15591);
and U15742 (N_15742,N_15524,N_15331);
nor U15743 (N_15743,N_15366,N_15538);
or U15744 (N_15744,N_15585,N_15234);
nor U15745 (N_15745,N_15597,N_15518);
and U15746 (N_15746,N_15365,N_15594);
nor U15747 (N_15747,N_15522,N_15275);
xor U15748 (N_15748,N_15337,N_15450);
nand U15749 (N_15749,N_15290,N_15253);
nand U15750 (N_15750,N_15511,N_15371);
and U15751 (N_15751,N_15406,N_15300);
nand U15752 (N_15752,N_15551,N_15362);
and U15753 (N_15753,N_15498,N_15425);
and U15754 (N_15754,N_15341,N_15434);
xor U15755 (N_15755,N_15240,N_15378);
xnor U15756 (N_15756,N_15266,N_15282);
nand U15757 (N_15757,N_15586,N_15327);
xnor U15758 (N_15758,N_15554,N_15384);
and U15759 (N_15759,N_15247,N_15249);
and U15760 (N_15760,N_15569,N_15548);
nor U15761 (N_15761,N_15333,N_15543);
nand U15762 (N_15762,N_15357,N_15413);
xnor U15763 (N_15763,N_15417,N_15446);
nor U15764 (N_15764,N_15203,N_15393);
and U15765 (N_15765,N_15528,N_15310);
nor U15766 (N_15766,N_15403,N_15285);
xor U15767 (N_15767,N_15283,N_15443);
or U15768 (N_15768,N_15592,N_15361);
and U15769 (N_15769,N_15401,N_15273);
xnor U15770 (N_15770,N_15459,N_15278);
and U15771 (N_15771,N_15462,N_15387);
and U15772 (N_15772,N_15209,N_15405);
nand U15773 (N_15773,N_15421,N_15302);
and U15774 (N_15774,N_15424,N_15558);
nor U15775 (N_15775,N_15409,N_15206);
or U15776 (N_15776,N_15370,N_15557);
and U15777 (N_15777,N_15363,N_15386);
nand U15778 (N_15778,N_15598,N_15248);
and U15779 (N_15779,N_15432,N_15367);
nor U15780 (N_15780,N_15328,N_15563);
xor U15781 (N_15781,N_15416,N_15414);
and U15782 (N_15782,N_15488,N_15219);
and U15783 (N_15783,N_15293,N_15339);
xnor U15784 (N_15784,N_15235,N_15468);
nor U15785 (N_15785,N_15379,N_15358);
nor U15786 (N_15786,N_15541,N_15223);
and U15787 (N_15787,N_15343,N_15494);
xnor U15788 (N_15788,N_15397,N_15404);
and U15789 (N_15789,N_15395,N_15228);
nand U15790 (N_15790,N_15474,N_15419);
nand U15791 (N_15791,N_15352,N_15338);
xnor U15792 (N_15792,N_15436,N_15316);
xnor U15793 (N_15793,N_15200,N_15281);
nand U15794 (N_15794,N_15527,N_15437);
nor U15795 (N_15795,N_15429,N_15418);
xnor U15796 (N_15796,N_15353,N_15445);
xnor U15797 (N_15797,N_15523,N_15519);
nand U15798 (N_15798,N_15329,N_15208);
and U15799 (N_15799,N_15514,N_15422);
and U15800 (N_15800,N_15514,N_15487);
nand U15801 (N_15801,N_15590,N_15530);
and U15802 (N_15802,N_15559,N_15599);
and U15803 (N_15803,N_15479,N_15524);
xnor U15804 (N_15804,N_15254,N_15473);
or U15805 (N_15805,N_15325,N_15263);
and U15806 (N_15806,N_15388,N_15323);
or U15807 (N_15807,N_15386,N_15553);
xnor U15808 (N_15808,N_15209,N_15444);
nor U15809 (N_15809,N_15445,N_15438);
and U15810 (N_15810,N_15293,N_15263);
and U15811 (N_15811,N_15434,N_15311);
nand U15812 (N_15812,N_15358,N_15437);
nor U15813 (N_15813,N_15539,N_15535);
xnor U15814 (N_15814,N_15392,N_15382);
nor U15815 (N_15815,N_15321,N_15205);
nand U15816 (N_15816,N_15304,N_15536);
nor U15817 (N_15817,N_15578,N_15215);
nand U15818 (N_15818,N_15462,N_15385);
xnor U15819 (N_15819,N_15358,N_15545);
or U15820 (N_15820,N_15238,N_15279);
nand U15821 (N_15821,N_15430,N_15284);
nand U15822 (N_15822,N_15279,N_15451);
or U15823 (N_15823,N_15401,N_15344);
nand U15824 (N_15824,N_15571,N_15595);
xnor U15825 (N_15825,N_15227,N_15574);
or U15826 (N_15826,N_15442,N_15361);
nand U15827 (N_15827,N_15272,N_15576);
nor U15828 (N_15828,N_15280,N_15566);
or U15829 (N_15829,N_15348,N_15269);
xnor U15830 (N_15830,N_15351,N_15314);
or U15831 (N_15831,N_15362,N_15392);
or U15832 (N_15832,N_15378,N_15583);
or U15833 (N_15833,N_15272,N_15398);
xor U15834 (N_15834,N_15258,N_15587);
and U15835 (N_15835,N_15422,N_15209);
and U15836 (N_15836,N_15279,N_15281);
xnor U15837 (N_15837,N_15200,N_15309);
xnor U15838 (N_15838,N_15574,N_15537);
nand U15839 (N_15839,N_15526,N_15530);
or U15840 (N_15840,N_15344,N_15296);
or U15841 (N_15841,N_15305,N_15546);
or U15842 (N_15842,N_15479,N_15588);
or U15843 (N_15843,N_15520,N_15448);
and U15844 (N_15844,N_15522,N_15412);
and U15845 (N_15845,N_15215,N_15488);
nor U15846 (N_15846,N_15467,N_15456);
nor U15847 (N_15847,N_15301,N_15587);
xor U15848 (N_15848,N_15387,N_15481);
xor U15849 (N_15849,N_15472,N_15500);
nor U15850 (N_15850,N_15504,N_15570);
or U15851 (N_15851,N_15480,N_15511);
xor U15852 (N_15852,N_15243,N_15250);
xnor U15853 (N_15853,N_15346,N_15384);
nand U15854 (N_15854,N_15362,N_15585);
nand U15855 (N_15855,N_15346,N_15590);
or U15856 (N_15856,N_15370,N_15375);
and U15857 (N_15857,N_15469,N_15308);
or U15858 (N_15858,N_15590,N_15584);
nand U15859 (N_15859,N_15208,N_15537);
nor U15860 (N_15860,N_15439,N_15440);
or U15861 (N_15861,N_15224,N_15487);
or U15862 (N_15862,N_15291,N_15333);
nand U15863 (N_15863,N_15383,N_15407);
xnor U15864 (N_15864,N_15230,N_15356);
and U15865 (N_15865,N_15400,N_15433);
xnor U15866 (N_15866,N_15544,N_15335);
xor U15867 (N_15867,N_15526,N_15488);
or U15868 (N_15868,N_15342,N_15466);
and U15869 (N_15869,N_15298,N_15371);
and U15870 (N_15870,N_15384,N_15229);
and U15871 (N_15871,N_15502,N_15456);
xor U15872 (N_15872,N_15425,N_15262);
or U15873 (N_15873,N_15431,N_15266);
and U15874 (N_15874,N_15243,N_15233);
and U15875 (N_15875,N_15402,N_15362);
and U15876 (N_15876,N_15217,N_15216);
or U15877 (N_15877,N_15402,N_15463);
nand U15878 (N_15878,N_15290,N_15541);
nor U15879 (N_15879,N_15305,N_15209);
nor U15880 (N_15880,N_15253,N_15380);
nand U15881 (N_15881,N_15314,N_15576);
nand U15882 (N_15882,N_15203,N_15462);
or U15883 (N_15883,N_15235,N_15554);
nand U15884 (N_15884,N_15398,N_15205);
xnor U15885 (N_15885,N_15493,N_15300);
xnor U15886 (N_15886,N_15226,N_15570);
nand U15887 (N_15887,N_15364,N_15547);
nor U15888 (N_15888,N_15486,N_15371);
nor U15889 (N_15889,N_15470,N_15315);
nand U15890 (N_15890,N_15343,N_15314);
and U15891 (N_15891,N_15502,N_15450);
nand U15892 (N_15892,N_15455,N_15357);
and U15893 (N_15893,N_15389,N_15505);
xor U15894 (N_15894,N_15449,N_15349);
xnor U15895 (N_15895,N_15501,N_15323);
nor U15896 (N_15896,N_15435,N_15297);
xor U15897 (N_15897,N_15446,N_15326);
or U15898 (N_15898,N_15482,N_15271);
xnor U15899 (N_15899,N_15285,N_15348);
xor U15900 (N_15900,N_15227,N_15383);
xnor U15901 (N_15901,N_15231,N_15562);
and U15902 (N_15902,N_15308,N_15325);
nor U15903 (N_15903,N_15269,N_15247);
nor U15904 (N_15904,N_15505,N_15477);
nand U15905 (N_15905,N_15273,N_15286);
or U15906 (N_15906,N_15247,N_15281);
nor U15907 (N_15907,N_15586,N_15241);
and U15908 (N_15908,N_15343,N_15576);
nand U15909 (N_15909,N_15499,N_15458);
or U15910 (N_15910,N_15266,N_15319);
and U15911 (N_15911,N_15518,N_15407);
or U15912 (N_15912,N_15595,N_15409);
and U15913 (N_15913,N_15558,N_15267);
and U15914 (N_15914,N_15528,N_15307);
nand U15915 (N_15915,N_15565,N_15424);
and U15916 (N_15916,N_15445,N_15589);
and U15917 (N_15917,N_15519,N_15202);
nand U15918 (N_15918,N_15412,N_15419);
and U15919 (N_15919,N_15233,N_15313);
and U15920 (N_15920,N_15528,N_15283);
nand U15921 (N_15921,N_15550,N_15575);
or U15922 (N_15922,N_15552,N_15375);
xnor U15923 (N_15923,N_15599,N_15336);
nand U15924 (N_15924,N_15570,N_15287);
xnor U15925 (N_15925,N_15483,N_15423);
nor U15926 (N_15926,N_15407,N_15470);
and U15927 (N_15927,N_15373,N_15204);
or U15928 (N_15928,N_15390,N_15470);
nor U15929 (N_15929,N_15345,N_15597);
and U15930 (N_15930,N_15302,N_15542);
nor U15931 (N_15931,N_15366,N_15336);
nand U15932 (N_15932,N_15466,N_15555);
or U15933 (N_15933,N_15443,N_15465);
nand U15934 (N_15934,N_15395,N_15288);
and U15935 (N_15935,N_15416,N_15285);
nor U15936 (N_15936,N_15417,N_15274);
xnor U15937 (N_15937,N_15219,N_15351);
nor U15938 (N_15938,N_15448,N_15289);
or U15939 (N_15939,N_15311,N_15491);
nor U15940 (N_15940,N_15343,N_15535);
nor U15941 (N_15941,N_15422,N_15223);
nand U15942 (N_15942,N_15588,N_15340);
xnor U15943 (N_15943,N_15410,N_15320);
nor U15944 (N_15944,N_15243,N_15229);
nand U15945 (N_15945,N_15405,N_15452);
and U15946 (N_15946,N_15520,N_15264);
xnor U15947 (N_15947,N_15392,N_15396);
nand U15948 (N_15948,N_15525,N_15263);
and U15949 (N_15949,N_15547,N_15398);
xor U15950 (N_15950,N_15210,N_15301);
nor U15951 (N_15951,N_15302,N_15359);
nor U15952 (N_15952,N_15242,N_15361);
nor U15953 (N_15953,N_15313,N_15557);
nor U15954 (N_15954,N_15549,N_15215);
or U15955 (N_15955,N_15253,N_15362);
and U15956 (N_15956,N_15525,N_15299);
nand U15957 (N_15957,N_15518,N_15458);
or U15958 (N_15958,N_15256,N_15480);
xor U15959 (N_15959,N_15340,N_15317);
nand U15960 (N_15960,N_15216,N_15400);
nand U15961 (N_15961,N_15235,N_15237);
and U15962 (N_15962,N_15323,N_15274);
or U15963 (N_15963,N_15460,N_15418);
nor U15964 (N_15964,N_15256,N_15567);
xor U15965 (N_15965,N_15442,N_15222);
nor U15966 (N_15966,N_15327,N_15535);
xnor U15967 (N_15967,N_15336,N_15433);
xnor U15968 (N_15968,N_15471,N_15369);
xor U15969 (N_15969,N_15247,N_15218);
nand U15970 (N_15970,N_15399,N_15593);
and U15971 (N_15971,N_15479,N_15412);
nand U15972 (N_15972,N_15532,N_15431);
or U15973 (N_15973,N_15535,N_15537);
nor U15974 (N_15974,N_15262,N_15395);
and U15975 (N_15975,N_15215,N_15536);
nand U15976 (N_15976,N_15254,N_15397);
and U15977 (N_15977,N_15505,N_15303);
xnor U15978 (N_15978,N_15403,N_15239);
nor U15979 (N_15979,N_15450,N_15211);
or U15980 (N_15980,N_15401,N_15407);
or U15981 (N_15981,N_15228,N_15332);
xor U15982 (N_15982,N_15541,N_15285);
or U15983 (N_15983,N_15427,N_15389);
xor U15984 (N_15984,N_15533,N_15213);
and U15985 (N_15985,N_15389,N_15494);
or U15986 (N_15986,N_15481,N_15326);
xor U15987 (N_15987,N_15502,N_15588);
nor U15988 (N_15988,N_15326,N_15529);
nand U15989 (N_15989,N_15257,N_15568);
and U15990 (N_15990,N_15310,N_15327);
and U15991 (N_15991,N_15585,N_15414);
nand U15992 (N_15992,N_15547,N_15584);
or U15993 (N_15993,N_15402,N_15385);
nand U15994 (N_15994,N_15293,N_15347);
and U15995 (N_15995,N_15318,N_15459);
or U15996 (N_15996,N_15355,N_15351);
or U15997 (N_15997,N_15239,N_15262);
or U15998 (N_15998,N_15457,N_15482);
xor U15999 (N_15999,N_15247,N_15554);
and U16000 (N_16000,N_15686,N_15935);
and U16001 (N_16001,N_15978,N_15796);
nand U16002 (N_16002,N_15690,N_15962);
xnor U16003 (N_16003,N_15741,N_15871);
nand U16004 (N_16004,N_15841,N_15735);
nand U16005 (N_16005,N_15863,N_15865);
xor U16006 (N_16006,N_15625,N_15763);
xnor U16007 (N_16007,N_15820,N_15626);
and U16008 (N_16008,N_15639,N_15613);
xnor U16009 (N_16009,N_15753,N_15859);
and U16010 (N_16010,N_15862,N_15842);
or U16011 (N_16011,N_15998,N_15986);
xor U16012 (N_16012,N_15891,N_15948);
and U16013 (N_16013,N_15929,N_15825);
xnor U16014 (N_16014,N_15600,N_15901);
and U16015 (N_16015,N_15621,N_15821);
and U16016 (N_16016,N_15839,N_15805);
and U16017 (N_16017,N_15630,N_15791);
xor U16018 (N_16018,N_15882,N_15816);
nor U16019 (N_16019,N_15977,N_15797);
and U16020 (N_16020,N_15781,N_15971);
nand U16021 (N_16021,N_15720,N_15730);
or U16022 (N_16022,N_15954,N_15666);
or U16023 (N_16023,N_15785,N_15910);
and U16024 (N_16024,N_15644,N_15773);
xnor U16025 (N_16025,N_15632,N_15677);
nor U16026 (N_16026,N_15965,N_15936);
xor U16027 (N_16027,N_15804,N_15780);
or U16028 (N_16028,N_15856,N_15744);
nor U16029 (N_16029,N_15667,N_15673);
and U16030 (N_16030,N_15790,N_15900);
xnor U16031 (N_16031,N_15895,N_15991);
xor U16032 (N_16032,N_15643,N_15757);
or U16033 (N_16033,N_15961,N_15736);
nor U16034 (N_16034,N_15828,N_15810);
and U16035 (N_16035,N_15803,N_15758);
nor U16036 (N_16036,N_15680,N_15890);
and U16037 (N_16037,N_15843,N_15619);
or U16038 (N_16038,N_15949,N_15792);
and U16039 (N_16039,N_15671,N_15762);
or U16040 (N_16040,N_15854,N_15649);
nand U16041 (N_16041,N_15684,N_15692);
nor U16042 (N_16042,N_15624,N_15605);
and U16043 (N_16043,N_15798,N_15727);
xnor U16044 (N_16044,N_15884,N_15618);
or U16045 (N_16045,N_15958,N_15653);
xnor U16046 (N_16046,N_15951,N_15628);
nor U16047 (N_16047,N_15722,N_15654);
and U16048 (N_16048,N_15990,N_15989);
or U16049 (N_16049,N_15725,N_15824);
xnor U16050 (N_16050,N_15728,N_15620);
and U16051 (N_16051,N_15745,N_15709);
or U16052 (N_16052,N_15918,N_15885);
and U16053 (N_16053,N_15999,N_15964);
xnor U16054 (N_16054,N_15658,N_15633);
xnor U16055 (N_16055,N_15738,N_15729);
nor U16056 (N_16056,N_15631,N_15661);
or U16057 (N_16057,N_15907,N_15768);
and U16058 (N_16058,N_15703,N_15855);
xor U16059 (N_16059,N_15813,N_15892);
and U16060 (N_16060,N_15778,N_15637);
or U16061 (N_16061,N_15887,N_15923);
nand U16062 (N_16062,N_15953,N_15646);
and U16063 (N_16063,N_15877,N_15934);
and U16064 (N_16064,N_15717,N_15611);
nand U16065 (N_16065,N_15732,N_15601);
or U16066 (N_16066,N_15919,N_15761);
nor U16067 (N_16067,N_15715,N_15849);
nand U16068 (N_16068,N_15636,N_15966);
nand U16069 (N_16069,N_15922,N_15615);
xnor U16070 (N_16070,N_15903,N_15694);
and U16071 (N_16071,N_15880,N_15604);
nor U16072 (N_16072,N_15784,N_15809);
nand U16073 (N_16073,N_15844,N_15648);
xnor U16074 (N_16074,N_15817,N_15875);
and U16075 (N_16075,N_15893,N_15852);
or U16076 (N_16076,N_15932,N_15651);
and U16077 (N_16077,N_15950,N_15876);
nor U16078 (N_16078,N_15984,N_15808);
or U16079 (N_16079,N_15988,N_15656);
nand U16080 (N_16080,N_15705,N_15731);
and U16081 (N_16081,N_15623,N_15603);
and U16082 (N_16082,N_15858,N_15898);
nor U16083 (N_16083,N_15664,N_15724);
or U16084 (N_16084,N_15838,N_15826);
or U16085 (N_16085,N_15723,N_15924);
xnor U16086 (N_16086,N_15967,N_15607);
and U16087 (N_16087,N_15827,N_15627);
or U16088 (N_16088,N_15739,N_15867);
xor U16089 (N_16089,N_15695,N_15756);
or U16090 (N_16090,N_15927,N_15851);
and U16091 (N_16091,N_15740,N_15629);
nor U16092 (N_16092,N_15814,N_15716);
nand U16093 (N_16093,N_15788,N_15748);
nor U16094 (N_16094,N_15972,N_15874);
nand U16095 (N_16095,N_15710,N_15952);
nand U16096 (N_16096,N_15946,N_15712);
or U16097 (N_16097,N_15767,N_15926);
and U16098 (N_16098,N_15771,N_15807);
xor U16099 (N_16099,N_15719,N_15879);
nand U16100 (N_16100,N_15789,N_15794);
and U16101 (N_16101,N_15714,N_15665);
or U16102 (N_16102,N_15845,N_15883);
xor U16103 (N_16103,N_15939,N_15755);
nor U16104 (N_16104,N_15764,N_15681);
and U16105 (N_16105,N_15645,N_15806);
or U16106 (N_16106,N_15802,N_15945);
nor U16107 (N_16107,N_15672,N_15749);
and U16108 (N_16108,N_15995,N_15691);
nand U16109 (N_16109,N_15905,N_15947);
or U16110 (N_16110,N_15641,N_15864);
nor U16111 (N_16111,N_15674,N_15669);
nor U16112 (N_16112,N_15920,N_15668);
or U16113 (N_16113,N_15683,N_15969);
xnor U16114 (N_16114,N_15996,N_15693);
or U16115 (N_16115,N_15957,N_15676);
and U16116 (N_16116,N_15751,N_15869);
and U16117 (N_16117,N_15622,N_15894);
or U16118 (N_16118,N_15793,N_15857);
and U16119 (N_16119,N_15787,N_15868);
and U16120 (N_16120,N_15979,N_15706);
or U16121 (N_16121,N_15993,N_15795);
or U16122 (N_16122,N_15878,N_15608);
nand U16123 (N_16123,N_15747,N_15870);
xnor U16124 (N_16124,N_15610,N_15769);
and U16125 (N_16125,N_15897,N_15702);
xnor U16126 (N_16126,N_15886,N_15963);
and U16127 (N_16127,N_15783,N_15997);
or U16128 (N_16128,N_15612,N_15733);
or U16129 (N_16129,N_15909,N_15888);
nor U16130 (N_16130,N_15635,N_15678);
or U16131 (N_16131,N_15687,N_15616);
nand U16132 (N_16132,N_15765,N_15960);
or U16133 (N_16133,N_15675,N_15742);
xor U16134 (N_16134,N_15896,N_15976);
or U16135 (N_16135,N_15743,N_15911);
nor U16136 (N_16136,N_15970,N_15662);
nor U16137 (N_16137,N_15663,N_15737);
and U16138 (N_16138,N_15861,N_15655);
nor U16139 (N_16139,N_15746,N_15779);
xor U16140 (N_16140,N_15602,N_15718);
nand U16141 (N_16141,N_15983,N_15698);
nand U16142 (N_16142,N_15754,N_15913);
nor U16143 (N_16143,N_15707,N_15899);
nand U16144 (N_16144,N_15638,N_15904);
nor U16145 (N_16145,N_15642,N_15938);
and U16146 (N_16146,N_15679,N_15614);
xnor U16147 (N_16147,N_15850,N_15943);
nor U16148 (N_16148,N_15959,N_15822);
or U16149 (N_16149,N_15609,N_15834);
xnor U16150 (N_16150,N_15928,N_15657);
nand U16151 (N_16151,N_15818,N_15786);
nand U16152 (N_16152,N_15914,N_15606);
nand U16153 (N_16153,N_15915,N_15873);
and U16154 (N_16154,N_15650,N_15982);
nand U16155 (N_16155,N_15881,N_15846);
nor U16156 (N_16156,N_15955,N_15974);
nor U16157 (N_16157,N_15829,N_15975);
nand U16158 (N_16158,N_15697,N_15734);
nand U16159 (N_16159,N_15713,N_15912);
or U16160 (N_16160,N_15685,N_15752);
and U16161 (N_16161,N_15640,N_15835);
nor U16162 (N_16162,N_15908,N_15688);
or U16163 (N_16163,N_15872,N_15985);
or U16164 (N_16164,N_15917,N_15775);
xor U16165 (N_16165,N_15940,N_15925);
xor U16166 (N_16166,N_15921,N_15774);
and U16167 (N_16167,N_15837,N_15832);
xor U16168 (N_16168,N_15906,N_15902);
nand U16169 (N_16169,N_15956,N_15889);
nor U16170 (N_16170,N_15647,N_15812);
and U16171 (N_16171,N_15726,N_15696);
or U16172 (N_16172,N_15973,N_15660);
xnor U16173 (N_16173,N_15670,N_15782);
nor U16174 (N_16174,N_15689,N_15811);
nand U16175 (N_16175,N_15860,N_15701);
and U16176 (N_16176,N_15981,N_15777);
or U16177 (N_16177,N_15848,N_15931);
xnor U16178 (N_16178,N_15866,N_15659);
nand U16179 (N_16179,N_15711,N_15704);
xnor U16180 (N_16180,N_15823,N_15799);
xor U16181 (N_16181,N_15916,N_15833);
xor U16182 (N_16182,N_15776,N_15847);
nand U16183 (N_16183,N_15801,N_15819);
or U16184 (N_16184,N_15652,N_15853);
nor U16185 (N_16185,N_15708,N_15760);
nand U16186 (N_16186,N_15750,N_15930);
or U16187 (N_16187,N_15700,N_15759);
nand U16188 (N_16188,N_15933,N_15830);
nor U16189 (N_16189,N_15987,N_15994);
and U16190 (N_16190,N_15766,N_15815);
nand U16191 (N_16191,N_15937,N_15617);
and U16192 (N_16192,N_15699,N_15634);
or U16193 (N_16193,N_15941,N_15772);
xor U16194 (N_16194,N_15770,N_15682);
or U16195 (N_16195,N_15944,N_15942);
or U16196 (N_16196,N_15721,N_15968);
and U16197 (N_16197,N_15840,N_15836);
and U16198 (N_16198,N_15992,N_15980);
and U16199 (N_16199,N_15831,N_15800);
nor U16200 (N_16200,N_15883,N_15787);
nand U16201 (N_16201,N_15831,N_15656);
or U16202 (N_16202,N_15952,N_15867);
xor U16203 (N_16203,N_15808,N_15669);
and U16204 (N_16204,N_15681,N_15867);
nor U16205 (N_16205,N_15950,N_15938);
nor U16206 (N_16206,N_15678,N_15870);
xor U16207 (N_16207,N_15604,N_15701);
and U16208 (N_16208,N_15881,N_15781);
xnor U16209 (N_16209,N_15683,N_15764);
nand U16210 (N_16210,N_15612,N_15851);
nor U16211 (N_16211,N_15813,N_15609);
nand U16212 (N_16212,N_15915,N_15716);
and U16213 (N_16213,N_15707,N_15790);
nor U16214 (N_16214,N_15979,N_15827);
nor U16215 (N_16215,N_15634,N_15609);
and U16216 (N_16216,N_15971,N_15994);
xnor U16217 (N_16217,N_15954,N_15672);
or U16218 (N_16218,N_15792,N_15785);
nand U16219 (N_16219,N_15640,N_15745);
nand U16220 (N_16220,N_15859,N_15696);
nor U16221 (N_16221,N_15734,N_15649);
and U16222 (N_16222,N_15915,N_15674);
nand U16223 (N_16223,N_15823,N_15696);
nand U16224 (N_16224,N_15818,N_15607);
and U16225 (N_16225,N_15850,N_15955);
and U16226 (N_16226,N_15735,N_15881);
and U16227 (N_16227,N_15665,N_15618);
nand U16228 (N_16228,N_15943,N_15778);
nand U16229 (N_16229,N_15845,N_15946);
or U16230 (N_16230,N_15958,N_15933);
nor U16231 (N_16231,N_15720,N_15859);
nand U16232 (N_16232,N_15866,N_15997);
nor U16233 (N_16233,N_15912,N_15809);
nor U16234 (N_16234,N_15926,N_15774);
and U16235 (N_16235,N_15801,N_15926);
nor U16236 (N_16236,N_15712,N_15743);
and U16237 (N_16237,N_15956,N_15708);
nor U16238 (N_16238,N_15632,N_15854);
or U16239 (N_16239,N_15628,N_15881);
xor U16240 (N_16240,N_15653,N_15785);
or U16241 (N_16241,N_15686,N_15627);
xnor U16242 (N_16242,N_15754,N_15921);
and U16243 (N_16243,N_15842,N_15974);
or U16244 (N_16244,N_15846,N_15976);
or U16245 (N_16245,N_15758,N_15892);
and U16246 (N_16246,N_15784,N_15729);
nor U16247 (N_16247,N_15632,N_15709);
xnor U16248 (N_16248,N_15642,N_15703);
nand U16249 (N_16249,N_15959,N_15899);
or U16250 (N_16250,N_15860,N_15726);
or U16251 (N_16251,N_15756,N_15856);
nor U16252 (N_16252,N_15723,N_15950);
nand U16253 (N_16253,N_15833,N_15699);
nand U16254 (N_16254,N_15722,N_15936);
nor U16255 (N_16255,N_15745,N_15945);
nor U16256 (N_16256,N_15993,N_15956);
and U16257 (N_16257,N_15745,N_15868);
and U16258 (N_16258,N_15996,N_15757);
nor U16259 (N_16259,N_15872,N_15935);
and U16260 (N_16260,N_15684,N_15970);
xor U16261 (N_16261,N_15924,N_15677);
xor U16262 (N_16262,N_15767,N_15771);
and U16263 (N_16263,N_15696,N_15668);
xor U16264 (N_16264,N_15966,N_15845);
nor U16265 (N_16265,N_15818,N_15755);
xor U16266 (N_16266,N_15781,N_15726);
xnor U16267 (N_16267,N_15728,N_15862);
or U16268 (N_16268,N_15775,N_15910);
nor U16269 (N_16269,N_15745,N_15980);
and U16270 (N_16270,N_15906,N_15978);
and U16271 (N_16271,N_15667,N_15619);
nand U16272 (N_16272,N_15617,N_15775);
or U16273 (N_16273,N_15733,N_15677);
or U16274 (N_16274,N_15789,N_15747);
nand U16275 (N_16275,N_15786,N_15916);
or U16276 (N_16276,N_15858,N_15915);
xor U16277 (N_16277,N_15618,N_15894);
nand U16278 (N_16278,N_15637,N_15910);
xnor U16279 (N_16279,N_15678,N_15819);
xnor U16280 (N_16280,N_15791,N_15895);
and U16281 (N_16281,N_15733,N_15903);
or U16282 (N_16282,N_15840,N_15620);
and U16283 (N_16283,N_15695,N_15977);
nor U16284 (N_16284,N_15918,N_15774);
or U16285 (N_16285,N_15758,N_15651);
nor U16286 (N_16286,N_15904,N_15924);
xnor U16287 (N_16287,N_15901,N_15604);
and U16288 (N_16288,N_15925,N_15612);
or U16289 (N_16289,N_15997,N_15657);
or U16290 (N_16290,N_15680,N_15703);
nor U16291 (N_16291,N_15743,N_15901);
nand U16292 (N_16292,N_15849,N_15622);
and U16293 (N_16293,N_15654,N_15612);
xor U16294 (N_16294,N_15875,N_15745);
or U16295 (N_16295,N_15657,N_15903);
or U16296 (N_16296,N_15984,N_15649);
nor U16297 (N_16297,N_15807,N_15778);
and U16298 (N_16298,N_15953,N_15649);
or U16299 (N_16299,N_15882,N_15773);
or U16300 (N_16300,N_15993,N_15695);
and U16301 (N_16301,N_15764,N_15857);
nor U16302 (N_16302,N_15792,N_15608);
xor U16303 (N_16303,N_15742,N_15747);
nor U16304 (N_16304,N_15950,N_15978);
nand U16305 (N_16305,N_15942,N_15600);
nor U16306 (N_16306,N_15717,N_15872);
nor U16307 (N_16307,N_15763,N_15692);
and U16308 (N_16308,N_15828,N_15904);
and U16309 (N_16309,N_15949,N_15872);
or U16310 (N_16310,N_15866,N_15868);
xor U16311 (N_16311,N_15818,N_15884);
or U16312 (N_16312,N_15870,N_15632);
xnor U16313 (N_16313,N_15720,N_15985);
xnor U16314 (N_16314,N_15644,N_15830);
or U16315 (N_16315,N_15669,N_15752);
nor U16316 (N_16316,N_15802,N_15899);
xor U16317 (N_16317,N_15821,N_15625);
nand U16318 (N_16318,N_15983,N_15761);
nand U16319 (N_16319,N_15945,N_15873);
and U16320 (N_16320,N_15636,N_15948);
xor U16321 (N_16321,N_15720,N_15869);
or U16322 (N_16322,N_15610,N_15825);
nand U16323 (N_16323,N_15652,N_15674);
nand U16324 (N_16324,N_15914,N_15713);
nand U16325 (N_16325,N_15866,N_15817);
and U16326 (N_16326,N_15894,N_15791);
xnor U16327 (N_16327,N_15855,N_15820);
and U16328 (N_16328,N_15799,N_15705);
nand U16329 (N_16329,N_15639,N_15622);
nand U16330 (N_16330,N_15846,N_15649);
xnor U16331 (N_16331,N_15641,N_15786);
nor U16332 (N_16332,N_15905,N_15993);
and U16333 (N_16333,N_15812,N_15950);
or U16334 (N_16334,N_15860,N_15830);
or U16335 (N_16335,N_15855,N_15697);
nand U16336 (N_16336,N_15958,N_15797);
and U16337 (N_16337,N_15997,N_15789);
or U16338 (N_16338,N_15703,N_15691);
or U16339 (N_16339,N_15980,N_15996);
xnor U16340 (N_16340,N_15759,N_15829);
nor U16341 (N_16341,N_15767,N_15600);
nor U16342 (N_16342,N_15620,N_15989);
and U16343 (N_16343,N_15712,N_15821);
nor U16344 (N_16344,N_15938,N_15719);
xnor U16345 (N_16345,N_15935,N_15827);
nor U16346 (N_16346,N_15695,N_15765);
or U16347 (N_16347,N_15944,N_15865);
or U16348 (N_16348,N_15789,N_15996);
and U16349 (N_16349,N_15666,N_15625);
nor U16350 (N_16350,N_15771,N_15808);
nand U16351 (N_16351,N_15847,N_15798);
nand U16352 (N_16352,N_15823,N_15894);
or U16353 (N_16353,N_15833,N_15653);
nand U16354 (N_16354,N_15850,N_15716);
or U16355 (N_16355,N_15789,N_15847);
xor U16356 (N_16356,N_15635,N_15649);
nor U16357 (N_16357,N_15999,N_15699);
and U16358 (N_16358,N_15844,N_15766);
nand U16359 (N_16359,N_15637,N_15957);
nor U16360 (N_16360,N_15614,N_15784);
and U16361 (N_16361,N_15661,N_15784);
nor U16362 (N_16362,N_15860,N_15772);
nor U16363 (N_16363,N_15636,N_15689);
nor U16364 (N_16364,N_15781,N_15844);
and U16365 (N_16365,N_15830,N_15885);
nor U16366 (N_16366,N_15837,N_15640);
xnor U16367 (N_16367,N_15957,N_15722);
xnor U16368 (N_16368,N_15650,N_15793);
xnor U16369 (N_16369,N_15799,N_15913);
and U16370 (N_16370,N_15691,N_15732);
nand U16371 (N_16371,N_15670,N_15897);
nor U16372 (N_16372,N_15942,N_15856);
or U16373 (N_16373,N_15849,N_15677);
xnor U16374 (N_16374,N_15751,N_15691);
nand U16375 (N_16375,N_15897,N_15712);
or U16376 (N_16376,N_15787,N_15683);
xor U16377 (N_16377,N_15644,N_15929);
nor U16378 (N_16378,N_15721,N_15610);
xnor U16379 (N_16379,N_15601,N_15989);
xor U16380 (N_16380,N_15935,N_15647);
or U16381 (N_16381,N_15611,N_15849);
and U16382 (N_16382,N_15986,N_15613);
nor U16383 (N_16383,N_15853,N_15813);
nand U16384 (N_16384,N_15835,N_15657);
nor U16385 (N_16385,N_15886,N_15930);
or U16386 (N_16386,N_15913,N_15723);
nor U16387 (N_16387,N_15608,N_15746);
or U16388 (N_16388,N_15700,N_15979);
or U16389 (N_16389,N_15759,N_15745);
and U16390 (N_16390,N_15750,N_15848);
and U16391 (N_16391,N_15647,N_15803);
nor U16392 (N_16392,N_15729,N_15908);
or U16393 (N_16393,N_15775,N_15714);
or U16394 (N_16394,N_15949,N_15901);
nor U16395 (N_16395,N_15864,N_15662);
xor U16396 (N_16396,N_15669,N_15892);
or U16397 (N_16397,N_15622,N_15655);
xor U16398 (N_16398,N_15649,N_15657);
and U16399 (N_16399,N_15822,N_15987);
and U16400 (N_16400,N_16122,N_16385);
nand U16401 (N_16401,N_16372,N_16176);
xnor U16402 (N_16402,N_16104,N_16160);
xnor U16403 (N_16403,N_16349,N_16155);
xor U16404 (N_16404,N_16261,N_16388);
xor U16405 (N_16405,N_16288,N_16259);
nor U16406 (N_16406,N_16082,N_16298);
and U16407 (N_16407,N_16101,N_16100);
nand U16408 (N_16408,N_16250,N_16293);
nor U16409 (N_16409,N_16084,N_16199);
nand U16410 (N_16410,N_16281,N_16369);
nor U16411 (N_16411,N_16395,N_16257);
xor U16412 (N_16412,N_16336,N_16269);
xor U16413 (N_16413,N_16152,N_16211);
xor U16414 (N_16414,N_16182,N_16297);
or U16415 (N_16415,N_16347,N_16060);
nor U16416 (N_16416,N_16076,N_16093);
nor U16417 (N_16417,N_16071,N_16179);
xor U16418 (N_16418,N_16364,N_16322);
xnor U16419 (N_16419,N_16241,N_16119);
or U16420 (N_16420,N_16196,N_16080);
xor U16421 (N_16421,N_16230,N_16058);
nor U16422 (N_16422,N_16099,N_16073);
nor U16423 (N_16423,N_16235,N_16392);
nor U16424 (N_16424,N_16150,N_16205);
or U16425 (N_16425,N_16217,N_16329);
xor U16426 (N_16426,N_16110,N_16353);
nand U16427 (N_16427,N_16394,N_16198);
nor U16428 (N_16428,N_16344,N_16022);
xor U16429 (N_16429,N_16292,N_16171);
or U16430 (N_16430,N_16024,N_16303);
nand U16431 (N_16431,N_16363,N_16126);
nor U16432 (N_16432,N_16277,N_16044);
nand U16433 (N_16433,N_16075,N_16214);
nand U16434 (N_16434,N_16328,N_16033);
nand U16435 (N_16435,N_16308,N_16262);
nor U16436 (N_16436,N_16190,N_16346);
nor U16437 (N_16437,N_16275,N_16129);
xnor U16438 (N_16438,N_16301,N_16354);
xnor U16439 (N_16439,N_16026,N_16059);
nand U16440 (N_16440,N_16371,N_16365);
nand U16441 (N_16441,N_16046,N_16186);
nor U16442 (N_16442,N_16227,N_16234);
and U16443 (N_16443,N_16002,N_16373);
nor U16444 (N_16444,N_16207,N_16156);
nand U16445 (N_16445,N_16131,N_16249);
or U16446 (N_16446,N_16089,N_16051);
nor U16447 (N_16447,N_16307,N_16218);
and U16448 (N_16448,N_16064,N_16181);
nand U16449 (N_16449,N_16192,N_16177);
or U16450 (N_16450,N_16352,N_16113);
or U16451 (N_16451,N_16115,N_16345);
nand U16452 (N_16452,N_16027,N_16017);
or U16453 (N_16453,N_16057,N_16013);
xor U16454 (N_16454,N_16007,N_16351);
xnor U16455 (N_16455,N_16374,N_16341);
nand U16456 (N_16456,N_16379,N_16109);
nand U16457 (N_16457,N_16128,N_16286);
and U16458 (N_16458,N_16135,N_16355);
and U16459 (N_16459,N_16054,N_16123);
nand U16460 (N_16460,N_16278,N_16220);
and U16461 (N_16461,N_16244,N_16103);
xnor U16462 (N_16462,N_16092,N_16312);
and U16463 (N_16463,N_16049,N_16197);
nand U16464 (N_16464,N_16117,N_16368);
or U16465 (N_16465,N_16136,N_16048);
nand U16466 (N_16466,N_16006,N_16132);
nand U16467 (N_16467,N_16139,N_16021);
xnor U16468 (N_16468,N_16065,N_16304);
or U16469 (N_16469,N_16321,N_16212);
nor U16470 (N_16470,N_16254,N_16223);
nand U16471 (N_16471,N_16360,N_16085);
and U16472 (N_16472,N_16225,N_16342);
and U16473 (N_16473,N_16087,N_16023);
xnor U16474 (N_16474,N_16072,N_16018);
nor U16475 (N_16475,N_16189,N_16224);
nand U16476 (N_16476,N_16034,N_16050);
nand U16477 (N_16477,N_16055,N_16173);
xor U16478 (N_16478,N_16037,N_16273);
and U16479 (N_16479,N_16012,N_16290);
nor U16480 (N_16480,N_16299,N_16195);
or U16481 (N_16481,N_16140,N_16141);
nand U16482 (N_16482,N_16145,N_16382);
xor U16483 (N_16483,N_16039,N_16170);
xor U16484 (N_16484,N_16338,N_16291);
xnor U16485 (N_16485,N_16094,N_16398);
nand U16486 (N_16486,N_16314,N_16053);
and U16487 (N_16487,N_16216,N_16316);
xnor U16488 (N_16488,N_16201,N_16063);
or U16489 (N_16489,N_16161,N_16175);
nand U16490 (N_16490,N_16003,N_16108);
nor U16491 (N_16491,N_16062,N_16289);
nand U16492 (N_16492,N_16266,N_16069);
nand U16493 (N_16493,N_16095,N_16020);
xnor U16494 (N_16494,N_16118,N_16383);
nor U16495 (N_16495,N_16004,N_16105);
and U16496 (N_16496,N_16294,N_16317);
xor U16497 (N_16497,N_16284,N_16031);
nor U16498 (N_16498,N_16200,N_16238);
and U16499 (N_16499,N_16239,N_16378);
xor U16500 (N_16500,N_16172,N_16384);
or U16501 (N_16501,N_16125,N_16138);
nand U16502 (N_16502,N_16265,N_16283);
xor U16503 (N_16503,N_16120,N_16300);
nor U16504 (N_16504,N_16019,N_16148);
xor U16505 (N_16505,N_16061,N_16319);
and U16506 (N_16506,N_16240,N_16334);
and U16507 (N_16507,N_16133,N_16246);
and U16508 (N_16508,N_16337,N_16107);
xor U16509 (N_16509,N_16130,N_16245);
and U16510 (N_16510,N_16014,N_16335);
nor U16511 (N_16511,N_16232,N_16208);
nor U16512 (N_16512,N_16295,N_16361);
nor U16513 (N_16513,N_16399,N_16008);
nand U16514 (N_16514,N_16121,N_16167);
and U16515 (N_16515,N_16011,N_16077);
and U16516 (N_16516,N_16040,N_16114);
and U16517 (N_16517,N_16358,N_16070);
or U16518 (N_16518,N_16124,N_16215);
and U16519 (N_16519,N_16134,N_16271);
nand U16520 (N_16520,N_16330,N_16256);
xor U16521 (N_16521,N_16315,N_16111);
nor U16522 (N_16522,N_16362,N_16083);
xnor U16523 (N_16523,N_16380,N_16390);
and U16524 (N_16524,N_16168,N_16228);
nor U16525 (N_16525,N_16397,N_16237);
nand U16526 (N_16526,N_16000,N_16035);
nor U16527 (N_16527,N_16268,N_16305);
xnor U16528 (N_16528,N_16203,N_16209);
and U16529 (N_16529,N_16356,N_16030);
xor U16530 (N_16530,N_16009,N_16274);
nand U16531 (N_16531,N_16016,N_16042);
nor U16532 (N_16532,N_16206,N_16178);
xnor U16533 (N_16533,N_16047,N_16086);
or U16534 (N_16534,N_16159,N_16067);
xnor U16535 (N_16535,N_16193,N_16323);
nand U16536 (N_16536,N_16376,N_16366);
xor U16537 (N_16537,N_16010,N_16096);
xnor U16538 (N_16538,N_16068,N_16210);
xor U16539 (N_16539,N_16306,N_16090);
and U16540 (N_16540,N_16045,N_16313);
or U16541 (N_16541,N_16276,N_16147);
xor U16542 (N_16542,N_16270,N_16252);
nand U16543 (N_16543,N_16157,N_16264);
and U16544 (N_16544,N_16028,N_16296);
nor U16545 (N_16545,N_16332,N_16112);
nor U16546 (N_16546,N_16106,N_16339);
nor U16547 (N_16547,N_16253,N_16185);
xor U16548 (N_16548,N_16285,N_16143);
xor U16549 (N_16549,N_16375,N_16343);
and U16550 (N_16550,N_16098,N_16183);
and U16551 (N_16551,N_16248,N_16279);
nor U16552 (N_16552,N_16043,N_16079);
nand U16553 (N_16553,N_16247,N_16309);
nor U16554 (N_16554,N_16005,N_16226);
and U16555 (N_16555,N_16377,N_16184);
nand U16556 (N_16556,N_16191,N_16162);
or U16557 (N_16557,N_16154,N_16153);
nand U16558 (N_16558,N_16097,N_16164);
xnor U16559 (N_16559,N_16081,N_16163);
xor U16560 (N_16560,N_16127,N_16015);
nand U16561 (N_16561,N_16263,N_16091);
nand U16562 (N_16562,N_16116,N_16267);
or U16563 (N_16563,N_16251,N_16327);
xor U16564 (N_16564,N_16204,N_16165);
or U16565 (N_16565,N_16038,N_16169);
and U16566 (N_16566,N_16386,N_16282);
nor U16567 (N_16567,N_16174,N_16137);
nand U16568 (N_16568,N_16310,N_16396);
nor U16569 (N_16569,N_16348,N_16236);
xnor U16570 (N_16570,N_16025,N_16233);
xor U16571 (N_16571,N_16333,N_16001);
nor U16572 (N_16572,N_16142,N_16287);
and U16573 (N_16573,N_16272,N_16188);
or U16574 (N_16574,N_16229,N_16221);
nor U16575 (N_16575,N_16357,N_16324);
and U16576 (N_16576,N_16146,N_16029);
xor U16577 (N_16577,N_16381,N_16367);
and U16578 (N_16578,N_16340,N_16387);
and U16579 (N_16579,N_16222,N_16180);
or U16580 (N_16580,N_16393,N_16158);
or U16581 (N_16581,N_16052,N_16331);
nand U16582 (N_16582,N_16302,N_16149);
nand U16583 (N_16583,N_16391,N_16151);
and U16584 (N_16584,N_16325,N_16213);
xnor U16585 (N_16585,N_16258,N_16255);
xnor U16586 (N_16586,N_16144,N_16187);
and U16587 (N_16587,N_16102,N_16088);
and U16588 (N_16588,N_16280,N_16326);
nor U16589 (N_16589,N_16350,N_16318);
nor U16590 (N_16590,N_16074,N_16231);
or U16591 (N_16591,N_16202,N_16359);
and U16592 (N_16592,N_16242,N_16166);
nand U16593 (N_16593,N_16078,N_16032);
and U16594 (N_16594,N_16194,N_16243);
and U16595 (N_16595,N_16260,N_16066);
or U16596 (N_16596,N_16041,N_16389);
xnor U16597 (N_16597,N_16320,N_16370);
nor U16598 (N_16598,N_16056,N_16219);
nor U16599 (N_16599,N_16311,N_16036);
or U16600 (N_16600,N_16265,N_16228);
nand U16601 (N_16601,N_16391,N_16289);
xor U16602 (N_16602,N_16288,N_16110);
or U16603 (N_16603,N_16120,N_16375);
or U16604 (N_16604,N_16123,N_16300);
nor U16605 (N_16605,N_16313,N_16003);
xnor U16606 (N_16606,N_16377,N_16229);
xnor U16607 (N_16607,N_16037,N_16104);
xor U16608 (N_16608,N_16257,N_16303);
or U16609 (N_16609,N_16108,N_16046);
or U16610 (N_16610,N_16377,N_16324);
nor U16611 (N_16611,N_16021,N_16063);
and U16612 (N_16612,N_16220,N_16310);
or U16613 (N_16613,N_16359,N_16085);
xor U16614 (N_16614,N_16163,N_16037);
nand U16615 (N_16615,N_16214,N_16158);
or U16616 (N_16616,N_16161,N_16369);
or U16617 (N_16617,N_16135,N_16191);
nand U16618 (N_16618,N_16167,N_16324);
nor U16619 (N_16619,N_16115,N_16332);
nor U16620 (N_16620,N_16328,N_16271);
and U16621 (N_16621,N_16155,N_16080);
or U16622 (N_16622,N_16161,N_16262);
nand U16623 (N_16623,N_16189,N_16241);
and U16624 (N_16624,N_16249,N_16272);
xor U16625 (N_16625,N_16047,N_16065);
or U16626 (N_16626,N_16111,N_16329);
and U16627 (N_16627,N_16170,N_16098);
xnor U16628 (N_16628,N_16276,N_16292);
nand U16629 (N_16629,N_16240,N_16280);
nor U16630 (N_16630,N_16388,N_16180);
and U16631 (N_16631,N_16107,N_16209);
nand U16632 (N_16632,N_16216,N_16359);
and U16633 (N_16633,N_16349,N_16129);
nand U16634 (N_16634,N_16263,N_16259);
xnor U16635 (N_16635,N_16238,N_16090);
and U16636 (N_16636,N_16015,N_16183);
nand U16637 (N_16637,N_16309,N_16053);
and U16638 (N_16638,N_16196,N_16030);
nor U16639 (N_16639,N_16237,N_16197);
nand U16640 (N_16640,N_16363,N_16004);
or U16641 (N_16641,N_16352,N_16102);
and U16642 (N_16642,N_16197,N_16010);
xor U16643 (N_16643,N_16290,N_16058);
or U16644 (N_16644,N_16357,N_16046);
xor U16645 (N_16645,N_16080,N_16131);
nor U16646 (N_16646,N_16375,N_16234);
and U16647 (N_16647,N_16153,N_16225);
nor U16648 (N_16648,N_16052,N_16245);
nor U16649 (N_16649,N_16069,N_16178);
nor U16650 (N_16650,N_16074,N_16353);
nand U16651 (N_16651,N_16237,N_16060);
and U16652 (N_16652,N_16169,N_16099);
xnor U16653 (N_16653,N_16072,N_16096);
or U16654 (N_16654,N_16374,N_16053);
nand U16655 (N_16655,N_16155,N_16104);
and U16656 (N_16656,N_16006,N_16192);
nor U16657 (N_16657,N_16223,N_16329);
xor U16658 (N_16658,N_16123,N_16261);
nand U16659 (N_16659,N_16029,N_16062);
nor U16660 (N_16660,N_16163,N_16217);
and U16661 (N_16661,N_16180,N_16154);
xnor U16662 (N_16662,N_16124,N_16048);
or U16663 (N_16663,N_16289,N_16236);
nand U16664 (N_16664,N_16149,N_16048);
nor U16665 (N_16665,N_16254,N_16048);
and U16666 (N_16666,N_16355,N_16253);
xnor U16667 (N_16667,N_16118,N_16056);
or U16668 (N_16668,N_16039,N_16100);
nand U16669 (N_16669,N_16226,N_16197);
nand U16670 (N_16670,N_16108,N_16287);
and U16671 (N_16671,N_16028,N_16140);
or U16672 (N_16672,N_16316,N_16135);
nand U16673 (N_16673,N_16365,N_16361);
and U16674 (N_16674,N_16264,N_16036);
xor U16675 (N_16675,N_16219,N_16147);
nand U16676 (N_16676,N_16032,N_16154);
xnor U16677 (N_16677,N_16372,N_16295);
nand U16678 (N_16678,N_16288,N_16050);
or U16679 (N_16679,N_16244,N_16251);
xor U16680 (N_16680,N_16058,N_16304);
or U16681 (N_16681,N_16150,N_16249);
and U16682 (N_16682,N_16343,N_16169);
xnor U16683 (N_16683,N_16332,N_16203);
nor U16684 (N_16684,N_16179,N_16365);
or U16685 (N_16685,N_16079,N_16152);
or U16686 (N_16686,N_16367,N_16357);
xnor U16687 (N_16687,N_16097,N_16203);
and U16688 (N_16688,N_16367,N_16310);
and U16689 (N_16689,N_16288,N_16150);
nand U16690 (N_16690,N_16231,N_16327);
xor U16691 (N_16691,N_16232,N_16198);
or U16692 (N_16692,N_16160,N_16172);
or U16693 (N_16693,N_16332,N_16072);
or U16694 (N_16694,N_16371,N_16293);
or U16695 (N_16695,N_16308,N_16013);
nand U16696 (N_16696,N_16058,N_16121);
xnor U16697 (N_16697,N_16351,N_16237);
xor U16698 (N_16698,N_16022,N_16139);
or U16699 (N_16699,N_16127,N_16219);
nor U16700 (N_16700,N_16099,N_16143);
nor U16701 (N_16701,N_16150,N_16344);
nand U16702 (N_16702,N_16372,N_16067);
nor U16703 (N_16703,N_16076,N_16216);
nor U16704 (N_16704,N_16387,N_16032);
and U16705 (N_16705,N_16396,N_16115);
xnor U16706 (N_16706,N_16144,N_16288);
or U16707 (N_16707,N_16223,N_16019);
and U16708 (N_16708,N_16083,N_16208);
or U16709 (N_16709,N_16132,N_16375);
or U16710 (N_16710,N_16390,N_16198);
nor U16711 (N_16711,N_16382,N_16077);
xor U16712 (N_16712,N_16067,N_16000);
or U16713 (N_16713,N_16170,N_16234);
or U16714 (N_16714,N_16199,N_16382);
xnor U16715 (N_16715,N_16271,N_16296);
nand U16716 (N_16716,N_16326,N_16256);
or U16717 (N_16717,N_16003,N_16147);
and U16718 (N_16718,N_16093,N_16216);
nand U16719 (N_16719,N_16080,N_16229);
xnor U16720 (N_16720,N_16205,N_16100);
xor U16721 (N_16721,N_16393,N_16117);
or U16722 (N_16722,N_16372,N_16336);
nor U16723 (N_16723,N_16217,N_16367);
nand U16724 (N_16724,N_16105,N_16034);
or U16725 (N_16725,N_16310,N_16292);
or U16726 (N_16726,N_16241,N_16307);
or U16727 (N_16727,N_16113,N_16134);
and U16728 (N_16728,N_16374,N_16001);
and U16729 (N_16729,N_16043,N_16228);
xnor U16730 (N_16730,N_16314,N_16080);
and U16731 (N_16731,N_16217,N_16112);
nand U16732 (N_16732,N_16016,N_16236);
xnor U16733 (N_16733,N_16211,N_16094);
xnor U16734 (N_16734,N_16105,N_16313);
and U16735 (N_16735,N_16335,N_16011);
nor U16736 (N_16736,N_16210,N_16360);
nor U16737 (N_16737,N_16029,N_16008);
nor U16738 (N_16738,N_16160,N_16054);
and U16739 (N_16739,N_16191,N_16157);
xor U16740 (N_16740,N_16155,N_16029);
or U16741 (N_16741,N_16087,N_16119);
or U16742 (N_16742,N_16063,N_16006);
or U16743 (N_16743,N_16392,N_16059);
or U16744 (N_16744,N_16298,N_16274);
nor U16745 (N_16745,N_16324,N_16037);
xor U16746 (N_16746,N_16073,N_16340);
or U16747 (N_16747,N_16214,N_16377);
xor U16748 (N_16748,N_16194,N_16199);
nor U16749 (N_16749,N_16145,N_16324);
nor U16750 (N_16750,N_16387,N_16085);
nor U16751 (N_16751,N_16371,N_16050);
nand U16752 (N_16752,N_16302,N_16116);
and U16753 (N_16753,N_16014,N_16137);
nand U16754 (N_16754,N_16247,N_16012);
or U16755 (N_16755,N_16165,N_16261);
or U16756 (N_16756,N_16019,N_16315);
and U16757 (N_16757,N_16201,N_16152);
and U16758 (N_16758,N_16330,N_16237);
and U16759 (N_16759,N_16356,N_16039);
and U16760 (N_16760,N_16249,N_16287);
or U16761 (N_16761,N_16006,N_16270);
or U16762 (N_16762,N_16287,N_16387);
nand U16763 (N_16763,N_16013,N_16060);
nor U16764 (N_16764,N_16176,N_16129);
or U16765 (N_16765,N_16270,N_16093);
nor U16766 (N_16766,N_16117,N_16057);
xor U16767 (N_16767,N_16312,N_16155);
xor U16768 (N_16768,N_16095,N_16326);
or U16769 (N_16769,N_16337,N_16044);
nor U16770 (N_16770,N_16115,N_16147);
nand U16771 (N_16771,N_16326,N_16010);
and U16772 (N_16772,N_16067,N_16390);
nand U16773 (N_16773,N_16210,N_16344);
xnor U16774 (N_16774,N_16351,N_16348);
or U16775 (N_16775,N_16387,N_16197);
nand U16776 (N_16776,N_16191,N_16111);
and U16777 (N_16777,N_16385,N_16157);
xnor U16778 (N_16778,N_16372,N_16015);
or U16779 (N_16779,N_16236,N_16156);
nand U16780 (N_16780,N_16385,N_16084);
nor U16781 (N_16781,N_16234,N_16220);
nor U16782 (N_16782,N_16108,N_16357);
and U16783 (N_16783,N_16245,N_16063);
or U16784 (N_16784,N_16145,N_16375);
nor U16785 (N_16785,N_16231,N_16300);
nor U16786 (N_16786,N_16132,N_16079);
xor U16787 (N_16787,N_16056,N_16209);
and U16788 (N_16788,N_16326,N_16276);
nor U16789 (N_16789,N_16023,N_16131);
or U16790 (N_16790,N_16376,N_16369);
xnor U16791 (N_16791,N_16388,N_16326);
xnor U16792 (N_16792,N_16058,N_16278);
nor U16793 (N_16793,N_16309,N_16112);
nand U16794 (N_16794,N_16063,N_16367);
nor U16795 (N_16795,N_16327,N_16068);
nor U16796 (N_16796,N_16108,N_16235);
xnor U16797 (N_16797,N_16357,N_16320);
nor U16798 (N_16798,N_16222,N_16162);
and U16799 (N_16799,N_16383,N_16130);
and U16800 (N_16800,N_16537,N_16746);
or U16801 (N_16801,N_16753,N_16479);
and U16802 (N_16802,N_16795,N_16695);
and U16803 (N_16803,N_16546,N_16644);
nor U16804 (N_16804,N_16666,N_16413);
nand U16805 (N_16805,N_16430,N_16400);
nor U16806 (N_16806,N_16453,N_16415);
or U16807 (N_16807,N_16733,N_16514);
xnor U16808 (N_16808,N_16759,N_16602);
and U16809 (N_16809,N_16445,N_16704);
nand U16810 (N_16810,N_16771,N_16507);
xor U16811 (N_16811,N_16788,N_16411);
and U16812 (N_16812,N_16767,N_16585);
nand U16813 (N_16813,N_16719,N_16655);
or U16814 (N_16814,N_16543,N_16576);
and U16815 (N_16815,N_16758,N_16451);
nor U16816 (N_16816,N_16611,N_16671);
nand U16817 (N_16817,N_16572,N_16559);
xnor U16818 (N_16818,N_16412,N_16799);
nor U16819 (N_16819,N_16423,N_16684);
xor U16820 (N_16820,N_16665,N_16631);
nand U16821 (N_16821,N_16701,N_16482);
nand U16822 (N_16822,N_16568,N_16716);
xnor U16823 (N_16823,N_16635,N_16551);
nand U16824 (N_16824,N_16553,N_16764);
and U16825 (N_16825,N_16567,N_16760);
xor U16826 (N_16826,N_16628,N_16427);
and U16827 (N_16827,N_16779,N_16691);
or U16828 (N_16828,N_16747,N_16683);
and U16829 (N_16829,N_16649,N_16639);
and U16830 (N_16830,N_16528,N_16680);
nand U16831 (N_16831,N_16774,N_16645);
and U16832 (N_16832,N_16539,N_16535);
or U16833 (N_16833,N_16452,N_16439);
xnor U16834 (N_16834,N_16506,N_16624);
nor U16835 (N_16835,N_16420,N_16679);
and U16836 (N_16836,N_16470,N_16501);
and U16837 (N_16837,N_16579,N_16401);
and U16838 (N_16838,N_16480,N_16474);
nand U16839 (N_16839,N_16563,N_16652);
nor U16840 (N_16840,N_16418,N_16743);
or U16841 (N_16841,N_16510,N_16626);
nor U16842 (N_16842,N_16486,N_16610);
nor U16843 (N_16843,N_16433,N_16462);
nor U16844 (N_16844,N_16589,N_16519);
or U16845 (N_16845,N_16773,N_16678);
xor U16846 (N_16846,N_16436,N_16662);
and U16847 (N_16847,N_16447,N_16698);
nand U16848 (N_16848,N_16722,N_16750);
nand U16849 (N_16849,N_16632,N_16521);
or U16850 (N_16850,N_16627,N_16775);
or U16851 (N_16851,N_16677,N_16581);
and U16852 (N_16852,N_16518,N_16545);
xor U16853 (N_16853,N_16598,N_16748);
xor U16854 (N_16854,N_16660,N_16573);
nor U16855 (N_16855,N_16755,N_16424);
or U16856 (N_16856,N_16772,N_16739);
nand U16857 (N_16857,N_16769,N_16527);
xor U16858 (N_16858,N_16570,N_16763);
xor U16859 (N_16859,N_16477,N_16650);
and U16860 (N_16860,N_16464,N_16475);
nor U16861 (N_16861,N_16577,N_16657);
nand U16862 (N_16862,N_16720,N_16777);
or U16863 (N_16863,N_16596,N_16600);
nor U16864 (N_16864,N_16571,N_16615);
nand U16865 (N_16865,N_16529,N_16580);
xnor U16866 (N_16866,N_16731,N_16786);
xor U16867 (N_16867,N_16497,N_16738);
xor U16868 (N_16868,N_16565,N_16637);
or U16869 (N_16869,N_16469,N_16736);
or U16870 (N_16870,N_16547,N_16508);
nand U16871 (N_16871,N_16406,N_16478);
nand U16872 (N_16872,N_16421,N_16766);
or U16873 (N_16873,N_16422,N_16450);
nand U16874 (N_16874,N_16703,N_16648);
nor U16875 (N_16875,N_16595,N_16560);
nor U16876 (N_16876,N_16597,N_16569);
nor U16877 (N_16877,N_16734,N_16705);
nand U16878 (N_16878,N_16416,N_16548);
nor U16879 (N_16879,N_16562,N_16647);
or U16880 (N_16880,N_16534,N_16793);
and U16881 (N_16881,N_16740,N_16667);
nor U16882 (N_16882,N_16414,N_16552);
xor U16883 (N_16883,N_16606,N_16756);
and U16884 (N_16884,N_16431,N_16604);
xor U16885 (N_16885,N_16781,N_16538);
nor U16886 (N_16886,N_16457,N_16710);
xnor U16887 (N_16887,N_16685,N_16690);
xnor U16888 (N_16888,N_16732,N_16664);
xnor U16889 (N_16889,N_16642,N_16785);
and U16890 (N_16890,N_16605,N_16542);
nand U16891 (N_16891,N_16646,N_16702);
xor U16892 (N_16892,N_16481,N_16409);
xnor U16893 (N_16893,N_16621,N_16455);
and U16894 (N_16894,N_16712,N_16717);
xnor U16895 (N_16895,N_16620,N_16643);
nand U16896 (N_16896,N_16540,N_16438);
nand U16897 (N_16897,N_16656,N_16728);
nor U16898 (N_16898,N_16511,N_16446);
nor U16899 (N_16899,N_16520,N_16417);
xor U16900 (N_16900,N_16517,N_16556);
nor U16901 (N_16901,N_16609,N_16599);
nand U16902 (N_16902,N_16493,N_16512);
or U16903 (N_16903,N_16454,N_16500);
and U16904 (N_16904,N_16762,N_16778);
and U16905 (N_16905,N_16724,N_16432);
xor U16906 (N_16906,N_16694,N_16798);
and U16907 (N_16907,N_16407,N_16640);
nor U16908 (N_16908,N_16531,N_16776);
nand U16909 (N_16909,N_16495,N_16711);
nor U16910 (N_16910,N_16752,N_16783);
xor U16911 (N_16911,N_16526,N_16471);
or U16912 (N_16912,N_16630,N_16532);
nor U16913 (N_16913,N_16434,N_16574);
nand U16914 (N_16914,N_16718,N_16437);
xnor U16915 (N_16915,N_16443,N_16663);
or U16916 (N_16916,N_16488,N_16670);
and U16917 (N_16917,N_16735,N_16463);
or U16918 (N_16918,N_16681,N_16582);
nor U16919 (N_16919,N_16715,N_16668);
nand U16920 (N_16920,N_16714,N_16588);
xnor U16921 (N_16921,N_16700,N_16402);
and U16922 (N_16922,N_16410,N_16513);
nand U16923 (N_16923,N_16460,N_16721);
xnor U16924 (N_16924,N_16654,N_16504);
nand U16925 (N_16925,N_16485,N_16601);
xor U16926 (N_16926,N_16692,N_16561);
nand U16927 (N_16927,N_16794,N_16614);
nor U16928 (N_16928,N_16675,N_16689);
nor U16929 (N_16929,N_16616,N_16564);
nand U16930 (N_16930,N_16708,N_16498);
xnor U16931 (N_16931,N_16603,N_16744);
nor U16932 (N_16932,N_16575,N_16676);
nand U16933 (N_16933,N_16405,N_16566);
nor U16934 (N_16934,N_16499,N_16403);
or U16935 (N_16935,N_16555,N_16673);
xnor U16936 (N_16936,N_16687,N_16522);
or U16937 (N_16937,N_16483,N_16709);
or U16938 (N_16938,N_16688,N_16473);
and U16939 (N_16939,N_16707,N_16404);
and U16940 (N_16940,N_16458,N_16792);
or U16941 (N_16941,N_16608,N_16490);
nand U16942 (N_16942,N_16465,N_16780);
or U16943 (N_16943,N_16787,N_16797);
and U16944 (N_16944,N_16737,N_16726);
nor U16945 (N_16945,N_16554,N_16784);
xor U16946 (N_16946,N_16651,N_16586);
nand U16947 (N_16947,N_16658,N_16425);
nand U16948 (N_16948,N_16461,N_16686);
or U16949 (N_16949,N_16557,N_16674);
or U16950 (N_16950,N_16730,N_16622);
or U16951 (N_16951,N_16741,N_16693);
xor U16952 (N_16952,N_16516,N_16444);
nand U16953 (N_16953,N_16593,N_16619);
nor U16954 (N_16954,N_16491,N_16549);
xnor U16955 (N_16955,N_16448,N_16487);
and U16956 (N_16956,N_16754,N_16796);
and U16957 (N_16957,N_16791,N_16629);
and U16958 (N_16958,N_16727,N_16697);
nand U16959 (N_16959,N_16441,N_16476);
xor U16960 (N_16960,N_16428,N_16623);
and U16961 (N_16961,N_16468,N_16713);
or U16962 (N_16962,N_16489,N_16789);
xor U16963 (N_16963,N_16590,N_16583);
xnor U16964 (N_16964,N_16533,N_16699);
and U16965 (N_16965,N_16633,N_16536);
xor U16966 (N_16966,N_16587,N_16496);
nand U16967 (N_16967,N_16653,N_16509);
nor U16968 (N_16968,N_16426,N_16558);
or U16969 (N_16969,N_16749,N_16523);
nor U16970 (N_16970,N_16617,N_16530);
xor U16971 (N_16971,N_16768,N_16550);
xnor U16972 (N_16972,N_16466,N_16419);
or U16973 (N_16973,N_16636,N_16467);
or U16974 (N_16974,N_16456,N_16525);
or U16975 (N_16975,N_16641,N_16429);
nor U16976 (N_16976,N_16442,N_16696);
nor U16977 (N_16977,N_16782,N_16659);
or U16978 (N_16978,N_16459,N_16492);
nor U16979 (N_16979,N_16751,N_16682);
or U16980 (N_16980,N_16790,N_16612);
xor U16981 (N_16981,N_16484,N_16505);
nand U16982 (N_16982,N_16672,N_16723);
or U16983 (N_16983,N_16669,N_16625);
nor U16984 (N_16984,N_16578,N_16770);
or U16985 (N_16985,N_16761,N_16706);
or U16986 (N_16986,N_16745,N_16618);
or U16987 (N_16987,N_16449,N_16494);
and U16988 (N_16988,N_16638,N_16757);
or U16989 (N_16989,N_16592,N_16594);
nor U16990 (N_16990,N_16591,N_16502);
and U16991 (N_16991,N_16634,N_16613);
or U16992 (N_16992,N_16408,N_16607);
or U16993 (N_16993,N_16544,N_16541);
nor U16994 (N_16994,N_16661,N_16584);
xor U16995 (N_16995,N_16524,N_16440);
nand U16996 (N_16996,N_16725,N_16515);
and U16997 (N_16997,N_16765,N_16742);
nor U16998 (N_16998,N_16435,N_16729);
nor U16999 (N_16999,N_16503,N_16472);
nand U17000 (N_17000,N_16786,N_16751);
or U17001 (N_17001,N_16628,N_16428);
and U17002 (N_17002,N_16421,N_16463);
or U17003 (N_17003,N_16681,N_16531);
xor U17004 (N_17004,N_16445,N_16722);
nand U17005 (N_17005,N_16736,N_16446);
nand U17006 (N_17006,N_16669,N_16629);
nor U17007 (N_17007,N_16550,N_16679);
nor U17008 (N_17008,N_16515,N_16564);
and U17009 (N_17009,N_16423,N_16732);
xor U17010 (N_17010,N_16422,N_16554);
nand U17011 (N_17011,N_16575,N_16442);
nor U17012 (N_17012,N_16589,N_16402);
nand U17013 (N_17013,N_16718,N_16781);
nor U17014 (N_17014,N_16425,N_16645);
xor U17015 (N_17015,N_16415,N_16488);
and U17016 (N_17016,N_16533,N_16423);
xnor U17017 (N_17017,N_16687,N_16506);
or U17018 (N_17018,N_16660,N_16753);
xnor U17019 (N_17019,N_16639,N_16442);
or U17020 (N_17020,N_16578,N_16711);
nand U17021 (N_17021,N_16504,N_16480);
or U17022 (N_17022,N_16734,N_16516);
or U17023 (N_17023,N_16493,N_16766);
nor U17024 (N_17024,N_16606,N_16496);
and U17025 (N_17025,N_16402,N_16443);
xnor U17026 (N_17026,N_16692,N_16702);
and U17027 (N_17027,N_16577,N_16747);
nand U17028 (N_17028,N_16782,N_16589);
xnor U17029 (N_17029,N_16466,N_16529);
and U17030 (N_17030,N_16514,N_16748);
nor U17031 (N_17031,N_16665,N_16591);
nor U17032 (N_17032,N_16598,N_16650);
nor U17033 (N_17033,N_16765,N_16745);
and U17034 (N_17034,N_16405,N_16730);
nor U17035 (N_17035,N_16498,N_16762);
or U17036 (N_17036,N_16597,N_16591);
nand U17037 (N_17037,N_16699,N_16478);
nand U17038 (N_17038,N_16590,N_16439);
nand U17039 (N_17039,N_16448,N_16638);
nand U17040 (N_17040,N_16662,N_16566);
or U17041 (N_17041,N_16615,N_16686);
and U17042 (N_17042,N_16494,N_16568);
xnor U17043 (N_17043,N_16573,N_16494);
xor U17044 (N_17044,N_16439,N_16664);
nand U17045 (N_17045,N_16787,N_16589);
or U17046 (N_17046,N_16406,N_16546);
nor U17047 (N_17047,N_16677,N_16470);
and U17048 (N_17048,N_16665,N_16667);
nand U17049 (N_17049,N_16550,N_16710);
and U17050 (N_17050,N_16632,N_16610);
and U17051 (N_17051,N_16442,N_16709);
nor U17052 (N_17052,N_16763,N_16566);
xnor U17053 (N_17053,N_16449,N_16583);
nor U17054 (N_17054,N_16652,N_16757);
or U17055 (N_17055,N_16654,N_16591);
xor U17056 (N_17056,N_16783,N_16724);
nand U17057 (N_17057,N_16746,N_16737);
and U17058 (N_17058,N_16501,N_16421);
and U17059 (N_17059,N_16602,N_16406);
and U17060 (N_17060,N_16649,N_16782);
and U17061 (N_17061,N_16599,N_16501);
or U17062 (N_17062,N_16480,N_16566);
and U17063 (N_17063,N_16656,N_16415);
nor U17064 (N_17064,N_16423,N_16442);
nand U17065 (N_17065,N_16499,N_16688);
and U17066 (N_17066,N_16454,N_16696);
nor U17067 (N_17067,N_16509,N_16536);
nor U17068 (N_17068,N_16723,N_16634);
xor U17069 (N_17069,N_16470,N_16706);
nor U17070 (N_17070,N_16779,N_16595);
xor U17071 (N_17071,N_16697,N_16533);
or U17072 (N_17072,N_16411,N_16794);
xor U17073 (N_17073,N_16486,N_16489);
or U17074 (N_17074,N_16703,N_16749);
nor U17075 (N_17075,N_16774,N_16731);
nor U17076 (N_17076,N_16709,N_16460);
or U17077 (N_17077,N_16547,N_16661);
and U17078 (N_17078,N_16673,N_16726);
nor U17079 (N_17079,N_16437,N_16696);
and U17080 (N_17080,N_16504,N_16701);
xnor U17081 (N_17081,N_16717,N_16484);
or U17082 (N_17082,N_16694,N_16517);
nor U17083 (N_17083,N_16621,N_16734);
and U17084 (N_17084,N_16718,N_16711);
and U17085 (N_17085,N_16405,N_16458);
or U17086 (N_17086,N_16508,N_16781);
xnor U17087 (N_17087,N_16744,N_16679);
and U17088 (N_17088,N_16655,N_16581);
nand U17089 (N_17089,N_16732,N_16702);
and U17090 (N_17090,N_16569,N_16553);
nor U17091 (N_17091,N_16583,N_16606);
nand U17092 (N_17092,N_16507,N_16656);
and U17093 (N_17093,N_16546,N_16444);
nand U17094 (N_17094,N_16527,N_16446);
nor U17095 (N_17095,N_16685,N_16753);
or U17096 (N_17096,N_16657,N_16779);
nor U17097 (N_17097,N_16587,N_16757);
or U17098 (N_17098,N_16683,N_16404);
or U17099 (N_17099,N_16422,N_16743);
and U17100 (N_17100,N_16481,N_16694);
xor U17101 (N_17101,N_16407,N_16726);
and U17102 (N_17102,N_16675,N_16754);
and U17103 (N_17103,N_16556,N_16510);
or U17104 (N_17104,N_16484,N_16612);
and U17105 (N_17105,N_16784,N_16781);
and U17106 (N_17106,N_16716,N_16495);
or U17107 (N_17107,N_16519,N_16534);
xor U17108 (N_17108,N_16707,N_16623);
and U17109 (N_17109,N_16469,N_16639);
or U17110 (N_17110,N_16606,N_16539);
and U17111 (N_17111,N_16561,N_16771);
xor U17112 (N_17112,N_16407,N_16461);
and U17113 (N_17113,N_16546,N_16704);
nand U17114 (N_17114,N_16588,N_16716);
and U17115 (N_17115,N_16415,N_16464);
nor U17116 (N_17116,N_16451,N_16464);
nor U17117 (N_17117,N_16498,N_16590);
nor U17118 (N_17118,N_16701,N_16711);
nand U17119 (N_17119,N_16501,N_16647);
nand U17120 (N_17120,N_16687,N_16669);
nand U17121 (N_17121,N_16541,N_16421);
or U17122 (N_17122,N_16435,N_16657);
nand U17123 (N_17123,N_16512,N_16563);
xor U17124 (N_17124,N_16687,N_16580);
nand U17125 (N_17125,N_16500,N_16522);
xnor U17126 (N_17126,N_16538,N_16564);
nand U17127 (N_17127,N_16455,N_16596);
nand U17128 (N_17128,N_16564,N_16721);
nand U17129 (N_17129,N_16410,N_16482);
or U17130 (N_17130,N_16452,N_16556);
nor U17131 (N_17131,N_16412,N_16784);
and U17132 (N_17132,N_16410,N_16701);
xnor U17133 (N_17133,N_16756,N_16546);
or U17134 (N_17134,N_16428,N_16645);
nor U17135 (N_17135,N_16773,N_16649);
nand U17136 (N_17136,N_16715,N_16568);
and U17137 (N_17137,N_16711,N_16777);
xnor U17138 (N_17138,N_16615,N_16472);
nor U17139 (N_17139,N_16482,N_16666);
and U17140 (N_17140,N_16614,N_16474);
nand U17141 (N_17141,N_16647,N_16565);
xnor U17142 (N_17142,N_16495,N_16706);
nand U17143 (N_17143,N_16620,N_16555);
xor U17144 (N_17144,N_16782,N_16477);
and U17145 (N_17145,N_16701,N_16671);
xnor U17146 (N_17146,N_16615,N_16545);
or U17147 (N_17147,N_16635,N_16643);
and U17148 (N_17148,N_16726,N_16413);
nand U17149 (N_17149,N_16734,N_16692);
xnor U17150 (N_17150,N_16605,N_16615);
nor U17151 (N_17151,N_16400,N_16644);
and U17152 (N_17152,N_16486,N_16403);
nor U17153 (N_17153,N_16670,N_16797);
nor U17154 (N_17154,N_16645,N_16771);
nor U17155 (N_17155,N_16776,N_16705);
nor U17156 (N_17156,N_16540,N_16617);
xnor U17157 (N_17157,N_16529,N_16409);
xnor U17158 (N_17158,N_16492,N_16497);
nor U17159 (N_17159,N_16703,N_16562);
or U17160 (N_17160,N_16455,N_16556);
nand U17161 (N_17161,N_16415,N_16692);
xor U17162 (N_17162,N_16484,N_16525);
and U17163 (N_17163,N_16753,N_16794);
nand U17164 (N_17164,N_16446,N_16623);
or U17165 (N_17165,N_16510,N_16536);
xnor U17166 (N_17166,N_16441,N_16606);
nand U17167 (N_17167,N_16606,N_16595);
or U17168 (N_17168,N_16661,N_16694);
xor U17169 (N_17169,N_16420,N_16536);
or U17170 (N_17170,N_16497,N_16548);
nor U17171 (N_17171,N_16512,N_16500);
and U17172 (N_17172,N_16720,N_16611);
and U17173 (N_17173,N_16572,N_16787);
xnor U17174 (N_17174,N_16541,N_16689);
nor U17175 (N_17175,N_16715,N_16618);
nor U17176 (N_17176,N_16615,N_16449);
and U17177 (N_17177,N_16639,N_16603);
and U17178 (N_17178,N_16526,N_16474);
nor U17179 (N_17179,N_16435,N_16773);
nand U17180 (N_17180,N_16572,N_16521);
or U17181 (N_17181,N_16688,N_16748);
xnor U17182 (N_17182,N_16658,N_16523);
and U17183 (N_17183,N_16453,N_16707);
or U17184 (N_17184,N_16727,N_16546);
and U17185 (N_17185,N_16568,N_16617);
nand U17186 (N_17186,N_16700,N_16721);
or U17187 (N_17187,N_16550,N_16662);
nor U17188 (N_17188,N_16454,N_16515);
nand U17189 (N_17189,N_16427,N_16623);
nand U17190 (N_17190,N_16577,N_16575);
nor U17191 (N_17191,N_16685,N_16686);
nand U17192 (N_17192,N_16412,N_16713);
nor U17193 (N_17193,N_16728,N_16744);
or U17194 (N_17194,N_16488,N_16774);
and U17195 (N_17195,N_16544,N_16492);
xor U17196 (N_17196,N_16669,N_16607);
nand U17197 (N_17197,N_16648,N_16410);
nand U17198 (N_17198,N_16495,N_16453);
nor U17199 (N_17199,N_16725,N_16612);
nand U17200 (N_17200,N_17143,N_17186);
and U17201 (N_17201,N_16884,N_16978);
nand U17202 (N_17202,N_16959,N_17179);
and U17203 (N_17203,N_16829,N_17164);
nand U17204 (N_17204,N_17198,N_16801);
or U17205 (N_17205,N_17194,N_17131);
xnor U17206 (N_17206,N_17112,N_16872);
and U17207 (N_17207,N_16891,N_16973);
xnor U17208 (N_17208,N_16949,N_16927);
nor U17209 (N_17209,N_17170,N_17012);
xor U17210 (N_17210,N_17081,N_16860);
nor U17211 (N_17211,N_17140,N_17197);
xnor U17212 (N_17212,N_16934,N_16844);
nor U17213 (N_17213,N_17003,N_16868);
or U17214 (N_17214,N_16996,N_16956);
nand U17215 (N_17215,N_17133,N_16822);
or U17216 (N_17216,N_16988,N_17106);
nor U17217 (N_17217,N_17006,N_16987);
xor U17218 (N_17218,N_17145,N_17155);
and U17219 (N_17219,N_16813,N_16857);
or U17220 (N_17220,N_17093,N_17068);
or U17221 (N_17221,N_16904,N_16933);
nor U17222 (N_17222,N_16853,N_16804);
xnor U17223 (N_17223,N_16869,N_17138);
and U17224 (N_17224,N_16885,N_16808);
and U17225 (N_17225,N_16895,N_17168);
or U17226 (N_17226,N_16858,N_16907);
xor U17227 (N_17227,N_17027,N_17064);
or U17228 (N_17228,N_17049,N_17117);
nor U17229 (N_17229,N_17094,N_16991);
nor U17230 (N_17230,N_16981,N_17090);
xnor U17231 (N_17231,N_16964,N_17084);
nor U17232 (N_17232,N_16923,N_16871);
xnor U17233 (N_17233,N_17128,N_16943);
or U17234 (N_17234,N_16993,N_16986);
and U17235 (N_17235,N_16824,N_17142);
or U17236 (N_17236,N_16831,N_17000);
nand U17237 (N_17237,N_16818,N_17134);
and U17238 (N_17238,N_17120,N_16913);
xor U17239 (N_17239,N_17125,N_17004);
nor U17240 (N_17240,N_17111,N_16870);
nand U17241 (N_17241,N_16819,N_17022);
and U17242 (N_17242,N_16952,N_16836);
and U17243 (N_17243,N_16873,N_16947);
and U17244 (N_17244,N_17100,N_17102);
nand U17245 (N_17245,N_16977,N_17113);
nand U17246 (N_17246,N_16916,N_16917);
nand U17247 (N_17247,N_17173,N_16851);
nor U17248 (N_17248,N_16866,N_17048);
nand U17249 (N_17249,N_16906,N_17051);
xor U17250 (N_17250,N_17074,N_17028);
xnor U17251 (N_17251,N_17174,N_16982);
and U17252 (N_17252,N_17129,N_16969);
nand U17253 (N_17253,N_16816,N_17137);
nand U17254 (N_17254,N_16825,N_17038);
nand U17255 (N_17255,N_17045,N_17165);
nor U17256 (N_17256,N_16837,N_16841);
xnor U17257 (N_17257,N_17024,N_16856);
xnor U17258 (N_17258,N_16854,N_17160);
xor U17259 (N_17259,N_16892,N_16838);
nor U17260 (N_17260,N_16879,N_16821);
nor U17261 (N_17261,N_17036,N_16963);
and U17262 (N_17262,N_16897,N_17053);
and U17263 (N_17263,N_16814,N_16939);
or U17264 (N_17264,N_17020,N_17069);
or U17265 (N_17265,N_17077,N_16887);
and U17266 (N_17266,N_17033,N_17055);
and U17267 (N_17267,N_16859,N_17144);
nand U17268 (N_17268,N_17035,N_17196);
nor U17269 (N_17269,N_16955,N_17147);
nand U17270 (N_17270,N_16984,N_17044);
nand U17271 (N_17271,N_17096,N_16863);
nor U17272 (N_17272,N_16881,N_16846);
xnor U17273 (N_17273,N_16840,N_17052);
xnor U17274 (N_17274,N_16985,N_17110);
and U17275 (N_17275,N_16890,N_17118);
and U17276 (N_17276,N_17149,N_17091);
or U17277 (N_17277,N_17030,N_17159);
or U17278 (N_17278,N_16979,N_17010);
nand U17279 (N_17279,N_16889,N_16929);
and U17280 (N_17280,N_16826,N_16926);
xnor U17281 (N_17281,N_17157,N_17065);
and U17282 (N_17282,N_17127,N_16850);
or U17283 (N_17283,N_17150,N_16880);
xor U17284 (N_17284,N_16997,N_16867);
nor U17285 (N_17285,N_16918,N_16928);
xor U17286 (N_17286,N_17178,N_17086);
xnor U17287 (N_17287,N_17104,N_17115);
xor U17288 (N_17288,N_17095,N_16875);
xor U17289 (N_17289,N_16864,N_16876);
nand U17290 (N_17290,N_17187,N_16886);
and U17291 (N_17291,N_16849,N_17021);
or U17292 (N_17292,N_17087,N_16883);
nand U17293 (N_17293,N_17067,N_17080);
and U17294 (N_17294,N_17002,N_16852);
nand U17295 (N_17295,N_16905,N_16970);
and U17296 (N_17296,N_16811,N_16954);
or U17297 (N_17297,N_16820,N_17025);
xor U17298 (N_17298,N_16896,N_17169);
and U17299 (N_17299,N_16805,N_17119);
nor U17300 (N_17300,N_17183,N_16835);
and U17301 (N_17301,N_16877,N_16810);
and U17302 (N_17302,N_17058,N_17177);
or U17303 (N_17303,N_17109,N_17114);
and U17304 (N_17304,N_16930,N_17008);
nand U17305 (N_17305,N_17031,N_17124);
xor U17306 (N_17306,N_16874,N_17063);
nand U17307 (N_17307,N_17188,N_16899);
nand U17308 (N_17308,N_16953,N_16999);
xor U17309 (N_17309,N_16800,N_17151);
xor U17310 (N_17310,N_17088,N_17189);
and U17311 (N_17311,N_17017,N_16976);
nand U17312 (N_17312,N_16834,N_17066);
and U17313 (N_17313,N_16862,N_17013);
nor U17314 (N_17314,N_16839,N_16998);
nand U17315 (N_17315,N_16902,N_17139);
or U17316 (N_17316,N_16971,N_17018);
or U17317 (N_17317,N_16915,N_17032);
nand U17318 (N_17318,N_16878,N_16968);
or U17319 (N_17319,N_16922,N_17016);
or U17320 (N_17320,N_16847,N_16803);
or U17321 (N_17321,N_17007,N_17073);
or U17322 (N_17322,N_17141,N_17029);
nand U17323 (N_17323,N_16957,N_17123);
and U17324 (N_17324,N_17156,N_17101);
or U17325 (N_17325,N_17199,N_17135);
nor U17326 (N_17326,N_16966,N_17043);
and U17327 (N_17327,N_16914,N_16924);
nand U17328 (N_17328,N_17009,N_17092);
nand U17329 (N_17329,N_16848,N_16830);
xnor U17330 (N_17330,N_17057,N_16936);
xor U17331 (N_17331,N_16843,N_16946);
nor U17332 (N_17332,N_17005,N_17099);
or U17333 (N_17333,N_17107,N_16961);
or U17334 (N_17334,N_17136,N_16812);
nor U17335 (N_17335,N_17116,N_17050);
nor U17336 (N_17336,N_17089,N_16932);
or U17337 (N_17337,N_16833,N_17108);
and U17338 (N_17338,N_17076,N_17132);
xnor U17339 (N_17339,N_17001,N_16865);
nor U17340 (N_17340,N_16958,N_17122);
or U17341 (N_17341,N_16941,N_17042);
or U17342 (N_17342,N_17072,N_16975);
or U17343 (N_17343,N_17166,N_16909);
or U17344 (N_17344,N_17130,N_17182);
or U17345 (N_17345,N_17191,N_16898);
nor U17346 (N_17346,N_16828,N_17158);
xnor U17347 (N_17347,N_17047,N_17172);
and U17348 (N_17348,N_17171,N_17019);
nand U17349 (N_17349,N_17059,N_17079);
nor U17350 (N_17350,N_16940,N_16855);
or U17351 (N_17351,N_16925,N_17026);
nand U17352 (N_17352,N_17148,N_17071);
or U17353 (N_17353,N_16980,N_16832);
and U17354 (N_17354,N_17195,N_16861);
nand U17355 (N_17355,N_17054,N_16983);
xor U17356 (N_17356,N_17023,N_17083);
and U17357 (N_17357,N_16823,N_16806);
nor U17358 (N_17358,N_17181,N_16901);
or U17359 (N_17359,N_16893,N_17190);
nor U17360 (N_17360,N_17060,N_17046);
nor U17361 (N_17361,N_16882,N_17167);
xnor U17362 (N_17362,N_16911,N_16967);
or U17363 (N_17363,N_17037,N_16960);
nand U17364 (N_17364,N_16908,N_17075);
and U17365 (N_17365,N_16994,N_17180);
and U17366 (N_17366,N_17014,N_17161);
and U17367 (N_17367,N_17034,N_16809);
or U17368 (N_17368,N_17015,N_17175);
and U17369 (N_17369,N_17192,N_16948);
nor U17370 (N_17370,N_16888,N_16965);
xor U17371 (N_17371,N_16817,N_16807);
or U17372 (N_17372,N_17070,N_16992);
nor U17373 (N_17373,N_17078,N_16845);
nand U17374 (N_17374,N_16974,N_17011);
nor U17375 (N_17375,N_17185,N_17193);
and U17376 (N_17376,N_17056,N_17184);
or U17377 (N_17377,N_16972,N_16950);
nor U17378 (N_17378,N_17176,N_16931);
nand U17379 (N_17379,N_16912,N_16900);
and U17380 (N_17380,N_16802,N_16995);
nor U17381 (N_17381,N_17126,N_16919);
and U17382 (N_17382,N_16921,N_17162);
nor U17383 (N_17383,N_16944,N_16962);
nand U17384 (N_17384,N_17154,N_16920);
and U17385 (N_17385,N_17163,N_16842);
or U17386 (N_17386,N_16942,N_17146);
xor U17387 (N_17387,N_17061,N_17152);
or U17388 (N_17388,N_17085,N_16945);
or U17389 (N_17389,N_16990,N_16815);
nand U17390 (N_17390,N_16937,N_17121);
and U17391 (N_17391,N_16989,N_17098);
xnor U17392 (N_17392,N_16951,N_17097);
xnor U17393 (N_17393,N_17039,N_16910);
nand U17394 (N_17394,N_17082,N_17041);
nand U17395 (N_17395,N_17062,N_16827);
and U17396 (N_17396,N_17103,N_17105);
and U17397 (N_17397,N_17040,N_16894);
nor U17398 (N_17398,N_16903,N_16935);
or U17399 (N_17399,N_17153,N_16938);
nand U17400 (N_17400,N_16802,N_17191);
or U17401 (N_17401,N_17081,N_16910);
or U17402 (N_17402,N_17118,N_16981);
nand U17403 (N_17403,N_17052,N_17165);
xor U17404 (N_17404,N_16835,N_17116);
and U17405 (N_17405,N_16884,N_16973);
nand U17406 (N_17406,N_17026,N_17068);
xor U17407 (N_17407,N_16887,N_17138);
nor U17408 (N_17408,N_17044,N_17167);
xnor U17409 (N_17409,N_16805,N_16975);
xor U17410 (N_17410,N_16893,N_16902);
xnor U17411 (N_17411,N_17159,N_17095);
nand U17412 (N_17412,N_16914,N_16806);
nor U17413 (N_17413,N_17011,N_16973);
and U17414 (N_17414,N_17182,N_17149);
xnor U17415 (N_17415,N_16818,N_17030);
nor U17416 (N_17416,N_16884,N_17021);
and U17417 (N_17417,N_16848,N_17155);
nor U17418 (N_17418,N_17033,N_16904);
or U17419 (N_17419,N_16944,N_16905);
nor U17420 (N_17420,N_16852,N_17037);
nor U17421 (N_17421,N_17046,N_17199);
or U17422 (N_17422,N_17040,N_16803);
nand U17423 (N_17423,N_16917,N_16868);
and U17424 (N_17424,N_16828,N_16936);
nor U17425 (N_17425,N_16800,N_16942);
and U17426 (N_17426,N_16864,N_16870);
and U17427 (N_17427,N_17184,N_16952);
or U17428 (N_17428,N_16834,N_17051);
and U17429 (N_17429,N_17133,N_17039);
nand U17430 (N_17430,N_16971,N_17096);
or U17431 (N_17431,N_17152,N_17086);
and U17432 (N_17432,N_16901,N_16944);
and U17433 (N_17433,N_17150,N_17047);
nor U17434 (N_17434,N_17101,N_17185);
xnor U17435 (N_17435,N_17192,N_16887);
nand U17436 (N_17436,N_16839,N_16851);
or U17437 (N_17437,N_16904,N_16914);
or U17438 (N_17438,N_16888,N_17092);
or U17439 (N_17439,N_17092,N_17133);
xor U17440 (N_17440,N_16913,N_16835);
nand U17441 (N_17441,N_17009,N_16813);
or U17442 (N_17442,N_17078,N_17043);
nand U17443 (N_17443,N_17027,N_17035);
nand U17444 (N_17444,N_17101,N_16800);
nand U17445 (N_17445,N_16982,N_17063);
and U17446 (N_17446,N_17014,N_17020);
xor U17447 (N_17447,N_17070,N_16952);
nor U17448 (N_17448,N_17024,N_16824);
nand U17449 (N_17449,N_16950,N_17169);
xor U17450 (N_17450,N_17032,N_17165);
nor U17451 (N_17451,N_17158,N_17073);
nor U17452 (N_17452,N_17095,N_16999);
nor U17453 (N_17453,N_17183,N_16868);
nor U17454 (N_17454,N_16836,N_17064);
nor U17455 (N_17455,N_16908,N_17197);
xnor U17456 (N_17456,N_16849,N_17036);
xor U17457 (N_17457,N_16869,N_16934);
xor U17458 (N_17458,N_17058,N_16941);
and U17459 (N_17459,N_16807,N_17062);
xnor U17460 (N_17460,N_16932,N_17057);
nand U17461 (N_17461,N_16957,N_16854);
nand U17462 (N_17462,N_17133,N_17163);
xnor U17463 (N_17463,N_17129,N_17051);
nor U17464 (N_17464,N_16905,N_17135);
xnor U17465 (N_17465,N_16836,N_17170);
and U17466 (N_17466,N_17120,N_16894);
nor U17467 (N_17467,N_17152,N_17078);
nand U17468 (N_17468,N_17152,N_16879);
or U17469 (N_17469,N_17021,N_17161);
or U17470 (N_17470,N_16879,N_17058);
xor U17471 (N_17471,N_16961,N_16811);
and U17472 (N_17472,N_16923,N_17138);
or U17473 (N_17473,N_17092,N_16882);
xor U17474 (N_17474,N_16944,N_17122);
or U17475 (N_17475,N_17132,N_16911);
xor U17476 (N_17476,N_16905,N_17042);
nor U17477 (N_17477,N_17168,N_16938);
nor U17478 (N_17478,N_17025,N_17167);
nor U17479 (N_17479,N_17022,N_17125);
and U17480 (N_17480,N_17191,N_17112);
xnor U17481 (N_17481,N_17125,N_17147);
and U17482 (N_17482,N_17174,N_17141);
and U17483 (N_17483,N_16881,N_16843);
nand U17484 (N_17484,N_17020,N_16836);
nor U17485 (N_17485,N_16848,N_17057);
and U17486 (N_17486,N_17077,N_16929);
or U17487 (N_17487,N_16866,N_16867);
or U17488 (N_17488,N_16832,N_17053);
nand U17489 (N_17489,N_17008,N_16887);
nor U17490 (N_17490,N_17182,N_16800);
xnor U17491 (N_17491,N_16971,N_17152);
nand U17492 (N_17492,N_17020,N_17165);
nor U17493 (N_17493,N_16843,N_17139);
or U17494 (N_17494,N_16950,N_17095);
and U17495 (N_17495,N_17055,N_16958);
nand U17496 (N_17496,N_16993,N_17077);
and U17497 (N_17497,N_17172,N_17152);
xnor U17498 (N_17498,N_17090,N_16918);
or U17499 (N_17499,N_17153,N_16846);
nor U17500 (N_17500,N_17004,N_16800);
nor U17501 (N_17501,N_16892,N_16815);
nor U17502 (N_17502,N_16806,N_16812);
nand U17503 (N_17503,N_16919,N_16913);
nand U17504 (N_17504,N_16950,N_17029);
xnor U17505 (N_17505,N_16949,N_16911);
and U17506 (N_17506,N_17145,N_16863);
and U17507 (N_17507,N_17156,N_17095);
nor U17508 (N_17508,N_16924,N_16895);
or U17509 (N_17509,N_17071,N_17159);
and U17510 (N_17510,N_16822,N_16992);
or U17511 (N_17511,N_17179,N_17198);
nor U17512 (N_17512,N_17166,N_17037);
nor U17513 (N_17513,N_16981,N_17186);
or U17514 (N_17514,N_16971,N_16998);
and U17515 (N_17515,N_17050,N_17144);
or U17516 (N_17516,N_17008,N_17003);
nor U17517 (N_17517,N_16833,N_17102);
xor U17518 (N_17518,N_16894,N_16961);
and U17519 (N_17519,N_16976,N_16882);
nor U17520 (N_17520,N_17128,N_16988);
or U17521 (N_17521,N_16827,N_17153);
xor U17522 (N_17522,N_17077,N_17098);
or U17523 (N_17523,N_16872,N_16948);
nand U17524 (N_17524,N_16898,N_17002);
nor U17525 (N_17525,N_16836,N_16948);
nor U17526 (N_17526,N_16954,N_17198);
nor U17527 (N_17527,N_16972,N_16880);
xor U17528 (N_17528,N_17085,N_16827);
nand U17529 (N_17529,N_17032,N_16804);
xnor U17530 (N_17530,N_17191,N_16957);
xor U17531 (N_17531,N_16913,N_16944);
or U17532 (N_17532,N_17094,N_17039);
nand U17533 (N_17533,N_16917,N_17038);
and U17534 (N_17534,N_17044,N_17136);
and U17535 (N_17535,N_16906,N_16819);
xnor U17536 (N_17536,N_17082,N_16832);
xor U17537 (N_17537,N_17120,N_17017);
xnor U17538 (N_17538,N_16949,N_16832);
xor U17539 (N_17539,N_17140,N_16817);
nand U17540 (N_17540,N_16934,N_16992);
and U17541 (N_17541,N_17164,N_16934);
nand U17542 (N_17542,N_16923,N_17024);
xor U17543 (N_17543,N_16962,N_17081);
xnor U17544 (N_17544,N_17153,N_16984);
or U17545 (N_17545,N_17148,N_16981);
or U17546 (N_17546,N_16964,N_16958);
nor U17547 (N_17547,N_17005,N_17114);
nor U17548 (N_17548,N_16845,N_17080);
nor U17549 (N_17549,N_17001,N_17149);
nand U17550 (N_17550,N_17158,N_16959);
or U17551 (N_17551,N_16974,N_17103);
xor U17552 (N_17552,N_16982,N_16875);
and U17553 (N_17553,N_17059,N_17188);
and U17554 (N_17554,N_16902,N_17191);
nor U17555 (N_17555,N_17144,N_17065);
nand U17556 (N_17556,N_16961,N_16854);
or U17557 (N_17557,N_16827,N_17100);
nand U17558 (N_17558,N_17186,N_17121);
nand U17559 (N_17559,N_17176,N_16856);
nor U17560 (N_17560,N_16963,N_17051);
nand U17561 (N_17561,N_16899,N_17036);
and U17562 (N_17562,N_17137,N_16939);
xor U17563 (N_17563,N_16833,N_17079);
or U17564 (N_17564,N_17002,N_17133);
or U17565 (N_17565,N_17112,N_16948);
xor U17566 (N_17566,N_17178,N_16995);
or U17567 (N_17567,N_17159,N_16817);
nor U17568 (N_17568,N_16848,N_16829);
or U17569 (N_17569,N_17083,N_17073);
nand U17570 (N_17570,N_17070,N_16823);
and U17571 (N_17571,N_17183,N_16957);
and U17572 (N_17572,N_16958,N_16806);
or U17573 (N_17573,N_17086,N_16950);
nor U17574 (N_17574,N_16926,N_16981);
nor U17575 (N_17575,N_16912,N_16913);
nor U17576 (N_17576,N_16940,N_16884);
or U17577 (N_17577,N_16800,N_16856);
xnor U17578 (N_17578,N_17170,N_16977);
xor U17579 (N_17579,N_16992,N_16946);
xor U17580 (N_17580,N_16841,N_16976);
nand U17581 (N_17581,N_17065,N_17001);
nand U17582 (N_17582,N_17127,N_17109);
nor U17583 (N_17583,N_17137,N_17193);
and U17584 (N_17584,N_17137,N_16887);
xor U17585 (N_17585,N_17167,N_16876);
or U17586 (N_17586,N_17038,N_17139);
xor U17587 (N_17587,N_17018,N_16802);
xor U17588 (N_17588,N_16803,N_17004);
xor U17589 (N_17589,N_17094,N_16982);
and U17590 (N_17590,N_16878,N_17165);
nor U17591 (N_17591,N_16979,N_17179);
or U17592 (N_17592,N_17106,N_17166);
xor U17593 (N_17593,N_16950,N_16910);
nor U17594 (N_17594,N_17091,N_17080);
xnor U17595 (N_17595,N_17025,N_17123);
nor U17596 (N_17596,N_17068,N_16921);
nand U17597 (N_17597,N_17086,N_16999);
xnor U17598 (N_17598,N_17097,N_17092);
and U17599 (N_17599,N_17153,N_17130);
nand U17600 (N_17600,N_17296,N_17501);
or U17601 (N_17601,N_17349,N_17593);
nand U17602 (N_17602,N_17285,N_17270);
or U17603 (N_17603,N_17509,N_17469);
nand U17604 (N_17604,N_17395,N_17209);
and U17605 (N_17605,N_17314,N_17399);
and U17606 (N_17606,N_17241,N_17466);
nand U17607 (N_17607,N_17313,N_17563);
or U17608 (N_17608,N_17362,N_17441);
nand U17609 (N_17609,N_17481,N_17398);
and U17610 (N_17610,N_17424,N_17586);
or U17611 (N_17611,N_17384,N_17453);
or U17612 (N_17612,N_17365,N_17476);
nor U17613 (N_17613,N_17576,N_17345);
nor U17614 (N_17614,N_17344,N_17248);
or U17615 (N_17615,N_17472,N_17213);
nand U17616 (N_17616,N_17369,N_17530);
nand U17617 (N_17617,N_17340,N_17376);
nand U17618 (N_17618,N_17432,N_17403);
nand U17619 (N_17619,N_17330,N_17503);
xor U17620 (N_17620,N_17238,N_17565);
and U17621 (N_17621,N_17416,N_17323);
nor U17622 (N_17622,N_17276,N_17236);
xor U17623 (N_17623,N_17474,N_17315);
and U17624 (N_17624,N_17326,N_17450);
nor U17625 (N_17625,N_17597,N_17214);
and U17626 (N_17626,N_17247,N_17320);
or U17627 (N_17627,N_17380,N_17310);
nor U17628 (N_17628,N_17298,N_17587);
nand U17629 (N_17629,N_17373,N_17363);
or U17630 (N_17630,N_17533,N_17378);
or U17631 (N_17631,N_17538,N_17516);
nand U17632 (N_17632,N_17559,N_17510);
or U17633 (N_17633,N_17351,N_17311);
or U17634 (N_17634,N_17519,N_17488);
or U17635 (N_17635,N_17451,N_17435);
or U17636 (N_17636,N_17583,N_17278);
and U17637 (N_17637,N_17419,N_17318);
and U17638 (N_17638,N_17402,N_17212);
nor U17639 (N_17639,N_17383,N_17551);
nand U17640 (N_17640,N_17341,N_17361);
nand U17641 (N_17641,N_17396,N_17337);
and U17642 (N_17642,N_17571,N_17391);
xor U17643 (N_17643,N_17215,N_17288);
nor U17644 (N_17644,N_17425,N_17271);
nor U17645 (N_17645,N_17377,N_17492);
nor U17646 (N_17646,N_17580,N_17226);
or U17647 (N_17647,N_17590,N_17521);
and U17648 (N_17648,N_17442,N_17431);
nand U17649 (N_17649,N_17397,N_17475);
or U17650 (N_17650,N_17568,N_17303);
or U17651 (N_17651,N_17459,N_17542);
nor U17652 (N_17652,N_17536,N_17591);
xor U17653 (N_17653,N_17302,N_17307);
or U17654 (N_17654,N_17232,N_17294);
nand U17655 (N_17655,N_17467,N_17452);
nor U17656 (N_17656,N_17550,N_17389);
xor U17657 (N_17657,N_17347,N_17287);
xnor U17658 (N_17658,N_17529,N_17532);
xor U17659 (N_17659,N_17350,N_17444);
nor U17660 (N_17660,N_17228,N_17418);
xnor U17661 (N_17661,N_17234,N_17443);
or U17662 (N_17662,N_17406,N_17566);
or U17663 (N_17663,N_17211,N_17574);
nor U17664 (N_17664,N_17581,N_17219);
and U17665 (N_17665,N_17308,N_17266);
and U17666 (N_17666,N_17272,N_17242);
xor U17667 (N_17667,N_17306,N_17421);
or U17668 (N_17668,N_17371,N_17561);
and U17669 (N_17669,N_17374,N_17372);
or U17670 (N_17670,N_17407,N_17237);
and U17671 (N_17671,N_17460,N_17355);
nor U17672 (N_17672,N_17200,N_17412);
nand U17673 (N_17673,N_17417,N_17358);
nor U17674 (N_17674,N_17375,N_17235);
and U17675 (N_17675,N_17484,N_17495);
and U17676 (N_17676,N_17217,N_17202);
nand U17677 (N_17677,N_17524,N_17410);
and U17678 (N_17678,N_17553,N_17342);
and U17679 (N_17679,N_17497,N_17392);
nor U17680 (N_17680,N_17269,N_17301);
and U17681 (N_17681,N_17390,N_17394);
xor U17682 (N_17682,N_17292,N_17539);
nand U17683 (N_17683,N_17253,N_17393);
and U17684 (N_17684,N_17336,N_17534);
nor U17685 (N_17685,N_17557,N_17487);
xor U17686 (N_17686,N_17227,N_17367);
and U17687 (N_17687,N_17449,N_17579);
nand U17688 (N_17688,N_17496,N_17368);
xor U17689 (N_17689,N_17327,N_17427);
and U17690 (N_17690,N_17457,N_17258);
nor U17691 (N_17691,N_17468,N_17598);
nor U17692 (N_17692,N_17325,N_17423);
nor U17693 (N_17693,N_17456,N_17562);
nand U17694 (N_17694,N_17319,N_17331);
and U17695 (N_17695,N_17520,N_17295);
xnor U17696 (N_17696,N_17429,N_17360);
or U17697 (N_17697,N_17245,N_17354);
or U17698 (N_17698,N_17494,N_17352);
xnor U17699 (N_17699,N_17246,N_17477);
and U17700 (N_17700,N_17277,N_17401);
or U17701 (N_17701,N_17317,N_17531);
and U17702 (N_17702,N_17312,N_17366);
or U17703 (N_17703,N_17414,N_17556);
nor U17704 (N_17704,N_17259,N_17305);
nor U17705 (N_17705,N_17458,N_17430);
xnor U17706 (N_17706,N_17502,N_17233);
xnor U17707 (N_17707,N_17518,N_17517);
and U17708 (N_17708,N_17426,N_17386);
nand U17709 (N_17709,N_17405,N_17223);
and U17710 (N_17710,N_17282,N_17229);
xnor U17711 (N_17711,N_17499,N_17493);
and U17712 (N_17712,N_17263,N_17387);
or U17713 (N_17713,N_17445,N_17244);
nand U17714 (N_17714,N_17257,N_17498);
and U17715 (N_17715,N_17549,N_17504);
and U17716 (N_17716,N_17290,N_17478);
xnor U17717 (N_17717,N_17230,N_17274);
nand U17718 (N_17718,N_17348,N_17379);
and U17719 (N_17719,N_17275,N_17221);
and U17720 (N_17720,N_17512,N_17514);
nor U17721 (N_17721,N_17413,N_17588);
or U17722 (N_17722,N_17555,N_17224);
nor U17723 (N_17723,N_17334,N_17385);
xnor U17724 (N_17724,N_17578,N_17511);
nand U17725 (N_17725,N_17268,N_17322);
nand U17726 (N_17726,N_17438,N_17515);
xor U17727 (N_17727,N_17255,N_17210);
xnor U17728 (N_17728,N_17283,N_17338);
or U17729 (N_17729,N_17505,N_17582);
or U17730 (N_17730,N_17465,N_17273);
nand U17731 (N_17731,N_17231,N_17299);
nor U17732 (N_17732,N_17250,N_17381);
and U17733 (N_17733,N_17206,N_17528);
or U17734 (N_17734,N_17463,N_17415);
nand U17735 (N_17735,N_17400,N_17490);
xor U17736 (N_17736,N_17324,N_17473);
or U17737 (N_17737,N_17541,N_17316);
and U17738 (N_17738,N_17329,N_17594);
nor U17739 (N_17739,N_17291,N_17500);
xor U17740 (N_17740,N_17267,N_17470);
or U17741 (N_17741,N_17569,N_17300);
and U17742 (N_17742,N_17454,N_17261);
xnor U17743 (N_17743,N_17422,N_17483);
and U17744 (N_17744,N_17409,N_17225);
xor U17745 (N_17745,N_17265,N_17522);
or U17746 (N_17746,N_17552,N_17222);
or U17747 (N_17747,N_17204,N_17356);
nand U17748 (N_17748,N_17526,N_17548);
nor U17749 (N_17749,N_17535,N_17353);
nand U17750 (N_17750,N_17508,N_17343);
nor U17751 (N_17751,N_17596,N_17260);
xor U17752 (N_17752,N_17359,N_17364);
or U17753 (N_17753,N_17558,N_17464);
xor U17754 (N_17754,N_17437,N_17346);
nor U17755 (N_17755,N_17370,N_17592);
nand U17756 (N_17756,N_17433,N_17544);
and U17757 (N_17757,N_17448,N_17585);
or U17758 (N_17758,N_17220,N_17575);
xnor U17759 (N_17759,N_17485,N_17527);
nand U17760 (N_17760,N_17280,N_17207);
and U17761 (N_17761,N_17599,N_17297);
nor U17762 (N_17762,N_17262,N_17335);
nand U17763 (N_17763,N_17545,N_17289);
or U17764 (N_17764,N_17554,N_17357);
nand U17765 (N_17765,N_17428,N_17480);
nor U17766 (N_17766,N_17491,N_17332);
nor U17767 (N_17767,N_17339,N_17279);
or U17768 (N_17768,N_17573,N_17404);
nor U17769 (N_17769,N_17537,N_17328);
and U17770 (N_17770,N_17281,N_17560);
xnor U17771 (N_17771,N_17201,N_17420);
nor U17772 (N_17772,N_17208,N_17525);
nand U17773 (N_17773,N_17572,N_17507);
or U17774 (N_17774,N_17479,N_17388);
xor U17775 (N_17775,N_17309,N_17203);
nand U17776 (N_17776,N_17304,N_17440);
nand U17777 (N_17777,N_17216,N_17252);
or U17778 (N_17778,N_17446,N_17589);
or U17779 (N_17779,N_17408,N_17254);
and U17780 (N_17780,N_17239,N_17436);
xnor U17781 (N_17781,N_17486,N_17577);
and U17782 (N_17782,N_17462,N_17570);
xor U17783 (N_17783,N_17455,N_17205);
nand U17784 (N_17784,N_17264,N_17240);
nor U17785 (N_17785,N_17243,N_17471);
or U17786 (N_17786,N_17434,N_17546);
or U17787 (N_17787,N_17333,N_17461);
nor U17788 (N_17788,N_17382,N_17321);
nand U17789 (N_17789,N_17543,N_17411);
or U17790 (N_17790,N_17595,N_17482);
nor U17791 (N_17791,N_17286,N_17584);
and U17792 (N_17792,N_17564,N_17540);
xor U17793 (N_17793,N_17523,N_17447);
xor U17794 (N_17794,N_17567,N_17513);
nor U17795 (N_17795,N_17439,N_17489);
nand U17796 (N_17796,N_17251,N_17218);
nand U17797 (N_17797,N_17256,N_17547);
or U17798 (N_17798,N_17284,N_17293);
nor U17799 (N_17799,N_17249,N_17506);
and U17800 (N_17800,N_17268,N_17569);
or U17801 (N_17801,N_17396,N_17280);
nand U17802 (N_17802,N_17569,N_17453);
and U17803 (N_17803,N_17364,N_17467);
nor U17804 (N_17804,N_17374,N_17258);
nand U17805 (N_17805,N_17407,N_17486);
and U17806 (N_17806,N_17343,N_17421);
xor U17807 (N_17807,N_17358,N_17339);
nor U17808 (N_17808,N_17585,N_17493);
and U17809 (N_17809,N_17224,N_17521);
nand U17810 (N_17810,N_17430,N_17517);
or U17811 (N_17811,N_17361,N_17253);
xor U17812 (N_17812,N_17347,N_17491);
xnor U17813 (N_17813,N_17507,N_17513);
xor U17814 (N_17814,N_17472,N_17437);
xor U17815 (N_17815,N_17353,N_17474);
or U17816 (N_17816,N_17315,N_17360);
and U17817 (N_17817,N_17553,N_17216);
xor U17818 (N_17818,N_17235,N_17244);
nand U17819 (N_17819,N_17540,N_17293);
and U17820 (N_17820,N_17357,N_17581);
nor U17821 (N_17821,N_17413,N_17306);
and U17822 (N_17822,N_17426,N_17482);
or U17823 (N_17823,N_17249,N_17521);
xnor U17824 (N_17824,N_17327,N_17218);
and U17825 (N_17825,N_17269,N_17320);
or U17826 (N_17826,N_17377,N_17531);
and U17827 (N_17827,N_17345,N_17243);
and U17828 (N_17828,N_17379,N_17333);
and U17829 (N_17829,N_17416,N_17501);
nand U17830 (N_17830,N_17411,N_17447);
nand U17831 (N_17831,N_17290,N_17590);
or U17832 (N_17832,N_17575,N_17354);
nor U17833 (N_17833,N_17546,N_17598);
nor U17834 (N_17834,N_17231,N_17323);
xnor U17835 (N_17835,N_17597,N_17306);
xnor U17836 (N_17836,N_17452,N_17592);
and U17837 (N_17837,N_17381,N_17574);
or U17838 (N_17838,N_17484,N_17532);
or U17839 (N_17839,N_17326,N_17283);
and U17840 (N_17840,N_17214,N_17348);
xnor U17841 (N_17841,N_17427,N_17520);
nand U17842 (N_17842,N_17260,N_17342);
nand U17843 (N_17843,N_17445,N_17227);
xnor U17844 (N_17844,N_17325,N_17206);
or U17845 (N_17845,N_17213,N_17527);
nor U17846 (N_17846,N_17499,N_17483);
xor U17847 (N_17847,N_17537,N_17279);
nor U17848 (N_17848,N_17228,N_17202);
nor U17849 (N_17849,N_17303,N_17569);
or U17850 (N_17850,N_17352,N_17245);
nor U17851 (N_17851,N_17537,N_17346);
nor U17852 (N_17852,N_17544,N_17200);
nor U17853 (N_17853,N_17479,N_17305);
and U17854 (N_17854,N_17581,N_17497);
nand U17855 (N_17855,N_17260,N_17465);
or U17856 (N_17856,N_17487,N_17286);
and U17857 (N_17857,N_17244,N_17358);
nor U17858 (N_17858,N_17285,N_17371);
or U17859 (N_17859,N_17390,N_17576);
nor U17860 (N_17860,N_17584,N_17578);
nor U17861 (N_17861,N_17570,N_17213);
nor U17862 (N_17862,N_17396,N_17361);
xor U17863 (N_17863,N_17320,N_17371);
and U17864 (N_17864,N_17513,N_17358);
and U17865 (N_17865,N_17407,N_17310);
nand U17866 (N_17866,N_17415,N_17263);
nor U17867 (N_17867,N_17467,N_17465);
and U17868 (N_17868,N_17431,N_17522);
or U17869 (N_17869,N_17293,N_17340);
and U17870 (N_17870,N_17296,N_17290);
or U17871 (N_17871,N_17360,N_17530);
nand U17872 (N_17872,N_17398,N_17446);
nor U17873 (N_17873,N_17228,N_17550);
nor U17874 (N_17874,N_17410,N_17538);
nand U17875 (N_17875,N_17319,N_17394);
or U17876 (N_17876,N_17587,N_17282);
or U17877 (N_17877,N_17217,N_17398);
or U17878 (N_17878,N_17306,N_17382);
nand U17879 (N_17879,N_17333,N_17313);
nand U17880 (N_17880,N_17308,N_17446);
and U17881 (N_17881,N_17483,N_17341);
and U17882 (N_17882,N_17573,N_17334);
nor U17883 (N_17883,N_17485,N_17456);
or U17884 (N_17884,N_17514,N_17274);
and U17885 (N_17885,N_17395,N_17285);
and U17886 (N_17886,N_17526,N_17465);
or U17887 (N_17887,N_17401,N_17519);
nand U17888 (N_17888,N_17216,N_17380);
nand U17889 (N_17889,N_17489,N_17227);
nand U17890 (N_17890,N_17462,N_17223);
and U17891 (N_17891,N_17214,N_17547);
nor U17892 (N_17892,N_17494,N_17580);
and U17893 (N_17893,N_17504,N_17249);
nor U17894 (N_17894,N_17526,N_17515);
xnor U17895 (N_17895,N_17509,N_17319);
xor U17896 (N_17896,N_17583,N_17407);
nor U17897 (N_17897,N_17264,N_17571);
or U17898 (N_17898,N_17475,N_17279);
nor U17899 (N_17899,N_17487,N_17409);
xor U17900 (N_17900,N_17509,N_17580);
and U17901 (N_17901,N_17531,N_17414);
xor U17902 (N_17902,N_17437,N_17429);
nand U17903 (N_17903,N_17532,N_17494);
nor U17904 (N_17904,N_17259,N_17210);
xor U17905 (N_17905,N_17438,N_17267);
xor U17906 (N_17906,N_17462,N_17324);
xnor U17907 (N_17907,N_17539,N_17565);
xor U17908 (N_17908,N_17556,N_17572);
or U17909 (N_17909,N_17387,N_17301);
and U17910 (N_17910,N_17398,N_17394);
xor U17911 (N_17911,N_17597,N_17582);
or U17912 (N_17912,N_17577,N_17497);
or U17913 (N_17913,N_17371,N_17393);
nand U17914 (N_17914,N_17390,N_17569);
xor U17915 (N_17915,N_17331,N_17335);
nor U17916 (N_17916,N_17458,N_17529);
or U17917 (N_17917,N_17242,N_17548);
and U17918 (N_17918,N_17330,N_17303);
or U17919 (N_17919,N_17208,N_17443);
and U17920 (N_17920,N_17445,N_17374);
or U17921 (N_17921,N_17554,N_17431);
nor U17922 (N_17922,N_17573,N_17418);
nand U17923 (N_17923,N_17419,N_17380);
xor U17924 (N_17924,N_17540,N_17421);
nand U17925 (N_17925,N_17280,N_17544);
nand U17926 (N_17926,N_17214,N_17347);
nor U17927 (N_17927,N_17433,N_17517);
and U17928 (N_17928,N_17329,N_17314);
nand U17929 (N_17929,N_17376,N_17530);
nor U17930 (N_17930,N_17243,N_17393);
xor U17931 (N_17931,N_17353,N_17449);
nor U17932 (N_17932,N_17266,N_17423);
nor U17933 (N_17933,N_17561,N_17244);
nor U17934 (N_17934,N_17341,N_17386);
xnor U17935 (N_17935,N_17460,N_17293);
xnor U17936 (N_17936,N_17407,N_17580);
or U17937 (N_17937,N_17287,N_17270);
nor U17938 (N_17938,N_17442,N_17210);
nor U17939 (N_17939,N_17351,N_17380);
and U17940 (N_17940,N_17470,N_17511);
nand U17941 (N_17941,N_17459,N_17349);
and U17942 (N_17942,N_17509,N_17298);
nand U17943 (N_17943,N_17324,N_17572);
nand U17944 (N_17944,N_17474,N_17530);
xor U17945 (N_17945,N_17237,N_17378);
nand U17946 (N_17946,N_17327,N_17535);
nand U17947 (N_17947,N_17549,N_17443);
xor U17948 (N_17948,N_17246,N_17454);
nor U17949 (N_17949,N_17235,N_17274);
and U17950 (N_17950,N_17496,N_17255);
xnor U17951 (N_17951,N_17324,N_17318);
xor U17952 (N_17952,N_17479,N_17549);
and U17953 (N_17953,N_17557,N_17570);
and U17954 (N_17954,N_17283,N_17267);
nor U17955 (N_17955,N_17361,N_17372);
or U17956 (N_17956,N_17495,N_17202);
nand U17957 (N_17957,N_17241,N_17593);
xor U17958 (N_17958,N_17450,N_17347);
or U17959 (N_17959,N_17559,N_17545);
or U17960 (N_17960,N_17235,N_17424);
nor U17961 (N_17961,N_17436,N_17340);
xnor U17962 (N_17962,N_17459,N_17362);
xor U17963 (N_17963,N_17317,N_17484);
xnor U17964 (N_17964,N_17206,N_17563);
nor U17965 (N_17965,N_17598,N_17451);
and U17966 (N_17966,N_17311,N_17391);
and U17967 (N_17967,N_17350,N_17270);
and U17968 (N_17968,N_17273,N_17494);
nor U17969 (N_17969,N_17517,N_17586);
nor U17970 (N_17970,N_17546,N_17301);
nor U17971 (N_17971,N_17255,N_17559);
xor U17972 (N_17972,N_17546,N_17268);
or U17973 (N_17973,N_17350,N_17592);
nor U17974 (N_17974,N_17478,N_17294);
or U17975 (N_17975,N_17331,N_17333);
nand U17976 (N_17976,N_17251,N_17572);
and U17977 (N_17977,N_17548,N_17348);
and U17978 (N_17978,N_17311,N_17598);
nand U17979 (N_17979,N_17393,N_17409);
nand U17980 (N_17980,N_17209,N_17454);
and U17981 (N_17981,N_17550,N_17449);
or U17982 (N_17982,N_17254,N_17487);
and U17983 (N_17983,N_17394,N_17239);
xor U17984 (N_17984,N_17264,N_17267);
xor U17985 (N_17985,N_17352,N_17407);
and U17986 (N_17986,N_17290,N_17491);
and U17987 (N_17987,N_17547,N_17340);
and U17988 (N_17988,N_17477,N_17213);
or U17989 (N_17989,N_17424,N_17489);
xor U17990 (N_17990,N_17320,N_17571);
or U17991 (N_17991,N_17213,N_17313);
xor U17992 (N_17992,N_17350,N_17516);
xor U17993 (N_17993,N_17234,N_17569);
or U17994 (N_17994,N_17355,N_17447);
and U17995 (N_17995,N_17538,N_17568);
xor U17996 (N_17996,N_17492,N_17260);
and U17997 (N_17997,N_17316,N_17271);
xnor U17998 (N_17998,N_17364,N_17275);
nor U17999 (N_17999,N_17500,N_17441);
or U18000 (N_18000,N_17812,N_17694);
and U18001 (N_18001,N_17933,N_17729);
nand U18002 (N_18002,N_17703,N_17761);
nand U18003 (N_18003,N_17604,N_17633);
or U18004 (N_18004,N_17940,N_17914);
nand U18005 (N_18005,N_17774,N_17639);
nand U18006 (N_18006,N_17712,N_17759);
or U18007 (N_18007,N_17810,N_17615);
or U18008 (N_18008,N_17884,N_17936);
and U18009 (N_18009,N_17800,N_17885);
nand U18010 (N_18010,N_17726,N_17880);
nand U18011 (N_18011,N_17620,N_17609);
or U18012 (N_18012,N_17792,N_17765);
nor U18013 (N_18013,N_17887,N_17695);
nor U18014 (N_18014,N_17938,N_17777);
nor U18015 (N_18015,N_17716,N_17822);
or U18016 (N_18016,N_17986,N_17912);
or U18017 (N_18017,N_17809,N_17919);
and U18018 (N_18018,N_17966,N_17668);
nand U18019 (N_18019,N_17814,N_17913);
xnor U18020 (N_18020,N_17920,N_17711);
nand U18021 (N_18021,N_17956,N_17975);
and U18022 (N_18022,N_17652,N_17926);
nor U18023 (N_18023,N_17861,N_17798);
nor U18024 (N_18024,N_17826,N_17917);
and U18025 (N_18025,N_17793,N_17728);
xor U18026 (N_18026,N_17710,N_17719);
and U18027 (N_18027,N_17803,N_17746);
or U18028 (N_18028,N_17757,N_17795);
xor U18029 (N_18029,N_17611,N_17631);
or U18030 (N_18030,N_17907,N_17738);
nor U18031 (N_18031,N_17651,N_17752);
xor U18032 (N_18032,N_17829,N_17871);
xor U18033 (N_18033,N_17808,N_17960);
and U18034 (N_18034,N_17699,N_17778);
and U18035 (N_18035,N_17982,N_17863);
xor U18036 (N_18036,N_17762,N_17906);
or U18037 (N_18037,N_17649,N_17794);
or U18038 (N_18038,N_17613,N_17769);
nor U18039 (N_18039,N_17819,N_17655);
nand U18040 (N_18040,N_17721,N_17677);
nand U18041 (N_18041,N_17605,N_17980);
and U18042 (N_18042,N_17953,N_17689);
xnor U18043 (N_18043,N_17748,N_17916);
and U18044 (N_18044,N_17663,N_17676);
nand U18045 (N_18045,N_17805,N_17678);
xor U18046 (N_18046,N_17867,N_17709);
and U18047 (N_18047,N_17976,N_17790);
and U18048 (N_18048,N_17934,N_17755);
or U18049 (N_18049,N_17847,N_17999);
or U18050 (N_18050,N_17931,N_17944);
and U18051 (N_18051,N_17619,N_17600);
nor U18052 (N_18052,N_17828,N_17618);
nand U18053 (N_18053,N_17879,N_17830);
nor U18054 (N_18054,N_17942,N_17791);
nand U18055 (N_18055,N_17891,N_17985);
nand U18056 (N_18056,N_17993,N_17606);
or U18057 (N_18057,N_17905,N_17693);
or U18058 (N_18058,N_17969,N_17626);
and U18059 (N_18059,N_17722,N_17915);
nor U18060 (N_18060,N_17687,N_17742);
xnor U18061 (N_18061,N_17786,N_17804);
and U18062 (N_18062,N_17700,N_17785);
or U18063 (N_18063,N_17967,N_17799);
nor U18064 (N_18064,N_17839,N_17682);
and U18065 (N_18065,N_17691,N_17841);
or U18066 (N_18066,N_17674,N_17856);
nor U18067 (N_18067,N_17997,N_17852);
and U18068 (N_18068,N_17770,N_17753);
and U18069 (N_18069,N_17834,N_17971);
and U18070 (N_18070,N_17987,N_17702);
nor U18071 (N_18071,N_17869,N_17989);
nor U18072 (N_18072,N_17662,N_17882);
nand U18073 (N_18073,N_17837,N_17959);
or U18074 (N_18074,N_17733,N_17947);
or U18075 (N_18075,N_17961,N_17789);
and U18076 (N_18076,N_17876,N_17925);
or U18077 (N_18077,N_17634,N_17801);
nor U18078 (N_18078,N_17815,N_17763);
or U18079 (N_18079,N_17945,N_17979);
or U18080 (N_18080,N_17610,N_17771);
nand U18081 (N_18081,N_17889,N_17664);
nand U18082 (N_18082,N_17675,N_17918);
nor U18083 (N_18083,N_17602,N_17783);
or U18084 (N_18084,N_17843,N_17737);
nor U18085 (N_18085,N_17855,N_17653);
nand U18086 (N_18086,N_17624,N_17643);
nand U18087 (N_18087,N_17892,N_17622);
xnor U18088 (N_18088,N_17696,N_17990);
xor U18089 (N_18089,N_17848,N_17977);
nand U18090 (N_18090,N_17734,N_17706);
or U18091 (N_18091,N_17921,N_17740);
nor U18092 (N_18092,N_17928,N_17692);
nand U18093 (N_18093,N_17648,N_17788);
xnor U18094 (N_18094,N_17645,N_17779);
xor U18095 (N_18095,N_17948,N_17909);
xnor U18096 (N_18096,N_17661,N_17628);
nor U18097 (N_18097,N_17608,N_17806);
nand U18098 (N_18098,N_17713,N_17784);
or U18099 (N_18099,N_17875,N_17756);
xor U18100 (N_18100,N_17900,N_17881);
xnor U18101 (N_18101,N_17865,N_17883);
and U18102 (N_18102,N_17923,N_17950);
or U18103 (N_18103,N_17686,N_17911);
xnor U18104 (N_18104,N_17717,N_17616);
or U18105 (N_18105,N_17660,N_17886);
or U18106 (N_18106,N_17874,N_17854);
or U18107 (N_18107,N_17954,N_17750);
and U18108 (N_18108,N_17970,N_17864);
or U18109 (N_18109,N_17817,N_17782);
xnor U18110 (N_18110,N_17772,N_17902);
nand U18111 (N_18111,N_17644,N_17690);
xnor U18112 (N_18112,N_17893,N_17813);
or U18113 (N_18113,N_17701,N_17858);
or U18114 (N_18114,N_17768,N_17868);
or U18115 (N_18115,N_17727,N_17697);
nor U18116 (N_18116,N_17603,N_17908);
xor U18117 (N_18117,N_17894,N_17866);
and U18118 (N_18118,N_17995,N_17963);
and U18119 (N_18119,N_17787,N_17637);
and U18120 (N_18120,N_17983,N_17988);
or U18121 (N_18121,N_17650,N_17705);
and U18122 (N_18122,N_17601,N_17898);
or U18123 (N_18123,N_17679,N_17965);
or U18124 (N_18124,N_17978,N_17922);
xnor U18125 (N_18125,N_17846,N_17754);
nor U18126 (N_18126,N_17932,N_17835);
nor U18127 (N_18127,N_17924,N_17658);
xnor U18128 (N_18128,N_17903,N_17941);
nor U18129 (N_18129,N_17635,N_17743);
nand U18130 (N_18130,N_17760,N_17665);
nor U18131 (N_18131,N_17910,N_17720);
and U18132 (N_18132,N_17897,N_17758);
nor U18133 (N_18133,N_17850,N_17797);
and U18134 (N_18134,N_17824,N_17952);
nand U18135 (N_18135,N_17998,N_17974);
or U18136 (N_18136,N_17838,N_17749);
and U18137 (N_18137,N_17968,N_17972);
or U18138 (N_18138,N_17832,N_17935);
nor U18139 (N_18139,N_17672,N_17816);
nand U18140 (N_18140,N_17849,N_17831);
and U18141 (N_18141,N_17642,N_17714);
nor U18142 (N_18142,N_17811,N_17647);
nor U18143 (N_18143,N_17825,N_17707);
or U18144 (N_18144,N_17612,N_17853);
nor U18145 (N_18145,N_17641,N_17764);
nor U18146 (N_18146,N_17607,N_17833);
or U18147 (N_18147,N_17736,N_17984);
and U18148 (N_18148,N_17827,N_17957);
xnor U18149 (N_18149,N_17745,N_17636);
nor U18150 (N_18150,N_17870,N_17654);
nand U18151 (N_18151,N_17730,N_17646);
or U18152 (N_18152,N_17860,N_17776);
and U18153 (N_18153,N_17739,N_17895);
or U18154 (N_18154,N_17890,N_17981);
nand U18155 (N_18155,N_17684,N_17669);
or U18156 (N_18156,N_17878,N_17704);
and U18157 (N_18157,N_17766,N_17751);
and U18158 (N_18158,N_17623,N_17744);
or U18159 (N_18159,N_17996,N_17741);
and U18160 (N_18160,N_17630,N_17773);
and U18161 (N_18161,N_17943,N_17632);
or U18162 (N_18162,N_17873,N_17946);
and U18163 (N_18163,N_17735,N_17780);
nand U18164 (N_18164,N_17899,N_17930);
or U18165 (N_18165,N_17857,N_17617);
or U18166 (N_18166,N_17964,N_17877);
or U18167 (N_18167,N_17939,N_17724);
nand U18168 (N_18168,N_17973,N_17732);
nand U18169 (N_18169,N_17802,N_17680);
or U18170 (N_18170,N_17842,N_17821);
nor U18171 (N_18171,N_17656,N_17851);
nand U18172 (N_18172,N_17673,N_17951);
nand U18173 (N_18173,N_17614,N_17796);
nor U18174 (N_18174,N_17807,N_17955);
and U18175 (N_18175,N_17823,N_17991);
nor U18176 (N_18176,N_17725,N_17767);
nor U18177 (N_18177,N_17840,N_17698);
and U18178 (N_18178,N_17671,N_17992);
and U18179 (N_18179,N_17901,N_17844);
or U18180 (N_18180,N_17775,N_17927);
or U18181 (N_18181,N_17627,N_17888);
xnor U18182 (N_18182,N_17681,N_17929);
xor U18183 (N_18183,N_17862,N_17949);
nand U18184 (N_18184,N_17820,N_17638);
and U18185 (N_18185,N_17708,N_17781);
and U18186 (N_18186,N_17621,N_17629);
or U18187 (N_18187,N_17625,N_17688);
nand U18188 (N_18188,N_17723,N_17937);
or U18189 (N_18189,N_17872,N_17896);
and U18190 (N_18190,N_17715,N_17845);
or U18191 (N_18191,N_17718,N_17670);
or U18192 (N_18192,N_17666,N_17994);
and U18193 (N_18193,N_17685,N_17657);
and U18194 (N_18194,N_17659,N_17683);
nor U18195 (N_18195,N_17859,N_17747);
nor U18196 (N_18196,N_17836,N_17731);
nand U18197 (N_18197,N_17640,N_17818);
xnor U18198 (N_18198,N_17962,N_17667);
or U18199 (N_18199,N_17958,N_17904);
nor U18200 (N_18200,N_17711,N_17627);
nor U18201 (N_18201,N_17770,N_17784);
nand U18202 (N_18202,N_17755,N_17705);
xor U18203 (N_18203,N_17671,N_17676);
and U18204 (N_18204,N_17906,N_17671);
and U18205 (N_18205,N_17879,N_17612);
nor U18206 (N_18206,N_17684,N_17774);
nor U18207 (N_18207,N_17880,N_17785);
nor U18208 (N_18208,N_17816,N_17779);
or U18209 (N_18209,N_17738,N_17649);
nor U18210 (N_18210,N_17874,N_17803);
nor U18211 (N_18211,N_17865,N_17712);
and U18212 (N_18212,N_17693,N_17708);
nor U18213 (N_18213,N_17775,N_17854);
nor U18214 (N_18214,N_17977,N_17726);
and U18215 (N_18215,N_17789,N_17705);
or U18216 (N_18216,N_17718,N_17706);
nand U18217 (N_18217,N_17709,N_17835);
and U18218 (N_18218,N_17905,N_17959);
nand U18219 (N_18219,N_17867,N_17647);
and U18220 (N_18220,N_17769,N_17829);
or U18221 (N_18221,N_17604,N_17895);
or U18222 (N_18222,N_17810,N_17898);
nand U18223 (N_18223,N_17612,N_17674);
or U18224 (N_18224,N_17871,N_17959);
or U18225 (N_18225,N_17659,N_17965);
xor U18226 (N_18226,N_17873,N_17966);
nor U18227 (N_18227,N_17610,N_17676);
and U18228 (N_18228,N_17662,N_17625);
nand U18229 (N_18229,N_17836,N_17789);
xor U18230 (N_18230,N_17762,N_17895);
and U18231 (N_18231,N_17644,N_17840);
or U18232 (N_18232,N_17957,N_17787);
or U18233 (N_18233,N_17812,N_17829);
nand U18234 (N_18234,N_17621,N_17854);
or U18235 (N_18235,N_17642,N_17946);
nand U18236 (N_18236,N_17792,N_17672);
xnor U18237 (N_18237,N_17973,N_17759);
nor U18238 (N_18238,N_17795,N_17664);
nor U18239 (N_18239,N_17938,N_17941);
xor U18240 (N_18240,N_17907,N_17960);
xnor U18241 (N_18241,N_17957,N_17613);
nor U18242 (N_18242,N_17738,N_17679);
or U18243 (N_18243,N_17912,N_17875);
nor U18244 (N_18244,N_17776,N_17830);
xnor U18245 (N_18245,N_17892,N_17739);
nor U18246 (N_18246,N_17977,N_17644);
and U18247 (N_18247,N_17673,N_17911);
nor U18248 (N_18248,N_17882,N_17664);
xnor U18249 (N_18249,N_17609,N_17782);
nor U18250 (N_18250,N_17603,N_17824);
or U18251 (N_18251,N_17853,N_17872);
nor U18252 (N_18252,N_17890,N_17864);
or U18253 (N_18253,N_17934,N_17992);
nor U18254 (N_18254,N_17959,N_17976);
xnor U18255 (N_18255,N_17697,N_17716);
nor U18256 (N_18256,N_17742,N_17927);
nand U18257 (N_18257,N_17642,N_17890);
nand U18258 (N_18258,N_17624,N_17877);
xor U18259 (N_18259,N_17791,N_17649);
and U18260 (N_18260,N_17721,N_17748);
xor U18261 (N_18261,N_17603,N_17877);
xnor U18262 (N_18262,N_17957,N_17820);
or U18263 (N_18263,N_17786,N_17907);
or U18264 (N_18264,N_17800,N_17742);
or U18265 (N_18265,N_17643,N_17605);
and U18266 (N_18266,N_17845,N_17641);
and U18267 (N_18267,N_17734,N_17827);
nor U18268 (N_18268,N_17876,N_17737);
nand U18269 (N_18269,N_17964,N_17952);
and U18270 (N_18270,N_17851,N_17711);
and U18271 (N_18271,N_17711,N_17988);
or U18272 (N_18272,N_17726,N_17997);
nand U18273 (N_18273,N_17852,N_17637);
xnor U18274 (N_18274,N_17668,N_17918);
nor U18275 (N_18275,N_17828,N_17678);
xor U18276 (N_18276,N_17699,N_17697);
xnor U18277 (N_18277,N_17929,N_17634);
nor U18278 (N_18278,N_17816,N_17634);
and U18279 (N_18279,N_17788,N_17740);
nand U18280 (N_18280,N_17671,N_17990);
xor U18281 (N_18281,N_17610,N_17795);
and U18282 (N_18282,N_17980,N_17937);
nor U18283 (N_18283,N_17669,N_17861);
nand U18284 (N_18284,N_17915,N_17601);
xor U18285 (N_18285,N_17933,N_17777);
xor U18286 (N_18286,N_17649,N_17686);
xnor U18287 (N_18287,N_17965,N_17948);
or U18288 (N_18288,N_17906,N_17760);
nand U18289 (N_18289,N_17925,N_17619);
xor U18290 (N_18290,N_17858,N_17865);
or U18291 (N_18291,N_17848,N_17858);
xor U18292 (N_18292,N_17731,N_17637);
and U18293 (N_18293,N_17728,N_17979);
nor U18294 (N_18294,N_17728,N_17743);
xor U18295 (N_18295,N_17944,N_17930);
or U18296 (N_18296,N_17653,N_17939);
xor U18297 (N_18297,N_17939,N_17980);
nand U18298 (N_18298,N_17752,N_17634);
or U18299 (N_18299,N_17686,N_17679);
nand U18300 (N_18300,N_17934,N_17665);
and U18301 (N_18301,N_17759,N_17772);
and U18302 (N_18302,N_17665,N_17870);
or U18303 (N_18303,N_17674,N_17959);
nor U18304 (N_18304,N_17818,N_17616);
and U18305 (N_18305,N_17753,N_17734);
or U18306 (N_18306,N_17944,N_17811);
xnor U18307 (N_18307,N_17959,N_17737);
or U18308 (N_18308,N_17802,N_17949);
and U18309 (N_18309,N_17676,N_17935);
and U18310 (N_18310,N_17683,N_17705);
xor U18311 (N_18311,N_17972,N_17948);
nor U18312 (N_18312,N_17608,N_17918);
and U18313 (N_18313,N_17649,N_17736);
nand U18314 (N_18314,N_17731,N_17953);
and U18315 (N_18315,N_17762,N_17809);
or U18316 (N_18316,N_17751,N_17842);
or U18317 (N_18317,N_17661,N_17741);
xnor U18318 (N_18318,N_17893,N_17640);
nand U18319 (N_18319,N_17718,N_17973);
and U18320 (N_18320,N_17854,N_17980);
xor U18321 (N_18321,N_17959,N_17966);
or U18322 (N_18322,N_17811,N_17737);
or U18323 (N_18323,N_17662,N_17981);
or U18324 (N_18324,N_17795,N_17612);
xor U18325 (N_18325,N_17993,N_17726);
nor U18326 (N_18326,N_17915,N_17712);
xnor U18327 (N_18327,N_17954,N_17843);
xor U18328 (N_18328,N_17671,N_17761);
xor U18329 (N_18329,N_17688,N_17994);
or U18330 (N_18330,N_17677,N_17899);
nor U18331 (N_18331,N_17793,N_17637);
nor U18332 (N_18332,N_17977,N_17732);
nor U18333 (N_18333,N_17829,N_17996);
nand U18334 (N_18334,N_17632,N_17627);
and U18335 (N_18335,N_17832,N_17877);
and U18336 (N_18336,N_17817,N_17652);
xnor U18337 (N_18337,N_17970,N_17626);
xor U18338 (N_18338,N_17985,N_17864);
nor U18339 (N_18339,N_17782,N_17850);
or U18340 (N_18340,N_17617,N_17791);
nor U18341 (N_18341,N_17644,N_17946);
nand U18342 (N_18342,N_17715,N_17731);
nand U18343 (N_18343,N_17921,N_17745);
xor U18344 (N_18344,N_17968,N_17641);
or U18345 (N_18345,N_17625,N_17717);
or U18346 (N_18346,N_17691,N_17975);
nand U18347 (N_18347,N_17626,N_17745);
or U18348 (N_18348,N_17775,N_17801);
xnor U18349 (N_18349,N_17753,N_17769);
or U18350 (N_18350,N_17885,N_17922);
xnor U18351 (N_18351,N_17781,N_17930);
nand U18352 (N_18352,N_17965,N_17747);
and U18353 (N_18353,N_17636,N_17948);
and U18354 (N_18354,N_17744,N_17826);
and U18355 (N_18355,N_17611,N_17889);
nor U18356 (N_18356,N_17620,N_17777);
nor U18357 (N_18357,N_17608,N_17683);
xor U18358 (N_18358,N_17942,N_17871);
or U18359 (N_18359,N_17617,N_17953);
xor U18360 (N_18360,N_17880,N_17664);
or U18361 (N_18361,N_17738,N_17905);
and U18362 (N_18362,N_17848,N_17647);
xnor U18363 (N_18363,N_17861,N_17865);
or U18364 (N_18364,N_17655,N_17931);
or U18365 (N_18365,N_17756,N_17991);
nor U18366 (N_18366,N_17877,N_17916);
or U18367 (N_18367,N_17837,N_17807);
nand U18368 (N_18368,N_17782,N_17858);
xnor U18369 (N_18369,N_17920,N_17780);
xnor U18370 (N_18370,N_17684,N_17843);
or U18371 (N_18371,N_17900,N_17722);
or U18372 (N_18372,N_17658,N_17618);
nand U18373 (N_18373,N_17729,N_17725);
or U18374 (N_18374,N_17870,N_17854);
or U18375 (N_18375,N_17745,N_17809);
and U18376 (N_18376,N_17657,N_17956);
nand U18377 (N_18377,N_17680,N_17681);
or U18378 (N_18378,N_17641,N_17636);
nor U18379 (N_18379,N_17663,N_17798);
and U18380 (N_18380,N_17679,N_17972);
nand U18381 (N_18381,N_17853,N_17755);
or U18382 (N_18382,N_17888,N_17620);
and U18383 (N_18383,N_17684,N_17787);
and U18384 (N_18384,N_17851,N_17664);
nor U18385 (N_18385,N_17928,N_17662);
nor U18386 (N_18386,N_17623,N_17841);
xor U18387 (N_18387,N_17936,N_17650);
xor U18388 (N_18388,N_17806,N_17935);
nor U18389 (N_18389,N_17903,N_17759);
nor U18390 (N_18390,N_17696,N_17655);
xor U18391 (N_18391,N_17657,N_17887);
and U18392 (N_18392,N_17940,N_17728);
xor U18393 (N_18393,N_17747,N_17947);
and U18394 (N_18394,N_17732,N_17853);
xor U18395 (N_18395,N_17647,N_17791);
xnor U18396 (N_18396,N_17685,N_17686);
and U18397 (N_18397,N_17772,N_17973);
nand U18398 (N_18398,N_17903,N_17790);
nor U18399 (N_18399,N_17626,N_17912);
or U18400 (N_18400,N_18278,N_18204);
or U18401 (N_18401,N_18324,N_18337);
nor U18402 (N_18402,N_18057,N_18352);
xor U18403 (N_18403,N_18085,N_18111);
xor U18404 (N_18404,N_18081,N_18275);
nand U18405 (N_18405,N_18092,N_18136);
and U18406 (N_18406,N_18163,N_18312);
or U18407 (N_18407,N_18225,N_18280);
and U18408 (N_18408,N_18130,N_18331);
nor U18409 (N_18409,N_18372,N_18226);
xnor U18410 (N_18410,N_18082,N_18314);
xnor U18411 (N_18411,N_18313,N_18380);
nor U18412 (N_18412,N_18270,N_18018);
or U18413 (N_18413,N_18129,N_18320);
nand U18414 (N_18414,N_18151,N_18247);
or U18415 (N_18415,N_18044,N_18309);
or U18416 (N_18416,N_18118,N_18393);
and U18417 (N_18417,N_18308,N_18124);
xor U18418 (N_18418,N_18268,N_18282);
and U18419 (N_18419,N_18015,N_18119);
nor U18420 (N_18420,N_18233,N_18166);
and U18421 (N_18421,N_18104,N_18061);
nand U18422 (N_18422,N_18031,N_18169);
or U18423 (N_18423,N_18115,N_18367);
and U18424 (N_18424,N_18388,N_18302);
nor U18425 (N_18425,N_18060,N_18279);
and U18426 (N_18426,N_18301,N_18340);
and U18427 (N_18427,N_18284,N_18200);
nand U18428 (N_18428,N_18055,N_18250);
nor U18429 (N_18429,N_18028,N_18013);
nand U18430 (N_18430,N_18235,N_18298);
nand U18431 (N_18431,N_18207,N_18223);
xor U18432 (N_18432,N_18170,N_18229);
nand U18433 (N_18433,N_18135,N_18276);
nor U18434 (N_18434,N_18287,N_18106);
nor U18435 (N_18435,N_18215,N_18024);
nor U18436 (N_18436,N_18142,N_18096);
nor U18437 (N_18437,N_18358,N_18160);
nor U18438 (N_18438,N_18064,N_18232);
and U18439 (N_18439,N_18213,N_18152);
or U18440 (N_18440,N_18334,N_18330);
nand U18441 (N_18441,N_18240,N_18054);
nand U18442 (N_18442,N_18265,N_18019);
xnor U18443 (N_18443,N_18214,N_18039);
nor U18444 (N_18444,N_18267,N_18147);
and U18445 (N_18445,N_18362,N_18156);
and U18446 (N_18446,N_18040,N_18212);
or U18447 (N_18447,N_18183,N_18059);
or U18448 (N_18448,N_18333,N_18236);
xor U18449 (N_18449,N_18074,N_18038);
and U18450 (N_18450,N_18006,N_18237);
and U18451 (N_18451,N_18153,N_18255);
or U18452 (N_18452,N_18014,N_18037);
and U18453 (N_18453,N_18205,N_18101);
nand U18454 (N_18454,N_18084,N_18264);
nor U18455 (N_18455,N_18016,N_18231);
or U18456 (N_18456,N_18257,N_18043);
nor U18457 (N_18457,N_18272,N_18379);
and U18458 (N_18458,N_18385,N_18297);
or U18459 (N_18459,N_18188,N_18208);
nor U18460 (N_18460,N_18258,N_18290);
nor U18461 (N_18461,N_18179,N_18194);
nor U18462 (N_18462,N_18398,N_18149);
and U18463 (N_18463,N_18004,N_18027);
nand U18464 (N_18464,N_18088,N_18274);
and U18465 (N_18465,N_18002,N_18076);
nor U18466 (N_18466,N_18343,N_18198);
nor U18467 (N_18467,N_18116,N_18351);
nand U18468 (N_18468,N_18220,N_18306);
xor U18469 (N_18469,N_18349,N_18000);
nand U18470 (N_18470,N_18245,N_18269);
xnor U18471 (N_18471,N_18359,N_18080);
nand U18472 (N_18472,N_18023,N_18341);
nand U18473 (N_18473,N_18300,N_18020);
nor U18474 (N_18474,N_18346,N_18374);
nand U18475 (N_18475,N_18176,N_18067);
xnor U18476 (N_18476,N_18056,N_18286);
and U18477 (N_18477,N_18073,N_18174);
or U18478 (N_18478,N_18065,N_18012);
and U18479 (N_18479,N_18053,N_18354);
nor U18480 (N_18480,N_18097,N_18386);
nand U18481 (N_18481,N_18253,N_18008);
xor U18482 (N_18482,N_18103,N_18172);
and U18483 (N_18483,N_18248,N_18397);
xnor U18484 (N_18484,N_18100,N_18140);
nand U18485 (N_18485,N_18090,N_18036);
and U18486 (N_18486,N_18357,N_18191);
and U18487 (N_18487,N_18126,N_18078);
or U18488 (N_18488,N_18001,N_18178);
nor U18489 (N_18489,N_18234,N_18102);
and U18490 (N_18490,N_18022,N_18339);
nand U18491 (N_18491,N_18062,N_18161);
and U18492 (N_18492,N_18109,N_18068);
xor U18493 (N_18493,N_18224,N_18238);
and U18494 (N_18494,N_18157,N_18295);
xor U18495 (N_18495,N_18009,N_18291);
or U18496 (N_18496,N_18273,N_18182);
xor U18497 (N_18497,N_18026,N_18196);
and U18498 (N_18498,N_18158,N_18221);
nor U18499 (N_18499,N_18377,N_18294);
xnor U18500 (N_18500,N_18303,N_18107);
xnor U18501 (N_18501,N_18353,N_18370);
nand U18502 (N_18502,N_18148,N_18384);
xnor U18503 (N_18503,N_18190,N_18133);
xor U18504 (N_18504,N_18378,N_18335);
or U18505 (N_18505,N_18243,N_18112);
and U18506 (N_18506,N_18329,N_18373);
or U18507 (N_18507,N_18350,N_18021);
or U18508 (N_18508,N_18093,N_18193);
nor U18509 (N_18509,N_18391,N_18167);
nor U18510 (N_18510,N_18371,N_18277);
nand U18511 (N_18511,N_18171,N_18177);
and U18512 (N_18512,N_18033,N_18134);
nand U18513 (N_18513,N_18047,N_18241);
or U18514 (N_18514,N_18260,N_18363);
nand U18515 (N_18515,N_18222,N_18077);
and U18516 (N_18516,N_18396,N_18328);
xnor U18517 (N_18517,N_18127,N_18387);
nor U18518 (N_18518,N_18010,N_18089);
and U18519 (N_18519,N_18360,N_18262);
and U18520 (N_18520,N_18138,N_18035);
nor U18521 (N_18521,N_18128,N_18319);
nor U18522 (N_18522,N_18311,N_18304);
nand U18523 (N_18523,N_18154,N_18338);
nand U18524 (N_18524,N_18075,N_18123);
xor U18525 (N_18525,N_18117,N_18283);
nor U18526 (N_18526,N_18095,N_18189);
and U18527 (N_18527,N_18246,N_18389);
nor U18528 (N_18528,N_18249,N_18292);
nor U18529 (N_18529,N_18087,N_18228);
nand U18530 (N_18530,N_18361,N_18242);
xnor U18531 (N_18531,N_18293,N_18121);
and U18532 (N_18532,N_18072,N_18356);
or U18533 (N_18533,N_18239,N_18227);
xor U18534 (N_18534,N_18321,N_18390);
nand U18535 (N_18535,N_18203,N_18155);
nand U18536 (N_18536,N_18098,N_18299);
and U18537 (N_18537,N_18122,N_18165);
and U18538 (N_18538,N_18305,N_18187);
nand U18539 (N_18539,N_18323,N_18144);
and U18540 (N_18540,N_18162,N_18394);
nor U18541 (N_18541,N_18114,N_18046);
xor U18542 (N_18542,N_18066,N_18316);
nor U18543 (N_18543,N_18281,N_18355);
nand U18544 (N_18544,N_18288,N_18184);
nor U18545 (N_18545,N_18254,N_18108);
or U18546 (N_18546,N_18086,N_18164);
nor U18547 (N_18547,N_18202,N_18342);
nor U18548 (N_18548,N_18141,N_18201);
xnor U18549 (N_18549,N_18199,N_18327);
nand U18550 (N_18550,N_18375,N_18345);
and U18551 (N_18551,N_18271,N_18218);
xnor U18552 (N_18552,N_18094,N_18381);
or U18553 (N_18553,N_18105,N_18051);
nand U18554 (N_18554,N_18025,N_18261);
and U18555 (N_18555,N_18139,N_18326);
nor U18556 (N_18556,N_18070,N_18091);
or U18557 (N_18557,N_18307,N_18083);
or U18558 (N_18558,N_18052,N_18071);
or U18559 (N_18559,N_18192,N_18173);
and U18560 (N_18560,N_18206,N_18315);
and U18561 (N_18561,N_18032,N_18244);
and U18562 (N_18562,N_18211,N_18181);
and U18563 (N_18563,N_18030,N_18079);
or U18564 (N_18564,N_18034,N_18366);
nand U18565 (N_18565,N_18058,N_18132);
or U18566 (N_18566,N_18364,N_18150);
nand U18567 (N_18567,N_18063,N_18125);
nand U18568 (N_18568,N_18318,N_18003);
xor U18569 (N_18569,N_18344,N_18365);
nand U18570 (N_18570,N_18099,N_18113);
xor U18571 (N_18571,N_18143,N_18263);
xnor U18572 (N_18572,N_18145,N_18131);
nand U18573 (N_18573,N_18029,N_18209);
or U18574 (N_18574,N_18042,N_18045);
xor U18575 (N_18575,N_18168,N_18219);
xnor U18576 (N_18576,N_18050,N_18399);
xnor U18577 (N_18577,N_18383,N_18216);
nor U18578 (N_18578,N_18069,N_18317);
or U18579 (N_18579,N_18146,N_18252);
or U18580 (N_18580,N_18049,N_18266);
nor U18581 (N_18581,N_18048,N_18382);
nand U18582 (N_18582,N_18348,N_18336);
and U18583 (N_18583,N_18137,N_18011);
or U18584 (N_18584,N_18322,N_18180);
or U18585 (N_18585,N_18175,N_18259);
xnor U18586 (N_18586,N_18392,N_18251);
xor U18587 (N_18587,N_18368,N_18159);
and U18588 (N_18588,N_18007,N_18195);
nand U18589 (N_18589,N_18017,N_18296);
nor U18590 (N_18590,N_18120,N_18332);
or U18591 (N_18591,N_18041,N_18395);
nand U18592 (N_18592,N_18197,N_18376);
and U18593 (N_18593,N_18005,N_18210);
nor U18594 (N_18594,N_18285,N_18325);
xor U18595 (N_18595,N_18289,N_18186);
or U18596 (N_18596,N_18185,N_18110);
xor U18597 (N_18597,N_18230,N_18217);
nor U18598 (N_18598,N_18369,N_18310);
xnor U18599 (N_18599,N_18256,N_18347);
nor U18600 (N_18600,N_18365,N_18369);
xor U18601 (N_18601,N_18032,N_18214);
and U18602 (N_18602,N_18299,N_18352);
nor U18603 (N_18603,N_18044,N_18343);
xnor U18604 (N_18604,N_18326,N_18327);
xor U18605 (N_18605,N_18029,N_18327);
and U18606 (N_18606,N_18171,N_18367);
nand U18607 (N_18607,N_18291,N_18347);
or U18608 (N_18608,N_18314,N_18109);
nand U18609 (N_18609,N_18103,N_18038);
xor U18610 (N_18610,N_18014,N_18363);
nor U18611 (N_18611,N_18030,N_18000);
nor U18612 (N_18612,N_18292,N_18296);
nor U18613 (N_18613,N_18019,N_18157);
or U18614 (N_18614,N_18384,N_18294);
and U18615 (N_18615,N_18134,N_18119);
and U18616 (N_18616,N_18300,N_18136);
or U18617 (N_18617,N_18232,N_18211);
xnor U18618 (N_18618,N_18281,N_18186);
nor U18619 (N_18619,N_18280,N_18356);
xnor U18620 (N_18620,N_18322,N_18109);
nand U18621 (N_18621,N_18296,N_18378);
or U18622 (N_18622,N_18219,N_18171);
nand U18623 (N_18623,N_18150,N_18191);
xor U18624 (N_18624,N_18190,N_18358);
or U18625 (N_18625,N_18168,N_18174);
nand U18626 (N_18626,N_18238,N_18048);
nand U18627 (N_18627,N_18307,N_18100);
or U18628 (N_18628,N_18126,N_18363);
and U18629 (N_18629,N_18021,N_18318);
xnor U18630 (N_18630,N_18133,N_18340);
nand U18631 (N_18631,N_18281,N_18153);
nor U18632 (N_18632,N_18162,N_18110);
nor U18633 (N_18633,N_18268,N_18278);
xor U18634 (N_18634,N_18089,N_18121);
nor U18635 (N_18635,N_18365,N_18384);
xor U18636 (N_18636,N_18262,N_18006);
or U18637 (N_18637,N_18301,N_18335);
and U18638 (N_18638,N_18283,N_18378);
or U18639 (N_18639,N_18061,N_18108);
xor U18640 (N_18640,N_18366,N_18179);
xor U18641 (N_18641,N_18317,N_18050);
xor U18642 (N_18642,N_18381,N_18133);
xor U18643 (N_18643,N_18112,N_18382);
nor U18644 (N_18644,N_18024,N_18139);
or U18645 (N_18645,N_18165,N_18281);
nand U18646 (N_18646,N_18202,N_18104);
or U18647 (N_18647,N_18343,N_18084);
or U18648 (N_18648,N_18068,N_18060);
and U18649 (N_18649,N_18139,N_18111);
and U18650 (N_18650,N_18259,N_18181);
and U18651 (N_18651,N_18396,N_18299);
or U18652 (N_18652,N_18302,N_18268);
and U18653 (N_18653,N_18106,N_18102);
or U18654 (N_18654,N_18138,N_18384);
or U18655 (N_18655,N_18080,N_18132);
nand U18656 (N_18656,N_18368,N_18033);
nor U18657 (N_18657,N_18301,N_18154);
nand U18658 (N_18658,N_18383,N_18333);
nor U18659 (N_18659,N_18320,N_18072);
nor U18660 (N_18660,N_18205,N_18095);
or U18661 (N_18661,N_18270,N_18086);
or U18662 (N_18662,N_18248,N_18297);
or U18663 (N_18663,N_18309,N_18022);
nor U18664 (N_18664,N_18289,N_18315);
and U18665 (N_18665,N_18340,N_18079);
nand U18666 (N_18666,N_18114,N_18379);
nor U18667 (N_18667,N_18058,N_18161);
or U18668 (N_18668,N_18148,N_18214);
and U18669 (N_18669,N_18339,N_18261);
nand U18670 (N_18670,N_18168,N_18261);
nor U18671 (N_18671,N_18375,N_18370);
or U18672 (N_18672,N_18297,N_18342);
or U18673 (N_18673,N_18020,N_18010);
xor U18674 (N_18674,N_18056,N_18204);
nor U18675 (N_18675,N_18304,N_18392);
xnor U18676 (N_18676,N_18332,N_18090);
or U18677 (N_18677,N_18204,N_18025);
nand U18678 (N_18678,N_18061,N_18263);
xnor U18679 (N_18679,N_18209,N_18336);
nand U18680 (N_18680,N_18005,N_18004);
or U18681 (N_18681,N_18383,N_18208);
nand U18682 (N_18682,N_18080,N_18229);
xnor U18683 (N_18683,N_18190,N_18163);
nor U18684 (N_18684,N_18098,N_18018);
and U18685 (N_18685,N_18362,N_18174);
nand U18686 (N_18686,N_18225,N_18089);
nor U18687 (N_18687,N_18190,N_18165);
nand U18688 (N_18688,N_18374,N_18370);
nand U18689 (N_18689,N_18137,N_18047);
nand U18690 (N_18690,N_18262,N_18037);
nor U18691 (N_18691,N_18001,N_18367);
and U18692 (N_18692,N_18079,N_18347);
nand U18693 (N_18693,N_18332,N_18284);
nor U18694 (N_18694,N_18300,N_18256);
and U18695 (N_18695,N_18379,N_18241);
and U18696 (N_18696,N_18147,N_18248);
nand U18697 (N_18697,N_18139,N_18014);
nor U18698 (N_18698,N_18301,N_18166);
nor U18699 (N_18699,N_18104,N_18249);
nand U18700 (N_18700,N_18250,N_18312);
or U18701 (N_18701,N_18289,N_18200);
or U18702 (N_18702,N_18029,N_18175);
and U18703 (N_18703,N_18289,N_18394);
and U18704 (N_18704,N_18398,N_18236);
or U18705 (N_18705,N_18001,N_18073);
or U18706 (N_18706,N_18172,N_18293);
xor U18707 (N_18707,N_18032,N_18057);
nand U18708 (N_18708,N_18295,N_18228);
xnor U18709 (N_18709,N_18097,N_18211);
or U18710 (N_18710,N_18228,N_18227);
xnor U18711 (N_18711,N_18240,N_18208);
nor U18712 (N_18712,N_18358,N_18140);
xnor U18713 (N_18713,N_18303,N_18227);
xnor U18714 (N_18714,N_18290,N_18392);
xor U18715 (N_18715,N_18311,N_18055);
or U18716 (N_18716,N_18337,N_18339);
nand U18717 (N_18717,N_18022,N_18328);
nor U18718 (N_18718,N_18351,N_18313);
nand U18719 (N_18719,N_18320,N_18378);
nand U18720 (N_18720,N_18297,N_18176);
xor U18721 (N_18721,N_18329,N_18270);
or U18722 (N_18722,N_18170,N_18226);
xnor U18723 (N_18723,N_18360,N_18217);
nand U18724 (N_18724,N_18223,N_18009);
nor U18725 (N_18725,N_18351,N_18057);
xor U18726 (N_18726,N_18354,N_18317);
or U18727 (N_18727,N_18205,N_18137);
or U18728 (N_18728,N_18311,N_18334);
xnor U18729 (N_18729,N_18067,N_18213);
and U18730 (N_18730,N_18137,N_18397);
nand U18731 (N_18731,N_18361,N_18077);
or U18732 (N_18732,N_18164,N_18229);
and U18733 (N_18733,N_18141,N_18080);
nand U18734 (N_18734,N_18043,N_18028);
and U18735 (N_18735,N_18287,N_18208);
nand U18736 (N_18736,N_18325,N_18234);
xnor U18737 (N_18737,N_18202,N_18261);
nand U18738 (N_18738,N_18299,N_18084);
xor U18739 (N_18739,N_18265,N_18164);
and U18740 (N_18740,N_18069,N_18357);
xor U18741 (N_18741,N_18167,N_18206);
xnor U18742 (N_18742,N_18068,N_18156);
or U18743 (N_18743,N_18331,N_18150);
xnor U18744 (N_18744,N_18185,N_18317);
and U18745 (N_18745,N_18176,N_18330);
and U18746 (N_18746,N_18293,N_18301);
xor U18747 (N_18747,N_18160,N_18132);
or U18748 (N_18748,N_18213,N_18187);
nand U18749 (N_18749,N_18037,N_18043);
and U18750 (N_18750,N_18062,N_18374);
or U18751 (N_18751,N_18224,N_18176);
or U18752 (N_18752,N_18038,N_18012);
nor U18753 (N_18753,N_18038,N_18309);
or U18754 (N_18754,N_18206,N_18076);
or U18755 (N_18755,N_18199,N_18003);
xnor U18756 (N_18756,N_18298,N_18126);
nand U18757 (N_18757,N_18211,N_18303);
nand U18758 (N_18758,N_18257,N_18399);
or U18759 (N_18759,N_18300,N_18108);
nand U18760 (N_18760,N_18342,N_18175);
nor U18761 (N_18761,N_18149,N_18331);
nand U18762 (N_18762,N_18358,N_18376);
or U18763 (N_18763,N_18031,N_18103);
xnor U18764 (N_18764,N_18336,N_18207);
and U18765 (N_18765,N_18261,N_18177);
nor U18766 (N_18766,N_18056,N_18067);
or U18767 (N_18767,N_18339,N_18249);
xnor U18768 (N_18768,N_18283,N_18040);
nor U18769 (N_18769,N_18358,N_18032);
nand U18770 (N_18770,N_18043,N_18053);
xnor U18771 (N_18771,N_18298,N_18165);
nand U18772 (N_18772,N_18123,N_18127);
and U18773 (N_18773,N_18113,N_18044);
and U18774 (N_18774,N_18309,N_18399);
and U18775 (N_18775,N_18109,N_18369);
xor U18776 (N_18776,N_18373,N_18395);
nor U18777 (N_18777,N_18033,N_18001);
nand U18778 (N_18778,N_18012,N_18244);
xnor U18779 (N_18779,N_18008,N_18296);
or U18780 (N_18780,N_18015,N_18236);
or U18781 (N_18781,N_18157,N_18154);
nor U18782 (N_18782,N_18044,N_18019);
xnor U18783 (N_18783,N_18182,N_18082);
or U18784 (N_18784,N_18267,N_18046);
nor U18785 (N_18785,N_18313,N_18220);
nand U18786 (N_18786,N_18316,N_18389);
or U18787 (N_18787,N_18115,N_18387);
and U18788 (N_18788,N_18202,N_18350);
or U18789 (N_18789,N_18111,N_18220);
xnor U18790 (N_18790,N_18359,N_18274);
nand U18791 (N_18791,N_18272,N_18011);
nor U18792 (N_18792,N_18097,N_18041);
xnor U18793 (N_18793,N_18323,N_18271);
or U18794 (N_18794,N_18121,N_18225);
nand U18795 (N_18795,N_18041,N_18234);
xnor U18796 (N_18796,N_18169,N_18376);
nor U18797 (N_18797,N_18188,N_18075);
nand U18798 (N_18798,N_18311,N_18343);
and U18799 (N_18799,N_18132,N_18025);
xor U18800 (N_18800,N_18418,N_18565);
xnor U18801 (N_18801,N_18653,N_18505);
nand U18802 (N_18802,N_18544,N_18726);
and U18803 (N_18803,N_18623,N_18710);
nand U18804 (N_18804,N_18468,N_18508);
or U18805 (N_18805,N_18717,N_18546);
xnor U18806 (N_18806,N_18563,N_18682);
nand U18807 (N_18807,N_18756,N_18687);
xnor U18808 (N_18808,N_18621,N_18777);
xnor U18809 (N_18809,N_18643,N_18734);
xor U18810 (N_18810,N_18600,N_18690);
nor U18811 (N_18811,N_18752,N_18470);
nor U18812 (N_18812,N_18666,N_18438);
and U18813 (N_18813,N_18521,N_18665);
nor U18814 (N_18814,N_18591,N_18489);
or U18815 (N_18815,N_18780,N_18748);
nand U18816 (N_18816,N_18555,N_18564);
nor U18817 (N_18817,N_18675,N_18459);
xnor U18818 (N_18818,N_18608,N_18631);
nand U18819 (N_18819,N_18523,N_18495);
nor U18820 (N_18820,N_18624,N_18746);
nor U18821 (N_18821,N_18498,N_18609);
nand U18822 (N_18822,N_18703,N_18541);
nor U18823 (N_18823,N_18730,N_18688);
xnor U18824 (N_18824,N_18640,N_18674);
or U18825 (N_18825,N_18502,N_18437);
nor U18826 (N_18826,N_18434,N_18407);
nand U18827 (N_18827,N_18693,N_18751);
or U18828 (N_18828,N_18798,N_18700);
xnor U18829 (N_18829,N_18651,N_18558);
and U18830 (N_18830,N_18614,N_18712);
or U18831 (N_18831,N_18694,N_18663);
nand U18832 (N_18832,N_18709,N_18695);
nor U18833 (N_18833,N_18552,N_18528);
nand U18834 (N_18834,N_18644,N_18585);
xor U18835 (N_18835,N_18778,N_18457);
or U18836 (N_18836,N_18629,N_18618);
nand U18837 (N_18837,N_18739,N_18537);
or U18838 (N_18838,N_18536,N_18602);
nor U18839 (N_18839,N_18707,N_18765);
nand U18840 (N_18840,N_18613,N_18701);
nand U18841 (N_18841,N_18553,N_18714);
xnor U18842 (N_18842,N_18641,N_18500);
or U18843 (N_18843,N_18779,N_18401);
or U18844 (N_18844,N_18454,N_18477);
xor U18845 (N_18845,N_18603,N_18652);
or U18846 (N_18846,N_18622,N_18711);
and U18847 (N_18847,N_18584,N_18781);
xnor U18848 (N_18848,N_18415,N_18556);
and U18849 (N_18849,N_18636,N_18784);
nand U18850 (N_18850,N_18607,N_18706);
and U18851 (N_18851,N_18638,N_18503);
nor U18852 (N_18852,N_18554,N_18429);
nand U18853 (N_18853,N_18460,N_18642);
xor U18854 (N_18854,N_18490,N_18514);
nand U18855 (N_18855,N_18594,N_18569);
and U18856 (N_18856,N_18443,N_18557);
or U18857 (N_18857,N_18635,N_18626);
nand U18858 (N_18858,N_18518,N_18658);
nand U18859 (N_18859,N_18743,N_18462);
nand U18860 (N_18860,N_18672,N_18504);
nor U18861 (N_18861,N_18705,N_18562);
nand U18862 (N_18862,N_18661,N_18570);
and U18863 (N_18863,N_18450,N_18561);
and U18864 (N_18864,N_18577,N_18659);
nor U18865 (N_18865,N_18439,N_18704);
and U18866 (N_18866,N_18729,N_18794);
or U18867 (N_18867,N_18491,N_18595);
xnor U18868 (N_18868,N_18582,N_18680);
and U18869 (N_18869,N_18573,N_18479);
xnor U18870 (N_18870,N_18417,N_18435);
nand U18871 (N_18871,N_18612,N_18493);
or U18872 (N_18872,N_18539,N_18551);
and U18873 (N_18873,N_18416,N_18755);
nand U18874 (N_18874,N_18764,N_18782);
or U18875 (N_18875,N_18722,N_18534);
and U18876 (N_18876,N_18409,N_18408);
nor U18877 (N_18877,N_18689,N_18447);
xnor U18878 (N_18878,N_18678,N_18766);
nand U18879 (N_18879,N_18444,N_18797);
nor U18880 (N_18880,N_18696,N_18630);
and U18881 (N_18881,N_18520,N_18679);
nand U18882 (N_18882,N_18719,N_18428);
nand U18883 (N_18883,N_18610,N_18749);
xnor U18884 (N_18884,N_18547,N_18527);
and U18885 (N_18885,N_18402,N_18483);
xnor U18886 (N_18886,N_18420,N_18458);
nand U18887 (N_18887,N_18436,N_18785);
and U18888 (N_18888,N_18583,N_18526);
nand U18889 (N_18889,N_18725,N_18761);
and U18890 (N_18890,N_18512,N_18617);
nor U18891 (N_18891,N_18426,N_18686);
nand U18892 (N_18892,N_18519,N_18713);
or U18893 (N_18893,N_18799,N_18431);
nand U18894 (N_18894,N_18550,N_18627);
nand U18895 (N_18895,N_18720,N_18654);
or U18896 (N_18896,N_18571,N_18511);
nor U18897 (N_18897,N_18773,N_18501);
or U18898 (N_18898,N_18792,N_18646);
nor U18899 (N_18899,N_18474,N_18510);
or U18900 (N_18900,N_18593,N_18759);
nand U18901 (N_18901,N_18760,N_18795);
xor U18902 (N_18902,N_18545,N_18449);
xor U18903 (N_18903,N_18455,N_18716);
or U18904 (N_18904,N_18668,N_18422);
and U18905 (N_18905,N_18620,N_18586);
and U18906 (N_18906,N_18655,N_18667);
xor U18907 (N_18907,N_18715,N_18403);
and U18908 (N_18908,N_18669,N_18647);
xor U18909 (N_18909,N_18513,N_18763);
or U18910 (N_18910,N_18578,N_18699);
or U18911 (N_18911,N_18522,N_18660);
or U18912 (N_18912,N_18702,N_18619);
or U18913 (N_18913,N_18517,N_18531);
nand U18914 (N_18914,N_18588,N_18597);
or U18915 (N_18915,N_18639,N_18440);
nor U18916 (N_18916,N_18697,N_18737);
nand U18917 (N_18917,N_18463,N_18579);
and U18918 (N_18918,N_18492,N_18718);
or U18919 (N_18919,N_18676,N_18506);
or U18920 (N_18920,N_18405,N_18775);
xnor U18921 (N_18921,N_18538,N_18671);
nand U18922 (N_18922,N_18472,N_18615);
xnor U18923 (N_18923,N_18733,N_18411);
or U18924 (N_18924,N_18410,N_18776);
nand U18925 (N_18925,N_18721,N_18406);
or U18926 (N_18926,N_18736,N_18657);
nand U18927 (N_18927,N_18485,N_18587);
and U18928 (N_18928,N_18482,N_18762);
nor U18929 (N_18929,N_18633,N_18589);
xnor U18930 (N_18930,N_18632,N_18580);
nor U18931 (N_18931,N_18499,N_18481);
xnor U18932 (N_18932,N_18559,N_18464);
nor U18933 (N_18933,N_18576,N_18480);
nand U18934 (N_18934,N_18788,N_18413);
xor U18935 (N_18935,N_18745,N_18423);
nand U18936 (N_18936,N_18786,N_18471);
nor U18937 (N_18937,N_18724,N_18598);
nand U18938 (N_18938,N_18771,N_18461);
or U18939 (N_18939,N_18656,N_18533);
and U18940 (N_18940,N_18476,N_18441);
nor U18941 (N_18941,N_18478,N_18758);
nand U18942 (N_18942,N_18601,N_18445);
or U18943 (N_18943,N_18497,N_18708);
xnor U18944 (N_18944,N_18685,N_18516);
and U18945 (N_18945,N_18424,N_18590);
or U18946 (N_18946,N_18469,N_18728);
and U18947 (N_18947,N_18404,N_18494);
xnor U18948 (N_18948,N_18525,N_18419);
xor U18949 (N_18949,N_18540,N_18684);
xor U18950 (N_18950,N_18560,N_18484);
nand U18951 (N_18951,N_18543,N_18496);
or U18952 (N_18952,N_18548,N_18448);
nor U18953 (N_18953,N_18568,N_18605);
nor U18954 (N_18954,N_18466,N_18670);
and U18955 (N_18955,N_18524,N_18787);
nor U18956 (N_18956,N_18673,N_18731);
nand U18957 (N_18957,N_18465,N_18599);
nand U18958 (N_18958,N_18529,N_18637);
and U18959 (N_18959,N_18427,N_18768);
and U18960 (N_18960,N_18430,N_18453);
nor U18961 (N_18961,N_18698,N_18446);
xor U18962 (N_18962,N_18604,N_18596);
nand U18963 (N_18963,N_18475,N_18488);
nor U18964 (N_18964,N_18509,N_18634);
or U18965 (N_18965,N_18772,N_18515);
nand U18966 (N_18966,N_18451,N_18567);
nand U18967 (N_18967,N_18467,N_18606);
xnor U18968 (N_18968,N_18433,N_18796);
nand U18969 (N_18969,N_18432,N_18683);
nand U18970 (N_18970,N_18611,N_18425);
nor U18971 (N_18971,N_18753,N_18592);
xnor U18972 (N_18972,N_18532,N_18530);
nor U18973 (N_18973,N_18727,N_18645);
xnor U18974 (N_18974,N_18616,N_18790);
nand U18975 (N_18975,N_18648,N_18757);
or U18976 (N_18976,N_18750,N_18754);
and U18977 (N_18977,N_18791,N_18740);
xor U18978 (N_18978,N_18662,N_18649);
xor U18979 (N_18979,N_18507,N_18770);
xor U18980 (N_18980,N_18542,N_18572);
or U18981 (N_18981,N_18723,N_18677);
nor U18982 (N_18982,N_18783,N_18735);
xnor U18983 (N_18983,N_18625,N_18774);
or U18984 (N_18984,N_18575,N_18793);
nand U18985 (N_18985,N_18566,N_18664);
nor U18986 (N_18986,N_18628,N_18442);
nand U18987 (N_18987,N_18747,N_18581);
nand U18988 (N_18988,N_18412,N_18742);
nand U18989 (N_18989,N_18744,N_18414);
nand U18990 (N_18990,N_18769,N_18486);
nor U18991 (N_18991,N_18452,N_18535);
nand U18992 (N_18992,N_18681,N_18421);
or U18993 (N_18993,N_18456,N_18741);
xnor U18994 (N_18994,N_18738,N_18549);
or U18995 (N_18995,N_18650,N_18487);
nor U18996 (N_18996,N_18767,N_18400);
xnor U18997 (N_18997,N_18574,N_18732);
and U18998 (N_18998,N_18692,N_18789);
nor U18999 (N_18999,N_18473,N_18691);
nand U19000 (N_19000,N_18659,N_18562);
xnor U19001 (N_19001,N_18785,N_18454);
xor U19002 (N_19002,N_18727,N_18730);
and U19003 (N_19003,N_18570,N_18471);
and U19004 (N_19004,N_18408,N_18663);
nor U19005 (N_19005,N_18494,N_18684);
and U19006 (N_19006,N_18476,N_18505);
xor U19007 (N_19007,N_18505,N_18432);
nor U19008 (N_19008,N_18498,N_18544);
nor U19009 (N_19009,N_18420,N_18691);
nand U19010 (N_19010,N_18787,N_18516);
xor U19011 (N_19011,N_18446,N_18460);
nand U19012 (N_19012,N_18521,N_18490);
and U19013 (N_19013,N_18694,N_18659);
xnor U19014 (N_19014,N_18477,N_18754);
nor U19015 (N_19015,N_18656,N_18400);
nor U19016 (N_19016,N_18635,N_18652);
xor U19017 (N_19017,N_18683,N_18720);
xnor U19018 (N_19018,N_18475,N_18473);
or U19019 (N_19019,N_18474,N_18490);
nor U19020 (N_19020,N_18763,N_18538);
xor U19021 (N_19021,N_18639,N_18467);
nor U19022 (N_19022,N_18589,N_18425);
and U19023 (N_19023,N_18718,N_18523);
nand U19024 (N_19024,N_18693,N_18432);
nand U19025 (N_19025,N_18405,N_18487);
nand U19026 (N_19026,N_18714,N_18508);
nor U19027 (N_19027,N_18526,N_18773);
and U19028 (N_19028,N_18544,N_18612);
nand U19029 (N_19029,N_18770,N_18615);
or U19030 (N_19030,N_18708,N_18553);
nor U19031 (N_19031,N_18441,N_18760);
or U19032 (N_19032,N_18760,N_18474);
xnor U19033 (N_19033,N_18778,N_18667);
nor U19034 (N_19034,N_18576,N_18443);
and U19035 (N_19035,N_18501,N_18706);
xnor U19036 (N_19036,N_18771,N_18619);
nor U19037 (N_19037,N_18554,N_18567);
and U19038 (N_19038,N_18631,N_18667);
or U19039 (N_19039,N_18455,N_18608);
or U19040 (N_19040,N_18581,N_18432);
xnor U19041 (N_19041,N_18693,N_18673);
nor U19042 (N_19042,N_18499,N_18466);
nor U19043 (N_19043,N_18682,N_18754);
nand U19044 (N_19044,N_18492,N_18665);
nand U19045 (N_19045,N_18587,N_18627);
and U19046 (N_19046,N_18794,N_18727);
nor U19047 (N_19047,N_18588,N_18771);
nor U19048 (N_19048,N_18696,N_18451);
xnor U19049 (N_19049,N_18637,N_18619);
nor U19050 (N_19050,N_18690,N_18530);
and U19051 (N_19051,N_18609,N_18728);
nand U19052 (N_19052,N_18550,N_18559);
xnor U19053 (N_19053,N_18529,N_18798);
nand U19054 (N_19054,N_18611,N_18498);
nor U19055 (N_19055,N_18572,N_18594);
xor U19056 (N_19056,N_18734,N_18613);
or U19057 (N_19057,N_18430,N_18770);
nor U19058 (N_19058,N_18560,N_18491);
xnor U19059 (N_19059,N_18757,N_18769);
and U19060 (N_19060,N_18512,N_18580);
nor U19061 (N_19061,N_18672,N_18698);
and U19062 (N_19062,N_18428,N_18796);
or U19063 (N_19063,N_18749,N_18475);
or U19064 (N_19064,N_18481,N_18554);
or U19065 (N_19065,N_18476,N_18784);
xnor U19066 (N_19066,N_18512,N_18716);
nand U19067 (N_19067,N_18627,N_18501);
or U19068 (N_19068,N_18625,N_18415);
xor U19069 (N_19069,N_18625,N_18649);
nor U19070 (N_19070,N_18743,N_18736);
nor U19071 (N_19071,N_18680,N_18665);
xnor U19072 (N_19072,N_18605,N_18612);
nand U19073 (N_19073,N_18557,N_18593);
and U19074 (N_19074,N_18539,N_18607);
nand U19075 (N_19075,N_18635,N_18729);
and U19076 (N_19076,N_18677,N_18513);
nand U19077 (N_19077,N_18685,N_18586);
and U19078 (N_19078,N_18483,N_18646);
or U19079 (N_19079,N_18595,N_18498);
nand U19080 (N_19080,N_18785,N_18570);
or U19081 (N_19081,N_18738,N_18620);
or U19082 (N_19082,N_18463,N_18679);
nor U19083 (N_19083,N_18407,N_18595);
xnor U19084 (N_19084,N_18529,N_18611);
nand U19085 (N_19085,N_18426,N_18501);
nand U19086 (N_19086,N_18714,N_18692);
or U19087 (N_19087,N_18759,N_18493);
or U19088 (N_19088,N_18769,N_18699);
xnor U19089 (N_19089,N_18450,N_18686);
or U19090 (N_19090,N_18753,N_18563);
nor U19091 (N_19091,N_18543,N_18706);
xor U19092 (N_19092,N_18449,N_18463);
xnor U19093 (N_19093,N_18604,N_18762);
xor U19094 (N_19094,N_18725,N_18713);
nand U19095 (N_19095,N_18499,N_18441);
and U19096 (N_19096,N_18420,N_18537);
nand U19097 (N_19097,N_18439,N_18731);
and U19098 (N_19098,N_18553,N_18690);
or U19099 (N_19099,N_18550,N_18720);
xor U19100 (N_19100,N_18627,N_18412);
or U19101 (N_19101,N_18754,N_18727);
nand U19102 (N_19102,N_18468,N_18611);
xor U19103 (N_19103,N_18407,N_18693);
nand U19104 (N_19104,N_18724,N_18455);
and U19105 (N_19105,N_18509,N_18458);
nor U19106 (N_19106,N_18727,N_18692);
nand U19107 (N_19107,N_18560,N_18414);
nand U19108 (N_19108,N_18416,N_18438);
nand U19109 (N_19109,N_18463,N_18481);
or U19110 (N_19110,N_18706,N_18764);
and U19111 (N_19111,N_18463,N_18733);
nand U19112 (N_19112,N_18621,N_18552);
xnor U19113 (N_19113,N_18592,N_18674);
or U19114 (N_19114,N_18464,N_18415);
and U19115 (N_19115,N_18541,N_18583);
xor U19116 (N_19116,N_18777,N_18693);
or U19117 (N_19117,N_18745,N_18519);
or U19118 (N_19118,N_18630,N_18570);
nand U19119 (N_19119,N_18640,N_18410);
nor U19120 (N_19120,N_18526,N_18635);
nand U19121 (N_19121,N_18517,N_18461);
or U19122 (N_19122,N_18479,N_18518);
nor U19123 (N_19123,N_18637,N_18729);
xor U19124 (N_19124,N_18690,N_18418);
nor U19125 (N_19125,N_18555,N_18569);
nand U19126 (N_19126,N_18486,N_18421);
xor U19127 (N_19127,N_18513,N_18787);
nand U19128 (N_19128,N_18590,N_18749);
nand U19129 (N_19129,N_18799,N_18726);
and U19130 (N_19130,N_18405,N_18771);
nor U19131 (N_19131,N_18611,N_18713);
nor U19132 (N_19132,N_18762,N_18661);
xnor U19133 (N_19133,N_18623,N_18741);
xnor U19134 (N_19134,N_18675,N_18799);
and U19135 (N_19135,N_18750,N_18576);
nor U19136 (N_19136,N_18588,N_18492);
and U19137 (N_19137,N_18500,N_18790);
nand U19138 (N_19138,N_18640,N_18505);
xor U19139 (N_19139,N_18457,N_18515);
and U19140 (N_19140,N_18428,N_18679);
nor U19141 (N_19141,N_18668,N_18484);
nand U19142 (N_19142,N_18672,N_18474);
xnor U19143 (N_19143,N_18533,N_18799);
xnor U19144 (N_19144,N_18797,N_18700);
or U19145 (N_19145,N_18662,N_18573);
nand U19146 (N_19146,N_18645,N_18631);
nor U19147 (N_19147,N_18542,N_18632);
or U19148 (N_19148,N_18575,N_18788);
nor U19149 (N_19149,N_18435,N_18485);
nor U19150 (N_19150,N_18446,N_18555);
and U19151 (N_19151,N_18636,N_18797);
nor U19152 (N_19152,N_18654,N_18556);
nand U19153 (N_19153,N_18711,N_18792);
and U19154 (N_19154,N_18591,N_18708);
and U19155 (N_19155,N_18515,N_18639);
or U19156 (N_19156,N_18445,N_18571);
or U19157 (N_19157,N_18400,N_18654);
nand U19158 (N_19158,N_18689,N_18703);
and U19159 (N_19159,N_18507,N_18591);
nand U19160 (N_19160,N_18533,N_18743);
nand U19161 (N_19161,N_18505,N_18478);
xor U19162 (N_19162,N_18714,N_18763);
or U19163 (N_19163,N_18408,N_18642);
and U19164 (N_19164,N_18476,N_18554);
nand U19165 (N_19165,N_18587,N_18471);
nor U19166 (N_19166,N_18623,N_18731);
nor U19167 (N_19167,N_18621,N_18699);
or U19168 (N_19168,N_18734,N_18648);
nor U19169 (N_19169,N_18521,N_18428);
or U19170 (N_19170,N_18439,N_18595);
nor U19171 (N_19171,N_18512,N_18430);
nor U19172 (N_19172,N_18645,N_18558);
nand U19173 (N_19173,N_18593,N_18796);
nor U19174 (N_19174,N_18601,N_18636);
nand U19175 (N_19175,N_18546,N_18593);
and U19176 (N_19176,N_18404,N_18731);
nand U19177 (N_19177,N_18646,N_18602);
nor U19178 (N_19178,N_18402,N_18407);
xnor U19179 (N_19179,N_18519,N_18799);
xor U19180 (N_19180,N_18556,N_18535);
and U19181 (N_19181,N_18662,N_18424);
xnor U19182 (N_19182,N_18707,N_18703);
nand U19183 (N_19183,N_18454,N_18715);
or U19184 (N_19184,N_18486,N_18733);
or U19185 (N_19185,N_18501,N_18781);
or U19186 (N_19186,N_18451,N_18440);
and U19187 (N_19187,N_18793,N_18751);
and U19188 (N_19188,N_18401,N_18776);
and U19189 (N_19189,N_18631,N_18724);
xor U19190 (N_19190,N_18550,N_18527);
nor U19191 (N_19191,N_18664,N_18595);
or U19192 (N_19192,N_18631,N_18415);
nor U19193 (N_19193,N_18624,N_18737);
nand U19194 (N_19194,N_18717,N_18507);
nor U19195 (N_19195,N_18488,N_18601);
nor U19196 (N_19196,N_18679,N_18518);
nor U19197 (N_19197,N_18722,N_18705);
xnor U19198 (N_19198,N_18440,N_18689);
xor U19199 (N_19199,N_18760,N_18627);
nand U19200 (N_19200,N_18873,N_19185);
and U19201 (N_19201,N_19001,N_18838);
or U19202 (N_19202,N_18827,N_19018);
nor U19203 (N_19203,N_18918,N_19186);
xor U19204 (N_19204,N_18969,N_19003);
nor U19205 (N_19205,N_18829,N_19140);
or U19206 (N_19206,N_18915,N_19089);
nor U19207 (N_19207,N_18992,N_18893);
or U19208 (N_19208,N_18804,N_18878);
nor U19209 (N_19209,N_18930,N_18863);
nand U19210 (N_19210,N_19025,N_18976);
or U19211 (N_19211,N_19170,N_19154);
nand U19212 (N_19212,N_18919,N_18937);
or U19213 (N_19213,N_19180,N_18948);
and U19214 (N_19214,N_18834,N_19147);
nor U19215 (N_19215,N_18995,N_19118);
or U19216 (N_19216,N_19188,N_18996);
or U19217 (N_19217,N_19100,N_19066);
nor U19218 (N_19218,N_19120,N_19062);
nor U19219 (N_19219,N_19189,N_19004);
and U19220 (N_19220,N_18901,N_18910);
or U19221 (N_19221,N_19096,N_19164);
and U19222 (N_19222,N_19023,N_18843);
nand U19223 (N_19223,N_18860,N_19184);
and U19224 (N_19224,N_19115,N_18884);
nor U19225 (N_19225,N_18891,N_19121);
xnor U19226 (N_19226,N_18876,N_18942);
xor U19227 (N_19227,N_19011,N_18984);
nor U19228 (N_19228,N_19074,N_18896);
nand U19229 (N_19229,N_19132,N_18957);
xnor U19230 (N_19230,N_19103,N_18862);
and U19231 (N_19231,N_19000,N_18831);
or U19232 (N_19232,N_18872,N_18926);
and U19233 (N_19233,N_19002,N_19080);
xor U19234 (N_19234,N_19053,N_18861);
xnor U19235 (N_19235,N_18908,N_18805);
xnor U19236 (N_19236,N_18857,N_19014);
or U19237 (N_19237,N_19171,N_19111);
nand U19238 (N_19238,N_19119,N_19155);
nor U19239 (N_19239,N_18979,N_19076);
or U19240 (N_19240,N_19077,N_19195);
xor U19241 (N_19241,N_19141,N_19144);
or U19242 (N_19242,N_18965,N_18989);
or U19243 (N_19243,N_19044,N_19050);
xor U19244 (N_19244,N_19047,N_19153);
nand U19245 (N_19245,N_19124,N_19090);
or U19246 (N_19246,N_18934,N_19084);
and U19247 (N_19247,N_18883,N_19095);
nor U19248 (N_19248,N_19159,N_19073);
nand U19249 (N_19249,N_19177,N_18801);
and U19250 (N_19250,N_19010,N_19058);
xnor U19251 (N_19251,N_18904,N_19085);
xnor U19252 (N_19252,N_19108,N_19029);
xor U19253 (N_19253,N_19143,N_18866);
nor U19254 (N_19254,N_19157,N_18899);
xnor U19255 (N_19255,N_18816,N_19190);
xnor U19256 (N_19256,N_18981,N_18824);
nand U19257 (N_19257,N_18837,N_18869);
xor U19258 (N_19258,N_18892,N_19040);
or U19259 (N_19259,N_19031,N_19110);
and U19260 (N_19260,N_19036,N_19021);
nand U19261 (N_19261,N_19113,N_18935);
nand U19262 (N_19262,N_18932,N_18875);
and U19263 (N_19263,N_19028,N_19024);
nand U19264 (N_19264,N_18975,N_18941);
nor U19265 (N_19265,N_19046,N_18944);
or U19266 (N_19266,N_18810,N_18821);
nor U19267 (N_19267,N_18972,N_18909);
nand U19268 (N_19268,N_18851,N_19160);
or U19269 (N_19269,N_18811,N_19032);
and U19270 (N_19270,N_18927,N_19105);
or U19271 (N_19271,N_18809,N_18895);
or U19272 (N_19272,N_18947,N_19059);
and U19273 (N_19273,N_18819,N_19161);
xor U19274 (N_19274,N_19052,N_19106);
nor U19275 (N_19275,N_18881,N_18840);
nor U19276 (N_19276,N_19149,N_19122);
or U19277 (N_19277,N_18980,N_19104);
and U19278 (N_19278,N_19199,N_19039);
and U19279 (N_19279,N_18839,N_18847);
nor U19280 (N_19280,N_18952,N_18822);
and U19281 (N_19281,N_18986,N_18897);
nand U19282 (N_19282,N_19043,N_19130);
xor U19283 (N_19283,N_19069,N_18983);
xnor U19284 (N_19284,N_19181,N_19131);
or U19285 (N_19285,N_18905,N_19087);
nand U19286 (N_19286,N_18921,N_18855);
and U19287 (N_19287,N_19129,N_19086);
and U19288 (N_19288,N_18998,N_18887);
or U19289 (N_19289,N_18939,N_18830);
and U19290 (N_19290,N_18828,N_18845);
xnor U19291 (N_19291,N_18867,N_18848);
and U19292 (N_19292,N_19030,N_19163);
nor U19293 (N_19293,N_18955,N_19006);
and U19294 (N_19294,N_19048,N_19051);
xor U19295 (N_19295,N_19166,N_18953);
xor U19296 (N_19296,N_19167,N_18880);
nor U19297 (N_19297,N_19126,N_19152);
nand U19298 (N_19298,N_19009,N_18886);
nor U19299 (N_19299,N_18920,N_18900);
and U19300 (N_19300,N_18958,N_19178);
and U19301 (N_19301,N_19027,N_19099);
nor U19302 (N_19302,N_19042,N_18987);
xnor U19303 (N_19303,N_19107,N_19198);
nand U19304 (N_19304,N_18999,N_19123);
or U19305 (N_19305,N_18945,N_18938);
nand U19306 (N_19306,N_19055,N_19102);
and U19307 (N_19307,N_19112,N_18817);
nor U19308 (N_19308,N_18968,N_19109);
nor U19309 (N_19309,N_19063,N_19156);
xor U19310 (N_19310,N_19019,N_19005);
or U19311 (N_19311,N_18967,N_18841);
xnor U19312 (N_19312,N_18929,N_18852);
nand U19313 (N_19313,N_18850,N_18990);
nor U19314 (N_19314,N_19127,N_19151);
and U19315 (N_19315,N_19088,N_19091);
and U19316 (N_19316,N_18991,N_18970);
nor U19317 (N_19317,N_18865,N_19182);
or U19318 (N_19318,N_19013,N_19081);
and U19319 (N_19319,N_18988,N_18823);
or U19320 (N_19320,N_19142,N_19070);
xor U19321 (N_19321,N_19192,N_18813);
or U19322 (N_19322,N_18913,N_19092);
nand U19323 (N_19323,N_18864,N_18936);
nor U19324 (N_19324,N_18960,N_18931);
nor U19325 (N_19325,N_19094,N_19012);
or U19326 (N_19326,N_18943,N_18885);
xor U19327 (N_19327,N_19056,N_19135);
nand U19328 (N_19328,N_18812,N_18868);
xor U19329 (N_19329,N_18923,N_19168);
xor U19330 (N_19330,N_19017,N_18907);
xnor U19331 (N_19331,N_18894,N_18903);
nor U19332 (N_19332,N_18808,N_18959);
and U19333 (N_19333,N_18914,N_18877);
nand U19334 (N_19334,N_19125,N_19150);
and U19335 (N_19335,N_18815,N_18835);
or U19336 (N_19336,N_19093,N_18853);
or U19337 (N_19337,N_18966,N_19060);
or U19338 (N_19338,N_19061,N_19179);
xor U19339 (N_19339,N_18950,N_19197);
and U19340 (N_19340,N_19183,N_19169);
and U19341 (N_19341,N_19101,N_19174);
nand U19342 (N_19342,N_19065,N_19193);
or U19343 (N_19343,N_19139,N_19097);
nand U19344 (N_19344,N_19158,N_19172);
nand U19345 (N_19345,N_19075,N_18917);
nor U19346 (N_19346,N_19196,N_19187);
xnor U19347 (N_19347,N_19136,N_19041);
or U19348 (N_19348,N_18993,N_18902);
and U19349 (N_19349,N_19138,N_18888);
nand U19350 (N_19350,N_18997,N_19057);
nand U19351 (N_19351,N_18974,N_18963);
xnor U19352 (N_19352,N_19083,N_18916);
and U19353 (N_19353,N_19148,N_19038);
nor U19354 (N_19354,N_18849,N_18807);
xor U19355 (N_19355,N_19054,N_18858);
nor U19356 (N_19356,N_18889,N_18825);
xor U19357 (N_19357,N_18946,N_19049);
nor U19358 (N_19358,N_18800,N_19145);
nand U19359 (N_19359,N_19082,N_18846);
nand U19360 (N_19360,N_18940,N_18879);
and U19361 (N_19361,N_19026,N_19020);
xnor U19362 (N_19362,N_18971,N_19176);
or U19363 (N_19363,N_18912,N_18922);
nor U19364 (N_19364,N_19114,N_18973);
and U19365 (N_19365,N_19037,N_18985);
or U19366 (N_19366,N_18949,N_18826);
nor U19367 (N_19367,N_18833,N_19173);
xor U19368 (N_19368,N_18954,N_19033);
or U19369 (N_19369,N_19137,N_18836);
or U19370 (N_19370,N_18924,N_19008);
nand U19371 (N_19371,N_19045,N_19068);
xor U19372 (N_19372,N_18882,N_18820);
and U19373 (N_19373,N_19064,N_18832);
nor U19374 (N_19374,N_19128,N_18978);
xor U19375 (N_19375,N_18911,N_19175);
nor U19376 (N_19376,N_19016,N_19015);
nor U19377 (N_19377,N_19116,N_18844);
or U19378 (N_19378,N_19162,N_19007);
nand U19379 (N_19379,N_18977,N_18964);
or U19380 (N_19380,N_18806,N_18933);
nor U19381 (N_19381,N_18925,N_18802);
and U19382 (N_19382,N_18956,N_18870);
and U19383 (N_19383,N_18874,N_19191);
or U19384 (N_19384,N_19072,N_19194);
and U19385 (N_19385,N_18906,N_19078);
and U19386 (N_19386,N_18871,N_18859);
or U19387 (N_19387,N_18854,N_18814);
nor U19388 (N_19388,N_19165,N_19034);
nor U19389 (N_19389,N_18982,N_19035);
and U19390 (N_19390,N_19071,N_19134);
nand U19391 (N_19391,N_18818,N_18898);
or U19392 (N_19392,N_19022,N_19098);
xor U19393 (N_19393,N_18928,N_18962);
and U19394 (N_19394,N_19079,N_19067);
or U19395 (N_19395,N_18951,N_18842);
or U19396 (N_19396,N_18803,N_18890);
nor U19397 (N_19397,N_18856,N_18961);
nand U19398 (N_19398,N_18994,N_19117);
or U19399 (N_19399,N_19133,N_19146);
or U19400 (N_19400,N_18846,N_18811);
xnor U19401 (N_19401,N_19014,N_18848);
nand U19402 (N_19402,N_19035,N_18877);
and U19403 (N_19403,N_18824,N_19153);
and U19404 (N_19404,N_18944,N_18903);
and U19405 (N_19405,N_18871,N_19198);
or U19406 (N_19406,N_19053,N_18901);
xnor U19407 (N_19407,N_18872,N_18871);
nand U19408 (N_19408,N_18898,N_19084);
and U19409 (N_19409,N_19029,N_19031);
xor U19410 (N_19410,N_18957,N_18944);
nor U19411 (N_19411,N_18965,N_19100);
or U19412 (N_19412,N_18839,N_19072);
nand U19413 (N_19413,N_19126,N_18973);
nor U19414 (N_19414,N_18991,N_19094);
and U19415 (N_19415,N_18871,N_18868);
nand U19416 (N_19416,N_19080,N_19017);
xor U19417 (N_19417,N_18991,N_19141);
or U19418 (N_19418,N_19134,N_18812);
nor U19419 (N_19419,N_18954,N_18818);
or U19420 (N_19420,N_19155,N_18929);
nor U19421 (N_19421,N_18852,N_19114);
or U19422 (N_19422,N_19107,N_19045);
nand U19423 (N_19423,N_18966,N_19185);
and U19424 (N_19424,N_18899,N_19001);
or U19425 (N_19425,N_18953,N_18948);
xnor U19426 (N_19426,N_19140,N_19057);
xor U19427 (N_19427,N_19158,N_18920);
xnor U19428 (N_19428,N_18887,N_18962);
xor U19429 (N_19429,N_19128,N_19031);
xor U19430 (N_19430,N_18804,N_18816);
or U19431 (N_19431,N_19102,N_19098);
and U19432 (N_19432,N_18892,N_19093);
nor U19433 (N_19433,N_18939,N_18977);
or U19434 (N_19434,N_18900,N_19029);
nor U19435 (N_19435,N_18948,N_19008);
nor U19436 (N_19436,N_19020,N_19107);
and U19437 (N_19437,N_18925,N_19096);
nor U19438 (N_19438,N_18807,N_18892);
nor U19439 (N_19439,N_19192,N_18806);
nand U19440 (N_19440,N_19038,N_19104);
and U19441 (N_19441,N_18808,N_18926);
and U19442 (N_19442,N_19136,N_18837);
nor U19443 (N_19443,N_18942,N_18936);
nor U19444 (N_19444,N_18901,N_19190);
or U19445 (N_19445,N_19132,N_19045);
or U19446 (N_19446,N_18996,N_19196);
and U19447 (N_19447,N_19050,N_19007);
xnor U19448 (N_19448,N_19143,N_19166);
or U19449 (N_19449,N_18883,N_19030);
and U19450 (N_19450,N_19174,N_18920);
or U19451 (N_19451,N_19054,N_19127);
nor U19452 (N_19452,N_18831,N_19133);
nor U19453 (N_19453,N_19176,N_19111);
or U19454 (N_19454,N_19129,N_19034);
or U19455 (N_19455,N_19072,N_18847);
nor U19456 (N_19456,N_18914,N_18803);
nand U19457 (N_19457,N_19163,N_19005);
nor U19458 (N_19458,N_18918,N_19037);
nand U19459 (N_19459,N_19160,N_18895);
nor U19460 (N_19460,N_19027,N_18912);
or U19461 (N_19461,N_18875,N_18819);
and U19462 (N_19462,N_19113,N_18881);
and U19463 (N_19463,N_19049,N_19140);
xor U19464 (N_19464,N_18976,N_18827);
and U19465 (N_19465,N_18819,N_19065);
xor U19466 (N_19466,N_19062,N_19113);
nor U19467 (N_19467,N_19106,N_19050);
or U19468 (N_19468,N_18850,N_19133);
xor U19469 (N_19469,N_19020,N_18893);
nand U19470 (N_19470,N_19188,N_18935);
xnor U19471 (N_19471,N_19022,N_18876);
nor U19472 (N_19472,N_18911,N_18870);
and U19473 (N_19473,N_19060,N_19068);
nand U19474 (N_19474,N_18928,N_19113);
nand U19475 (N_19475,N_19101,N_19156);
or U19476 (N_19476,N_18811,N_19040);
and U19477 (N_19477,N_18937,N_18968);
xor U19478 (N_19478,N_18851,N_19138);
nor U19479 (N_19479,N_18802,N_19024);
xor U19480 (N_19480,N_19033,N_19051);
and U19481 (N_19481,N_18873,N_19149);
xor U19482 (N_19482,N_18803,N_19037);
and U19483 (N_19483,N_18823,N_19063);
and U19484 (N_19484,N_19088,N_19137);
nor U19485 (N_19485,N_18968,N_18962);
or U19486 (N_19486,N_18812,N_19139);
nor U19487 (N_19487,N_18980,N_19020);
and U19488 (N_19488,N_19004,N_18955);
nor U19489 (N_19489,N_18829,N_18946);
nor U19490 (N_19490,N_18930,N_18984);
xnor U19491 (N_19491,N_18999,N_19050);
or U19492 (N_19492,N_19043,N_18835);
xor U19493 (N_19493,N_18863,N_18843);
and U19494 (N_19494,N_19034,N_19055);
nand U19495 (N_19495,N_19124,N_18858);
or U19496 (N_19496,N_18890,N_19099);
and U19497 (N_19497,N_19019,N_19191);
xnor U19498 (N_19498,N_18827,N_19189);
nor U19499 (N_19499,N_18960,N_19096);
nand U19500 (N_19500,N_18887,N_18860);
or U19501 (N_19501,N_18973,N_18891);
and U19502 (N_19502,N_18820,N_18841);
nand U19503 (N_19503,N_19075,N_19090);
and U19504 (N_19504,N_19157,N_18965);
nor U19505 (N_19505,N_19131,N_18874);
xnor U19506 (N_19506,N_19005,N_18899);
and U19507 (N_19507,N_19031,N_19182);
or U19508 (N_19508,N_19003,N_19131);
nand U19509 (N_19509,N_18878,N_18842);
and U19510 (N_19510,N_19082,N_19042);
or U19511 (N_19511,N_19136,N_18881);
or U19512 (N_19512,N_19099,N_19183);
and U19513 (N_19513,N_19002,N_19194);
xnor U19514 (N_19514,N_19139,N_18904);
xnor U19515 (N_19515,N_18812,N_18928);
and U19516 (N_19516,N_18952,N_19189);
nor U19517 (N_19517,N_18926,N_18968);
and U19518 (N_19518,N_18895,N_19188);
nor U19519 (N_19519,N_19089,N_18927);
xor U19520 (N_19520,N_19079,N_18880);
or U19521 (N_19521,N_18816,N_18940);
nor U19522 (N_19522,N_18985,N_18921);
nor U19523 (N_19523,N_18823,N_19153);
or U19524 (N_19524,N_19192,N_19037);
nor U19525 (N_19525,N_18835,N_18843);
nand U19526 (N_19526,N_19117,N_18968);
nand U19527 (N_19527,N_18962,N_18876);
nor U19528 (N_19528,N_19180,N_19183);
and U19529 (N_19529,N_19094,N_19130);
or U19530 (N_19530,N_18872,N_18934);
and U19531 (N_19531,N_18837,N_18994);
or U19532 (N_19532,N_19187,N_18847);
nand U19533 (N_19533,N_19126,N_19014);
nor U19534 (N_19534,N_19157,N_19183);
xnor U19535 (N_19535,N_18952,N_18928);
nor U19536 (N_19536,N_18976,N_18911);
or U19537 (N_19537,N_19123,N_19167);
and U19538 (N_19538,N_18827,N_18859);
xor U19539 (N_19539,N_19102,N_19010);
nand U19540 (N_19540,N_19019,N_18884);
nor U19541 (N_19541,N_19072,N_18981);
nand U19542 (N_19542,N_18913,N_19194);
or U19543 (N_19543,N_18908,N_18909);
xnor U19544 (N_19544,N_18888,N_18964);
nand U19545 (N_19545,N_18962,N_19023);
nor U19546 (N_19546,N_18933,N_19167);
and U19547 (N_19547,N_19103,N_19073);
nor U19548 (N_19548,N_18970,N_18957);
or U19549 (N_19549,N_19024,N_19075);
and U19550 (N_19550,N_18897,N_18823);
xnor U19551 (N_19551,N_18831,N_18915);
nor U19552 (N_19552,N_19083,N_19004);
xnor U19553 (N_19553,N_18837,N_19159);
nand U19554 (N_19554,N_19105,N_19096);
and U19555 (N_19555,N_18829,N_18931);
or U19556 (N_19556,N_19058,N_18947);
or U19557 (N_19557,N_18871,N_19144);
or U19558 (N_19558,N_19004,N_19125);
xnor U19559 (N_19559,N_18923,N_18871);
and U19560 (N_19560,N_19112,N_18953);
or U19561 (N_19561,N_18978,N_18971);
nor U19562 (N_19562,N_19094,N_19038);
and U19563 (N_19563,N_18848,N_18989);
or U19564 (N_19564,N_18962,N_19082);
or U19565 (N_19565,N_19022,N_18854);
and U19566 (N_19566,N_19034,N_18886);
and U19567 (N_19567,N_18871,N_19136);
and U19568 (N_19568,N_18854,N_19128);
nor U19569 (N_19569,N_18939,N_19152);
xor U19570 (N_19570,N_19109,N_19142);
nor U19571 (N_19571,N_19192,N_19111);
and U19572 (N_19572,N_18971,N_19171);
or U19573 (N_19573,N_19196,N_18998);
xnor U19574 (N_19574,N_19104,N_19101);
xnor U19575 (N_19575,N_19171,N_18917);
nor U19576 (N_19576,N_18846,N_19043);
xor U19577 (N_19577,N_19026,N_19037);
or U19578 (N_19578,N_19083,N_18880);
xnor U19579 (N_19579,N_19159,N_19155);
xor U19580 (N_19580,N_19007,N_19049);
and U19581 (N_19581,N_19133,N_18906);
xnor U19582 (N_19582,N_19031,N_18994);
xnor U19583 (N_19583,N_19052,N_18848);
or U19584 (N_19584,N_18835,N_18987);
or U19585 (N_19585,N_18944,N_19165);
nand U19586 (N_19586,N_18881,N_19004);
nor U19587 (N_19587,N_18949,N_18850);
and U19588 (N_19588,N_18972,N_19066);
or U19589 (N_19589,N_19022,N_19133);
xor U19590 (N_19590,N_18977,N_18944);
or U19591 (N_19591,N_18881,N_18883);
nand U19592 (N_19592,N_18891,N_18945);
and U19593 (N_19593,N_19198,N_19024);
nor U19594 (N_19594,N_19196,N_18852);
nand U19595 (N_19595,N_19033,N_19021);
and U19596 (N_19596,N_19076,N_18804);
nand U19597 (N_19597,N_18937,N_19169);
nor U19598 (N_19598,N_19043,N_18830);
or U19599 (N_19599,N_19082,N_18929);
nand U19600 (N_19600,N_19311,N_19474);
nor U19601 (N_19601,N_19280,N_19565);
nand U19602 (N_19602,N_19589,N_19300);
or U19603 (N_19603,N_19504,N_19418);
xor U19604 (N_19604,N_19314,N_19431);
or U19605 (N_19605,N_19224,N_19371);
nand U19606 (N_19606,N_19265,N_19454);
and U19607 (N_19607,N_19271,N_19452);
or U19608 (N_19608,N_19357,N_19342);
and U19609 (N_19609,N_19460,N_19451);
or U19610 (N_19610,N_19248,N_19385);
nand U19611 (N_19611,N_19550,N_19554);
nand U19612 (N_19612,N_19487,N_19365);
or U19613 (N_19613,N_19345,N_19448);
nor U19614 (N_19614,N_19313,N_19576);
and U19615 (N_19615,N_19330,N_19476);
xnor U19616 (N_19616,N_19536,N_19564);
and U19617 (N_19617,N_19307,N_19363);
xor U19618 (N_19618,N_19478,N_19470);
nor U19619 (N_19619,N_19329,N_19347);
and U19620 (N_19620,N_19333,N_19226);
and U19621 (N_19621,N_19569,N_19406);
nand U19622 (N_19622,N_19533,N_19320);
or U19623 (N_19623,N_19309,N_19350);
or U19624 (N_19624,N_19362,N_19259);
nor U19625 (N_19625,N_19257,N_19272);
nor U19626 (N_19626,N_19223,N_19207);
xor U19627 (N_19627,N_19425,N_19377);
xnor U19628 (N_19628,N_19530,N_19441);
xor U19629 (N_19629,N_19518,N_19368);
nand U19630 (N_19630,N_19408,N_19279);
nor U19631 (N_19631,N_19402,N_19570);
nand U19632 (N_19632,N_19228,N_19484);
and U19633 (N_19633,N_19281,N_19493);
or U19634 (N_19634,N_19278,N_19239);
nand U19635 (N_19635,N_19323,N_19409);
and U19636 (N_19636,N_19293,N_19415);
nor U19637 (N_19637,N_19359,N_19205);
nor U19638 (N_19638,N_19566,N_19219);
nor U19639 (N_19639,N_19541,N_19497);
nand U19640 (N_19640,N_19496,N_19430);
nor U19641 (N_19641,N_19232,N_19374);
nor U19642 (N_19642,N_19482,N_19260);
or U19643 (N_19643,N_19503,N_19417);
nor U19644 (N_19644,N_19584,N_19549);
nand U19645 (N_19645,N_19546,N_19521);
nor U19646 (N_19646,N_19514,N_19412);
xnor U19647 (N_19647,N_19535,N_19354);
xor U19648 (N_19648,N_19398,N_19594);
and U19649 (N_19649,N_19339,N_19305);
and U19650 (N_19650,N_19435,N_19466);
xor U19651 (N_19651,N_19446,N_19407);
nor U19652 (N_19652,N_19388,N_19560);
nand U19653 (N_19653,N_19526,N_19575);
nor U19654 (N_19654,N_19577,N_19447);
nand U19655 (N_19655,N_19432,N_19225);
and U19656 (N_19656,N_19250,N_19439);
and U19657 (N_19657,N_19264,N_19251);
or U19658 (N_19658,N_19203,N_19332);
and U19659 (N_19659,N_19310,N_19218);
and U19660 (N_19660,N_19472,N_19277);
nand U19661 (N_19661,N_19210,N_19324);
and U19662 (N_19662,N_19587,N_19539);
and U19663 (N_19663,N_19591,N_19289);
or U19664 (N_19664,N_19491,N_19302);
or U19665 (N_19665,N_19258,N_19369);
and U19666 (N_19666,N_19298,N_19282);
or U19667 (N_19667,N_19519,N_19284);
or U19668 (N_19668,N_19410,N_19352);
nor U19669 (N_19669,N_19364,N_19241);
and U19670 (N_19670,N_19586,N_19580);
nor U19671 (N_19671,N_19489,N_19465);
nand U19672 (N_19672,N_19548,N_19304);
nand U19673 (N_19673,N_19348,N_19341);
and U19674 (N_19674,N_19469,N_19552);
or U19675 (N_19675,N_19276,N_19331);
and U19676 (N_19676,N_19413,N_19319);
and U19677 (N_19677,N_19442,N_19467);
xnor U19678 (N_19678,N_19375,N_19567);
and U19679 (N_19679,N_19574,N_19557);
xnor U19680 (N_19680,N_19438,N_19367);
and U19681 (N_19681,N_19488,N_19527);
nand U19682 (N_19682,N_19543,N_19243);
xnor U19683 (N_19683,N_19273,N_19502);
or U19684 (N_19684,N_19286,N_19372);
or U19685 (N_19685,N_19501,N_19202);
xor U19686 (N_19686,N_19249,N_19595);
nor U19687 (N_19687,N_19340,N_19414);
or U19688 (N_19688,N_19401,N_19433);
xor U19689 (N_19689,N_19295,N_19321);
nand U19690 (N_19690,N_19582,N_19532);
or U19691 (N_19691,N_19204,N_19326);
or U19692 (N_19692,N_19351,N_19598);
nor U19693 (N_19693,N_19394,N_19421);
nor U19694 (N_19694,N_19547,N_19434);
or U19695 (N_19695,N_19424,N_19209);
or U19696 (N_19696,N_19395,N_19509);
nor U19697 (N_19697,N_19562,N_19328);
nor U19698 (N_19698,N_19392,N_19393);
and U19699 (N_19699,N_19573,N_19361);
nor U19700 (N_19700,N_19349,N_19338);
xnor U19701 (N_19701,N_19471,N_19390);
and U19702 (N_19702,N_19422,N_19237);
and U19703 (N_19703,N_19429,N_19444);
nor U19704 (N_19704,N_19544,N_19212);
nand U19705 (N_19705,N_19563,N_19531);
nand U19706 (N_19706,N_19515,N_19525);
xnor U19707 (N_19707,N_19461,N_19379);
nor U19708 (N_19708,N_19353,N_19599);
or U19709 (N_19709,N_19381,N_19268);
nor U19710 (N_19710,N_19510,N_19294);
and U19711 (N_19711,N_19366,N_19597);
xnor U19712 (N_19712,N_19383,N_19308);
or U19713 (N_19713,N_19522,N_19581);
and U19714 (N_19714,N_19490,N_19358);
or U19715 (N_19715,N_19200,N_19235);
or U19716 (N_19716,N_19245,N_19222);
or U19717 (N_19717,N_19336,N_19495);
or U19718 (N_19718,N_19585,N_19318);
nor U19719 (N_19719,N_19356,N_19456);
xor U19720 (N_19720,N_19337,N_19578);
xor U19721 (N_19721,N_19457,N_19556);
nand U19722 (N_19722,N_19481,N_19261);
nor U19723 (N_19723,N_19238,N_19391);
nor U19724 (N_19724,N_19483,N_19303);
or U19725 (N_19725,N_19485,N_19206);
and U19726 (N_19726,N_19215,N_19559);
nand U19727 (N_19727,N_19463,N_19274);
nand U19728 (N_19728,N_19427,N_19397);
nand U19729 (N_19729,N_19380,N_19299);
xnor U19730 (N_19730,N_19384,N_19396);
nand U19731 (N_19731,N_19568,N_19520);
nand U19732 (N_19732,N_19312,N_19459);
and U19733 (N_19733,N_19233,N_19437);
xor U19734 (N_19734,N_19419,N_19505);
and U19735 (N_19735,N_19344,N_19517);
nor U19736 (N_19736,N_19376,N_19378);
and U19737 (N_19737,N_19211,N_19247);
nand U19738 (N_19738,N_19229,N_19382);
xor U19739 (N_19739,N_19267,N_19227);
and U19740 (N_19740,N_19492,N_19389);
xnor U19741 (N_19741,N_19360,N_19499);
or U19742 (N_19742,N_19240,N_19387);
nand U19743 (N_19743,N_19480,N_19426);
nor U19744 (N_19744,N_19334,N_19473);
nand U19745 (N_19745,N_19399,N_19416);
nand U19746 (N_19746,N_19553,N_19445);
nand U19747 (N_19747,N_19252,N_19475);
and U19748 (N_19748,N_19523,N_19327);
nand U19749 (N_19749,N_19287,N_19275);
xnor U19750 (N_19750,N_19440,N_19283);
nand U19751 (N_19751,N_19593,N_19458);
or U19752 (N_19752,N_19464,N_19325);
nand U19753 (N_19753,N_19449,N_19558);
and U19754 (N_19754,N_19500,N_19524);
nor U19755 (N_19755,N_19253,N_19290);
and U19756 (N_19756,N_19404,N_19511);
and U19757 (N_19757,N_19234,N_19400);
xor U19758 (N_19758,N_19486,N_19528);
and U19759 (N_19759,N_19285,N_19588);
and U19760 (N_19760,N_19443,N_19590);
nor U19761 (N_19761,N_19370,N_19512);
or U19762 (N_19762,N_19579,N_19571);
nand U19763 (N_19763,N_19583,N_19317);
and U19764 (N_19764,N_19255,N_19405);
nor U19765 (N_19765,N_19538,N_19201);
nand U19766 (N_19766,N_19297,N_19296);
and U19767 (N_19767,N_19420,N_19498);
and U19768 (N_19768,N_19316,N_19572);
and U19769 (N_19769,N_19423,N_19508);
nand U19770 (N_19770,N_19306,N_19221);
and U19771 (N_19771,N_19428,N_19355);
xnor U19772 (N_19772,N_19230,N_19322);
and U19773 (N_19773,N_19477,N_19213);
nand U19774 (N_19774,N_19254,N_19537);
and U19775 (N_19775,N_19291,N_19270);
nand U19776 (N_19776,N_19513,N_19494);
or U19777 (N_19777,N_19373,N_19506);
or U19778 (N_19778,N_19214,N_19545);
and U19779 (N_19779,N_19269,N_19220);
nand U19780 (N_19780,N_19507,N_19217);
nand U19781 (N_19781,N_19561,N_19242);
nand U19782 (N_19782,N_19479,N_19542);
xnor U19783 (N_19783,N_19534,N_19386);
and U19784 (N_19784,N_19244,N_19343);
xnor U19785 (N_19785,N_19246,N_19301);
xor U19786 (N_19786,N_19468,N_19236);
nand U19787 (N_19787,N_19263,N_19266);
or U19788 (N_19788,N_19462,N_19436);
xnor U19789 (N_19789,N_19411,N_19455);
xor U19790 (N_19790,N_19555,N_19450);
xnor U19791 (N_19791,N_19529,N_19231);
nor U19792 (N_19792,N_19288,N_19208);
or U19793 (N_19793,N_19346,N_19540);
and U19794 (N_19794,N_19216,N_19596);
nand U19795 (N_19795,N_19551,N_19292);
xor U19796 (N_19796,N_19335,N_19453);
xor U19797 (N_19797,N_19592,N_19315);
and U19798 (N_19798,N_19403,N_19516);
nor U19799 (N_19799,N_19256,N_19262);
nor U19800 (N_19800,N_19480,N_19515);
nand U19801 (N_19801,N_19429,N_19517);
nor U19802 (N_19802,N_19511,N_19307);
nand U19803 (N_19803,N_19466,N_19542);
nand U19804 (N_19804,N_19219,N_19581);
nand U19805 (N_19805,N_19203,N_19321);
xor U19806 (N_19806,N_19514,N_19376);
xor U19807 (N_19807,N_19278,N_19549);
nand U19808 (N_19808,N_19338,N_19362);
and U19809 (N_19809,N_19266,N_19234);
nor U19810 (N_19810,N_19211,N_19388);
and U19811 (N_19811,N_19271,N_19357);
and U19812 (N_19812,N_19491,N_19349);
xor U19813 (N_19813,N_19446,N_19577);
nand U19814 (N_19814,N_19288,N_19559);
nor U19815 (N_19815,N_19330,N_19234);
or U19816 (N_19816,N_19473,N_19536);
and U19817 (N_19817,N_19323,N_19421);
nand U19818 (N_19818,N_19369,N_19585);
xnor U19819 (N_19819,N_19425,N_19547);
and U19820 (N_19820,N_19290,N_19476);
and U19821 (N_19821,N_19453,N_19226);
nand U19822 (N_19822,N_19221,N_19232);
nor U19823 (N_19823,N_19206,N_19461);
or U19824 (N_19824,N_19576,N_19529);
and U19825 (N_19825,N_19282,N_19477);
nand U19826 (N_19826,N_19214,N_19573);
nand U19827 (N_19827,N_19229,N_19575);
xor U19828 (N_19828,N_19516,N_19278);
or U19829 (N_19829,N_19417,N_19541);
and U19830 (N_19830,N_19230,N_19487);
nor U19831 (N_19831,N_19529,N_19515);
xor U19832 (N_19832,N_19353,N_19290);
xnor U19833 (N_19833,N_19297,N_19420);
nor U19834 (N_19834,N_19484,N_19433);
and U19835 (N_19835,N_19475,N_19499);
xnor U19836 (N_19836,N_19284,N_19527);
or U19837 (N_19837,N_19540,N_19454);
nor U19838 (N_19838,N_19444,N_19257);
nor U19839 (N_19839,N_19599,N_19428);
nor U19840 (N_19840,N_19466,N_19256);
or U19841 (N_19841,N_19524,N_19291);
xnor U19842 (N_19842,N_19412,N_19512);
or U19843 (N_19843,N_19461,N_19251);
nand U19844 (N_19844,N_19396,N_19480);
or U19845 (N_19845,N_19530,N_19527);
xnor U19846 (N_19846,N_19351,N_19566);
xor U19847 (N_19847,N_19582,N_19430);
and U19848 (N_19848,N_19348,N_19362);
or U19849 (N_19849,N_19457,N_19340);
xnor U19850 (N_19850,N_19504,N_19330);
or U19851 (N_19851,N_19512,N_19545);
and U19852 (N_19852,N_19200,N_19538);
nor U19853 (N_19853,N_19371,N_19597);
nor U19854 (N_19854,N_19433,N_19313);
xnor U19855 (N_19855,N_19419,N_19511);
nand U19856 (N_19856,N_19472,N_19447);
nor U19857 (N_19857,N_19568,N_19328);
and U19858 (N_19858,N_19572,N_19268);
xnor U19859 (N_19859,N_19387,N_19210);
xor U19860 (N_19860,N_19212,N_19569);
nor U19861 (N_19861,N_19306,N_19421);
or U19862 (N_19862,N_19372,N_19209);
xor U19863 (N_19863,N_19416,N_19446);
and U19864 (N_19864,N_19265,N_19236);
and U19865 (N_19865,N_19475,N_19532);
or U19866 (N_19866,N_19541,N_19342);
or U19867 (N_19867,N_19304,N_19374);
nand U19868 (N_19868,N_19410,N_19388);
xnor U19869 (N_19869,N_19415,N_19489);
nand U19870 (N_19870,N_19386,N_19226);
or U19871 (N_19871,N_19486,N_19506);
and U19872 (N_19872,N_19306,N_19255);
xor U19873 (N_19873,N_19331,N_19564);
or U19874 (N_19874,N_19356,N_19550);
xnor U19875 (N_19875,N_19327,N_19479);
nor U19876 (N_19876,N_19407,N_19359);
nand U19877 (N_19877,N_19290,N_19543);
nand U19878 (N_19878,N_19331,N_19260);
and U19879 (N_19879,N_19417,N_19513);
xor U19880 (N_19880,N_19265,N_19201);
and U19881 (N_19881,N_19559,N_19404);
or U19882 (N_19882,N_19439,N_19321);
and U19883 (N_19883,N_19254,N_19483);
nor U19884 (N_19884,N_19530,N_19553);
or U19885 (N_19885,N_19445,N_19202);
nand U19886 (N_19886,N_19314,N_19445);
or U19887 (N_19887,N_19242,N_19228);
or U19888 (N_19888,N_19229,N_19433);
or U19889 (N_19889,N_19364,N_19557);
or U19890 (N_19890,N_19240,N_19531);
xor U19891 (N_19891,N_19564,N_19516);
or U19892 (N_19892,N_19383,N_19578);
xor U19893 (N_19893,N_19393,N_19210);
nor U19894 (N_19894,N_19473,N_19386);
xnor U19895 (N_19895,N_19537,N_19279);
or U19896 (N_19896,N_19421,N_19324);
nand U19897 (N_19897,N_19586,N_19440);
xor U19898 (N_19898,N_19474,N_19445);
xor U19899 (N_19899,N_19396,N_19234);
nor U19900 (N_19900,N_19235,N_19548);
nand U19901 (N_19901,N_19476,N_19228);
xor U19902 (N_19902,N_19274,N_19489);
xnor U19903 (N_19903,N_19319,N_19213);
xnor U19904 (N_19904,N_19475,N_19349);
and U19905 (N_19905,N_19238,N_19439);
and U19906 (N_19906,N_19549,N_19528);
nand U19907 (N_19907,N_19540,N_19292);
nor U19908 (N_19908,N_19290,N_19330);
xor U19909 (N_19909,N_19446,N_19202);
or U19910 (N_19910,N_19562,N_19369);
and U19911 (N_19911,N_19385,N_19230);
or U19912 (N_19912,N_19286,N_19298);
xor U19913 (N_19913,N_19466,N_19348);
or U19914 (N_19914,N_19526,N_19450);
and U19915 (N_19915,N_19316,N_19513);
nor U19916 (N_19916,N_19208,N_19396);
nor U19917 (N_19917,N_19428,N_19375);
nor U19918 (N_19918,N_19383,N_19246);
nand U19919 (N_19919,N_19223,N_19337);
or U19920 (N_19920,N_19282,N_19520);
and U19921 (N_19921,N_19390,N_19286);
nor U19922 (N_19922,N_19252,N_19341);
and U19923 (N_19923,N_19310,N_19278);
or U19924 (N_19924,N_19524,N_19280);
or U19925 (N_19925,N_19535,N_19279);
and U19926 (N_19926,N_19337,N_19284);
xor U19927 (N_19927,N_19441,N_19576);
nor U19928 (N_19928,N_19343,N_19485);
xor U19929 (N_19929,N_19267,N_19560);
nand U19930 (N_19930,N_19435,N_19234);
nand U19931 (N_19931,N_19532,N_19229);
and U19932 (N_19932,N_19218,N_19279);
nand U19933 (N_19933,N_19561,N_19406);
nand U19934 (N_19934,N_19320,N_19313);
or U19935 (N_19935,N_19212,N_19344);
nor U19936 (N_19936,N_19520,N_19342);
nor U19937 (N_19937,N_19431,N_19560);
or U19938 (N_19938,N_19492,N_19499);
nand U19939 (N_19939,N_19501,N_19552);
and U19940 (N_19940,N_19386,N_19410);
or U19941 (N_19941,N_19514,N_19426);
nand U19942 (N_19942,N_19391,N_19396);
and U19943 (N_19943,N_19438,N_19370);
and U19944 (N_19944,N_19255,N_19440);
and U19945 (N_19945,N_19393,N_19399);
nand U19946 (N_19946,N_19230,N_19266);
nand U19947 (N_19947,N_19358,N_19210);
nor U19948 (N_19948,N_19518,N_19267);
nor U19949 (N_19949,N_19261,N_19292);
xnor U19950 (N_19950,N_19353,N_19374);
xnor U19951 (N_19951,N_19243,N_19501);
nor U19952 (N_19952,N_19399,N_19583);
nand U19953 (N_19953,N_19222,N_19581);
nor U19954 (N_19954,N_19424,N_19355);
xor U19955 (N_19955,N_19349,N_19272);
nand U19956 (N_19956,N_19530,N_19503);
nand U19957 (N_19957,N_19386,N_19577);
nor U19958 (N_19958,N_19289,N_19393);
xnor U19959 (N_19959,N_19573,N_19380);
and U19960 (N_19960,N_19241,N_19431);
and U19961 (N_19961,N_19456,N_19446);
nand U19962 (N_19962,N_19368,N_19418);
and U19963 (N_19963,N_19488,N_19440);
xnor U19964 (N_19964,N_19549,N_19223);
and U19965 (N_19965,N_19384,N_19339);
nand U19966 (N_19966,N_19340,N_19259);
nand U19967 (N_19967,N_19517,N_19558);
nand U19968 (N_19968,N_19598,N_19272);
or U19969 (N_19969,N_19326,N_19534);
or U19970 (N_19970,N_19470,N_19258);
nor U19971 (N_19971,N_19311,N_19552);
nand U19972 (N_19972,N_19437,N_19432);
xnor U19973 (N_19973,N_19550,N_19330);
and U19974 (N_19974,N_19269,N_19485);
and U19975 (N_19975,N_19386,N_19466);
nor U19976 (N_19976,N_19519,N_19310);
or U19977 (N_19977,N_19230,N_19299);
and U19978 (N_19978,N_19567,N_19443);
or U19979 (N_19979,N_19560,N_19386);
or U19980 (N_19980,N_19286,N_19432);
nand U19981 (N_19981,N_19376,N_19419);
or U19982 (N_19982,N_19482,N_19506);
nor U19983 (N_19983,N_19319,N_19332);
and U19984 (N_19984,N_19464,N_19367);
nand U19985 (N_19985,N_19303,N_19560);
nor U19986 (N_19986,N_19319,N_19381);
nand U19987 (N_19987,N_19510,N_19267);
nand U19988 (N_19988,N_19212,N_19227);
or U19989 (N_19989,N_19531,N_19305);
nor U19990 (N_19990,N_19269,N_19379);
nor U19991 (N_19991,N_19288,N_19567);
nor U19992 (N_19992,N_19352,N_19560);
and U19993 (N_19993,N_19226,N_19306);
nor U19994 (N_19994,N_19505,N_19595);
xnor U19995 (N_19995,N_19440,N_19384);
and U19996 (N_19996,N_19417,N_19221);
nand U19997 (N_19997,N_19503,N_19591);
and U19998 (N_19998,N_19202,N_19490);
nand U19999 (N_19999,N_19593,N_19273);
and UO_0 (O_0,N_19882,N_19845);
and UO_1 (O_1,N_19772,N_19911);
or UO_2 (O_2,N_19895,N_19636);
and UO_3 (O_3,N_19902,N_19690);
xnor UO_4 (O_4,N_19719,N_19939);
nor UO_5 (O_5,N_19989,N_19816);
nand UO_6 (O_6,N_19774,N_19763);
nand UO_7 (O_7,N_19940,N_19853);
nand UO_8 (O_8,N_19838,N_19963);
xnor UO_9 (O_9,N_19986,N_19937);
or UO_10 (O_10,N_19642,N_19696);
and UO_11 (O_11,N_19996,N_19835);
nand UO_12 (O_12,N_19914,N_19977);
or UO_13 (O_13,N_19625,N_19701);
or UO_14 (O_14,N_19910,N_19828);
or UO_15 (O_15,N_19757,N_19775);
or UO_16 (O_16,N_19703,N_19707);
and UO_17 (O_17,N_19614,N_19605);
xor UO_18 (O_18,N_19741,N_19734);
nand UO_19 (O_19,N_19821,N_19639);
or UO_20 (O_20,N_19618,N_19724);
and UO_21 (O_21,N_19922,N_19941);
xnor UO_22 (O_22,N_19736,N_19817);
nand UO_23 (O_23,N_19744,N_19990);
xor UO_24 (O_24,N_19607,N_19924);
and UO_25 (O_25,N_19799,N_19795);
nand UO_26 (O_26,N_19779,N_19766);
nor UO_27 (O_27,N_19824,N_19920);
or UO_28 (O_28,N_19800,N_19968);
nand UO_29 (O_29,N_19967,N_19749);
or UO_30 (O_30,N_19826,N_19848);
and UO_31 (O_31,N_19679,N_19930);
and UO_32 (O_32,N_19641,N_19851);
nor UO_33 (O_33,N_19698,N_19776);
nand UO_34 (O_34,N_19601,N_19712);
nor UO_35 (O_35,N_19889,N_19718);
xnor UO_36 (O_36,N_19648,N_19926);
xor UO_37 (O_37,N_19833,N_19946);
nand UO_38 (O_38,N_19938,N_19808);
nand UO_39 (O_39,N_19862,N_19794);
or UO_40 (O_40,N_19945,N_19888);
xnor UO_41 (O_41,N_19691,N_19656);
and UO_42 (O_42,N_19747,N_19982);
xor UO_43 (O_43,N_19704,N_19907);
or UO_44 (O_44,N_19886,N_19723);
xnor UO_45 (O_45,N_19847,N_19952);
nand UO_46 (O_46,N_19603,N_19832);
xor UO_47 (O_47,N_19602,N_19675);
xor UO_48 (O_48,N_19767,N_19745);
xnor UO_49 (O_49,N_19658,N_19975);
xnor UO_50 (O_50,N_19830,N_19765);
and UO_51 (O_51,N_19849,N_19604);
nand UO_52 (O_52,N_19633,N_19773);
xnor UO_53 (O_53,N_19970,N_19836);
nor UO_54 (O_54,N_19873,N_19993);
nand UO_55 (O_55,N_19667,N_19842);
nand UO_56 (O_56,N_19740,N_19655);
nor UO_57 (O_57,N_19730,N_19610);
xnor UO_58 (O_58,N_19643,N_19927);
nand UO_59 (O_59,N_19887,N_19791);
and UO_60 (O_60,N_19709,N_19634);
or UO_61 (O_61,N_19657,N_19620);
xor UO_62 (O_62,N_19969,N_19874);
and UO_63 (O_63,N_19864,N_19872);
or UO_64 (O_64,N_19735,N_19615);
and UO_65 (O_65,N_19796,N_19829);
xor UO_66 (O_66,N_19819,N_19743);
or UO_67 (O_67,N_19805,N_19646);
and UO_68 (O_68,N_19664,N_19960);
and UO_69 (O_69,N_19725,N_19687);
or UO_70 (O_70,N_19798,N_19890);
nand UO_71 (O_71,N_19733,N_19622);
xor UO_72 (O_72,N_19613,N_19962);
nand UO_73 (O_73,N_19943,N_19632);
or UO_74 (O_74,N_19992,N_19869);
or UO_75 (O_75,N_19801,N_19844);
xnor UO_76 (O_76,N_19971,N_19978);
nor UO_77 (O_77,N_19681,N_19893);
nor UO_78 (O_78,N_19955,N_19715);
nor UO_79 (O_79,N_19668,N_19822);
and UO_80 (O_80,N_19860,N_19731);
xor UO_81 (O_81,N_19883,N_19891);
and UO_82 (O_82,N_19637,N_19769);
nor UO_83 (O_83,N_19640,N_19998);
nor UO_84 (O_84,N_19793,N_19854);
nor UO_85 (O_85,N_19789,N_19997);
nor UO_86 (O_86,N_19953,N_19617);
nor UO_87 (O_87,N_19980,N_19797);
and UO_88 (O_88,N_19818,N_19780);
xor UO_89 (O_89,N_19739,N_19981);
or UO_90 (O_90,N_19635,N_19760);
nand UO_91 (O_91,N_19964,N_19693);
nor UO_92 (O_92,N_19954,N_19630);
or UO_93 (O_93,N_19683,N_19959);
nand UO_94 (O_94,N_19688,N_19958);
nor UO_95 (O_95,N_19965,N_19647);
and UO_96 (O_96,N_19689,N_19699);
or UO_97 (O_97,N_19863,N_19752);
nand UO_98 (O_98,N_19810,N_19686);
nor UO_99 (O_99,N_19843,N_19881);
and UO_100 (O_100,N_19645,N_19777);
xor UO_101 (O_101,N_19803,N_19961);
nand UO_102 (O_102,N_19976,N_19995);
nor UO_103 (O_103,N_19714,N_19729);
nand UO_104 (O_104,N_19823,N_19758);
and UO_105 (O_105,N_19612,N_19624);
or UO_106 (O_106,N_19680,N_19901);
xor UO_107 (O_107,N_19852,N_19855);
nand UO_108 (O_108,N_19820,N_19792);
nand UO_109 (O_109,N_19831,N_19606);
and UO_110 (O_110,N_19616,N_19721);
and UO_111 (O_111,N_19933,N_19700);
nor UO_112 (O_112,N_19942,N_19827);
or UO_113 (O_113,N_19627,N_19850);
or UO_114 (O_114,N_19650,N_19754);
or UO_115 (O_115,N_19732,N_19770);
and UO_116 (O_116,N_19786,N_19979);
or UO_117 (O_117,N_19841,N_19629);
or UO_118 (O_118,N_19807,N_19812);
nand UO_119 (O_119,N_19726,N_19814);
nor UO_120 (O_120,N_19949,N_19751);
nand UO_121 (O_121,N_19677,N_19894);
nor UO_122 (O_122,N_19611,N_19985);
or UO_123 (O_123,N_19662,N_19972);
nand UO_124 (O_124,N_19935,N_19755);
or UO_125 (O_125,N_19856,N_19802);
or UO_126 (O_126,N_19759,N_19896);
xor UO_127 (O_127,N_19884,N_19875);
nand UO_128 (O_128,N_19900,N_19925);
nor UO_129 (O_129,N_19957,N_19837);
or UO_130 (O_130,N_19878,N_19892);
or UO_131 (O_131,N_19934,N_19778);
nand UO_132 (O_132,N_19950,N_19834);
or UO_133 (O_133,N_19705,N_19917);
nor UO_134 (O_134,N_19684,N_19840);
nor UO_135 (O_135,N_19999,N_19905);
xnor UO_136 (O_136,N_19644,N_19694);
nand UO_137 (O_137,N_19988,N_19931);
or UO_138 (O_138,N_19669,N_19682);
or UO_139 (O_139,N_19991,N_19638);
and UO_140 (O_140,N_19654,N_19784);
nand UO_141 (O_141,N_19720,N_19738);
nor UO_142 (O_142,N_19947,N_19876);
xnor UO_143 (O_143,N_19932,N_19727);
xnor UO_144 (O_144,N_19813,N_19708);
and UO_145 (O_145,N_19659,N_19706);
xor UO_146 (O_146,N_19748,N_19631);
or UO_147 (O_147,N_19717,N_19861);
nand UO_148 (O_148,N_19877,N_19804);
or UO_149 (O_149,N_19600,N_19742);
nand UO_150 (O_150,N_19762,N_19919);
or UO_151 (O_151,N_19787,N_19913);
xor UO_152 (O_152,N_19653,N_19809);
or UO_153 (O_153,N_19663,N_19661);
and UO_154 (O_154,N_19753,N_19858);
nor UO_155 (O_155,N_19673,N_19923);
xnor UO_156 (O_156,N_19966,N_19652);
and UO_157 (O_157,N_19728,N_19660);
and UO_158 (O_158,N_19761,N_19626);
nor UO_159 (O_159,N_19665,N_19771);
xnor UO_160 (O_160,N_19974,N_19839);
nand UO_161 (O_161,N_19783,N_19870);
nand UO_162 (O_162,N_19904,N_19929);
nand UO_163 (O_163,N_19948,N_19951);
xnor UO_164 (O_164,N_19912,N_19746);
nor UO_165 (O_165,N_19750,N_19666);
or UO_166 (O_166,N_19782,N_19908);
nand UO_167 (O_167,N_19764,N_19983);
nor UO_168 (O_168,N_19678,N_19722);
xnor UO_169 (O_169,N_19649,N_19806);
nor UO_170 (O_170,N_19713,N_19885);
nand UO_171 (O_171,N_19903,N_19936);
nand UO_172 (O_172,N_19692,N_19623);
nand UO_173 (O_173,N_19899,N_19711);
nand UO_174 (O_174,N_19871,N_19898);
xor UO_175 (O_175,N_19768,N_19619);
xnor UO_176 (O_176,N_19609,N_19716);
or UO_177 (O_177,N_19859,N_19790);
nor UO_178 (O_178,N_19811,N_19984);
xor UO_179 (O_179,N_19921,N_19973);
or UO_180 (O_180,N_19756,N_19628);
nor UO_181 (O_181,N_19987,N_19918);
or UO_182 (O_182,N_19670,N_19788);
xor UO_183 (O_183,N_19857,N_19815);
nor UO_184 (O_184,N_19956,N_19915);
and UO_185 (O_185,N_19621,N_19785);
nor UO_186 (O_186,N_19737,N_19651);
nand UO_187 (O_187,N_19676,N_19781);
nand UO_188 (O_188,N_19671,N_19880);
nor UO_189 (O_189,N_19825,N_19674);
nand UO_190 (O_190,N_19866,N_19702);
xor UO_191 (O_191,N_19879,N_19695);
and UO_192 (O_192,N_19897,N_19685);
nor UO_193 (O_193,N_19865,N_19916);
nand UO_194 (O_194,N_19906,N_19710);
xnor UO_195 (O_195,N_19867,N_19868);
nor UO_196 (O_196,N_19909,N_19697);
or UO_197 (O_197,N_19944,N_19928);
or UO_198 (O_198,N_19994,N_19672);
and UO_199 (O_199,N_19846,N_19608);
nor UO_200 (O_200,N_19982,N_19618);
or UO_201 (O_201,N_19688,N_19736);
xor UO_202 (O_202,N_19836,N_19930);
nor UO_203 (O_203,N_19898,N_19816);
nand UO_204 (O_204,N_19826,N_19673);
and UO_205 (O_205,N_19634,N_19891);
or UO_206 (O_206,N_19972,N_19606);
or UO_207 (O_207,N_19838,N_19796);
or UO_208 (O_208,N_19998,N_19891);
xor UO_209 (O_209,N_19765,N_19666);
nand UO_210 (O_210,N_19815,N_19632);
or UO_211 (O_211,N_19729,N_19717);
and UO_212 (O_212,N_19917,N_19707);
or UO_213 (O_213,N_19725,N_19836);
and UO_214 (O_214,N_19956,N_19674);
xor UO_215 (O_215,N_19671,N_19615);
xor UO_216 (O_216,N_19685,N_19809);
and UO_217 (O_217,N_19926,N_19767);
and UO_218 (O_218,N_19919,N_19856);
nand UO_219 (O_219,N_19815,N_19828);
nand UO_220 (O_220,N_19983,N_19996);
xnor UO_221 (O_221,N_19665,N_19833);
nand UO_222 (O_222,N_19998,N_19892);
xor UO_223 (O_223,N_19602,N_19910);
and UO_224 (O_224,N_19980,N_19813);
and UO_225 (O_225,N_19914,N_19885);
or UO_226 (O_226,N_19789,N_19846);
and UO_227 (O_227,N_19947,N_19958);
nand UO_228 (O_228,N_19739,N_19978);
nand UO_229 (O_229,N_19881,N_19760);
nor UO_230 (O_230,N_19977,N_19690);
or UO_231 (O_231,N_19609,N_19752);
xor UO_232 (O_232,N_19811,N_19759);
or UO_233 (O_233,N_19930,N_19738);
xnor UO_234 (O_234,N_19992,N_19827);
and UO_235 (O_235,N_19912,N_19932);
xor UO_236 (O_236,N_19799,N_19774);
nand UO_237 (O_237,N_19978,N_19692);
nor UO_238 (O_238,N_19831,N_19748);
nand UO_239 (O_239,N_19904,N_19999);
or UO_240 (O_240,N_19628,N_19738);
or UO_241 (O_241,N_19987,N_19831);
or UO_242 (O_242,N_19805,N_19618);
nor UO_243 (O_243,N_19757,N_19865);
xnor UO_244 (O_244,N_19667,N_19819);
and UO_245 (O_245,N_19764,N_19936);
nor UO_246 (O_246,N_19829,N_19727);
and UO_247 (O_247,N_19626,N_19929);
or UO_248 (O_248,N_19959,N_19796);
xor UO_249 (O_249,N_19724,N_19822);
nor UO_250 (O_250,N_19692,N_19836);
and UO_251 (O_251,N_19690,N_19803);
nor UO_252 (O_252,N_19701,N_19994);
or UO_253 (O_253,N_19739,N_19883);
nor UO_254 (O_254,N_19822,N_19748);
nand UO_255 (O_255,N_19916,N_19884);
nand UO_256 (O_256,N_19718,N_19988);
and UO_257 (O_257,N_19866,N_19833);
or UO_258 (O_258,N_19684,N_19730);
xor UO_259 (O_259,N_19861,N_19668);
or UO_260 (O_260,N_19715,N_19926);
or UO_261 (O_261,N_19891,N_19833);
xor UO_262 (O_262,N_19641,N_19636);
nor UO_263 (O_263,N_19974,N_19852);
nor UO_264 (O_264,N_19831,N_19647);
xnor UO_265 (O_265,N_19865,N_19720);
or UO_266 (O_266,N_19756,N_19835);
xnor UO_267 (O_267,N_19832,N_19951);
nand UO_268 (O_268,N_19942,N_19750);
nor UO_269 (O_269,N_19645,N_19828);
and UO_270 (O_270,N_19952,N_19812);
xor UO_271 (O_271,N_19916,N_19636);
or UO_272 (O_272,N_19896,N_19858);
nor UO_273 (O_273,N_19981,N_19702);
or UO_274 (O_274,N_19905,N_19939);
or UO_275 (O_275,N_19821,N_19892);
and UO_276 (O_276,N_19895,N_19761);
xnor UO_277 (O_277,N_19649,N_19749);
or UO_278 (O_278,N_19760,N_19865);
or UO_279 (O_279,N_19660,N_19849);
xor UO_280 (O_280,N_19722,N_19924);
xor UO_281 (O_281,N_19970,N_19947);
nand UO_282 (O_282,N_19938,N_19681);
nor UO_283 (O_283,N_19615,N_19727);
xor UO_284 (O_284,N_19932,N_19661);
and UO_285 (O_285,N_19915,N_19847);
xnor UO_286 (O_286,N_19813,N_19918);
xor UO_287 (O_287,N_19919,N_19646);
nor UO_288 (O_288,N_19859,N_19975);
or UO_289 (O_289,N_19823,N_19880);
nand UO_290 (O_290,N_19992,N_19815);
xor UO_291 (O_291,N_19933,N_19738);
nand UO_292 (O_292,N_19727,N_19904);
nand UO_293 (O_293,N_19672,N_19880);
nor UO_294 (O_294,N_19608,N_19843);
and UO_295 (O_295,N_19967,N_19857);
and UO_296 (O_296,N_19723,N_19770);
xor UO_297 (O_297,N_19714,N_19668);
nand UO_298 (O_298,N_19682,N_19973);
xor UO_299 (O_299,N_19978,N_19892);
xnor UO_300 (O_300,N_19946,N_19615);
nor UO_301 (O_301,N_19751,N_19826);
and UO_302 (O_302,N_19954,N_19930);
nand UO_303 (O_303,N_19678,N_19661);
nor UO_304 (O_304,N_19680,N_19645);
nor UO_305 (O_305,N_19677,N_19709);
and UO_306 (O_306,N_19737,N_19650);
xor UO_307 (O_307,N_19914,N_19608);
xor UO_308 (O_308,N_19950,N_19766);
and UO_309 (O_309,N_19698,N_19959);
xor UO_310 (O_310,N_19986,N_19991);
nor UO_311 (O_311,N_19827,N_19601);
nor UO_312 (O_312,N_19602,N_19788);
xor UO_313 (O_313,N_19736,N_19968);
nand UO_314 (O_314,N_19800,N_19602);
and UO_315 (O_315,N_19827,N_19762);
nand UO_316 (O_316,N_19719,N_19808);
and UO_317 (O_317,N_19628,N_19888);
xor UO_318 (O_318,N_19659,N_19767);
nor UO_319 (O_319,N_19835,N_19719);
and UO_320 (O_320,N_19650,N_19666);
and UO_321 (O_321,N_19789,N_19717);
and UO_322 (O_322,N_19949,N_19793);
nand UO_323 (O_323,N_19906,N_19981);
nor UO_324 (O_324,N_19848,N_19735);
nor UO_325 (O_325,N_19890,N_19856);
nor UO_326 (O_326,N_19648,N_19628);
xnor UO_327 (O_327,N_19845,N_19770);
and UO_328 (O_328,N_19768,N_19679);
nor UO_329 (O_329,N_19653,N_19745);
or UO_330 (O_330,N_19878,N_19722);
nand UO_331 (O_331,N_19798,N_19987);
or UO_332 (O_332,N_19762,N_19931);
or UO_333 (O_333,N_19671,N_19715);
nor UO_334 (O_334,N_19930,N_19812);
nor UO_335 (O_335,N_19757,N_19658);
nand UO_336 (O_336,N_19867,N_19666);
or UO_337 (O_337,N_19674,N_19845);
or UO_338 (O_338,N_19876,N_19677);
nor UO_339 (O_339,N_19742,N_19616);
and UO_340 (O_340,N_19865,N_19920);
nor UO_341 (O_341,N_19895,N_19609);
or UO_342 (O_342,N_19731,N_19611);
nand UO_343 (O_343,N_19938,N_19668);
nand UO_344 (O_344,N_19642,N_19745);
or UO_345 (O_345,N_19836,N_19666);
nor UO_346 (O_346,N_19767,N_19722);
nand UO_347 (O_347,N_19813,N_19863);
and UO_348 (O_348,N_19994,N_19825);
xnor UO_349 (O_349,N_19659,N_19648);
nand UO_350 (O_350,N_19843,N_19647);
xnor UO_351 (O_351,N_19601,N_19977);
xor UO_352 (O_352,N_19605,N_19999);
and UO_353 (O_353,N_19859,N_19901);
and UO_354 (O_354,N_19990,N_19720);
nand UO_355 (O_355,N_19698,N_19838);
or UO_356 (O_356,N_19607,N_19811);
nor UO_357 (O_357,N_19616,N_19810);
or UO_358 (O_358,N_19946,N_19935);
and UO_359 (O_359,N_19708,N_19996);
and UO_360 (O_360,N_19997,N_19658);
and UO_361 (O_361,N_19811,N_19926);
or UO_362 (O_362,N_19830,N_19625);
or UO_363 (O_363,N_19812,N_19773);
or UO_364 (O_364,N_19979,N_19923);
xnor UO_365 (O_365,N_19987,N_19875);
or UO_366 (O_366,N_19852,N_19850);
or UO_367 (O_367,N_19624,N_19757);
xor UO_368 (O_368,N_19808,N_19616);
nor UO_369 (O_369,N_19679,N_19663);
nor UO_370 (O_370,N_19905,N_19940);
and UO_371 (O_371,N_19883,N_19806);
and UO_372 (O_372,N_19640,N_19849);
and UO_373 (O_373,N_19962,N_19611);
or UO_374 (O_374,N_19941,N_19796);
nand UO_375 (O_375,N_19900,N_19988);
and UO_376 (O_376,N_19633,N_19688);
nor UO_377 (O_377,N_19685,N_19818);
nand UO_378 (O_378,N_19791,N_19698);
and UO_379 (O_379,N_19997,N_19623);
or UO_380 (O_380,N_19844,N_19933);
xnor UO_381 (O_381,N_19975,N_19700);
nand UO_382 (O_382,N_19843,N_19938);
nor UO_383 (O_383,N_19966,N_19611);
and UO_384 (O_384,N_19934,N_19841);
or UO_385 (O_385,N_19623,N_19765);
or UO_386 (O_386,N_19758,N_19852);
and UO_387 (O_387,N_19702,N_19758);
or UO_388 (O_388,N_19883,N_19899);
nand UO_389 (O_389,N_19605,N_19840);
and UO_390 (O_390,N_19875,N_19701);
or UO_391 (O_391,N_19964,N_19826);
nor UO_392 (O_392,N_19624,N_19771);
nor UO_393 (O_393,N_19701,N_19709);
and UO_394 (O_394,N_19963,N_19911);
nor UO_395 (O_395,N_19943,N_19946);
or UO_396 (O_396,N_19659,N_19969);
nor UO_397 (O_397,N_19783,N_19679);
nor UO_398 (O_398,N_19624,N_19792);
nor UO_399 (O_399,N_19684,N_19789);
and UO_400 (O_400,N_19900,N_19817);
xor UO_401 (O_401,N_19842,N_19975);
nor UO_402 (O_402,N_19685,N_19738);
and UO_403 (O_403,N_19839,N_19672);
or UO_404 (O_404,N_19982,N_19702);
or UO_405 (O_405,N_19823,N_19905);
nand UO_406 (O_406,N_19638,N_19734);
nand UO_407 (O_407,N_19618,N_19789);
nand UO_408 (O_408,N_19818,N_19724);
nor UO_409 (O_409,N_19788,N_19781);
xor UO_410 (O_410,N_19821,N_19974);
xnor UO_411 (O_411,N_19670,N_19926);
xnor UO_412 (O_412,N_19744,N_19629);
and UO_413 (O_413,N_19616,N_19907);
nand UO_414 (O_414,N_19623,N_19970);
xor UO_415 (O_415,N_19794,N_19832);
or UO_416 (O_416,N_19751,N_19726);
xor UO_417 (O_417,N_19619,N_19711);
or UO_418 (O_418,N_19856,N_19629);
and UO_419 (O_419,N_19815,N_19874);
or UO_420 (O_420,N_19661,N_19844);
and UO_421 (O_421,N_19767,N_19725);
nand UO_422 (O_422,N_19837,N_19686);
xnor UO_423 (O_423,N_19728,N_19723);
nand UO_424 (O_424,N_19856,N_19685);
nand UO_425 (O_425,N_19873,N_19757);
or UO_426 (O_426,N_19878,N_19617);
and UO_427 (O_427,N_19836,N_19611);
or UO_428 (O_428,N_19947,N_19898);
xnor UO_429 (O_429,N_19704,N_19888);
nand UO_430 (O_430,N_19655,N_19903);
nor UO_431 (O_431,N_19617,N_19600);
and UO_432 (O_432,N_19648,N_19612);
and UO_433 (O_433,N_19748,N_19909);
and UO_434 (O_434,N_19715,N_19805);
nand UO_435 (O_435,N_19616,N_19896);
xnor UO_436 (O_436,N_19749,N_19943);
or UO_437 (O_437,N_19619,N_19740);
xor UO_438 (O_438,N_19622,N_19889);
or UO_439 (O_439,N_19788,N_19797);
and UO_440 (O_440,N_19895,N_19973);
or UO_441 (O_441,N_19981,N_19666);
or UO_442 (O_442,N_19622,N_19772);
and UO_443 (O_443,N_19898,N_19770);
nor UO_444 (O_444,N_19712,N_19783);
or UO_445 (O_445,N_19749,N_19761);
nor UO_446 (O_446,N_19801,N_19889);
and UO_447 (O_447,N_19940,N_19981);
or UO_448 (O_448,N_19910,N_19681);
or UO_449 (O_449,N_19667,N_19762);
nand UO_450 (O_450,N_19959,N_19996);
nor UO_451 (O_451,N_19774,N_19986);
and UO_452 (O_452,N_19952,N_19654);
nand UO_453 (O_453,N_19947,N_19919);
or UO_454 (O_454,N_19700,N_19651);
xnor UO_455 (O_455,N_19882,N_19732);
and UO_456 (O_456,N_19948,N_19667);
or UO_457 (O_457,N_19791,N_19779);
xnor UO_458 (O_458,N_19663,N_19952);
nor UO_459 (O_459,N_19685,N_19671);
nor UO_460 (O_460,N_19831,N_19872);
or UO_461 (O_461,N_19876,N_19780);
nand UO_462 (O_462,N_19786,N_19817);
xnor UO_463 (O_463,N_19957,N_19687);
and UO_464 (O_464,N_19635,N_19795);
and UO_465 (O_465,N_19932,N_19854);
xor UO_466 (O_466,N_19719,N_19952);
nor UO_467 (O_467,N_19812,N_19754);
xnor UO_468 (O_468,N_19886,N_19996);
nand UO_469 (O_469,N_19852,N_19711);
nand UO_470 (O_470,N_19834,N_19641);
or UO_471 (O_471,N_19811,N_19639);
and UO_472 (O_472,N_19871,N_19761);
nand UO_473 (O_473,N_19758,N_19896);
xor UO_474 (O_474,N_19686,N_19869);
or UO_475 (O_475,N_19802,N_19943);
or UO_476 (O_476,N_19912,N_19744);
or UO_477 (O_477,N_19902,N_19685);
nand UO_478 (O_478,N_19720,N_19967);
nand UO_479 (O_479,N_19603,N_19909);
nand UO_480 (O_480,N_19784,N_19825);
nor UO_481 (O_481,N_19631,N_19830);
and UO_482 (O_482,N_19658,N_19717);
nor UO_483 (O_483,N_19654,N_19881);
nor UO_484 (O_484,N_19601,N_19990);
nor UO_485 (O_485,N_19811,N_19932);
nand UO_486 (O_486,N_19970,N_19635);
nand UO_487 (O_487,N_19929,N_19903);
xor UO_488 (O_488,N_19782,N_19986);
or UO_489 (O_489,N_19617,N_19831);
nor UO_490 (O_490,N_19805,N_19808);
and UO_491 (O_491,N_19809,N_19965);
xor UO_492 (O_492,N_19798,N_19707);
nor UO_493 (O_493,N_19807,N_19988);
or UO_494 (O_494,N_19723,N_19962);
nor UO_495 (O_495,N_19912,N_19639);
or UO_496 (O_496,N_19913,N_19836);
and UO_497 (O_497,N_19736,N_19910);
xor UO_498 (O_498,N_19903,N_19652);
and UO_499 (O_499,N_19932,N_19853);
xor UO_500 (O_500,N_19718,N_19964);
nor UO_501 (O_501,N_19991,N_19712);
or UO_502 (O_502,N_19617,N_19950);
xnor UO_503 (O_503,N_19760,N_19697);
and UO_504 (O_504,N_19688,N_19954);
nor UO_505 (O_505,N_19729,N_19783);
xnor UO_506 (O_506,N_19786,N_19985);
nor UO_507 (O_507,N_19662,N_19802);
nor UO_508 (O_508,N_19793,N_19750);
xor UO_509 (O_509,N_19784,N_19785);
xor UO_510 (O_510,N_19791,N_19805);
and UO_511 (O_511,N_19783,N_19615);
nand UO_512 (O_512,N_19965,N_19668);
nor UO_513 (O_513,N_19995,N_19906);
nand UO_514 (O_514,N_19819,N_19680);
and UO_515 (O_515,N_19993,N_19746);
or UO_516 (O_516,N_19678,N_19972);
nor UO_517 (O_517,N_19927,N_19802);
nand UO_518 (O_518,N_19674,N_19724);
nor UO_519 (O_519,N_19625,N_19745);
and UO_520 (O_520,N_19699,N_19679);
nor UO_521 (O_521,N_19601,N_19896);
xnor UO_522 (O_522,N_19948,N_19796);
and UO_523 (O_523,N_19637,N_19607);
nor UO_524 (O_524,N_19946,N_19651);
or UO_525 (O_525,N_19788,N_19809);
and UO_526 (O_526,N_19898,N_19711);
or UO_527 (O_527,N_19961,N_19845);
nor UO_528 (O_528,N_19689,N_19899);
or UO_529 (O_529,N_19829,N_19846);
xnor UO_530 (O_530,N_19916,N_19689);
nand UO_531 (O_531,N_19956,N_19806);
xnor UO_532 (O_532,N_19773,N_19926);
or UO_533 (O_533,N_19868,N_19689);
nand UO_534 (O_534,N_19781,N_19926);
and UO_535 (O_535,N_19989,N_19725);
and UO_536 (O_536,N_19730,N_19612);
nor UO_537 (O_537,N_19774,N_19794);
and UO_538 (O_538,N_19666,N_19661);
and UO_539 (O_539,N_19940,N_19975);
nand UO_540 (O_540,N_19699,N_19655);
nand UO_541 (O_541,N_19911,N_19771);
xor UO_542 (O_542,N_19941,N_19703);
nand UO_543 (O_543,N_19606,N_19861);
xor UO_544 (O_544,N_19703,N_19705);
xnor UO_545 (O_545,N_19705,N_19672);
nand UO_546 (O_546,N_19813,N_19789);
nor UO_547 (O_547,N_19981,N_19870);
nand UO_548 (O_548,N_19879,N_19691);
nor UO_549 (O_549,N_19805,N_19622);
and UO_550 (O_550,N_19628,N_19863);
nor UO_551 (O_551,N_19742,N_19812);
nor UO_552 (O_552,N_19948,N_19601);
nand UO_553 (O_553,N_19808,N_19726);
or UO_554 (O_554,N_19761,N_19693);
xnor UO_555 (O_555,N_19831,N_19784);
nand UO_556 (O_556,N_19693,N_19973);
nor UO_557 (O_557,N_19970,N_19974);
nor UO_558 (O_558,N_19722,N_19984);
and UO_559 (O_559,N_19799,N_19843);
and UO_560 (O_560,N_19917,N_19681);
nor UO_561 (O_561,N_19639,N_19844);
and UO_562 (O_562,N_19826,N_19889);
xnor UO_563 (O_563,N_19813,N_19916);
nand UO_564 (O_564,N_19976,N_19709);
xor UO_565 (O_565,N_19601,N_19978);
nor UO_566 (O_566,N_19745,N_19954);
and UO_567 (O_567,N_19764,N_19870);
or UO_568 (O_568,N_19871,N_19601);
nor UO_569 (O_569,N_19835,N_19891);
and UO_570 (O_570,N_19935,N_19624);
nand UO_571 (O_571,N_19693,N_19701);
nor UO_572 (O_572,N_19757,N_19656);
nor UO_573 (O_573,N_19634,N_19760);
or UO_574 (O_574,N_19986,N_19999);
or UO_575 (O_575,N_19945,N_19908);
and UO_576 (O_576,N_19762,N_19726);
xor UO_577 (O_577,N_19653,N_19824);
xnor UO_578 (O_578,N_19717,N_19852);
nor UO_579 (O_579,N_19657,N_19655);
or UO_580 (O_580,N_19890,N_19739);
nor UO_581 (O_581,N_19649,N_19686);
nand UO_582 (O_582,N_19942,N_19713);
or UO_583 (O_583,N_19640,N_19905);
or UO_584 (O_584,N_19632,N_19997);
and UO_585 (O_585,N_19815,N_19818);
nor UO_586 (O_586,N_19621,N_19634);
or UO_587 (O_587,N_19806,N_19959);
and UO_588 (O_588,N_19835,N_19787);
nand UO_589 (O_589,N_19813,N_19958);
nor UO_590 (O_590,N_19605,N_19775);
nor UO_591 (O_591,N_19952,N_19912);
or UO_592 (O_592,N_19866,N_19748);
xor UO_593 (O_593,N_19852,N_19995);
or UO_594 (O_594,N_19955,N_19993);
nor UO_595 (O_595,N_19621,N_19954);
xnor UO_596 (O_596,N_19805,N_19743);
or UO_597 (O_597,N_19902,N_19957);
xor UO_598 (O_598,N_19906,N_19619);
xnor UO_599 (O_599,N_19617,N_19894);
xnor UO_600 (O_600,N_19934,N_19860);
and UO_601 (O_601,N_19907,N_19891);
and UO_602 (O_602,N_19964,N_19930);
xor UO_603 (O_603,N_19771,N_19985);
and UO_604 (O_604,N_19965,N_19764);
nor UO_605 (O_605,N_19665,N_19957);
or UO_606 (O_606,N_19795,N_19923);
nand UO_607 (O_607,N_19956,N_19668);
nand UO_608 (O_608,N_19914,N_19823);
nor UO_609 (O_609,N_19928,N_19618);
xor UO_610 (O_610,N_19886,N_19893);
and UO_611 (O_611,N_19682,N_19701);
or UO_612 (O_612,N_19916,N_19701);
nand UO_613 (O_613,N_19981,N_19834);
xnor UO_614 (O_614,N_19746,N_19861);
xor UO_615 (O_615,N_19644,N_19821);
and UO_616 (O_616,N_19801,N_19668);
xnor UO_617 (O_617,N_19729,N_19994);
xor UO_618 (O_618,N_19641,N_19710);
nand UO_619 (O_619,N_19750,N_19649);
or UO_620 (O_620,N_19746,N_19957);
or UO_621 (O_621,N_19861,N_19739);
nor UO_622 (O_622,N_19885,N_19949);
nand UO_623 (O_623,N_19916,N_19784);
nand UO_624 (O_624,N_19777,N_19677);
xnor UO_625 (O_625,N_19878,N_19629);
or UO_626 (O_626,N_19721,N_19782);
xnor UO_627 (O_627,N_19784,N_19883);
and UO_628 (O_628,N_19771,N_19744);
xor UO_629 (O_629,N_19803,N_19743);
or UO_630 (O_630,N_19884,N_19841);
nand UO_631 (O_631,N_19962,N_19889);
or UO_632 (O_632,N_19611,N_19834);
nand UO_633 (O_633,N_19820,N_19910);
or UO_634 (O_634,N_19893,N_19904);
nor UO_635 (O_635,N_19671,N_19963);
xnor UO_636 (O_636,N_19964,N_19909);
nor UO_637 (O_637,N_19947,N_19965);
nand UO_638 (O_638,N_19702,N_19899);
or UO_639 (O_639,N_19624,N_19995);
nor UO_640 (O_640,N_19689,N_19770);
or UO_641 (O_641,N_19987,N_19858);
nor UO_642 (O_642,N_19934,N_19788);
nor UO_643 (O_643,N_19715,N_19631);
and UO_644 (O_644,N_19743,N_19739);
nand UO_645 (O_645,N_19635,N_19993);
nor UO_646 (O_646,N_19600,N_19921);
and UO_647 (O_647,N_19842,N_19670);
nand UO_648 (O_648,N_19803,N_19716);
and UO_649 (O_649,N_19810,N_19956);
xnor UO_650 (O_650,N_19757,N_19818);
nor UO_651 (O_651,N_19717,N_19837);
xnor UO_652 (O_652,N_19881,N_19655);
nand UO_653 (O_653,N_19906,N_19606);
and UO_654 (O_654,N_19640,N_19954);
nor UO_655 (O_655,N_19914,N_19799);
or UO_656 (O_656,N_19986,N_19715);
and UO_657 (O_657,N_19973,N_19823);
or UO_658 (O_658,N_19703,N_19748);
and UO_659 (O_659,N_19883,N_19778);
xnor UO_660 (O_660,N_19688,N_19714);
and UO_661 (O_661,N_19690,N_19662);
nand UO_662 (O_662,N_19738,N_19828);
or UO_663 (O_663,N_19799,N_19766);
and UO_664 (O_664,N_19685,N_19618);
nand UO_665 (O_665,N_19605,N_19752);
or UO_666 (O_666,N_19650,N_19608);
or UO_667 (O_667,N_19691,N_19904);
or UO_668 (O_668,N_19893,N_19704);
nand UO_669 (O_669,N_19631,N_19955);
or UO_670 (O_670,N_19920,N_19761);
xor UO_671 (O_671,N_19836,N_19790);
nand UO_672 (O_672,N_19911,N_19622);
nor UO_673 (O_673,N_19873,N_19834);
and UO_674 (O_674,N_19631,N_19803);
xor UO_675 (O_675,N_19738,N_19730);
or UO_676 (O_676,N_19725,N_19829);
xnor UO_677 (O_677,N_19923,N_19874);
nand UO_678 (O_678,N_19937,N_19713);
xor UO_679 (O_679,N_19673,N_19751);
nand UO_680 (O_680,N_19869,N_19893);
nand UO_681 (O_681,N_19907,N_19924);
or UO_682 (O_682,N_19769,N_19761);
nand UO_683 (O_683,N_19936,N_19756);
or UO_684 (O_684,N_19918,N_19605);
nand UO_685 (O_685,N_19928,N_19829);
and UO_686 (O_686,N_19841,N_19972);
nand UO_687 (O_687,N_19883,N_19759);
nand UO_688 (O_688,N_19980,N_19708);
nor UO_689 (O_689,N_19808,N_19884);
nor UO_690 (O_690,N_19972,N_19736);
and UO_691 (O_691,N_19852,N_19915);
and UO_692 (O_692,N_19672,N_19830);
or UO_693 (O_693,N_19627,N_19866);
and UO_694 (O_694,N_19870,N_19868);
xnor UO_695 (O_695,N_19957,N_19873);
nor UO_696 (O_696,N_19741,N_19611);
nand UO_697 (O_697,N_19921,N_19711);
nor UO_698 (O_698,N_19729,N_19713);
or UO_699 (O_699,N_19694,N_19754);
or UO_700 (O_700,N_19818,N_19787);
and UO_701 (O_701,N_19687,N_19758);
or UO_702 (O_702,N_19871,N_19748);
nor UO_703 (O_703,N_19699,N_19795);
or UO_704 (O_704,N_19771,N_19874);
nor UO_705 (O_705,N_19719,N_19999);
nand UO_706 (O_706,N_19754,N_19619);
and UO_707 (O_707,N_19961,N_19749);
or UO_708 (O_708,N_19990,N_19933);
and UO_709 (O_709,N_19892,N_19873);
nand UO_710 (O_710,N_19888,N_19871);
nor UO_711 (O_711,N_19739,N_19679);
nor UO_712 (O_712,N_19820,N_19662);
nor UO_713 (O_713,N_19872,N_19900);
nor UO_714 (O_714,N_19722,N_19978);
nand UO_715 (O_715,N_19980,N_19906);
and UO_716 (O_716,N_19952,N_19976);
nor UO_717 (O_717,N_19689,N_19762);
and UO_718 (O_718,N_19969,N_19733);
nand UO_719 (O_719,N_19790,N_19772);
nand UO_720 (O_720,N_19773,N_19754);
nor UO_721 (O_721,N_19982,N_19958);
xor UO_722 (O_722,N_19761,N_19813);
or UO_723 (O_723,N_19887,N_19706);
or UO_724 (O_724,N_19807,N_19754);
and UO_725 (O_725,N_19776,N_19863);
xor UO_726 (O_726,N_19696,N_19870);
nor UO_727 (O_727,N_19690,N_19795);
nor UO_728 (O_728,N_19732,N_19673);
and UO_729 (O_729,N_19653,N_19934);
and UO_730 (O_730,N_19685,N_19973);
xor UO_731 (O_731,N_19613,N_19801);
xnor UO_732 (O_732,N_19630,N_19621);
nand UO_733 (O_733,N_19849,N_19844);
nand UO_734 (O_734,N_19710,N_19901);
or UO_735 (O_735,N_19720,N_19833);
xor UO_736 (O_736,N_19912,N_19713);
and UO_737 (O_737,N_19944,N_19833);
or UO_738 (O_738,N_19620,N_19625);
and UO_739 (O_739,N_19791,N_19775);
nor UO_740 (O_740,N_19865,N_19840);
or UO_741 (O_741,N_19665,N_19647);
or UO_742 (O_742,N_19910,N_19986);
or UO_743 (O_743,N_19615,N_19841);
nor UO_744 (O_744,N_19664,N_19815);
or UO_745 (O_745,N_19979,N_19977);
xnor UO_746 (O_746,N_19682,N_19915);
xor UO_747 (O_747,N_19745,N_19611);
nand UO_748 (O_748,N_19804,N_19896);
xnor UO_749 (O_749,N_19883,N_19983);
and UO_750 (O_750,N_19616,N_19911);
nor UO_751 (O_751,N_19975,N_19953);
nor UO_752 (O_752,N_19626,N_19665);
xor UO_753 (O_753,N_19812,N_19631);
nand UO_754 (O_754,N_19783,N_19784);
xnor UO_755 (O_755,N_19805,N_19842);
and UO_756 (O_756,N_19808,N_19932);
nand UO_757 (O_757,N_19954,N_19600);
and UO_758 (O_758,N_19629,N_19817);
xnor UO_759 (O_759,N_19815,N_19622);
nor UO_760 (O_760,N_19810,N_19919);
and UO_761 (O_761,N_19952,N_19874);
nor UO_762 (O_762,N_19831,N_19687);
nand UO_763 (O_763,N_19823,N_19966);
and UO_764 (O_764,N_19915,N_19861);
or UO_765 (O_765,N_19777,N_19742);
nor UO_766 (O_766,N_19865,N_19813);
nand UO_767 (O_767,N_19826,N_19908);
or UO_768 (O_768,N_19609,N_19995);
nor UO_769 (O_769,N_19756,N_19966);
nor UO_770 (O_770,N_19875,N_19889);
or UO_771 (O_771,N_19985,N_19879);
nand UO_772 (O_772,N_19696,N_19624);
xnor UO_773 (O_773,N_19858,N_19693);
nor UO_774 (O_774,N_19845,N_19900);
nand UO_775 (O_775,N_19926,N_19760);
xor UO_776 (O_776,N_19948,N_19725);
nor UO_777 (O_777,N_19823,N_19868);
nand UO_778 (O_778,N_19911,N_19818);
nor UO_779 (O_779,N_19906,N_19975);
xor UO_780 (O_780,N_19742,N_19955);
nor UO_781 (O_781,N_19969,N_19845);
and UO_782 (O_782,N_19941,N_19698);
and UO_783 (O_783,N_19933,N_19714);
and UO_784 (O_784,N_19767,N_19995);
or UO_785 (O_785,N_19863,N_19864);
xor UO_786 (O_786,N_19806,N_19808);
nand UO_787 (O_787,N_19658,N_19905);
nor UO_788 (O_788,N_19771,N_19883);
or UO_789 (O_789,N_19780,N_19827);
or UO_790 (O_790,N_19836,N_19899);
and UO_791 (O_791,N_19974,N_19954);
or UO_792 (O_792,N_19811,N_19883);
or UO_793 (O_793,N_19810,N_19682);
nor UO_794 (O_794,N_19668,N_19684);
nor UO_795 (O_795,N_19975,N_19662);
or UO_796 (O_796,N_19710,N_19786);
and UO_797 (O_797,N_19674,N_19640);
nor UO_798 (O_798,N_19912,N_19611);
nor UO_799 (O_799,N_19976,N_19625);
xnor UO_800 (O_800,N_19862,N_19685);
or UO_801 (O_801,N_19655,N_19909);
nor UO_802 (O_802,N_19892,N_19832);
xor UO_803 (O_803,N_19792,N_19896);
nand UO_804 (O_804,N_19744,N_19752);
nor UO_805 (O_805,N_19978,N_19687);
or UO_806 (O_806,N_19799,N_19699);
or UO_807 (O_807,N_19675,N_19853);
or UO_808 (O_808,N_19837,N_19939);
nor UO_809 (O_809,N_19860,N_19963);
xnor UO_810 (O_810,N_19772,N_19731);
xor UO_811 (O_811,N_19884,N_19756);
or UO_812 (O_812,N_19949,N_19993);
nor UO_813 (O_813,N_19966,N_19771);
nand UO_814 (O_814,N_19625,N_19601);
nand UO_815 (O_815,N_19777,N_19636);
nand UO_816 (O_816,N_19600,N_19667);
and UO_817 (O_817,N_19776,N_19668);
nor UO_818 (O_818,N_19658,N_19798);
and UO_819 (O_819,N_19665,N_19610);
nor UO_820 (O_820,N_19744,N_19995);
or UO_821 (O_821,N_19798,N_19873);
or UO_822 (O_822,N_19885,N_19736);
and UO_823 (O_823,N_19686,N_19669);
xnor UO_824 (O_824,N_19992,N_19980);
nand UO_825 (O_825,N_19966,N_19603);
xor UO_826 (O_826,N_19912,N_19619);
and UO_827 (O_827,N_19634,N_19846);
nand UO_828 (O_828,N_19770,N_19800);
xnor UO_829 (O_829,N_19696,N_19718);
and UO_830 (O_830,N_19993,N_19855);
nand UO_831 (O_831,N_19972,N_19665);
nand UO_832 (O_832,N_19700,N_19612);
nor UO_833 (O_833,N_19842,N_19865);
nand UO_834 (O_834,N_19796,N_19901);
nand UO_835 (O_835,N_19652,N_19661);
nor UO_836 (O_836,N_19987,N_19978);
or UO_837 (O_837,N_19624,N_19781);
nand UO_838 (O_838,N_19655,N_19813);
or UO_839 (O_839,N_19660,N_19930);
nor UO_840 (O_840,N_19956,N_19823);
xor UO_841 (O_841,N_19606,N_19676);
and UO_842 (O_842,N_19638,N_19835);
and UO_843 (O_843,N_19744,N_19734);
or UO_844 (O_844,N_19809,N_19895);
nor UO_845 (O_845,N_19703,N_19640);
xor UO_846 (O_846,N_19892,N_19952);
and UO_847 (O_847,N_19828,N_19808);
nand UO_848 (O_848,N_19725,N_19960);
nand UO_849 (O_849,N_19662,N_19792);
or UO_850 (O_850,N_19853,N_19852);
xor UO_851 (O_851,N_19852,N_19991);
nor UO_852 (O_852,N_19980,N_19993);
and UO_853 (O_853,N_19737,N_19986);
nor UO_854 (O_854,N_19827,N_19859);
and UO_855 (O_855,N_19875,N_19828);
xor UO_856 (O_856,N_19642,N_19715);
and UO_857 (O_857,N_19747,N_19989);
nand UO_858 (O_858,N_19671,N_19926);
and UO_859 (O_859,N_19874,N_19656);
xnor UO_860 (O_860,N_19805,N_19875);
nor UO_861 (O_861,N_19894,N_19640);
nand UO_862 (O_862,N_19704,N_19887);
nor UO_863 (O_863,N_19940,N_19868);
or UO_864 (O_864,N_19927,N_19976);
nor UO_865 (O_865,N_19780,N_19795);
or UO_866 (O_866,N_19707,N_19741);
nand UO_867 (O_867,N_19871,N_19927);
xnor UO_868 (O_868,N_19819,N_19763);
xor UO_869 (O_869,N_19725,N_19794);
nand UO_870 (O_870,N_19696,N_19781);
or UO_871 (O_871,N_19694,N_19964);
xor UO_872 (O_872,N_19883,N_19842);
nand UO_873 (O_873,N_19934,N_19846);
nor UO_874 (O_874,N_19693,N_19821);
xnor UO_875 (O_875,N_19829,N_19880);
nand UO_876 (O_876,N_19935,N_19857);
nand UO_877 (O_877,N_19610,N_19950);
and UO_878 (O_878,N_19766,N_19810);
nand UO_879 (O_879,N_19661,N_19879);
xnor UO_880 (O_880,N_19888,N_19759);
nand UO_881 (O_881,N_19843,N_19676);
xor UO_882 (O_882,N_19797,N_19886);
or UO_883 (O_883,N_19796,N_19921);
or UO_884 (O_884,N_19876,N_19782);
nor UO_885 (O_885,N_19717,N_19766);
and UO_886 (O_886,N_19889,N_19818);
and UO_887 (O_887,N_19663,N_19900);
and UO_888 (O_888,N_19867,N_19755);
nor UO_889 (O_889,N_19906,N_19617);
and UO_890 (O_890,N_19669,N_19773);
xor UO_891 (O_891,N_19641,N_19721);
nor UO_892 (O_892,N_19855,N_19713);
or UO_893 (O_893,N_19891,N_19950);
and UO_894 (O_894,N_19947,N_19655);
and UO_895 (O_895,N_19917,N_19656);
nor UO_896 (O_896,N_19602,N_19968);
xor UO_897 (O_897,N_19600,N_19688);
and UO_898 (O_898,N_19894,N_19698);
and UO_899 (O_899,N_19790,N_19717);
nand UO_900 (O_900,N_19840,N_19949);
nor UO_901 (O_901,N_19708,N_19620);
xnor UO_902 (O_902,N_19801,N_19756);
nand UO_903 (O_903,N_19890,N_19907);
xor UO_904 (O_904,N_19681,N_19684);
nor UO_905 (O_905,N_19699,N_19895);
or UO_906 (O_906,N_19659,N_19813);
and UO_907 (O_907,N_19819,N_19858);
and UO_908 (O_908,N_19704,N_19817);
or UO_909 (O_909,N_19892,N_19754);
or UO_910 (O_910,N_19650,N_19738);
and UO_911 (O_911,N_19722,N_19711);
or UO_912 (O_912,N_19857,N_19851);
nor UO_913 (O_913,N_19657,N_19746);
nor UO_914 (O_914,N_19935,N_19715);
and UO_915 (O_915,N_19944,N_19760);
nand UO_916 (O_916,N_19937,N_19914);
nor UO_917 (O_917,N_19652,N_19739);
nand UO_918 (O_918,N_19693,N_19686);
and UO_919 (O_919,N_19793,N_19934);
xor UO_920 (O_920,N_19832,N_19954);
nand UO_921 (O_921,N_19886,N_19943);
or UO_922 (O_922,N_19683,N_19834);
and UO_923 (O_923,N_19943,N_19727);
or UO_924 (O_924,N_19689,N_19980);
nor UO_925 (O_925,N_19668,N_19870);
or UO_926 (O_926,N_19923,N_19848);
nand UO_927 (O_927,N_19686,N_19788);
or UO_928 (O_928,N_19934,N_19858);
or UO_929 (O_929,N_19860,N_19942);
nor UO_930 (O_930,N_19799,N_19681);
or UO_931 (O_931,N_19844,N_19901);
nand UO_932 (O_932,N_19650,N_19743);
or UO_933 (O_933,N_19685,N_19752);
xnor UO_934 (O_934,N_19809,N_19828);
xnor UO_935 (O_935,N_19943,N_19888);
xor UO_936 (O_936,N_19769,N_19629);
nor UO_937 (O_937,N_19967,N_19658);
and UO_938 (O_938,N_19701,N_19937);
and UO_939 (O_939,N_19805,N_19676);
xnor UO_940 (O_940,N_19851,N_19872);
or UO_941 (O_941,N_19650,N_19698);
xor UO_942 (O_942,N_19783,N_19791);
and UO_943 (O_943,N_19930,N_19668);
nor UO_944 (O_944,N_19806,N_19717);
or UO_945 (O_945,N_19786,N_19840);
or UO_946 (O_946,N_19848,N_19672);
nand UO_947 (O_947,N_19607,N_19928);
nor UO_948 (O_948,N_19679,N_19875);
nor UO_949 (O_949,N_19865,N_19662);
nor UO_950 (O_950,N_19770,N_19965);
and UO_951 (O_951,N_19650,N_19840);
nand UO_952 (O_952,N_19843,N_19612);
nand UO_953 (O_953,N_19645,N_19793);
xnor UO_954 (O_954,N_19746,N_19929);
or UO_955 (O_955,N_19615,N_19719);
and UO_956 (O_956,N_19961,N_19747);
and UO_957 (O_957,N_19828,N_19713);
or UO_958 (O_958,N_19768,N_19864);
nor UO_959 (O_959,N_19919,N_19874);
and UO_960 (O_960,N_19839,N_19851);
or UO_961 (O_961,N_19938,N_19780);
nor UO_962 (O_962,N_19943,N_19761);
or UO_963 (O_963,N_19706,N_19657);
nor UO_964 (O_964,N_19866,N_19802);
xor UO_965 (O_965,N_19882,N_19667);
or UO_966 (O_966,N_19864,N_19990);
nor UO_967 (O_967,N_19884,N_19664);
xnor UO_968 (O_968,N_19692,N_19917);
or UO_969 (O_969,N_19791,N_19700);
and UO_970 (O_970,N_19683,N_19719);
and UO_971 (O_971,N_19850,N_19724);
or UO_972 (O_972,N_19970,N_19842);
or UO_973 (O_973,N_19947,N_19906);
nand UO_974 (O_974,N_19760,N_19960);
xor UO_975 (O_975,N_19933,N_19783);
or UO_976 (O_976,N_19681,N_19775);
xnor UO_977 (O_977,N_19830,N_19851);
and UO_978 (O_978,N_19743,N_19686);
xor UO_979 (O_979,N_19662,N_19766);
xnor UO_980 (O_980,N_19798,N_19688);
and UO_981 (O_981,N_19973,N_19817);
or UO_982 (O_982,N_19709,N_19973);
or UO_983 (O_983,N_19944,N_19832);
nor UO_984 (O_984,N_19731,N_19878);
xnor UO_985 (O_985,N_19685,N_19697);
and UO_986 (O_986,N_19697,N_19696);
or UO_987 (O_987,N_19942,N_19958);
nand UO_988 (O_988,N_19607,N_19740);
nor UO_989 (O_989,N_19708,N_19738);
or UO_990 (O_990,N_19739,N_19616);
or UO_991 (O_991,N_19845,N_19963);
xor UO_992 (O_992,N_19963,N_19772);
nand UO_993 (O_993,N_19676,N_19973);
nor UO_994 (O_994,N_19941,N_19729);
nand UO_995 (O_995,N_19847,N_19742);
and UO_996 (O_996,N_19732,N_19961);
xnor UO_997 (O_997,N_19673,N_19915);
xor UO_998 (O_998,N_19917,N_19778);
xnor UO_999 (O_999,N_19806,N_19782);
and UO_1000 (O_1000,N_19947,N_19972);
or UO_1001 (O_1001,N_19848,N_19821);
nor UO_1002 (O_1002,N_19715,N_19740);
nand UO_1003 (O_1003,N_19795,N_19662);
nand UO_1004 (O_1004,N_19798,N_19636);
nor UO_1005 (O_1005,N_19950,N_19872);
nand UO_1006 (O_1006,N_19757,N_19814);
nor UO_1007 (O_1007,N_19646,N_19698);
nand UO_1008 (O_1008,N_19852,N_19998);
or UO_1009 (O_1009,N_19702,N_19897);
xnor UO_1010 (O_1010,N_19917,N_19841);
nand UO_1011 (O_1011,N_19831,N_19866);
nand UO_1012 (O_1012,N_19976,N_19918);
and UO_1013 (O_1013,N_19818,N_19814);
nand UO_1014 (O_1014,N_19686,N_19720);
xor UO_1015 (O_1015,N_19628,N_19844);
xor UO_1016 (O_1016,N_19623,N_19633);
nor UO_1017 (O_1017,N_19883,N_19949);
and UO_1018 (O_1018,N_19794,N_19951);
xnor UO_1019 (O_1019,N_19931,N_19627);
and UO_1020 (O_1020,N_19856,N_19648);
nand UO_1021 (O_1021,N_19759,N_19907);
nor UO_1022 (O_1022,N_19692,N_19803);
or UO_1023 (O_1023,N_19853,N_19837);
nor UO_1024 (O_1024,N_19800,N_19852);
nand UO_1025 (O_1025,N_19800,N_19724);
or UO_1026 (O_1026,N_19900,N_19665);
xor UO_1027 (O_1027,N_19773,N_19676);
xor UO_1028 (O_1028,N_19631,N_19675);
xor UO_1029 (O_1029,N_19631,N_19848);
or UO_1030 (O_1030,N_19841,N_19753);
nor UO_1031 (O_1031,N_19887,N_19908);
and UO_1032 (O_1032,N_19600,N_19830);
nor UO_1033 (O_1033,N_19796,N_19759);
nand UO_1034 (O_1034,N_19877,N_19771);
nand UO_1035 (O_1035,N_19673,N_19729);
xor UO_1036 (O_1036,N_19740,N_19714);
nor UO_1037 (O_1037,N_19997,N_19814);
and UO_1038 (O_1038,N_19995,N_19713);
and UO_1039 (O_1039,N_19858,N_19869);
xnor UO_1040 (O_1040,N_19839,N_19788);
nor UO_1041 (O_1041,N_19906,N_19928);
and UO_1042 (O_1042,N_19672,N_19674);
xnor UO_1043 (O_1043,N_19941,N_19830);
or UO_1044 (O_1044,N_19965,N_19606);
nor UO_1045 (O_1045,N_19841,N_19768);
nand UO_1046 (O_1046,N_19628,N_19666);
or UO_1047 (O_1047,N_19625,N_19796);
nor UO_1048 (O_1048,N_19941,N_19900);
nor UO_1049 (O_1049,N_19655,N_19762);
nand UO_1050 (O_1050,N_19772,N_19924);
or UO_1051 (O_1051,N_19877,N_19655);
nor UO_1052 (O_1052,N_19893,N_19918);
nor UO_1053 (O_1053,N_19605,N_19882);
xor UO_1054 (O_1054,N_19912,N_19968);
and UO_1055 (O_1055,N_19991,N_19918);
and UO_1056 (O_1056,N_19946,N_19679);
nor UO_1057 (O_1057,N_19837,N_19736);
and UO_1058 (O_1058,N_19899,N_19829);
or UO_1059 (O_1059,N_19712,N_19860);
nor UO_1060 (O_1060,N_19632,N_19809);
nand UO_1061 (O_1061,N_19822,N_19721);
and UO_1062 (O_1062,N_19928,N_19797);
nor UO_1063 (O_1063,N_19928,N_19957);
nand UO_1064 (O_1064,N_19731,N_19850);
or UO_1065 (O_1065,N_19776,N_19621);
xor UO_1066 (O_1066,N_19724,N_19813);
nor UO_1067 (O_1067,N_19713,N_19663);
nand UO_1068 (O_1068,N_19639,N_19872);
xnor UO_1069 (O_1069,N_19761,N_19796);
and UO_1070 (O_1070,N_19992,N_19998);
xnor UO_1071 (O_1071,N_19749,N_19686);
nand UO_1072 (O_1072,N_19731,N_19867);
nand UO_1073 (O_1073,N_19786,N_19958);
and UO_1074 (O_1074,N_19777,N_19833);
or UO_1075 (O_1075,N_19708,N_19682);
or UO_1076 (O_1076,N_19987,N_19759);
nand UO_1077 (O_1077,N_19802,N_19604);
xnor UO_1078 (O_1078,N_19832,N_19733);
xnor UO_1079 (O_1079,N_19672,N_19876);
xor UO_1080 (O_1080,N_19626,N_19890);
or UO_1081 (O_1081,N_19975,N_19721);
nor UO_1082 (O_1082,N_19635,N_19910);
nor UO_1083 (O_1083,N_19660,N_19780);
nor UO_1084 (O_1084,N_19874,N_19809);
nand UO_1085 (O_1085,N_19728,N_19749);
nor UO_1086 (O_1086,N_19922,N_19643);
nand UO_1087 (O_1087,N_19615,N_19966);
or UO_1088 (O_1088,N_19676,N_19941);
xor UO_1089 (O_1089,N_19836,N_19780);
and UO_1090 (O_1090,N_19732,N_19691);
nand UO_1091 (O_1091,N_19965,N_19669);
nor UO_1092 (O_1092,N_19806,N_19934);
nand UO_1093 (O_1093,N_19707,N_19954);
nand UO_1094 (O_1094,N_19754,N_19776);
and UO_1095 (O_1095,N_19729,N_19824);
nor UO_1096 (O_1096,N_19796,N_19630);
nand UO_1097 (O_1097,N_19871,N_19739);
nor UO_1098 (O_1098,N_19974,N_19837);
nor UO_1099 (O_1099,N_19985,N_19877);
or UO_1100 (O_1100,N_19970,N_19810);
xnor UO_1101 (O_1101,N_19934,N_19999);
or UO_1102 (O_1102,N_19927,N_19973);
or UO_1103 (O_1103,N_19834,N_19941);
and UO_1104 (O_1104,N_19810,N_19693);
and UO_1105 (O_1105,N_19764,N_19828);
or UO_1106 (O_1106,N_19613,N_19741);
nor UO_1107 (O_1107,N_19746,N_19925);
nand UO_1108 (O_1108,N_19917,N_19908);
or UO_1109 (O_1109,N_19641,N_19778);
or UO_1110 (O_1110,N_19840,N_19713);
xor UO_1111 (O_1111,N_19919,N_19977);
or UO_1112 (O_1112,N_19607,N_19674);
xnor UO_1113 (O_1113,N_19665,N_19864);
nand UO_1114 (O_1114,N_19623,N_19645);
and UO_1115 (O_1115,N_19984,N_19790);
nand UO_1116 (O_1116,N_19655,N_19835);
or UO_1117 (O_1117,N_19977,N_19658);
nor UO_1118 (O_1118,N_19869,N_19615);
and UO_1119 (O_1119,N_19820,N_19897);
and UO_1120 (O_1120,N_19604,N_19741);
xor UO_1121 (O_1121,N_19837,N_19673);
and UO_1122 (O_1122,N_19878,N_19849);
nand UO_1123 (O_1123,N_19945,N_19738);
or UO_1124 (O_1124,N_19836,N_19990);
nand UO_1125 (O_1125,N_19943,N_19926);
xor UO_1126 (O_1126,N_19858,N_19769);
nor UO_1127 (O_1127,N_19636,N_19688);
or UO_1128 (O_1128,N_19897,N_19662);
or UO_1129 (O_1129,N_19900,N_19710);
xor UO_1130 (O_1130,N_19716,N_19898);
xor UO_1131 (O_1131,N_19899,N_19962);
nor UO_1132 (O_1132,N_19855,N_19792);
nor UO_1133 (O_1133,N_19652,N_19750);
or UO_1134 (O_1134,N_19659,N_19917);
xnor UO_1135 (O_1135,N_19671,N_19819);
or UO_1136 (O_1136,N_19753,N_19771);
nor UO_1137 (O_1137,N_19690,N_19610);
or UO_1138 (O_1138,N_19976,N_19816);
or UO_1139 (O_1139,N_19905,N_19874);
and UO_1140 (O_1140,N_19805,N_19640);
or UO_1141 (O_1141,N_19719,N_19888);
xor UO_1142 (O_1142,N_19695,N_19731);
nand UO_1143 (O_1143,N_19802,N_19777);
or UO_1144 (O_1144,N_19663,N_19684);
nand UO_1145 (O_1145,N_19693,N_19882);
nand UO_1146 (O_1146,N_19699,N_19789);
xor UO_1147 (O_1147,N_19685,N_19935);
and UO_1148 (O_1148,N_19731,N_19965);
nor UO_1149 (O_1149,N_19829,N_19621);
nand UO_1150 (O_1150,N_19969,N_19883);
xor UO_1151 (O_1151,N_19761,N_19668);
and UO_1152 (O_1152,N_19775,N_19833);
nand UO_1153 (O_1153,N_19656,N_19803);
nor UO_1154 (O_1154,N_19807,N_19753);
and UO_1155 (O_1155,N_19643,N_19835);
and UO_1156 (O_1156,N_19995,N_19968);
xnor UO_1157 (O_1157,N_19938,N_19867);
nand UO_1158 (O_1158,N_19882,N_19653);
nand UO_1159 (O_1159,N_19858,N_19963);
or UO_1160 (O_1160,N_19802,N_19911);
and UO_1161 (O_1161,N_19811,N_19770);
and UO_1162 (O_1162,N_19840,N_19712);
xor UO_1163 (O_1163,N_19654,N_19779);
and UO_1164 (O_1164,N_19928,N_19772);
nand UO_1165 (O_1165,N_19626,N_19985);
nor UO_1166 (O_1166,N_19738,N_19971);
xnor UO_1167 (O_1167,N_19993,N_19776);
nand UO_1168 (O_1168,N_19793,N_19695);
xnor UO_1169 (O_1169,N_19646,N_19609);
xnor UO_1170 (O_1170,N_19674,N_19635);
xor UO_1171 (O_1171,N_19657,N_19753);
or UO_1172 (O_1172,N_19828,N_19620);
nor UO_1173 (O_1173,N_19714,N_19674);
xor UO_1174 (O_1174,N_19702,N_19672);
or UO_1175 (O_1175,N_19875,N_19718);
nand UO_1176 (O_1176,N_19935,N_19864);
xnor UO_1177 (O_1177,N_19707,N_19647);
nor UO_1178 (O_1178,N_19830,N_19886);
nand UO_1179 (O_1179,N_19953,N_19685);
nor UO_1180 (O_1180,N_19915,N_19879);
xor UO_1181 (O_1181,N_19754,N_19770);
nor UO_1182 (O_1182,N_19791,N_19927);
and UO_1183 (O_1183,N_19723,N_19670);
or UO_1184 (O_1184,N_19770,N_19878);
nor UO_1185 (O_1185,N_19811,N_19807);
nand UO_1186 (O_1186,N_19706,N_19857);
or UO_1187 (O_1187,N_19948,N_19661);
and UO_1188 (O_1188,N_19922,N_19616);
xor UO_1189 (O_1189,N_19614,N_19955);
nand UO_1190 (O_1190,N_19628,N_19878);
nand UO_1191 (O_1191,N_19755,N_19700);
nand UO_1192 (O_1192,N_19968,N_19643);
xor UO_1193 (O_1193,N_19768,N_19831);
xnor UO_1194 (O_1194,N_19644,N_19717);
and UO_1195 (O_1195,N_19741,N_19998);
and UO_1196 (O_1196,N_19775,N_19993);
nor UO_1197 (O_1197,N_19835,N_19764);
xnor UO_1198 (O_1198,N_19889,N_19879);
nand UO_1199 (O_1199,N_19842,N_19792);
nor UO_1200 (O_1200,N_19931,N_19976);
nor UO_1201 (O_1201,N_19977,N_19767);
and UO_1202 (O_1202,N_19685,N_19887);
nand UO_1203 (O_1203,N_19768,N_19843);
nor UO_1204 (O_1204,N_19995,N_19769);
or UO_1205 (O_1205,N_19715,N_19901);
and UO_1206 (O_1206,N_19648,N_19864);
nand UO_1207 (O_1207,N_19685,N_19929);
nand UO_1208 (O_1208,N_19942,N_19855);
nand UO_1209 (O_1209,N_19935,N_19881);
xnor UO_1210 (O_1210,N_19992,N_19918);
nor UO_1211 (O_1211,N_19621,N_19611);
xor UO_1212 (O_1212,N_19991,N_19814);
and UO_1213 (O_1213,N_19712,N_19827);
or UO_1214 (O_1214,N_19739,N_19683);
and UO_1215 (O_1215,N_19695,N_19653);
nand UO_1216 (O_1216,N_19617,N_19748);
or UO_1217 (O_1217,N_19784,N_19850);
nor UO_1218 (O_1218,N_19982,N_19939);
nand UO_1219 (O_1219,N_19844,N_19739);
xor UO_1220 (O_1220,N_19656,N_19851);
nor UO_1221 (O_1221,N_19769,N_19693);
and UO_1222 (O_1222,N_19975,N_19895);
xnor UO_1223 (O_1223,N_19929,N_19829);
xnor UO_1224 (O_1224,N_19801,N_19828);
xor UO_1225 (O_1225,N_19906,N_19627);
and UO_1226 (O_1226,N_19692,N_19628);
and UO_1227 (O_1227,N_19976,N_19963);
and UO_1228 (O_1228,N_19915,N_19768);
and UO_1229 (O_1229,N_19613,N_19933);
and UO_1230 (O_1230,N_19846,N_19758);
xnor UO_1231 (O_1231,N_19697,N_19882);
xor UO_1232 (O_1232,N_19680,N_19702);
xor UO_1233 (O_1233,N_19725,N_19637);
xor UO_1234 (O_1234,N_19787,N_19788);
nor UO_1235 (O_1235,N_19705,N_19849);
nor UO_1236 (O_1236,N_19918,N_19710);
nand UO_1237 (O_1237,N_19983,N_19991);
or UO_1238 (O_1238,N_19934,N_19938);
nand UO_1239 (O_1239,N_19634,N_19946);
and UO_1240 (O_1240,N_19760,N_19703);
xor UO_1241 (O_1241,N_19947,N_19680);
nor UO_1242 (O_1242,N_19624,N_19640);
nand UO_1243 (O_1243,N_19805,N_19829);
and UO_1244 (O_1244,N_19924,N_19615);
xnor UO_1245 (O_1245,N_19872,N_19636);
and UO_1246 (O_1246,N_19686,N_19990);
nand UO_1247 (O_1247,N_19609,N_19759);
xor UO_1248 (O_1248,N_19992,N_19838);
and UO_1249 (O_1249,N_19806,N_19770);
or UO_1250 (O_1250,N_19608,N_19788);
xnor UO_1251 (O_1251,N_19685,N_19873);
and UO_1252 (O_1252,N_19639,N_19892);
xnor UO_1253 (O_1253,N_19824,N_19921);
and UO_1254 (O_1254,N_19657,N_19607);
nand UO_1255 (O_1255,N_19906,N_19987);
and UO_1256 (O_1256,N_19756,N_19736);
nor UO_1257 (O_1257,N_19966,N_19831);
nor UO_1258 (O_1258,N_19968,N_19627);
nand UO_1259 (O_1259,N_19747,N_19668);
and UO_1260 (O_1260,N_19608,N_19754);
nand UO_1261 (O_1261,N_19698,N_19881);
nand UO_1262 (O_1262,N_19658,N_19774);
or UO_1263 (O_1263,N_19760,N_19728);
or UO_1264 (O_1264,N_19921,N_19652);
and UO_1265 (O_1265,N_19957,N_19721);
xnor UO_1266 (O_1266,N_19838,N_19853);
nor UO_1267 (O_1267,N_19652,N_19671);
xor UO_1268 (O_1268,N_19805,N_19801);
nand UO_1269 (O_1269,N_19746,N_19921);
and UO_1270 (O_1270,N_19988,N_19746);
or UO_1271 (O_1271,N_19927,N_19707);
xor UO_1272 (O_1272,N_19934,N_19639);
nor UO_1273 (O_1273,N_19928,N_19884);
and UO_1274 (O_1274,N_19780,N_19851);
and UO_1275 (O_1275,N_19993,N_19722);
and UO_1276 (O_1276,N_19956,N_19608);
xnor UO_1277 (O_1277,N_19984,N_19648);
or UO_1278 (O_1278,N_19778,N_19748);
or UO_1279 (O_1279,N_19719,N_19966);
or UO_1280 (O_1280,N_19898,N_19886);
nor UO_1281 (O_1281,N_19929,N_19670);
and UO_1282 (O_1282,N_19734,N_19696);
nor UO_1283 (O_1283,N_19975,N_19630);
xor UO_1284 (O_1284,N_19959,N_19971);
and UO_1285 (O_1285,N_19827,N_19840);
nand UO_1286 (O_1286,N_19784,N_19986);
or UO_1287 (O_1287,N_19868,N_19780);
nor UO_1288 (O_1288,N_19784,N_19834);
nand UO_1289 (O_1289,N_19801,N_19724);
and UO_1290 (O_1290,N_19692,N_19983);
xor UO_1291 (O_1291,N_19825,N_19829);
nor UO_1292 (O_1292,N_19975,N_19723);
xor UO_1293 (O_1293,N_19649,N_19760);
xor UO_1294 (O_1294,N_19663,N_19912);
nor UO_1295 (O_1295,N_19945,N_19712);
and UO_1296 (O_1296,N_19665,N_19653);
or UO_1297 (O_1297,N_19881,N_19961);
nor UO_1298 (O_1298,N_19610,N_19746);
xnor UO_1299 (O_1299,N_19774,N_19905);
and UO_1300 (O_1300,N_19761,N_19785);
or UO_1301 (O_1301,N_19647,N_19892);
xnor UO_1302 (O_1302,N_19855,N_19630);
and UO_1303 (O_1303,N_19605,N_19988);
xnor UO_1304 (O_1304,N_19968,N_19796);
xor UO_1305 (O_1305,N_19752,N_19694);
or UO_1306 (O_1306,N_19752,N_19976);
xor UO_1307 (O_1307,N_19877,N_19872);
nor UO_1308 (O_1308,N_19871,N_19732);
or UO_1309 (O_1309,N_19865,N_19682);
and UO_1310 (O_1310,N_19696,N_19993);
nand UO_1311 (O_1311,N_19779,N_19900);
or UO_1312 (O_1312,N_19651,N_19652);
nand UO_1313 (O_1313,N_19887,N_19659);
or UO_1314 (O_1314,N_19858,N_19995);
and UO_1315 (O_1315,N_19705,N_19989);
nor UO_1316 (O_1316,N_19719,N_19613);
or UO_1317 (O_1317,N_19961,N_19891);
or UO_1318 (O_1318,N_19830,N_19679);
nand UO_1319 (O_1319,N_19840,N_19878);
nand UO_1320 (O_1320,N_19680,N_19674);
xnor UO_1321 (O_1321,N_19814,N_19704);
nand UO_1322 (O_1322,N_19893,N_19666);
xnor UO_1323 (O_1323,N_19664,N_19911);
or UO_1324 (O_1324,N_19831,N_19973);
nor UO_1325 (O_1325,N_19624,N_19827);
or UO_1326 (O_1326,N_19787,N_19847);
xnor UO_1327 (O_1327,N_19758,N_19706);
or UO_1328 (O_1328,N_19608,N_19850);
xor UO_1329 (O_1329,N_19762,N_19626);
and UO_1330 (O_1330,N_19864,N_19622);
nand UO_1331 (O_1331,N_19785,N_19997);
or UO_1332 (O_1332,N_19788,N_19942);
or UO_1333 (O_1333,N_19681,N_19734);
nor UO_1334 (O_1334,N_19755,N_19817);
and UO_1335 (O_1335,N_19946,N_19863);
nand UO_1336 (O_1336,N_19868,N_19718);
xnor UO_1337 (O_1337,N_19874,N_19715);
and UO_1338 (O_1338,N_19666,N_19931);
and UO_1339 (O_1339,N_19792,N_19673);
xor UO_1340 (O_1340,N_19669,N_19731);
nand UO_1341 (O_1341,N_19814,N_19688);
and UO_1342 (O_1342,N_19937,N_19860);
nand UO_1343 (O_1343,N_19619,N_19818);
xor UO_1344 (O_1344,N_19740,N_19870);
xor UO_1345 (O_1345,N_19947,N_19823);
or UO_1346 (O_1346,N_19882,N_19860);
xor UO_1347 (O_1347,N_19666,N_19847);
xnor UO_1348 (O_1348,N_19974,N_19607);
or UO_1349 (O_1349,N_19859,N_19833);
and UO_1350 (O_1350,N_19940,N_19677);
xor UO_1351 (O_1351,N_19676,N_19779);
nand UO_1352 (O_1352,N_19744,N_19706);
or UO_1353 (O_1353,N_19785,N_19851);
nand UO_1354 (O_1354,N_19718,N_19805);
and UO_1355 (O_1355,N_19636,N_19997);
nor UO_1356 (O_1356,N_19927,N_19964);
or UO_1357 (O_1357,N_19933,N_19934);
or UO_1358 (O_1358,N_19717,N_19761);
xor UO_1359 (O_1359,N_19889,N_19790);
and UO_1360 (O_1360,N_19816,N_19746);
or UO_1361 (O_1361,N_19844,N_19980);
or UO_1362 (O_1362,N_19722,N_19854);
or UO_1363 (O_1363,N_19616,N_19667);
nand UO_1364 (O_1364,N_19996,N_19795);
nand UO_1365 (O_1365,N_19923,N_19658);
xnor UO_1366 (O_1366,N_19800,N_19746);
or UO_1367 (O_1367,N_19846,N_19956);
nand UO_1368 (O_1368,N_19783,N_19772);
nor UO_1369 (O_1369,N_19857,N_19922);
xnor UO_1370 (O_1370,N_19610,N_19662);
or UO_1371 (O_1371,N_19695,N_19685);
xor UO_1372 (O_1372,N_19617,N_19869);
nand UO_1373 (O_1373,N_19968,N_19987);
nand UO_1374 (O_1374,N_19711,N_19812);
xor UO_1375 (O_1375,N_19728,N_19792);
or UO_1376 (O_1376,N_19888,N_19840);
or UO_1377 (O_1377,N_19649,N_19655);
or UO_1378 (O_1378,N_19796,N_19720);
nor UO_1379 (O_1379,N_19958,N_19671);
and UO_1380 (O_1380,N_19616,N_19764);
or UO_1381 (O_1381,N_19890,N_19998);
xnor UO_1382 (O_1382,N_19955,N_19692);
xor UO_1383 (O_1383,N_19720,N_19736);
and UO_1384 (O_1384,N_19893,N_19713);
and UO_1385 (O_1385,N_19624,N_19608);
xor UO_1386 (O_1386,N_19802,N_19728);
nand UO_1387 (O_1387,N_19800,N_19772);
and UO_1388 (O_1388,N_19853,N_19966);
nor UO_1389 (O_1389,N_19856,N_19801);
nand UO_1390 (O_1390,N_19895,N_19727);
or UO_1391 (O_1391,N_19720,N_19821);
nand UO_1392 (O_1392,N_19636,N_19813);
and UO_1393 (O_1393,N_19659,N_19739);
or UO_1394 (O_1394,N_19921,N_19822);
xnor UO_1395 (O_1395,N_19877,N_19677);
xor UO_1396 (O_1396,N_19948,N_19964);
and UO_1397 (O_1397,N_19632,N_19729);
nand UO_1398 (O_1398,N_19622,N_19863);
and UO_1399 (O_1399,N_19932,N_19791);
or UO_1400 (O_1400,N_19956,N_19863);
nand UO_1401 (O_1401,N_19729,N_19788);
and UO_1402 (O_1402,N_19863,N_19679);
nor UO_1403 (O_1403,N_19686,N_19790);
nor UO_1404 (O_1404,N_19752,N_19755);
and UO_1405 (O_1405,N_19721,N_19689);
and UO_1406 (O_1406,N_19962,N_19789);
nand UO_1407 (O_1407,N_19918,N_19763);
nor UO_1408 (O_1408,N_19773,N_19832);
xor UO_1409 (O_1409,N_19677,N_19721);
nor UO_1410 (O_1410,N_19937,N_19732);
xnor UO_1411 (O_1411,N_19844,N_19896);
or UO_1412 (O_1412,N_19674,N_19611);
nor UO_1413 (O_1413,N_19783,N_19778);
nor UO_1414 (O_1414,N_19840,N_19776);
xnor UO_1415 (O_1415,N_19726,N_19802);
xor UO_1416 (O_1416,N_19992,N_19850);
and UO_1417 (O_1417,N_19639,N_19690);
nand UO_1418 (O_1418,N_19943,N_19682);
nand UO_1419 (O_1419,N_19647,N_19743);
nand UO_1420 (O_1420,N_19841,N_19924);
or UO_1421 (O_1421,N_19825,N_19656);
nor UO_1422 (O_1422,N_19984,N_19772);
nand UO_1423 (O_1423,N_19611,N_19754);
xnor UO_1424 (O_1424,N_19888,N_19857);
or UO_1425 (O_1425,N_19963,N_19886);
nand UO_1426 (O_1426,N_19950,N_19946);
or UO_1427 (O_1427,N_19890,N_19975);
xor UO_1428 (O_1428,N_19981,N_19989);
nand UO_1429 (O_1429,N_19917,N_19764);
or UO_1430 (O_1430,N_19606,N_19644);
xnor UO_1431 (O_1431,N_19989,N_19861);
and UO_1432 (O_1432,N_19644,N_19665);
nand UO_1433 (O_1433,N_19754,N_19993);
or UO_1434 (O_1434,N_19630,N_19794);
xor UO_1435 (O_1435,N_19668,N_19846);
and UO_1436 (O_1436,N_19754,N_19647);
and UO_1437 (O_1437,N_19793,N_19871);
and UO_1438 (O_1438,N_19879,N_19623);
xnor UO_1439 (O_1439,N_19740,N_19792);
and UO_1440 (O_1440,N_19784,N_19644);
nand UO_1441 (O_1441,N_19864,N_19645);
or UO_1442 (O_1442,N_19618,N_19663);
nor UO_1443 (O_1443,N_19886,N_19879);
xor UO_1444 (O_1444,N_19611,N_19903);
nor UO_1445 (O_1445,N_19659,N_19888);
nor UO_1446 (O_1446,N_19942,N_19785);
nand UO_1447 (O_1447,N_19676,N_19730);
nor UO_1448 (O_1448,N_19735,N_19674);
nor UO_1449 (O_1449,N_19840,N_19761);
nand UO_1450 (O_1450,N_19833,N_19849);
nand UO_1451 (O_1451,N_19916,N_19664);
and UO_1452 (O_1452,N_19779,N_19758);
or UO_1453 (O_1453,N_19793,N_19849);
nor UO_1454 (O_1454,N_19852,N_19685);
nor UO_1455 (O_1455,N_19676,N_19902);
nor UO_1456 (O_1456,N_19987,N_19966);
nand UO_1457 (O_1457,N_19754,N_19798);
nor UO_1458 (O_1458,N_19850,N_19748);
and UO_1459 (O_1459,N_19706,N_19796);
and UO_1460 (O_1460,N_19829,N_19704);
xnor UO_1461 (O_1461,N_19733,N_19953);
xor UO_1462 (O_1462,N_19998,N_19975);
or UO_1463 (O_1463,N_19623,N_19705);
xnor UO_1464 (O_1464,N_19806,N_19783);
or UO_1465 (O_1465,N_19640,N_19736);
and UO_1466 (O_1466,N_19915,N_19939);
nand UO_1467 (O_1467,N_19940,N_19631);
or UO_1468 (O_1468,N_19909,N_19647);
xor UO_1469 (O_1469,N_19693,N_19772);
or UO_1470 (O_1470,N_19804,N_19929);
or UO_1471 (O_1471,N_19826,N_19837);
nand UO_1472 (O_1472,N_19932,N_19713);
or UO_1473 (O_1473,N_19688,N_19676);
nor UO_1474 (O_1474,N_19962,N_19812);
xnor UO_1475 (O_1475,N_19627,N_19772);
nand UO_1476 (O_1476,N_19849,N_19681);
xor UO_1477 (O_1477,N_19870,N_19996);
nand UO_1478 (O_1478,N_19780,N_19635);
or UO_1479 (O_1479,N_19668,N_19666);
nor UO_1480 (O_1480,N_19807,N_19910);
nor UO_1481 (O_1481,N_19845,N_19902);
nor UO_1482 (O_1482,N_19839,N_19947);
and UO_1483 (O_1483,N_19958,N_19678);
nor UO_1484 (O_1484,N_19873,N_19860);
and UO_1485 (O_1485,N_19650,N_19700);
or UO_1486 (O_1486,N_19969,N_19956);
and UO_1487 (O_1487,N_19855,N_19901);
and UO_1488 (O_1488,N_19836,N_19882);
nand UO_1489 (O_1489,N_19654,N_19706);
and UO_1490 (O_1490,N_19845,N_19803);
nand UO_1491 (O_1491,N_19944,N_19705);
or UO_1492 (O_1492,N_19681,N_19728);
nand UO_1493 (O_1493,N_19704,N_19677);
or UO_1494 (O_1494,N_19731,N_19745);
nand UO_1495 (O_1495,N_19846,N_19932);
nor UO_1496 (O_1496,N_19988,N_19688);
or UO_1497 (O_1497,N_19974,N_19956);
xor UO_1498 (O_1498,N_19970,N_19689);
or UO_1499 (O_1499,N_19922,N_19762);
nand UO_1500 (O_1500,N_19868,N_19751);
xor UO_1501 (O_1501,N_19729,N_19900);
nand UO_1502 (O_1502,N_19602,N_19850);
and UO_1503 (O_1503,N_19888,N_19925);
nor UO_1504 (O_1504,N_19669,N_19764);
or UO_1505 (O_1505,N_19695,N_19746);
xor UO_1506 (O_1506,N_19641,N_19634);
and UO_1507 (O_1507,N_19716,N_19747);
xnor UO_1508 (O_1508,N_19855,N_19917);
xor UO_1509 (O_1509,N_19842,N_19762);
nand UO_1510 (O_1510,N_19653,N_19951);
xor UO_1511 (O_1511,N_19964,N_19628);
and UO_1512 (O_1512,N_19820,N_19871);
xor UO_1513 (O_1513,N_19864,N_19859);
nor UO_1514 (O_1514,N_19894,N_19665);
and UO_1515 (O_1515,N_19633,N_19640);
or UO_1516 (O_1516,N_19912,N_19696);
xnor UO_1517 (O_1517,N_19794,N_19798);
nor UO_1518 (O_1518,N_19625,N_19988);
and UO_1519 (O_1519,N_19903,N_19608);
nand UO_1520 (O_1520,N_19862,N_19653);
and UO_1521 (O_1521,N_19754,N_19758);
xnor UO_1522 (O_1522,N_19936,N_19642);
nand UO_1523 (O_1523,N_19600,N_19962);
or UO_1524 (O_1524,N_19659,N_19652);
nor UO_1525 (O_1525,N_19921,N_19795);
or UO_1526 (O_1526,N_19827,N_19804);
nand UO_1527 (O_1527,N_19605,N_19649);
nand UO_1528 (O_1528,N_19728,N_19933);
nor UO_1529 (O_1529,N_19733,N_19751);
nor UO_1530 (O_1530,N_19617,N_19815);
or UO_1531 (O_1531,N_19958,N_19956);
nand UO_1532 (O_1532,N_19683,N_19982);
or UO_1533 (O_1533,N_19976,N_19949);
and UO_1534 (O_1534,N_19894,N_19899);
and UO_1535 (O_1535,N_19882,N_19955);
nand UO_1536 (O_1536,N_19988,N_19732);
and UO_1537 (O_1537,N_19631,N_19992);
or UO_1538 (O_1538,N_19697,N_19982);
and UO_1539 (O_1539,N_19936,N_19606);
and UO_1540 (O_1540,N_19850,N_19655);
xor UO_1541 (O_1541,N_19659,N_19992);
nor UO_1542 (O_1542,N_19931,N_19886);
and UO_1543 (O_1543,N_19792,N_19659);
xnor UO_1544 (O_1544,N_19775,N_19616);
nand UO_1545 (O_1545,N_19996,N_19925);
or UO_1546 (O_1546,N_19634,N_19972);
or UO_1547 (O_1547,N_19884,N_19803);
and UO_1548 (O_1548,N_19601,N_19733);
xor UO_1549 (O_1549,N_19767,N_19972);
nand UO_1550 (O_1550,N_19953,N_19898);
or UO_1551 (O_1551,N_19898,N_19933);
or UO_1552 (O_1552,N_19921,N_19605);
xor UO_1553 (O_1553,N_19730,N_19939);
nor UO_1554 (O_1554,N_19671,N_19678);
nor UO_1555 (O_1555,N_19625,N_19851);
or UO_1556 (O_1556,N_19892,N_19635);
nor UO_1557 (O_1557,N_19894,N_19924);
and UO_1558 (O_1558,N_19736,N_19905);
and UO_1559 (O_1559,N_19842,N_19824);
or UO_1560 (O_1560,N_19856,N_19810);
nor UO_1561 (O_1561,N_19752,N_19690);
xnor UO_1562 (O_1562,N_19671,N_19951);
xor UO_1563 (O_1563,N_19879,N_19666);
or UO_1564 (O_1564,N_19759,N_19700);
nor UO_1565 (O_1565,N_19901,N_19695);
or UO_1566 (O_1566,N_19837,N_19780);
nand UO_1567 (O_1567,N_19937,N_19640);
xor UO_1568 (O_1568,N_19961,N_19807);
nand UO_1569 (O_1569,N_19747,N_19835);
xnor UO_1570 (O_1570,N_19861,N_19857);
nor UO_1571 (O_1571,N_19734,N_19634);
nor UO_1572 (O_1572,N_19739,N_19929);
nor UO_1573 (O_1573,N_19912,N_19779);
nor UO_1574 (O_1574,N_19656,N_19720);
and UO_1575 (O_1575,N_19648,N_19680);
nor UO_1576 (O_1576,N_19840,N_19785);
nor UO_1577 (O_1577,N_19965,N_19690);
xnor UO_1578 (O_1578,N_19902,N_19816);
and UO_1579 (O_1579,N_19854,N_19955);
and UO_1580 (O_1580,N_19769,N_19694);
or UO_1581 (O_1581,N_19785,N_19691);
xnor UO_1582 (O_1582,N_19734,N_19768);
or UO_1583 (O_1583,N_19936,N_19952);
and UO_1584 (O_1584,N_19734,N_19828);
nand UO_1585 (O_1585,N_19974,N_19830);
xor UO_1586 (O_1586,N_19980,N_19772);
xnor UO_1587 (O_1587,N_19938,N_19992);
xnor UO_1588 (O_1588,N_19964,N_19986);
xor UO_1589 (O_1589,N_19657,N_19761);
and UO_1590 (O_1590,N_19870,N_19808);
nand UO_1591 (O_1591,N_19605,N_19977);
nand UO_1592 (O_1592,N_19988,N_19702);
xor UO_1593 (O_1593,N_19608,N_19826);
nand UO_1594 (O_1594,N_19637,N_19885);
xor UO_1595 (O_1595,N_19963,N_19725);
nor UO_1596 (O_1596,N_19986,N_19687);
and UO_1597 (O_1597,N_19952,N_19835);
nor UO_1598 (O_1598,N_19758,N_19654);
nor UO_1599 (O_1599,N_19661,N_19982);
and UO_1600 (O_1600,N_19891,N_19657);
xnor UO_1601 (O_1601,N_19628,N_19611);
nor UO_1602 (O_1602,N_19724,N_19993);
and UO_1603 (O_1603,N_19894,N_19702);
nand UO_1604 (O_1604,N_19955,N_19713);
nand UO_1605 (O_1605,N_19888,N_19781);
nand UO_1606 (O_1606,N_19771,N_19950);
and UO_1607 (O_1607,N_19654,N_19854);
xnor UO_1608 (O_1608,N_19711,N_19700);
and UO_1609 (O_1609,N_19856,N_19842);
and UO_1610 (O_1610,N_19789,N_19619);
xnor UO_1611 (O_1611,N_19835,N_19786);
and UO_1612 (O_1612,N_19818,N_19906);
nand UO_1613 (O_1613,N_19736,N_19710);
and UO_1614 (O_1614,N_19951,N_19776);
xor UO_1615 (O_1615,N_19767,N_19718);
xnor UO_1616 (O_1616,N_19668,N_19842);
nand UO_1617 (O_1617,N_19916,N_19768);
and UO_1618 (O_1618,N_19726,N_19954);
nand UO_1619 (O_1619,N_19735,N_19857);
xor UO_1620 (O_1620,N_19910,N_19687);
nor UO_1621 (O_1621,N_19826,N_19811);
or UO_1622 (O_1622,N_19766,N_19904);
nor UO_1623 (O_1623,N_19843,N_19782);
nand UO_1624 (O_1624,N_19842,N_19664);
or UO_1625 (O_1625,N_19855,N_19922);
and UO_1626 (O_1626,N_19826,N_19648);
xnor UO_1627 (O_1627,N_19738,N_19910);
and UO_1628 (O_1628,N_19858,N_19977);
xor UO_1629 (O_1629,N_19964,N_19682);
nand UO_1630 (O_1630,N_19689,N_19704);
nand UO_1631 (O_1631,N_19686,N_19714);
nor UO_1632 (O_1632,N_19857,N_19707);
nand UO_1633 (O_1633,N_19621,N_19784);
nand UO_1634 (O_1634,N_19882,N_19863);
nor UO_1635 (O_1635,N_19954,N_19677);
xnor UO_1636 (O_1636,N_19841,N_19785);
and UO_1637 (O_1637,N_19716,N_19822);
and UO_1638 (O_1638,N_19606,N_19788);
or UO_1639 (O_1639,N_19918,N_19609);
nor UO_1640 (O_1640,N_19785,N_19632);
nand UO_1641 (O_1641,N_19747,N_19662);
nand UO_1642 (O_1642,N_19700,N_19837);
xor UO_1643 (O_1643,N_19625,N_19724);
and UO_1644 (O_1644,N_19930,N_19750);
and UO_1645 (O_1645,N_19726,N_19789);
and UO_1646 (O_1646,N_19890,N_19957);
xor UO_1647 (O_1647,N_19931,N_19850);
nand UO_1648 (O_1648,N_19775,N_19753);
or UO_1649 (O_1649,N_19904,N_19836);
or UO_1650 (O_1650,N_19874,N_19843);
and UO_1651 (O_1651,N_19925,N_19601);
xor UO_1652 (O_1652,N_19901,N_19835);
xnor UO_1653 (O_1653,N_19621,N_19975);
nand UO_1654 (O_1654,N_19705,N_19857);
xnor UO_1655 (O_1655,N_19641,N_19822);
nand UO_1656 (O_1656,N_19995,N_19604);
or UO_1657 (O_1657,N_19822,N_19872);
nand UO_1658 (O_1658,N_19814,N_19961);
xor UO_1659 (O_1659,N_19654,N_19979);
and UO_1660 (O_1660,N_19824,N_19922);
xor UO_1661 (O_1661,N_19899,N_19691);
nand UO_1662 (O_1662,N_19888,N_19953);
and UO_1663 (O_1663,N_19989,N_19820);
nor UO_1664 (O_1664,N_19873,N_19716);
and UO_1665 (O_1665,N_19767,N_19830);
nand UO_1666 (O_1666,N_19710,N_19997);
xor UO_1667 (O_1667,N_19813,N_19903);
nor UO_1668 (O_1668,N_19774,N_19692);
nand UO_1669 (O_1669,N_19791,N_19800);
xnor UO_1670 (O_1670,N_19945,N_19868);
nor UO_1671 (O_1671,N_19778,N_19959);
xor UO_1672 (O_1672,N_19647,N_19752);
nor UO_1673 (O_1673,N_19703,N_19624);
nor UO_1674 (O_1674,N_19819,N_19642);
xnor UO_1675 (O_1675,N_19763,N_19841);
nand UO_1676 (O_1676,N_19647,N_19938);
and UO_1677 (O_1677,N_19681,N_19692);
nand UO_1678 (O_1678,N_19662,N_19893);
nand UO_1679 (O_1679,N_19982,N_19787);
nor UO_1680 (O_1680,N_19726,N_19930);
xnor UO_1681 (O_1681,N_19667,N_19654);
and UO_1682 (O_1682,N_19755,N_19783);
nand UO_1683 (O_1683,N_19632,N_19904);
nor UO_1684 (O_1684,N_19611,N_19892);
xor UO_1685 (O_1685,N_19940,N_19911);
nor UO_1686 (O_1686,N_19758,N_19659);
and UO_1687 (O_1687,N_19743,N_19612);
xor UO_1688 (O_1688,N_19984,N_19601);
or UO_1689 (O_1689,N_19906,N_19826);
or UO_1690 (O_1690,N_19927,N_19720);
nor UO_1691 (O_1691,N_19876,N_19778);
nor UO_1692 (O_1692,N_19701,N_19954);
nand UO_1693 (O_1693,N_19703,N_19871);
and UO_1694 (O_1694,N_19946,N_19928);
nand UO_1695 (O_1695,N_19813,N_19999);
xnor UO_1696 (O_1696,N_19839,N_19956);
nand UO_1697 (O_1697,N_19713,N_19712);
and UO_1698 (O_1698,N_19644,N_19797);
xor UO_1699 (O_1699,N_19625,N_19896);
or UO_1700 (O_1700,N_19798,N_19988);
xnor UO_1701 (O_1701,N_19686,N_19694);
or UO_1702 (O_1702,N_19802,N_19753);
nand UO_1703 (O_1703,N_19694,N_19863);
or UO_1704 (O_1704,N_19970,N_19756);
and UO_1705 (O_1705,N_19711,N_19603);
nand UO_1706 (O_1706,N_19713,N_19629);
nand UO_1707 (O_1707,N_19772,N_19939);
nand UO_1708 (O_1708,N_19629,N_19826);
nand UO_1709 (O_1709,N_19926,N_19639);
nor UO_1710 (O_1710,N_19947,N_19889);
xor UO_1711 (O_1711,N_19756,N_19635);
and UO_1712 (O_1712,N_19731,N_19664);
nor UO_1713 (O_1713,N_19967,N_19958);
nand UO_1714 (O_1714,N_19882,N_19812);
nor UO_1715 (O_1715,N_19944,N_19725);
and UO_1716 (O_1716,N_19867,N_19709);
xnor UO_1717 (O_1717,N_19674,N_19965);
xor UO_1718 (O_1718,N_19769,N_19880);
nor UO_1719 (O_1719,N_19831,N_19805);
xor UO_1720 (O_1720,N_19837,N_19794);
nor UO_1721 (O_1721,N_19814,N_19747);
nand UO_1722 (O_1722,N_19750,N_19974);
and UO_1723 (O_1723,N_19997,N_19794);
xor UO_1724 (O_1724,N_19870,N_19687);
nor UO_1725 (O_1725,N_19637,N_19858);
nor UO_1726 (O_1726,N_19658,N_19684);
xnor UO_1727 (O_1727,N_19651,N_19619);
nor UO_1728 (O_1728,N_19751,N_19861);
and UO_1729 (O_1729,N_19696,N_19739);
or UO_1730 (O_1730,N_19857,N_19678);
xnor UO_1731 (O_1731,N_19973,N_19930);
and UO_1732 (O_1732,N_19856,N_19907);
nand UO_1733 (O_1733,N_19982,N_19666);
xor UO_1734 (O_1734,N_19690,N_19982);
nand UO_1735 (O_1735,N_19859,N_19909);
nor UO_1736 (O_1736,N_19835,N_19668);
or UO_1737 (O_1737,N_19786,N_19929);
nand UO_1738 (O_1738,N_19816,N_19813);
and UO_1739 (O_1739,N_19836,N_19686);
or UO_1740 (O_1740,N_19655,N_19887);
nand UO_1741 (O_1741,N_19991,N_19623);
nor UO_1742 (O_1742,N_19791,N_19899);
or UO_1743 (O_1743,N_19998,N_19902);
nor UO_1744 (O_1744,N_19602,N_19773);
xnor UO_1745 (O_1745,N_19853,N_19740);
nor UO_1746 (O_1746,N_19745,N_19987);
nor UO_1747 (O_1747,N_19754,N_19970);
and UO_1748 (O_1748,N_19939,N_19685);
and UO_1749 (O_1749,N_19777,N_19621);
and UO_1750 (O_1750,N_19992,N_19625);
xnor UO_1751 (O_1751,N_19850,N_19997);
xnor UO_1752 (O_1752,N_19970,N_19980);
nor UO_1753 (O_1753,N_19976,N_19829);
or UO_1754 (O_1754,N_19990,N_19886);
nand UO_1755 (O_1755,N_19953,N_19630);
nor UO_1756 (O_1756,N_19684,N_19639);
nor UO_1757 (O_1757,N_19831,N_19843);
and UO_1758 (O_1758,N_19672,N_19851);
or UO_1759 (O_1759,N_19813,N_19614);
or UO_1760 (O_1760,N_19964,N_19685);
nand UO_1761 (O_1761,N_19620,N_19732);
and UO_1762 (O_1762,N_19673,N_19725);
nand UO_1763 (O_1763,N_19761,N_19979);
or UO_1764 (O_1764,N_19800,N_19948);
xnor UO_1765 (O_1765,N_19608,N_19978);
and UO_1766 (O_1766,N_19753,N_19945);
and UO_1767 (O_1767,N_19902,N_19932);
or UO_1768 (O_1768,N_19957,N_19756);
or UO_1769 (O_1769,N_19953,N_19673);
xnor UO_1770 (O_1770,N_19935,N_19931);
nor UO_1771 (O_1771,N_19861,N_19722);
nor UO_1772 (O_1772,N_19675,N_19987);
nor UO_1773 (O_1773,N_19680,N_19979);
nor UO_1774 (O_1774,N_19938,N_19886);
nand UO_1775 (O_1775,N_19855,N_19991);
or UO_1776 (O_1776,N_19751,N_19737);
and UO_1777 (O_1777,N_19899,N_19910);
and UO_1778 (O_1778,N_19985,N_19874);
and UO_1779 (O_1779,N_19732,N_19995);
xnor UO_1780 (O_1780,N_19637,N_19852);
xor UO_1781 (O_1781,N_19759,N_19729);
xor UO_1782 (O_1782,N_19941,N_19665);
nor UO_1783 (O_1783,N_19624,N_19616);
nand UO_1784 (O_1784,N_19714,N_19769);
nand UO_1785 (O_1785,N_19944,N_19759);
nand UO_1786 (O_1786,N_19639,N_19792);
or UO_1787 (O_1787,N_19918,N_19897);
nor UO_1788 (O_1788,N_19606,N_19747);
nand UO_1789 (O_1789,N_19613,N_19944);
or UO_1790 (O_1790,N_19657,N_19663);
or UO_1791 (O_1791,N_19690,N_19705);
nor UO_1792 (O_1792,N_19658,N_19879);
or UO_1793 (O_1793,N_19966,N_19847);
or UO_1794 (O_1794,N_19916,N_19639);
nand UO_1795 (O_1795,N_19887,N_19632);
nand UO_1796 (O_1796,N_19823,N_19891);
or UO_1797 (O_1797,N_19895,N_19898);
xnor UO_1798 (O_1798,N_19909,N_19870);
nor UO_1799 (O_1799,N_19772,N_19764);
nand UO_1800 (O_1800,N_19960,N_19849);
nand UO_1801 (O_1801,N_19893,N_19978);
and UO_1802 (O_1802,N_19979,N_19899);
nor UO_1803 (O_1803,N_19752,N_19781);
xnor UO_1804 (O_1804,N_19647,N_19763);
or UO_1805 (O_1805,N_19760,N_19650);
nor UO_1806 (O_1806,N_19879,N_19917);
nor UO_1807 (O_1807,N_19902,N_19893);
and UO_1808 (O_1808,N_19856,N_19768);
and UO_1809 (O_1809,N_19814,N_19803);
nand UO_1810 (O_1810,N_19677,N_19915);
nor UO_1811 (O_1811,N_19876,N_19895);
xor UO_1812 (O_1812,N_19789,N_19727);
and UO_1813 (O_1813,N_19971,N_19722);
or UO_1814 (O_1814,N_19756,N_19788);
or UO_1815 (O_1815,N_19986,N_19698);
xnor UO_1816 (O_1816,N_19980,N_19723);
xor UO_1817 (O_1817,N_19820,N_19746);
nand UO_1818 (O_1818,N_19742,N_19995);
xnor UO_1819 (O_1819,N_19838,N_19650);
nand UO_1820 (O_1820,N_19600,N_19927);
or UO_1821 (O_1821,N_19866,N_19893);
or UO_1822 (O_1822,N_19994,N_19810);
xnor UO_1823 (O_1823,N_19790,N_19796);
or UO_1824 (O_1824,N_19778,N_19954);
xor UO_1825 (O_1825,N_19962,N_19771);
or UO_1826 (O_1826,N_19814,N_19685);
xor UO_1827 (O_1827,N_19943,N_19959);
xor UO_1828 (O_1828,N_19715,N_19982);
or UO_1829 (O_1829,N_19898,N_19843);
nand UO_1830 (O_1830,N_19641,N_19635);
or UO_1831 (O_1831,N_19612,N_19779);
and UO_1832 (O_1832,N_19861,N_19830);
nor UO_1833 (O_1833,N_19733,N_19895);
or UO_1834 (O_1834,N_19689,N_19634);
nor UO_1835 (O_1835,N_19787,N_19732);
and UO_1836 (O_1836,N_19722,N_19868);
nor UO_1837 (O_1837,N_19631,N_19971);
xor UO_1838 (O_1838,N_19911,N_19796);
and UO_1839 (O_1839,N_19619,N_19837);
or UO_1840 (O_1840,N_19935,N_19677);
and UO_1841 (O_1841,N_19851,N_19837);
or UO_1842 (O_1842,N_19674,N_19828);
nor UO_1843 (O_1843,N_19707,N_19831);
xor UO_1844 (O_1844,N_19893,N_19669);
xnor UO_1845 (O_1845,N_19840,N_19871);
nor UO_1846 (O_1846,N_19988,N_19907);
nand UO_1847 (O_1847,N_19707,N_19694);
xnor UO_1848 (O_1848,N_19997,N_19622);
nor UO_1849 (O_1849,N_19729,N_19936);
nand UO_1850 (O_1850,N_19816,N_19909);
or UO_1851 (O_1851,N_19959,N_19721);
nor UO_1852 (O_1852,N_19714,N_19689);
and UO_1853 (O_1853,N_19814,N_19875);
or UO_1854 (O_1854,N_19692,N_19673);
and UO_1855 (O_1855,N_19881,N_19744);
xnor UO_1856 (O_1856,N_19662,N_19668);
and UO_1857 (O_1857,N_19723,N_19754);
or UO_1858 (O_1858,N_19708,N_19668);
and UO_1859 (O_1859,N_19905,N_19910);
and UO_1860 (O_1860,N_19825,N_19735);
nor UO_1861 (O_1861,N_19956,N_19835);
nor UO_1862 (O_1862,N_19950,N_19733);
xnor UO_1863 (O_1863,N_19711,N_19975);
and UO_1864 (O_1864,N_19717,N_19804);
and UO_1865 (O_1865,N_19950,N_19893);
or UO_1866 (O_1866,N_19909,N_19994);
nor UO_1867 (O_1867,N_19989,N_19865);
xnor UO_1868 (O_1868,N_19761,N_19954);
nand UO_1869 (O_1869,N_19796,N_19805);
or UO_1870 (O_1870,N_19942,N_19611);
and UO_1871 (O_1871,N_19962,N_19852);
nor UO_1872 (O_1872,N_19919,N_19744);
or UO_1873 (O_1873,N_19721,N_19826);
xor UO_1874 (O_1874,N_19995,N_19927);
xor UO_1875 (O_1875,N_19646,N_19817);
xnor UO_1876 (O_1876,N_19696,N_19986);
xor UO_1877 (O_1877,N_19610,N_19736);
xnor UO_1878 (O_1878,N_19977,N_19714);
or UO_1879 (O_1879,N_19633,N_19941);
or UO_1880 (O_1880,N_19839,N_19769);
nor UO_1881 (O_1881,N_19850,N_19945);
nor UO_1882 (O_1882,N_19857,N_19713);
nor UO_1883 (O_1883,N_19641,N_19991);
or UO_1884 (O_1884,N_19919,N_19931);
xnor UO_1885 (O_1885,N_19986,N_19845);
nor UO_1886 (O_1886,N_19898,N_19808);
and UO_1887 (O_1887,N_19949,N_19965);
xnor UO_1888 (O_1888,N_19710,N_19798);
or UO_1889 (O_1889,N_19691,N_19774);
nor UO_1890 (O_1890,N_19944,N_19777);
xor UO_1891 (O_1891,N_19830,N_19751);
nand UO_1892 (O_1892,N_19794,N_19812);
nand UO_1893 (O_1893,N_19639,N_19785);
xnor UO_1894 (O_1894,N_19875,N_19752);
or UO_1895 (O_1895,N_19670,N_19966);
nand UO_1896 (O_1896,N_19836,N_19734);
and UO_1897 (O_1897,N_19644,N_19898);
xor UO_1898 (O_1898,N_19961,N_19997);
nor UO_1899 (O_1899,N_19635,N_19719);
xnor UO_1900 (O_1900,N_19894,N_19774);
or UO_1901 (O_1901,N_19851,N_19927);
nand UO_1902 (O_1902,N_19827,N_19956);
nor UO_1903 (O_1903,N_19974,N_19779);
nand UO_1904 (O_1904,N_19648,N_19713);
and UO_1905 (O_1905,N_19664,N_19773);
or UO_1906 (O_1906,N_19959,N_19710);
nand UO_1907 (O_1907,N_19946,N_19664);
and UO_1908 (O_1908,N_19611,N_19959);
nand UO_1909 (O_1909,N_19833,N_19639);
and UO_1910 (O_1910,N_19803,N_19889);
nand UO_1911 (O_1911,N_19835,N_19991);
nand UO_1912 (O_1912,N_19889,N_19686);
or UO_1913 (O_1913,N_19779,N_19898);
nor UO_1914 (O_1914,N_19693,N_19634);
and UO_1915 (O_1915,N_19870,N_19650);
nand UO_1916 (O_1916,N_19905,N_19932);
nor UO_1917 (O_1917,N_19764,N_19689);
nor UO_1918 (O_1918,N_19626,N_19938);
xor UO_1919 (O_1919,N_19845,N_19898);
nor UO_1920 (O_1920,N_19894,N_19804);
nor UO_1921 (O_1921,N_19772,N_19930);
nor UO_1922 (O_1922,N_19813,N_19613);
nor UO_1923 (O_1923,N_19972,N_19802);
or UO_1924 (O_1924,N_19810,N_19883);
nor UO_1925 (O_1925,N_19955,N_19751);
nor UO_1926 (O_1926,N_19606,N_19613);
and UO_1927 (O_1927,N_19884,N_19963);
xnor UO_1928 (O_1928,N_19628,N_19721);
or UO_1929 (O_1929,N_19772,N_19747);
or UO_1930 (O_1930,N_19911,N_19789);
xor UO_1931 (O_1931,N_19708,N_19628);
or UO_1932 (O_1932,N_19773,N_19886);
nand UO_1933 (O_1933,N_19692,N_19805);
and UO_1934 (O_1934,N_19762,N_19710);
xnor UO_1935 (O_1935,N_19630,N_19815);
nand UO_1936 (O_1936,N_19780,N_19967);
nand UO_1937 (O_1937,N_19792,N_19947);
nand UO_1938 (O_1938,N_19699,N_19982);
or UO_1939 (O_1939,N_19854,N_19933);
or UO_1940 (O_1940,N_19721,N_19814);
nor UO_1941 (O_1941,N_19614,N_19990);
nor UO_1942 (O_1942,N_19821,N_19773);
xnor UO_1943 (O_1943,N_19971,N_19827);
xor UO_1944 (O_1944,N_19922,N_19634);
or UO_1945 (O_1945,N_19835,N_19731);
xor UO_1946 (O_1946,N_19693,N_19948);
and UO_1947 (O_1947,N_19962,N_19838);
nor UO_1948 (O_1948,N_19742,N_19674);
and UO_1949 (O_1949,N_19684,N_19903);
or UO_1950 (O_1950,N_19622,N_19836);
and UO_1951 (O_1951,N_19613,N_19672);
and UO_1952 (O_1952,N_19800,N_19912);
xor UO_1953 (O_1953,N_19851,N_19606);
nor UO_1954 (O_1954,N_19728,N_19747);
and UO_1955 (O_1955,N_19791,N_19919);
or UO_1956 (O_1956,N_19986,N_19942);
or UO_1957 (O_1957,N_19775,N_19761);
xor UO_1958 (O_1958,N_19784,N_19608);
nand UO_1959 (O_1959,N_19800,N_19694);
xor UO_1960 (O_1960,N_19915,N_19725);
nand UO_1961 (O_1961,N_19890,N_19665);
or UO_1962 (O_1962,N_19873,N_19950);
nor UO_1963 (O_1963,N_19988,N_19976);
or UO_1964 (O_1964,N_19694,N_19774);
nor UO_1965 (O_1965,N_19740,N_19766);
nand UO_1966 (O_1966,N_19924,N_19608);
and UO_1967 (O_1967,N_19842,N_19740);
nor UO_1968 (O_1968,N_19734,N_19775);
nor UO_1969 (O_1969,N_19859,N_19953);
or UO_1970 (O_1970,N_19849,N_19703);
xor UO_1971 (O_1971,N_19875,N_19966);
xor UO_1972 (O_1972,N_19974,N_19709);
xnor UO_1973 (O_1973,N_19895,N_19925);
nor UO_1974 (O_1974,N_19705,N_19864);
nor UO_1975 (O_1975,N_19734,N_19927);
nand UO_1976 (O_1976,N_19621,N_19873);
nor UO_1977 (O_1977,N_19968,N_19715);
or UO_1978 (O_1978,N_19706,N_19943);
or UO_1979 (O_1979,N_19826,N_19881);
xnor UO_1980 (O_1980,N_19969,N_19855);
xor UO_1981 (O_1981,N_19671,N_19718);
nand UO_1982 (O_1982,N_19956,N_19939);
nand UO_1983 (O_1983,N_19746,N_19745);
nor UO_1984 (O_1984,N_19769,N_19998);
nor UO_1985 (O_1985,N_19921,N_19846);
nand UO_1986 (O_1986,N_19935,N_19699);
nor UO_1987 (O_1987,N_19723,N_19782);
xor UO_1988 (O_1988,N_19689,N_19954);
or UO_1989 (O_1989,N_19738,N_19732);
nor UO_1990 (O_1990,N_19752,N_19767);
nand UO_1991 (O_1991,N_19900,N_19901);
or UO_1992 (O_1992,N_19998,N_19830);
and UO_1993 (O_1993,N_19674,N_19669);
and UO_1994 (O_1994,N_19884,N_19858);
or UO_1995 (O_1995,N_19734,N_19797);
and UO_1996 (O_1996,N_19606,N_19870);
and UO_1997 (O_1997,N_19839,N_19946);
nand UO_1998 (O_1998,N_19860,N_19749);
or UO_1999 (O_1999,N_19724,N_19909);
or UO_2000 (O_2000,N_19790,N_19623);
nand UO_2001 (O_2001,N_19911,N_19971);
xnor UO_2002 (O_2002,N_19784,N_19753);
or UO_2003 (O_2003,N_19669,N_19990);
nand UO_2004 (O_2004,N_19968,N_19848);
xnor UO_2005 (O_2005,N_19626,N_19957);
nor UO_2006 (O_2006,N_19963,N_19601);
and UO_2007 (O_2007,N_19745,N_19814);
or UO_2008 (O_2008,N_19673,N_19640);
or UO_2009 (O_2009,N_19883,N_19750);
or UO_2010 (O_2010,N_19905,N_19696);
xnor UO_2011 (O_2011,N_19888,N_19828);
or UO_2012 (O_2012,N_19974,N_19870);
xor UO_2013 (O_2013,N_19729,N_19867);
nand UO_2014 (O_2014,N_19607,N_19904);
or UO_2015 (O_2015,N_19902,N_19992);
nor UO_2016 (O_2016,N_19929,N_19986);
nand UO_2017 (O_2017,N_19764,N_19822);
nor UO_2018 (O_2018,N_19628,N_19809);
and UO_2019 (O_2019,N_19792,N_19828);
and UO_2020 (O_2020,N_19843,N_19699);
and UO_2021 (O_2021,N_19838,N_19667);
and UO_2022 (O_2022,N_19834,N_19891);
nor UO_2023 (O_2023,N_19897,N_19762);
nor UO_2024 (O_2024,N_19700,N_19710);
or UO_2025 (O_2025,N_19944,N_19797);
nand UO_2026 (O_2026,N_19765,N_19818);
xnor UO_2027 (O_2027,N_19822,N_19749);
nor UO_2028 (O_2028,N_19682,N_19676);
or UO_2029 (O_2029,N_19854,N_19970);
nand UO_2030 (O_2030,N_19647,N_19659);
and UO_2031 (O_2031,N_19788,N_19913);
nor UO_2032 (O_2032,N_19770,N_19608);
nand UO_2033 (O_2033,N_19973,N_19989);
and UO_2034 (O_2034,N_19891,N_19767);
nand UO_2035 (O_2035,N_19626,N_19930);
nor UO_2036 (O_2036,N_19944,N_19699);
nor UO_2037 (O_2037,N_19601,N_19614);
nand UO_2038 (O_2038,N_19775,N_19972);
nor UO_2039 (O_2039,N_19871,N_19715);
and UO_2040 (O_2040,N_19772,N_19769);
and UO_2041 (O_2041,N_19790,N_19804);
xnor UO_2042 (O_2042,N_19910,N_19686);
nor UO_2043 (O_2043,N_19867,N_19613);
xnor UO_2044 (O_2044,N_19791,N_19739);
or UO_2045 (O_2045,N_19926,N_19629);
xor UO_2046 (O_2046,N_19731,N_19775);
xor UO_2047 (O_2047,N_19651,N_19932);
and UO_2048 (O_2048,N_19787,N_19873);
nor UO_2049 (O_2049,N_19759,N_19947);
nand UO_2050 (O_2050,N_19933,N_19655);
or UO_2051 (O_2051,N_19902,N_19677);
or UO_2052 (O_2052,N_19688,N_19992);
or UO_2053 (O_2053,N_19665,N_19759);
or UO_2054 (O_2054,N_19882,N_19813);
nand UO_2055 (O_2055,N_19734,N_19984);
or UO_2056 (O_2056,N_19755,N_19634);
nand UO_2057 (O_2057,N_19955,N_19853);
nor UO_2058 (O_2058,N_19686,N_19654);
or UO_2059 (O_2059,N_19633,N_19723);
and UO_2060 (O_2060,N_19958,N_19660);
and UO_2061 (O_2061,N_19688,N_19979);
and UO_2062 (O_2062,N_19775,N_19835);
and UO_2063 (O_2063,N_19876,N_19849);
nand UO_2064 (O_2064,N_19941,N_19992);
nor UO_2065 (O_2065,N_19776,N_19719);
or UO_2066 (O_2066,N_19972,N_19674);
or UO_2067 (O_2067,N_19864,N_19812);
and UO_2068 (O_2068,N_19624,N_19894);
and UO_2069 (O_2069,N_19946,N_19842);
and UO_2070 (O_2070,N_19951,N_19644);
or UO_2071 (O_2071,N_19838,N_19830);
nand UO_2072 (O_2072,N_19694,N_19706);
nor UO_2073 (O_2073,N_19846,N_19902);
nor UO_2074 (O_2074,N_19645,N_19884);
nor UO_2075 (O_2075,N_19976,N_19801);
and UO_2076 (O_2076,N_19975,N_19800);
xor UO_2077 (O_2077,N_19950,N_19945);
xor UO_2078 (O_2078,N_19643,N_19930);
and UO_2079 (O_2079,N_19873,N_19866);
and UO_2080 (O_2080,N_19881,N_19692);
nand UO_2081 (O_2081,N_19764,N_19624);
nor UO_2082 (O_2082,N_19832,N_19659);
and UO_2083 (O_2083,N_19672,N_19960);
nor UO_2084 (O_2084,N_19941,N_19710);
and UO_2085 (O_2085,N_19635,N_19945);
nand UO_2086 (O_2086,N_19859,N_19676);
or UO_2087 (O_2087,N_19613,N_19892);
xor UO_2088 (O_2088,N_19626,N_19602);
and UO_2089 (O_2089,N_19837,N_19940);
or UO_2090 (O_2090,N_19992,N_19982);
nand UO_2091 (O_2091,N_19620,N_19627);
nor UO_2092 (O_2092,N_19733,N_19697);
and UO_2093 (O_2093,N_19861,N_19841);
or UO_2094 (O_2094,N_19847,N_19778);
and UO_2095 (O_2095,N_19958,N_19765);
or UO_2096 (O_2096,N_19617,N_19945);
nand UO_2097 (O_2097,N_19657,N_19668);
and UO_2098 (O_2098,N_19950,N_19982);
nand UO_2099 (O_2099,N_19801,N_19829);
nor UO_2100 (O_2100,N_19808,N_19796);
or UO_2101 (O_2101,N_19634,N_19815);
xor UO_2102 (O_2102,N_19733,N_19944);
xnor UO_2103 (O_2103,N_19845,N_19745);
or UO_2104 (O_2104,N_19930,N_19831);
nand UO_2105 (O_2105,N_19905,N_19921);
xnor UO_2106 (O_2106,N_19672,N_19809);
nor UO_2107 (O_2107,N_19753,N_19926);
or UO_2108 (O_2108,N_19787,N_19664);
nand UO_2109 (O_2109,N_19941,N_19773);
and UO_2110 (O_2110,N_19726,N_19691);
and UO_2111 (O_2111,N_19923,N_19961);
nand UO_2112 (O_2112,N_19786,N_19612);
nand UO_2113 (O_2113,N_19828,N_19946);
nand UO_2114 (O_2114,N_19932,N_19863);
nor UO_2115 (O_2115,N_19912,N_19818);
or UO_2116 (O_2116,N_19625,N_19907);
nand UO_2117 (O_2117,N_19612,N_19714);
or UO_2118 (O_2118,N_19614,N_19902);
and UO_2119 (O_2119,N_19743,N_19796);
nor UO_2120 (O_2120,N_19889,N_19605);
or UO_2121 (O_2121,N_19817,N_19922);
xor UO_2122 (O_2122,N_19794,N_19720);
and UO_2123 (O_2123,N_19886,N_19826);
xor UO_2124 (O_2124,N_19794,N_19773);
and UO_2125 (O_2125,N_19977,N_19769);
and UO_2126 (O_2126,N_19741,N_19839);
xor UO_2127 (O_2127,N_19838,N_19999);
and UO_2128 (O_2128,N_19903,N_19736);
and UO_2129 (O_2129,N_19792,N_19917);
xnor UO_2130 (O_2130,N_19757,N_19823);
xnor UO_2131 (O_2131,N_19957,N_19941);
and UO_2132 (O_2132,N_19945,N_19855);
and UO_2133 (O_2133,N_19819,N_19690);
nor UO_2134 (O_2134,N_19865,N_19762);
nand UO_2135 (O_2135,N_19862,N_19640);
nand UO_2136 (O_2136,N_19984,N_19751);
nand UO_2137 (O_2137,N_19669,N_19650);
or UO_2138 (O_2138,N_19863,N_19857);
or UO_2139 (O_2139,N_19603,N_19729);
and UO_2140 (O_2140,N_19903,N_19828);
nor UO_2141 (O_2141,N_19962,N_19615);
or UO_2142 (O_2142,N_19974,N_19665);
or UO_2143 (O_2143,N_19863,N_19621);
and UO_2144 (O_2144,N_19778,N_19884);
and UO_2145 (O_2145,N_19734,N_19685);
nor UO_2146 (O_2146,N_19737,N_19769);
nand UO_2147 (O_2147,N_19862,N_19733);
xor UO_2148 (O_2148,N_19896,N_19707);
nand UO_2149 (O_2149,N_19908,N_19956);
or UO_2150 (O_2150,N_19887,N_19754);
or UO_2151 (O_2151,N_19871,N_19967);
and UO_2152 (O_2152,N_19746,N_19864);
xnor UO_2153 (O_2153,N_19788,N_19691);
xnor UO_2154 (O_2154,N_19845,N_19836);
nor UO_2155 (O_2155,N_19624,N_19682);
or UO_2156 (O_2156,N_19894,N_19850);
and UO_2157 (O_2157,N_19844,N_19754);
nor UO_2158 (O_2158,N_19786,N_19708);
or UO_2159 (O_2159,N_19809,N_19800);
and UO_2160 (O_2160,N_19851,N_19850);
nand UO_2161 (O_2161,N_19615,N_19797);
nand UO_2162 (O_2162,N_19600,N_19908);
or UO_2163 (O_2163,N_19721,N_19788);
and UO_2164 (O_2164,N_19836,N_19781);
xor UO_2165 (O_2165,N_19684,N_19991);
and UO_2166 (O_2166,N_19751,N_19939);
and UO_2167 (O_2167,N_19759,N_19672);
or UO_2168 (O_2168,N_19911,N_19610);
xor UO_2169 (O_2169,N_19797,N_19757);
nor UO_2170 (O_2170,N_19896,N_19666);
nor UO_2171 (O_2171,N_19710,N_19989);
or UO_2172 (O_2172,N_19723,N_19658);
nor UO_2173 (O_2173,N_19809,N_19789);
xor UO_2174 (O_2174,N_19817,N_19894);
nor UO_2175 (O_2175,N_19602,N_19738);
nand UO_2176 (O_2176,N_19724,N_19831);
or UO_2177 (O_2177,N_19958,N_19629);
xnor UO_2178 (O_2178,N_19708,N_19983);
and UO_2179 (O_2179,N_19952,N_19863);
xor UO_2180 (O_2180,N_19652,N_19648);
nor UO_2181 (O_2181,N_19946,N_19642);
xor UO_2182 (O_2182,N_19607,N_19611);
or UO_2183 (O_2183,N_19783,N_19654);
nor UO_2184 (O_2184,N_19991,N_19715);
xnor UO_2185 (O_2185,N_19600,N_19726);
or UO_2186 (O_2186,N_19937,N_19960);
nor UO_2187 (O_2187,N_19853,N_19994);
and UO_2188 (O_2188,N_19650,N_19656);
xnor UO_2189 (O_2189,N_19695,N_19965);
or UO_2190 (O_2190,N_19921,N_19696);
nor UO_2191 (O_2191,N_19985,N_19872);
or UO_2192 (O_2192,N_19730,N_19814);
and UO_2193 (O_2193,N_19944,N_19632);
xor UO_2194 (O_2194,N_19748,N_19747);
nor UO_2195 (O_2195,N_19670,N_19657);
xor UO_2196 (O_2196,N_19711,N_19814);
nand UO_2197 (O_2197,N_19713,N_19780);
nand UO_2198 (O_2198,N_19649,N_19969);
or UO_2199 (O_2199,N_19763,N_19734);
and UO_2200 (O_2200,N_19723,N_19929);
or UO_2201 (O_2201,N_19850,N_19932);
or UO_2202 (O_2202,N_19998,N_19970);
xor UO_2203 (O_2203,N_19607,N_19972);
nor UO_2204 (O_2204,N_19645,N_19629);
nor UO_2205 (O_2205,N_19864,N_19631);
nor UO_2206 (O_2206,N_19908,N_19619);
and UO_2207 (O_2207,N_19820,N_19810);
nand UO_2208 (O_2208,N_19701,N_19886);
nand UO_2209 (O_2209,N_19653,N_19764);
and UO_2210 (O_2210,N_19741,N_19831);
or UO_2211 (O_2211,N_19643,N_19876);
nand UO_2212 (O_2212,N_19648,N_19666);
nand UO_2213 (O_2213,N_19680,N_19882);
nor UO_2214 (O_2214,N_19864,N_19618);
or UO_2215 (O_2215,N_19881,N_19799);
nor UO_2216 (O_2216,N_19679,N_19738);
and UO_2217 (O_2217,N_19734,N_19995);
nand UO_2218 (O_2218,N_19793,N_19786);
or UO_2219 (O_2219,N_19941,N_19863);
xor UO_2220 (O_2220,N_19627,N_19810);
xor UO_2221 (O_2221,N_19824,N_19873);
or UO_2222 (O_2222,N_19868,N_19980);
xor UO_2223 (O_2223,N_19637,N_19701);
or UO_2224 (O_2224,N_19708,N_19728);
or UO_2225 (O_2225,N_19818,N_19866);
or UO_2226 (O_2226,N_19684,N_19924);
nand UO_2227 (O_2227,N_19878,N_19967);
nor UO_2228 (O_2228,N_19696,N_19931);
xnor UO_2229 (O_2229,N_19974,N_19632);
nand UO_2230 (O_2230,N_19651,N_19669);
or UO_2231 (O_2231,N_19670,N_19887);
xor UO_2232 (O_2232,N_19766,N_19704);
xor UO_2233 (O_2233,N_19682,N_19929);
and UO_2234 (O_2234,N_19737,N_19764);
and UO_2235 (O_2235,N_19831,N_19696);
and UO_2236 (O_2236,N_19807,N_19897);
nand UO_2237 (O_2237,N_19957,N_19940);
nor UO_2238 (O_2238,N_19819,N_19837);
xor UO_2239 (O_2239,N_19661,N_19849);
nand UO_2240 (O_2240,N_19933,N_19626);
or UO_2241 (O_2241,N_19625,N_19734);
nor UO_2242 (O_2242,N_19694,N_19992);
and UO_2243 (O_2243,N_19934,N_19701);
xor UO_2244 (O_2244,N_19833,N_19956);
and UO_2245 (O_2245,N_19835,N_19837);
and UO_2246 (O_2246,N_19674,N_19969);
nand UO_2247 (O_2247,N_19917,N_19965);
nand UO_2248 (O_2248,N_19952,N_19761);
nand UO_2249 (O_2249,N_19620,N_19835);
nand UO_2250 (O_2250,N_19870,N_19636);
xor UO_2251 (O_2251,N_19793,N_19872);
xor UO_2252 (O_2252,N_19843,N_19668);
nor UO_2253 (O_2253,N_19614,N_19882);
xor UO_2254 (O_2254,N_19878,N_19776);
nor UO_2255 (O_2255,N_19869,N_19641);
and UO_2256 (O_2256,N_19823,N_19879);
nor UO_2257 (O_2257,N_19815,N_19802);
nor UO_2258 (O_2258,N_19737,N_19973);
nor UO_2259 (O_2259,N_19834,N_19915);
nand UO_2260 (O_2260,N_19607,N_19693);
or UO_2261 (O_2261,N_19688,N_19641);
or UO_2262 (O_2262,N_19960,N_19645);
nor UO_2263 (O_2263,N_19998,N_19916);
or UO_2264 (O_2264,N_19759,N_19950);
nor UO_2265 (O_2265,N_19815,N_19946);
nor UO_2266 (O_2266,N_19682,N_19658);
nand UO_2267 (O_2267,N_19954,N_19609);
xor UO_2268 (O_2268,N_19894,N_19901);
or UO_2269 (O_2269,N_19935,N_19865);
nand UO_2270 (O_2270,N_19871,N_19636);
nand UO_2271 (O_2271,N_19874,N_19852);
or UO_2272 (O_2272,N_19656,N_19983);
and UO_2273 (O_2273,N_19946,N_19668);
nand UO_2274 (O_2274,N_19620,N_19783);
nor UO_2275 (O_2275,N_19764,N_19852);
and UO_2276 (O_2276,N_19700,N_19805);
nand UO_2277 (O_2277,N_19641,N_19944);
and UO_2278 (O_2278,N_19762,N_19696);
nor UO_2279 (O_2279,N_19771,N_19674);
and UO_2280 (O_2280,N_19948,N_19950);
or UO_2281 (O_2281,N_19926,N_19698);
xnor UO_2282 (O_2282,N_19953,N_19783);
nor UO_2283 (O_2283,N_19762,N_19834);
nor UO_2284 (O_2284,N_19861,N_19804);
nor UO_2285 (O_2285,N_19954,N_19841);
and UO_2286 (O_2286,N_19709,N_19902);
nor UO_2287 (O_2287,N_19715,N_19971);
and UO_2288 (O_2288,N_19984,N_19739);
xor UO_2289 (O_2289,N_19914,N_19739);
or UO_2290 (O_2290,N_19840,N_19784);
and UO_2291 (O_2291,N_19947,N_19666);
or UO_2292 (O_2292,N_19973,N_19699);
or UO_2293 (O_2293,N_19856,N_19963);
xor UO_2294 (O_2294,N_19786,N_19643);
nor UO_2295 (O_2295,N_19737,N_19883);
and UO_2296 (O_2296,N_19662,N_19687);
or UO_2297 (O_2297,N_19764,N_19944);
nand UO_2298 (O_2298,N_19778,N_19761);
nor UO_2299 (O_2299,N_19941,N_19961);
xnor UO_2300 (O_2300,N_19638,N_19701);
nor UO_2301 (O_2301,N_19810,N_19754);
nor UO_2302 (O_2302,N_19948,N_19675);
xnor UO_2303 (O_2303,N_19639,N_19813);
or UO_2304 (O_2304,N_19786,N_19608);
nor UO_2305 (O_2305,N_19879,N_19636);
and UO_2306 (O_2306,N_19905,N_19946);
xnor UO_2307 (O_2307,N_19682,N_19816);
and UO_2308 (O_2308,N_19972,N_19609);
xor UO_2309 (O_2309,N_19789,N_19746);
nand UO_2310 (O_2310,N_19795,N_19971);
nor UO_2311 (O_2311,N_19734,N_19920);
and UO_2312 (O_2312,N_19849,N_19887);
and UO_2313 (O_2313,N_19909,N_19666);
nand UO_2314 (O_2314,N_19754,N_19743);
nor UO_2315 (O_2315,N_19763,N_19758);
xnor UO_2316 (O_2316,N_19711,N_19971);
nor UO_2317 (O_2317,N_19610,N_19726);
or UO_2318 (O_2318,N_19617,N_19812);
and UO_2319 (O_2319,N_19950,N_19695);
nor UO_2320 (O_2320,N_19605,N_19788);
or UO_2321 (O_2321,N_19707,N_19922);
nor UO_2322 (O_2322,N_19821,N_19659);
and UO_2323 (O_2323,N_19856,N_19927);
or UO_2324 (O_2324,N_19951,N_19714);
nor UO_2325 (O_2325,N_19858,N_19659);
nand UO_2326 (O_2326,N_19772,N_19736);
nand UO_2327 (O_2327,N_19707,N_19966);
nand UO_2328 (O_2328,N_19712,N_19721);
and UO_2329 (O_2329,N_19869,N_19829);
nor UO_2330 (O_2330,N_19846,N_19823);
and UO_2331 (O_2331,N_19989,N_19717);
or UO_2332 (O_2332,N_19946,N_19819);
nand UO_2333 (O_2333,N_19932,N_19754);
nor UO_2334 (O_2334,N_19961,N_19888);
xnor UO_2335 (O_2335,N_19758,N_19778);
or UO_2336 (O_2336,N_19708,N_19922);
xnor UO_2337 (O_2337,N_19849,N_19946);
and UO_2338 (O_2338,N_19657,N_19774);
nand UO_2339 (O_2339,N_19890,N_19962);
xnor UO_2340 (O_2340,N_19729,N_19701);
nand UO_2341 (O_2341,N_19884,N_19697);
nor UO_2342 (O_2342,N_19906,N_19865);
and UO_2343 (O_2343,N_19926,N_19636);
xnor UO_2344 (O_2344,N_19871,N_19990);
nor UO_2345 (O_2345,N_19837,N_19956);
xnor UO_2346 (O_2346,N_19928,N_19729);
and UO_2347 (O_2347,N_19746,N_19772);
nor UO_2348 (O_2348,N_19691,N_19843);
and UO_2349 (O_2349,N_19924,N_19747);
nand UO_2350 (O_2350,N_19720,N_19786);
nand UO_2351 (O_2351,N_19634,N_19796);
and UO_2352 (O_2352,N_19779,N_19828);
xnor UO_2353 (O_2353,N_19658,N_19690);
xor UO_2354 (O_2354,N_19678,N_19796);
xor UO_2355 (O_2355,N_19777,N_19672);
nand UO_2356 (O_2356,N_19675,N_19804);
or UO_2357 (O_2357,N_19927,N_19900);
or UO_2358 (O_2358,N_19646,N_19777);
and UO_2359 (O_2359,N_19941,N_19831);
xor UO_2360 (O_2360,N_19919,N_19950);
and UO_2361 (O_2361,N_19992,N_19772);
xor UO_2362 (O_2362,N_19710,N_19734);
xor UO_2363 (O_2363,N_19826,N_19719);
nand UO_2364 (O_2364,N_19605,N_19883);
xor UO_2365 (O_2365,N_19940,N_19711);
nand UO_2366 (O_2366,N_19988,N_19696);
or UO_2367 (O_2367,N_19696,N_19740);
xnor UO_2368 (O_2368,N_19916,N_19717);
or UO_2369 (O_2369,N_19926,N_19860);
nand UO_2370 (O_2370,N_19693,N_19752);
xor UO_2371 (O_2371,N_19959,N_19978);
and UO_2372 (O_2372,N_19756,N_19879);
xnor UO_2373 (O_2373,N_19686,N_19696);
and UO_2374 (O_2374,N_19914,N_19603);
or UO_2375 (O_2375,N_19998,N_19749);
and UO_2376 (O_2376,N_19932,N_19707);
xnor UO_2377 (O_2377,N_19907,N_19607);
xnor UO_2378 (O_2378,N_19806,N_19738);
and UO_2379 (O_2379,N_19728,N_19624);
nand UO_2380 (O_2380,N_19960,N_19708);
xnor UO_2381 (O_2381,N_19966,N_19845);
xnor UO_2382 (O_2382,N_19677,N_19815);
or UO_2383 (O_2383,N_19893,N_19968);
nor UO_2384 (O_2384,N_19616,N_19873);
nor UO_2385 (O_2385,N_19990,N_19641);
and UO_2386 (O_2386,N_19892,N_19895);
or UO_2387 (O_2387,N_19749,N_19945);
and UO_2388 (O_2388,N_19723,N_19955);
or UO_2389 (O_2389,N_19909,N_19720);
nand UO_2390 (O_2390,N_19787,N_19766);
xnor UO_2391 (O_2391,N_19749,N_19807);
nand UO_2392 (O_2392,N_19957,N_19943);
xnor UO_2393 (O_2393,N_19749,N_19802);
xor UO_2394 (O_2394,N_19972,N_19791);
or UO_2395 (O_2395,N_19706,N_19672);
nor UO_2396 (O_2396,N_19960,N_19976);
and UO_2397 (O_2397,N_19675,N_19772);
xor UO_2398 (O_2398,N_19846,N_19938);
and UO_2399 (O_2399,N_19889,N_19966);
nand UO_2400 (O_2400,N_19836,N_19849);
xnor UO_2401 (O_2401,N_19804,N_19706);
xor UO_2402 (O_2402,N_19670,N_19834);
nor UO_2403 (O_2403,N_19872,N_19672);
nor UO_2404 (O_2404,N_19775,N_19871);
or UO_2405 (O_2405,N_19828,N_19803);
nand UO_2406 (O_2406,N_19631,N_19787);
nand UO_2407 (O_2407,N_19978,N_19899);
or UO_2408 (O_2408,N_19624,N_19676);
and UO_2409 (O_2409,N_19790,N_19710);
xnor UO_2410 (O_2410,N_19604,N_19916);
nand UO_2411 (O_2411,N_19719,N_19747);
and UO_2412 (O_2412,N_19888,N_19962);
or UO_2413 (O_2413,N_19908,N_19837);
xor UO_2414 (O_2414,N_19648,N_19998);
nand UO_2415 (O_2415,N_19718,N_19857);
xor UO_2416 (O_2416,N_19910,N_19739);
or UO_2417 (O_2417,N_19775,N_19828);
nor UO_2418 (O_2418,N_19896,N_19886);
nor UO_2419 (O_2419,N_19895,N_19957);
nand UO_2420 (O_2420,N_19949,N_19998);
xor UO_2421 (O_2421,N_19979,N_19842);
or UO_2422 (O_2422,N_19939,N_19848);
xnor UO_2423 (O_2423,N_19630,N_19797);
nor UO_2424 (O_2424,N_19664,N_19793);
and UO_2425 (O_2425,N_19749,N_19827);
or UO_2426 (O_2426,N_19878,N_19861);
and UO_2427 (O_2427,N_19640,N_19866);
and UO_2428 (O_2428,N_19891,N_19602);
nor UO_2429 (O_2429,N_19768,N_19607);
nand UO_2430 (O_2430,N_19861,N_19748);
nand UO_2431 (O_2431,N_19602,N_19631);
and UO_2432 (O_2432,N_19942,N_19686);
nand UO_2433 (O_2433,N_19667,N_19872);
nor UO_2434 (O_2434,N_19682,N_19766);
and UO_2435 (O_2435,N_19766,N_19669);
or UO_2436 (O_2436,N_19755,N_19872);
nor UO_2437 (O_2437,N_19930,N_19809);
and UO_2438 (O_2438,N_19741,N_19861);
nor UO_2439 (O_2439,N_19937,N_19805);
and UO_2440 (O_2440,N_19925,N_19899);
nor UO_2441 (O_2441,N_19753,N_19994);
or UO_2442 (O_2442,N_19851,N_19654);
nor UO_2443 (O_2443,N_19962,N_19660);
nor UO_2444 (O_2444,N_19743,N_19830);
xnor UO_2445 (O_2445,N_19865,N_19660);
xor UO_2446 (O_2446,N_19962,N_19863);
nor UO_2447 (O_2447,N_19987,N_19984);
and UO_2448 (O_2448,N_19797,N_19949);
or UO_2449 (O_2449,N_19743,N_19872);
nor UO_2450 (O_2450,N_19629,N_19997);
nand UO_2451 (O_2451,N_19773,N_19808);
nor UO_2452 (O_2452,N_19687,N_19782);
or UO_2453 (O_2453,N_19935,N_19841);
nor UO_2454 (O_2454,N_19995,N_19638);
nor UO_2455 (O_2455,N_19696,N_19852);
xnor UO_2456 (O_2456,N_19846,N_19822);
nand UO_2457 (O_2457,N_19786,N_19602);
or UO_2458 (O_2458,N_19912,N_19857);
nand UO_2459 (O_2459,N_19842,N_19882);
xnor UO_2460 (O_2460,N_19974,N_19622);
nor UO_2461 (O_2461,N_19607,N_19691);
nor UO_2462 (O_2462,N_19971,N_19825);
nor UO_2463 (O_2463,N_19956,N_19742);
and UO_2464 (O_2464,N_19692,N_19718);
xnor UO_2465 (O_2465,N_19861,N_19636);
nand UO_2466 (O_2466,N_19948,N_19998);
xnor UO_2467 (O_2467,N_19781,N_19974);
and UO_2468 (O_2468,N_19871,N_19702);
nor UO_2469 (O_2469,N_19819,N_19863);
or UO_2470 (O_2470,N_19765,N_19612);
and UO_2471 (O_2471,N_19672,N_19625);
nand UO_2472 (O_2472,N_19934,N_19907);
nor UO_2473 (O_2473,N_19867,N_19876);
nand UO_2474 (O_2474,N_19741,N_19669);
nand UO_2475 (O_2475,N_19910,N_19870);
or UO_2476 (O_2476,N_19906,N_19860);
and UO_2477 (O_2477,N_19936,N_19890);
and UO_2478 (O_2478,N_19725,N_19949);
nor UO_2479 (O_2479,N_19870,N_19749);
and UO_2480 (O_2480,N_19799,N_19936);
nor UO_2481 (O_2481,N_19962,N_19755);
nor UO_2482 (O_2482,N_19999,N_19739);
nand UO_2483 (O_2483,N_19793,N_19982);
or UO_2484 (O_2484,N_19904,N_19613);
xnor UO_2485 (O_2485,N_19991,N_19704);
and UO_2486 (O_2486,N_19629,N_19968);
and UO_2487 (O_2487,N_19711,N_19717);
or UO_2488 (O_2488,N_19697,N_19783);
or UO_2489 (O_2489,N_19963,N_19629);
nor UO_2490 (O_2490,N_19633,N_19677);
or UO_2491 (O_2491,N_19967,N_19963);
xnor UO_2492 (O_2492,N_19892,N_19913);
or UO_2493 (O_2493,N_19968,N_19766);
nand UO_2494 (O_2494,N_19835,N_19984);
nor UO_2495 (O_2495,N_19829,N_19941);
and UO_2496 (O_2496,N_19686,N_19833);
or UO_2497 (O_2497,N_19757,N_19609);
nand UO_2498 (O_2498,N_19827,N_19865);
or UO_2499 (O_2499,N_19864,N_19816);
endmodule