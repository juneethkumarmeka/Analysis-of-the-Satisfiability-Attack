module basic_1500_15000_2000_10_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xnor U0 (N_0,In_524,In_1064);
nand U1 (N_1,In_485,In_1361);
nand U2 (N_2,In_230,In_922);
or U3 (N_3,In_964,In_450);
nor U4 (N_4,In_71,In_965);
and U5 (N_5,In_340,In_1105);
xnor U6 (N_6,In_300,In_708);
xor U7 (N_7,In_445,In_1236);
xor U8 (N_8,In_1337,In_638);
or U9 (N_9,In_1014,In_1238);
or U10 (N_10,In_428,In_162);
and U11 (N_11,In_6,In_1195);
and U12 (N_12,In_420,In_1397);
or U13 (N_13,In_395,In_1487);
nand U14 (N_14,In_1191,In_725);
nand U15 (N_15,In_990,In_1327);
xor U16 (N_16,In_1297,In_957);
or U17 (N_17,In_532,In_1204);
and U18 (N_18,In_329,In_1112);
and U19 (N_19,In_493,In_347);
nand U20 (N_20,In_627,In_381);
or U21 (N_21,In_1248,In_260);
nand U22 (N_22,In_446,In_80);
or U23 (N_23,In_831,In_951);
or U24 (N_24,In_1109,In_938);
nand U25 (N_25,In_779,In_737);
or U26 (N_26,In_919,In_1442);
xor U27 (N_27,In_89,In_1070);
nor U28 (N_28,In_1063,In_860);
nor U29 (N_29,In_21,In_114);
and U30 (N_30,In_622,In_1004);
nand U31 (N_31,In_1072,In_1402);
or U32 (N_32,In_418,In_1246);
or U33 (N_33,In_661,In_1111);
nand U34 (N_34,In_1051,In_92);
or U35 (N_35,In_542,In_384);
nor U36 (N_36,In_1092,In_264);
nor U37 (N_37,In_787,In_1285);
xor U38 (N_38,In_15,In_1374);
nand U39 (N_39,In_291,In_647);
and U40 (N_40,In_1131,In_1179);
and U41 (N_41,In_253,In_1443);
or U42 (N_42,In_1229,In_43);
or U43 (N_43,In_753,In_175);
nor U44 (N_44,In_516,In_1349);
nand U45 (N_45,In_25,In_920);
nor U46 (N_46,In_392,In_839);
nor U47 (N_47,In_339,In_1161);
nand U48 (N_48,In_1037,In_668);
or U49 (N_49,In_734,In_274);
nand U50 (N_50,In_410,In_1061);
or U51 (N_51,In_121,In_663);
nand U52 (N_52,In_1360,In_491);
or U53 (N_53,In_746,In_1008);
and U54 (N_54,In_864,In_2);
or U55 (N_55,In_34,In_1416);
nand U56 (N_56,In_1068,In_1433);
nor U57 (N_57,In_605,In_214);
and U58 (N_58,In_413,In_750);
and U59 (N_59,In_45,In_947);
nand U60 (N_60,In_1371,In_1394);
xnor U61 (N_61,In_1233,In_197);
nand U62 (N_62,In_1197,In_874);
xnor U63 (N_63,In_1474,In_767);
or U64 (N_64,In_1107,In_348);
xor U65 (N_65,In_1138,In_1216);
nand U66 (N_66,In_807,In_936);
or U67 (N_67,In_99,In_1214);
xor U68 (N_68,In_1206,In_459);
nor U69 (N_69,In_1032,In_824);
nand U70 (N_70,In_960,In_18);
nor U71 (N_71,In_287,In_1029);
xnor U72 (N_72,In_1345,In_157);
or U73 (N_73,In_93,In_5);
xor U74 (N_74,In_1430,In_308);
nand U75 (N_75,In_177,In_703);
nand U76 (N_76,In_482,In_48);
or U77 (N_77,In_1099,In_204);
and U78 (N_78,In_820,In_1428);
and U79 (N_79,In_1380,In_1451);
and U80 (N_80,In_616,In_698);
xor U81 (N_81,In_1239,In_1299);
nor U82 (N_82,In_697,In_973);
or U83 (N_83,In_1024,In_1359);
nor U84 (N_84,In_1200,In_306);
or U85 (N_85,In_160,In_766);
xor U86 (N_86,In_265,In_945);
and U87 (N_87,In_46,In_1322);
nor U88 (N_88,In_512,In_1346);
nand U89 (N_89,In_907,In_758);
xor U90 (N_90,In_189,In_568);
xor U91 (N_91,In_588,In_1266);
nand U92 (N_92,In_1053,In_1336);
and U93 (N_93,In_1104,In_722);
and U94 (N_94,In_1088,In_1211);
nor U95 (N_95,In_1291,In_364);
xor U96 (N_96,In_1243,In_579);
or U97 (N_97,In_1413,In_1465);
or U98 (N_98,In_87,In_137);
nand U99 (N_99,In_517,In_222);
xor U100 (N_100,In_140,In_553);
nand U101 (N_101,In_1084,In_151);
xor U102 (N_102,In_138,In_1173);
and U103 (N_103,In_1282,In_59);
or U104 (N_104,In_959,In_161);
nand U105 (N_105,In_50,In_169);
or U106 (N_106,In_771,In_227);
xor U107 (N_107,In_360,In_321);
xnor U108 (N_108,In_501,In_449);
or U109 (N_109,In_1011,In_586);
nor U110 (N_110,In_603,In_408);
xnor U111 (N_111,In_1202,In_694);
xor U112 (N_112,In_712,In_64);
nor U113 (N_113,In_967,In_1375);
xnor U114 (N_114,In_1033,In_1106);
nor U115 (N_115,In_505,In_609);
xnor U116 (N_116,In_112,In_953);
nand U117 (N_117,In_1146,In_728);
xnor U118 (N_118,In_991,In_1101);
or U119 (N_119,In_1075,In_723);
or U120 (N_120,In_27,In_233);
nand U121 (N_121,In_856,In_271);
or U122 (N_122,In_1365,In_662);
or U123 (N_123,In_427,In_126);
xnor U124 (N_124,In_1208,In_1393);
nand U125 (N_125,In_254,In_809);
and U126 (N_126,In_475,In_16);
nor U127 (N_127,In_232,In_909);
and U128 (N_128,In_871,In_10);
and U129 (N_129,In_726,In_896);
xnor U130 (N_130,In_671,In_336);
and U131 (N_131,In_925,In_334);
or U132 (N_132,In_382,In_426);
xnor U133 (N_133,In_317,In_1143);
nor U134 (N_134,In_778,In_421);
xnor U135 (N_135,In_970,In_700);
nor U136 (N_136,In_660,In_368);
nor U137 (N_137,In_1093,In_432);
and U138 (N_138,In_486,In_76);
nor U139 (N_139,In_361,In_223);
or U140 (N_140,In_63,In_1135);
or U141 (N_141,In_1426,In_803);
xor U142 (N_142,In_1497,In_1218);
nor U143 (N_143,In_379,In_133);
nor U144 (N_144,In_640,In_1445);
nand U145 (N_145,In_1231,In_1312);
nand U146 (N_146,In_1020,In_1010);
or U147 (N_147,In_585,In_437);
nor U148 (N_148,In_424,In_1252);
nor U149 (N_149,In_966,In_66);
and U150 (N_150,In_1398,In_95);
nand U151 (N_151,In_213,In_1047);
xor U152 (N_152,In_794,In_207);
and U153 (N_153,In_139,In_1189);
or U154 (N_154,In_425,In_855);
xnor U155 (N_155,In_613,In_390);
nor U156 (N_156,In_467,In_1471);
and U157 (N_157,In_132,In_955);
xnor U158 (N_158,In_648,In_191);
nor U159 (N_159,In_288,In_240);
nor U160 (N_160,In_812,In_208);
nor U161 (N_161,In_178,In_1119);
xnor U162 (N_162,In_286,In_304);
and U163 (N_163,In_1254,In_1005);
xor U164 (N_164,In_1247,In_389);
nand U165 (N_165,In_1268,In_67);
nand U166 (N_166,In_780,In_1357);
nor U167 (N_167,In_236,In_396);
or U168 (N_168,In_1326,In_1155);
xnor U169 (N_169,In_309,In_101);
or U170 (N_170,In_544,In_623);
nand U171 (N_171,In_1,In_1355);
xnor U172 (N_172,In_943,In_1083);
xor U173 (N_173,In_1235,In_1320);
or U174 (N_174,In_356,In_536);
nor U175 (N_175,In_713,In_885);
or U176 (N_176,In_520,In_331);
xnor U177 (N_177,In_685,In_183);
xnor U178 (N_178,In_740,In_159);
or U179 (N_179,In_1097,In_301);
and U180 (N_180,In_198,In_124);
and U181 (N_181,In_370,In_1036);
and U182 (N_182,In_1126,In_910);
nor U183 (N_183,In_1491,In_1418);
nand U184 (N_184,In_111,In_1407);
nor U185 (N_185,In_634,In_73);
or U186 (N_186,In_678,In_1016);
xnor U187 (N_187,In_19,In_674);
or U188 (N_188,In_1453,In_689);
nand U189 (N_189,In_709,In_1158);
and U190 (N_190,In_937,In_1180);
nand U191 (N_191,In_914,In_838);
xnor U192 (N_192,In_894,In_1153);
and U193 (N_193,In_1294,In_983);
nand U194 (N_194,In_1108,In_1164);
or U195 (N_195,In_1116,In_65);
xor U196 (N_196,In_215,In_1241);
nor U197 (N_197,In_594,In_147);
and U198 (N_198,In_362,In_523);
xnor U199 (N_199,In_1492,In_377);
or U200 (N_200,In_367,In_455);
nor U201 (N_201,In_268,In_631);
nand U202 (N_202,In_719,In_399);
or U203 (N_203,In_515,In_980);
xnor U204 (N_204,In_1178,In_136);
or U205 (N_205,In_1421,In_715);
nand U206 (N_206,In_1415,In_262);
nand U207 (N_207,In_656,In_759);
nor U208 (N_208,In_996,In_565);
xnor U209 (N_209,In_851,In_174);
and U210 (N_210,In_688,In_13);
nor U211 (N_211,In_606,In_1048);
xor U212 (N_212,In_720,In_1201);
nand U213 (N_213,In_220,In_1270);
and U214 (N_214,In_352,In_120);
and U215 (N_215,In_884,In_1425);
nor U216 (N_216,In_1256,In_672);
and U217 (N_217,In_1103,In_1009);
and U218 (N_218,In_567,In_513);
xnor U219 (N_219,In_483,In_1427);
nor U220 (N_220,In_1102,In_701);
and U221 (N_221,In_745,In_590);
and U222 (N_222,In_571,In_252);
nand U223 (N_223,In_75,In_1262);
and U224 (N_224,In_514,In_448);
nor U225 (N_225,In_507,In_394);
nor U226 (N_226,In_1123,In_91);
and U227 (N_227,In_42,In_799);
and U228 (N_228,In_739,In_33);
and U229 (N_229,In_774,In_1403);
or U230 (N_230,In_714,In_1478);
nor U231 (N_231,In_742,In_504);
xor U232 (N_232,In_332,In_267);
nor U233 (N_233,In_1227,In_1187);
or U234 (N_234,In_155,In_108);
xnor U235 (N_235,In_1392,In_1333);
and U236 (N_236,In_70,In_1387);
or U237 (N_237,In_1076,In_30);
xor U238 (N_238,In_74,In_266);
xor U239 (N_239,In_60,In_429);
nor U240 (N_240,In_1376,In_61);
nor U241 (N_241,In_154,In_1279);
or U242 (N_242,In_889,In_1039);
or U243 (N_243,In_439,In_229);
nor U244 (N_244,In_1089,In_890);
and U245 (N_245,In_247,In_310);
nor U246 (N_246,In_351,In_1446);
or U247 (N_247,In_939,In_1001);
nand U248 (N_248,In_1452,In_573);
and U249 (N_249,In_679,In_1059);
xnor U250 (N_250,In_1196,In_1321);
nand U251 (N_251,In_1456,In_51);
and U252 (N_252,In_727,In_971);
nand U253 (N_253,In_217,In_1100);
or U254 (N_254,In_888,In_37);
nor U255 (N_255,In_813,In_433);
xnor U256 (N_256,In_805,In_1174);
nor U257 (N_257,In_77,In_158);
nand U258 (N_258,In_843,In_1269);
or U259 (N_259,In_570,In_1481);
or U260 (N_260,In_684,In_383);
xor U261 (N_261,In_950,In_582);
xor U262 (N_262,In_1385,In_366);
xor U263 (N_263,In_103,In_776);
nand U264 (N_264,In_1348,In_658);
xnor U265 (N_265,In_695,In_1364);
nand U266 (N_266,In_763,In_324);
xor U267 (N_267,In_284,In_273);
nand U268 (N_268,In_529,In_146);
nand U269 (N_269,In_302,In_1280);
xnor U270 (N_270,In_55,In_768);
nor U271 (N_271,In_447,In_562);
xnor U272 (N_272,In_1215,In_924);
nor U273 (N_273,In_531,In_201);
or U274 (N_274,In_591,In_1118);
or U275 (N_275,In_1461,In_113);
nor U276 (N_276,In_827,In_297);
nor U277 (N_277,In_1477,In_295);
nand U278 (N_278,In_850,In_928);
nor U279 (N_279,In_1017,In_1125);
nand U280 (N_280,In_869,In_858);
xnor U281 (N_281,In_354,In_1450);
and U282 (N_282,In_625,In_96);
nor U283 (N_283,In_600,In_875);
nand U284 (N_284,In_550,In_221);
and U285 (N_285,In_307,In_1475);
xor U286 (N_286,In_1171,In_604);
xor U287 (N_287,In_335,In_1226);
nor U288 (N_288,In_409,In_1205);
and U289 (N_289,In_985,In_1144);
and U290 (N_290,In_1275,In_338);
and U291 (N_291,In_211,In_235);
nand U292 (N_292,In_566,In_952);
xnor U293 (N_293,In_1352,In_202);
nand U294 (N_294,In_941,In_895);
nand U295 (N_295,In_577,In_682);
or U296 (N_296,In_1052,In_403);
or U297 (N_297,In_365,In_930);
xnor U298 (N_298,In_1486,In_1328);
nand U299 (N_299,In_692,In_393);
nand U300 (N_300,In_1133,In_1213);
or U301 (N_301,In_1021,In_496);
nand U302 (N_302,In_1259,In_163);
xor U303 (N_303,In_1002,In_974);
xnor U304 (N_304,In_330,In_1160);
nor U305 (N_305,In_1292,In_102);
xnor U306 (N_306,In_633,In_862);
nand U307 (N_307,In_918,In_1484);
and U308 (N_308,In_578,In_313);
xor U309 (N_309,In_276,In_1274);
nor U310 (N_310,In_1315,In_28);
and U311 (N_311,In_620,In_891);
or U312 (N_312,In_503,In_845);
nor U313 (N_313,In_86,In_643);
or U314 (N_314,In_1343,In_773);
or U315 (N_315,In_1354,In_690);
or U316 (N_316,In_107,In_817);
nand U317 (N_317,In_1168,In_312);
nand U318 (N_318,In_1234,In_1074);
nand U319 (N_319,In_23,In_411);
xor U320 (N_320,In_624,In_316);
xnor U321 (N_321,In_83,In_1124);
or U322 (N_322,In_1221,In_1080);
and U323 (N_323,In_1272,In_397);
or U324 (N_324,In_1082,In_628);
xor U325 (N_325,In_881,In_1495);
nand U326 (N_326,In_583,In_1490);
nor U327 (N_327,In_993,In_380);
or U328 (N_328,In_865,In_1183);
and U329 (N_329,In_593,In_328);
or U330 (N_330,In_1013,In_1289);
xnor U331 (N_331,In_1046,In_333);
xnor U332 (N_332,In_1431,In_1055);
xor U333 (N_333,In_1310,In_1399);
or U334 (N_334,In_1249,In_1018);
xor U335 (N_335,In_810,In_915);
nand U336 (N_336,In_842,In_88);
or U337 (N_337,In_1313,In_22);
or U338 (N_338,In_789,In_1341);
or U339 (N_339,In_462,In_1303);
nor U340 (N_340,In_664,In_675);
nor U341 (N_341,In_1309,In_1034);
nand U342 (N_342,In_314,In_533);
xor U343 (N_343,In_1258,In_704);
nand U344 (N_344,In_772,In_528);
or U345 (N_345,In_1412,In_1127);
or U346 (N_346,In_629,In_691);
xor U347 (N_347,In_829,In_463);
nand U348 (N_348,In_238,In_683);
or U349 (N_349,In_1145,In_555);
xnor U350 (N_350,In_441,In_785);
nor U351 (N_351,In_1237,In_1458);
nand U352 (N_352,In_849,In_168);
nor U353 (N_353,In_1261,In_3);
xnor U354 (N_354,In_1347,In_815);
nand U355 (N_355,In_1460,In_1007);
nor U356 (N_356,In_981,In_893);
nor U357 (N_357,In_944,In_357);
or U358 (N_358,In_1411,In_319);
nor U359 (N_359,In_755,In_181);
or U360 (N_360,In_12,In_0);
and U361 (N_361,In_1087,In_574);
and U362 (N_362,In_791,In_182);
nor U363 (N_363,In_749,In_1057);
xnor U364 (N_364,In_490,In_934);
xnor U365 (N_365,In_434,In_4);
xor U366 (N_366,In_68,In_1470);
nor U367 (N_367,In_1071,In_797);
or U368 (N_368,In_987,In_1283);
and U369 (N_369,In_1340,In_495);
nand U370 (N_370,In_1028,In_203);
nor U371 (N_371,In_1128,In_241);
or U372 (N_372,In_537,In_109);
xor U373 (N_373,In_134,In_1031);
nand U374 (N_374,In_552,In_469);
or U375 (N_375,In_1485,In_721);
xnor U376 (N_376,In_696,In_545);
or U377 (N_377,In_251,In_1467);
nor U378 (N_378,In_1194,In_747);
nand U379 (N_379,In_311,In_617);
nor U380 (N_380,In_1339,In_670);
nor U381 (N_381,In_632,In_1351);
nand U382 (N_382,In_1081,In_752);
nor U383 (N_383,In_775,In_461);
nand U384 (N_384,In_948,In_1225);
nor U385 (N_385,In_984,In_1366);
xor U386 (N_386,In_572,In_972);
or U387 (N_387,In_526,In_453);
nand U388 (N_388,In_770,In_917);
and U389 (N_389,In_818,In_901);
nand U390 (N_390,In_1113,In_1027);
nand U391 (N_391,In_886,In_857);
nor U392 (N_392,In_363,In_880);
and U393 (N_393,In_1260,In_1177);
and U394 (N_394,In_226,In_1382);
nor U395 (N_395,In_417,In_38);
or U396 (N_396,In_1219,In_1429);
or U397 (N_397,In_1157,In_116);
or U398 (N_398,In_1388,In_988);
xor U399 (N_399,In_318,In_1330);
nand U400 (N_400,In_584,In_1255);
or U401 (N_401,In_1190,In_873);
nor U402 (N_402,In_636,In_649);
or U403 (N_403,In_164,In_756);
nand U404 (N_404,In_748,In_601);
nor U405 (N_405,In_407,In_195);
xor U406 (N_406,In_1390,In_729);
and U407 (N_407,In_1163,In_466);
and U408 (N_408,In_497,In_724);
and U409 (N_409,In_800,In_968);
and U410 (N_410,In_1040,In_781);
nand U411 (N_411,In_1338,In_305);
xnor U412 (N_412,In_293,In_498);
nand U413 (N_413,In_196,In_595);
xor U414 (N_414,In_626,In_852);
or U415 (N_415,In_808,In_24);
nand U416 (N_416,In_206,In_1423);
and U417 (N_417,In_187,In_702);
xor U418 (N_418,In_956,In_1000);
nand U419 (N_419,In_190,In_510);
nand U420 (N_420,In_81,In_743);
or U421 (N_421,In_816,In_541);
and U422 (N_422,In_1245,In_777);
or U423 (N_423,In_1044,In_551);
nor U424 (N_424,In_927,In_298);
and U425 (N_425,In_1424,In_471);
nand U426 (N_426,In_1041,In_1149);
nand U427 (N_427,In_173,In_387);
and U428 (N_428,In_1316,In_110);
nand U429 (N_429,In_337,In_69);
nor U430 (N_430,In_769,In_419);
or U431 (N_431,In_961,In_35);
xor U432 (N_432,In_1134,In_1318);
and U433 (N_433,In_406,In_611);
nand U434 (N_434,In_958,In_472);
nand U435 (N_435,In_1420,In_1381);
or U436 (N_436,In_414,In_1401);
nand U437 (N_437,In_1367,In_599);
and U438 (N_438,In_615,In_608);
nor U439 (N_439,In_982,In_525);
nand U440 (N_440,In_470,In_1120);
nor U441 (N_441,In_1395,In_1496);
xor U442 (N_442,In_1409,In_557);
xnor U443 (N_443,In_476,In_156);
and U444 (N_444,In_693,In_7);
and U445 (N_445,In_846,In_994);
nor U446 (N_446,In_1483,In_706);
nand U447 (N_447,In_1482,In_14);
and U448 (N_448,In_563,In_1066);
nand U449 (N_449,In_144,In_1172);
nor U450 (N_450,In_1198,In_192);
nor U451 (N_451,In_841,In_1098);
and U452 (N_452,In_946,In_1265);
nand U453 (N_453,In_90,In_1045);
nor U454 (N_454,In_1410,In_404);
and U455 (N_455,In_761,In_989);
or U456 (N_456,In_20,In_833);
nor U457 (N_457,In_346,In_119);
nand U458 (N_458,In_320,In_653);
or U459 (N_459,In_373,In_569);
and U460 (N_460,In_258,In_659);
xnor U461 (N_461,In_677,In_979);
nand U462 (N_462,In_530,In_1078);
or U463 (N_463,In_710,In_166);
xnor U464 (N_464,In_508,In_738);
and U465 (N_465,In_1335,In_534);
nor U466 (N_466,In_1473,In_1073);
and U467 (N_467,In_630,In_995);
or U468 (N_468,In_152,In_853);
and U469 (N_469,In_54,In_883);
and U470 (N_470,In_484,In_741);
and U471 (N_471,In_430,In_296);
xnor U472 (N_472,In_1152,In_736);
or U473 (N_473,In_1244,In_442);
nand U474 (N_474,In_279,In_1408);
xnor U475 (N_475,In_1121,In_444);
xor U476 (N_476,In_145,In_194);
nor U477 (N_477,In_1181,In_281);
nor U478 (N_478,In_249,In_1166);
nor U479 (N_479,In_607,In_861);
or U480 (N_480,In_912,In_487);
xor U481 (N_481,In_1396,In_234);
and U482 (N_482,In_644,In_962);
or U483 (N_483,In_906,In_801);
nand U484 (N_484,In_1192,In_1379);
xnor U485 (N_485,In_511,In_921);
and U486 (N_486,In_451,In_1026);
or U487 (N_487,In_848,In_435);
nand U488 (N_488,In_506,In_478);
xnor U489 (N_489,In_1331,In_1447);
nand U490 (N_490,In_665,In_473);
nand U491 (N_491,In_1422,In_1184);
and U492 (N_492,In_1278,In_1488);
xor U493 (N_493,In_1095,In_1217);
or U494 (N_494,In_903,In_1466);
nand U495 (N_495,In_219,In_9);
nor U496 (N_496,In_543,In_500);
xnor U497 (N_497,In_997,In_795);
or U498 (N_498,In_402,In_1378);
nor U499 (N_499,In_244,In_376);
xnor U500 (N_500,In_602,In_1188);
xnor U501 (N_501,In_811,In_185);
xor U502 (N_502,In_1003,In_1372);
nand U503 (N_503,In_802,In_1077);
or U504 (N_504,In_125,In_1140);
and U505 (N_505,In_581,In_716);
nand U506 (N_506,In_1232,In_642);
or U507 (N_507,In_949,In_165);
xnor U508 (N_508,In_1440,In_468);
nand U509 (N_509,In_863,In_1096);
nand U510 (N_510,In_792,In_641);
nand U511 (N_511,In_47,In_153);
nor U512 (N_512,In_1295,In_1253);
and U513 (N_513,In_378,In_210);
or U514 (N_514,In_908,In_1454);
xnor U515 (N_515,In_242,In_290);
or U516 (N_516,In_1334,In_1267);
xnor U517 (N_517,In_1136,In_1368);
nor U518 (N_518,In_519,In_575);
nor U519 (N_519,In_1383,In_1298);
nor U520 (N_520,In_754,In_499);
or U521 (N_521,In_1193,In_1170);
and U522 (N_522,In_1043,In_1444);
xnor U523 (N_523,In_1350,In_1117);
xnor U524 (N_524,In_1094,In_122);
xnor U525 (N_525,In_1290,In_1449);
or U526 (N_526,In_1257,In_1147);
nor U527 (N_527,In_868,In_1223);
and U528 (N_528,In_782,In_294);
and U529 (N_529,In_245,In_913);
nand U530 (N_530,In_589,In_645);
nand U531 (N_531,In_11,In_892);
nor U532 (N_532,In_431,In_836);
nor U533 (N_533,In_148,In_452);
xnor U534 (N_534,In_285,In_1369);
or U535 (N_535,In_489,In_735);
nor U536 (N_536,In_592,In_902);
nor U537 (N_537,In_1284,In_744);
or U538 (N_538,In_904,In_1476);
or U539 (N_539,In_1353,In_877);
or U540 (N_540,In_186,In_1325);
xnor U541 (N_541,In_1494,In_176);
xor U542 (N_542,In_1150,In_1224);
nand U543 (N_543,In_558,In_976);
or U544 (N_544,In_1499,In_117);
and U545 (N_545,In_167,In_1023);
or U546 (N_546,In_39,In_707);
or U547 (N_547,In_1199,In_492);
and U548 (N_548,In_216,In_1463);
xnor U549 (N_549,In_1060,In_464);
or U550 (N_550,In_375,In_1030);
xor U551 (N_551,In_911,In_549);
or U552 (N_552,In_667,In_129);
or U553 (N_553,In_784,In_1176);
nand U554 (N_554,In_1302,In_1151);
xnor U555 (N_555,In_1251,In_932);
nand U556 (N_556,In_127,In_118);
and U557 (N_557,In_548,In_479);
or U558 (N_558,In_790,In_78);
nor U559 (N_559,In_1342,In_1207);
and U560 (N_560,In_303,In_458);
nor U561 (N_561,In_56,In_1271);
xor U562 (N_562,In_1035,In_32);
or U563 (N_563,In_933,In_731);
xor U564 (N_564,In_1319,In_1276);
and U565 (N_565,In_786,In_405);
or U566 (N_566,In_1356,In_57);
and U567 (N_567,In_1464,In_1228);
or U568 (N_568,In_977,In_854);
nor U569 (N_569,In_94,In_1050);
xor U570 (N_570,In_1438,In_1230);
or U571 (N_571,In_53,In_1242);
nand U572 (N_572,In_128,In_259);
and U573 (N_573,In_1344,In_228);
xor U574 (N_574,In_576,In_1414);
nand U575 (N_575,In_1468,In_170);
xnor U576 (N_576,In_277,In_876);
nor U577 (N_577,In_342,In_171);
nor U578 (N_578,In_243,In_872);
xnor U579 (N_579,In_1175,In_327);
xor U580 (N_580,In_1115,In_1263);
or U581 (N_581,In_8,In_527);
nor U582 (N_582,In_1286,In_1022);
xnor U583 (N_583,In_837,In_686);
nor U584 (N_584,In_1049,In_359);
or U585 (N_585,In_559,In_1086);
xnor U586 (N_586,In_699,In_765);
nand U587 (N_587,In_619,In_923);
nand U588 (N_588,In_1472,In_1090);
xnor U589 (N_589,In_456,In_454);
nor U590 (N_590,In_438,In_830);
xor U591 (N_591,In_1389,In_345);
and U592 (N_592,In_898,In_940);
nor U593 (N_593,In_283,In_184);
nand U594 (N_594,In_1110,In_926);
nand U595 (N_595,In_400,In_1306);
or U596 (N_596,In_255,In_832);
nand U597 (N_597,In_621,In_556);
nand U598 (N_598,In_1156,In_814);
and U599 (N_599,In_969,In_422);
nor U600 (N_600,In_358,In_374);
nand U601 (N_601,In_52,In_1363);
xnor U602 (N_602,In_538,In_278);
nor U603 (N_603,In_1240,In_1006);
or U604 (N_604,In_85,In_1159);
xor U605 (N_605,In_188,In_1362);
nand U606 (N_606,In_272,In_72);
or U607 (N_607,In_681,In_866);
or U608 (N_608,In_1489,In_651);
xnor U609 (N_609,In_385,In_823);
and U610 (N_610,In_199,In_1019);
nor U611 (N_611,In_494,In_31);
and U612 (N_612,In_261,In_539);
nand U613 (N_613,In_344,In_1185);
nand U614 (N_614,In_1304,In_1056);
or U615 (N_615,In_231,In_610);
and U616 (N_616,In_477,In_323);
nor U617 (N_617,In_1042,In_796);
or U618 (N_618,In_1287,In_900);
nand U619 (N_619,In_218,In_135);
and U620 (N_620,In_1384,In_1203);
xnor U621 (N_621,In_1169,In_1142);
nor U622 (N_622,In_123,In_986);
and U623 (N_623,In_718,In_929);
xnor U624 (N_624,In_1469,In_1165);
nand U625 (N_625,In_1358,In_460);
nor U626 (N_626,In_1436,In_205);
nor U627 (N_627,In_637,In_280);
xor U628 (N_628,In_1311,In_819);
nor U629 (N_629,In_369,In_1132);
xor U630 (N_630,In_1130,In_897);
nand U631 (N_631,In_349,In_547);
and U632 (N_632,In_669,In_521);
nand U633 (N_633,In_41,In_580);
and U634 (N_634,In_29,In_1308);
nor U635 (N_635,In_612,In_1281);
nor U636 (N_636,In_546,In_289);
nor U637 (N_637,In_1391,In_1058);
xor U638 (N_638,In_248,In_783);
and U639 (N_639,In_355,In_687);
and U640 (N_640,In_522,In_878);
and U641 (N_641,In_423,In_1129);
nand U642 (N_642,In_598,In_1137);
or U643 (N_643,In_416,In_1091);
xor U644 (N_644,In_680,In_353);
xor U645 (N_645,In_180,In_326);
nand U646 (N_646,In_751,In_540);
nor U647 (N_647,In_847,In_652);
or U648 (N_648,In_299,In_1212);
nand U649 (N_649,In_1154,In_762);
and U650 (N_650,In_554,In_1406);
and U651 (N_651,In_1448,In_179);
xnor U652 (N_652,In_1479,In_935);
xor U653 (N_653,In_666,In_415);
nor U654 (N_654,In_398,In_650);
xnor U655 (N_655,In_1434,In_518);
xnor U656 (N_656,In_646,In_760);
xor U657 (N_657,In_481,In_1437);
nor U658 (N_658,In_1012,In_711);
and U659 (N_659,In_256,In_825);
and U660 (N_660,In_1141,In_804);
nor U661 (N_661,In_931,In_535);
xnor U662 (N_662,In_341,In_1277);
xor U663 (N_663,In_62,In_1085);
nand U664 (N_664,In_733,In_879);
nor U665 (N_665,In_673,In_509);
and U666 (N_666,In_372,In_835);
and U667 (N_667,In_1480,In_1417);
or U668 (N_668,In_793,In_1148);
xor U669 (N_669,In_1065,In_1386);
nor U670 (N_670,In_1305,In_97);
nor U671 (N_671,In_597,In_457);
nand U672 (N_672,In_270,In_1186);
nor U673 (N_673,In_867,In_141);
or U674 (N_674,In_596,In_1264);
and U675 (N_675,In_106,In_1054);
or U676 (N_676,In_1296,In_1419);
nor U677 (N_677,In_36,In_1273);
nand U678 (N_678,In_1250,In_655);
or U679 (N_679,In_1167,In_1062);
and U680 (N_680,In_822,In_828);
or U681 (N_681,In_1400,In_730);
xor U682 (N_682,In_1370,In_26);
nor U683 (N_683,In_1329,In_840);
and U684 (N_684,In_992,In_826);
nor U685 (N_685,In_44,In_98);
nor U686 (N_686,In_1139,In_225);
and U687 (N_687,In_821,In_401);
nor U688 (N_688,In_322,In_1288);
and U689 (N_689,In_150,In_292);
and U690 (N_690,In_436,In_564);
and U691 (N_691,In_105,In_1122);
nand U692 (N_692,In_998,In_859);
and U693 (N_693,In_757,In_963);
xor U694 (N_694,In_104,In_488);
or U695 (N_695,In_788,In_1455);
or U696 (N_696,In_560,In_193);
nand U697 (N_697,In_58,In_388);
or U698 (N_698,In_172,In_440);
xnor U699 (N_699,In_1377,In_315);
xnor U700 (N_700,In_1220,In_224);
or U701 (N_701,In_1182,In_635);
nand U702 (N_702,In_1432,In_237);
nor U703 (N_703,In_732,In_200);
nor U704 (N_704,In_40,In_142);
nor U705 (N_705,In_561,In_412);
xnor U706 (N_706,In_1293,In_587);
nor U707 (N_707,In_1405,In_239);
xor U708 (N_708,In_257,In_1439);
nor U709 (N_709,In_899,In_844);
or U710 (N_710,In_209,In_1462);
nand U711 (N_711,In_350,In_905);
nor U712 (N_712,In_1314,In_502);
nor U713 (N_713,In_82,In_282);
or U714 (N_714,In_275,In_17);
nor U715 (N_715,In_942,In_657);
and U716 (N_716,In_1435,In_84);
nor U717 (N_717,In_246,In_1015);
or U718 (N_718,In_1222,In_343);
and U719 (N_719,In_1441,In_764);
and U720 (N_720,In_443,In_1210);
or U721 (N_721,In_325,In_999);
xnor U722 (N_722,In_1404,In_130);
or U723 (N_723,In_100,In_1457);
and U724 (N_724,In_386,In_1323);
nand U725 (N_725,In_1317,In_371);
nand U726 (N_726,In_1301,In_1332);
nor U727 (N_727,In_1493,In_798);
xor U728 (N_728,In_131,In_79);
and U729 (N_729,In_465,In_149);
xnor U730 (N_730,In_474,In_263);
xor U731 (N_731,In_212,In_676);
nor U732 (N_732,In_1162,In_1069);
or U733 (N_733,In_480,In_1324);
and U734 (N_734,In_705,In_978);
nor U735 (N_735,In_806,In_1498);
nor U736 (N_736,In_1300,In_639);
or U737 (N_737,In_269,In_115);
and U738 (N_738,In_1209,In_618);
nor U739 (N_739,In_391,In_49);
and U740 (N_740,In_954,In_1373);
or U741 (N_741,In_887,In_1079);
and U742 (N_742,In_614,In_975);
and U743 (N_743,In_250,In_1114);
and U744 (N_744,In_1025,In_143);
and U745 (N_745,In_882,In_916);
or U746 (N_746,In_834,In_1067);
or U747 (N_747,In_654,In_717);
nand U748 (N_748,In_1307,In_1038);
nor U749 (N_749,In_1459,In_870);
and U750 (N_750,In_448,In_511);
and U751 (N_751,In_885,In_1233);
nor U752 (N_752,In_1399,In_1396);
xor U753 (N_753,In_704,In_1054);
nor U754 (N_754,In_590,In_1193);
xor U755 (N_755,In_1265,In_660);
xnor U756 (N_756,In_689,In_952);
or U757 (N_757,In_1148,In_623);
xor U758 (N_758,In_163,In_511);
and U759 (N_759,In_1095,In_658);
nand U760 (N_760,In_732,In_816);
and U761 (N_761,In_582,In_1365);
xor U762 (N_762,In_490,In_7);
nand U763 (N_763,In_967,In_1120);
nor U764 (N_764,In_127,In_68);
nand U765 (N_765,In_358,In_662);
xor U766 (N_766,In_172,In_585);
nand U767 (N_767,In_1496,In_871);
xor U768 (N_768,In_168,In_207);
nor U769 (N_769,In_859,In_1208);
or U770 (N_770,In_508,In_335);
xnor U771 (N_771,In_764,In_863);
nor U772 (N_772,In_877,In_994);
xnor U773 (N_773,In_1153,In_314);
nand U774 (N_774,In_1333,In_716);
or U775 (N_775,In_1184,In_989);
xnor U776 (N_776,In_9,In_800);
xor U777 (N_777,In_52,In_390);
xor U778 (N_778,In_928,In_1087);
and U779 (N_779,In_840,In_937);
or U780 (N_780,In_1179,In_939);
nand U781 (N_781,In_193,In_610);
xnor U782 (N_782,In_7,In_965);
xnor U783 (N_783,In_869,In_414);
and U784 (N_784,In_330,In_133);
nand U785 (N_785,In_590,In_827);
nor U786 (N_786,In_280,In_591);
and U787 (N_787,In_490,In_1362);
and U788 (N_788,In_731,In_830);
and U789 (N_789,In_735,In_479);
nand U790 (N_790,In_28,In_421);
and U791 (N_791,In_1268,In_1065);
and U792 (N_792,In_9,In_1145);
and U793 (N_793,In_263,In_1229);
nor U794 (N_794,In_1310,In_725);
or U795 (N_795,In_586,In_248);
nand U796 (N_796,In_1250,In_1419);
nand U797 (N_797,In_823,In_1041);
nand U798 (N_798,In_9,In_501);
nand U799 (N_799,In_1242,In_284);
nand U800 (N_800,In_1339,In_1141);
and U801 (N_801,In_282,In_1074);
nor U802 (N_802,In_4,In_582);
and U803 (N_803,In_1079,In_173);
or U804 (N_804,In_22,In_1087);
nor U805 (N_805,In_502,In_948);
and U806 (N_806,In_456,In_1064);
xnor U807 (N_807,In_1434,In_827);
nor U808 (N_808,In_932,In_645);
and U809 (N_809,In_392,In_1152);
and U810 (N_810,In_906,In_1306);
nand U811 (N_811,In_596,In_232);
nor U812 (N_812,In_1473,In_703);
or U813 (N_813,In_1480,In_816);
and U814 (N_814,In_1150,In_287);
xnor U815 (N_815,In_1396,In_1030);
or U816 (N_816,In_1012,In_1000);
and U817 (N_817,In_55,In_1179);
nand U818 (N_818,In_1478,In_532);
or U819 (N_819,In_1435,In_398);
nor U820 (N_820,In_422,In_546);
and U821 (N_821,In_5,In_250);
xnor U822 (N_822,In_814,In_404);
xor U823 (N_823,In_1411,In_30);
xnor U824 (N_824,In_1485,In_866);
nand U825 (N_825,In_976,In_980);
or U826 (N_826,In_21,In_1448);
or U827 (N_827,In_995,In_1288);
or U828 (N_828,In_967,In_181);
nand U829 (N_829,In_824,In_458);
nor U830 (N_830,In_571,In_858);
nor U831 (N_831,In_886,In_155);
and U832 (N_832,In_924,In_1003);
nand U833 (N_833,In_1395,In_918);
nand U834 (N_834,In_1193,In_471);
nand U835 (N_835,In_578,In_1364);
or U836 (N_836,In_1007,In_97);
and U837 (N_837,In_301,In_220);
xor U838 (N_838,In_914,In_25);
or U839 (N_839,In_1017,In_256);
or U840 (N_840,In_582,In_963);
or U841 (N_841,In_417,In_370);
nand U842 (N_842,In_1421,In_1305);
nor U843 (N_843,In_13,In_342);
nor U844 (N_844,In_507,In_71);
nor U845 (N_845,In_478,In_562);
and U846 (N_846,In_870,In_226);
nand U847 (N_847,In_78,In_388);
and U848 (N_848,In_949,In_288);
xor U849 (N_849,In_689,In_947);
or U850 (N_850,In_72,In_995);
nor U851 (N_851,In_1322,In_234);
or U852 (N_852,In_1224,In_248);
nor U853 (N_853,In_115,In_1034);
nand U854 (N_854,In_622,In_996);
and U855 (N_855,In_1272,In_790);
and U856 (N_856,In_243,In_367);
nand U857 (N_857,In_154,In_161);
xnor U858 (N_858,In_1011,In_1227);
xnor U859 (N_859,In_1143,In_1415);
or U860 (N_860,In_254,In_179);
xor U861 (N_861,In_890,In_1145);
or U862 (N_862,In_552,In_726);
or U863 (N_863,In_584,In_186);
nor U864 (N_864,In_583,In_669);
xor U865 (N_865,In_82,In_696);
xor U866 (N_866,In_883,In_209);
or U867 (N_867,In_804,In_648);
and U868 (N_868,In_888,In_58);
or U869 (N_869,In_1013,In_793);
nand U870 (N_870,In_852,In_62);
xor U871 (N_871,In_986,In_465);
or U872 (N_872,In_687,In_1405);
nand U873 (N_873,In_605,In_754);
nor U874 (N_874,In_599,In_290);
or U875 (N_875,In_1222,In_11);
or U876 (N_876,In_401,In_538);
and U877 (N_877,In_142,In_446);
xnor U878 (N_878,In_996,In_1081);
nand U879 (N_879,In_1231,In_1454);
xnor U880 (N_880,In_628,In_470);
and U881 (N_881,In_773,In_593);
nand U882 (N_882,In_710,In_1307);
and U883 (N_883,In_81,In_1359);
nor U884 (N_884,In_1034,In_251);
and U885 (N_885,In_1389,In_451);
and U886 (N_886,In_859,In_98);
nor U887 (N_887,In_1395,In_574);
and U888 (N_888,In_525,In_444);
xnor U889 (N_889,In_1221,In_587);
nand U890 (N_890,In_444,In_1113);
and U891 (N_891,In_396,In_207);
xor U892 (N_892,In_635,In_429);
xor U893 (N_893,In_599,In_934);
and U894 (N_894,In_174,In_368);
or U895 (N_895,In_1205,In_1216);
xor U896 (N_896,In_576,In_879);
nor U897 (N_897,In_235,In_431);
nand U898 (N_898,In_1284,In_966);
nand U899 (N_899,In_1407,In_1049);
nor U900 (N_900,In_1140,In_754);
or U901 (N_901,In_504,In_202);
nor U902 (N_902,In_1105,In_401);
xnor U903 (N_903,In_1092,In_4);
nand U904 (N_904,In_196,In_252);
nor U905 (N_905,In_672,In_209);
nor U906 (N_906,In_890,In_69);
or U907 (N_907,In_510,In_349);
nand U908 (N_908,In_50,In_1477);
xor U909 (N_909,In_469,In_254);
xor U910 (N_910,In_784,In_621);
or U911 (N_911,In_1424,In_749);
and U912 (N_912,In_1007,In_117);
or U913 (N_913,In_1212,In_767);
and U914 (N_914,In_397,In_1259);
nand U915 (N_915,In_1475,In_163);
nand U916 (N_916,In_386,In_1448);
xnor U917 (N_917,In_957,In_1494);
nand U918 (N_918,In_321,In_1041);
nand U919 (N_919,In_433,In_485);
or U920 (N_920,In_17,In_186);
nor U921 (N_921,In_525,In_1131);
xnor U922 (N_922,In_1201,In_617);
xnor U923 (N_923,In_216,In_450);
xor U924 (N_924,In_26,In_443);
nand U925 (N_925,In_763,In_574);
xor U926 (N_926,In_440,In_232);
nor U927 (N_927,In_1032,In_326);
xnor U928 (N_928,In_901,In_900);
or U929 (N_929,In_924,In_1148);
nor U930 (N_930,In_1088,In_1093);
or U931 (N_931,In_113,In_441);
nor U932 (N_932,In_221,In_554);
or U933 (N_933,In_811,In_746);
xor U934 (N_934,In_1319,In_888);
or U935 (N_935,In_1488,In_719);
xor U936 (N_936,In_796,In_834);
and U937 (N_937,In_375,In_42);
or U938 (N_938,In_820,In_471);
nor U939 (N_939,In_256,In_545);
nand U940 (N_940,In_199,In_1315);
or U941 (N_941,In_198,In_777);
xnor U942 (N_942,In_905,In_97);
nor U943 (N_943,In_154,In_1217);
nand U944 (N_944,In_79,In_1257);
nand U945 (N_945,In_350,In_1241);
nand U946 (N_946,In_772,In_548);
or U947 (N_947,In_1083,In_1418);
and U948 (N_948,In_1249,In_1054);
or U949 (N_949,In_839,In_89);
nor U950 (N_950,In_502,In_914);
or U951 (N_951,In_1431,In_1094);
xor U952 (N_952,In_577,In_1259);
nand U953 (N_953,In_722,In_41);
xor U954 (N_954,In_752,In_712);
xnor U955 (N_955,In_503,In_1299);
nand U956 (N_956,In_608,In_611);
xor U957 (N_957,In_1350,In_741);
nor U958 (N_958,In_973,In_577);
nor U959 (N_959,In_799,In_625);
xor U960 (N_960,In_45,In_423);
or U961 (N_961,In_688,In_1431);
or U962 (N_962,In_625,In_328);
nor U963 (N_963,In_377,In_549);
or U964 (N_964,In_437,In_1045);
or U965 (N_965,In_1175,In_952);
xnor U966 (N_966,In_1358,In_324);
xnor U967 (N_967,In_430,In_582);
nand U968 (N_968,In_784,In_1111);
and U969 (N_969,In_1034,In_253);
and U970 (N_970,In_757,In_1434);
or U971 (N_971,In_1006,In_350);
nand U972 (N_972,In_1406,In_305);
or U973 (N_973,In_149,In_971);
nor U974 (N_974,In_487,In_1104);
nor U975 (N_975,In_407,In_268);
nand U976 (N_976,In_1203,In_905);
and U977 (N_977,In_1093,In_1213);
xor U978 (N_978,In_1472,In_404);
and U979 (N_979,In_666,In_634);
xor U980 (N_980,In_331,In_445);
xnor U981 (N_981,In_366,In_348);
nand U982 (N_982,In_799,In_124);
and U983 (N_983,In_809,In_1155);
nor U984 (N_984,In_998,In_7);
nand U985 (N_985,In_390,In_591);
xor U986 (N_986,In_1186,In_70);
and U987 (N_987,In_1161,In_1142);
nand U988 (N_988,In_1313,In_1382);
and U989 (N_989,In_554,In_906);
xor U990 (N_990,In_273,In_281);
nor U991 (N_991,In_741,In_994);
nand U992 (N_992,In_565,In_238);
or U993 (N_993,In_1270,In_889);
and U994 (N_994,In_451,In_730);
xor U995 (N_995,In_1356,In_1012);
and U996 (N_996,In_902,In_387);
xnor U997 (N_997,In_1005,In_557);
xor U998 (N_998,In_352,In_286);
xnor U999 (N_999,In_1497,In_1095);
nand U1000 (N_1000,In_581,In_1406);
and U1001 (N_1001,In_1115,In_522);
xor U1002 (N_1002,In_452,In_1170);
nand U1003 (N_1003,In_868,In_72);
or U1004 (N_1004,In_775,In_1002);
nor U1005 (N_1005,In_459,In_281);
xnor U1006 (N_1006,In_321,In_1045);
xor U1007 (N_1007,In_614,In_947);
nand U1008 (N_1008,In_171,In_744);
nand U1009 (N_1009,In_1463,In_989);
nand U1010 (N_1010,In_729,In_292);
or U1011 (N_1011,In_696,In_1410);
nor U1012 (N_1012,In_918,In_24);
or U1013 (N_1013,In_441,In_79);
nand U1014 (N_1014,In_330,In_1235);
or U1015 (N_1015,In_1434,In_1237);
and U1016 (N_1016,In_297,In_316);
nand U1017 (N_1017,In_764,In_1170);
nor U1018 (N_1018,In_833,In_717);
xnor U1019 (N_1019,In_238,In_706);
xnor U1020 (N_1020,In_906,In_190);
and U1021 (N_1021,In_1384,In_878);
nor U1022 (N_1022,In_1053,In_1124);
or U1023 (N_1023,In_741,In_1457);
xnor U1024 (N_1024,In_998,In_944);
and U1025 (N_1025,In_736,In_1337);
xor U1026 (N_1026,In_1287,In_1244);
or U1027 (N_1027,In_860,In_651);
nor U1028 (N_1028,In_856,In_610);
nand U1029 (N_1029,In_844,In_1013);
nand U1030 (N_1030,In_1304,In_204);
nor U1031 (N_1031,In_208,In_1310);
and U1032 (N_1032,In_1495,In_717);
nand U1033 (N_1033,In_1129,In_672);
nand U1034 (N_1034,In_988,In_1143);
nor U1035 (N_1035,In_247,In_885);
nand U1036 (N_1036,In_1488,In_1220);
or U1037 (N_1037,In_666,In_268);
or U1038 (N_1038,In_243,In_1016);
and U1039 (N_1039,In_440,In_635);
or U1040 (N_1040,In_1356,In_581);
or U1041 (N_1041,In_652,In_1485);
nor U1042 (N_1042,In_1338,In_289);
nor U1043 (N_1043,In_477,In_611);
or U1044 (N_1044,In_260,In_45);
nand U1045 (N_1045,In_367,In_591);
or U1046 (N_1046,In_708,In_1050);
or U1047 (N_1047,In_530,In_29);
nor U1048 (N_1048,In_753,In_1241);
and U1049 (N_1049,In_1450,In_265);
and U1050 (N_1050,In_1145,In_660);
and U1051 (N_1051,In_146,In_915);
or U1052 (N_1052,In_512,In_205);
or U1053 (N_1053,In_872,In_240);
nand U1054 (N_1054,In_139,In_1186);
nor U1055 (N_1055,In_1039,In_1125);
or U1056 (N_1056,In_405,In_63);
nand U1057 (N_1057,In_1478,In_906);
and U1058 (N_1058,In_914,In_639);
nand U1059 (N_1059,In_260,In_1341);
and U1060 (N_1060,In_1114,In_428);
nor U1061 (N_1061,In_261,In_290);
and U1062 (N_1062,In_918,In_185);
or U1063 (N_1063,In_509,In_395);
nand U1064 (N_1064,In_954,In_1073);
or U1065 (N_1065,In_6,In_496);
nor U1066 (N_1066,In_1101,In_1450);
and U1067 (N_1067,In_456,In_248);
nand U1068 (N_1068,In_920,In_1365);
or U1069 (N_1069,In_1400,In_207);
and U1070 (N_1070,In_91,In_841);
or U1071 (N_1071,In_1244,In_1371);
and U1072 (N_1072,In_1125,In_504);
nor U1073 (N_1073,In_1290,In_1417);
nand U1074 (N_1074,In_672,In_237);
xor U1075 (N_1075,In_750,In_1330);
and U1076 (N_1076,In_1315,In_603);
nand U1077 (N_1077,In_1203,In_1290);
nor U1078 (N_1078,In_390,In_302);
or U1079 (N_1079,In_1007,In_243);
nor U1080 (N_1080,In_967,In_1099);
nor U1081 (N_1081,In_1305,In_400);
nor U1082 (N_1082,In_508,In_831);
nand U1083 (N_1083,In_979,In_1279);
nand U1084 (N_1084,In_713,In_1475);
nand U1085 (N_1085,In_351,In_1258);
or U1086 (N_1086,In_910,In_412);
and U1087 (N_1087,In_1493,In_95);
and U1088 (N_1088,In_1166,In_29);
nand U1089 (N_1089,In_192,In_1466);
and U1090 (N_1090,In_84,In_209);
xor U1091 (N_1091,In_1259,In_259);
xor U1092 (N_1092,In_738,In_1321);
and U1093 (N_1093,In_1496,In_485);
and U1094 (N_1094,In_1488,In_1378);
or U1095 (N_1095,In_334,In_181);
nor U1096 (N_1096,In_1153,In_815);
nand U1097 (N_1097,In_397,In_322);
xor U1098 (N_1098,In_353,In_387);
xor U1099 (N_1099,In_391,In_840);
xor U1100 (N_1100,In_1292,In_1142);
xnor U1101 (N_1101,In_361,In_224);
nand U1102 (N_1102,In_516,In_605);
xor U1103 (N_1103,In_600,In_1369);
or U1104 (N_1104,In_980,In_766);
nand U1105 (N_1105,In_1192,In_791);
nand U1106 (N_1106,In_1393,In_285);
nor U1107 (N_1107,In_113,In_91);
xor U1108 (N_1108,In_1163,In_1353);
and U1109 (N_1109,In_814,In_717);
nand U1110 (N_1110,In_1477,In_142);
nand U1111 (N_1111,In_902,In_720);
nand U1112 (N_1112,In_1247,In_1377);
or U1113 (N_1113,In_1425,In_126);
nor U1114 (N_1114,In_264,In_1190);
or U1115 (N_1115,In_302,In_1073);
xnor U1116 (N_1116,In_781,In_729);
nor U1117 (N_1117,In_973,In_683);
nor U1118 (N_1118,In_1276,In_1255);
and U1119 (N_1119,In_757,In_695);
and U1120 (N_1120,In_1051,In_458);
nand U1121 (N_1121,In_1048,In_643);
nor U1122 (N_1122,In_757,In_1139);
or U1123 (N_1123,In_146,In_1069);
xor U1124 (N_1124,In_1122,In_148);
or U1125 (N_1125,In_983,In_170);
nor U1126 (N_1126,In_1462,In_743);
or U1127 (N_1127,In_1351,In_1310);
nand U1128 (N_1128,In_649,In_450);
xor U1129 (N_1129,In_725,In_1169);
nand U1130 (N_1130,In_250,In_1285);
and U1131 (N_1131,In_178,In_949);
nor U1132 (N_1132,In_988,In_1282);
nor U1133 (N_1133,In_1284,In_403);
nor U1134 (N_1134,In_345,In_893);
or U1135 (N_1135,In_37,In_325);
nor U1136 (N_1136,In_255,In_559);
and U1137 (N_1137,In_1115,In_363);
and U1138 (N_1138,In_390,In_170);
and U1139 (N_1139,In_482,In_1469);
or U1140 (N_1140,In_187,In_8);
nand U1141 (N_1141,In_976,In_1471);
or U1142 (N_1142,In_360,In_820);
xnor U1143 (N_1143,In_1205,In_1018);
or U1144 (N_1144,In_31,In_1265);
or U1145 (N_1145,In_493,In_1041);
or U1146 (N_1146,In_1102,In_470);
and U1147 (N_1147,In_640,In_798);
or U1148 (N_1148,In_1270,In_267);
and U1149 (N_1149,In_364,In_998);
xnor U1150 (N_1150,In_337,In_823);
or U1151 (N_1151,In_364,In_1349);
nor U1152 (N_1152,In_653,In_69);
nand U1153 (N_1153,In_194,In_130);
nor U1154 (N_1154,In_238,In_1147);
or U1155 (N_1155,In_269,In_798);
or U1156 (N_1156,In_1454,In_293);
nor U1157 (N_1157,In_446,In_1365);
or U1158 (N_1158,In_632,In_385);
or U1159 (N_1159,In_259,In_11);
nor U1160 (N_1160,In_183,In_831);
and U1161 (N_1161,In_1495,In_680);
nor U1162 (N_1162,In_499,In_623);
nand U1163 (N_1163,In_635,In_959);
nor U1164 (N_1164,In_671,In_419);
or U1165 (N_1165,In_995,In_1156);
nor U1166 (N_1166,In_998,In_37);
or U1167 (N_1167,In_74,In_1193);
and U1168 (N_1168,In_1328,In_1198);
xor U1169 (N_1169,In_1091,In_696);
nand U1170 (N_1170,In_1492,In_770);
nand U1171 (N_1171,In_1279,In_603);
and U1172 (N_1172,In_972,In_157);
xor U1173 (N_1173,In_337,In_16);
xor U1174 (N_1174,In_942,In_725);
or U1175 (N_1175,In_586,In_1159);
xnor U1176 (N_1176,In_89,In_1361);
xnor U1177 (N_1177,In_1398,In_418);
nor U1178 (N_1178,In_1260,In_821);
and U1179 (N_1179,In_253,In_1391);
nand U1180 (N_1180,In_836,In_628);
and U1181 (N_1181,In_357,In_1073);
or U1182 (N_1182,In_954,In_1412);
xnor U1183 (N_1183,In_1134,In_595);
nor U1184 (N_1184,In_1208,In_1304);
and U1185 (N_1185,In_884,In_56);
or U1186 (N_1186,In_1461,In_102);
xor U1187 (N_1187,In_1461,In_701);
and U1188 (N_1188,In_1121,In_1150);
nor U1189 (N_1189,In_1006,In_1428);
xor U1190 (N_1190,In_251,In_657);
or U1191 (N_1191,In_1230,In_978);
nor U1192 (N_1192,In_714,In_151);
nor U1193 (N_1193,In_40,In_1225);
and U1194 (N_1194,In_354,In_154);
nor U1195 (N_1195,In_1351,In_1442);
nor U1196 (N_1196,In_972,In_1020);
or U1197 (N_1197,In_698,In_341);
or U1198 (N_1198,In_489,In_797);
and U1199 (N_1199,In_299,In_928);
nand U1200 (N_1200,In_607,In_802);
nand U1201 (N_1201,In_598,In_465);
and U1202 (N_1202,In_1478,In_1345);
or U1203 (N_1203,In_1189,In_960);
nor U1204 (N_1204,In_950,In_94);
and U1205 (N_1205,In_275,In_1323);
nand U1206 (N_1206,In_276,In_743);
or U1207 (N_1207,In_1426,In_496);
or U1208 (N_1208,In_756,In_1299);
nor U1209 (N_1209,In_1170,In_1201);
or U1210 (N_1210,In_1300,In_1289);
nand U1211 (N_1211,In_1093,In_514);
xnor U1212 (N_1212,In_899,In_1471);
nand U1213 (N_1213,In_215,In_175);
nor U1214 (N_1214,In_1462,In_656);
nand U1215 (N_1215,In_1491,In_627);
or U1216 (N_1216,In_508,In_1278);
and U1217 (N_1217,In_1002,In_1258);
nor U1218 (N_1218,In_810,In_765);
and U1219 (N_1219,In_856,In_1061);
and U1220 (N_1220,In_1399,In_748);
or U1221 (N_1221,In_16,In_946);
nand U1222 (N_1222,In_18,In_287);
or U1223 (N_1223,In_1305,In_368);
and U1224 (N_1224,In_116,In_141);
and U1225 (N_1225,In_1030,In_261);
nand U1226 (N_1226,In_1417,In_365);
xnor U1227 (N_1227,In_747,In_662);
or U1228 (N_1228,In_1381,In_1210);
xnor U1229 (N_1229,In_851,In_640);
xor U1230 (N_1230,In_268,In_1479);
and U1231 (N_1231,In_1350,In_847);
or U1232 (N_1232,In_854,In_1002);
xor U1233 (N_1233,In_309,In_1175);
nor U1234 (N_1234,In_495,In_217);
nand U1235 (N_1235,In_1425,In_11);
nor U1236 (N_1236,In_1441,In_868);
nand U1237 (N_1237,In_953,In_1334);
nor U1238 (N_1238,In_17,In_902);
nand U1239 (N_1239,In_115,In_832);
and U1240 (N_1240,In_77,In_373);
or U1241 (N_1241,In_915,In_1073);
nand U1242 (N_1242,In_1284,In_81);
and U1243 (N_1243,In_174,In_1256);
or U1244 (N_1244,In_1321,In_420);
nand U1245 (N_1245,In_632,In_1027);
and U1246 (N_1246,In_956,In_1101);
and U1247 (N_1247,In_908,In_1195);
nor U1248 (N_1248,In_180,In_225);
nor U1249 (N_1249,In_242,In_1196);
or U1250 (N_1250,In_1135,In_132);
or U1251 (N_1251,In_609,In_821);
or U1252 (N_1252,In_583,In_403);
nand U1253 (N_1253,In_1450,In_999);
and U1254 (N_1254,In_323,In_744);
nor U1255 (N_1255,In_497,In_1259);
nand U1256 (N_1256,In_486,In_832);
xor U1257 (N_1257,In_33,In_223);
nor U1258 (N_1258,In_1372,In_645);
and U1259 (N_1259,In_1036,In_1167);
xnor U1260 (N_1260,In_670,In_42);
nand U1261 (N_1261,In_1049,In_311);
nor U1262 (N_1262,In_411,In_809);
and U1263 (N_1263,In_646,In_1010);
nand U1264 (N_1264,In_1316,In_1055);
xnor U1265 (N_1265,In_144,In_1389);
or U1266 (N_1266,In_92,In_840);
and U1267 (N_1267,In_295,In_496);
or U1268 (N_1268,In_885,In_397);
nor U1269 (N_1269,In_244,In_1135);
nor U1270 (N_1270,In_510,In_460);
xor U1271 (N_1271,In_1194,In_664);
xnor U1272 (N_1272,In_402,In_1206);
or U1273 (N_1273,In_625,In_233);
xor U1274 (N_1274,In_436,In_448);
nor U1275 (N_1275,In_821,In_1444);
nand U1276 (N_1276,In_968,In_376);
or U1277 (N_1277,In_963,In_1449);
nand U1278 (N_1278,In_446,In_255);
xor U1279 (N_1279,In_833,In_1330);
xnor U1280 (N_1280,In_1092,In_551);
nor U1281 (N_1281,In_762,In_687);
nor U1282 (N_1282,In_1079,In_345);
nor U1283 (N_1283,In_651,In_782);
nor U1284 (N_1284,In_282,In_523);
nand U1285 (N_1285,In_1391,In_862);
and U1286 (N_1286,In_36,In_780);
xnor U1287 (N_1287,In_768,In_362);
nand U1288 (N_1288,In_634,In_1218);
or U1289 (N_1289,In_1314,In_1029);
and U1290 (N_1290,In_1349,In_728);
nand U1291 (N_1291,In_350,In_858);
nand U1292 (N_1292,In_842,In_435);
and U1293 (N_1293,In_1032,In_1326);
nand U1294 (N_1294,In_761,In_1484);
and U1295 (N_1295,In_252,In_51);
nand U1296 (N_1296,In_910,In_1446);
and U1297 (N_1297,In_692,In_327);
nand U1298 (N_1298,In_768,In_102);
and U1299 (N_1299,In_345,In_968);
or U1300 (N_1300,In_631,In_825);
or U1301 (N_1301,In_1395,In_373);
or U1302 (N_1302,In_503,In_83);
xor U1303 (N_1303,In_670,In_613);
or U1304 (N_1304,In_921,In_39);
or U1305 (N_1305,In_84,In_1454);
xor U1306 (N_1306,In_1036,In_1354);
or U1307 (N_1307,In_1279,In_576);
xor U1308 (N_1308,In_312,In_1293);
xor U1309 (N_1309,In_771,In_1137);
nand U1310 (N_1310,In_1245,In_433);
or U1311 (N_1311,In_714,In_803);
or U1312 (N_1312,In_896,In_482);
nand U1313 (N_1313,In_378,In_412);
xnor U1314 (N_1314,In_22,In_1238);
nor U1315 (N_1315,In_582,In_698);
nand U1316 (N_1316,In_537,In_733);
or U1317 (N_1317,In_109,In_990);
xnor U1318 (N_1318,In_86,In_1063);
and U1319 (N_1319,In_996,In_199);
nor U1320 (N_1320,In_1459,In_299);
xor U1321 (N_1321,In_1379,In_513);
nor U1322 (N_1322,In_617,In_86);
nor U1323 (N_1323,In_633,In_191);
and U1324 (N_1324,In_900,In_228);
nor U1325 (N_1325,In_249,In_166);
and U1326 (N_1326,In_1354,In_569);
xnor U1327 (N_1327,In_518,In_606);
or U1328 (N_1328,In_102,In_1212);
or U1329 (N_1329,In_1232,In_960);
and U1330 (N_1330,In_841,In_1031);
nor U1331 (N_1331,In_744,In_849);
nor U1332 (N_1332,In_191,In_1456);
nor U1333 (N_1333,In_30,In_51);
and U1334 (N_1334,In_1214,In_640);
or U1335 (N_1335,In_869,In_1307);
xnor U1336 (N_1336,In_646,In_1396);
and U1337 (N_1337,In_937,In_11);
nor U1338 (N_1338,In_538,In_956);
and U1339 (N_1339,In_1477,In_478);
and U1340 (N_1340,In_1360,In_1115);
or U1341 (N_1341,In_380,In_747);
or U1342 (N_1342,In_1221,In_1032);
nor U1343 (N_1343,In_1128,In_1335);
and U1344 (N_1344,In_887,In_336);
nand U1345 (N_1345,In_1417,In_88);
xnor U1346 (N_1346,In_758,In_1398);
nor U1347 (N_1347,In_152,In_423);
nand U1348 (N_1348,In_832,In_1277);
or U1349 (N_1349,In_1218,In_731);
or U1350 (N_1350,In_18,In_643);
nor U1351 (N_1351,In_513,In_819);
nor U1352 (N_1352,In_1471,In_245);
nand U1353 (N_1353,In_330,In_799);
nand U1354 (N_1354,In_119,In_708);
xor U1355 (N_1355,In_138,In_1260);
or U1356 (N_1356,In_646,In_1202);
and U1357 (N_1357,In_804,In_1072);
xnor U1358 (N_1358,In_685,In_18);
or U1359 (N_1359,In_756,In_66);
or U1360 (N_1360,In_1122,In_1000);
and U1361 (N_1361,In_1297,In_1364);
xor U1362 (N_1362,In_770,In_551);
nor U1363 (N_1363,In_2,In_625);
nand U1364 (N_1364,In_879,In_1181);
or U1365 (N_1365,In_590,In_702);
nand U1366 (N_1366,In_172,In_1231);
and U1367 (N_1367,In_932,In_59);
xor U1368 (N_1368,In_348,In_547);
nor U1369 (N_1369,In_1078,In_817);
and U1370 (N_1370,In_158,In_753);
or U1371 (N_1371,In_1416,In_782);
nor U1372 (N_1372,In_149,In_1261);
xor U1373 (N_1373,In_920,In_1401);
or U1374 (N_1374,In_157,In_1119);
xor U1375 (N_1375,In_1154,In_1265);
xnor U1376 (N_1376,In_173,In_679);
nor U1377 (N_1377,In_1282,In_550);
or U1378 (N_1378,In_1485,In_163);
nand U1379 (N_1379,In_393,In_383);
nand U1380 (N_1380,In_777,In_163);
nand U1381 (N_1381,In_18,In_391);
xor U1382 (N_1382,In_272,In_421);
or U1383 (N_1383,In_1364,In_1193);
or U1384 (N_1384,In_987,In_777);
xnor U1385 (N_1385,In_141,In_598);
nor U1386 (N_1386,In_70,In_356);
or U1387 (N_1387,In_108,In_1115);
and U1388 (N_1388,In_166,In_1196);
and U1389 (N_1389,In_1339,In_936);
nor U1390 (N_1390,In_96,In_10);
and U1391 (N_1391,In_1148,In_11);
nand U1392 (N_1392,In_1195,In_516);
nor U1393 (N_1393,In_449,In_349);
xnor U1394 (N_1394,In_1076,In_574);
nor U1395 (N_1395,In_1003,In_1216);
xor U1396 (N_1396,In_299,In_1488);
nor U1397 (N_1397,In_507,In_278);
xor U1398 (N_1398,In_345,In_697);
nor U1399 (N_1399,In_872,In_404);
nand U1400 (N_1400,In_562,In_1147);
and U1401 (N_1401,In_1193,In_1231);
xor U1402 (N_1402,In_20,In_271);
and U1403 (N_1403,In_1262,In_646);
xor U1404 (N_1404,In_196,In_814);
xnor U1405 (N_1405,In_902,In_1434);
nor U1406 (N_1406,In_695,In_439);
and U1407 (N_1407,In_446,In_72);
nand U1408 (N_1408,In_153,In_1130);
and U1409 (N_1409,In_413,In_867);
nand U1410 (N_1410,In_97,In_549);
or U1411 (N_1411,In_803,In_679);
and U1412 (N_1412,In_822,In_490);
or U1413 (N_1413,In_72,In_927);
nand U1414 (N_1414,In_1104,In_1000);
or U1415 (N_1415,In_1454,In_609);
or U1416 (N_1416,In_763,In_319);
or U1417 (N_1417,In_1277,In_1387);
xor U1418 (N_1418,In_1496,In_1168);
xnor U1419 (N_1419,In_1485,In_112);
and U1420 (N_1420,In_496,In_925);
nor U1421 (N_1421,In_263,In_662);
and U1422 (N_1422,In_679,In_910);
or U1423 (N_1423,In_902,In_711);
and U1424 (N_1424,In_888,In_695);
or U1425 (N_1425,In_242,In_138);
or U1426 (N_1426,In_368,In_513);
xor U1427 (N_1427,In_1268,In_708);
nor U1428 (N_1428,In_1009,In_1106);
nor U1429 (N_1429,In_671,In_730);
xor U1430 (N_1430,In_1253,In_1037);
nor U1431 (N_1431,In_1459,In_1130);
nand U1432 (N_1432,In_1312,In_899);
nor U1433 (N_1433,In_447,In_1377);
xor U1434 (N_1434,In_161,In_53);
xor U1435 (N_1435,In_1107,In_1319);
and U1436 (N_1436,In_184,In_100);
nand U1437 (N_1437,In_646,In_73);
or U1438 (N_1438,In_766,In_1094);
and U1439 (N_1439,In_1387,In_643);
nand U1440 (N_1440,In_339,In_539);
nand U1441 (N_1441,In_762,In_452);
nor U1442 (N_1442,In_1462,In_379);
or U1443 (N_1443,In_136,In_90);
or U1444 (N_1444,In_892,In_711);
or U1445 (N_1445,In_914,In_698);
nor U1446 (N_1446,In_63,In_19);
or U1447 (N_1447,In_476,In_597);
and U1448 (N_1448,In_1354,In_927);
nor U1449 (N_1449,In_450,In_367);
and U1450 (N_1450,In_722,In_1435);
xnor U1451 (N_1451,In_1069,In_832);
nor U1452 (N_1452,In_1088,In_1399);
nand U1453 (N_1453,In_142,In_172);
nor U1454 (N_1454,In_1391,In_377);
nor U1455 (N_1455,In_71,In_761);
and U1456 (N_1456,In_563,In_524);
nor U1457 (N_1457,In_1119,In_1184);
xor U1458 (N_1458,In_744,In_1148);
and U1459 (N_1459,In_503,In_445);
nand U1460 (N_1460,In_1007,In_729);
nand U1461 (N_1461,In_397,In_572);
or U1462 (N_1462,In_1179,In_772);
nor U1463 (N_1463,In_1047,In_125);
nor U1464 (N_1464,In_40,In_1224);
xnor U1465 (N_1465,In_943,In_1126);
or U1466 (N_1466,In_1264,In_1357);
xor U1467 (N_1467,In_636,In_1139);
nor U1468 (N_1468,In_377,In_413);
xnor U1469 (N_1469,In_1394,In_782);
nand U1470 (N_1470,In_494,In_799);
and U1471 (N_1471,In_1217,In_499);
nand U1472 (N_1472,In_515,In_533);
nor U1473 (N_1473,In_1300,In_1376);
or U1474 (N_1474,In_389,In_211);
xnor U1475 (N_1475,In_919,In_337);
xnor U1476 (N_1476,In_368,In_1044);
and U1477 (N_1477,In_1396,In_420);
and U1478 (N_1478,In_1453,In_1329);
and U1479 (N_1479,In_842,In_1068);
xnor U1480 (N_1480,In_977,In_1062);
or U1481 (N_1481,In_653,In_91);
xnor U1482 (N_1482,In_457,In_1343);
xnor U1483 (N_1483,In_577,In_801);
or U1484 (N_1484,In_951,In_407);
or U1485 (N_1485,In_799,In_1370);
nand U1486 (N_1486,In_1118,In_774);
xnor U1487 (N_1487,In_228,In_406);
and U1488 (N_1488,In_288,In_280);
nand U1489 (N_1489,In_672,In_180);
xnor U1490 (N_1490,In_51,In_500);
and U1491 (N_1491,In_396,In_751);
and U1492 (N_1492,In_1441,In_810);
or U1493 (N_1493,In_385,In_1492);
nor U1494 (N_1494,In_603,In_1116);
nand U1495 (N_1495,In_1102,In_966);
xor U1496 (N_1496,In_227,In_769);
nand U1497 (N_1497,In_524,In_420);
and U1498 (N_1498,In_270,In_1416);
or U1499 (N_1499,In_273,In_952);
xnor U1500 (N_1500,N_305,N_515);
nand U1501 (N_1501,N_899,N_246);
nand U1502 (N_1502,N_284,N_248);
or U1503 (N_1503,N_429,N_718);
nor U1504 (N_1504,N_117,N_20);
nand U1505 (N_1505,N_894,N_462);
and U1506 (N_1506,N_957,N_1142);
or U1507 (N_1507,N_453,N_1354);
and U1508 (N_1508,N_1397,N_1026);
and U1509 (N_1509,N_714,N_1366);
or U1510 (N_1510,N_1433,N_1144);
or U1511 (N_1511,N_567,N_26);
xor U1512 (N_1512,N_177,N_1136);
and U1513 (N_1513,N_167,N_1118);
nand U1514 (N_1514,N_1303,N_766);
and U1515 (N_1515,N_1452,N_1025);
nand U1516 (N_1516,N_1086,N_962);
and U1517 (N_1517,N_858,N_1313);
or U1518 (N_1518,N_1199,N_768);
nand U1519 (N_1519,N_39,N_586);
and U1520 (N_1520,N_611,N_1390);
or U1521 (N_1521,N_1154,N_1063);
nor U1522 (N_1522,N_223,N_650);
or U1523 (N_1523,N_116,N_469);
or U1524 (N_1524,N_1043,N_1329);
or U1525 (N_1525,N_985,N_696);
nand U1526 (N_1526,N_1128,N_760);
or U1527 (N_1527,N_1445,N_986);
nor U1528 (N_1528,N_1141,N_336);
nor U1529 (N_1529,N_633,N_658);
nand U1530 (N_1530,N_511,N_813);
xor U1531 (N_1531,N_1006,N_1114);
and U1532 (N_1532,N_48,N_1258);
xor U1533 (N_1533,N_761,N_695);
and U1534 (N_1534,N_369,N_131);
or U1535 (N_1535,N_218,N_464);
nor U1536 (N_1536,N_1339,N_509);
nor U1537 (N_1537,N_1391,N_45);
xor U1538 (N_1538,N_876,N_1442);
xor U1539 (N_1539,N_179,N_1426);
xnor U1540 (N_1540,N_1305,N_428);
xnor U1541 (N_1541,N_1315,N_1472);
nor U1542 (N_1542,N_406,N_954);
or U1543 (N_1543,N_543,N_328);
and U1544 (N_1544,N_582,N_783);
or U1545 (N_1545,N_1069,N_1330);
or U1546 (N_1546,N_295,N_114);
and U1547 (N_1547,N_735,N_44);
nand U1548 (N_1548,N_1230,N_913);
and U1549 (N_1549,N_934,N_495);
and U1550 (N_1550,N_202,N_351);
xnor U1551 (N_1551,N_533,N_1236);
nand U1552 (N_1552,N_700,N_545);
xor U1553 (N_1553,N_1471,N_615);
nand U1554 (N_1554,N_657,N_212);
nand U1555 (N_1555,N_1115,N_589);
xnor U1556 (N_1556,N_283,N_1402);
nor U1557 (N_1557,N_1215,N_447);
xor U1558 (N_1558,N_332,N_1244);
nor U1559 (N_1559,N_1399,N_1385);
and U1560 (N_1560,N_775,N_301);
or U1561 (N_1561,N_1166,N_1485);
xor U1562 (N_1562,N_590,N_1148);
and U1563 (N_1563,N_1239,N_1386);
or U1564 (N_1564,N_414,N_879);
or U1565 (N_1565,N_163,N_949);
xor U1566 (N_1566,N_149,N_866);
nor U1567 (N_1567,N_877,N_747);
nor U1568 (N_1568,N_408,N_239);
nor U1569 (N_1569,N_420,N_1029);
or U1570 (N_1570,N_190,N_1207);
xnor U1571 (N_1571,N_1080,N_532);
nor U1572 (N_1572,N_551,N_952);
and U1573 (N_1573,N_180,N_267);
nand U1574 (N_1574,N_1159,N_405);
or U1575 (N_1575,N_882,N_561);
nand U1576 (N_1576,N_726,N_152);
xnor U1577 (N_1577,N_1035,N_519);
and U1578 (N_1578,N_878,N_651);
and U1579 (N_1579,N_1356,N_591);
or U1580 (N_1580,N_455,N_963);
or U1581 (N_1581,N_1211,N_374);
xnor U1582 (N_1582,N_965,N_702);
nor U1583 (N_1583,N_855,N_1235);
xor U1584 (N_1584,N_1217,N_1297);
and U1585 (N_1585,N_850,N_898);
nor U1586 (N_1586,N_132,N_268);
nor U1587 (N_1587,N_819,N_1374);
or U1588 (N_1588,N_839,N_194);
xnor U1589 (N_1589,N_1444,N_347);
nor U1590 (N_1590,N_778,N_397);
nor U1591 (N_1591,N_193,N_1285);
xnor U1592 (N_1592,N_412,N_1441);
xnor U1593 (N_1593,N_883,N_925);
nand U1594 (N_1594,N_1430,N_440);
nand U1595 (N_1595,N_1284,N_1240);
or U1596 (N_1596,N_1034,N_55);
nand U1597 (N_1597,N_300,N_477);
xnor U1598 (N_1598,N_1321,N_981);
nand U1599 (N_1599,N_227,N_1074);
or U1600 (N_1600,N_1406,N_181);
nand U1601 (N_1601,N_1047,N_265);
xnor U1602 (N_1602,N_786,N_376);
nor U1603 (N_1603,N_597,N_296);
or U1604 (N_1604,N_365,N_1408);
and U1605 (N_1605,N_30,N_262);
nor U1606 (N_1606,N_388,N_998);
xor U1607 (N_1607,N_1476,N_1295);
nor U1608 (N_1608,N_504,N_610);
xor U1609 (N_1609,N_1463,N_638);
nor U1610 (N_1610,N_356,N_1044);
nor U1611 (N_1611,N_780,N_238);
and U1612 (N_1612,N_929,N_410);
or U1613 (N_1613,N_708,N_1322);
nand U1614 (N_1614,N_770,N_587);
xor U1615 (N_1615,N_627,N_1486);
and U1616 (N_1616,N_1113,N_970);
nor U1617 (N_1617,N_662,N_531);
nor U1618 (N_1618,N_215,N_236);
nor U1619 (N_1619,N_1296,N_359);
nor U1620 (N_1620,N_1362,N_1394);
or U1621 (N_1621,N_632,N_1131);
or U1622 (N_1622,N_968,N_1410);
nand U1623 (N_1623,N_1060,N_422);
nand U1624 (N_1624,N_115,N_739);
and U1625 (N_1625,N_33,N_1010);
xnor U1626 (N_1626,N_1096,N_489);
xor U1627 (N_1627,N_844,N_1382);
and U1628 (N_1628,N_1238,N_886);
nand U1629 (N_1629,N_1138,N_903);
nand U1630 (N_1630,N_123,N_1245);
or U1631 (N_1631,N_908,N_105);
and U1632 (N_1632,N_624,N_1260);
and U1633 (N_1633,N_421,N_1040);
or U1634 (N_1634,N_643,N_917);
nor U1635 (N_1635,N_1254,N_921);
and U1636 (N_1636,N_1400,N_237);
nand U1637 (N_1637,N_357,N_698);
nor U1638 (N_1638,N_546,N_6);
or U1639 (N_1639,N_1048,N_743);
or U1640 (N_1640,N_1101,N_1451);
nor U1641 (N_1641,N_948,N_806);
nor U1642 (N_1642,N_1482,N_1023);
nor U1643 (N_1643,N_602,N_217);
xor U1644 (N_1644,N_373,N_1028);
nor U1645 (N_1645,N_555,N_541);
nor U1646 (N_1646,N_85,N_220);
xor U1647 (N_1647,N_1094,N_1062);
or U1648 (N_1648,N_128,N_1164);
nor U1649 (N_1649,N_297,N_1017);
nor U1650 (N_1650,N_690,N_1355);
or U1651 (N_1651,N_942,N_840);
or U1652 (N_1652,N_1484,N_481);
nand U1653 (N_1653,N_1090,N_787);
xnor U1654 (N_1654,N_506,N_1001);
xnor U1655 (N_1655,N_463,N_1181);
xnor U1656 (N_1656,N_199,N_1342);
nor U1657 (N_1657,N_1462,N_1294);
nor U1658 (N_1658,N_1083,N_607);
or U1659 (N_1659,N_185,N_725);
and U1660 (N_1660,N_1016,N_992);
or U1661 (N_1661,N_1450,N_1461);
xnor U1662 (N_1662,N_1468,N_130);
xor U1663 (N_1663,N_293,N_1184);
nand U1664 (N_1664,N_1020,N_315);
nor U1665 (N_1665,N_756,N_121);
nor U1666 (N_1666,N_868,N_314);
xnor U1667 (N_1667,N_1070,N_748);
or U1668 (N_1668,N_1483,N_1425);
xnor U1669 (N_1669,N_694,N_895);
nand U1670 (N_1670,N_316,N_873);
xnor U1671 (N_1671,N_794,N_1380);
xor U1672 (N_1672,N_192,N_1073);
nand U1673 (N_1673,N_922,N_528);
xnor U1674 (N_1674,N_1370,N_1229);
or U1675 (N_1675,N_678,N_1099);
and U1676 (N_1676,N_62,N_919);
xnor U1677 (N_1677,N_345,N_1378);
xnor U1678 (N_1678,N_272,N_460);
xor U1679 (N_1679,N_1171,N_1013);
or U1680 (N_1680,N_67,N_1190);
nor U1681 (N_1681,N_399,N_856);
nor U1682 (N_1682,N_111,N_618);
nor U1683 (N_1683,N_1210,N_427);
nor U1684 (N_1684,N_91,N_782);
nand U1685 (N_1685,N_859,N_604);
or U1686 (N_1686,N_752,N_941);
or U1687 (N_1687,N_304,N_423);
and U1688 (N_1688,N_892,N_285);
and U1689 (N_1689,N_1333,N_995);
nand U1690 (N_1690,N_955,N_1498);
nor U1691 (N_1691,N_1267,N_1404);
xor U1692 (N_1692,N_1431,N_1328);
xnor U1693 (N_1693,N_1122,N_57);
nand U1694 (N_1694,N_1352,N_523);
nand U1695 (N_1695,N_1496,N_885);
and U1696 (N_1696,N_1237,N_1111);
nor U1697 (N_1697,N_500,N_186);
or U1698 (N_1698,N_1107,N_11);
nor U1699 (N_1699,N_70,N_1130);
and U1700 (N_1700,N_645,N_540);
nand U1701 (N_1701,N_1156,N_1396);
and U1702 (N_1702,N_1413,N_796);
xor U1703 (N_1703,N_971,N_902);
and U1704 (N_1704,N_683,N_1266);
or U1705 (N_1705,N_1289,N_1341);
or U1706 (N_1706,N_671,N_975);
nand U1707 (N_1707,N_652,N_936);
nand U1708 (N_1708,N_1071,N_709);
and U1709 (N_1709,N_253,N_503);
xnor U1710 (N_1710,N_884,N_92);
nor U1711 (N_1711,N_795,N_631);
xnor U1712 (N_1712,N_165,N_150);
xnor U1713 (N_1713,N_807,N_145);
or U1714 (N_1714,N_355,N_1435);
nor U1715 (N_1715,N_584,N_1155);
nand U1716 (N_1716,N_572,N_299);
or U1717 (N_1717,N_1160,N_380);
nand U1718 (N_1718,N_1189,N_1493);
xnor U1719 (N_1719,N_349,N_309);
and U1720 (N_1720,N_334,N_209);
nor U1721 (N_1721,N_918,N_790);
nand U1722 (N_1722,N_901,N_1273);
and U1723 (N_1723,N_1310,N_1334);
nand U1724 (N_1724,N_15,N_153);
or U1725 (N_1725,N_1436,N_415);
nor U1726 (N_1726,N_684,N_1286);
xor U1727 (N_1727,N_433,N_802);
xnor U1728 (N_1728,N_581,N_213);
nor U1729 (N_1729,N_577,N_721);
or U1730 (N_1730,N_472,N_909);
or U1731 (N_1731,N_1077,N_784);
nand U1732 (N_1732,N_1124,N_53);
and U1733 (N_1733,N_1012,N_211);
nand U1734 (N_1734,N_1255,N_1403);
or U1735 (N_1735,N_291,N_874);
and U1736 (N_1736,N_573,N_751);
or U1737 (N_1737,N_1093,N_490);
nand U1738 (N_1738,N_1150,N_758);
and U1739 (N_1739,N_817,N_811);
or U1740 (N_1740,N_1458,N_978);
or U1741 (N_1741,N_1277,N_665);
or U1742 (N_1742,N_1401,N_197);
nand U1743 (N_1743,N_1018,N_976);
and U1744 (N_1744,N_980,N_263);
or U1745 (N_1745,N_446,N_1203);
nor U1746 (N_1746,N_703,N_303);
nor U1747 (N_1747,N_323,N_808);
nand U1748 (N_1748,N_842,N_852);
nor U1749 (N_1749,N_711,N_1068);
nand U1750 (N_1750,N_1358,N_73);
nand U1751 (N_1751,N_1337,N_1188);
nor U1752 (N_1752,N_256,N_413);
xnor U1753 (N_1753,N_548,N_505);
and U1754 (N_1754,N_734,N_64);
and U1755 (N_1755,N_84,N_867);
xor U1756 (N_1756,N_1216,N_547);
nand U1757 (N_1757,N_241,N_544);
or U1758 (N_1758,N_1365,N_1191);
nor U1759 (N_1759,N_372,N_516);
xnor U1760 (N_1760,N_810,N_745);
nor U1761 (N_1761,N_754,N_1357);
or U1762 (N_1762,N_1422,N_1209);
xnor U1763 (N_1763,N_550,N_527);
nand U1764 (N_1764,N_1293,N_1446);
and U1765 (N_1765,N_763,N_1416);
nand U1766 (N_1766,N_1106,N_996);
nor U1767 (N_1767,N_17,N_950);
nor U1768 (N_1768,N_1088,N_1299);
or U1769 (N_1769,N_442,N_319);
and U1770 (N_1770,N_933,N_1234);
xor U1771 (N_1771,N_1252,N_322);
nand U1772 (N_1772,N_367,N_109);
and U1773 (N_1773,N_308,N_1281);
xor U1774 (N_1774,N_475,N_189);
xnor U1775 (N_1775,N_843,N_360);
nand U1776 (N_1776,N_277,N_705);
nor U1777 (N_1777,N_287,N_333);
nor U1778 (N_1778,N_915,N_1173);
or U1779 (N_1779,N_71,N_822);
or U1780 (N_1780,N_375,N_1499);
xor U1781 (N_1781,N_914,N_330);
or U1782 (N_1782,N_497,N_385);
or U1783 (N_1783,N_689,N_1434);
and U1784 (N_1784,N_744,N_499);
nand U1785 (N_1785,N_348,N_767);
xnor U1786 (N_1786,N_788,N_340);
nor U1787 (N_1787,N_1112,N_1492);
or U1788 (N_1788,N_571,N_459);
nor U1789 (N_1789,N_264,N_321);
nor U1790 (N_1790,N_835,N_967);
nand U1791 (N_1791,N_655,N_1162);
or U1792 (N_1792,N_1343,N_445);
nor U1793 (N_1793,N_59,N_487);
nor U1794 (N_1794,N_77,N_1307);
and U1795 (N_1795,N_142,N_25);
nand U1796 (N_1796,N_729,N_1041);
nor U1797 (N_1797,N_753,N_520);
xnor U1798 (N_1798,N_1327,N_1146);
or U1799 (N_1799,N_609,N_588);
xnor U1800 (N_1800,N_1227,N_552);
xor U1801 (N_1801,N_812,N_1291);
nand U1802 (N_1802,N_1007,N_1477);
xnor U1803 (N_1803,N_723,N_1376);
nand U1804 (N_1804,N_622,N_654);
nor U1805 (N_1805,N_605,N_1172);
or U1806 (N_1806,N_219,N_1490);
nand U1807 (N_1807,N_95,N_361);
or U1808 (N_1808,N_1097,N_1470);
nand U1809 (N_1809,N_1000,N_260);
nor U1810 (N_1810,N_151,N_1176);
and U1811 (N_1811,N_498,N_419);
or U1812 (N_1812,N_827,N_851);
nand U1813 (N_1813,N_982,N_493);
or U1814 (N_1814,N_774,N_746);
xnor U1815 (N_1815,N_456,N_668);
nor U1816 (N_1816,N_5,N_742);
nand U1817 (N_1817,N_849,N_178);
or U1818 (N_1818,N_1423,N_997);
or U1819 (N_1819,N_424,N_407);
nor U1820 (N_1820,N_274,N_1116);
nor U1821 (N_1821,N_1186,N_88);
and U1822 (N_1822,N_988,N_1393);
or U1823 (N_1823,N_1479,N_89);
nand U1824 (N_1824,N_973,N_1046);
nand U1825 (N_1825,N_722,N_49);
nor U1826 (N_1826,N_1497,N_1197);
or U1827 (N_1827,N_635,N_906);
xor U1828 (N_1828,N_1361,N_101);
nand U1829 (N_1829,N_554,N_1031);
nand U1830 (N_1830,N_104,N_1491);
nand U1831 (N_1831,N_1271,N_66);
and U1832 (N_1832,N_1324,N_155);
nand U1833 (N_1833,N_1021,N_1250);
nand U1834 (N_1834,N_1087,N_1373);
and U1835 (N_1835,N_1264,N_1466);
nor U1836 (N_1836,N_344,N_1282);
or U1837 (N_1837,N_231,N_1249);
or U1838 (N_1838,N_430,N_232);
nor U1839 (N_1839,N_1481,N_118);
xnor U1840 (N_1840,N_821,N_1449);
or U1841 (N_1841,N_928,N_660);
xnor U1842 (N_1842,N_273,N_598);
and U1843 (N_1843,N_1359,N_1056);
xnor U1844 (N_1844,N_1169,N_1248);
and U1845 (N_1845,N_1200,N_1312);
and U1846 (N_1846,N_994,N_1439);
or U1847 (N_1847,N_1398,N_1495);
nor U1848 (N_1848,N_1121,N_869);
nand U1849 (N_1849,N_18,N_364);
nor U1850 (N_1850,N_1054,N_1278);
or U1851 (N_1851,N_1195,N_960);
or U1852 (N_1852,N_1015,N_110);
xor U1853 (N_1853,N_280,N_492);
and U1854 (N_1854,N_670,N_682);
nor U1855 (N_1855,N_140,N_486);
nand U1856 (N_1856,N_452,N_1432);
or U1857 (N_1857,N_688,N_522);
nand U1858 (N_1858,N_730,N_964);
nor U1859 (N_1859,N_19,N_259);
xnor U1860 (N_1860,N_488,N_1100);
xnor U1861 (N_1861,N_989,N_1319);
xor U1862 (N_1862,N_37,N_944);
or U1863 (N_1863,N_93,N_134);
or U1864 (N_1864,N_1182,N_52);
and U1865 (N_1865,N_1135,N_815);
and U1866 (N_1866,N_324,N_1102);
and U1867 (N_1867,N_1226,N_393);
nor U1868 (N_1868,N_182,N_210);
and U1869 (N_1869,N_983,N_496);
or U1870 (N_1870,N_932,N_1022);
nand U1871 (N_1871,N_733,N_628);
nor U1872 (N_1872,N_510,N_379);
or U1873 (N_1873,N_757,N_31);
nand U1874 (N_1874,N_1261,N_203);
nand U1875 (N_1875,N_853,N_436);
nand U1876 (N_1876,N_148,N_1473);
nor U1877 (N_1877,N_366,N_243);
or U1878 (N_1878,N_4,N_828);
nand U1879 (N_1879,N_630,N_1194);
xor U1880 (N_1880,N_378,N_426);
nor U1881 (N_1881,N_521,N_809);
and U1882 (N_1882,N_776,N_1340);
and U1883 (N_1883,N_390,N_720);
and U1884 (N_1884,N_371,N_1288);
nor U1885 (N_1885,N_1231,N_535);
nand U1886 (N_1886,N_1089,N_1371);
nor U1887 (N_1887,N_846,N_1387);
nor U1888 (N_1888,N_1405,N_8);
nand U1889 (N_1889,N_1233,N_1427);
nand U1890 (N_1890,N_438,N_1272);
or U1891 (N_1891,N_953,N_1045);
and U1892 (N_1892,N_1201,N_434);
nand U1893 (N_1893,N_1030,N_1268);
xor U1894 (N_1894,N_838,N_889);
nor U1895 (N_1895,N_1335,N_1318);
and U1896 (N_1896,N_391,N_599);
nand U1897 (N_1897,N_732,N_765);
and U1898 (N_1898,N_352,N_1407);
nand U1899 (N_1899,N_943,N_749);
and U1900 (N_1900,N_1208,N_1117);
nand U1901 (N_1901,N_1424,N_613);
nand U1902 (N_1902,N_1262,N_12);
xor U1903 (N_1903,N_875,N_482);
nor U1904 (N_1904,N_266,N_1153);
or U1905 (N_1905,N_1306,N_900);
or U1906 (N_1906,N_1152,N_830);
xor U1907 (N_1907,N_480,N_1187);
xnor U1908 (N_1908,N_1345,N_289);
nor U1909 (N_1909,N_890,N_1379);
nor U1910 (N_1910,N_789,N_229);
and U1911 (N_1911,N_108,N_454);
xor U1912 (N_1912,N_564,N_558);
xor U1913 (N_1913,N_320,N_1265);
nor U1914 (N_1914,N_579,N_617);
nand U1915 (N_1915,N_575,N_1253);
or U1916 (N_1916,N_649,N_206);
or U1917 (N_1917,N_777,N_98);
xnor U1918 (N_1918,N_1465,N_76);
xor U1919 (N_1919,N_36,N_1129);
nor U1920 (N_1920,N_741,N_619);
nand U1921 (N_1921,N_468,N_461);
nand U1922 (N_1922,N_930,N_78);
and U1923 (N_1923,N_1447,N_1437);
nand U1924 (N_1924,N_354,N_51);
or U1925 (N_1925,N_1414,N_162);
xnor U1926 (N_1926,N_553,N_634);
xnor U1927 (N_1927,N_1331,N_68);
nor U1928 (N_1928,N_513,N_724);
and U1929 (N_1929,N_431,N_1);
xnor U1930 (N_1930,N_805,N_43);
and U1931 (N_1931,N_443,N_126);
and U1932 (N_1932,N_1140,N_42);
nor U1933 (N_1933,N_1421,N_278);
nand U1934 (N_1934,N_1457,N_143);
nand U1935 (N_1935,N_1360,N_1344);
or U1936 (N_1936,N_100,N_841);
or U1937 (N_1937,N_1287,N_1158);
nor U1938 (N_1938,N_1232,N_1332);
or U1939 (N_1939,N_159,N_254);
xor U1940 (N_1940,N_501,N_946);
nor U1941 (N_1941,N_82,N_834);
or U1942 (N_1942,N_565,N_559);
nand U1943 (N_1943,N_1065,N_1078);
nand U1944 (N_1944,N_977,N_329);
xor U1945 (N_1945,N_1456,N_603);
or U1946 (N_1946,N_484,N_905);
and U1947 (N_1947,N_1145,N_401);
and U1948 (N_1948,N_233,N_294);
nor U1949 (N_1949,N_1301,N_312);
xor U1950 (N_1950,N_910,N_41);
nand U1951 (N_1951,N_158,N_1304);
xnor U1952 (N_1952,N_276,N_106);
nor U1953 (N_1953,N_1348,N_83);
and U1954 (N_1954,N_80,N_642);
nor U1955 (N_1955,N_993,N_666);
xor U1956 (N_1956,N_647,N_1459);
xor U1957 (N_1957,N_313,N_325);
nand U1958 (N_1958,N_1292,N_825);
xnor U1959 (N_1959,N_699,N_172);
and U1960 (N_1960,N_1347,N_1383);
or U1961 (N_1961,N_1049,N_269);
or U1962 (N_1962,N_1363,N_661);
nand U1963 (N_1963,N_823,N_1196);
and U1964 (N_1964,N_931,N_940);
or U1965 (N_1965,N_974,N_465);
or U1966 (N_1966,N_959,N_1147);
xor U1967 (N_1967,N_637,N_69);
and U1968 (N_1968,N_570,N_1257);
nand U1969 (N_1969,N_417,N_350);
nand U1970 (N_1970,N_279,N_1126);
xor U1971 (N_1971,N_920,N_1338);
and U1972 (N_1972,N_1066,N_1179);
and U1973 (N_1973,N_831,N_395);
nand U1974 (N_1974,N_317,N_1005);
nor U1975 (N_1975,N_338,N_341);
nand U1976 (N_1976,N_772,N_402);
and U1977 (N_1977,N_127,N_1350);
nor U1978 (N_1978,N_1036,N_1420);
xnor U1979 (N_1979,N_466,N_257);
nor U1980 (N_1980,N_737,N_1467);
nand U1981 (N_1981,N_435,N_96);
xnor U1982 (N_1982,N_801,N_563);
xor U1983 (N_1983,N_673,N_409);
nor U1984 (N_1984,N_1185,N_74);
nand U1985 (N_1985,N_1480,N_1019);
or U1986 (N_1986,N_1346,N_1027);
or U1987 (N_1987,N_1443,N_23);
xnor U1988 (N_1988,N_956,N_170);
nor U1989 (N_1989,N_1180,N_904);
xnor U1990 (N_1990,N_249,N_1193);
xnor U1991 (N_1991,N_814,N_537);
or U1992 (N_1992,N_75,N_224);
xor U1993 (N_1993,N_411,N_1137);
and U1994 (N_1994,N_534,N_594);
or U1995 (N_1995,N_255,N_458);
nor U1996 (N_1996,N_1108,N_1218);
nor U1997 (N_1997,N_383,N_1161);
nor U1998 (N_1998,N_24,N_389);
xnor U1999 (N_1999,N_384,N_691);
xnor U2000 (N_2000,N_1259,N_394);
nor U2001 (N_2001,N_1003,N_871);
or U2002 (N_2002,N_112,N_854);
xnor U2003 (N_2003,N_1214,N_228);
or U2004 (N_2004,N_120,N_595);
and U2005 (N_2005,N_1325,N_508);
nand U2006 (N_2006,N_353,N_494);
and U2007 (N_2007,N_755,N_154);
or U2008 (N_2008,N_240,N_1064);
xor U2009 (N_2009,N_425,N_1448);
nor U2010 (N_2010,N_958,N_61);
nor U2011 (N_2011,N_14,N_578);
and U2012 (N_2012,N_891,N_583);
and U2013 (N_2013,N_518,N_38);
nor U2014 (N_2014,N_1082,N_693);
xor U2015 (N_2015,N_614,N_3);
xor U2016 (N_2016,N_214,N_1228);
nand U2017 (N_2017,N_870,N_169);
nand U2018 (N_2018,N_1168,N_663);
or U2019 (N_2019,N_1167,N_569);
or U2020 (N_2020,N_512,N_1004);
nand U2021 (N_2021,N_99,N_1220);
xor U2022 (N_2022,N_1474,N_972);
xor U2023 (N_2023,N_1095,N_1454);
nand U2024 (N_2024,N_524,N_1219);
and U2025 (N_2025,N_225,N_863);
xnor U2026 (N_2026,N_592,N_147);
or U2027 (N_2027,N_636,N_833);
xnor U2028 (N_2028,N_750,N_864);
and U2029 (N_2029,N_1308,N_34);
or U2030 (N_2030,N_593,N_1388);
and U2031 (N_2031,N_1061,N_113);
or U2032 (N_2032,N_222,N_1139);
xnor U2033 (N_2033,N_912,N_927);
and U2034 (N_2034,N_200,N_1143);
nor U2035 (N_2035,N_1311,N_847);
nor U2036 (N_2036,N_1478,N_392);
or U2037 (N_2037,N_1269,N_32);
or U2038 (N_2038,N_1320,N_728);
nand U2039 (N_2039,N_188,N_740);
or U2040 (N_2040,N_793,N_1464);
and U2041 (N_2041,N_207,N_362);
nor U2042 (N_2042,N_1453,N_1163);
and U2043 (N_2043,N_820,N_1165);
and U2044 (N_2044,N_470,N_1149);
xnor U2045 (N_2045,N_230,N_865);
or U2046 (N_2046,N_646,N_318);
nor U2047 (N_2047,N_861,N_1368);
xor U2048 (N_2048,N_377,N_887);
or U2049 (N_2049,N_1381,N_144);
nor U2050 (N_2050,N_990,N_13);
or U2051 (N_2051,N_173,N_0);
and U2052 (N_2052,N_736,N_400);
nor U2053 (N_2053,N_1058,N_596);
or U2054 (N_2054,N_125,N_418);
or U2055 (N_2055,N_1243,N_529);
nand U2056 (N_2056,N_1279,N_398);
or U2057 (N_2057,N_138,N_103);
nand U2058 (N_2058,N_439,N_764);
xor U2059 (N_2059,N_1314,N_327);
xnor U2060 (N_2060,N_1247,N_97);
nand U2061 (N_2061,N_343,N_1290);
or U2062 (N_2062,N_204,N_608);
and U2063 (N_2063,N_1395,N_692);
and U2064 (N_2064,N_358,N_916);
nand U2065 (N_2065,N_987,N_161);
and U2066 (N_2066,N_880,N_467);
or U2067 (N_2067,N_860,N_644);
xnor U2068 (N_2068,N_832,N_1489);
nor U2069 (N_2069,N_1081,N_800);
nand U2070 (N_2070,N_198,N_669);
or U2071 (N_2071,N_1052,N_680);
xor U2072 (N_2072,N_1174,N_281);
or U2073 (N_2073,N_687,N_382);
or U2074 (N_2074,N_195,N_1317);
nor U2075 (N_2075,N_22,N_1316);
xor U2076 (N_2076,N_261,N_1494);
xnor U2077 (N_2077,N_872,N_601);
and U2078 (N_2078,N_47,N_1372);
or U2079 (N_2079,N_79,N_40);
and U2080 (N_2080,N_781,N_136);
xor U2081 (N_2081,N_245,N_56);
nand U2082 (N_2082,N_1075,N_1119);
nor U2083 (N_2083,N_947,N_1067);
nand U2084 (N_2084,N_966,N_1011);
xor U2085 (N_2085,N_568,N_771);
nor U2086 (N_2086,N_1323,N_999);
and U2087 (N_2087,N_1033,N_1298);
or U2088 (N_2088,N_1091,N_370);
or U2089 (N_2089,N_244,N_542);
xor U2090 (N_2090,N_1302,N_474);
and U2091 (N_2091,N_1205,N_1475);
nand U2092 (N_2092,N_311,N_27);
nor U2093 (N_2093,N_122,N_616);
or U2094 (N_2094,N_574,N_160);
nand U2095 (N_2095,N_183,N_969);
xor U2096 (N_2096,N_1072,N_1024);
and U2097 (N_2097,N_271,N_1055);
nor U2098 (N_2098,N_1127,N_86);
or U2099 (N_2099,N_1170,N_707);
nand U2100 (N_2100,N_346,N_600);
xor U2101 (N_2101,N_710,N_1270);
or U2102 (N_2102,N_769,N_1224);
and U2103 (N_2103,N_137,N_1057);
and U2104 (N_2104,N_845,N_1120);
nor U2105 (N_2105,N_1418,N_664);
or U2106 (N_2106,N_386,N_896);
and U2107 (N_2107,N_335,N_483);
and U2108 (N_2108,N_205,N_81);
or U2109 (N_2109,N_29,N_1326);
xnor U2110 (N_2110,N_201,N_606);
nand U2111 (N_2111,N_926,N_252);
or U2112 (N_2112,N_234,N_298);
and U2113 (N_2113,N_826,N_1256);
nand U2114 (N_2114,N_798,N_677);
nand U2115 (N_2115,N_704,N_485);
nor U2116 (N_2116,N_797,N_621);
xnor U2117 (N_2117,N_888,N_258);
nor U2118 (N_2118,N_681,N_1039);
xor U2119 (N_2119,N_247,N_403);
nand U2120 (N_2120,N_717,N_1002);
or U2121 (N_2121,N_641,N_907);
nand U2122 (N_2122,N_857,N_1242);
nor U2123 (N_2123,N_1037,N_1412);
xor U2124 (N_2124,N_16,N_803);
and U2125 (N_2125,N_1275,N_1104);
nand U2126 (N_2126,N_837,N_897);
nand U2127 (N_2127,N_1336,N_404);
nor U2128 (N_2128,N_881,N_1300);
nand U2129 (N_2129,N_779,N_1051);
nand U2130 (N_2130,N_164,N_275);
xnor U2131 (N_2131,N_290,N_270);
nand U2132 (N_2132,N_1157,N_102);
or U2133 (N_2133,N_1438,N_1377);
xor U2134 (N_2134,N_762,N_107);
or U2135 (N_2135,N_727,N_1084);
nand U2136 (N_2136,N_525,N_1367);
nand U2137 (N_2137,N_242,N_938);
or U2138 (N_2138,N_381,N_984);
xnor U2139 (N_2139,N_816,N_712);
and U2140 (N_2140,N_1109,N_530);
nand U2141 (N_2141,N_1283,N_457);
nor U2142 (N_2142,N_235,N_715);
nand U2143 (N_2143,N_476,N_1079);
xor U2144 (N_2144,N_502,N_1183);
nand U2145 (N_2145,N_1419,N_1032);
nor U2146 (N_2146,N_28,N_94);
nor U2147 (N_2147,N_1411,N_58);
or U2148 (N_2148,N_1050,N_1309);
xnor U2149 (N_2149,N_639,N_368);
or U2150 (N_2150,N_507,N_679);
or U2151 (N_2151,N_1469,N_221);
nand U2152 (N_2152,N_1085,N_63);
or U2153 (N_2153,N_9,N_396);
nor U2154 (N_2154,N_437,N_1212);
nand U2155 (N_2155,N_286,N_716);
nor U2156 (N_2156,N_566,N_72);
or U2157 (N_2157,N_65,N_157);
nor U2158 (N_2158,N_135,N_1014);
nand U2159 (N_2159,N_342,N_893);
nand U2160 (N_2160,N_935,N_667);
xor U2161 (N_2161,N_625,N_836);
or U2162 (N_2162,N_307,N_191);
nand U2163 (N_2163,N_451,N_60);
or U2164 (N_2164,N_292,N_331);
nand U2165 (N_2165,N_706,N_623);
or U2166 (N_2166,N_1123,N_1384);
nor U2167 (N_2167,N_1246,N_829);
xnor U2168 (N_2168,N_174,N_1192);
nand U2169 (N_2169,N_1274,N_656);
nor U2170 (N_2170,N_562,N_556);
or U2171 (N_2171,N_626,N_791);
xnor U2172 (N_2172,N_924,N_1349);
and U2173 (N_2173,N_1206,N_1133);
and U2174 (N_2174,N_1455,N_10);
or U2175 (N_2175,N_1460,N_1132);
nor U2176 (N_2176,N_337,N_1178);
or U2177 (N_2177,N_824,N_1375);
xnor U2178 (N_2178,N_282,N_1134);
and U2179 (N_2179,N_302,N_585);
nor U2180 (N_2180,N_432,N_124);
or U2181 (N_2181,N_1221,N_686);
or U2182 (N_2182,N_2,N_251);
nand U2183 (N_2183,N_1105,N_685);
nand U2184 (N_2184,N_187,N_675);
nand U2185 (N_2185,N_580,N_1417);
and U2186 (N_2186,N_471,N_526);
nand U2187 (N_2187,N_1076,N_441);
nor U2188 (N_2188,N_738,N_473);
xnor U2189 (N_2189,N_1225,N_54);
xor U2190 (N_2190,N_560,N_156);
nor U2191 (N_2191,N_536,N_448);
nand U2192 (N_2192,N_1223,N_168);
xnor U2193 (N_2193,N_216,N_119);
nand U2194 (N_2194,N_1198,N_1369);
nor U2195 (N_2195,N_196,N_288);
nor U2196 (N_2196,N_719,N_991);
nand U2197 (N_2197,N_310,N_363);
xnor U2198 (N_2198,N_697,N_146);
xnor U2199 (N_2199,N_1222,N_1392);
xnor U2200 (N_2200,N_339,N_1241);
nor U2201 (N_2201,N_792,N_1151);
or U2202 (N_2202,N_818,N_759);
nand U2203 (N_2203,N_1059,N_416);
xnor U2204 (N_2204,N_1389,N_1098);
or U2205 (N_2205,N_862,N_961);
nor U2206 (N_2206,N_848,N_576);
xor U2207 (N_2207,N_612,N_640);
and U2208 (N_2208,N_133,N_1488);
or U2209 (N_2209,N_129,N_557);
xnor U2210 (N_2210,N_1110,N_444);
or U2211 (N_2211,N_166,N_1202);
nand U2212 (N_2212,N_676,N_1487);
xor U2213 (N_2213,N_923,N_1364);
or U2214 (N_2214,N_450,N_731);
nand U2215 (N_2215,N_937,N_804);
nand U2216 (N_2216,N_538,N_87);
or U2217 (N_2217,N_449,N_549);
nor U2218 (N_2218,N_620,N_939);
xor U2219 (N_2219,N_1008,N_46);
nand U2220 (N_2220,N_517,N_479);
or U2221 (N_2221,N_1092,N_1429);
or U2222 (N_2222,N_648,N_674);
xor U2223 (N_2223,N_306,N_1428);
or U2224 (N_2224,N_139,N_514);
and U2225 (N_2225,N_171,N_478);
nand U2226 (N_2226,N_911,N_659);
or U2227 (N_2227,N_945,N_1038);
xnor U2228 (N_2228,N_1103,N_1351);
nand U2229 (N_2229,N_176,N_1177);
nand U2230 (N_2230,N_1204,N_1009);
nor U2231 (N_2231,N_141,N_713);
nand U2232 (N_2232,N_979,N_184);
nor U2233 (N_2233,N_90,N_539);
nor U2234 (N_2234,N_21,N_35);
or U2235 (N_2235,N_1415,N_250);
or U2236 (N_2236,N_1280,N_226);
nor U2237 (N_2237,N_1175,N_1353);
or U2238 (N_2238,N_208,N_1213);
or U2239 (N_2239,N_799,N_1409);
and U2240 (N_2240,N_175,N_672);
nand U2241 (N_2241,N_1251,N_653);
nor U2242 (N_2242,N_1125,N_1440);
xnor U2243 (N_2243,N_50,N_491);
and U2244 (N_2244,N_1276,N_701);
and U2245 (N_2245,N_629,N_951);
and U2246 (N_2246,N_326,N_1263);
nand U2247 (N_2247,N_1042,N_7);
nor U2248 (N_2248,N_773,N_1053);
xor U2249 (N_2249,N_785,N_387);
nand U2250 (N_2250,N_1356,N_1120);
nor U2251 (N_2251,N_1260,N_1296);
and U2252 (N_2252,N_158,N_552);
xor U2253 (N_2253,N_487,N_464);
or U2254 (N_2254,N_317,N_452);
and U2255 (N_2255,N_1103,N_1174);
nand U2256 (N_2256,N_173,N_581);
xor U2257 (N_2257,N_1169,N_495);
xor U2258 (N_2258,N_1498,N_1102);
xor U2259 (N_2259,N_1336,N_1073);
xnor U2260 (N_2260,N_745,N_689);
nor U2261 (N_2261,N_291,N_1450);
nand U2262 (N_2262,N_1145,N_221);
and U2263 (N_2263,N_90,N_1371);
and U2264 (N_2264,N_1373,N_541);
nand U2265 (N_2265,N_818,N_957);
and U2266 (N_2266,N_1469,N_201);
nor U2267 (N_2267,N_923,N_1417);
nor U2268 (N_2268,N_561,N_50);
nand U2269 (N_2269,N_1063,N_649);
xor U2270 (N_2270,N_354,N_507);
and U2271 (N_2271,N_924,N_1438);
and U2272 (N_2272,N_1063,N_1021);
nand U2273 (N_2273,N_332,N_778);
and U2274 (N_2274,N_456,N_586);
and U2275 (N_2275,N_532,N_334);
and U2276 (N_2276,N_555,N_437);
nand U2277 (N_2277,N_971,N_802);
and U2278 (N_2278,N_1389,N_1433);
nand U2279 (N_2279,N_1484,N_1041);
or U2280 (N_2280,N_1044,N_670);
nand U2281 (N_2281,N_559,N_947);
nor U2282 (N_2282,N_1342,N_869);
and U2283 (N_2283,N_467,N_398);
xor U2284 (N_2284,N_387,N_233);
and U2285 (N_2285,N_117,N_1268);
and U2286 (N_2286,N_1069,N_443);
or U2287 (N_2287,N_1267,N_628);
and U2288 (N_2288,N_933,N_139);
nand U2289 (N_2289,N_28,N_1181);
nand U2290 (N_2290,N_895,N_587);
xnor U2291 (N_2291,N_255,N_819);
nand U2292 (N_2292,N_486,N_1264);
or U2293 (N_2293,N_372,N_224);
nand U2294 (N_2294,N_862,N_517);
xnor U2295 (N_2295,N_1308,N_525);
nor U2296 (N_2296,N_864,N_421);
nand U2297 (N_2297,N_452,N_86);
nand U2298 (N_2298,N_122,N_1476);
and U2299 (N_2299,N_1256,N_1205);
xor U2300 (N_2300,N_1150,N_731);
and U2301 (N_2301,N_1325,N_835);
xor U2302 (N_2302,N_546,N_483);
or U2303 (N_2303,N_519,N_882);
and U2304 (N_2304,N_386,N_624);
xnor U2305 (N_2305,N_282,N_126);
xnor U2306 (N_2306,N_1171,N_821);
xnor U2307 (N_2307,N_74,N_546);
nor U2308 (N_2308,N_1159,N_87);
and U2309 (N_2309,N_1257,N_450);
and U2310 (N_2310,N_936,N_465);
and U2311 (N_2311,N_1030,N_1049);
xnor U2312 (N_2312,N_292,N_849);
and U2313 (N_2313,N_95,N_412);
or U2314 (N_2314,N_560,N_1131);
and U2315 (N_2315,N_116,N_1047);
nor U2316 (N_2316,N_541,N_1495);
and U2317 (N_2317,N_617,N_550);
nand U2318 (N_2318,N_145,N_837);
xor U2319 (N_2319,N_390,N_345);
xor U2320 (N_2320,N_489,N_806);
nor U2321 (N_2321,N_798,N_916);
xnor U2322 (N_2322,N_564,N_597);
and U2323 (N_2323,N_274,N_771);
or U2324 (N_2324,N_230,N_1443);
or U2325 (N_2325,N_26,N_807);
nor U2326 (N_2326,N_356,N_595);
and U2327 (N_2327,N_1267,N_87);
nand U2328 (N_2328,N_407,N_952);
and U2329 (N_2329,N_1196,N_842);
nand U2330 (N_2330,N_237,N_1266);
or U2331 (N_2331,N_1139,N_254);
or U2332 (N_2332,N_329,N_519);
xor U2333 (N_2333,N_602,N_882);
or U2334 (N_2334,N_186,N_605);
xnor U2335 (N_2335,N_1186,N_638);
nand U2336 (N_2336,N_1113,N_220);
and U2337 (N_2337,N_832,N_1143);
nor U2338 (N_2338,N_84,N_1000);
xor U2339 (N_2339,N_345,N_850);
nor U2340 (N_2340,N_637,N_1193);
or U2341 (N_2341,N_1269,N_281);
nor U2342 (N_2342,N_1318,N_1148);
or U2343 (N_2343,N_1208,N_41);
nand U2344 (N_2344,N_1390,N_260);
or U2345 (N_2345,N_1072,N_1246);
nor U2346 (N_2346,N_944,N_1007);
or U2347 (N_2347,N_1175,N_918);
nor U2348 (N_2348,N_860,N_535);
and U2349 (N_2349,N_1124,N_830);
nor U2350 (N_2350,N_1485,N_347);
nor U2351 (N_2351,N_1429,N_1395);
nand U2352 (N_2352,N_1266,N_224);
nand U2353 (N_2353,N_1268,N_314);
xnor U2354 (N_2354,N_677,N_412);
and U2355 (N_2355,N_887,N_1083);
nor U2356 (N_2356,N_317,N_1345);
and U2357 (N_2357,N_1345,N_1143);
nor U2358 (N_2358,N_616,N_472);
and U2359 (N_2359,N_1118,N_848);
xnor U2360 (N_2360,N_340,N_10);
nor U2361 (N_2361,N_190,N_542);
or U2362 (N_2362,N_499,N_893);
and U2363 (N_2363,N_1024,N_1090);
nand U2364 (N_2364,N_241,N_1203);
or U2365 (N_2365,N_860,N_1203);
nor U2366 (N_2366,N_971,N_373);
nor U2367 (N_2367,N_707,N_1426);
and U2368 (N_2368,N_112,N_944);
nor U2369 (N_2369,N_446,N_60);
xor U2370 (N_2370,N_494,N_1386);
nor U2371 (N_2371,N_1243,N_1400);
nand U2372 (N_2372,N_907,N_932);
and U2373 (N_2373,N_678,N_1219);
or U2374 (N_2374,N_385,N_973);
nor U2375 (N_2375,N_488,N_687);
xnor U2376 (N_2376,N_587,N_151);
nand U2377 (N_2377,N_1411,N_124);
or U2378 (N_2378,N_1487,N_1191);
nor U2379 (N_2379,N_732,N_714);
and U2380 (N_2380,N_92,N_999);
or U2381 (N_2381,N_1452,N_333);
nor U2382 (N_2382,N_828,N_564);
nand U2383 (N_2383,N_653,N_55);
xnor U2384 (N_2384,N_1135,N_1366);
or U2385 (N_2385,N_641,N_1478);
nand U2386 (N_2386,N_1325,N_114);
nand U2387 (N_2387,N_1089,N_785);
xor U2388 (N_2388,N_1172,N_1167);
or U2389 (N_2389,N_1284,N_299);
and U2390 (N_2390,N_497,N_134);
or U2391 (N_2391,N_727,N_571);
nor U2392 (N_2392,N_352,N_582);
xor U2393 (N_2393,N_857,N_317);
or U2394 (N_2394,N_1117,N_1366);
nand U2395 (N_2395,N_688,N_1259);
xor U2396 (N_2396,N_1001,N_58);
nand U2397 (N_2397,N_357,N_152);
xnor U2398 (N_2398,N_991,N_433);
and U2399 (N_2399,N_50,N_237);
xor U2400 (N_2400,N_10,N_1438);
nor U2401 (N_2401,N_497,N_424);
nor U2402 (N_2402,N_911,N_799);
nor U2403 (N_2403,N_1128,N_28);
nand U2404 (N_2404,N_241,N_1153);
or U2405 (N_2405,N_999,N_1314);
or U2406 (N_2406,N_1230,N_416);
xnor U2407 (N_2407,N_952,N_496);
nand U2408 (N_2408,N_1379,N_795);
xor U2409 (N_2409,N_146,N_980);
or U2410 (N_2410,N_146,N_125);
nor U2411 (N_2411,N_94,N_143);
nor U2412 (N_2412,N_305,N_260);
or U2413 (N_2413,N_1147,N_375);
nor U2414 (N_2414,N_414,N_936);
nand U2415 (N_2415,N_332,N_1273);
nand U2416 (N_2416,N_1447,N_1);
and U2417 (N_2417,N_611,N_1483);
nor U2418 (N_2418,N_1039,N_139);
xor U2419 (N_2419,N_1241,N_690);
or U2420 (N_2420,N_327,N_127);
or U2421 (N_2421,N_1354,N_369);
xor U2422 (N_2422,N_1181,N_455);
nand U2423 (N_2423,N_912,N_1005);
nand U2424 (N_2424,N_1118,N_64);
nand U2425 (N_2425,N_453,N_182);
nand U2426 (N_2426,N_220,N_1134);
and U2427 (N_2427,N_327,N_1096);
nand U2428 (N_2428,N_70,N_217);
nand U2429 (N_2429,N_1118,N_68);
and U2430 (N_2430,N_5,N_968);
nand U2431 (N_2431,N_729,N_1050);
and U2432 (N_2432,N_902,N_450);
xnor U2433 (N_2433,N_622,N_1285);
nor U2434 (N_2434,N_1446,N_245);
and U2435 (N_2435,N_541,N_1340);
nand U2436 (N_2436,N_526,N_674);
or U2437 (N_2437,N_451,N_1020);
nand U2438 (N_2438,N_1236,N_283);
nand U2439 (N_2439,N_1435,N_1404);
or U2440 (N_2440,N_1398,N_1156);
nand U2441 (N_2441,N_1203,N_1333);
xor U2442 (N_2442,N_238,N_322);
xor U2443 (N_2443,N_958,N_754);
and U2444 (N_2444,N_981,N_225);
xnor U2445 (N_2445,N_749,N_886);
nand U2446 (N_2446,N_1442,N_327);
nor U2447 (N_2447,N_75,N_528);
and U2448 (N_2448,N_619,N_688);
nand U2449 (N_2449,N_1240,N_418);
and U2450 (N_2450,N_414,N_1448);
or U2451 (N_2451,N_1234,N_752);
nor U2452 (N_2452,N_1291,N_1223);
nand U2453 (N_2453,N_166,N_923);
or U2454 (N_2454,N_1320,N_391);
or U2455 (N_2455,N_1122,N_652);
or U2456 (N_2456,N_1440,N_1051);
nor U2457 (N_2457,N_768,N_1437);
and U2458 (N_2458,N_1042,N_1106);
and U2459 (N_2459,N_305,N_1194);
or U2460 (N_2460,N_709,N_919);
nor U2461 (N_2461,N_303,N_178);
xor U2462 (N_2462,N_279,N_727);
nand U2463 (N_2463,N_1114,N_43);
nand U2464 (N_2464,N_591,N_309);
nand U2465 (N_2465,N_248,N_153);
and U2466 (N_2466,N_456,N_1285);
nor U2467 (N_2467,N_913,N_1028);
xnor U2468 (N_2468,N_1356,N_1219);
nor U2469 (N_2469,N_1333,N_1099);
nor U2470 (N_2470,N_1304,N_650);
nor U2471 (N_2471,N_1034,N_1499);
nor U2472 (N_2472,N_993,N_1009);
nor U2473 (N_2473,N_1262,N_128);
xor U2474 (N_2474,N_998,N_1420);
nand U2475 (N_2475,N_852,N_41);
and U2476 (N_2476,N_371,N_288);
or U2477 (N_2477,N_405,N_782);
or U2478 (N_2478,N_409,N_1306);
or U2479 (N_2479,N_26,N_408);
nor U2480 (N_2480,N_760,N_999);
nor U2481 (N_2481,N_1051,N_995);
nand U2482 (N_2482,N_446,N_486);
nand U2483 (N_2483,N_197,N_409);
or U2484 (N_2484,N_943,N_856);
nor U2485 (N_2485,N_410,N_842);
and U2486 (N_2486,N_1320,N_1196);
or U2487 (N_2487,N_1369,N_113);
or U2488 (N_2488,N_926,N_1123);
nand U2489 (N_2489,N_641,N_204);
xor U2490 (N_2490,N_46,N_709);
nor U2491 (N_2491,N_874,N_208);
or U2492 (N_2492,N_1157,N_380);
and U2493 (N_2493,N_467,N_947);
and U2494 (N_2494,N_395,N_1331);
and U2495 (N_2495,N_249,N_43);
xor U2496 (N_2496,N_391,N_833);
nor U2497 (N_2497,N_681,N_133);
nand U2498 (N_2498,N_246,N_1121);
nor U2499 (N_2499,N_811,N_363);
nor U2500 (N_2500,N_10,N_881);
or U2501 (N_2501,N_1412,N_132);
nor U2502 (N_2502,N_962,N_1015);
and U2503 (N_2503,N_1205,N_1222);
xnor U2504 (N_2504,N_1164,N_36);
nand U2505 (N_2505,N_1025,N_857);
or U2506 (N_2506,N_1292,N_298);
or U2507 (N_2507,N_392,N_290);
and U2508 (N_2508,N_1464,N_925);
and U2509 (N_2509,N_996,N_1399);
xnor U2510 (N_2510,N_777,N_389);
or U2511 (N_2511,N_1297,N_1181);
nand U2512 (N_2512,N_56,N_1408);
or U2513 (N_2513,N_1472,N_86);
xnor U2514 (N_2514,N_1338,N_801);
nor U2515 (N_2515,N_14,N_990);
or U2516 (N_2516,N_72,N_1357);
nand U2517 (N_2517,N_295,N_86);
or U2518 (N_2518,N_149,N_169);
xor U2519 (N_2519,N_842,N_582);
nor U2520 (N_2520,N_1197,N_1024);
xnor U2521 (N_2521,N_372,N_256);
xor U2522 (N_2522,N_1330,N_594);
nand U2523 (N_2523,N_958,N_72);
nand U2524 (N_2524,N_691,N_1160);
and U2525 (N_2525,N_1376,N_1167);
nand U2526 (N_2526,N_833,N_619);
or U2527 (N_2527,N_1186,N_1087);
xor U2528 (N_2528,N_1185,N_923);
and U2529 (N_2529,N_192,N_1348);
xor U2530 (N_2530,N_109,N_903);
xnor U2531 (N_2531,N_985,N_196);
xnor U2532 (N_2532,N_355,N_911);
and U2533 (N_2533,N_1061,N_68);
nor U2534 (N_2534,N_369,N_146);
and U2535 (N_2535,N_824,N_1236);
nand U2536 (N_2536,N_1128,N_1396);
nor U2537 (N_2537,N_32,N_853);
xnor U2538 (N_2538,N_514,N_879);
and U2539 (N_2539,N_667,N_1245);
nor U2540 (N_2540,N_1171,N_921);
nor U2541 (N_2541,N_544,N_1109);
xor U2542 (N_2542,N_810,N_320);
or U2543 (N_2543,N_979,N_567);
xnor U2544 (N_2544,N_671,N_228);
nand U2545 (N_2545,N_248,N_1074);
or U2546 (N_2546,N_601,N_740);
xnor U2547 (N_2547,N_777,N_14);
xnor U2548 (N_2548,N_401,N_406);
nand U2549 (N_2549,N_21,N_1310);
nor U2550 (N_2550,N_1327,N_955);
nand U2551 (N_2551,N_913,N_536);
and U2552 (N_2552,N_1203,N_19);
nand U2553 (N_2553,N_203,N_457);
nand U2554 (N_2554,N_701,N_717);
xor U2555 (N_2555,N_125,N_77);
nand U2556 (N_2556,N_284,N_319);
and U2557 (N_2557,N_616,N_674);
and U2558 (N_2558,N_672,N_1367);
or U2559 (N_2559,N_105,N_1382);
and U2560 (N_2560,N_24,N_995);
and U2561 (N_2561,N_1375,N_135);
nand U2562 (N_2562,N_263,N_1041);
xnor U2563 (N_2563,N_389,N_855);
and U2564 (N_2564,N_753,N_437);
nor U2565 (N_2565,N_724,N_1134);
nor U2566 (N_2566,N_1058,N_139);
nand U2567 (N_2567,N_190,N_900);
or U2568 (N_2568,N_916,N_738);
and U2569 (N_2569,N_362,N_1219);
nor U2570 (N_2570,N_766,N_1147);
or U2571 (N_2571,N_1013,N_92);
nand U2572 (N_2572,N_1268,N_604);
xnor U2573 (N_2573,N_276,N_586);
nand U2574 (N_2574,N_277,N_30);
xor U2575 (N_2575,N_829,N_842);
and U2576 (N_2576,N_707,N_325);
xnor U2577 (N_2577,N_149,N_645);
xor U2578 (N_2578,N_1086,N_180);
nand U2579 (N_2579,N_1037,N_94);
nor U2580 (N_2580,N_127,N_242);
xor U2581 (N_2581,N_1485,N_514);
xnor U2582 (N_2582,N_1066,N_697);
nand U2583 (N_2583,N_1376,N_1491);
or U2584 (N_2584,N_707,N_319);
xor U2585 (N_2585,N_520,N_219);
or U2586 (N_2586,N_362,N_868);
xnor U2587 (N_2587,N_1215,N_792);
nor U2588 (N_2588,N_331,N_536);
nand U2589 (N_2589,N_907,N_66);
nand U2590 (N_2590,N_1265,N_1340);
nor U2591 (N_2591,N_113,N_1462);
nor U2592 (N_2592,N_1335,N_883);
nand U2593 (N_2593,N_1290,N_855);
and U2594 (N_2594,N_1268,N_403);
nand U2595 (N_2595,N_207,N_1169);
and U2596 (N_2596,N_94,N_95);
nor U2597 (N_2597,N_1350,N_1108);
or U2598 (N_2598,N_388,N_208);
and U2599 (N_2599,N_1162,N_191);
nand U2600 (N_2600,N_579,N_460);
or U2601 (N_2601,N_623,N_273);
or U2602 (N_2602,N_598,N_490);
xnor U2603 (N_2603,N_1069,N_679);
or U2604 (N_2604,N_1452,N_389);
or U2605 (N_2605,N_173,N_93);
xnor U2606 (N_2606,N_1139,N_741);
nor U2607 (N_2607,N_203,N_296);
nand U2608 (N_2608,N_819,N_758);
or U2609 (N_2609,N_349,N_308);
xnor U2610 (N_2610,N_235,N_173);
xnor U2611 (N_2611,N_100,N_80);
and U2612 (N_2612,N_807,N_1428);
nor U2613 (N_2613,N_401,N_25);
xor U2614 (N_2614,N_1166,N_1285);
nand U2615 (N_2615,N_403,N_436);
nand U2616 (N_2616,N_345,N_771);
nor U2617 (N_2617,N_974,N_1347);
nor U2618 (N_2618,N_229,N_251);
and U2619 (N_2619,N_774,N_370);
or U2620 (N_2620,N_1271,N_1029);
nand U2621 (N_2621,N_1447,N_1221);
xnor U2622 (N_2622,N_1183,N_565);
or U2623 (N_2623,N_400,N_1058);
or U2624 (N_2624,N_1154,N_1497);
nand U2625 (N_2625,N_920,N_505);
nand U2626 (N_2626,N_939,N_920);
or U2627 (N_2627,N_753,N_1046);
nor U2628 (N_2628,N_265,N_334);
nor U2629 (N_2629,N_251,N_885);
and U2630 (N_2630,N_134,N_152);
xnor U2631 (N_2631,N_1489,N_712);
nor U2632 (N_2632,N_956,N_370);
xnor U2633 (N_2633,N_1067,N_397);
or U2634 (N_2634,N_240,N_1182);
nor U2635 (N_2635,N_207,N_615);
or U2636 (N_2636,N_418,N_544);
nand U2637 (N_2637,N_758,N_1325);
nand U2638 (N_2638,N_539,N_1236);
or U2639 (N_2639,N_504,N_1317);
nor U2640 (N_2640,N_1195,N_1303);
nand U2641 (N_2641,N_828,N_1417);
and U2642 (N_2642,N_819,N_332);
and U2643 (N_2643,N_1435,N_673);
or U2644 (N_2644,N_847,N_1151);
and U2645 (N_2645,N_391,N_1);
and U2646 (N_2646,N_165,N_455);
nand U2647 (N_2647,N_975,N_526);
nor U2648 (N_2648,N_893,N_1093);
xnor U2649 (N_2649,N_1127,N_1410);
nor U2650 (N_2650,N_1393,N_678);
or U2651 (N_2651,N_278,N_200);
nor U2652 (N_2652,N_64,N_660);
nor U2653 (N_2653,N_219,N_186);
nand U2654 (N_2654,N_84,N_653);
nor U2655 (N_2655,N_753,N_192);
nor U2656 (N_2656,N_931,N_876);
nand U2657 (N_2657,N_294,N_1497);
nor U2658 (N_2658,N_1496,N_265);
nor U2659 (N_2659,N_862,N_20);
xnor U2660 (N_2660,N_626,N_1121);
and U2661 (N_2661,N_557,N_1123);
or U2662 (N_2662,N_436,N_777);
xor U2663 (N_2663,N_917,N_976);
nand U2664 (N_2664,N_151,N_387);
xnor U2665 (N_2665,N_149,N_946);
and U2666 (N_2666,N_337,N_1042);
xor U2667 (N_2667,N_407,N_1328);
nand U2668 (N_2668,N_820,N_1030);
xor U2669 (N_2669,N_1078,N_655);
xor U2670 (N_2670,N_1236,N_311);
nor U2671 (N_2671,N_158,N_1258);
nor U2672 (N_2672,N_1193,N_314);
nor U2673 (N_2673,N_550,N_1387);
xor U2674 (N_2674,N_149,N_1273);
or U2675 (N_2675,N_930,N_842);
nand U2676 (N_2676,N_458,N_879);
xnor U2677 (N_2677,N_546,N_1265);
nor U2678 (N_2678,N_863,N_293);
nand U2679 (N_2679,N_150,N_705);
nor U2680 (N_2680,N_361,N_55);
nor U2681 (N_2681,N_502,N_1366);
nand U2682 (N_2682,N_1204,N_1195);
or U2683 (N_2683,N_267,N_1302);
and U2684 (N_2684,N_1345,N_832);
and U2685 (N_2685,N_546,N_334);
xor U2686 (N_2686,N_621,N_300);
and U2687 (N_2687,N_60,N_1260);
nor U2688 (N_2688,N_187,N_614);
nor U2689 (N_2689,N_240,N_279);
or U2690 (N_2690,N_340,N_955);
or U2691 (N_2691,N_35,N_56);
nor U2692 (N_2692,N_819,N_810);
or U2693 (N_2693,N_957,N_801);
nor U2694 (N_2694,N_1184,N_1011);
and U2695 (N_2695,N_775,N_1338);
nor U2696 (N_2696,N_787,N_119);
and U2697 (N_2697,N_249,N_598);
nor U2698 (N_2698,N_578,N_1244);
nor U2699 (N_2699,N_1123,N_792);
or U2700 (N_2700,N_1496,N_410);
nor U2701 (N_2701,N_669,N_1021);
and U2702 (N_2702,N_362,N_436);
or U2703 (N_2703,N_1071,N_1340);
and U2704 (N_2704,N_561,N_1316);
xnor U2705 (N_2705,N_74,N_707);
or U2706 (N_2706,N_906,N_1235);
nor U2707 (N_2707,N_437,N_645);
or U2708 (N_2708,N_286,N_37);
or U2709 (N_2709,N_984,N_674);
and U2710 (N_2710,N_1115,N_723);
or U2711 (N_2711,N_1127,N_1382);
xnor U2712 (N_2712,N_296,N_899);
or U2713 (N_2713,N_712,N_181);
nand U2714 (N_2714,N_1304,N_658);
and U2715 (N_2715,N_947,N_1424);
xor U2716 (N_2716,N_109,N_488);
and U2717 (N_2717,N_306,N_391);
nand U2718 (N_2718,N_1495,N_1345);
and U2719 (N_2719,N_217,N_812);
xor U2720 (N_2720,N_562,N_1317);
nor U2721 (N_2721,N_480,N_857);
nor U2722 (N_2722,N_1434,N_435);
xor U2723 (N_2723,N_748,N_1314);
or U2724 (N_2724,N_70,N_1402);
or U2725 (N_2725,N_1029,N_1378);
and U2726 (N_2726,N_83,N_903);
nand U2727 (N_2727,N_720,N_1293);
nand U2728 (N_2728,N_452,N_973);
or U2729 (N_2729,N_1096,N_1419);
and U2730 (N_2730,N_365,N_1230);
or U2731 (N_2731,N_755,N_729);
nor U2732 (N_2732,N_1425,N_452);
nand U2733 (N_2733,N_707,N_256);
xnor U2734 (N_2734,N_71,N_674);
or U2735 (N_2735,N_1195,N_1134);
nand U2736 (N_2736,N_1072,N_193);
and U2737 (N_2737,N_744,N_693);
nor U2738 (N_2738,N_613,N_641);
and U2739 (N_2739,N_781,N_692);
or U2740 (N_2740,N_866,N_1286);
or U2741 (N_2741,N_1245,N_827);
xor U2742 (N_2742,N_206,N_339);
xnor U2743 (N_2743,N_1123,N_817);
nand U2744 (N_2744,N_331,N_1393);
and U2745 (N_2745,N_1320,N_857);
nor U2746 (N_2746,N_104,N_737);
and U2747 (N_2747,N_559,N_1033);
or U2748 (N_2748,N_635,N_154);
nor U2749 (N_2749,N_729,N_1283);
nor U2750 (N_2750,N_1,N_661);
nor U2751 (N_2751,N_809,N_1423);
or U2752 (N_2752,N_279,N_1206);
xor U2753 (N_2753,N_1089,N_1036);
nor U2754 (N_2754,N_863,N_937);
or U2755 (N_2755,N_1407,N_297);
nand U2756 (N_2756,N_934,N_477);
or U2757 (N_2757,N_1093,N_82);
nor U2758 (N_2758,N_164,N_1192);
or U2759 (N_2759,N_199,N_466);
xor U2760 (N_2760,N_988,N_898);
and U2761 (N_2761,N_510,N_623);
nand U2762 (N_2762,N_908,N_1062);
nand U2763 (N_2763,N_9,N_128);
nor U2764 (N_2764,N_572,N_694);
nand U2765 (N_2765,N_711,N_147);
xor U2766 (N_2766,N_927,N_652);
nand U2767 (N_2767,N_1183,N_633);
xor U2768 (N_2768,N_1421,N_1206);
or U2769 (N_2769,N_0,N_1366);
nor U2770 (N_2770,N_184,N_879);
and U2771 (N_2771,N_1238,N_365);
nand U2772 (N_2772,N_244,N_201);
nand U2773 (N_2773,N_1091,N_1083);
nor U2774 (N_2774,N_172,N_494);
nand U2775 (N_2775,N_125,N_1496);
or U2776 (N_2776,N_155,N_1238);
nand U2777 (N_2777,N_191,N_1265);
and U2778 (N_2778,N_782,N_1035);
and U2779 (N_2779,N_1490,N_1099);
or U2780 (N_2780,N_234,N_138);
and U2781 (N_2781,N_1251,N_442);
xor U2782 (N_2782,N_949,N_229);
and U2783 (N_2783,N_1298,N_1260);
or U2784 (N_2784,N_1117,N_565);
or U2785 (N_2785,N_729,N_1347);
xnor U2786 (N_2786,N_294,N_1443);
xor U2787 (N_2787,N_774,N_781);
xnor U2788 (N_2788,N_491,N_1229);
and U2789 (N_2789,N_1203,N_868);
and U2790 (N_2790,N_860,N_546);
or U2791 (N_2791,N_364,N_995);
nand U2792 (N_2792,N_1289,N_748);
or U2793 (N_2793,N_109,N_847);
nor U2794 (N_2794,N_1227,N_1129);
and U2795 (N_2795,N_1286,N_1163);
xor U2796 (N_2796,N_1025,N_258);
or U2797 (N_2797,N_996,N_889);
xor U2798 (N_2798,N_1332,N_636);
nand U2799 (N_2799,N_516,N_1213);
and U2800 (N_2800,N_747,N_1206);
or U2801 (N_2801,N_195,N_289);
nand U2802 (N_2802,N_141,N_920);
nand U2803 (N_2803,N_355,N_1039);
nand U2804 (N_2804,N_1397,N_419);
and U2805 (N_2805,N_650,N_836);
xnor U2806 (N_2806,N_676,N_1378);
xnor U2807 (N_2807,N_744,N_833);
xnor U2808 (N_2808,N_871,N_1092);
nor U2809 (N_2809,N_319,N_1315);
and U2810 (N_2810,N_116,N_648);
or U2811 (N_2811,N_942,N_723);
xnor U2812 (N_2812,N_841,N_1368);
and U2813 (N_2813,N_801,N_217);
nor U2814 (N_2814,N_987,N_612);
xor U2815 (N_2815,N_1285,N_303);
nor U2816 (N_2816,N_1206,N_1255);
and U2817 (N_2817,N_856,N_228);
xnor U2818 (N_2818,N_394,N_254);
nor U2819 (N_2819,N_1265,N_840);
xor U2820 (N_2820,N_1444,N_681);
and U2821 (N_2821,N_367,N_29);
nand U2822 (N_2822,N_504,N_5);
nor U2823 (N_2823,N_1203,N_1198);
nor U2824 (N_2824,N_710,N_1077);
nor U2825 (N_2825,N_951,N_1158);
and U2826 (N_2826,N_952,N_143);
xnor U2827 (N_2827,N_777,N_553);
xnor U2828 (N_2828,N_550,N_1410);
nand U2829 (N_2829,N_1026,N_636);
or U2830 (N_2830,N_258,N_131);
or U2831 (N_2831,N_763,N_11);
nor U2832 (N_2832,N_993,N_957);
xor U2833 (N_2833,N_703,N_609);
or U2834 (N_2834,N_373,N_1347);
and U2835 (N_2835,N_336,N_195);
nand U2836 (N_2836,N_876,N_97);
nor U2837 (N_2837,N_934,N_444);
nor U2838 (N_2838,N_1051,N_801);
or U2839 (N_2839,N_719,N_1142);
or U2840 (N_2840,N_191,N_122);
or U2841 (N_2841,N_500,N_819);
nor U2842 (N_2842,N_819,N_1337);
or U2843 (N_2843,N_1063,N_17);
nand U2844 (N_2844,N_238,N_217);
xor U2845 (N_2845,N_748,N_549);
nor U2846 (N_2846,N_1084,N_1328);
or U2847 (N_2847,N_1470,N_266);
or U2848 (N_2848,N_825,N_869);
xor U2849 (N_2849,N_908,N_452);
nor U2850 (N_2850,N_704,N_659);
and U2851 (N_2851,N_485,N_208);
nand U2852 (N_2852,N_593,N_333);
xnor U2853 (N_2853,N_1399,N_1246);
nor U2854 (N_2854,N_145,N_407);
nor U2855 (N_2855,N_125,N_1023);
nand U2856 (N_2856,N_1114,N_52);
nand U2857 (N_2857,N_309,N_768);
and U2858 (N_2858,N_1492,N_993);
xor U2859 (N_2859,N_1061,N_522);
or U2860 (N_2860,N_211,N_1240);
and U2861 (N_2861,N_929,N_1149);
and U2862 (N_2862,N_1343,N_534);
nor U2863 (N_2863,N_357,N_850);
nor U2864 (N_2864,N_89,N_10);
or U2865 (N_2865,N_302,N_805);
xor U2866 (N_2866,N_1412,N_177);
nand U2867 (N_2867,N_630,N_957);
nand U2868 (N_2868,N_583,N_637);
nand U2869 (N_2869,N_1029,N_486);
or U2870 (N_2870,N_548,N_662);
and U2871 (N_2871,N_509,N_900);
or U2872 (N_2872,N_490,N_928);
and U2873 (N_2873,N_153,N_763);
or U2874 (N_2874,N_194,N_602);
or U2875 (N_2875,N_319,N_697);
xor U2876 (N_2876,N_1079,N_836);
xnor U2877 (N_2877,N_416,N_1212);
xor U2878 (N_2878,N_196,N_834);
and U2879 (N_2879,N_437,N_813);
nand U2880 (N_2880,N_1326,N_1339);
xor U2881 (N_2881,N_628,N_364);
nor U2882 (N_2882,N_815,N_38);
and U2883 (N_2883,N_895,N_421);
or U2884 (N_2884,N_516,N_39);
nor U2885 (N_2885,N_261,N_656);
or U2886 (N_2886,N_502,N_1364);
nor U2887 (N_2887,N_811,N_1109);
nor U2888 (N_2888,N_467,N_62);
xor U2889 (N_2889,N_382,N_853);
or U2890 (N_2890,N_922,N_622);
nand U2891 (N_2891,N_120,N_1072);
nor U2892 (N_2892,N_340,N_229);
nor U2893 (N_2893,N_1104,N_1225);
nand U2894 (N_2894,N_777,N_1415);
xor U2895 (N_2895,N_696,N_1352);
and U2896 (N_2896,N_1401,N_403);
or U2897 (N_2897,N_999,N_735);
nand U2898 (N_2898,N_1196,N_958);
nor U2899 (N_2899,N_134,N_674);
nor U2900 (N_2900,N_927,N_135);
and U2901 (N_2901,N_1357,N_1375);
nor U2902 (N_2902,N_693,N_509);
nand U2903 (N_2903,N_1357,N_115);
xnor U2904 (N_2904,N_299,N_1349);
xor U2905 (N_2905,N_933,N_532);
and U2906 (N_2906,N_1355,N_897);
nor U2907 (N_2907,N_1428,N_513);
nor U2908 (N_2908,N_1007,N_450);
or U2909 (N_2909,N_1180,N_392);
and U2910 (N_2910,N_281,N_425);
and U2911 (N_2911,N_725,N_590);
nand U2912 (N_2912,N_203,N_120);
or U2913 (N_2913,N_893,N_896);
and U2914 (N_2914,N_1310,N_1109);
xnor U2915 (N_2915,N_835,N_253);
nand U2916 (N_2916,N_1057,N_365);
nor U2917 (N_2917,N_827,N_520);
nor U2918 (N_2918,N_764,N_493);
and U2919 (N_2919,N_681,N_814);
or U2920 (N_2920,N_1308,N_839);
or U2921 (N_2921,N_892,N_1461);
and U2922 (N_2922,N_276,N_174);
xnor U2923 (N_2923,N_718,N_1298);
xnor U2924 (N_2924,N_1118,N_1289);
nor U2925 (N_2925,N_684,N_767);
xnor U2926 (N_2926,N_1265,N_645);
and U2927 (N_2927,N_700,N_593);
nor U2928 (N_2928,N_146,N_925);
and U2929 (N_2929,N_140,N_457);
nor U2930 (N_2930,N_83,N_1110);
nor U2931 (N_2931,N_61,N_571);
or U2932 (N_2932,N_1267,N_357);
and U2933 (N_2933,N_888,N_97);
nor U2934 (N_2934,N_915,N_1186);
xnor U2935 (N_2935,N_1155,N_498);
xor U2936 (N_2936,N_615,N_782);
nand U2937 (N_2937,N_114,N_803);
xor U2938 (N_2938,N_1188,N_548);
and U2939 (N_2939,N_474,N_1403);
xnor U2940 (N_2940,N_660,N_1259);
or U2941 (N_2941,N_324,N_1387);
or U2942 (N_2942,N_201,N_303);
and U2943 (N_2943,N_49,N_882);
nand U2944 (N_2944,N_1044,N_183);
or U2945 (N_2945,N_327,N_470);
nand U2946 (N_2946,N_202,N_1382);
and U2947 (N_2947,N_913,N_1118);
nor U2948 (N_2948,N_1149,N_961);
nor U2949 (N_2949,N_1259,N_668);
xnor U2950 (N_2950,N_325,N_668);
or U2951 (N_2951,N_765,N_1434);
nand U2952 (N_2952,N_1190,N_876);
and U2953 (N_2953,N_799,N_39);
and U2954 (N_2954,N_462,N_1446);
nand U2955 (N_2955,N_547,N_1274);
xor U2956 (N_2956,N_160,N_266);
or U2957 (N_2957,N_1485,N_386);
and U2958 (N_2958,N_657,N_938);
nor U2959 (N_2959,N_1321,N_1312);
and U2960 (N_2960,N_367,N_655);
xor U2961 (N_2961,N_687,N_36);
nand U2962 (N_2962,N_729,N_381);
nand U2963 (N_2963,N_1364,N_291);
xnor U2964 (N_2964,N_945,N_348);
xor U2965 (N_2965,N_705,N_1170);
nand U2966 (N_2966,N_337,N_818);
nor U2967 (N_2967,N_172,N_1428);
nand U2968 (N_2968,N_696,N_115);
nor U2969 (N_2969,N_1221,N_1031);
nand U2970 (N_2970,N_545,N_1359);
or U2971 (N_2971,N_282,N_190);
xnor U2972 (N_2972,N_803,N_562);
nor U2973 (N_2973,N_960,N_71);
xnor U2974 (N_2974,N_1442,N_1073);
nand U2975 (N_2975,N_444,N_700);
nor U2976 (N_2976,N_249,N_109);
xor U2977 (N_2977,N_232,N_119);
and U2978 (N_2978,N_1442,N_275);
or U2979 (N_2979,N_1311,N_1122);
xor U2980 (N_2980,N_286,N_924);
or U2981 (N_2981,N_909,N_1336);
nor U2982 (N_2982,N_133,N_809);
nor U2983 (N_2983,N_299,N_441);
nor U2984 (N_2984,N_900,N_139);
or U2985 (N_2985,N_982,N_932);
nor U2986 (N_2986,N_872,N_264);
nand U2987 (N_2987,N_1177,N_1470);
or U2988 (N_2988,N_1134,N_370);
nand U2989 (N_2989,N_1106,N_1299);
nand U2990 (N_2990,N_1172,N_943);
xnor U2991 (N_2991,N_1135,N_986);
nor U2992 (N_2992,N_1138,N_1116);
and U2993 (N_2993,N_23,N_666);
or U2994 (N_2994,N_171,N_531);
nand U2995 (N_2995,N_1061,N_391);
or U2996 (N_2996,N_1394,N_466);
nand U2997 (N_2997,N_1004,N_1488);
nand U2998 (N_2998,N_972,N_1488);
and U2999 (N_2999,N_157,N_693);
nand U3000 (N_3000,N_2188,N_2328);
nor U3001 (N_3001,N_1905,N_1895);
xor U3002 (N_3002,N_2797,N_2110);
nor U3003 (N_3003,N_2184,N_1919);
xor U3004 (N_3004,N_2627,N_2150);
nor U3005 (N_3005,N_2850,N_2487);
nor U3006 (N_3006,N_1553,N_2500);
and U3007 (N_3007,N_2421,N_2599);
and U3008 (N_3008,N_2633,N_2573);
xor U3009 (N_3009,N_2350,N_2557);
xor U3010 (N_3010,N_2751,N_2798);
xnor U3011 (N_3011,N_1943,N_2276);
xor U3012 (N_3012,N_2058,N_1954);
nor U3013 (N_3013,N_2274,N_2118);
and U3014 (N_3014,N_2712,N_2509);
and U3015 (N_3015,N_2539,N_2919);
nor U3016 (N_3016,N_2192,N_2843);
xnor U3017 (N_3017,N_2203,N_2194);
nand U3018 (N_3018,N_2742,N_1639);
xnor U3019 (N_3019,N_2607,N_2541);
nand U3020 (N_3020,N_1947,N_2172);
and U3021 (N_3021,N_2102,N_2068);
nor U3022 (N_3022,N_1876,N_2868);
or U3023 (N_3023,N_2445,N_2891);
or U3024 (N_3024,N_2206,N_1546);
nand U3025 (N_3025,N_2837,N_2855);
and U3026 (N_3026,N_1679,N_2489);
xor U3027 (N_3027,N_1501,N_1863);
nor U3028 (N_3028,N_2448,N_2444);
xor U3029 (N_3029,N_2610,N_1861);
xnor U3030 (N_3030,N_1759,N_2830);
nand U3031 (N_3031,N_1878,N_1978);
nand U3032 (N_3032,N_1793,N_2105);
nand U3033 (N_3033,N_2289,N_2481);
xor U3034 (N_3034,N_2637,N_1684);
and U3035 (N_3035,N_1825,N_2734);
nor U3036 (N_3036,N_2628,N_2364);
nor U3037 (N_3037,N_2251,N_2626);
nor U3038 (N_3038,N_2567,N_2312);
nor U3039 (N_3039,N_2848,N_1686);
nand U3040 (N_3040,N_2580,N_2208);
or U3041 (N_3041,N_2136,N_2993);
and U3042 (N_3042,N_2578,N_2072);
and U3043 (N_3043,N_1627,N_2323);
nand U3044 (N_3044,N_2232,N_2715);
and U3045 (N_3045,N_2317,N_1646);
or U3046 (N_3046,N_1768,N_2186);
nand U3047 (N_3047,N_1617,N_2763);
xor U3048 (N_3048,N_2882,N_2934);
and U3049 (N_3049,N_2017,N_2166);
and U3050 (N_3050,N_2080,N_2288);
xor U3051 (N_3051,N_1711,N_1915);
nand U3052 (N_3052,N_1827,N_2488);
nand U3053 (N_3053,N_1666,N_2769);
nand U3054 (N_3054,N_1846,N_2319);
and U3055 (N_3055,N_2320,N_2761);
or U3056 (N_3056,N_2051,N_2417);
nand U3057 (N_3057,N_2157,N_2684);
nand U3058 (N_3058,N_1875,N_2482);
nor U3059 (N_3059,N_2899,N_2402);
nor U3060 (N_3060,N_2461,N_2928);
or U3061 (N_3061,N_2505,N_1537);
or U3062 (N_3062,N_1731,N_2070);
nand U3063 (N_3063,N_2400,N_1688);
xnor U3064 (N_3064,N_2493,N_2059);
nor U3065 (N_3065,N_1693,N_1662);
nand U3066 (N_3066,N_1937,N_2237);
xnor U3067 (N_3067,N_1559,N_2268);
nand U3068 (N_3068,N_2191,N_2923);
nand U3069 (N_3069,N_1908,N_2709);
or U3070 (N_3070,N_1599,N_2249);
and U3071 (N_3071,N_2021,N_2254);
xnor U3072 (N_3072,N_2436,N_1916);
and U3073 (N_3073,N_1552,N_1841);
nor U3074 (N_3074,N_1555,N_2248);
nand U3075 (N_3075,N_1781,N_1900);
nor U3076 (N_3076,N_2643,N_1758);
nand U3077 (N_3077,N_2281,N_2615);
nor U3078 (N_3078,N_2373,N_2532);
xor U3079 (N_3079,N_2201,N_2877);
nand U3080 (N_3080,N_1609,N_2006);
nor U3081 (N_3081,N_2153,N_2949);
xnor U3082 (N_3082,N_2937,N_1565);
nor U3083 (N_3083,N_2778,N_2951);
xor U3084 (N_3084,N_1784,N_1745);
and U3085 (N_3085,N_1914,N_2936);
nand U3086 (N_3086,N_1574,N_2592);
nand U3087 (N_3087,N_2047,N_2329);
or U3088 (N_3088,N_1920,N_1749);
nand U3089 (N_3089,N_2696,N_1761);
and U3090 (N_3090,N_1587,N_2468);
nand U3091 (N_3091,N_2943,N_2990);
and U3092 (N_3092,N_2386,N_1635);
nor U3093 (N_3093,N_2008,N_1752);
xor U3094 (N_3094,N_2754,N_2512);
and U3095 (N_3095,N_1695,N_2681);
nand U3096 (N_3096,N_2087,N_2388);
or U3097 (N_3097,N_2605,N_2582);
or U3098 (N_3098,N_2563,N_1826);
and U3099 (N_3099,N_2521,N_1830);
nand U3100 (N_3100,N_2524,N_1692);
or U3101 (N_3101,N_2959,N_1787);
and U3102 (N_3102,N_2128,N_2978);
nor U3103 (N_3103,N_2939,N_2406);
nor U3104 (N_3104,N_1535,N_2679);
or U3105 (N_3105,N_2533,N_1691);
nor U3106 (N_3106,N_2915,N_1869);
nand U3107 (N_3107,N_2957,N_2473);
nor U3108 (N_3108,N_1655,N_2759);
and U3109 (N_3109,N_2829,N_2185);
or U3110 (N_3110,N_2429,N_2976);
xor U3111 (N_3111,N_1816,N_1744);
nor U3112 (N_3112,N_2921,N_2499);
nor U3113 (N_3113,N_1653,N_1969);
nor U3114 (N_3114,N_2093,N_2299);
nor U3115 (N_3115,N_1562,N_2897);
and U3116 (N_3116,N_2731,N_2062);
nand U3117 (N_3117,N_2716,N_2282);
xnor U3118 (N_3118,N_1677,N_1796);
nand U3119 (N_3119,N_2711,N_2974);
nand U3120 (N_3120,N_1697,N_1585);
nand U3121 (N_3121,N_2073,N_2480);
nor U3122 (N_3122,N_2581,N_2832);
nor U3123 (N_3123,N_2924,N_1897);
xor U3124 (N_3124,N_1614,N_2649);
or U3125 (N_3125,N_1853,N_2371);
or U3126 (N_3126,N_2361,N_2440);
or U3127 (N_3127,N_1851,N_1786);
nor U3128 (N_3128,N_1938,N_2700);
and U3129 (N_3129,N_2146,N_1959);
and U3130 (N_3130,N_2630,N_2587);
or U3131 (N_3131,N_2556,N_2728);
nand U3132 (N_3132,N_1933,N_1556);
nand U3133 (N_3133,N_1766,N_2652);
xnor U3134 (N_3134,N_2180,N_2531);
and U3135 (N_3135,N_2239,N_1723);
xor U3136 (N_3136,N_1712,N_2635);
nor U3137 (N_3137,N_1970,N_1683);
xor U3138 (N_3138,N_1868,N_1615);
nor U3139 (N_3139,N_2857,N_1531);
xnor U3140 (N_3140,N_2434,N_2562);
or U3141 (N_3141,N_2423,N_1660);
or U3142 (N_3142,N_2870,N_2253);
and U3143 (N_3143,N_2964,N_2694);
nand U3144 (N_3144,N_2106,N_2033);
nor U3145 (N_3145,N_1940,N_1981);
nand U3146 (N_3146,N_2397,N_1831);
nand U3147 (N_3147,N_1833,N_2977);
nor U3148 (N_3148,N_2376,N_1917);
or U3149 (N_3149,N_1586,N_2647);
or U3150 (N_3150,N_1772,N_2227);
and U3151 (N_3151,N_2243,N_2552);
nor U3152 (N_3152,N_2663,N_2796);
nor U3153 (N_3153,N_2139,N_2379);
nor U3154 (N_3154,N_2453,N_1631);
or U3155 (N_3155,N_2382,N_2534);
nand U3156 (N_3156,N_1945,N_1698);
and U3157 (N_3157,N_2902,N_2776);
xor U3158 (N_3158,N_2212,N_1626);
nor U3159 (N_3159,N_2967,N_2735);
and U3160 (N_3160,N_1799,N_2846);
xor U3161 (N_3161,N_2727,N_2875);
and U3162 (N_3162,N_2507,N_2931);
or U3163 (N_3163,N_2665,N_2876);
nor U3164 (N_3164,N_2634,N_2290);
or U3165 (N_3165,N_1946,N_2775);
xor U3166 (N_3166,N_2835,N_1887);
nor U3167 (N_3167,N_2001,N_2656);
or U3168 (N_3168,N_2218,N_2749);
nand U3169 (N_3169,N_2351,N_2654);
nand U3170 (N_3170,N_1742,N_2960);
nor U3171 (N_3171,N_2304,N_2571);
or U3172 (N_3172,N_1906,N_2321);
and U3173 (N_3173,N_2409,N_1505);
or U3174 (N_3174,N_2041,N_2045);
and U3175 (N_3175,N_2853,N_2660);
or U3176 (N_3176,N_2365,N_1973);
and U3177 (N_3177,N_2026,N_2081);
or U3178 (N_3178,N_2585,N_1873);
xor U3179 (N_3179,N_1608,N_2459);
or U3180 (N_3180,N_2173,N_2800);
nor U3181 (N_3181,N_1767,N_2447);
nor U3182 (N_3182,N_1707,N_2893);
or U3183 (N_3183,N_1950,N_1942);
xnor U3184 (N_3184,N_1842,N_1741);
xnor U3185 (N_3185,N_1771,N_2553);
xor U3186 (N_3186,N_2456,N_1699);
xnor U3187 (N_3187,N_2549,N_2820);
nor U3188 (N_3188,N_1650,N_2815);
nor U3189 (N_3189,N_2278,N_2662);
xnor U3190 (N_3190,N_1910,N_1717);
nand U3191 (N_3191,N_1704,N_2140);
nand U3192 (N_3192,N_2971,N_2529);
nand U3193 (N_3193,N_2123,N_2730);
nand U3194 (N_3194,N_2917,N_1618);
xnor U3195 (N_3195,N_2010,N_2392);
nand U3196 (N_3196,N_1719,N_2209);
xor U3197 (N_3197,N_1604,N_2852);
and U3198 (N_3198,N_1665,N_2104);
or U3199 (N_3199,N_2955,N_2819);
nand U3200 (N_3200,N_2393,N_2012);
nand U3201 (N_3201,N_2621,N_1814);
or U3202 (N_3202,N_2519,N_2762);
nand U3203 (N_3203,N_1746,N_2871);
or U3204 (N_3204,N_2043,N_2219);
and U3205 (N_3205,N_2141,N_1957);
nor U3206 (N_3206,N_1990,N_2407);
nand U3207 (N_3207,N_1748,N_2691);
or U3208 (N_3208,N_1648,N_2674);
xor U3209 (N_3209,N_2362,N_1934);
nand U3210 (N_3210,N_2925,N_1901);
xor U3211 (N_3211,N_2183,N_2619);
xnor U3212 (N_3212,N_1571,N_2739);
xnor U3213 (N_3213,N_1652,N_1611);
nand U3214 (N_3214,N_2903,N_2994);
nor U3215 (N_3215,N_2228,N_1857);
nor U3216 (N_3216,N_2119,N_2866);
nor U3217 (N_3217,N_1521,N_1867);
and U3218 (N_3218,N_2451,N_2551);
nand U3219 (N_3219,N_2314,N_2189);
and U3220 (N_3220,N_1638,N_2167);
nand U3221 (N_3221,N_1709,N_2113);
nor U3222 (N_3222,N_1924,N_2294);
xnor U3223 (N_3223,N_2432,N_1927);
nor U3224 (N_3224,N_2612,N_2344);
and U3225 (N_3225,N_2325,N_2296);
xnor U3226 (N_3226,N_1583,N_1725);
nor U3227 (N_3227,N_2358,N_2911);
nand U3228 (N_3228,N_2682,N_2544);
xor U3229 (N_3229,N_2063,N_2708);
and U3230 (N_3230,N_2992,N_1821);
nor U3231 (N_3231,N_2217,N_2530);
nand U3232 (N_3232,N_2300,N_2152);
nor U3233 (N_3233,N_2805,N_2211);
or U3234 (N_3234,N_1542,N_1909);
or U3235 (N_3235,N_2414,N_2190);
xnor U3236 (N_3236,N_2498,N_2442);
and U3237 (N_3237,N_2596,N_2437);
nand U3238 (N_3238,N_2623,N_2116);
xnor U3239 (N_3239,N_2604,N_2458);
nand U3240 (N_3240,N_1886,N_2287);
and U3241 (N_3241,N_2095,N_2618);
nor U3242 (N_3242,N_1925,N_2575);
xnor U3243 (N_3243,N_2168,N_2109);
and U3244 (N_3244,N_2540,N_2079);
and U3245 (N_3245,N_2688,N_1975);
nor U3246 (N_3246,N_1832,N_1534);
or U3247 (N_3247,N_1602,N_2035);
or U3248 (N_3248,N_2309,N_1680);
nor U3249 (N_3249,N_2395,N_2327);
xnor U3250 (N_3250,N_2983,N_2920);
nand U3251 (N_3251,N_2584,N_2678);
xor U3252 (N_3252,N_1507,N_2845);
nor U3253 (N_3253,N_1997,N_2375);
nor U3254 (N_3254,N_2881,N_2205);
and U3255 (N_3255,N_1852,N_1517);
nand U3256 (N_3256,N_2690,N_2069);
nor U3257 (N_3257,N_2947,N_2683);
and U3258 (N_3258,N_2018,N_2378);
nor U3259 (N_3259,N_1685,N_1949);
nor U3260 (N_3260,N_2611,N_2291);
and U3261 (N_3261,N_2600,N_1977);
nand U3262 (N_3262,N_2430,N_2965);
nand U3263 (N_3263,N_1613,N_2023);
or U3264 (N_3264,N_2394,N_1641);
nand U3265 (N_3265,N_2736,N_2779);
xnor U3266 (N_3266,N_1728,N_2616);
xor U3267 (N_3267,N_2638,N_2302);
xnor U3268 (N_3268,N_2435,N_2914);
nor U3269 (N_3269,N_1636,N_2096);
and U3270 (N_3270,N_2060,N_2197);
or U3271 (N_3271,N_2439,N_2367);
xor U3272 (N_3272,N_2280,N_2103);
nor U3273 (N_3273,N_1729,N_1865);
xor U3274 (N_3274,N_1808,N_2940);
xor U3275 (N_3275,N_1822,N_1502);
nor U3276 (N_3276,N_1656,N_2174);
or U3277 (N_3277,N_2339,N_1755);
or U3278 (N_3278,N_1563,N_1524);
nor U3279 (N_3279,N_1775,N_2066);
nand U3280 (N_3280,N_2804,N_1823);
or U3281 (N_3281,N_2120,N_2617);
nor U3282 (N_3282,N_1912,N_1770);
and U3283 (N_3283,N_1989,N_1893);
or U3284 (N_3284,N_2163,N_1840);
xnor U3285 (N_3285,N_2090,N_2518);
xnor U3286 (N_3286,N_1612,N_1575);
nor U3287 (N_3287,N_2029,N_2667);
nand U3288 (N_3288,N_2216,N_2037);
or U3289 (N_3289,N_1543,N_1667);
nor U3290 (N_3290,N_2181,N_2816);
nor U3291 (N_3291,N_1913,N_1762);
or U3292 (N_3292,N_1682,N_1750);
or U3293 (N_3293,N_1670,N_1918);
xnor U3294 (N_3294,N_2595,N_2858);
nand U3295 (N_3295,N_2740,N_1972);
or U3296 (N_3296,N_1804,N_2067);
nor U3297 (N_3297,N_1991,N_2420);
or U3298 (N_3298,N_2454,N_2865);
xor U3299 (N_3299,N_2396,N_2101);
xnor U3300 (N_3300,N_2622,N_2537);
nand U3301 (N_3301,N_1965,N_2520);
xnor U3302 (N_3302,N_2279,N_2810);
nor U3303 (N_3303,N_1928,N_1544);
nor U3304 (N_3304,N_1605,N_1738);
and U3305 (N_3305,N_2151,N_2833);
nand U3306 (N_3306,N_1883,N_2494);
and U3307 (N_3307,N_2391,N_2655);
nor U3308 (N_3308,N_2542,N_1603);
and U3309 (N_3309,N_2257,N_2705);
nor U3310 (N_3310,N_2071,N_2699);
xnor U3311 (N_3311,N_2464,N_2303);
and U3312 (N_3312,N_2515,N_1678);
or U3313 (N_3313,N_1760,N_2873);
nor U3314 (N_3314,N_1889,N_2545);
or U3315 (N_3315,N_2771,N_2024);
nor U3316 (N_3316,N_2286,N_2784);
xor U3317 (N_3317,N_1663,N_2252);
or U3318 (N_3318,N_2370,N_2020);
nand U3319 (N_3319,N_1545,N_2044);
and U3320 (N_3320,N_1668,N_2236);
xor U3321 (N_3321,N_1926,N_1547);
xor U3322 (N_3322,N_2813,N_2231);
xor U3323 (N_3323,N_1533,N_2221);
nand U3324 (N_3324,N_2295,N_2526);
xnor U3325 (N_3325,N_2441,N_1658);
or U3326 (N_3326,N_2854,N_2559);
nand U3327 (N_3327,N_1500,N_1952);
xor U3328 (N_3328,N_2117,N_1885);
and U3329 (N_3329,N_2648,N_1664);
or U3330 (N_3330,N_2111,N_2745);
and U3331 (N_3331,N_1736,N_1988);
xnor U3332 (N_3332,N_1982,N_2692);
nor U3333 (N_3333,N_1519,N_2210);
xnor U3334 (N_3334,N_2790,N_2415);
and U3335 (N_3335,N_1783,N_2410);
nand U3336 (N_3336,N_2952,N_2387);
nor U3337 (N_3337,N_1835,N_2591);
or U3338 (N_3338,N_1509,N_2015);
nor U3339 (N_3339,N_2326,N_1932);
nor U3340 (N_3340,N_1870,N_1862);
xor U3341 (N_3341,N_2603,N_2646);
nand U3342 (N_3342,N_2996,N_2277);
nor U3343 (N_3343,N_2298,N_2431);
xnor U3344 (N_3344,N_2213,N_1705);
xor U3345 (N_3345,N_2703,N_2478);
and U3346 (N_3346,N_2950,N_1856);
xor U3347 (N_3347,N_2697,N_2503);
nand U3348 (N_3348,N_2199,N_2476);
and U3349 (N_3349,N_1582,N_2527);
nor U3350 (N_3350,N_1721,N_2273);
nand U3351 (N_3351,N_2831,N_2910);
or U3352 (N_3352,N_2084,N_2864);
nor U3353 (N_3353,N_2786,N_2022);
or U3354 (N_3354,N_2668,N_2054);
and U3355 (N_3355,N_2650,N_2625);
and U3356 (N_3356,N_2064,N_2849);
and U3357 (N_3357,N_1961,N_2721);
nor U3358 (N_3358,N_2052,N_2789);
nand U3359 (N_3359,N_2474,N_1992);
nor U3360 (N_3360,N_2042,N_2972);
nand U3361 (N_3361,N_2985,N_2477);
and U3362 (N_3362,N_2177,N_1829);
nand U3363 (N_3363,N_2357,N_1795);
nand U3364 (N_3364,N_2270,N_2817);
nor U3365 (N_3365,N_2785,N_2133);
and U3366 (N_3366,N_2782,N_1813);
nor U3367 (N_3367,N_2196,N_2861);
and U3368 (N_3368,N_2672,N_2057);
xor U3369 (N_3369,N_1708,N_2982);
nor U3370 (N_3370,N_2859,N_2121);
xnor U3371 (N_3371,N_2510,N_2025);
xnor U3372 (N_3372,N_1568,N_2576);
and U3373 (N_3373,N_2872,N_2082);
and U3374 (N_3374,N_2412,N_1776);
and U3375 (N_3375,N_2718,N_2341);
nand U3376 (N_3376,N_2988,N_1706);
nand U3377 (N_3377,N_1740,N_2000);
nor U3378 (N_3378,N_2543,N_2536);
xnor U3379 (N_3379,N_2337,N_1577);
or U3380 (N_3380,N_1516,N_2258);
xnor U3381 (N_3381,N_2175,N_1642);
nor U3382 (N_3382,N_1894,N_2085);
nand U3383 (N_3383,N_2165,N_2200);
and U3384 (N_3384,N_2956,N_2124);
nand U3385 (N_3385,N_2061,N_1881);
nand U3386 (N_3386,N_1659,N_1751);
and U3387 (N_3387,N_1780,N_2313);
xor U3388 (N_3388,N_1737,N_2677);
nor U3389 (N_3389,N_1807,N_2701);
or U3390 (N_3390,N_2564,N_1790);
or U3391 (N_3391,N_1979,N_2094);
xnor U3392 (N_3392,N_1694,N_2879);
nand U3393 (N_3393,N_2132,N_1743);
xor U3394 (N_3394,N_2032,N_2342);
or U3395 (N_3395,N_2720,N_2787);
xnor U3396 (N_3396,N_1640,N_2267);
and U3397 (N_3397,N_2598,N_2687);
or U3398 (N_3398,N_2841,N_2307);
xor U3399 (N_3399,N_1960,N_2565);
nor U3400 (N_3400,N_2706,N_1968);
nand U3401 (N_3401,N_1994,N_2443);
or U3402 (N_3402,N_2310,N_2486);
or U3403 (N_3403,N_1936,N_2242);
nor U3404 (N_3404,N_2752,N_2896);
or U3405 (N_3405,N_2372,N_2568);
nor U3406 (N_3406,N_1904,N_2013);
nand U3407 (N_3407,N_2144,N_2572);
nand U3408 (N_3408,N_2159,N_2651);
or U3409 (N_3409,N_2457,N_2083);
or U3410 (N_3410,N_1733,N_2844);
and U3411 (N_3411,N_2698,N_2856);
or U3412 (N_3412,N_2097,N_2099);
and U3413 (N_3413,N_2331,N_2629);
or U3414 (N_3414,N_2970,N_2129);
or U3415 (N_3415,N_2946,N_2918);
xnor U3416 (N_3416,N_2220,N_1632);
xnor U3417 (N_3417,N_2352,N_2502);
and U3418 (N_3418,N_2422,N_1593);
nand U3419 (N_3419,N_2997,N_2424);
or U3420 (N_3420,N_2160,N_1566);
or U3421 (N_3421,N_2263,N_1657);
xnor U3422 (N_3422,N_2222,N_2377);
nand U3423 (N_3423,N_2538,N_2765);
xnor U3424 (N_3424,N_1690,N_2803);
and U3425 (N_3425,N_2380,N_2466);
xor U3426 (N_3426,N_2030,N_2636);
or U3427 (N_3427,N_1523,N_2385);
and U3428 (N_3428,N_1578,N_2156);
and U3429 (N_3429,N_2425,N_1896);
nand U3430 (N_3430,N_1864,N_2348);
nor U3431 (N_3431,N_1576,N_1844);
nand U3432 (N_3432,N_2704,N_2193);
nor U3433 (N_3433,N_2889,N_2075);
xnor U3434 (N_3434,N_2065,N_2034);
or U3435 (N_3435,N_1527,N_2399);
nand U3436 (N_3436,N_1675,N_1696);
nor U3437 (N_3437,N_2433,N_1782);
xor U3438 (N_3438,N_1956,N_2469);
nand U3439 (N_3439,N_1794,N_1701);
nand U3440 (N_3440,N_2586,N_2593);
and U3441 (N_3441,N_1600,N_2086);
xnor U3442 (N_3442,N_2485,N_1525);
xnor U3443 (N_3443,N_2301,N_2702);
nor U3444 (N_3444,N_1558,N_1763);
xor U3445 (N_3445,N_2491,N_2011);
nand U3446 (N_3446,N_2525,N_1929);
nor U3447 (N_3447,N_2574,N_2418);
or U3448 (N_3448,N_2463,N_2261);
and U3449 (N_3449,N_1518,N_1777);
and U3450 (N_3450,N_1859,N_2330);
and U3451 (N_3451,N_2948,N_2383);
or U3452 (N_3452,N_1998,N_2826);
nand U3453 (N_3453,N_1922,N_2641);
nor U3454 (N_3454,N_2675,N_2389);
xor U3455 (N_3455,N_2980,N_1958);
xnor U3456 (N_3456,N_2710,N_1597);
nand U3457 (N_3457,N_2570,N_1623);
xor U3458 (N_3458,N_1687,N_2031);
xnor U3459 (N_3459,N_1674,N_2398);
and U3460 (N_3460,N_2522,N_2901);
and U3461 (N_3461,N_1930,N_2359);
and U3462 (N_3462,N_2148,N_2941);
and U3463 (N_3463,N_1769,N_1986);
and U3464 (N_3464,N_1720,N_2100);
and U3465 (N_3465,N_2229,N_1724);
or U3466 (N_3466,N_2888,N_1515);
nand U3467 (N_3467,N_2091,N_1672);
nor U3468 (N_3468,N_1966,N_2164);
and U3469 (N_3469,N_2913,N_1860);
and U3470 (N_3470,N_1710,N_2986);
and U3471 (N_3471,N_2569,N_1681);
xor U3472 (N_3472,N_2014,N_2756);
nor U3473 (N_3473,N_1557,N_2860);
and U3474 (N_3474,N_2887,N_2723);
and U3475 (N_3475,N_2028,N_2046);
nor U3476 (N_3476,N_2601,N_1530);
nand U3477 (N_3477,N_2195,N_2460);
nand U3478 (N_3478,N_1753,N_2926);
nor U3479 (N_3479,N_2851,N_1734);
nand U3480 (N_3480,N_2606,N_2039);
nor U3481 (N_3481,N_2381,N_2411);
nor U3482 (N_3482,N_2155,N_1999);
or U3483 (N_3483,N_1980,N_2847);
and U3484 (N_3484,N_2269,N_1628);
xor U3485 (N_3485,N_2470,N_2973);
or U3486 (N_3486,N_2271,N_1564);
nor U3487 (N_3487,N_1561,N_2892);
and U3488 (N_3488,N_2811,N_1654);
nor U3489 (N_3489,N_1941,N_2802);
nand U3490 (N_3490,N_2732,N_2981);
nand U3491 (N_3491,N_2839,N_2142);
xnor U3492 (N_3492,N_1837,N_2126);
nand U3493 (N_3493,N_1824,N_2602);
and U3494 (N_3494,N_2535,N_2016);
and U3495 (N_3495,N_1884,N_2496);
or U3496 (N_3496,N_2260,N_2501);
xnor U3497 (N_3497,N_2332,N_2883);
and U3498 (N_3498,N_2202,N_2311);
and U3499 (N_3499,N_2547,N_1726);
and U3500 (N_3500,N_2516,N_1789);
nand U3501 (N_3501,N_2179,N_1645);
nand U3502 (N_3502,N_2235,N_2770);
and U3503 (N_3503,N_2416,N_1948);
or U3504 (N_3504,N_2597,N_1702);
nand U3505 (N_3505,N_1538,N_2945);
nor U3506 (N_3506,N_1774,N_2089);
nor U3507 (N_3507,N_2283,N_2589);
or U3508 (N_3508,N_1730,N_2842);
nor U3509 (N_3509,N_2895,N_2036);
nor U3510 (N_3510,N_1532,N_2475);
xor U3511 (N_3511,N_1797,N_2360);
xnor U3512 (N_3512,N_1669,N_2885);
xnor U3513 (N_3513,N_2640,N_1792);
xnor U3514 (N_3514,N_1625,N_2809);
or U3515 (N_3515,N_2369,N_2419);
and U3516 (N_3516,N_1882,N_2719);
and U3517 (N_3517,N_2078,N_1838);
and U3518 (N_3518,N_2513,N_2528);
nor U3519 (N_3519,N_2401,N_2426);
xor U3520 (N_3520,N_2878,N_2292);
and U3521 (N_3521,N_2867,N_1588);
nand U3522 (N_3522,N_2747,N_1620);
and U3523 (N_3523,N_2497,N_2561);
nand U3524 (N_3524,N_1847,N_2916);
nor U3525 (N_3525,N_2403,N_2255);
xnor U3526 (N_3526,N_2384,N_1570);
or U3527 (N_3527,N_1637,N_2158);
xnor U3528 (N_3528,N_2558,N_1732);
nand U3529 (N_3529,N_2349,N_2223);
or U3530 (N_3530,N_2483,N_2135);
and U3531 (N_3531,N_1963,N_1812);
or U3532 (N_3532,N_2822,N_2741);
xor U3533 (N_3533,N_1967,N_1508);
or U3534 (N_3534,N_1788,N_2056);
xor U3535 (N_3535,N_1747,N_2048);
xor U3536 (N_3536,N_2324,N_2256);
nor U3537 (N_3537,N_2588,N_2169);
or U3538 (N_3538,N_2812,N_2363);
xor U3539 (N_3539,N_2644,N_2673);
xor U3540 (N_3540,N_2695,N_2170);
nor U3541 (N_3541,N_2176,N_2661);
nor U3542 (N_3542,N_2471,N_1778);
nand U3543 (N_3543,N_2958,N_1673);
nor U3544 (N_3544,N_2149,N_2134);
nor U3545 (N_3545,N_1880,N_2262);
or U3546 (N_3546,N_2162,N_2963);
nor U3547 (N_3547,N_1935,N_2178);
nor U3548 (N_3548,N_2954,N_2098);
nor U3549 (N_3549,N_1809,N_1629);
nand U3550 (N_3550,N_1902,N_2297);
and U3551 (N_3551,N_1848,N_1722);
and U3552 (N_3552,N_1843,N_2750);
or U3553 (N_3553,N_2354,N_2777);
nand U3554 (N_3554,N_1594,N_2233);
xnor U3555 (N_3555,N_2807,N_2114);
xnor U3556 (N_3556,N_2620,N_2479);
nor U3557 (N_3557,N_1818,N_1836);
or U3558 (N_3558,N_1549,N_2658);
nor U3559 (N_3559,N_2131,N_2244);
nor U3560 (N_3560,N_1964,N_1536);
and U3561 (N_3561,N_2147,N_1596);
or U3562 (N_3562,N_1589,N_2161);
xnor U3563 (N_3563,N_2115,N_2138);
xor U3564 (N_3564,N_2438,N_2944);
nor U3565 (N_3565,N_1815,N_1805);
and U3566 (N_3566,N_1616,N_2998);
and U3567 (N_3567,N_2215,N_1871);
xnor U3568 (N_3568,N_2345,N_2259);
nor U3569 (N_3569,N_1700,N_2907);
nand U3570 (N_3570,N_2927,N_1572);
and U3571 (N_3571,N_1845,N_2984);
or U3572 (N_3572,N_1944,N_2725);
nand U3573 (N_3573,N_1540,N_2579);
nand U3574 (N_3574,N_1866,N_2315);
and U3575 (N_3575,N_2548,N_2005);
xor U3576 (N_3576,N_2108,N_2880);
or U3577 (N_3577,N_2107,N_2583);
nor U3578 (N_3578,N_2305,N_2226);
and U3579 (N_3579,N_2343,N_2693);
and U3580 (N_3580,N_1630,N_2886);
xor U3581 (N_3581,N_2717,N_2794);
xnor U3582 (N_3582,N_1962,N_1907);
or U3583 (N_3583,N_2686,N_2508);
nand U3584 (N_3584,N_2743,N_2366);
or U3585 (N_3585,N_2791,N_2241);
or U3586 (N_3586,N_1779,N_2356);
or U3587 (N_3587,N_2092,N_2657);
or U3588 (N_3588,N_2904,N_2799);
and U3589 (N_3589,N_1995,N_1526);
and U3590 (N_3590,N_2449,N_1606);
nand U3591 (N_3591,N_1985,N_2758);
xor U3592 (N_3592,N_2130,N_2293);
and U3593 (N_3593,N_1735,N_1898);
and U3594 (N_3594,N_2230,N_2659);
and U3595 (N_3595,N_2427,N_1579);
xnor U3596 (N_3596,N_2322,N_2038);
and U3597 (N_3597,N_1839,N_2609);
nor U3598 (N_3598,N_2207,N_1791);
xor U3599 (N_3599,N_1541,N_2922);
and U3600 (N_3600,N_1633,N_2989);
or U3601 (N_3601,N_1996,N_1671);
and U3602 (N_3602,N_1644,N_2053);
nand U3603 (N_3603,N_2368,N_2355);
nand U3604 (N_3604,N_1955,N_1624);
nand U3605 (N_3605,N_2019,N_2744);
nor U3606 (N_3606,N_2909,N_2225);
and U3607 (N_3607,N_2767,N_1560);
nand U3608 (N_3608,N_1858,N_2204);
or U3609 (N_3609,N_2143,N_2613);
or U3610 (N_3610,N_2737,N_1892);
or U3611 (N_3611,N_1512,N_1718);
nor U3612 (N_3612,N_1573,N_2550);
and U3613 (N_3613,N_2724,N_2793);
nand U3614 (N_3614,N_2265,N_2995);
nor U3615 (N_3615,N_2874,N_2506);
and U3616 (N_3616,N_2768,N_2465);
nor U3617 (N_3617,N_2374,N_2689);
or U3618 (N_3618,N_2801,N_2828);
or U3619 (N_3619,N_2780,N_2554);
or U3620 (N_3620,N_2795,N_2836);
xnor U3621 (N_3621,N_2766,N_2912);
or U3622 (N_3622,N_2590,N_1621);
nor U3623 (N_3623,N_2825,N_1714);
xnor U3624 (N_3624,N_1554,N_2760);
and U3625 (N_3625,N_2112,N_2346);
nand U3626 (N_3626,N_2755,N_1819);
and U3627 (N_3627,N_2467,N_2932);
nand U3628 (N_3628,N_1872,N_2318);
xor U3629 (N_3629,N_1580,N_2979);
and U3630 (N_3630,N_1911,N_2009);
and U3631 (N_3631,N_2821,N_2975);
xnor U3632 (N_3632,N_2338,N_2639);
xor U3633 (N_3633,N_1817,N_2306);
nand U3634 (N_3634,N_2333,N_1647);
or U3635 (N_3635,N_1739,N_1820);
and U3636 (N_3636,N_2224,N_2930);
and U3637 (N_3637,N_2900,N_2234);
xnor U3638 (N_3638,N_2908,N_1951);
nand U3639 (N_3639,N_2555,N_2285);
xnor U3640 (N_3640,N_1764,N_1984);
nor U3641 (N_3641,N_2335,N_2774);
or U3642 (N_3642,N_2546,N_2145);
xnor U3643 (N_3643,N_2666,N_2726);
and U3644 (N_3644,N_2840,N_2334);
xor U3645 (N_3645,N_2969,N_1643);
nor U3646 (N_3646,N_2714,N_2238);
nor U3647 (N_3647,N_2814,N_2834);
xnor U3648 (N_3648,N_2472,N_1584);
nand U3649 (N_3649,N_2240,N_2187);
nor U3650 (N_3650,N_2353,N_2608);
and U3651 (N_3651,N_2452,N_2631);
nand U3652 (N_3652,N_2748,N_2004);
or U3653 (N_3653,N_1890,N_2898);
nand U3654 (N_3654,N_1522,N_2055);
nor U3655 (N_3655,N_1601,N_1987);
nor U3656 (N_3656,N_2455,N_1939);
or U3657 (N_3657,N_2818,N_1854);
nor U3658 (N_3658,N_1651,N_2182);
nor U3659 (N_3659,N_2669,N_2773);
nor U3660 (N_3660,N_2890,N_1595);
and U3661 (N_3661,N_1551,N_1607);
nor U3662 (N_3662,N_2577,N_2808);
or U3663 (N_3663,N_1514,N_2806);
xor U3664 (N_3664,N_1828,N_2560);
and U3665 (N_3665,N_2781,N_1976);
and U3666 (N_3666,N_2390,N_1713);
xor U3667 (N_3667,N_2632,N_2198);
and U3668 (N_3668,N_2077,N_1591);
and U3669 (N_3669,N_2336,N_2645);
nand U3670 (N_3670,N_2746,N_1798);
nor U3671 (N_3671,N_2246,N_1765);
or U3672 (N_3672,N_1773,N_2824);
nand U3673 (N_3673,N_2999,N_1689);
or U3674 (N_3674,N_1511,N_2862);
xnor U3675 (N_3675,N_2929,N_2484);
nor U3676 (N_3676,N_1802,N_2968);
xor U3677 (N_3677,N_2738,N_2250);
xor U3678 (N_3678,N_1510,N_2137);
nand U3679 (N_3679,N_1503,N_2272);
xor U3680 (N_3680,N_2827,N_2566);
nor U3681 (N_3681,N_1953,N_1598);
or U3682 (N_3682,N_1974,N_1649);
nor U3683 (N_3683,N_2614,N_2792);
or U3684 (N_3684,N_2764,N_1874);
xnor U3685 (N_3685,N_1539,N_1806);
xor U3686 (N_3686,N_2125,N_1757);
nor U3687 (N_3687,N_2408,N_2027);
nand U3688 (N_3688,N_1529,N_2664);
nor U3689 (N_3689,N_1983,N_1971);
and U3690 (N_3690,N_2935,N_1801);
or U3691 (N_3691,N_1520,N_1567);
nand U3692 (N_3692,N_2753,N_2517);
xor U3693 (N_3693,N_1834,N_2347);
xor U3694 (N_3694,N_2514,N_2823);
nor U3695 (N_3695,N_2003,N_2428);
or U3696 (N_3696,N_2788,N_2007);
or U3697 (N_3697,N_2492,N_1622);
xor U3698 (N_3698,N_2284,N_2894);
xnor U3699 (N_3699,N_2966,N_2962);
or U3700 (N_3700,N_2707,N_1513);
xor U3701 (N_3701,N_2266,N_1715);
and U3702 (N_3702,N_2680,N_2713);
nand U3703 (N_3703,N_1923,N_1756);
nor U3704 (N_3704,N_2316,N_1877);
nand U3705 (N_3705,N_1785,N_1569);
and U3706 (N_3706,N_2490,N_1528);
xnor U3707 (N_3707,N_2122,N_2772);
nand U3708 (N_3708,N_2987,N_2214);
nand U3709 (N_3709,N_2991,N_1610);
and U3710 (N_3710,N_1891,N_1548);
or U3711 (N_3711,N_2938,N_2733);
and U3712 (N_3712,N_2729,N_2245);
nand U3713 (N_3713,N_1849,N_1800);
or U3714 (N_3714,N_1903,N_2088);
nand U3715 (N_3715,N_2783,N_1550);
nand U3716 (N_3716,N_2905,N_1921);
and U3717 (N_3717,N_1703,N_2942);
nor U3718 (N_3718,N_1716,N_2450);
xor U3719 (N_3719,N_2446,N_1899);
nor U3720 (N_3720,N_1850,N_1727);
nor U3721 (N_3721,N_2405,N_2961);
and U3722 (N_3722,N_2275,N_1581);
or U3723 (N_3723,N_2340,N_1592);
or U3724 (N_3724,N_2863,N_2050);
and U3725 (N_3725,N_1879,N_2404);
xnor U3726 (N_3726,N_2624,N_1676);
nor U3727 (N_3727,N_1931,N_2653);
nand U3728 (N_3728,N_2676,N_2523);
and U3729 (N_3729,N_2074,N_2906);
xnor U3730 (N_3730,N_1888,N_2154);
nor U3731 (N_3731,N_2076,N_2002);
nor U3732 (N_3732,N_2308,N_2933);
xnor U3733 (N_3733,N_2264,N_1993);
and U3734 (N_3734,N_2504,N_2685);
xor U3735 (N_3735,N_2671,N_1590);
or U3736 (N_3736,N_2838,N_2511);
nor U3737 (N_3737,N_2670,N_2594);
xnor U3738 (N_3738,N_1810,N_1661);
nand U3739 (N_3739,N_1855,N_2642);
nor U3740 (N_3740,N_2049,N_2495);
and U3741 (N_3741,N_2171,N_2953);
nor U3742 (N_3742,N_1506,N_1619);
and U3743 (N_3743,N_2127,N_1811);
or U3744 (N_3744,N_1754,N_2884);
nand U3745 (N_3745,N_2462,N_2722);
and U3746 (N_3746,N_1504,N_1634);
nand U3747 (N_3747,N_2869,N_2757);
nand U3748 (N_3748,N_2247,N_2040);
nor U3749 (N_3749,N_2413,N_1803);
nor U3750 (N_3750,N_2999,N_1859);
nor U3751 (N_3751,N_2346,N_2716);
and U3752 (N_3752,N_1663,N_2993);
or U3753 (N_3753,N_2395,N_2555);
nor U3754 (N_3754,N_2886,N_2372);
nor U3755 (N_3755,N_2240,N_1507);
xor U3756 (N_3756,N_2711,N_2248);
nand U3757 (N_3757,N_2296,N_1571);
and U3758 (N_3758,N_1951,N_2516);
xor U3759 (N_3759,N_2631,N_2797);
nand U3760 (N_3760,N_1535,N_2150);
and U3761 (N_3761,N_1517,N_2543);
nand U3762 (N_3762,N_2384,N_2438);
and U3763 (N_3763,N_2276,N_1862);
and U3764 (N_3764,N_2719,N_2753);
xor U3765 (N_3765,N_2462,N_2896);
nand U3766 (N_3766,N_2169,N_2802);
xnor U3767 (N_3767,N_2712,N_1660);
or U3768 (N_3768,N_1596,N_2146);
nand U3769 (N_3769,N_1634,N_2493);
or U3770 (N_3770,N_2762,N_1707);
or U3771 (N_3771,N_2468,N_2007);
nor U3772 (N_3772,N_2184,N_2479);
nand U3773 (N_3773,N_1685,N_2915);
xnor U3774 (N_3774,N_2921,N_2392);
xor U3775 (N_3775,N_1874,N_2652);
xor U3776 (N_3776,N_2238,N_1772);
nand U3777 (N_3777,N_2602,N_2977);
nor U3778 (N_3778,N_2655,N_2680);
xor U3779 (N_3779,N_2800,N_1592);
and U3780 (N_3780,N_2729,N_1954);
nand U3781 (N_3781,N_2061,N_1633);
or U3782 (N_3782,N_1638,N_2621);
nand U3783 (N_3783,N_2913,N_1723);
nor U3784 (N_3784,N_2010,N_2837);
or U3785 (N_3785,N_1658,N_2200);
or U3786 (N_3786,N_2604,N_1983);
and U3787 (N_3787,N_2103,N_2794);
xnor U3788 (N_3788,N_2209,N_1529);
and U3789 (N_3789,N_2200,N_2185);
nand U3790 (N_3790,N_2808,N_1608);
nor U3791 (N_3791,N_1899,N_2484);
or U3792 (N_3792,N_2967,N_2618);
xnor U3793 (N_3793,N_1635,N_1900);
nand U3794 (N_3794,N_2317,N_1923);
nor U3795 (N_3795,N_2599,N_2319);
xnor U3796 (N_3796,N_2820,N_2090);
or U3797 (N_3797,N_1560,N_2104);
nor U3798 (N_3798,N_2518,N_2969);
or U3799 (N_3799,N_2099,N_2438);
nor U3800 (N_3800,N_1607,N_2753);
xnor U3801 (N_3801,N_2643,N_1639);
xnor U3802 (N_3802,N_1665,N_2181);
or U3803 (N_3803,N_2419,N_1988);
nor U3804 (N_3804,N_2617,N_2023);
xor U3805 (N_3805,N_1934,N_1718);
or U3806 (N_3806,N_2341,N_2262);
and U3807 (N_3807,N_2337,N_2015);
xnor U3808 (N_3808,N_1896,N_2809);
nor U3809 (N_3809,N_1884,N_1895);
or U3810 (N_3810,N_1864,N_2114);
and U3811 (N_3811,N_1738,N_2661);
nand U3812 (N_3812,N_1935,N_2642);
and U3813 (N_3813,N_2379,N_2830);
or U3814 (N_3814,N_2397,N_2271);
and U3815 (N_3815,N_2497,N_2346);
xnor U3816 (N_3816,N_2356,N_2639);
nor U3817 (N_3817,N_1699,N_2045);
xnor U3818 (N_3818,N_2017,N_1793);
xor U3819 (N_3819,N_2640,N_2907);
and U3820 (N_3820,N_2029,N_1859);
nand U3821 (N_3821,N_1843,N_2402);
xor U3822 (N_3822,N_2152,N_2600);
xnor U3823 (N_3823,N_1960,N_2476);
and U3824 (N_3824,N_2321,N_2497);
nor U3825 (N_3825,N_2407,N_2349);
nor U3826 (N_3826,N_1863,N_2722);
or U3827 (N_3827,N_1642,N_1865);
nand U3828 (N_3828,N_2946,N_1601);
or U3829 (N_3829,N_1648,N_2124);
nand U3830 (N_3830,N_1739,N_1955);
or U3831 (N_3831,N_2144,N_2450);
xnor U3832 (N_3832,N_1852,N_1708);
or U3833 (N_3833,N_2258,N_1913);
nor U3834 (N_3834,N_1949,N_2909);
or U3835 (N_3835,N_2850,N_2074);
xnor U3836 (N_3836,N_2933,N_2558);
nand U3837 (N_3837,N_2476,N_2718);
nand U3838 (N_3838,N_2415,N_2233);
nor U3839 (N_3839,N_1691,N_1885);
and U3840 (N_3840,N_2723,N_1634);
xnor U3841 (N_3841,N_2360,N_2054);
and U3842 (N_3842,N_1506,N_1885);
xor U3843 (N_3843,N_1568,N_2608);
and U3844 (N_3844,N_2358,N_2750);
or U3845 (N_3845,N_2491,N_2679);
xnor U3846 (N_3846,N_2723,N_1830);
nand U3847 (N_3847,N_2003,N_2924);
xnor U3848 (N_3848,N_2071,N_2463);
xor U3849 (N_3849,N_1915,N_2571);
or U3850 (N_3850,N_1808,N_1636);
and U3851 (N_3851,N_2439,N_2580);
nand U3852 (N_3852,N_2325,N_1960);
and U3853 (N_3853,N_2034,N_2268);
nor U3854 (N_3854,N_1899,N_1658);
xnor U3855 (N_3855,N_2017,N_1648);
nor U3856 (N_3856,N_2562,N_1860);
nor U3857 (N_3857,N_2979,N_1969);
or U3858 (N_3858,N_2179,N_2115);
nand U3859 (N_3859,N_2263,N_2700);
nand U3860 (N_3860,N_2752,N_2285);
nand U3861 (N_3861,N_2536,N_2892);
nand U3862 (N_3862,N_2343,N_1709);
and U3863 (N_3863,N_2597,N_2276);
xor U3864 (N_3864,N_2290,N_2269);
nor U3865 (N_3865,N_1527,N_2625);
xor U3866 (N_3866,N_2349,N_2602);
and U3867 (N_3867,N_1806,N_2083);
or U3868 (N_3868,N_2496,N_2962);
xor U3869 (N_3869,N_1948,N_2320);
xnor U3870 (N_3870,N_2112,N_1670);
nand U3871 (N_3871,N_2777,N_2539);
nor U3872 (N_3872,N_2743,N_1868);
nand U3873 (N_3873,N_2431,N_2803);
xor U3874 (N_3874,N_2270,N_2799);
and U3875 (N_3875,N_1598,N_2112);
nand U3876 (N_3876,N_2201,N_2982);
xnor U3877 (N_3877,N_1752,N_2723);
xor U3878 (N_3878,N_2955,N_1817);
and U3879 (N_3879,N_2639,N_2317);
and U3880 (N_3880,N_2863,N_1965);
nor U3881 (N_3881,N_2392,N_2616);
nor U3882 (N_3882,N_1668,N_2486);
and U3883 (N_3883,N_2964,N_2313);
or U3884 (N_3884,N_2572,N_2303);
nand U3885 (N_3885,N_2304,N_2702);
or U3886 (N_3886,N_2964,N_1734);
or U3887 (N_3887,N_2763,N_2394);
xnor U3888 (N_3888,N_1622,N_2652);
xnor U3889 (N_3889,N_1703,N_2296);
nor U3890 (N_3890,N_2190,N_2718);
xnor U3891 (N_3891,N_2508,N_2608);
nor U3892 (N_3892,N_2808,N_1536);
xnor U3893 (N_3893,N_2768,N_1709);
or U3894 (N_3894,N_2239,N_1704);
and U3895 (N_3895,N_2765,N_1666);
nor U3896 (N_3896,N_2128,N_2256);
nand U3897 (N_3897,N_1512,N_1985);
nand U3898 (N_3898,N_2099,N_2839);
and U3899 (N_3899,N_1591,N_2199);
nand U3900 (N_3900,N_2514,N_2490);
nand U3901 (N_3901,N_2534,N_2008);
nand U3902 (N_3902,N_2166,N_2258);
xnor U3903 (N_3903,N_2206,N_2806);
xor U3904 (N_3904,N_2720,N_1728);
nor U3905 (N_3905,N_2754,N_2854);
or U3906 (N_3906,N_1971,N_2844);
nand U3907 (N_3907,N_1867,N_2341);
nand U3908 (N_3908,N_2318,N_1674);
nand U3909 (N_3909,N_2019,N_1711);
or U3910 (N_3910,N_1704,N_2548);
nor U3911 (N_3911,N_2420,N_2443);
xnor U3912 (N_3912,N_1898,N_2237);
and U3913 (N_3913,N_1695,N_1811);
nor U3914 (N_3914,N_2358,N_2474);
nor U3915 (N_3915,N_2393,N_2628);
and U3916 (N_3916,N_2199,N_1865);
xnor U3917 (N_3917,N_2761,N_1841);
xor U3918 (N_3918,N_2315,N_1808);
and U3919 (N_3919,N_2334,N_1934);
nor U3920 (N_3920,N_1619,N_2073);
nand U3921 (N_3921,N_1862,N_1839);
and U3922 (N_3922,N_2737,N_2871);
nand U3923 (N_3923,N_2044,N_1640);
and U3924 (N_3924,N_1729,N_1807);
nor U3925 (N_3925,N_2363,N_2336);
nand U3926 (N_3926,N_2261,N_1727);
nand U3927 (N_3927,N_2988,N_2811);
xnor U3928 (N_3928,N_2260,N_2314);
and U3929 (N_3929,N_2951,N_1552);
nor U3930 (N_3930,N_1872,N_1811);
nand U3931 (N_3931,N_2730,N_1874);
xnor U3932 (N_3932,N_1818,N_2144);
nand U3933 (N_3933,N_2025,N_1599);
xor U3934 (N_3934,N_2974,N_2936);
nor U3935 (N_3935,N_2799,N_1886);
nand U3936 (N_3936,N_2640,N_2312);
nand U3937 (N_3937,N_2347,N_2825);
and U3938 (N_3938,N_2065,N_2133);
or U3939 (N_3939,N_2248,N_2002);
nor U3940 (N_3940,N_2880,N_1938);
and U3941 (N_3941,N_1767,N_2907);
xnor U3942 (N_3942,N_1517,N_2008);
and U3943 (N_3943,N_2070,N_2114);
and U3944 (N_3944,N_1903,N_2795);
nor U3945 (N_3945,N_1715,N_1719);
and U3946 (N_3946,N_2204,N_1671);
and U3947 (N_3947,N_1542,N_2222);
nand U3948 (N_3948,N_2202,N_2551);
or U3949 (N_3949,N_1860,N_2446);
nor U3950 (N_3950,N_2348,N_2530);
nand U3951 (N_3951,N_2710,N_2107);
nor U3952 (N_3952,N_2497,N_2803);
or U3953 (N_3953,N_2618,N_2361);
xor U3954 (N_3954,N_1749,N_1978);
nor U3955 (N_3955,N_2896,N_2181);
nor U3956 (N_3956,N_2049,N_1933);
or U3957 (N_3957,N_1500,N_2301);
or U3958 (N_3958,N_2868,N_1649);
nand U3959 (N_3959,N_2371,N_2994);
nor U3960 (N_3960,N_1573,N_2656);
nand U3961 (N_3961,N_2201,N_1829);
and U3962 (N_3962,N_2883,N_1783);
xor U3963 (N_3963,N_2690,N_1569);
xor U3964 (N_3964,N_1961,N_1693);
and U3965 (N_3965,N_1756,N_1983);
nor U3966 (N_3966,N_2930,N_2030);
nor U3967 (N_3967,N_2690,N_1986);
nand U3968 (N_3968,N_1550,N_2324);
nor U3969 (N_3969,N_2502,N_2423);
and U3970 (N_3970,N_2290,N_2715);
and U3971 (N_3971,N_2424,N_2417);
and U3972 (N_3972,N_2512,N_2127);
and U3973 (N_3973,N_2294,N_2611);
nor U3974 (N_3974,N_1907,N_1858);
and U3975 (N_3975,N_2663,N_1630);
nand U3976 (N_3976,N_2921,N_1659);
nand U3977 (N_3977,N_1566,N_2791);
and U3978 (N_3978,N_1536,N_2124);
xor U3979 (N_3979,N_2961,N_2456);
or U3980 (N_3980,N_2276,N_2160);
nor U3981 (N_3981,N_2551,N_2172);
nor U3982 (N_3982,N_2583,N_2373);
nand U3983 (N_3983,N_2836,N_2374);
or U3984 (N_3984,N_2379,N_2276);
nor U3985 (N_3985,N_2852,N_2451);
and U3986 (N_3986,N_2181,N_2471);
and U3987 (N_3987,N_2310,N_2628);
xnor U3988 (N_3988,N_2516,N_2024);
and U3989 (N_3989,N_1673,N_2169);
xnor U3990 (N_3990,N_2181,N_2656);
xor U3991 (N_3991,N_1608,N_2551);
or U3992 (N_3992,N_1779,N_2311);
nor U3993 (N_3993,N_2529,N_1717);
nor U3994 (N_3994,N_1663,N_2764);
xor U3995 (N_3995,N_2816,N_2225);
nand U3996 (N_3996,N_1728,N_2955);
or U3997 (N_3997,N_2197,N_1985);
nand U3998 (N_3998,N_2271,N_1629);
and U3999 (N_3999,N_1778,N_1691);
nor U4000 (N_4000,N_2366,N_2387);
and U4001 (N_4001,N_2395,N_1765);
nand U4002 (N_4002,N_2561,N_1617);
nand U4003 (N_4003,N_2791,N_2407);
or U4004 (N_4004,N_1906,N_1972);
nand U4005 (N_4005,N_2424,N_2480);
or U4006 (N_4006,N_2562,N_2662);
nand U4007 (N_4007,N_2974,N_2446);
and U4008 (N_4008,N_2898,N_1934);
nor U4009 (N_4009,N_2501,N_2614);
and U4010 (N_4010,N_2872,N_1571);
or U4011 (N_4011,N_2438,N_1684);
nand U4012 (N_4012,N_2945,N_2172);
or U4013 (N_4013,N_2756,N_1696);
and U4014 (N_4014,N_2032,N_2970);
xnor U4015 (N_4015,N_2988,N_1685);
nor U4016 (N_4016,N_2798,N_2905);
nor U4017 (N_4017,N_2447,N_2277);
or U4018 (N_4018,N_2919,N_2717);
nor U4019 (N_4019,N_2705,N_1842);
nand U4020 (N_4020,N_1820,N_2845);
and U4021 (N_4021,N_1576,N_2552);
or U4022 (N_4022,N_1682,N_2920);
xor U4023 (N_4023,N_1679,N_1633);
nand U4024 (N_4024,N_1504,N_2216);
nand U4025 (N_4025,N_2353,N_1570);
and U4026 (N_4026,N_1656,N_2907);
xnor U4027 (N_4027,N_2003,N_2832);
or U4028 (N_4028,N_1925,N_2168);
nand U4029 (N_4029,N_2475,N_1695);
xor U4030 (N_4030,N_1613,N_2158);
xor U4031 (N_4031,N_2705,N_2607);
and U4032 (N_4032,N_2889,N_1587);
xor U4033 (N_4033,N_2200,N_2183);
and U4034 (N_4034,N_1693,N_1836);
and U4035 (N_4035,N_2873,N_2759);
nor U4036 (N_4036,N_2013,N_1501);
or U4037 (N_4037,N_2974,N_2162);
nand U4038 (N_4038,N_2743,N_1924);
or U4039 (N_4039,N_2619,N_1925);
nor U4040 (N_4040,N_1698,N_2528);
xnor U4041 (N_4041,N_1928,N_2524);
nor U4042 (N_4042,N_2279,N_2321);
nand U4043 (N_4043,N_2674,N_1890);
and U4044 (N_4044,N_2845,N_2336);
nand U4045 (N_4045,N_2146,N_2113);
xnor U4046 (N_4046,N_1602,N_2448);
xnor U4047 (N_4047,N_2071,N_2404);
and U4048 (N_4048,N_2860,N_1847);
nand U4049 (N_4049,N_2919,N_2772);
or U4050 (N_4050,N_1971,N_2791);
and U4051 (N_4051,N_1729,N_1589);
nand U4052 (N_4052,N_2368,N_2448);
nor U4053 (N_4053,N_2142,N_2200);
nor U4054 (N_4054,N_1757,N_1672);
nor U4055 (N_4055,N_2373,N_1717);
and U4056 (N_4056,N_2146,N_2718);
and U4057 (N_4057,N_1657,N_1767);
nor U4058 (N_4058,N_2276,N_2446);
nor U4059 (N_4059,N_2035,N_1987);
nor U4060 (N_4060,N_1634,N_1920);
and U4061 (N_4061,N_2272,N_2993);
nor U4062 (N_4062,N_1530,N_2461);
xnor U4063 (N_4063,N_2011,N_1938);
nand U4064 (N_4064,N_1966,N_2886);
and U4065 (N_4065,N_2703,N_2498);
nand U4066 (N_4066,N_1601,N_2997);
xnor U4067 (N_4067,N_2990,N_1994);
nand U4068 (N_4068,N_2714,N_2938);
xnor U4069 (N_4069,N_2555,N_1912);
xor U4070 (N_4070,N_2311,N_2933);
or U4071 (N_4071,N_1759,N_1957);
nor U4072 (N_4072,N_1933,N_2384);
or U4073 (N_4073,N_2849,N_2777);
or U4074 (N_4074,N_1563,N_1790);
xor U4075 (N_4075,N_2352,N_1783);
nor U4076 (N_4076,N_1811,N_1501);
nor U4077 (N_4077,N_1970,N_2159);
or U4078 (N_4078,N_2195,N_1669);
xor U4079 (N_4079,N_2247,N_2166);
and U4080 (N_4080,N_2810,N_1575);
nand U4081 (N_4081,N_2730,N_1784);
nand U4082 (N_4082,N_1746,N_2042);
or U4083 (N_4083,N_2863,N_2347);
or U4084 (N_4084,N_2318,N_2966);
nand U4085 (N_4085,N_2425,N_2505);
and U4086 (N_4086,N_2362,N_1819);
or U4087 (N_4087,N_1749,N_1541);
nor U4088 (N_4088,N_2965,N_2827);
and U4089 (N_4089,N_1576,N_1692);
and U4090 (N_4090,N_1794,N_2919);
nand U4091 (N_4091,N_1782,N_2734);
nand U4092 (N_4092,N_2945,N_2511);
and U4093 (N_4093,N_1930,N_2660);
nand U4094 (N_4094,N_1549,N_2304);
or U4095 (N_4095,N_1801,N_1536);
and U4096 (N_4096,N_2839,N_1835);
and U4097 (N_4097,N_2578,N_1539);
nand U4098 (N_4098,N_1694,N_2598);
xnor U4099 (N_4099,N_1904,N_2879);
or U4100 (N_4100,N_1689,N_2572);
or U4101 (N_4101,N_2664,N_1721);
nand U4102 (N_4102,N_2564,N_2783);
or U4103 (N_4103,N_2470,N_2452);
and U4104 (N_4104,N_1681,N_2937);
nor U4105 (N_4105,N_2870,N_1543);
nor U4106 (N_4106,N_2499,N_2931);
or U4107 (N_4107,N_2569,N_2107);
nor U4108 (N_4108,N_2814,N_2235);
nand U4109 (N_4109,N_2680,N_1894);
nand U4110 (N_4110,N_1939,N_1888);
and U4111 (N_4111,N_1693,N_2318);
or U4112 (N_4112,N_2737,N_1703);
nand U4113 (N_4113,N_1968,N_2639);
or U4114 (N_4114,N_1509,N_2835);
and U4115 (N_4115,N_2574,N_2563);
xnor U4116 (N_4116,N_1938,N_1992);
or U4117 (N_4117,N_2813,N_2146);
and U4118 (N_4118,N_1725,N_2376);
or U4119 (N_4119,N_2155,N_1871);
and U4120 (N_4120,N_2144,N_2382);
nor U4121 (N_4121,N_2151,N_2082);
xnor U4122 (N_4122,N_1678,N_2059);
and U4123 (N_4123,N_1904,N_2918);
or U4124 (N_4124,N_2906,N_2188);
nand U4125 (N_4125,N_1738,N_2209);
or U4126 (N_4126,N_2998,N_1539);
nand U4127 (N_4127,N_2195,N_2157);
xnor U4128 (N_4128,N_1784,N_2501);
or U4129 (N_4129,N_2901,N_2442);
or U4130 (N_4130,N_2485,N_2104);
xor U4131 (N_4131,N_2075,N_2791);
nor U4132 (N_4132,N_2330,N_1615);
and U4133 (N_4133,N_2901,N_2140);
nand U4134 (N_4134,N_2814,N_1791);
nand U4135 (N_4135,N_1865,N_2878);
nand U4136 (N_4136,N_2514,N_1883);
and U4137 (N_4137,N_2925,N_2880);
nor U4138 (N_4138,N_1577,N_1726);
xnor U4139 (N_4139,N_1501,N_2715);
xor U4140 (N_4140,N_2177,N_2582);
nand U4141 (N_4141,N_1542,N_1768);
and U4142 (N_4142,N_1530,N_1615);
xnor U4143 (N_4143,N_2849,N_1982);
nor U4144 (N_4144,N_2336,N_2041);
nor U4145 (N_4145,N_1902,N_1916);
nor U4146 (N_4146,N_2799,N_1847);
xor U4147 (N_4147,N_2164,N_1922);
and U4148 (N_4148,N_2412,N_1734);
xor U4149 (N_4149,N_1508,N_2273);
and U4150 (N_4150,N_1703,N_2533);
nor U4151 (N_4151,N_2050,N_2332);
xnor U4152 (N_4152,N_1810,N_2383);
nand U4153 (N_4153,N_2908,N_2811);
xor U4154 (N_4154,N_2178,N_2885);
xor U4155 (N_4155,N_2053,N_2533);
xor U4156 (N_4156,N_2974,N_2422);
and U4157 (N_4157,N_2494,N_2094);
nor U4158 (N_4158,N_1986,N_1896);
xor U4159 (N_4159,N_2518,N_2900);
or U4160 (N_4160,N_1991,N_2036);
nor U4161 (N_4161,N_1685,N_2701);
or U4162 (N_4162,N_1582,N_2450);
and U4163 (N_4163,N_2629,N_1643);
nor U4164 (N_4164,N_2734,N_2868);
or U4165 (N_4165,N_1560,N_2882);
nor U4166 (N_4166,N_2554,N_2647);
nand U4167 (N_4167,N_1506,N_1909);
xor U4168 (N_4168,N_2770,N_2113);
and U4169 (N_4169,N_2217,N_2050);
and U4170 (N_4170,N_2423,N_1970);
xor U4171 (N_4171,N_2724,N_2632);
nand U4172 (N_4172,N_2236,N_2729);
xnor U4173 (N_4173,N_2736,N_1571);
nor U4174 (N_4174,N_2995,N_2023);
nor U4175 (N_4175,N_2717,N_2303);
and U4176 (N_4176,N_1709,N_2742);
xnor U4177 (N_4177,N_1590,N_1635);
or U4178 (N_4178,N_1783,N_2110);
nor U4179 (N_4179,N_2520,N_2431);
nand U4180 (N_4180,N_2555,N_2826);
nor U4181 (N_4181,N_2276,N_2299);
and U4182 (N_4182,N_2488,N_1897);
xor U4183 (N_4183,N_2144,N_2308);
xnor U4184 (N_4184,N_1777,N_2931);
and U4185 (N_4185,N_2143,N_1650);
or U4186 (N_4186,N_2372,N_2678);
and U4187 (N_4187,N_2887,N_1753);
nor U4188 (N_4188,N_2908,N_2483);
nand U4189 (N_4189,N_2043,N_1516);
or U4190 (N_4190,N_2290,N_2830);
nor U4191 (N_4191,N_1709,N_2417);
and U4192 (N_4192,N_2432,N_2605);
nand U4193 (N_4193,N_2425,N_2265);
or U4194 (N_4194,N_2290,N_2212);
nand U4195 (N_4195,N_2170,N_1905);
nand U4196 (N_4196,N_2179,N_1565);
xnor U4197 (N_4197,N_1842,N_2054);
xnor U4198 (N_4198,N_2829,N_2575);
nor U4199 (N_4199,N_2579,N_1671);
xnor U4200 (N_4200,N_1572,N_2414);
and U4201 (N_4201,N_2140,N_1502);
nor U4202 (N_4202,N_1979,N_1607);
nor U4203 (N_4203,N_2600,N_2819);
and U4204 (N_4204,N_2260,N_2788);
xor U4205 (N_4205,N_2083,N_2473);
or U4206 (N_4206,N_1625,N_2344);
or U4207 (N_4207,N_2690,N_2881);
or U4208 (N_4208,N_1833,N_2116);
and U4209 (N_4209,N_1788,N_1741);
nor U4210 (N_4210,N_1941,N_2675);
nor U4211 (N_4211,N_2780,N_2955);
nand U4212 (N_4212,N_2751,N_2094);
nor U4213 (N_4213,N_2763,N_2969);
nor U4214 (N_4214,N_2067,N_1758);
or U4215 (N_4215,N_2122,N_2333);
nand U4216 (N_4216,N_2012,N_1516);
xor U4217 (N_4217,N_1765,N_2286);
and U4218 (N_4218,N_1815,N_1693);
or U4219 (N_4219,N_1594,N_2757);
nand U4220 (N_4220,N_2093,N_2807);
xnor U4221 (N_4221,N_1547,N_2836);
and U4222 (N_4222,N_1989,N_2473);
nor U4223 (N_4223,N_2455,N_1584);
xor U4224 (N_4224,N_2872,N_2179);
or U4225 (N_4225,N_2409,N_2068);
and U4226 (N_4226,N_2756,N_1748);
xor U4227 (N_4227,N_2600,N_2590);
nor U4228 (N_4228,N_2369,N_1678);
nor U4229 (N_4229,N_1736,N_2816);
and U4230 (N_4230,N_1730,N_2200);
or U4231 (N_4231,N_2901,N_1622);
and U4232 (N_4232,N_2344,N_2811);
nor U4233 (N_4233,N_2237,N_1556);
nand U4234 (N_4234,N_1956,N_2106);
and U4235 (N_4235,N_1585,N_2420);
xnor U4236 (N_4236,N_2666,N_2299);
or U4237 (N_4237,N_2156,N_2948);
and U4238 (N_4238,N_2518,N_1631);
and U4239 (N_4239,N_2382,N_2540);
xor U4240 (N_4240,N_1748,N_2580);
or U4241 (N_4241,N_2527,N_1657);
nand U4242 (N_4242,N_2861,N_1902);
nand U4243 (N_4243,N_1712,N_2427);
nand U4244 (N_4244,N_2026,N_2445);
and U4245 (N_4245,N_2799,N_2160);
nand U4246 (N_4246,N_2918,N_2673);
or U4247 (N_4247,N_2379,N_2253);
nor U4248 (N_4248,N_2661,N_2909);
xnor U4249 (N_4249,N_2784,N_2578);
nand U4250 (N_4250,N_2767,N_2709);
nand U4251 (N_4251,N_2629,N_2132);
nor U4252 (N_4252,N_2771,N_2398);
nand U4253 (N_4253,N_1594,N_1708);
nand U4254 (N_4254,N_1755,N_2291);
nor U4255 (N_4255,N_1905,N_1851);
xor U4256 (N_4256,N_2977,N_2415);
xor U4257 (N_4257,N_2189,N_1681);
or U4258 (N_4258,N_1970,N_2950);
nand U4259 (N_4259,N_2857,N_2139);
nand U4260 (N_4260,N_1698,N_2087);
and U4261 (N_4261,N_1671,N_1903);
xnor U4262 (N_4262,N_2332,N_1604);
and U4263 (N_4263,N_2362,N_2274);
or U4264 (N_4264,N_1867,N_2039);
nor U4265 (N_4265,N_1976,N_2231);
nand U4266 (N_4266,N_2075,N_2395);
xnor U4267 (N_4267,N_1644,N_2530);
nor U4268 (N_4268,N_1615,N_2120);
nor U4269 (N_4269,N_1946,N_2268);
nand U4270 (N_4270,N_1733,N_2624);
nor U4271 (N_4271,N_2712,N_2541);
nor U4272 (N_4272,N_2805,N_1825);
xor U4273 (N_4273,N_2881,N_2629);
and U4274 (N_4274,N_2513,N_1709);
nor U4275 (N_4275,N_1891,N_2098);
xnor U4276 (N_4276,N_2552,N_1959);
and U4277 (N_4277,N_2424,N_1843);
nand U4278 (N_4278,N_2574,N_2497);
and U4279 (N_4279,N_1789,N_2003);
nand U4280 (N_4280,N_2549,N_2597);
or U4281 (N_4281,N_2574,N_1838);
nor U4282 (N_4282,N_1993,N_2419);
nand U4283 (N_4283,N_1878,N_1722);
xor U4284 (N_4284,N_2290,N_2097);
nand U4285 (N_4285,N_2525,N_1835);
xor U4286 (N_4286,N_1613,N_1778);
or U4287 (N_4287,N_2422,N_2945);
and U4288 (N_4288,N_2870,N_1942);
nand U4289 (N_4289,N_2890,N_2461);
or U4290 (N_4290,N_1840,N_2089);
nand U4291 (N_4291,N_1549,N_2165);
nand U4292 (N_4292,N_1740,N_2128);
nand U4293 (N_4293,N_1820,N_2152);
and U4294 (N_4294,N_2005,N_2964);
and U4295 (N_4295,N_1554,N_2164);
nand U4296 (N_4296,N_2723,N_2810);
or U4297 (N_4297,N_2968,N_1816);
xnor U4298 (N_4298,N_1675,N_2661);
nor U4299 (N_4299,N_2182,N_2814);
and U4300 (N_4300,N_1546,N_1971);
or U4301 (N_4301,N_1688,N_1610);
or U4302 (N_4302,N_2604,N_2706);
or U4303 (N_4303,N_2165,N_1917);
and U4304 (N_4304,N_1900,N_2273);
xor U4305 (N_4305,N_2660,N_2891);
nand U4306 (N_4306,N_2165,N_2300);
nand U4307 (N_4307,N_2134,N_2456);
and U4308 (N_4308,N_2108,N_2730);
and U4309 (N_4309,N_1724,N_2289);
xor U4310 (N_4310,N_2262,N_2217);
and U4311 (N_4311,N_2759,N_2160);
nand U4312 (N_4312,N_2669,N_2198);
or U4313 (N_4313,N_2918,N_1546);
nor U4314 (N_4314,N_2097,N_1990);
and U4315 (N_4315,N_2201,N_2789);
or U4316 (N_4316,N_2965,N_1933);
nor U4317 (N_4317,N_2102,N_2872);
and U4318 (N_4318,N_2645,N_1636);
and U4319 (N_4319,N_2325,N_2241);
xnor U4320 (N_4320,N_2645,N_1528);
xnor U4321 (N_4321,N_1760,N_2672);
xor U4322 (N_4322,N_1710,N_2560);
nand U4323 (N_4323,N_2070,N_1683);
xnor U4324 (N_4324,N_2109,N_2144);
or U4325 (N_4325,N_2625,N_2981);
xnor U4326 (N_4326,N_1811,N_2141);
xnor U4327 (N_4327,N_2630,N_2423);
nor U4328 (N_4328,N_2853,N_1949);
and U4329 (N_4329,N_2589,N_2623);
nand U4330 (N_4330,N_1618,N_1827);
xnor U4331 (N_4331,N_2681,N_1576);
or U4332 (N_4332,N_1906,N_2756);
or U4333 (N_4333,N_1540,N_2919);
xnor U4334 (N_4334,N_2130,N_2242);
nor U4335 (N_4335,N_2404,N_1671);
or U4336 (N_4336,N_1735,N_2112);
xnor U4337 (N_4337,N_2520,N_1501);
or U4338 (N_4338,N_1957,N_2028);
or U4339 (N_4339,N_1977,N_2529);
xnor U4340 (N_4340,N_1606,N_2604);
nand U4341 (N_4341,N_2522,N_2395);
or U4342 (N_4342,N_2448,N_2494);
nor U4343 (N_4343,N_2215,N_2833);
nand U4344 (N_4344,N_1771,N_2296);
nand U4345 (N_4345,N_2725,N_2203);
and U4346 (N_4346,N_1515,N_2765);
or U4347 (N_4347,N_1654,N_1698);
xor U4348 (N_4348,N_2132,N_2324);
and U4349 (N_4349,N_1611,N_2589);
xnor U4350 (N_4350,N_2987,N_2328);
xnor U4351 (N_4351,N_1824,N_1798);
nor U4352 (N_4352,N_1891,N_2515);
nor U4353 (N_4353,N_2786,N_1807);
and U4354 (N_4354,N_1725,N_2135);
nor U4355 (N_4355,N_2966,N_2385);
nand U4356 (N_4356,N_2571,N_1865);
xor U4357 (N_4357,N_2293,N_1501);
or U4358 (N_4358,N_1647,N_1530);
xor U4359 (N_4359,N_2396,N_2563);
nor U4360 (N_4360,N_2932,N_2521);
nand U4361 (N_4361,N_2088,N_1791);
and U4362 (N_4362,N_2240,N_1732);
or U4363 (N_4363,N_2838,N_2395);
and U4364 (N_4364,N_2525,N_1650);
nand U4365 (N_4365,N_2585,N_1579);
xor U4366 (N_4366,N_2358,N_1776);
nand U4367 (N_4367,N_2616,N_1989);
and U4368 (N_4368,N_2665,N_2995);
nor U4369 (N_4369,N_2451,N_2002);
or U4370 (N_4370,N_2218,N_1842);
or U4371 (N_4371,N_2573,N_2065);
or U4372 (N_4372,N_2004,N_2508);
nand U4373 (N_4373,N_2667,N_2911);
xnor U4374 (N_4374,N_2314,N_1672);
nand U4375 (N_4375,N_2933,N_2025);
xor U4376 (N_4376,N_1767,N_2553);
xnor U4377 (N_4377,N_2813,N_2041);
xor U4378 (N_4378,N_2162,N_2203);
or U4379 (N_4379,N_2279,N_2588);
or U4380 (N_4380,N_2332,N_2331);
or U4381 (N_4381,N_2147,N_2073);
or U4382 (N_4382,N_2852,N_2204);
and U4383 (N_4383,N_1859,N_2218);
and U4384 (N_4384,N_2517,N_2675);
xnor U4385 (N_4385,N_2045,N_1507);
and U4386 (N_4386,N_1638,N_1568);
and U4387 (N_4387,N_2573,N_2645);
and U4388 (N_4388,N_1813,N_2814);
and U4389 (N_4389,N_2637,N_2827);
nor U4390 (N_4390,N_1644,N_1577);
or U4391 (N_4391,N_2125,N_2407);
and U4392 (N_4392,N_2080,N_1707);
xnor U4393 (N_4393,N_2920,N_1817);
xnor U4394 (N_4394,N_2469,N_1839);
and U4395 (N_4395,N_2426,N_1841);
nor U4396 (N_4396,N_1662,N_2559);
or U4397 (N_4397,N_1779,N_2480);
or U4398 (N_4398,N_2471,N_2660);
nand U4399 (N_4399,N_1686,N_2202);
nand U4400 (N_4400,N_2581,N_2785);
nor U4401 (N_4401,N_2877,N_1932);
and U4402 (N_4402,N_2943,N_2477);
xor U4403 (N_4403,N_2881,N_1526);
nor U4404 (N_4404,N_2051,N_1773);
nor U4405 (N_4405,N_1651,N_2107);
xor U4406 (N_4406,N_2646,N_2577);
or U4407 (N_4407,N_2968,N_1541);
nor U4408 (N_4408,N_2087,N_1849);
nand U4409 (N_4409,N_2523,N_1971);
or U4410 (N_4410,N_1707,N_2283);
xnor U4411 (N_4411,N_1961,N_2142);
xor U4412 (N_4412,N_1860,N_2290);
xnor U4413 (N_4413,N_1713,N_2164);
and U4414 (N_4414,N_1683,N_2125);
xnor U4415 (N_4415,N_2099,N_2368);
or U4416 (N_4416,N_2822,N_2572);
or U4417 (N_4417,N_1707,N_2119);
xnor U4418 (N_4418,N_1693,N_2332);
and U4419 (N_4419,N_2677,N_2899);
xor U4420 (N_4420,N_1592,N_1541);
nand U4421 (N_4421,N_1543,N_2462);
or U4422 (N_4422,N_2643,N_1783);
xor U4423 (N_4423,N_1782,N_1944);
and U4424 (N_4424,N_1767,N_1947);
nand U4425 (N_4425,N_2522,N_2002);
nor U4426 (N_4426,N_1555,N_2344);
and U4427 (N_4427,N_1598,N_2868);
or U4428 (N_4428,N_2977,N_1736);
or U4429 (N_4429,N_1636,N_1696);
or U4430 (N_4430,N_1726,N_1651);
nand U4431 (N_4431,N_1983,N_2878);
xor U4432 (N_4432,N_1518,N_2440);
nand U4433 (N_4433,N_1733,N_2710);
or U4434 (N_4434,N_2253,N_1824);
xor U4435 (N_4435,N_2968,N_2788);
nor U4436 (N_4436,N_1869,N_1904);
nor U4437 (N_4437,N_1514,N_2383);
xnor U4438 (N_4438,N_2063,N_2881);
nand U4439 (N_4439,N_2345,N_2976);
or U4440 (N_4440,N_1536,N_2607);
or U4441 (N_4441,N_2387,N_1827);
nor U4442 (N_4442,N_1754,N_2699);
or U4443 (N_4443,N_2609,N_1810);
xor U4444 (N_4444,N_2494,N_2541);
nand U4445 (N_4445,N_1587,N_1785);
nor U4446 (N_4446,N_2005,N_1893);
xor U4447 (N_4447,N_2382,N_2628);
xor U4448 (N_4448,N_2305,N_1759);
or U4449 (N_4449,N_2894,N_2247);
nand U4450 (N_4450,N_2793,N_2875);
nand U4451 (N_4451,N_1921,N_2073);
or U4452 (N_4452,N_2978,N_2465);
nor U4453 (N_4453,N_2981,N_1911);
nor U4454 (N_4454,N_1680,N_1632);
nor U4455 (N_4455,N_2059,N_2831);
or U4456 (N_4456,N_2411,N_1692);
nor U4457 (N_4457,N_2818,N_2330);
nor U4458 (N_4458,N_2376,N_2239);
nand U4459 (N_4459,N_1880,N_1912);
or U4460 (N_4460,N_1722,N_1968);
xor U4461 (N_4461,N_2407,N_2924);
nand U4462 (N_4462,N_1732,N_2043);
xor U4463 (N_4463,N_2504,N_2112);
xor U4464 (N_4464,N_2232,N_1956);
and U4465 (N_4465,N_2276,N_2627);
nor U4466 (N_4466,N_1782,N_1987);
and U4467 (N_4467,N_2023,N_2507);
nor U4468 (N_4468,N_1795,N_2311);
or U4469 (N_4469,N_2376,N_1527);
xor U4470 (N_4470,N_1962,N_2310);
and U4471 (N_4471,N_2306,N_2320);
or U4472 (N_4472,N_1575,N_2493);
nor U4473 (N_4473,N_2159,N_1639);
nor U4474 (N_4474,N_1607,N_1591);
and U4475 (N_4475,N_1625,N_2038);
nand U4476 (N_4476,N_2852,N_2472);
nand U4477 (N_4477,N_1983,N_2063);
or U4478 (N_4478,N_1557,N_1864);
nor U4479 (N_4479,N_1593,N_2964);
and U4480 (N_4480,N_1534,N_1654);
or U4481 (N_4481,N_2436,N_1509);
and U4482 (N_4482,N_1997,N_1711);
or U4483 (N_4483,N_1729,N_2087);
nor U4484 (N_4484,N_1524,N_2116);
and U4485 (N_4485,N_2714,N_2975);
nand U4486 (N_4486,N_1616,N_1571);
nand U4487 (N_4487,N_2886,N_1759);
and U4488 (N_4488,N_1900,N_1525);
and U4489 (N_4489,N_1577,N_1732);
xnor U4490 (N_4490,N_2161,N_2750);
or U4491 (N_4491,N_1920,N_1665);
nand U4492 (N_4492,N_2217,N_2410);
and U4493 (N_4493,N_2439,N_2416);
or U4494 (N_4494,N_1520,N_2099);
nor U4495 (N_4495,N_2778,N_2881);
xnor U4496 (N_4496,N_1750,N_2020);
or U4497 (N_4497,N_2368,N_1559);
xnor U4498 (N_4498,N_2196,N_1904);
and U4499 (N_4499,N_2892,N_1775);
nor U4500 (N_4500,N_4318,N_3448);
nor U4501 (N_4501,N_4078,N_4200);
nor U4502 (N_4502,N_3522,N_4455);
or U4503 (N_4503,N_3700,N_4283);
or U4504 (N_4504,N_4257,N_3598);
xor U4505 (N_4505,N_3758,N_3046);
and U4506 (N_4506,N_4055,N_3604);
nor U4507 (N_4507,N_3180,N_3312);
nor U4508 (N_4508,N_4392,N_3354);
and U4509 (N_4509,N_3630,N_4271);
xnor U4510 (N_4510,N_3652,N_3768);
xor U4511 (N_4511,N_3192,N_4029);
nor U4512 (N_4512,N_3791,N_3508);
or U4513 (N_4513,N_4143,N_3589);
or U4514 (N_4514,N_3455,N_4415);
nor U4515 (N_4515,N_4281,N_3644);
nor U4516 (N_4516,N_3707,N_3394);
nand U4517 (N_4517,N_3268,N_3492);
nand U4518 (N_4518,N_4052,N_4256);
xor U4519 (N_4519,N_4491,N_3078);
xnor U4520 (N_4520,N_3682,N_3495);
or U4521 (N_4521,N_3244,N_3490);
and U4522 (N_4522,N_4490,N_3882);
xor U4523 (N_4523,N_4049,N_3562);
or U4524 (N_4524,N_3405,N_3410);
and U4525 (N_4525,N_4195,N_3294);
xor U4526 (N_4526,N_3436,N_3311);
and U4527 (N_4527,N_3272,N_4298);
xnor U4528 (N_4528,N_3478,N_4126);
nor U4529 (N_4529,N_3327,N_4028);
or U4530 (N_4530,N_3142,N_3947);
xor U4531 (N_4531,N_4227,N_4310);
or U4532 (N_4532,N_3989,N_3524);
nand U4533 (N_4533,N_4158,N_3325);
nor U4534 (N_4534,N_3717,N_3109);
nand U4535 (N_4535,N_3107,N_3377);
or U4536 (N_4536,N_4290,N_4097);
xnor U4537 (N_4537,N_3952,N_3494);
nand U4538 (N_4538,N_4347,N_4407);
nor U4539 (N_4539,N_3526,N_3854);
xnor U4540 (N_4540,N_3629,N_4246);
nand U4541 (N_4541,N_3292,N_3452);
nand U4542 (N_4542,N_3211,N_3486);
nand U4543 (N_4543,N_3510,N_4367);
xnor U4544 (N_4544,N_3266,N_4332);
nor U4545 (N_4545,N_3259,N_3550);
xor U4546 (N_4546,N_4149,N_3050);
and U4547 (N_4547,N_3641,N_3970);
nand U4548 (N_4548,N_4082,N_4353);
xnor U4549 (N_4549,N_4448,N_3428);
and U4550 (N_4550,N_3156,N_3541);
nand U4551 (N_4551,N_3442,N_3305);
xor U4552 (N_4552,N_3673,N_3333);
xor U4553 (N_4553,N_3485,N_3565);
nand U4554 (N_4554,N_4285,N_4348);
and U4555 (N_4555,N_3302,N_3561);
xor U4556 (N_4556,N_3875,N_3661);
and U4557 (N_4557,N_3537,N_4156);
and U4558 (N_4558,N_3197,N_3348);
or U4559 (N_4559,N_3191,N_3146);
nand U4560 (N_4560,N_3218,N_4184);
or U4561 (N_4561,N_4008,N_3850);
nand U4562 (N_4562,N_4007,N_3162);
nor U4563 (N_4563,N_3577,N_3179);
xnor U4564 (N_4564,N_4027,N_4245);
or U4565 (N_4565,N_3543,N_4408);
nand U4566 (N_4566,N_3934,N_3602);
nand U4567 (N_4567,N_3297,N_3461);
nor U4568 (N_4568,N_4327,N_3027);
nor U4569 (N_4569,N_3400,N_3463);
or U4570 (N_4570,N_4425,N_4030);
and U4571 (N_4571,N_3987,N_3527);
nor U4572 (N_4572,N_3030,N_4094);
nand U4573 (N_4573,N_3624,N_3320);
or U4574 (N_4574,N_3118,N_3077);
and U4575 (N_4575,N_4215,N_3141);
xnor U4576 (N_4576,N_3065,N_3221);
and U4577 (N_4577,N_3806,N_4228);
nand U4578 (N_4578,N_3099,N_4239);
and U4579 (N_4579,N_3957,N_3429);
xnor U4580 (N_4580,N_4032,N_3597);
xor U4581 (N_4581,N_4344,N_3376);
nor U4582 (N_4582,N_4066,N_3942);
nor U4583 (N_4583,N_3190,N_3496);
xor U4584 (N_4584,N_3096,N_3069);
nor U4585 (N_4585,N_4289,N_3997);
nand U4586 (N_4586,N_3224,N_3977);
and U4587 (N_4587,N_3827,N_3434);
nand U4588 (N_4588,N_3135,N_3532);
and U4589 (N_4589,N_4462,N_3293);
xor U4590 (N_4590,N_4307,N_3631);
nand U4591 (N_4591,N_3176,N_4213);
and U4592 (N_4592,N_3481,N_3688);
and U4593 (N_4593,N_3672,N_4370);
xor U4594 (N_4594,N_4450,N_4087);
and U4595 (N_4595,N_4287,N_3164);
and U4596 (N_4596,N_3219,N_4266);
nand U4597 (N_4597,N_3450,N_3435);
xnor U4598 (N_4598,N_3445,N_4336);
nor U4599 (N_4599,N_3001,N_4105);
xnor U4600 (N_4600,N_3073,N_3122);
nand U4601 (N_4601,N_4489,N_4122);
and U4602 (N_4602,N_4207,N_3782);
nor U4603 (N_4603,N_4333,N_4135);
or U4604 (N_4604,N_3599,N_3385);
nor U4605 (N_4605,N_3796,N_3034);
nand U4606 (N_4606,N_3674,N_3012);
nor U4607 (N_4607,N_3205,N_3169);
and U4608 (N_4608,N_3476,N_3759);
nand U4609 (N_4609,N_3131,N_3343);
xor U4610 (N_4610,N_3919,N_3147);
and U4611 (N_4611,N_3229,N_3780);
or U4612 (N_4612,N_3043,N_4042);
and U4613 (N_4613,N_4026,N_3699);
or U4614 (N_4614,N_3255,N_3430);
nor U4615 (N_4615,N_3324,N_3844);
nor U4616 (N_4616,N_3412,N_3613);
nor U4617 (N_4617,N_3714,N_3225);
xnor U4618 (N_4618,N_4282,N_3881);
nor U4619 (N_4619,N_4437,N_4388);
and U4620 (N_4620,N_4403,N_4361);
and U4621 (N_4621,N_3424,N_3254);
and U4622 (N_4622,N_4124,N_3004);
nor U4623 (N_4623,N_3667,N_3581);
nand U4624 (N_4624,N_4494,N_3896);
or U4625 (N_4625,N_4335,N_3587);
nor U4626 (N_4626,N_3912,N_4334);
or U4627 (N_4627,N_3359,N_3848);
nand U4628 (N_4628,N_3217,N_3372);
nand U4629 (N_4629,N_3468,N_4234);
and U4630 (N_4630,N_3625,N_3095);
or U4631 (N_4631,N_4410,N_4005);
xor U4632 (N_4632,N_3969,N_4064);
xnor U4633 (N_4633,N_3698,N_3584);
or U4634 (N_4634,N_3009,N_3238);
xor U4635 (N_4635,N_4165,N_3940);
xor U4636 (N_4636,N_3763,N_4473);
or U4637 (N_4637,N_4360,N_4365);
nand U4638 (N_4638,N_3016,N_3570);
nor U4639 (N_4639,N_4059,N_3276);
nor U4640 (N_4640,N_3145,N_3057);
and U4641 (N_4641,N_3684,N_3132);
nand U4642 (N_4642,N_3928,N_3222);
nand U4643 (N_4643,N_4401,N_3635);
nor U4644 (N_4644,N_3234,N_3766);
xor U4645 (N_4645,N_4169,N_3816);
xnor U4646 (N_4646,N_3396,N_3418);
or U4647 (N_4647,N_3188,N_3946);
or U4648 (N_4648,N_4436,N_3513);
nand U4649 (N_4649,N_3511,N_3512);
nor U4650 (N_4650,N_4349,N_3863);
nand U4651 (N_4651,N_3499,N_3313);
xnor U4652 (N_4652,N_4373,N_4311);
nor U4653 (N_4653,N_4286,N_3163);
and U4654 (N_4654,N_3299,N_3540);
and U4655 (N_4655,N_3675,N_4208);
or U4656 (N_4656,N_4421,N_3263);
nand U4657 (N_4657,N_3640,N_3756);
nor U4658 (N_4658,N_3264,N_3925);
nor U4659 (N_4659,N_3319,N_3159);
xor U4660 (N_4660,N_3458,N_4134);
nor U4661 (N_4661,N_3045,N_3964);
nor U4662 (N_4662,N_3195,N_3639);
nor U4663 (N_4663,N_4181,N_3194);
or U4664 (N_4664,N_3733,N_4118);
or U4665 (N_4665,N_4383,N_4019);
nor U4666 (N_4666,N_4247,N_3341);
nor U4667 (N_4667,N_4018,N_3828);
nor U4668 (N_4668,N_4154,N_4002);
nor U4669 (N_4669,N_3826,N_4420);
and U4670 (N_4670,N_4251,N_3612);
nor U4671 (N_4671,N_3465,N_3220);
nor U4672 (N_4672,N_3975,N_3172);
nor U4673 (N_4673,N_4446,N_4166);
and U4674 (N_4674,N_3545,N_4268);
nand U4675 (N_4675,N_4080,N_4101);
and U4676 (N_4676,N_4369,N_3460);
and U4677 (N_4677,N_4442,N_3185);
or U4678 (N_4678,N_3008,N_3965);
xor U4679 (N_4679,N_3817,N_4261);
or U4680 (N_4680,N_3849,N_3566);
nand U4681 (N_4681,N_3271,N_3905);
nor U4682 (N_4682,N_3295,N_3535);
xor U4683 (N_4683,N_3923,N_4299);
nor U4684 (N_4684,N_3559,N_4352);
and U4685 (N_4685,N_3867,N_3249);
or U4686 (N_4686,N_4468,N_3678);
and U4687 (N_4687,N_3835,N_4453);
and U4688 (N_4688,N_4481,N_3127);
nand U4689 (N_4689,N_3838,N_3748);
xnor U4690 (N_4690,N_4113,N_3885);
nor U4691 (N_4691,N_3308,N_3974);
nand U4692 (N_4692,N_4021,N_4389);
xor U4693 (N_4693,N_4477,N_4045);
xnor U4694 (N_4694,N_4157,N_3167);
xnor U4695 (N_4695,N_3938,N_3709);
xor U4696 (N_4696,N_4302,N_3807);
nor U4697 (N_4697,N_4241,N_4233);
xor U4698 (N_4698,N_3871,N_3764);
and U4699 (N_4699,N_3544,N_4277);
nand U4700 (N_4700,N_4356,N_4212);
or U4701 (N_4701,N_4293,N_4306);
and U4702 (N_4702,N_4148,N_3967);
nor U4703 (N_4703,N_3151,N_4387);
and U4704 (N_4704,N_3775,N_3280);
xor U4705 (N_4705,N_3315,N_4482);
xor U4706 (N_4706,N_4395,N_4366);
xnor U4707 (N_4707,N_4036,N_4186);
and U4708 (N_4708,N_3591,N_4449);
xnor U4709 (N_4709,N_3466,N_4168);
nor U4710 (N_4710,N_4423,N_3277);
or U4711 (N_4711,N_3039,N_4003);
nor U4712 (N_4712,N_3284,N_3841);
nand U4713 (N_4713,N_4191,N_3323);
nor U4714 (N_4714,N_3471,N_4121);
and U4715 (N_4715,N_3557,N_3393);
xor U4716 (N_4716,N_3388,N_4140);
nor U4717 (N_4717,N_3206,N_3389);
nor U4718 (N_4718,N_3419,N_4465);
nand U4719 (N_4719,N_3011,N_4294);
and U4720 (N_4720,N_3752,N_4153);
xor U4721 (N_4721,N_4398,N_3110);
nor U4722 (N_4722,N_3797,N_3772);
or U4723 (N_4723,N_4432,N_3334);
and U4724 (N_4724,N_3747,N_3979);
nand U4725 (N_4725,N_3770,N_3322);
nand U4726 (N_4726,N_4229,N_4350);
or U4727 (N_4727,N_3335,N_3047);
xor U4728 (N_4728,N_3529,N_3380);
xnor U4729 (N_4729,N_3798,N_4372);
and U4730 (N_4730,N_3178,N_3130);
xor U4731 (N_4731,N_4033,N_3628);
xnor U4732 (N_4732,N_3339,N_3754);
nor U4733 (N_4733,N_4196,N_3618);
or U4734 (N_4734,N_3409,N_3825);
and U4735 (N_4735,N_3262,N_3836);
or U4736 (N_4736,N_3647,N_3993);
nor U4737 (N_4737,N_4136,N_3392);
nand U4738 (N_4738,N_3745,N_3955);
nand U4739 (N_4739,N_3250,N_3983);
or U4740 (N_4740,N_4484,N_3596);
xnor U4741 (N_4741,N_4120,N_3906);
nand U4742 (N_4742,N_3711,N_4230);
xor U4743 (N_4743,N_3068,N_3852);
nor U4744 (N_4744,N_3901,N_4272);
nor U4745 (N_4745,N_3856,N_3382);
xor U4746 (N_4746,N_4204,N_3801);
or U4747 (N_4747,N_3858,N_3677);
or U4748 (N_4748,N_3013,N_3310);
nor U4749 (N_4749,N_3075,N_4061);
xnor U4750 (N_4750,N_3866,N_4071);
and U4751 (N_4751,N_4024,N_3546);
xnor U4752 (N_4752,N_3232,N_4378);
or U4753 (N_4753,N_4109,N_4434);
or U4754 (N_4754,N_3171,N_4456);
and U4755 (N_4755,N_3988,N_3365);
xnor U4756 (N_4756,N_4133,N_3799);
nand U4757 (N_4757,N_3257,N_3051);
xnor U4758 (N_4758,N_4131,N_3100);
nor U4759 (N_4759,N_4471,N_3088);
xnor U4760 (N_4760,N_4428,N_3976);
nor U4761 (N_4761,N_4412,N_3152);
nor U4762 (N_4762,N_3744,N_3133);
nand U4763 (N_4763,N_4072,N_3692);
xor U4764 (N_4764,N_3336,N_3715);
or U4765 (N_4765,N_3571,N_3098);
or U4766 (N_4766,N_4235,N_3873);
nand U4767 (N_4767,N_3981,N_3862);
and U4768 (N_4768,N_4377,N_4390);
nand U4769 (N_4769,N_4357,N_3153);
nor U4770 (N_4770,N_3531,N_3658);
nand U4771 (N_4771,N_4117,N_3681);
and U4772 (N_4772,N_4062,N_3776);
nand U4773 (N_4773,N_3921,N_3116);
xnor U4774 (N_4774,N_3144,N_4433);
or U4775 (N_4775,N_3421,N_4180);
nand U4776 (N_4776,N_3615,N_4321);
or U4777 (N_4777,N_3017,N_4265);
and U4778 (N_4778,N_3632,N_4253);
xor U4779 (N_4779,N_3793,N_3374);
and U4780 (N_4780,N_4457,N_3564);
nor U4781 (N_4781,N_4031,N_3114);
and U4782 (N_4782,N_3353,N_4254);
nor U4783 (N_4783,N_4313,N_4380);
or U4784 (N_4784,N_3583,N_3340);
or U4785 (N_4785,N_3137,N_4331);
nor U4786 (N_4786,N_3578,N_3815);
and U4787 (N_4787,N_3554,N_3306);
or U4788 (N_4788,N_3833,N_4221);
or U4789 (N_4789,N_3911,N_4106);
xnor U4790 (N_4790,N_3203,N_3845);
nand U4791 (N_4791,N_3083,N_3304);
nor U4792 (N_4792,N_3651,N_3035);
xnor U4793 (N_4793,N_3755,N_3586);
nand U4794 (N_4794,N_3683,N_3290);
or U4795 (N_4795,N_4260,N_4142);
nand U4796 (N_4796,N_3992,N_3722);
or U4797 (N_4797,N_3187,N_3884);
nor U4798 (N_4798,N_3309,N_3636);
nand U4799 (N_4799,N_3737,N_3746);
nor U4800 (N_4800,N_3732,N_3433);
or U4801 (N_4801,N_3182,N_3175);
xor U4802 (N_4802,N_4201,N_3018);
nor U4803 (N_4803,N_3665,N_3379);
xor U4804 (N_4804,N_3605,N_3660);
nor U4805 (N_4805,N_3804,N_3237);
or U4806 (N_4806,N_3278,N_4190);
xor U4807 (N_4807,N_3106,N_4044);
or U4808 (N_4808,N_3761,N_4279);
and U4809 (N_4809,N_3019,N_4319);
nor U4810 (N_4810,N_4466,N_4047);
nand U4811 (N_4811,N_3910,N_3252);
nor U4812 (N_4812,N_3959,N_3378);
nand U4813 (N_4813,N_4079,N_4362);
or U4814 (N_4814,N_3814,N_3242);
and U4815 (N_4815,N_4292,N_3381);
nand U4816 (N_4816,N_3781,N_3346);
and U4817 (N_4817,N_3369,N_3580);
nor U4818 (N_4818,N_4363,N_3139);
or U4819 (N_4819,N_3129,N_3403);
and U4820 (N_4820,N_4155,N_3456);
xnor U4821 (N_4821,N_4038,N_3534);
and U4822 (N_4822,N_3489,N_4385);
and U4823 (N_4823,N_3402,N_3549);
xor U4824 (N_4824,N_3861,N_4162);
nor U4825 (N_4825,N_3506,N_3444);
xor U4826 (N_4826,N_4478,N_3656);
and U4827 (N_4827,N_3935,N_3742);
nor U4828 (N_4828,N_3502,N_3670);
xor U4829 (N_4829,N_4351,N_3820);
nor U4830 (N_4830,N_4431,N_3834);
and U4831 (N_4831,N_3480,N_3767);
and U4832 (N_4832,N_4023,N_3783);
nor U4833 (N_4833,N_4053,N_4391);
xnor U4834 (N_4834,N_4000,N_4070);
nand U4835 (N_4835,N_4375,N_3880);
or U4836 (N_4836,N_3398,N_3859);
nand U4837 (N_4837,N_4161,N_4404);
or U4838 (N_4838,N_4288,N_3966);
nor U4839 (N_4839,N_4259,N_3572);
xnor U4840 (N_4840,N_4009,N_3680);
or U4841 (N_4841,N_4050,N_3044);
or U4842 (N_4842,N_3842,N_4341);
xor U4843 (N_4843,N_4130,N_3113);
nor U4844 (N_4844,N_3857,N_3364);
nand U4845 (N_4845,N_3939,N_4339);
and U4846 (N_4846,N_4382,N_4056);
nor U4847 (N_4847,N_3041,N_3762);
nand U4848 (N_4848,N_3633,N_3666);
nand U4849 (N_4849,N_3671,N_3962);
or U4850 (N_4850,N_3922,N_4240);
nand U4851 (N_4851,N_3467,N_4326);
and U4852 (N_4852,N_4496,N_3990);
xor U4853 (N_4853,N_3548,N_3607);
and U4854 (N_4854,N_4474,N_4076);
or U4855 (N_4855,N_4427,N_4296);
xor U4856 (N_4856,N_4090,N_3240);
xor U4857 (N_4857,N_3415,N_3738);
xnor U4858 (N_4858,N_3813,N_4107);
or U4859 (N_4859,N_3091,N_3081);
xnor U4860 (N_4860,N_4400,N_4188);
and U4861 (N_4861,N_4419,N_3235);
nand U4862 (N_4862,N_3691,N_4262);
nand U4863 (N_4863,N_4416,N_3005);
xnor U4864 (N_4864,N_3089,N_4499);
xnor U4865 (N_4865,N_3594,N_3283);
or U4866 (N_4866,N_4252,N_3941);
xor U4867 (N_4867,N_3757,N_3387);
xor U4868 (N_4868,N_3637,N_3654);
or U4869 (N_4869,N_3148,N_4051);
xor U4870 (N_4870,N_3918,N_4010);
or U4871 (N_4871,N_3477,N_3840);
nand U4872 (N_4872,N_3702,N_3360);
nand U4873 (N_4873,N_3634,N_4202);
or U4874 (N_4874,N_4170,N_4138);
nor U4875 (N_4875,N_4402,N_3803);
nor U4876 (N_4876,N_4236,N_3904);
nor U4877 (N_4877,N_3097,N_3422);
and U4878 (N_4878,N_4376,N_3573);
xnor U4879 (N_4879,N_3556,N_3251);
or U4880 (N_4880,N_4443,N_4152);
or U4881 (N_4881,N_3503,N_3080);
nor U4882 (N_4882,N_3473,N_3662);
or U4883 (N_4883,N_3610,N_3507);
and U4884 (N_4884,N_3337,N_3208);
xor U4885 (N_4885,N_3120,N_4183);
xnor U4886 (N_4886,N_4399,N_4337);
xnor U4887 (N_4887,N_3860,N_3869);
or U4888 (N_4888,N_3887,N_4128);
and U4889 (N_4889,N_3567,N_3879);
nand U4890 (N_4890,N_3972,N_4238);
nand U4891 (N_4891,N_3831,N_3248);
nor U4892 (N_4892,N_3085,N_4086);
nor U4893 (N_4893,N_3425,N_3427);
or U4894 (N_4894,N_4173,N_3855);
xor U4895 (N_4895,N_3223,N_4264);
nand U4896 (N_4896,N_3706,N_3014);
and U4897 (N_4897,N_3846,N_4480);
nand U4898 (N_4898,N_3128,N_3464);
xnor U4899 (N_4899,N_3563,N_3181);
and U4900 (N_4900,N_3138,N_3676);
and U4901 (N_4901,N_4393,N_3112);
and U4902 (N_4902,N_4020,N_4025);
nand U4903 (N_4903,N_3287,N_3288);
nand U4904 (N_4904,N_3719,N_3937);
nor U4905 (N_4905,N_3411,N_4275);
and U4906 (N_4906,N_3273,N_4438);
and U4907 (N_4907,N_3498,N_3518);
xnor U4908 (N_4908,N_3207,N_3201);
and U4909 (N_4909,N_3161,N_4119);
nand U4910 (N_4910,N_3479,N_3600);
nand U4911 (N_4911,N_3054,N_3995);
nand U4912 (N_4912,N_4151,N_4100);
xnor U4913 (N_4913,N_3200,N_3713);
nand U4914 (N_4914,N_4248,N_3291);
nor U4915 (N_4915,N_4185,N_3822);
nor U4916 (N_4916,N_3279,N_3832);
and U4917 (N_4917,N_3101,N_3617);
and U4918 (N_4918,N_3328,N_3611);
nand U4919 (N_4919,N_3483,N_3712);
and U4920 (N_4920,N_3202,N_4217);
or U4921 (N_4921,N_3943,N_3285);
and U4922 (N_4922,N_3547,N_3892);
xor U4923 (N_4923,N_3620,N_3214);
nand U4924 (N_4924,N_3727,N_3493);
or U4925 (N_4925,N_3542,N_4315);
or U4926 (N_4926,N_4014,N_3007);
or U4927 (N_4927,N_4301,N_3576);
nand U4928 (N_4928,N_4074,N_3784);
nor U4929 (N_4929,N_3991,N_3451);
xnor U4930 (N_4930,N_4314,N_4013);
nor U4931 (N_4931,N_3420,N_4461);
nand U4932 (N_4932,N_3999,N_4127);
xnor U4933 (N_4933,N_4067,N_4269);
nand U4934 (N_4934,N_3245,N_4258);
nand U4935 (N_4935,N_3270,N_3318);
xnor U4936 (N_4936,N_3794,N_4325);
and U4937 (N_4937,N_3504,N_3914);
or U4938 (N_4938,N_3036,N_3800);
and U4939 (N_4939,N_4479,N_4330);
xor U4940 (N_4940,N_3903,N_3150);
and U4941 (N_4941,N_3391,N_3643);
and U4942 (N_4942,N_3094,N_3160);
xor U4943 (N_4943,N_3040,N_4340);
and U4944 (N_4944,N_3802,N_3345);
or U4945 (N_4945,N_3984,N_3760);
nand U4946 (N_4946,N_4096,N_4475);
xor U4947 (N_4947,N_4469,N_4214);
nor U4948 (N_4948,N_3210,N_3978);
or U4949 (N_4949,N_3743,N_3177);
and U4950 (N_4950,N_4276,N_3482);
or U4951 (N_4951,N_3718,N_4034);
or U4952 (N_4952,N_4171,N_3771);
and U4953 (N_4953,N_4129,N_4312);
nor U4954 (N_4954,N_3853,N_3487);
nor U4955 (N_4955,N_4329,N_3355);
nor U4956 (N_4956,N_4406,N_3053);
and U4957 (N_4957,N_3298,N_3031);
xnor U4958 (N_4958,N_3447,N_3316);
nand U4959 (N_4959,N_4394,N_3694);
nor U4960 (N_4960,N_3553,N_3948);
xor U4961 (N_4961,N_3063,N_4384);
xnor U4962 (N_4962,N_3693,N_3659);
nor U4963 (N_4963,N_3183,N_3818);
or U4964 (N_4964,N_4304,N_3552);
or U4965 (N_4965,N_4374,N_4041);
or U4966 (N_4966,N_4150,N_4163);
nor U4967 (N_4967,N_4065,N_3663);
nor U4968 (N_4968,N_4274,N_3533);
or U4969 (N_4969,N_3728,N_4464);
nand U4970 (N_4970,N_3621,N_3716);
or U4971 (N_4971,N_4343,N_3648);
nand U4972 (N_4972,N_3087,N_3689);
and U4973 (N_4973,N_4194,N_3741);
or U4974 (N_4974,N_3616,N_3908);
xor U4975 (N_4975,N_3119,N_3125);
nor U4976 (N_4976,N_4141,N_3404);
nand U4977 (N_4977,N_4498,N_3890);
nor U4978 (N_4978,N_3363,N_3189);
nand U4979 (N_4979,N_3623,N_3705);
or U4980 (N_4980,N_3358,N_3084);
xor U4981 (N_4981,N_3307,N_3500);
and U4982 (N_4982,N_3126,N_4177);
or U4983 (N_4983,N_4016,N_3514);
and U4984 (N_4984,N_3423,N_3876);
or U4985 (N_4985,N_3929,N_3601);
xnor U4986 (N_4986,N_4172,N_3449);
nand U4987 (N_4987,N_3893,N_3029);
nand U4988 (N_4988,N_4418,N_3439);
and U4989 (N_4989,N_4405,N_4081);
and U4990 (N_4990,N_3123,N_3703);
nor U4991 (N_4991,N_4458,N_3950);
nand U4992 (N_4992,N_3157,N_3143);
and U4993 (N_4993,N_3399,N_4411);
nor U4994 (N_4994,N_4077,N_3216);
xnor U4995 (N_4995,N_4112,N_3710);
xnor U4996 (N_4996,N_3174,N_3314);
and U4997 (N_4997,N_3949,N_3645);
xnor U4998 (N_4998,N_3082,N_3275);
nand U4999 (N_4999,N_3592,N_3021);
nand U5000 (N_5000,N_4263,N_4409);
nor U5001 (N_5001,N_3895,N_3198);
xor U5002 (N_5002,N_3370,N_3383);
or U5003 (N_5003,N_4358,N_3154);
xnor U5004 (N_5004,N_3265,N_3723);
xnor U5005 (N_5005,N_3555,N_3551);
and U5006 (N_5006,N_3258,N_4328);
and U5007 (N_5007,N_3437,N_4278);
and U5008 (N_5008,N_3406,N_4223);
and U5009 (N_5009,N_4192,N_4085);
nor U5010 (N_5010,N_3296,N_3236);
and U5011 (N_5011,N_3475,N_3347);
nor U5012 (N_5012,N_3792,N_3331);
xnor U5013 (N_5013,N_4459,N_3932);
nor U5014 (N_5014,N_4379,N_3212);
and U5015 (N_5015,N_3401,N_3668);
nand U5016 (N_5016,N_3704,N_3915);
or U5017 (N_5017,N_3664,N_3246);
and U5018 (N_5018,N_3256,N_3769);
or U5019 (N_5019,N_4476,N_3985);
nand U5020 (N_5020,N_3971,N_4322);
and U5021 (N_5021,N_4209,N_3536);
nor U5022 (N_5022,N_4338,N_3686);
or U5023 (N_5023,N_4486,N_3158);
xnor U5024 (N_5024,N_3134,N_3963);
nand U5025 (N_5025,N_4291,N_4284);
or U5026 (N_5026,N_4123,N_3375);
xnor U5027 (N_5027,N_4309,N_4199);
nand U5028 (N_5028,N_3520,N_3994);
or U5029 (N_5029,N_3821,N_3173);
nand U5030 (N_5030,N_4102,N_3982);
and U5031 (N_5031,N_3996,N_3779);
nand U5032 (N_5032,N_3326,N_3239);
and U5033 (N_5033,N_3459,N_3777);
nor U5034 (N_5034,N_4203,N_3883);
or U5035 (N_5035,N_4004,N_3539);
nand U5036 (N_5036,N_3260,N_4280);
or U5037 (N_5037,N_4139,N_4493);
or U5038 (N_5038,N_3973,N_3350);
nor U5039 (N_5039,N_4303,N_4060);
nor U5040 (N_5040,N_3627,N_4430);
and U5041 (N_5041,N_3386,N_3209);
and U5042 (N_5042,N_4058,N_4182);
nor U5043 (N_5043,N_4110,N_3575);
and U5044 (N_5044,N_3300,N_4093);
and U5045 (N_5045,N_3805,N_4206);
xnor U5046 (N_5046,N_3199,N_3945);
nor U5047 (N_5047,N_3614,N_3000);
or U5048 (N_5048,N_3843,N_3361);
or U5049 (N_5049,N_4222,N_3124);
and U5050 (N_5050,N_3917,N_4483);
xnor U5051 (N_5051,N_4006,N_3371);
and U5052 (N_5052,N_4472,N_3140);
or U5053 (N_5053,N_4037,N_3149);
nor U5054 (N_5054,N_4220,N_4011);
and U5055 (N_5055,N_3669,N_3810);
nor U5056 (N_5056,N_4355,N_3070);
or U5057 (N_5057,N_3497,N_3491);
and U5058 (N_5058,N_4320,N_3585);
and U5059 (N_5059,N_3790,N_3488);
nand U5060 (N_5060,N_4224,N_3695);
nor U5061 (N_5061,N_4323,N_4063);
nand U5062 (N_5062,N_4174,N_3899);
nand U5063 (N_5063,N_3438,N_4445);
xor U5064 (N_5064,N_4164,N_3090);
and U5065 (N_5065,N_4297,N_3368);
or U5066 (N_5066,N_4083,N_3015);
and U5067 (N_5067,N_3342,N_3453);
or U5068 (N_5068,N_3568,N_4175);
nor U5069 (N_5069,N_3384,N_4422);
xor U5070 (N_5070,N_3117,N_4167);
or U5071 (N_5071,N_3373,N_3525);
xnor U5072 (N_5072,N_3788,N_3753);
xnor U5073 (N_5073,N_3517,N_3227);
nand U5074 (N_5074,N_3735,N_4043);
xor U5075 (N_5075,N_4159,N_3724);
and U5076 (N_5076,N_3062,N_3523);
nand U5077 (N_5077,N_4435,N_4046);
nor U5078 (N_5078,N_4178,N_3267);
and U5079 (N_5079,N_3609,N_3913);
xor U5080 (N_5080,N_3872,N_3907);
nor U5081 (N_5081,N_3739,N_4295);
xor U5082 (N_5082,N_3344,N_3367);
xor U5083 (N_5083,N_3936,N_3115);
nor U5084 (N_5084,N_3329,N_4069);
and U5085 (N_5085,N_3058,N_4242);
nor U5086 (N_5086,N_3301,N_4452);
or U5087 (N_5087,N_3795,N_3352);
or U5088 (N_5088,N_3956,N_4232);
nor U5089 (N_5089,N_3002,N_3193);
nand U5090 (N_5090,N_3072,N_3730);
nand U5091 (N_5091,N_3916,N_4470);
and U5092 (N_5092,N_4099,N_4424);
nor U5093 (N_5093,N_3213,N_4488);
nor U5094 (N_5094,N_4015,N_4371);
and U5095 (N_5095,N_3944,N_4179);
or U5096 (N_5096,N_4439,N_3093);
and U5097 (N_5097,N_4022,N_3897);
nand U5098 (N_5098,N_4137,N_3593);
or U5099 (N_5099,N_4231,N_3060);
nor U5100 (N_5100,N_3685,N_3274);
nand U5101 (N_5101,N_4487,N_3516);
and U5102 (N_5102,N_3049,N_3519);
xor U5103 (N_5103,N_4210,N_4346);
nor U5104 (N_5104,N_3408,N_3281);
and U5105 (N_5105,N_3066,N_3356);
or U5106 (N_5106,N_4273,N_3909);
nand U5107 (N_5107,N_4160,N_3032);
and U5108 (N_5108,N_3509,N_3441);
nand U5109 (N_5109,N_3823,N_3186);
and U5110 (N_5110,N_3170,N_3655);
or U5111 (N_5111,N_3056,N_3864);
xnor U5112 (N_5112,N_4255,N_4414);
xor U5113 (N_5113,N_4441,N_3111);
xnor U5114 (N_5114,N_3968,N_3679);
xor U5115 (N_5115,N_4485,N_4115);
nor U5116 (N_5116,N_4211,N_4111);
and U5117 (N_5117,N_3765,N_3261);
or U5118 (N_5118,N_3958,N_3390);
xor U5119 (N_5119,N_4463,N_3734);
nand U5120 (N_5120,N_4057,N_3282);
xnor U5121 (N_5121,N_3076,N_3588);
and U5122 (N_5122,N_3010,N_3332);
xor U5123 (N_5123,N_3022,N_4017);
and U5124 (N_5124,N_4187,N_3808);
or U5125 (N_5125,N_3638,N_3560);
or U5126 (N_5126,N_4091,N_3064);
or U5127 (N_5127,N_4075,N_4413);
and U5128 (N_5128,N_3657,N_3426);
nor U5129 (N_5129,N_4237,N_4001);
nand U5130 (N_5130,N_3886,N_3824);
xor U5131 (N_5131,N_3569,N_3690);
xor U5132 (N_5132,N_3105,N_3839);
nor U5133 (N_5133,N_3931,N_3530);
xnor U5134 (N_5134,N_3233,N_3052);
or U5135 (N_5135,N_3961,N_3474);
nand U5136 (N_5136,N_3902,N_4354);
and U5137 (N_5137,N_3431,N_3619);
and U5138 (N_5138,N_3443,N_4054);
nand U5139 (N_5139,N_3025,N_3457);
and U5140 (N_5140,N_3231,N_3595);
and U5141 (N_5141,N_3868,N_3321);
and U5142 (N_5142,N_4205,N_3121);
nand U5143 (N_5143,N_3184,N_4098);
xnor U5144 (N_5144,N_3042,N_4364);
and U5145 (N_5145,N_4219,N_3061);
or U5146 (N_5146,N_3933,N_4249);
and U5147 (N_5147,N_3608,N_3888);
xor U5148 (N_5148,N_3558,N_3020);
nand U5149 (N_5149,N_4084,N_4397);
nor U5150 (N_5150,N_3472,N_3751);
or U5151 (N_5151,N_3582,N_4417);
and U5152 (N_5152,N_3454,N_3247);
and U5153 (N_5153,N_3785,N_4495);
and U5154 (N_5154,N_3515,N_4048);
and U5155 (N_5155,N_4116,N_4359);
and U5156 (N_5156,N_3006,N_4342);
nand U5157 (N_5157,N_3074,N_4088);
and U5158 (N_5158,N_4381,N_3646);
nor U5159 (N_5159,N_4270,N_3366);
or U5160 (N_5160,N_3878,N_3720);
xnor U5161 (N_5161,N_3847,N_3196);
nor U5162 (N_5162,N_3462,N_3926);
nor U5163 (N_5163,N_3697,N_4012);
or U5164 (N_5164,N_3407,N_3230);
nand U5165 (N_5165,N_4092,N_3877);
or U5166 (N_5166,N_4308,N_3155);
nand U5167 (N_5167,N_3528,N_3446);
or U5168 (N_5168,N_4176,N_4189);
nand U5169 (N_5169,N_4108,N_3998);
and U5170 (N_5170,N_3484,N_3898);
xnor U5171 (N_5171,N_3642,N_4317);
and U5172 (N_5172,N_3851,N_4426);
or U5173 (N_5173,N_3432,N_3108);
xnor U5174 (N_5174,N_3136,N_3330);
nand U5175 (N_5175,N_3048,N_3696);
nor U5176 (N_5176,N_4243,N_4440);
nor U5177 (N_5177,N_4250,N_3574);
nor U5178 (N_5178,N_3215,N_3870);
or U5179 (N_5179,N_3924,N_3440);
nor U5180 (N_5180,N_3003,N_3395);
xor U5181 (N_5181,N_3086,N_3059);
nand U5182 (N_5182,N_3317,N_4035);
nand U5183 (N_5183,N_3079,N_3749);
and U5184 (N_5184,N_3773,N_4460);
and U5185 (N_5185,N_4068,N_4103);
nand U5186 (N_5186,N_3338,N_3874);
nor U5187 (N_5187,N_3243,N_4226);
nand U5188 (N_5188,N_3960,N_3253);
xor U5189 (N_5189,N_3092,N_3024);
and U5190 (N_5190,N_4429,N_4396);
or U5191 (N_5191,N_3357,N_3067);
or U5192 (N_5192,N_3812,N_4492);
xor U5193 (N_5193,N_4324,N_3033);
or U5194 (N_5194,N_3303,N_4144);
nor U5195 (N_5195,N_3953,N_3351);
nor U5196 (N_5196,N_3104,N_3789);
nand U5197 (N_5197,N_3725,N_3416);
xnor U5198 (N_5198,N_3102,N_3649);
and U5199 (N_5199,N_4216,N_4451);
xnor U5200 (N_5200,N_3920,N_4040);
nor U5201 (N_5201,N_3269,N_3731);
nand U5202 (N_5202,N_3986,N_3590);
nor U5203 (N_5203,N_3837,N_3778);
and U5204 (N_5204,N_4368,N_4146);
nor U5205 (N_5205,N_3786,N_3606);
or U5206 (N_5206,N_4316,N_3740);
nor U5207 (N_5207,N_3362,N_3286);
and U5208 (N_5208,N_3037,N_3166);
nand U5209 (N_5209,N_3469,N_3026);
xor U5210 (N_5210,N_3819,N_3787);
or U5211 (N_5211,N_3900,N_4497);
and U5212 (N_5212,N_4095,N_3071);
nand U5213 (N_5213,N_3501,N_3865);
nand U5214 (N_5214,N_3204,N_4305);
or U5215 (N_5215,N_3397,N_4132);
xnor U5216 (N_5216,N_3028,N_3023);
xor U5217 (N_5217,N_3289,N_3729);
and U5218 (N_5218,N_3811,N_3521);
xor U5219 (N_5219,N_4089,N_3168);
or U5220 (N_5220,N_4125,N_3538);
nand U5221 (N_5221,N_4218,N_3750);
or U5222 (N_5222,N_3980,N_4198);
xnor U5223 (N_5223,N_3038,N_3626);
nand U5224 (N_5224,N_3927,N_3951);
nor U5225 (N_5225,N_4104,N_4197);
nor U5226 (N_5226,N_3470,N_3726);
or U5227 (N_5227,N_3505,N_3650);
or U5228 (N_5228,N_3413,N_4114);
nor U5229 (N_5229,N_3103,N_4073);
nor U5230 (N_5230,N_4444,N_4244);
xor U5231 (N_5231,N_4145,N_3721);
xor U5232 (N_5232,N_4345,N_3809);
or U5233 (N_5233,N_3687,N_4147);
xnor U5234 (N_5234,N_3774,N_4225);
nor U5235 (N_5235,N_3954,N_4267);
nand U5236 (N_5236,N_4300,N_3830);
nor U5237 (N_5237,N_3417,N_3701);
xnor U5238 (N_5238,N_4467,N_3891);
and U5239 (N_5239,N_3349,N_3226);
xor U5240 (N_5240,N_3708,N_4039);
and U5241 (N_5241,N_3165,N_4454);
nor U5242 (N_5242,N_3622,N_3889);
xnor U5243 (N_5243,N_3930,N_4386);
nor U5244 (N_5244,N_3603,N_3579);
or U5245 (N_5245,N_3228,N_3829);
or U5246 (N_5246,N_3414,N_4193);
and U5247 (N_5247,N_4447,N_3055);
and U5248 (N_5248,N_3241,N_3736);
nand U5249 (N_5249,N_3653,N_3894);
and U5250 (N_5250,N_4298,N_4106);
nor U5251 (N_5251,N_4203,N_3562);
nand U5252 (N_5252,N_3089,N_3827);
nand U5253 (N_5253,N_3795,N_3686);
nand U5254 (N_5254,N_3754,N_3260);
nand U5255 (N_5255,N_3238,N_4404);
or U5256 (N_5256,N_4271,N_3863);
and U5257 (N_5257,N_3537,N_3433);
and U5258 (N_5258,N_4352,N_4284);
or U5259 (N_5259,N_4144,N_3352);
or U5260 (N_5260,N_3644,N_3830);
nand U5261 (N_5261,N_3290,N_3693);
nor U5262 (N_5262,N_3600,N_3005);
nor U5263 (N_5263,N_3498,N_4144);
or U5264 (N_5264,N_3760,N_4201);
nor U5265 (N_5265,N_4280,N_4403);
and U5266 (N_5266,N_4050,N_4091);
xor U5267 (N_5267,N_3406,N_3023);
and U5268 (N_5268,N_4379,N_3003);
nand U5269 (N_5269,N_3084,N_4346);
nand U5270 (N_5270,N_3622,N_3953);
nand U5271 (N_5271,N_4099,N_4059);
nand U5272 (N_5272,N_4419,N_4471);
xor U5273 (N_5273,N_3410,N_3781);
or U5274 (N_5274,N_4036,N_3497);
nor U5275 (N_5275,N_3842,N_3414);
and U5276 (N_5276,N_4100,N_3849);
nor U5277 (N_5277,N_4337,N_4446);
nand U5278 (N_5278,N_3760,N_3828);
xor U5279 (N_5279,N_3491,N_4368);
nand U5280 (N_5280,N_3648,N_4216);
nor U5281 (N_5281,N_3833,N_3660);
nor U5282 (N_5282,N_3625,N_3290);
nand U5283 (N_5283,N_3935,N_4353);
nand U5284 (N_5284,N_3732,N_3529);
nor U5285 (N_5285,N_3828,N_4418);
xnor U5286 (N_5286,N_3010,N_3060);
or U5287 (N_5287,N_3374,N_3347);
nor U5288 (N_5288,N_3264,N_3350);
xnor U5289 (N_5289,N_3563,N_3505);
and U5290 (N_5290,N_3755,N_3389);
and U5291 (N_5291,N_3205,N_3931);
xor U5292 (N_5292,N_3884,N_4415);
or U5293 (N_5293,N_4201,N_3240);
or U5294 (N_5294,N_3743,N_4103);
and U5295 (N_5295,N_3858,N_3605);
and U5296 (N_5296,N_4084,N_3210);
xor U5297 (N_5297,N_4018,N_4030);
xor U5298 (N_5298,N_3529,N_3118);
nand U5299 (N_5299,N_3992,N_3660);
or U5300 (N_5300,N_3227,N_3172);
and U5301 (N_5301,N_3198,N_3174);
and U5302 (N_5302,N_3660,N_4144);
xor U5303 (N_5303,N_3325,N_4305);
xnor U5304 (N_5304,N_3754,N_4193);
xnor U5305 (N_5305,N_3117,N_3980);
nor U5306 (N_5306,N_3877,N_4408);
and U5307 (N_5307,N_3009,N_4446);
nor U5308 (N_5308,N_4218,N_3225);
nor U5309 (N_5309,N_3427,N_3836);
nor U5310 (N_5310,N_3292,N_4261);
or U5311 (N_5311,N_3875,N_3331);
nand U5312 (N_5312,N_3860,N_3012);
and U5313 (N_5313,N_3465,N_4171);
nand U5314 (N_5314,N_3649,N_3037);
and U5315 (N_5315,N_3198,N_3456);
nor U5316 (N_5316,N_3969,N_3871);
xor U5317 (N_5317,N_4268,N_4474);
nor U5318 (N_5318,N_4041,N_4476);
nand U5319 (N_5319,N_3202,N_4256);
or U5320 (N_5320,N_4495,N_3782);
or U5321 (N_5321,N_4117,N_3184);
and U5322 (N_5322,N_3554,N_3065);
nand U5323 (N_5323,N_3052,N_3392);
nand U5324 (N_5324,N_3067,N_4294);
or U5325 (N_5325,N_3480,N_3157);
or U5326 (N_5326,N_3567,N_4445);
nor U5327 (N_5327,N_3675,N_3938);
nor U5328 (N_5328,N_3664,N_4171);
nand U5329 (N_5329,N_3960,N_4430);
nor U5330 (N_5330,N_3598,N_3596);
nor U5331 (N_5331,N_4257,N_3776);
nand U5332 (N_5332,N_3282,N_3220);
xnor U5333 (N_5333,N_3411,N_4052);
xor U5334 (N_5334,N_3026,N_4124);
nor U5335 (N_5335,N_4369,N_3110);
or U5336 (N_5336,N_4106,N_3198);
nor U5337 (N_5337,N_3975,N_3592);
nor U5338 (N_5338,N_3632,N_3177);
and U5339 (N_5339,N_3036,N_3308);
nor U5340 (N_5340,N_4089,N_3300);
nand U5341 (N_5341,N_4043,N_3706);
xor U5342 (N_5342,N_3106,N_3292);
or U5343 (N_5343,N_3811,N_3444);
nor U5344 (N_5344,N_3868,N_4163);
xnor U5345 (N_5345,N_3096,N_4496);
or U5346 (N_5346,N_3564,N_4247);
nand U5347 (N_5347,N_4260,N_3391);
and U5348 (N_5348,N_3732,N_3916);
and U5349 (N_5349,N_3328,N_3716);
xor U5350 (N_5350,N_3438,N_4226);
xnor U5351 (N_5351,N_3173,N_4387);
or U5352 (N_5352,N_3004,N_4392);
nand U5353 (N_5353,N_3244,N_3251);
and U5354 (N_5354,N_3857,N_4381);
and U5355 (N_5355,N_3521,N_4217);
or U5356 (N_5356,N_4092,N_4390);
and U5357 (N_5357,N_3769,N_3371);
and U5358 (N_5358,N_4362,N_3431);
nor U5359 (N_5359,N_3079,N_3017);
xnor U5360 (N_5360,N_3799,N_4157);
nor U5361 (N_5361,N_3274,N_4355);
nand U5362 (N_5362,N_3909,N_3040);
nor U5363 (N_5363,N_3443,N_4166);
and U5364 (N_5364,N_4373,N_4429);
or U5365 (N_5365,N_3592,N_4082);
and U5366 (N_5366,N_3276,N_3688);
nand U5367 (N_5367,N_3828,N_3355);
and U5368 (N_5368,N_4428,N_3743);
nand U5369 (N_5369,N_3075,N_3087);
or U5370 (N_5370,N_3177,N_3017);
and U5371 (N_5371,N_4196,N_3762);
nand U5372 (N_5372,N_4355,N_4378);
nor U5373 (N_5373,N_3759,N_3619);
nand U5374 (N_5374,N_3063,N_4216);
and U5375 (N_5375,N_3257,N_3206);
nor U5376 (N_5376,N_3552,N_3535);
nor U5377 (N_5377,N_3324,N_3358);
nor U5378 (N_5378,N_3160,N_3091);
xor U5379 (N_5379,N_4429,N_3111);
xor U5380 (N_5380,N_3638,N_3156);
or U5381 (N_5381,N_3070,N_3361);
and U5382 (N_5382,N_3624,N_3412);
or U5383 (N_5383,N_3385,N_4030);
and U5384 (N_5384,N_3943,N_3556);
or U5385 (N_5385,N_4122,N_3412);
nand U5386 (N_5386,N_3450,N_3475);
xnor U5387 (N_5387,N_4304,N_3410);
xor U5388 (N_5388,N_3018,N_4199);
nand U5389 (N_5389,N_3606,N_3792);
and U5390 (N_5390,N_3834,N_3822);
nand U5391 (N_5391,N_3697,N_3726);
and U5392 (N_5392,N_3530,N_4414);
nand U5393 (N_5393,N_4496,N_4386);
or U5394 (N_5394,N_4427,N_4207);
nor U5395 (N_5395,N_4292,N_3203);
and U5396 (N_5396,N_3675,N_3702);
xnor U5397 (N_5397,N_3291,N_4373);
or U5398 (N_5398,N_3070,N_4336);
xor U5399 (N_5399,N_3517,N_4281);
and U5400 (N_5400,N_3413,N_3124);
nand U5401 (N_5401,N_3184,N_3361);
nand U5402 (N_5402,N_4447,N_3442);
nand U5403 (N_5403,N_3569,N_3911);
nand U5404 (N_5404,N_3260,N_3968);
nand U5405 (N_5405,N_3486,N_3738);
and U5406 (N_5406,N_3333,N_3796);
nor U5407 (N_5407,N_3708,N_4483);
xnor U5408 (N_5408,N_4035,N_3577);
nor U5409 (N_5409,N_3652,N_3589);
nand U5410 (N_5410,N_4247,N_4322);
xnor U5411 (N_5411,N_4409,N_3029);
and U5412 (N_5412,N_3192,N_4289);
xnor U5413 (N_5413,N_3023,N_3314);
or U5414 (N_5414,N_4261,N_3340);
xor U5415 (N_5415,N_3460,N_3036);
nand U5416 (N_5416,N_3557,N_4318);
nand U5417 (N_5417,N_3572,N_3874);
nand U5418 (N_5418,N_3743,N_3331);
and U5419 (N_5419,N_4498,N_4425);
nand U5420 (N_5420,N_4428,N_3984);
xor U5421 (N_5421,N_3907,N_4198);
or U5422 (N_5422,N_3468,N_3847);
xnor U5423 (N_5423,N_4169,N_4353);
and U5424 (N_5424,N_3221,N_4203);
and U5425 (N_5425,N_4143,N_3198);
nor U5426 (N_5426,N_4015,N_3940);
xnor U5427 (N_5427,N_4414,N_4234);
and U5428 (N_5428,N_3782,N_4324);
or U5429 (N_5429,N_3644,N_4473);
and U5430 (N_5430,N_3477,N_4172);
xnor U5431 (N_5431,N_3579,N_3676);
nor U5432 (N_5432,N_3606,N_3563);
xnor U5433 (N_5433,N_3001,N_3391);
nand U5434 (N_5434,N_3302,N_4285);
nor U5435 (N_5435,N_3226,N_3389);
nor U5436 (N_5436,N_3560,N_3907);
xnor U5437 (N_5437,N_3174,N_4333);
and U5438 (N_5438,N_3728,N_4087);
or U5439 (N_5439,N_3157,N_3500);
and U5440 (N_5440,N_4439,N_4042);
or U5441 (N_5441,N_3291,N_3535);
and U5442 (N_5442,N_4194,N_3850);
and U5443 (N_5443,N_3044,N_4173);
nand U5444 (N_5444,N_3679,N_3214);
and U5445 (N_5445,N_3795,N_3771);
or U5446 (N_5446,N_3169,N_3288);
nand U5447 (N_5447,N_3998,N_3308);
and U5448 (N_5448,N_4404,N_3257);
xnor U5449 (N_5449,N_3391,N_3406);
or U5450 (N_5450,N_3082,N_4368);
nand U5451 (N_5451,N_3804,N_3862);
xnor U5452 (N_5452,N_3061,N_3396);
and U5453 (N_5453,N_4325,N_3338);
nor U5454 (N_5454,N_3081,N_3066);
xor U5455 (N_5455,N_4133,N_3825);
nand U5456 (N_5456,N_4077,N_3897);
nor U5457 (N_5457,N_4041,N_3538);
and U5458 (N_5458,N_3818,N_3417);
or U5459 (N_5459,N_3376,N_3933);
xnor U5460 (N_5460,N_3252,N_3935);
nor U5461 (N_5461,N_3762,N_3295);
nand U5462 (N_5462,N_3533,N_3659);
nor U5463 (N_5463,N_3846,N_3394);
and U5464 (N_5464,N_3584,N_4479);
nand U5465 (N_5465,N_3457,N_3047);
nor U5466 (N_5466,N_3048,N_3938);
and U5467 (N_5467,N_3940,N_3327);
nor U5468 (N_5468,N_4131,N_3064);
xor U5469 (N_5469,N_4246,N_4105);
xnor U5470 (N_5470,N_3932,N_3525);
or U5471 (N_5471,N_3346,N_3441);
and U5472 (N_5472,N_3748,N_4265);
nand U5473 (N_5473,N_4108,N_4449);
and U5474 (N_5474,N_4298,N_4152);
xnor U5475 (N_5475,N_4324,N_3859);
xor U5476 (N_5476,N_3870,N_4490);
xor U5477 (N_5477,N_3128,N_3163);
or U5478 (N_5478,N_4218,N_3582);
or U5479 (N_5479,N_4356,N_3546);
nand U5480 (N_5480,N_3196,N_3572);
or U5481 (N_5481,N_4094,N_3985);
nand U5482 (N_5482,N_4112,N_3137);
and U5483 (N_5483,N_3741,N_3779);
xor U5484 (N_5484,N_3343,N_4452);
xnor U5485 (N_5485,N_3978,N_3878);
nand U5486 (N_5486,N_4293,N_3701);
or U5487 (N_5487,N_4481,N_4185);
or U5488 (N_5488,N_3241,N_3403);
and U5489 (N_5489,N_3692,N_3779);
or U5490 (N_5490,N_4331,N_3439);
nor U5491 (N_5491,N_4275,N_3840);
and U5492 (N_5492,N_4173,N_4450);
xor U5493 (N_5493,N_3339,N_4109);
xor U5494 (N_5494,N_3656,N_3149);
and U5495 (N_5495,N_3368,N_3471);
or U5496 (N_5496,N_3428,N_4280);
and U5497 (N_5497,N_4147,N_4249);
xnor U5498 (N_5498,N_3067,N_4426);
nand U5499 (N_5499,N_3079,N_3856);
and U5500 (N_5500,N_4462,N_3814);
and U5501 (N_5501,N_4138,N_3286);
nand U5502 (N_5502,N_3433,N_4126);
nor U5503 (N_5503,N_3607,N_4042);
and U5504 (N_5504,N_4113,N_3130);
nand U5505 (N_5505,N_3680,N_4427);
nor U5506 (N_5506,N_4285,N_4233);
nand U5507 (N_5507,N_3012,N_3306);
nand U5508 (N_5508,N_3324,N_4361);
xnor U5509 (N_5509,N_4282,N_3079);
xnor U5510 (N_5510,N_3094,N_4341);
or U5511 (N_5511,N_3118,N_4144);
and U5512 (N_5512,N_4328,N_3323);
nor U5513 (N_5513,N_3010,N_4052);
xnor U5514 (N_5514,N_3554,N_4393);
nand U5515 (N_5515,N_3062,N_4441);
nor U5516 (N_5516,N_3539,N_3123);
nor U5517 (N_5517,N_4427,N_4311);
xnor U5518 (N_5518,N_3183,N_3575);
or U5519 (N_5519,N_3450,N_4413);
nand U5520 (N_5520,N_4188,N_3109);
xor U5521 (N_5521,N_4461,N_4332);
or U5522 (N_5522,N_3934,N_3002);
nand U5523 (N_5523,N_3749,N_3557);
and U5524 (N_5524,N_4438,N_3769);
or U5525 (N_5525,N_3959,N_3285);
and U5526 (N_5526,N_4197,N_3278);
or U5527 (N_5527,N_3669,N_3815);
nor U5528 (N_5528,N_3422,N_3604);
nand U5529 (N_5529,N_3158,N_3860);
nand U5530 (N_5530,N_3176,N_3005);
xor U5531 (N_5531,N_3061,N_4194);
or U5532 (N_5532,N_4418,N_3252);
xnor U5533 (N_5533,N_3087,N_4201);
and U5534 (N_5534,N_4247,N_3054);
and U5535 (N_5535,N_3505,N_4016);
nor U5536 (N_5536,N_3843,N_4478);
or U5537 (N_5537,N_4331,N_3391);
xor U5538 (N_5538,N_3759,N_3871);
xor U5539 (N_5539,N_4089,N_4235);
and U5540 (N_5540,N_3576,N_3815);
xor U5541 (N_5541,N_3574,N_4209);
xor U5542 (N_5542,N_3645,N_4131);
xnor U5543 (N_5543,N_4027,N_3696);
and U5544 (N_5544,N_3234,N_3209);
xor U5545 (N_5545,N_4227,N_3611);
or U5546 (N_5546,N_3459,N_3660);
xnor U5547 (N_5547,N_3273,N_3057);
nor U5548 (N_5548,N_3801,N_3405);
nor U5549 (N_5549,N_3832,N_3379);
or U5550 (N_5550,N_3831,N_4231);
and U5551 (N_5551,N_3750,N_3717);
or U5552 (N_5552,N_3148,N_3735);
or U5553 (N_5553,N_4012,N_3263);
xor U5554 (N_5554,N_4367,N_3415);
nor U5555 (N_5555,N_4043,N_3760);
and U5556 (N_5556,N_3847,N_3688);
xor U5557 (N_5557,N_3602,N_3186);
xnor U5558 (N_5558,N_3019,N_4046);
nor U5559 (N_5559,N_3228,N_4044);
and U5560 (N_5560,N_3716,N_3744);
nor U5561 (N_5561,N_3178,N_3671);
and U5562 (N_5562,N_4382,N_3321);
and U5563 (N_5563,N_3990,N_3459);
or U5564 (N_5564,N_4254,N_3786);
or U5565 (N_5565,N_4474,N_4164);
nand U5566 (N_5566,N_4329,N_3882);
nand U5567 (N_5567,N_3047,N_3157);
and U5568 (N_5568,N_3290,N_3104);
nor U5569 (N_5569,N_3993,N_3530);
and U5570 (N_5570,N_3946,N_4155);
or U5571 (N_5571,N_3369,N_3447);
and U5572 (N_5572,N_3686,N_3081);
nand U5573 (N_5573,N_3300,N_3349);
and U5574 (N_5574,N_3837,N_4135);
and U5575 (N_5575,N_3735,N_3335);
xor U5576 (N_5576,N_3315,N_4178);
nor U5577 (N_5577,N_3410,N_4285);
nor U5578 (N_5578,N_4271,N_3749);
nand U5579 (N_5579,N_4014,N_3716);
nand U5580 (N_5580,N_4270,N_4091);
or U5581 (N_5581,N_3573,N_4428);
xnor U5582 (N_5582,N_4020,N_3560);
nor U5583 (N_5583,N_3804,N_3364);
or U5584 (N_5584,N_4178,N_4003);
nand U5585 (N_5585,N_3510,N_4306);
and U5586 (N_5586,N_3039,N_3316);
and U5587 (N_5587,N_3311,N_3162);
and U5588 (N_5588,N_3478,N_4480);
and U5589 (N_5589,N_4206,N_3589);
and U5590 (N_5590,N_3518,N_3557);
nand U5591 (N_5591,N_3252,N_4108);
nor U5592 (N_5592,N_3915,N_3788);
and U5593 (N_5593,N_4224,N_3456);
xor U5594 (N_5594,N_3136,N_3558);
or U5595 (N_5595,N_4032,N_3780);
nand U5596 (N_5596,N_3278,N_3803);
and U5597 (N_5597,N_3668,N_3852);
xnor U5598 (N_5598,N_3798,N_4367);
nor U5599 (N_5599,N_4082,N_3648);
and U5600 (N_5600,N_3223,N_3934);
nor U5601 (N_5601,N_3762,N_3348);
nor U5602 (N_5602,N_3313,N_4421);
nor U5603 (N_5603,N_3812,N_4373);
or U5604 (N_5604,N_4270,N_4169);
or U5605 (N_5605,N_4381,N_3053);
and U5606 (N_5606,N_3452,N_3488);
xor U5607 (N_5607,N_3261,N_4444);
nand U5608 (N_5608,N_4186,N_3296);
or U5609 (N_5609,N_3919,N_3607);
xor U5610 (N_5610,N_3324,N_3554);
xor U5611 (N_5611,N_3425,N_3766);
nand U5612 (N_5612,N_4248,N_4498);
or U5613 (N_5613,N_3303,N_3362);
nand U5614 (N_5614,N_3836,N_3189);
xor U5615 (N_5615,N_3459,N_4102);
and U5616 (N_5616,N_3216,N_3387);
nor U5617 (N_5617,N_4360,N_3683);
nand U5618 (N_5618,N_3950,N_3521);
xor U5619 (N_5619,N_3895,N_4318);
and U5620 (N_5620,N_3738,N_3138);
nand U5621 (N_5621,N_4460,N_4248);
and U5622 (N_5622,N_3590,N_3199);
nor U5623 (N_5623,N_3962,N_4304);
and U5624 (N_5624,N_4465,N_3284);
xor U5625 (N_5625,N_3133,N_3608);
xor U5626 (N_5626,N_3707,N_3700);
nor U5627 (N_5627,N_4369,N_3409);
and U5628 (N_5628,N_3754,N_4176);
xnor U5629 (N_5629,N_4404,N_3162);
nor U5630 (N_5630,N_4385,N_3286);
nand U5631 (N_5631,N_4285,N_4056);
xor U5632 (N_5632,N_3090,N_3135);
or U5633 (N_5633,N_4329,N_3625);
nor U5634 (N_5634,N_3612,N_3562);
nor U5635 (N_5635,N_3008,N_3403);
xor U5636 (N_5636,N_4115,N_3846);
nor U5637 (N_5637,N_3864,N_3798);
nand U5638 (N_5638,N_3493,N_3886);
and U5639 (N_5639,N_3889,N_3936);
nand U5640 (N_5640,N_3649,N_3974);
xnor U5641 (N_5641,N_3189,N_3081);
nand U5642 (N_5642,N_3219,N_4213);
xnor U5643 (N_5643,N_3115,N_3140);
xnor U5644 (N_5644,N_4063,N_3404);
nor U5645 (N_5645,N_3491,N_3966);
and U5646 (N_5646,N_3836,N_3894);
or U5647 (N_5647,N_3350,N_3229);
or U5648 (N_5648,N_4036,N_3418);
or U5649 (N_5649,N_3677,N_3133);
nor U5650 (N_5650,N_4398,N_4031);
nor U5651 (N_5651,N_4207,N_4304);
nand U5652 (N_5652,N_3162,N_3887);
nor U5653 (N_5653,N_4370,N_4151);
nand U5654 (N_5654,N_3358,N_4111);
and U5655 (N_5655,N_4247,N_3491);
and U5656 (N_5656,N_3703,N_3059);
and U5657 (N_5657,N_3899,N_4043);
or U5658 (N_5658,N_3298,N_4340);
or U5659 (N_5659,N_4241,N_4230);
nor U5660 (N_5660,N_3897,N_3613);
xnor U5661 (N_5661,N_4460,N_3324);
and U5662 (N_5662,N_4298,N_3103);
nor U5663 (N_5663,N_3134,N_3307);
nand U5664 (N_5664,N_4377,N_4392);
and U5665 (N_5665,N_4456,N_3659);
nor U5666 (N_5666,N_3276,N_3087);
or U5667 (N_5667,N_3683,N_3366);
nand U5668 (N_5668,N_4163,N_4476);
nand U5669 (N_5669,N_3326,N_3097);
or U5670 (N_5670,N_3942,N_3310);
nor U5671 (N_5671,N_3231,N_3914);
xnor U5672 (N_5672,N_3706,N_4359);
and U5673 (N_5673,N_4274,N_3974);
or U5674 (N_5674,N_3898,N_3429);
and U5675 (N_5675,N_4140,N_3996);
or U5676 (N_5676,N_3378,N_3365);
and U5677 (N_5677,N_3246,N_3204);
and U5678 (N_5678,N_3734,N_3416);
and U5679 (N_5679,N_3933,N_4048);
nor U5680 (N_5680,N_4037,N_3834);
and U5681 (N_5681,N_3219,N_4435);
nor U5682 (N_5682,N_4367,N_3879);
nand U5683 (N_5683,N_3590,N_3601);
and U5684 (N_5684,N_3166,N_3112);
nand U5685 (N_5685,N_3207,N_4323);
nand U5686 (N_5686,N_3538,N_3180);
nand U5687 (N_5687,N_4122,N_3199);
and U5688 (N_5688,N_3799,N_3410);
and U5689 (N_5689,N_3070,N_4437);
xor U5690 (N_5690,N_4426,N_3792);
nor U5691 (N_5691,N_3921,N_4469);
and U5692 (N_5692,N_3123,N_3824);
nor U5693 (N_5693,N_4170,N_3794);
and U5694 (N_5694,N_4178,N_3945);
or U5695 (N_5695,N_3248,N_3138);
xor U5696 (N_5696,N_3156,N_3223);
and U5697 (N_5697,N_3158,N_3022);
nor U5698 (N_5698,N_3802,N_4013);
and U5699 (N_5699,N_3300,N_4244);
or U5700 (N_5700,N_3681,N_4240);
nand U5701 (N_5701,N_3082,N_4476);
or U5702 (N_5702,N_3267,N_4024);
and U5703 (N_5703,N_4380,N_4397);
xor U5704 (N_5704,N_4156,N_3249);
nor U5705 (N_5705,N_3964,N_4014);
and U5706 (N_5706,N_3713,N_3123);
and U5707 (N_5707,N_3827,N_3313);
or U5708 (N_5708,N_4045,N_4012);
and U5709 (N_5709,N_3241,N_3556);
nor U5710 (N_5710,N_3896,N_3109);
nand U5711 (N_5711,N_3016,N_4209);
nor U5712 (N_5712,N_3170,N_3647);
and U5713 (N_5713,N_3291,N_3480);
nor U5714 (N_5714,N_3484,N_3414);
or U5715 (N_5715,N_3243,N_4178);
and U5716 (N_5716,N_3010,N_3218);
or U5717 (N_5717,N_3045,N_3888);
nor U5718 (N_5718,N_3232,N_3841);
and U5719 (N_5719,N_3617,N_3313);
or U5720 (N_5720,N_4205,N_3403);
and U5721 (N_5721,N_4438,N_3812);
nand U5722 (N_5722,N_4417,N_3422);
or U5723 (N_5723,N_3311,N_4011);
and U5724 (N_5724,N_4181,N_4303);
and U5725 (N_5725,N_4167,N_3120);
nor U5726 (N_5726,N_3083,N_3275);
and U5727 (N_5727,N_4091,N_3230);
or U5728 (N_5728,N_3867,N_4388);
xor U5729 (N_5729,N_3282,N_4231);
nand U5730 (N_5730,N_3087,N_3096);
nor U5731 (N_5731,N_3298,N_3244);
nand U5732 (N_5732,N_3933,N_3909);
nor U5733 (N_5733,N_3057,N_4298);
and U5734 (N_5734,N_3934,N_4339);
nor U5735 (N_5735,N_3635,N_3257);
nor U5736 (N_5736,N_3822,N_3417);
nor U5737 (N_5737,N_3797,N_4035);
and U5738 (N_5738,N_3834,N_3688);
nor U5739 (N_5739,N_3098,N_3908);
nand U5740 (N_5740,N_4186,N_3948);
nand U5741 (N_5741,N_3540,N_3271);
or U5742 (N_5742,N_3146,N_4095);
or U5743 (N_5743,N_3279,N_3567);
nand U5744 (N_5744,N_3914,N_3752);
or U5745 (N_5745,N_4129,N_4124);
or U5746 (N_5746,N_3536,N_3728);
nand U5747 (N_5747,N_4486,N_3722);
xor U5748 (N_5748,N_3493,N_3530);
or U5749 (N_5749,N_4131,N_4481);
and U5750 (N_5750,N_3949,N_3154);
nand U5751 (N_5751,N_3275,N_4239);
xnor U5752 (N_5752,N_3322,N_3645);
nand U5753 (N_5753,N_3806,N_3589);
or U5754 (N_5754,N_4118,N_4080);
nor U5755 (N_5755,N_3756,N_3314);
nor U5756 (N_5756,N_4453,N_3796);
nand U5757 (N_5757,N_4084,N_4115);
nand U5758 (N_5758,N_3876,N_3590);
nor U5759 (N_5759,N_3766,N_3492);
nand U5760 (N_5760,N_3389,N_3138);
nor U5761 (N_5761,N_3867,N_3001);
or U5762 (N_5762,N_3133,N_3405);
and U5763 (N_5763,N_3596,N_4294);
nand U5764 (N_5764,N_4280,N_3626);
nor U5765 (N_5765,N_3855,N_3945);
xnor U5766 (N_5766,N_3587,N_3091);
and U5767 (N_5767,N_4100,N_4486);
xnor U5768 (N_5768,N_3448,N_4462);
nor U5769 (N_5769,N_3259,N_3914);
nor U5770 (N_5770,N_3398,N_4208);
or U5771 (N_5771,N_3877,N_4416);
and U5772 (N_5772,N_3042,N_4238);
nor U5773 (N_5773,N_3457,N_4115);
nand U5774 (N_5774,N_3765,N_3350);
nor U5775 (N_5775,N_4325,N_3137);
or U5776 (N_5776,N_3367,N_3763);
nor U5777 (N_5777,N_4013,N_3219);
nor U5778 (N_5778,N_3342,N_3358);
nor U5779 (N_5779,N_4157,N_4354);
xor U5780 (N_5780,N_4038,N_3976);
or U5781 (N_5781,N_4068,N_3832);
nor U5782 (N_5782,N_3173,N_4449);
and U5783 (N_5783,N_4021,N_4379);
nor U5784 (N_5784,N_4493,N_3613);
and U5785 (N_5785,N_3534,N_3822);
nor U5786 (N_5786,N_3630,N_4338);
nor U5787 (N_5787,N_3966,N_4376);
and U5788 (N_5788,N_4002,N_4078);
xnor U5789 (N_5789,N_3084,N_3149);
nor U5790 (N_5790,N_4086,N_3522);
nand U5791 (N_5791,N_4226,N_3356);
or U5792 (N_5792,N_4451,N_3149);
nand U5793 (N_5793,N_3832,N_4177);
or U5794 (N_5794,N_4327,N_4032);
xnor U5795 (N_5795,N_3283,N_4407);
xor U5796 (N_5796,N_3811,N_3963);
nor U5797 (N_5797,N_3855,N_3648);
nand U5798 (N_5798,N_3662,N_3033);
or U5799 (N_5799,N_3433,N_4468);
xnor U5800 (N_5800,N_3627,N_3012);
nand U5801 (N_5801,N_4422,N_3538);
nand U5802 (N_5802,N_4344,N_4332);
nand U5803 (N_5803,N_4165,N_3406);
nor U5804 (N_5804,N_4126,N_4192);
xor U5805 (N_5805,N_3148,N_4037);
nor U5806 (N_5806,N_3339,N_3831);
xor U5807 (N_5807,N_3639,N_3024);
nand U5808 (N_5808,N_3653,N_3082);
nand U5809 (N_5809,N_4356,N_3840);
nand U5810 (N_5810,N_3471,N_3911);
and U5811 (N_5811,N_3638,N_3748);
nor U5812 (N_5812,N_4484,N_3343);
and U5813 (N_5813,N_3409,N_4496);
nand U5814 (N_5814,N_4038,N_3649);
nand U5815 (N_5815,N_4493,N_3896);
nand U5816 (N_5816,N_3609,N_3396);
or U5817 (N_5817,N_4362,N_4267);
nor U5818 (N_5818,N_4358,N_4490);
and U5819 (N_5819,N_4020,N_3035);
xnor U5820 (N_5820,N_3609,N_4338);
or U5821 (N_5821,N_4185,N_4043);
or U5822 (N_5822,N_3507,N_3100);
nand U5823 (N_5823,N_4321,N_4342);
or U5824 (N_5824,N_4275,N_3994);
xor U5825 (N_5825,N_3852,N_3957);
or U5826 (N_5826,N_3117,N_3243);
nor U5827 (N_5827,N_3683,N_3680);
nand U5828 (N_5828,N_3055,N_3480);
nor U5829 (N_5829,N_3544,N_3125);
xor U5830 (N_5830,N_4234,N_3655);
xnor U5831 (N_5831,N_3080,N_4140);
nand U5832 (N_5832,N_4436,N_4484);
nand U5833 (N_5833,N_4455,N_3880);
or U5834 (N_5834,N_3319,N_3188);
nand U5835 (N_5835,N_4446,N_3526);
xor U5836 (N_5836,N_3743,N_3293);
nand U5837 (N_5837,N_4203,N_3265);
nand U5838 (N_5838,N_3098,N_4457);
nor U5839 (N_5839,N_3448,N_4402);
nor U5840 (N_5840,N_3643,N_3948);
nand U5841 (N_5841,N_3005,N_3538);
nor U5842 (N_5842,N_4432,N_4209);
nand U5843 (N_5843,N_3269,N_3215);
and U5844 (N_5844,N_4422,N_3143);
xnor U5845 (N_5845,N_4061,N_3334);
nor U5846 (N_5846,N_3797,N_3896);
xor U5847 (N_5847,N_3207,N_3507);
xor U5848 (N_5848,N_3020,N_4084);
and U5849 (N_5849,N_4280,N_3388);
nor U5850 (N_5850,N_3050,N_3051);
xnor U5851 (N_5851,N_3268,N_3248);
nor U5852 (N_5852,N_4256,N_3714);
xor U5853 (N_5853,N_3719,N_3683);
nor U5854 (N_5854,N_4251,N_3319);
nor U5855 (N_5855,N_3664,N_3959);
or U5856 (N_5856,N_4246,N_4286);
or U5857 (N_5857,N_3735,N_3476);
nor U5858 (N_5858,N_3123,N_3851);
nor U5859 (N_5859,N_3269,N_3232);
or U5860 (N_5860,N_3057,N_3443);
xor U5861 (N_5861,N_3079,N_3775);
xor U5862 (N_5862,N_3948,N_4091);
nand U5863 (N_5863,N_3836,N_3870);
nor U5864 (N_5864,N_4446,N_3634);
nand U5865 (N_5865,N_3055,N_3102);
and U5866 (N_5866,N_4047,N_3542);
xor U5867 (N_5867,N_3947,N_3571);
nand U5868 (N_5868,N_4438,N_3981);
xnor U5869 (N_5869,N_3384,N_3876);
and U5870 (N_5870,N_4163,N_3727);
nor U5871 (N_5871,N_3085,N_3576);
nand U5872 (N_5872,N_3027,N_4379);
or U5873 (N_5873,N_4144,N_4405);
xnor U5874 (N_5874,N_3648,N_3419);
nand U5875 (N_5875,N_3794,N_3140);
nor U5876 (N_5876,N_3077,N_4169);
and U5877 (N_5877,N_3931,N_3007);
nor U5878 (N_5878,N_4079,N_3672);
nand U5879 (N_5879,N_4126,N_3203);
or U5880 (N_5880,N_3256,N_3177);
or U5881 (N_5881,N_3784,N_3609);
or U5882 (N_5882,N_4377,N_4048);
or U5883 (N_5883,N_3837,N_3659);
nor U5884 (N_5884,N_3022,N_3249);
and U5885 (N_5885,N_4456,N_4265);
nor U5886 (N_5886,N_3961,N_3284);
xor U5887 (N_5887,N_3724,N_3662);
nand U5888 (N_5888,N_4189,N_3249);
nor U5889 (N_5889,N_3997,N_3482);
nor U5890 (N_5890,N_3668,N_3160);
nor U5891 (N_5891,N_3342,N_4081);
or U5892 (N_5892,N_4436,N_3299);
and U5893 (N_5893,N_4084,N_4015);
xor U5894 (N_5894,N_3369,N_4111);
nand U5895 (N_5895,N_3948,N_3106);
nand U5896 (N_5896,N_3627,N_3389);
nand U5897 (N_5897,N_4448,N_4350);
nor U5898 (N_5898,N_3870,N_3546);
or U5899 (N_5899,N_3590,N_3096);
or U5900 (N_5900,N_3132,N_3557);
and U5901 (N_5901,N_3863,N_3350);
xnor U5902 (N_5902,N_3892,N_3197);
nand U5903 (N_5903,N_3207,N_4191);
or U5904 (N_5904,N_3093,N_3052);
nor U5905 (N_5905,N_3660,N_3525);
nor U5906 (N_5906,N_3985,N_4288);
xor U5907 (N_5907,N_3220,N_3606);
and U5908 (N_5908,N_3553,N_4017);
or U5909 (N_5909,N_3350,N_4248);
or U5910 (N_5910,N_3564,N_4019);
and U5911 (N_5911,N_3397,N_3477);
nor U5912 (N_5912,N_3139,N_3499);
and U5913 (N_5913,N_3182,N_3027);
and U5914 (N_5914,N_4002,N_3077);
and U5915 (N_5915,N_3556,N_3447);
or U5916 (N_5916,N_3706,N_4010);
and U5917 (N_5917,N_3306,N_4385);
or U5918 (N_5918,N_3364,N_3220);
nor U5919 (N_5919,N_4044,N_3493);
nand U5920 (N_5920,N_3944,N_4355);
nor U5921 (N_5921,N_3004,N_3851);
or U5922 (N_5922,N_4279,N_3116);
or U5923 (N_5923,N_3318,N_4217);
or U5924 (N_5924,N_3061,N_3701);
or U5925 (N_5925,N_3432,N_4441);
nor U5926 (N_5926,N_4392,N_3022);
or U5927 (N_5927,N_3607,N_3879);
or U5928 (N_5928,N_4115,N_3625);
nor U5929 (N_5929,N_3434,N_3746);
nand U5930 (N_5930,N_3639,N_4448);
nand U5931 (N_5931,N_3890,N_3931);
nor U5932 (N_5932,N_3528,N_3215);
nand U5933 (N_5933,N_4011,N_3262);
nor U5934 (N_5934,N_4003,N_4060);
and U5935 (N_5935,N_3569,N_4417);
and U5936 (N_5936,N_4190,N_4058);
or U5937 (N_5937,N_3549,N_3345);
nand U5938 (N_5938,N_4117,N_3491);
or U5939 (N_5939,N_4063,N_3956);
nor U5940 (N_5940,N_4374,N_4471);
nor U5941 (N_5941,N_3215,N_4231);
xnor U5942 (N_5942,N_3157,N_4260);
or U5943 (N_5943,N_4092,N_3017);
and U5944 (N_5944,N_4265,N_4134);
nand U5945 (N_5945,N_3052,N_3203);
or U5946 (N_5946,N_4204,N_4088);
nand U5947 (N_5947,N_4245,N_3309);
nand U5948 (N_5948,N_3792,N_4467);
nor U5949 (N_5949,N_3559,N_4281);
or U5950 (N_5950,N_3243,N_3289);
and U5951 (N_5951,N_3012,N_3158);
or U5952 (N_5952,N_4052,N_3387);
nand U5953 (N_5953,N_3811,N_3059);
xor U5954 (N_5954,N_3446,N_3190);
or U5955 (N_5955,N_3260,N_4197);
nand U5956 (N_5956,N_3557,N_3490);
and U5957 (N_5957,N_3164,N_3816);
xnor U5958 (N_5958,N_3886,N_4442);
nand U5959 (N_5959,N_3523,N_4327);
or U5960 (N_5960,N_3903,N_3625);
nor U5961 (N_5961,N_3806,N_3029);
nand U5962 (N_5962,N_3682,N_3608);
or U5963 (N_5963,N_4313,N_4455);
and U5964 (N_5964,N_4141,N_4355);
and U5965 (N_5965,N_3598,N_3169);
nand U5966 (N_5966,N_3856,N_3151);
nand U5967 (N_5967,N_3568,N_3120);
and U5968 (N_5968,N_4067,N_3387);
nor U5969 (N_5969,N_4250,N_3681);
nand U5970 (N_5970,N_3360,N_3091);
or U5971 (N_5971,N_4039,N_3902);
nand U5972 (N_5972,N_3884,N_3449);
nand U5973 (N_5973,N_3729,N_3231);
nor U5974 (N_5974,N_3570,N_3421);
nand U5975 (N_5975,N_3757,N_4014);
and U5976 (N_5976,N_3013,N_3962);
xor U5977 (N_5977,N_3146,N_4403);
xnor U5978 (N_5978,N_4247,N_4459);
xnor U5979 (N_5979,N_3333,N_3283);
or U5980 (N_5980,N_4305,N_3551);
nor U5981 (N_5981,N_4295,N_3884);
xor U5982 (N_5982,N_3937,N_4276);
nor U5983 (N_5983,N_4146,N_3409);
nand U5984 (N_5984,N_3391,N_3399);
nor U5985 (N_5985,N_3426,N_4475);
or U5986 (N_5986,N_4348,N_4388);
xnor U5987 (N_5987,N_3087,N_3609);
nor U5988 (N_5988,N_4251,N_3384);
and U5989 (N_5989,N_4096,N_4414);
xnor U5990 (N_5990,N_4027,N_4024);
xor U5991 (N_5991,N_3275,N_3136);
nor U5992 (N_5992,N_3410,N_3591);
nand U5993 (N_5993,N_3369,N_3968);
xnor U5994 (N_5994,N_3660,N_4375);
nor U5995 (N_5995,N_4115,N_3957);
or U5996 (N_5996,N_4087,N_4154);
or U5997 (N_5997,N_3394,N_4338);
or U5998 (N_5998,N_3906,N_3347);
nor U5999 (N_5999,N_4149,N_3708);
or U6000 (N_6000,N_5797,N_5520);
xor U6001 (N_6001,N_4734,N_5214);
and U6002 (N_6002,N_5044,N_4895);
or U6003 (N_6003,N_4668,N_4636);
or U6004 (N_6004,N_5069,N_4696);
and U6005 (N_6005,N_4924,N_5896);
or U6006 (N_6006,N_5762,N_5800);
or U6007 (N_6007,N_4915,N_4969);
or U6008 (N_6008,N_5879,N_5273);
nand U6009 (N_6009,N_4960,N_4842);
and U6010 (N_6010,N_5009,N_5497);
or U6011 (N_6011,N_4680,N_5733);
and U6012 (N_6012,N_5112,N_4580);
and U6013 (N_6013,N_5739,N_4747);
and U6014 (N_6014,N_4635,N_5300);
nand U6015 (N_6015,N_5967,N_5758);
and U6016 (N_6016,N_5564,N_5351);
nand U6017 (N_6017,N_5054,N_4810);
nand U6018 (N_6018,N_4932,N_4574);
or U6019 (N_6019,N_5996,N_4869);
or U6020 (N_6020,N_5597,N_5663);
nand U6021 (N_6021,N_5901,N_5842);
and U6022 (N_6022,N_5659,N_4703);
or U6023 (N_6023,N_5642,N_5122);
or U6024 (N_6024,N_4772,N_5827);
nand U6025 (N_6025,N_4971,N_5518);
or U6026 (N_6026,N_4504,N_5360);
nand U6027 (N_6027,N_5655,N_4846);
and U6028 (N_6028,N_5860,N_5265);
or U6029 (N_6029,N_4594,N_5899);
nor U6030 (N_6030,N_5324,N_5319);
or U6031 (N_6031,N_5923,N_4847);
xor U6032 (N_6032,N_5403,N_4687);
nand U6033 (N_6033,N_4515,N_4914);
xor U6034 (N_6034,N_5169,N_5666);
or U6035 (N_6035,N_5257,N_4547);
or U6036 (N_6036,N_5230,N_5181);
nand U6037 (N_6037,N_5085,N_5333);
xnor U6038 (N_6038,N_5955,N_5872);
xnor U6039 (N_6039,N_5960,N_5378);
xor U6040 (N_6040,N_5455,N_5315);
and U6041 (N_6041,N_4795,N_5250);
nand U6042 (N_6042,N_5660,N_5185);
or U6043 (N_6043,N_5845,N_4959);
xnor U6044 (N_6044,N_5502,N_5920);
nand U6045 (N_6045,N_5875,N_5201);
nand U6046 (N_6046,N_5880,N_4714);
nor U6047 (N_6047,N_4566,N_4723);
xor U6048 (N_6048,N_5462,N_4508);
and U6049 (N_6049,N_4667,N_4642);
nand U6050 (N_6050,N_5825,N_4849);
xnor U6051 (N_6051,N_5893,N_5486);
nand U6052 (N_6052,N_5843,N_5386);
and U6053 (N_6053,N_4964,N_5368);
or U6054 (N_6054,N_5523,N_5033);
and U6055 (N_6055,N_4740,N_5638);
nand U6056 (N_6056,N_5195,N_4627);
or U6057 (N_6057,N_4792,N_4682);
and U6058 (N_6058,N_4560,N_5731);
nor U6059 (N_6059,N_5219,N_5567);
nand U6060 (N_6060,N_4608,N_5534);
or U6061 (N_6061,N_4856,N_5939);
or U6062 (N_6062,N_4808,N_5090);
and U6063 (N_6063,N_4735,N_4709);
and U6064 (N_6064,N_5260,N_5695);
or U6065 (N_6065,N_5709,N_5191);
or U6066 (N_6066,N_5808,N_4602);
or U6067 (N_6067,N_4758,N_5132);
nor U6068 (N_6068,N_5237,N_4596);
nor U6069 (N_6069,N_5989,N_5473);
or U6070 (N_6070,N_5010,N_5743);
or U6071 (N_6071,N_5160,N_5051);
xor U6072 (N_6072,N_5590,N_5352);
xnor U6073 (N_6073,N_4748,N_5463);
xnor U6074 (N_6074,N_5392,N_5116);
xor U6075 (N_6075,N_5376,N_4834);
nand U6076 (N_6076,N_5513,N_5287);
xor U6077 (N_6077,N_5938,N_5338);
nor U6078 (N_6078,N_5772,N_5350);
and U6079 (N_6079,N_4841,N_4939);
or U6080 (N_6080,N_4633,N_5754);
xnor U6081 (N_6081,N_5434,N_4955);
nor U6082 (N_6082,N_5080,N_5226);
and U6083 (N_6083,N_5799,N_5504);
nor U6084 (N_6084,N_5173,N_5970);
or U6085 (N_6085,N_5027,N_4943);
or U6086 (N_6086,N_5373,N_5865);
and U6087 (N_6087,N_5339,N_5117);
xnor U6088 (N_6088,N_5038,N_5328);
nor U6089 (N_6089,N_5714,N_5838);
nand U6090 (N_6090,N_5212,N_4870);
xor U6091 (N_6091,N_4835,N_5482);
nor U6092 (N_6092,N_4880,N_4718);
or U6093 (N_6093,N_5229,N_5929);
and U6094 (N_6094,N_5785,N_5423);
nand U6095 (N_6095,N_4876,N_5162);
nor U6096 (N_6096,N_4579,N_5442);
nand U6097 (N_6097,N_5438,N_5947);
xor U6098 (N_6098,N_5425,N_5064);
xnor U6099 (N_6099,N_5533,N_5798);
and U6100 (N_6100,N_5544,N_4889);
or U6101 (N_6101,N_5917,N_4698);
or U6102 (N_6102,N_5562,N_5952);
or U6103 (N_6103,N_5632,N_5155);
nor U6104 (N_6104,N_4583,N_5735);
xor U6105 (N_6105,N_5458,N_4770);
xnor U6106 (N_6106,N_5493,N_5599);
and U6107 (N_6107,N_5634,N_5931);
nand U6108 (N_6108,N_5956,N_4956);
nand U6109 (N_6109,N_5016,N_5720);
or U6110 (N_6110,N_5013,N_4991);
and U6111 (N_6111,N_5428,N_5427);
or U6112 (N_6112,N_4710,N_4731);
nand U6113 (N_6113,N_4637,N_5586);
or U6114 (N_6114,N_5248,N_4818);
or U6115 (N_6115,N_4521,N_4700);
nand U6116 (N_6116,N_4541,N_5715);
or U6117 (N_6117,N_5857,N_5503);
and U6118 (N_6118,N_5026,N_4858);
and U6119 (N_6119,N_4564,N_4517);
nand U6120 (N_6120,N_4581,N_5318);
or U6121 (N_6121,N_4561,N_4715);
nor U6122 (N_6122,N_5813,N_4528);
and U6123 (N_6123,N_4985,N_5224);
and U6124 (N_6124,N_5167,N_5252);
or U6125 (N_6125,N_4706,N_5949);
xor U6126 (N_6126,N_4823,N_5959);
nand U6127 (N_6127,N_5142,N_5835);
and U6128 (N_6128,N_4685,N_4609);
and U6129 (N_6129,N_5271,N_5419);
or U6130 (N_6130,N_4957,N_5579);
or U6131 (N_6131,N_4669,N_5216);
or U6132 (N_6132,N_5646,N_5820);
nor U6133 (N_6133,N_5873,N_4540);
or U6134 (N_6134,N_4712,N_5700);
nand U6135 (N_6135,N_5496,N_5344);
nand U6136 (N_6136,N_5672,N_5969);
nand U6137 (N_6137,N_5306,N_4514);
xnor U6138 (N_6138,N_5778,N_4784);
xor U6139 (N_6139,N_5537,N_5490);
xor U6140 (N_6140,N_4606,N_5029);
and U6141 (N_6141,N_4752,N_4531);
xor U6142 (N_6142,N_5926,N_4844);
nor U6143 (N_6143,N_4942,N_5635);
or U6144 (N_6144,N_5810,N_5187);
or U6145 (N_6145,N_5558,N_5043);
or U6146 (N_6146,N_5450,N_5833);
and U6147 (N_6147,N_5974,N_4790);
and U6148 (N_6148,N_5134,N_5035);
or U6149 (N_6149,N_5601,N_4916);
or U6150 (N_6150,N_5584,N_5102);
and U6151 (N_6151,N_4989,N_4565);
or U6152 (N_6152,N_5980,N_5846);
xor U6153 (N_6153,N_4645,N_5329);
nand U6154 (N_6154,N_5128,N_5449);
xor U6155 (N_6155,N_5528,N_5748);
xnor U6156 (N_6156,N_5270,N_5359);
and U6157 (N_6157,N_5998,N_4995);
or U6158 (N_6158,N_5478,N_4953);
or U6159 (N_6159,N_4587,N_5760);
and U6160 (N_6160,N_4891,N_5943);
and U6161 (N_6161,N_5574,N_5815);
and U6162 (N_6162,N_5406,N_5559);
xnor U6163 (N_6163,N_5025,N_5105);
or U6164 (N_6164,N_5445,N_4607);
nand U6165 (N_6165,N_5023,N_4569);
nand U6166 (N_6166,N_5501,N_5078);
nand U6167 (N_6167,N_5118,N_5147);
or U6168 (N_6168,N_4549,N_4526);
nor U6169 (N_6169,N_5942,N_5763);
xnor U6170 (N_6170,N_5750,N_5217);
nand U6171 (N_6171,N_5231,N_5653);
xnor U6172 (N_6172,N_5531,N_5258);
nor U6173 (N_6173,N_4997,N_5305);
nor U6174 (N_6174,N_5005,N_5578);
nor U6175 (N_6175,N_5603,N_5380);
and U6176 (N_6176,N_5232,N_4918);
nor U6177 (N_6177,N_5674,N_5809);
and U6178 (N_6178,N_5079,N_4763);
and U6179 (N_6179,N_5281,N_4940);
or U6180 (N_6180,N_5919,N_5288);
nor U6181 (N_6181,N_5247,N_5383);
and U6182 (N_6182,N_4728,N_5855);
xor U6183 (N_6183,N_5417,N_4611);
xnor U6184 (N_6184,N_5312,N_5277);
nand U6185 (N_6185,N_4807,N_5859);
nand U6186 (N_6186,N_4542,N_5264);
xor U6187 (N_6187,N_5510,N_4831);
nor U6188 (N_6188,N_5021,N_4513);
nor U6189 (N_6189,N_5215,N_5261);
or U6190 (N_6190,N_4769,N_5190);
and U6191 (N_6191,N_4644,N_5057);
xnor U6192 (N_6192,N_5335,N_5032);
nand U6193 (N_6193,N_5592,N_5863);
nor U6194 (N_6194,N_5936,N_5734);
nand U6195 (N_6195,N_5325,N_5067);
nor U6196 (N_6196,N_4934,N_5717);
or U6197 (N_6197,N_5506,N_5183);
and U6198 (N_6198,N_4737,N_5072);
nand U6199 (N_6199,N_5397,N_5178);
or U6200 (N_6200,N_5151,N_4791);
or U6201 (N_6201,N_5088,N_4716);
nor U6202 (N_6202,N_4990,N_5149);
or U6203 (N_6203,N_5961,N_5153);
nand U6204 (N_6204,N_4738,N_5727);
nor U6205 (N_6205,N_4519,N_4927);
nor U6206 (N_6206,N_4988,N_5805);
nor U6207 (N_6207,N_5157,N_5196);
nand U6208 (N_6208,N_5255,N_4938);
nor U6209 (N_6209,N_4979,N_4773);
and U6210 (N_6210,N_5984,N_5630);
nand U6211 (N_6211,N_4825,N_5911);
nor U6212 (N_6212,N_4872,N_5227);
nand U6213 (N_6213,N_4548,N_5158);
xor U6214 (N_6214,N_4648,N_4967);
nand U6215 (N_6215,N_4653,N_5882);
or U6216 (N_6216,N_4892,N_4518);
nor U6217 (N_6217,N_4638,N_5432);
nor U6218 (N_6218,N_5457,N_5436);
and U6219 (N_6219,N_4605,N_5823);
and U6220 (N_6220,N_4705,N_5404);
and U6221 (N_6221,N_5168,N_4701);
nor U6222 (N_6222,N_5588,N_5172);
or U6223 (N_6223,N_4659,N_4978);
and U6224 (N_6224,N_5652,N_4588);
xnor U6225 (N_6225,N_4983,N_4708);
nor U6226 (N_6226,N_4501,N_5240);
xnor U6227 (N_6227,N_5516,N_5055);
nor U6228 (N_6228,N_5332,N_5140);
or U6229 (N_6229,N_4597,N_4742);
xnor U6230 (N_6230,N_4720,N_4570);
or U6231 (N_6231,N_5096,N_5916);
nor U6232 (N_6232,N_4984,N_5444);
or U6233 (N_6233,N_4759,N_5017);
nor U6234 (N_6234,N_4593,N_5821);
and U6235 (N_6235,N_5362,N_5767);
or U6236 (N_6236,N_5795,N_5235);
nor U6237 (N_6237,N_5789,N_5806);
nor U6238 (N_6238,N_5964,N_4907);
nor U6239 (N_6239,N_5934,N_4655);
xnor U6240 (N_6240,N_5527,N_5909);
nor U6241 (N_6241,N_4950,N_5670);
nor U6242 (N_6242,N_5207,N_5613);
and U6243 (N_6243,N_4875,N_5186);
nand U6244 (N_6244,N_5243,N_4658);
or U6245 (N_6245,N_4800,N_4536);
nand U6246 (N_6246,N_4545,N_5782);
xnor U6247 (N_6247,N_4801,N_5651);
nand U6248 (N_6248,N_5278,N_4717);
and U6249 (N_6249,N_5361,N_5256);
xor U6250 (N_6250,N_4503,N_4539);
and U6251 (N_6251,N_5507,N_5125);
or U6252 (N_6252,N_4894,N_4704);
nor U6253 (N_6253,N_5978,N_5034);
nor U6254 (N_6254,N_4817,N_5903);
nand U6255 (N_6255,N_5020,N_4951);
nor U6256 (N_6256,N_5294,N_4511);
nand U6257 (N_6257,N_5794,N_5557);
or U6258 (N_6258,N_5259,N_5414);
xor U6259 (N_6259,N_5616,N_4629);
xnor U6260 (N_6260,N_4762,N_5648);
and U6261 (N_6261,N_5852,N_4600);
nor U6262 (N_6262,N_5894,N_5712);
and U6263 (N_6263,N_5921,N_4890);
xnor U6264 (N_6264,N_5114,N_4931);
nor U6265 (N_6265,N_4917,N_4502);
or U6266 (N_6266,N_5440,N_5394);
and U6267 (N_6267,N_5469,N_5776);
nor U6268 (N_6268,N_5885,N_5111);
or U6269 (N_6269,N_5460,N_5728);
nor U6270 (N_6270,N_5529,N_4903);
nor U6271 (N_6271,N_5900,N_5669);
and U6272 (N_6272,N_4986,N_4505);
xnor U6273 (N_6273,N_4603,N_5494);
and U6274 (N_6274,N_5089,N_4525);
xnor U6275 (N_6275,N_5566,N_5348);
xnor U6276 (N_6276,N_4778,N_4866);
and U6277 (N_6277,N_4885,N_5565);
nor U6278 (N_6278,N_4530,N_5738);
or U6279 (N_6279,N_4965,N_4524);
and U6280 (N_6280,N_5199,N_4838);
nand U6281 (N_6281,N_4908,N_5891);
nand U6282 (N_6282,N_5014,N_4584);
nand U6283 (N_6283,N_5621,N_5568);
nand U6284 (N_6284,N_5979,N_5757);
xnor U6285 (N_6285,N_5405,N_5365);
nor U6286 (N_6286,N_4722,N_5213);
and U6287 (N_6287,N_5127,N_5656);
and U6288 (N_6288,N_5550,N_5087);
or U6289 (N_6289,N_4725,N_5930);
xnor U6290 (N_6290,N_5391,N_5861);
or U6291 (N_6291,N_4992,N_4640);
nor U6292 (N_6292,N_5696,N_4905);
xnor U6293 (N_6293,N_4578,N_5103);
xor U6294 (N_6294,N_4557,N_5699);
and U6295 (N_6295,N_5123,N_4794);
nand U6296 (N_6296,N_4881,N_4516);
nor U6297 (N_6297,N_4688,N_5246);
nor U6298 (N_6298,N_5120,N_5161);
nor U6299 (N_6299,N_5729,N_5220);
and U6300 (N_6300,N_4961,N_4553);
nor U6301 (N_6301,N_5612,N_5992);
or U6302 (N_6302,N_4789,N_4532);
or U6303 (N_6303,N_4661,N_5316);
nor U6304 (N_6304,N_5061,N_5336);
or U6305 (N_6305,N_5596,N_5620);
nand U6306 (N_6306,N_5274,N_4973);
nor U6307 (N_6307,N_5390,N_5171);
nand U6308 (N_6308,N_5685,N_4904);
nand U6309 (N_6309,N_5965,N_4727);
or U6310 (N_6310,N_4601,N_5317);
xnor U6311 (N_6311,N_5396,N_5399);
nor U6312 (N_6312,N_4756,N_5184);
nand U6313 (N_6313,N_4691,N_5710);
nor U6314 (N_6314,N_4860,N_5000);
xor U6315 (N_6315,N_5472,N_4820);
and U6316 (N_6316,N_4926,N_5045);
and U6317 (N_6317,N_5898,N_5814);
xnor U6318 (N_6318,N_4780,N_5740);
nor U6319 (N_6319,N_5532,N_5517);
or U6320 (N_6320,N_4833,N_5234);
xor U6321 (N_6321,N_4863,N_5225);
nand U6322 (N_6322,N_4861,N_5573);
xor U6323 (N_6323,N_5293,N_4746);
nor U6324 (N_6324,N_5345,N_4686);
nor U6325 (N_6325,N_5349,N_5751);
and U6326 (N_6326,N_5869,N_5692);
or U6327 (N_6327,N_4862,N_5844);
and U6328 (N_6328,N_5137,N_5945);
and U6329 (N_6329,N_4556,N_5119);
xor U6330 (N_6330,N_4672,N_4976);
nor U6331 (N_6331,N_4851,N_5447);
and U6332 (N_6332,N_5953,N_5415);
or U6333 (N_6333,N_5571,N_4572);
or U6334 (N_6334,N_5704,N_5049);
nand U6335 (N_6335,N_5662,N_5115);
nand U6336 (N_6336,N_5951,N_4854);
xnor U6337 (N_6337,N_5487,N_4912);
nand U6338 (N_6338,N_5617,N_5824);
and U6339 (N_6339,N_4897,N_5966);
and U6340 (N_6340,N_4523,N_4814);
nor U6341 (N_6341,N_4966,N_5356);
xnor U6342 (N_6342,N_5585,N_5705);
nand U6343 (N_6343,N_4946,N_5176);
nor U6344 (N_6344,N_4981,N_4726);
and U6345 (N_6345,N_5492,N_5876);
and U6346 (N_6346,N_5847,N_4836);
or U6347 (N_6347,N_5985,N_4887);
or U6348 (N_6348,N_4647,N_5540);
or U6349 (N_6349,N_4510,N_5702);
and U6350 (N_6350,N_5976,N_4850);
nand U6351 (N_6351,N_5193,N_5320);
xor U6352 (N_6352,N_4848,N_5831);
and U6353 (N_6353,N_5222,N_5295);
nand U6354 (N_6354,N_5104,N_4567);
xor U6355 (N_6355,N_5605,N_5836);
and U6356 (N_6356,N_5622,N_5525);
nor U6357 (N_6357,N_5145,N_4628);
or U6358 (N_6358,N_4804,N_5628);
nor U6359 (N_6359,N_5107,N_5884);
or U6360 (N_6360,N_4512,N_4527);
or U6361 (N_6361,N_5221,N_5547);
nor U6362 (N_6362,N_5665,N_5680);
xor U6363 (N_6363,N_4744,N_5924);
xor U6364 (N_6364,N_5777,N_5242);
or U6365 (N_6365,N_5626,N_5047);
nand U6366 (N_6366,N_5548,N_5279);
or U6367 (N_6367,N_5488,N_5437);
or U6368 (N_6368,N_5389,N_5498);
or U6369 (N_6369,N_5522,N_5286);
xnor U6370 (N_6370,N_5515,N_5897);
or U6371 (N_6371,N_5546,N_4692);
xor U6372 (N_6372,N_5367,N_5888);
nor U6373 (N_6373,N_5770,N_5986);
nor U6374 (N_6374,N_5807,N_4520);
nand U6375 (N_6375,N_5086,N_5299);
nand U6376 (N_6376,N_5643,N_5615);
or U6377 (N_6377,N_5511,N_5402);
and U6378 (N_6378,N_4534,N_5041);
and U6379 (N_6379,N_5377,N_5902);
and U6380 (N_6380,N_5830,N_5707);
and U6381 (N_6381,N_4782,N_4879);
xnor U6382 (N_6382,N_5937,N_5591);
and U6383 (N_6383,N_4900,N_5963);
xor U6384 (N_6384,N_4613,N_4948);
or U6385 (N_6385,N_4767,N_5101);
nor U6386 (N_6386,N_4626,N_4673);
xnor U6387 (N_6387,N_4529,N_5791);
and U6388 (N_6388,N_4975,N_5291);
nor U6389 (N_6389,N_5802,N_5796);
or U6390 (N_6390,N_5113,N_5408);
or U6391 (N_6391,N_4674,N_5954);
and U6392 (N_6392,N_4577,N_5200);
and U6393 (N_6393,N_5701,N_5988);
or U6394 (N_6394,N_4568,N_5594);
or U6395 (N_6395,N_4676,N_5780);
nand U6396 (N_6396,N_4506,N_5732);
nand U6397 (N_6397,N_5092,N_4972);
nor U6398 (N_6398,N_5790,N_5866);
nand U6399 (N_6399,N_4745,N_5907);
nand U6400 (N_6400,N_4788,N_4592);
xnor U6401 (N_6401,N_4630,N_5703);
nand U6402 (N_6402,N_4922,N_5188);
nor U6403 (N_6403,N_5143,N_5280);
nor U6404 (N_6404,N_4650,N_5012);
nor U6405 (N_6405,N_5721,N_4987);
and U6406 (N_6406,N_5309,N_5822);
xor U6407 (N_6407,N_5410,N_5456);
xor U6408 (N_6408,N_4641,N_4779);
nor U6409 (N_6409,N_4677,N_5688);
nor U6410 (N_6410,N_5787,N_5563);
and U6411 (N_6411,N_4551,N_4697);
nor U6412 (N_6412,N_4585,N_5950);
nand U6413 (N_6413,N_5290,N_5684);
xor U6414 (N_6414,N_5283,N_5036);
xor U6415 (N_6415,N_4910,N_5204);
nor U6416 (N_6416,N_5895,N_5040);
or U6417 (N_6417,N_5355,N_4617);
and U6418 (N_6418,N_4877,N_5587);
xor U6419 (N_6419,N_5337,N_5412);
xnor U6420 (N_6420,N_4840,N_5433);
or U6421 (N_6421,N_5205,N_5485);
and U6422 (N_6422,N_4554,N_5491);
nand U6423 (N_6423,N_4925,N_5874);
nor U6424 (N_6424,N_5453,N_5244);
and U6425 (N_6425,N_5289,N_5285);
and U6426 (N_6426,N_5766,N_5121);
xnor U6427 (N_6427,N_5129,N_4913);
and U6428 (N_6428,N_4947,N_5133);
nor U6429 (N_6429,N_4816,N_5625);
or U6430 (N_6430,N_5495,N_4670);
nor U6431 (N_6431,N_5915,N_5679);
xnor U6432 (N_6432,N_5542,N_5435);
or U6433 (N_6433,N_5071,N_5644);
xnor U6434 (N_6434,N_5509,N_5060);
nand U6435 (N_6435,N_5551,N_5995);
or U6436 (N_6436,N_4970,N_5892);
nor U6437 (N_6437,N_4589,N_4828);
xor U6438 (N_6438,N_5788,N_5607);
nor U6439 (N_6439,N_5253,N_5817);
or U6440 (N_6440,N_5686,N_5858);
nand U6441 (N_6441,N_5354,N_5159);
xor U6442 (N_6442,N_5311,N_5282);
nor U6443 (N_6443,N_5850,N_5993);
xnor U6444 (N_6444,N_4711,N_5239);
and U6445 (N_6445,N_4802,N_5326);
nor U6446 (N_6446,N_5514,N_5228);
xnor U6447 (N_6447,N_5812,N_4736);
nor U6448 (N_6448,N_5479,N_4811);
xor U6449 (N_6449,N_4535,N_5177);
nand U6450 (N_6450,N_4852,N_5683);
nor U6451 (N_6451,N_5755,N_5868);
nand U6452 (N_6452,N_5851,N_5983);
and U6453 (N_6453,N_4797,N_5334);
xnor U6454 (N_6454,N_4622,N_5331);
nand U6455 (N_6455,N_5677,N_4998);
nor U6456 (N_6456,N_4883,N_5595);
xor U6457 (N_6457,N_5649,N_5973);
xor U6458 (N_6458,N_4552,N_4787);
nor U6459 (N_6459,N_4886,N_5657);
or U6460 (N_6460,N_4766,N_5371);
and U6461 (N_6461,N_5914,N_4821);
nor U6462 (N_6462,N_5761,N_5972);
and U6463 (N_6463,N_5004,N_5381);
nor U6464 (N_6464,N_5308,N_5002);
and U6465 (N_6465,N_5958,N_4757);
and U6466 (N_6466,N_5582,N_5146);
and U6467 (N_6467,N_5420,N_5725);
xor U6468 (N_6468,N_4809,N_4805);
and U6469 (N_6469,N_5210,N_5801);
and U6470 (N_6470,N_5179,N_5053);
or U6471 (N_6471,N_4599,N_5687);
or U6472 (N_6472,N_4812,N_5304);
nand U6473 (N_6473,N_4544,N_5424);
nand U6474 (N_6474,N_5928,N_5711);
and U6475 (N_6475,N_4819,N_5690);
xnor U6476 (N_6476,N_4537,N_5039);
or U6477 (N_6477,N_5608,N_4619);
or U6478 (N_6478,N_5610,N_5639);
or U6479 (N_6479,N_5618,N_4873);
or U6480 (N_6480,N_5742,N_4571);
nor U6481 (N_6481,N_4660,N_5726);
xnor U6482 (N_6482,N_5097,N_5619);
xnor U6483 (N_6483,N_5681,N_4796);
nand U6484 (N_6484,N_4899,N_4941);
or U6485 (N_6485,N_5059,N_5007);
or U6486 (N_6486,N_4586,N_5614);
and U6487 (N_6487,N_4857,N_5081);
nor U6488 (N_6488,N_5175,N_5991);
xnor U6489 (N_6489,N_4830,N_5481);
nand U6490 (N_6490,N_5918,N_5569);
nor U6491 (N_6491,N_4935,N_4707);
nor U6492 (N_6492,N_5358,N_5461);
and U6493 (N_6493,N_5971,N_5292);
and U6494 (N_6494,N_5675,N_5627);
and U6495 (N_6495,N_4730,N_5395);
xor U6496 (N_6496,N_4573,N_5130);
nor U6497 (N_6497,N_5267,N_5296);
nand U6498 (N_6498,N_5864,N_5019);
nand U6499 (N_6499,N_4827,N_5471);
or U6500 (N_6500,N_5932,N_5962);
and U6501 (N_6501,N_4590,N_4771);
xnor U6502 (N_6502,N_4996,N_5301);
or U6503 (N_6503,N_5393,N_5340);
xnor U6504 (N_6504,N_5136,N_5837);
xor U6505 (N_6505,N_5374,N_5091);
and U6506 (N_6506,N_4786,N_5570);
nand U6507 (N_6507,N_5241,N_5223);
xnor U6508 (N_6508,N_4949,N_5262);
nor U6509 (N_6509,N_5541,N_4882);
and U6510 (N_6510,N_4621,N_4952);
and U6511 (N_6511,N_5946,N_5957);
nor U6512 (N_6512,N_5877,N_4936);
nand U6513 (N_6513,N_5165,N_5126);
nand U6514 (N_6514,N_5779,N_4776);
or U6515 (N_6515,N_5724,N_5609);
or U6516 (N_6516,N_5008,N_4625);
nor U6517 (N_6517,N_5298,N_5465);
xnor U6518 (N_6518,N_4678,N_4760);
nor U6519 (N_6519,N_5095,N_4665);
nand U6520 (N_6520,N_5862,N_4614);
or U6521 (N_6521,N_5364,N_5834);
nand U6522 (N_6522,N_4675,N_5249);
nand U6523 (N_6523,N_5430,N_5624);
nand U6524 (N_6524,N_4559,N_5106);
nor U6525 (N_6525,N_4871,N_5284);
xor U6526 (N_6526,N_5135,N_5429);
xor U6527 (N_6527,N_5313,N_4743);
and U6528 (N_6528,N_5327,N_5723);
xnor U6529 (N_6529,N_5182,N_5912);
or U6530 (N_6530,N_5131,N_5881);
xnor U6531 (N_6531,N_5056,N_5475);
nand U6532 (N_6532,N_5545,N_5254);
nand U6533 (N_6533,N_5110,N_5583);
or U6534 (N_6534,N_4729,N_5968);
xnor U6535 (N_6535,N_4822,N_4664);
nand U6536 (N_6536,N_5667,N_4694);
nand U6537 (N_6537,N_5303,N_5816);
xnor U6538 (N_6538,N_4826,N_5561);
xnor U6539 (N_6539,N_5046,N_5074);
xor U6540 (N_6540,N_5948,N_5003);
nand U6541 (N_6541,N_5611,N_5853);
nand U6542 (N_6542,N_5856,N_5068);
nor U6543 (N_6543,N_5388,N_5058);
nor U6544 (N_6544,N_5218,N_4884);
nand U6545 (N_6545,N_4774,N_4563);
xor U6546 (N_6546,N_5658,N_5910);
xor U6547 (N_6547,N_5150,N_4654);
or U6548 (N_6548,N_5575,N_4945);
xnor U6549 (N_6549,N_5661,N_4896);
xor U6550 (N_6550,N_5606,N_4930);
or U6551 (N_6551,N_5066,N_4944);
xnor U6552 (N_6552,N_4624,N_4754);
nor U6553 (N_6553,N_5828,N_5623);
or U6554 (N_6554,N_5421,N_4639);
nor U6555 (N_6555,N_5192,N_4533);
nand U6556 (N_6556,N_5752,N_4865);
xnor U6557 (N_6557,N_5431,N_5098);
xnor U6558 (N_6558,N_4646,N_5170);
xnor U6559 (N_6559,N_5297,N_5321);
xor U6560 (N_6560,N_5792,N_4777);
or U6561 (N_6561,N_5382,N_4901);
nor U6562 (N_6562,N_5369,N_4562);
nor U6563 (N_6563,N_5341,N_5769);
nor U6564 (N_6564,N_4618,N_5401);
and U6565 (N_6565,N_5076,N_4911);
xor U6566 (N_6566,N_5357,N_5268);
nand U6567 (N_6567,N_5276,N_5483);
xor U6568 (N_6568,N_4543,N_5841);
nor U6569 (N_6569,N_5689,N_5307);
or U6570 (N_6570,N_5314,N_5443);
nor U6571 (N_6571,N_4963,N_4761);
nor U6572 (N_6572,N_4878,N_5018);
and U6573 (N_6573,N_4999,N_4906);
or U6574 (N_6574,N_5889,N_5100);
nor U6575 (N_6575,N_5398,N_5906);
nor U6576 (N_6576,N_5713,N_5272);
nor U6577 (N_6577,N_5600,N_4902);
xor U6578 (N_6578,N_4689,N_4853);
nor U6579 (N_6579,N_5987,N_4929);
nor U6580 (N_6580,N_5682,N_5581);
or U6581 (N_6581,N_5749,N_4803);
nor U6582 (N_6582,N_5693,N_5730);
and U6583 (N_6583,N_4977,N_5746);
and U6584 (N_6584,N_4733,N_5543);
xnor U6585 (N_6585,N_5413,N_4974);
nor U6586 (N_6586,N_5454,N_4652);
nor U6587 (N_6587,N_4663,N_5839);
nor U6588 (N_6588,N_4632,N_4923);
nand U6589 (N_6589,N_5353,N_4765);
and U6590 (N_6590,N_4829,N_4909);
or U6591 (N_6591,N_5141,N_5556);
or U6592 (N_6592,N_4781,N_5981);
nor U6593 (N_6593,N_5031,N_5640);
nand U6594 (N_6594,N_4749,N_4868);
nor U6595 (N_6595,N_4968,N_5678);
nor U6596 (N_6596,N_5997,N_4684);
or U6597 (N_6597,N_4575,N_4755);
nor U6598 (N_6598,N_5741,N_5577);
and U6599 (N_6599,N_5908,N_4954);
xor U6600 (N_6600,N_4558,N_5166);
and U6601 (N_6601,N_5459,N_5941);
and U6602 (N_6602,N_5375,N_5466);
nand U6603 (N_6603,N_5786,N_5671);
or U6604 (N_6604,N_5099,N_4764);
xor U6605 (N_6605,N_5645,N_5999);
nor U6606 (N_6606,N_5553,N_5826);
xnor U6607 (N_6607,N_5722,N_5633);
nand U6608 (N_6608,N_5524,N_5526);
nor U6609 (N_6609,N_5484,N_4509);
or U6610 (N_6610,N_5209,N_5927);
nor U6611 (N_6611,N_5198,N_5535);
xnor U6612 (N_6612,N_5589,N_5940);
or U6613 (N_6613,N_4994,N_4546);
or U6614 (N_6614,N_5082,N_5904);
xor U6615 (N_6615,N_4815,N_5124);
and U6616 (N_6616,N_5886,N_5370);
or U6617 (N_6617,N_5774,N_5194);
and U6618 (N_6618,N_5015,N_5407);
or U6619 (N_6619,N_5022,N_4937);
or U6620 (N_6620,N_5164,N_5251);
nor U6621 (N_6621,N_5775,N_4679);
xor U6622 (N_6622,N_4610,N_5342);
nand U6623 (N_6623,N_5539,N_5768);
nor U6624 (N_6624,N_5753,N_5347);
or U6625 (N_6625,N_4741,N_4598);
xor U6626 (N_6626,N_5468,N_5001);
and U6627 (N_6627,N_5654,N_5152);
nand U6628 (N_6628,N_5781,N_5676);
nor U6629 (N_6629,N_5148,N_5451);
nor U6630 (N_6630,N_5275,N_5764);
nand U6631 (N_6631,N_5922,N_4699);
nor U6632 (N_6632,N_5773,N_5206);
nand U6633 (N_6633,N_5977,N_5197);
or U6634 (N_6634,N_5549,N_5464);
nand U6635 (N_6635,N_5602,N_5804);
nand U6636 (N_6636,N_5387,N_5694);
or U6637 (N_6637,N_5083,N_4666);
nor U6638 (N_6638,N_4837,N_5650);
nand U6639 (N_6639,N_5028,N_4623);
nor U6640 (N_6640,N_4753,N_5042);
nand U6641 (N_6641,N_5878,N_5048);
xor U6642 (N_6642,N_5848,N_5994);
nand U6643 (N_6643,N_5593,N_5905);
xor U6644 (N_6644,N_5343,N_5363);
or U6645 (N_6645,N_4919,N_4612);
xor U6646 (N_6646,N_5933,N_4683);
nor U6647 (N_6647,N_4888,N_5935);
xor U6648 (N_6648,N_5138,N_5189);
nor U6649 (N_6649,N_4649,N_4507);
nand U6650 (N_6650,N_4982,N_4832);
nand U6651 (N_6651,N_4631,N_5416);
or U6652 (N_6652,N_5452,N_5508);
xnor U6653 (N_6653,N_5990,N_5384);
nand U6654 (N_6654,N_4662,N_4864);
or U6655 (N_6655,N_5441,N_5302);
or U6656 (N_6656,N_4855,N_5024);
and U6657 (N_6657,N_5512,N_4799);
and U6658 (N_6658,N_5576,N_4591);
xnor U6659 (N_6659,N_4750,N_5784);
nor U6660 (N_6660,N_5385,N_5505);
nor U6661 (N_6661,N_4604,N_5673);
or U6662 (N_6662,N_5637,N_5030);
nor U6663 (N_6663,N_5238,N_5521);
nor U6664 (N_6664,N_5854,N_4671);
nand U6665 (N_6665,N_5803,N_5409);
or U6666 (N_6666,N_5366,N_4693);
nand U6667 (N_6667,N_5745,N_4845);
and U6668 (N_6668,N_5819,N_5944);
or U6669 (N_6669,N_5736,N_5975);
nand U6670 (N_6670,N_5084,N_5411);
xnor U6671 (N_6671,N_5580,N_5793);
nor U6672 (N_6672,N_5467,N_5536);
and U6673 (N_6673,N_5477,N_4768);
nor U6674 (N_6674,N_5718,N_4656);
and U6675 (N_6675,N_5759,N_5245);
and U6676 (N_6676,N_5744,N_5697);
nand U6677 (N_6677,N_4616,N_5050);
or U6678 (N_6678,N_4681,N_5631);
nor U6679 (N_6679,N_4713,N_5783);
or U6680 (N_6680,N_5418,N_5075);
nor U6681 (N_6681,N_5552,N_5011);
or U6682 (N_6682,N_4793,N_4724);
or U6683 (N_6683,N_4928,N_5203);
nor U6684 (N_6684,N_4775,N_4933);
nand U6685 (N_6685,N_5310,N_5829);
nand U6686 (N_6686,N_5400,N_5636);
xor U6687 (N_6687,N_5263,N_5500);
and U6688 (N_6688,N_5719,N_5849);
nand U6689 (N_6689,N_5422,N_5698);
and U6690 (N_6690,N_5598,N_5647);
and U6691 (N_6691,N_5323,N_5629);
xnor U6692 (N_6692,N_5073,N_5109);
or U6693 (N_6693,N_5765,N_4522);
nor U6694 (N_6694,N_5070,N_4582);
nor U6695 (N_6695,N_5139,N_4721);
xnor U6696 (N_6696,N_5747,N_5330);
and U6697 (N_6697,N_4920,N_5037);
nor U6698 (N_6698,N_5756,N_5867);
and U6699 (N_6699,N_4500,N_4839);
nand U6700 (N_6700,N_5208,N_5093);
or U6701 (N_6701,N_5379,N_5269);
or U6702 (N_6702,N_5233,N_4690);
and U6703 (N_6703,N_4867,N_5811);
nand U6704 (N_6704,N_5913,N_5887);
xor U6705 (N_6705,N_5771,N_4813);
nor U6706 (N_6706,N_5832,N_5560);
nand U6707 (N_6707,N_4719,N_5925);
or U6708 (N_6708,N_5691,N_4958);
xnor U6709 (N_6709,N_5174,N_5202);
xor U6710 (N_6710,N_5094,N_4657);
nand U6711 (N_6711,N_5555,N_5737);
nor U6712 (N_6712,N_4732,N_5144);
or U6713 (N_6713,N_4874,N_4785);
xor U6714 (N_6714,N_5664,N_4898);
nand U6715 (N_6715,N_4783,N_4620);
nor U6716 (N_6716,N_5604,N_4824);
xor U6717 (N_6717,N_5446,N_5708);
and U6718 (N_6718,N_4751,N_5470);
nor U6719 (N_6719,N_5108,N_4980);
xnor U6720 (N_6720,N_5322,N_4576);
xnor U6721 (N_6721,N_5890,N_5372);
nand U6722 (N_6722,N_4702,N_5530);
xnor U6723 (N_6723,N_5052,N_5346);
xnor U6724 (N_6724,N_5870,N_5982);
nand U6725 (N_6725,N_5062,N_4643);
and U6726 (N_6726,N_5641,N_5871);
nor U6727 (N_6727,N_5668,N_4806);
xor U6728 (N_6728,N_4555,N_5154);
xnor U6729 (N_6729,N_5554,N_4595);
nor U6730 (N_6730,N_5716,N_5706);
and U6731 (N_6731,N_5480,N_5448);
xnor U6732 (N_6732,N_5180,N_5211);
and U6733 (N_6733,N_4962,N_4634);
nor U6734 (N_6734,N_5476,N_4993);
nand U6735 (N_6735,N_4651,N_4739);
xnor U6736 (N_6736,N_5883,N_5163);
nor U6737 (N_6737,N_5572,N_5006);
nand U6738 (N_6738,N_5266,N_5065);
nor U6739 (N_6739,N_4615,N_5489);
nand U6740 (N_6740,N_5519,N_5077);
nor U6741 (N_6741,N_5156,N_4921);
or U6742 (N_6742,N_4893,N_5499);
nor U6743 (N_6743,N_5236,N_5474);
xor U6744 (N_6744,N_5426,N_4798);
or U6745 (N_6745,N_4550,N_5840);
nand U6746 (N_6746,N_5538,N_5439);
nand U6747 (N_6747,N_4538,N_5818);
xor U6748 (N_6748,N_5063,N_4695);
and U6749 (N_6749,N_4843,N_4859);
and U6750 (N_6750,N_5098,N_5169);
and U6751 (N_6751,N_4642,N_5792);
nor U6752 (N_6752,N_4612,N_4724);
nor U6753 (N_6753,N_4872,N_5333);
nor U6754 (N_6754,N_4580,N_5364);
xor U6755 (N_6755,N_4972,N_5658);
nor U6756 (N_6756,N_5454,N_4729);
nor U6757 (N_6757,N_5305,N_4741);
or U6758 (N_6758,N_4915,N_5141);
and U6759 (N_6759,N_5023,N_5076);
and U6760 (N_6760,N_4521,N_4520);
and U6761 (N_6761,N_5840,N_5235);
and U6762 (N_6762,N_5879,N_5887);
or U6763 (N_6763,N_5091,N_4578);
or U6764 (N_6764,N_5542,N_4649);
nand U6765 (N_6765,N_5595,N_5130);
or U6766 (N_6766,N_5018,N_5035);
xor U6767 (N_6767,N_4517,N_4910);
or U6768 (N_6768,N_4825,N_5052);
xnor U6769 (N_6769,N_4907,N_5809);
xor U6770 (N_6770,N_4971,N_5307);
xor U6771 (N_6771,N_4832,N_4895);
nor U6772 (N_6772,N_5171,N_4666);
or U6773 (N_6773,N_5607,N_5680);
nor U6774 (N_6774,N_4650,N_5812);
and U6775 (N_6775,N_4740,N_5373);
nand U6776 (N_6776,N_5091,N_5693);
nor U6777 (N_6777,N_5010,N_5355);
or U6778 (N_6778,N_5735,N_5482);
xnor U6779 (N_6779,N_4519,N_5261);
nand U6780 (N_6780,N_5613,N_5049);
xor U6781 (N_6781,N_5338,N_5539);
nor U6782 (N_6782,N_5961,N_5610);
and U6783 (N_6783,N_4880,N_5615);
xnor U6784 (N_6784,N_5167,N_5393);
or U6785 (N_6785,N_5985,N_5548);
nand U6786 (N_6786,N_5635,N_5415);
nor U6787 (N_6787,N_5208,N_5505);
nand U6788 (N_6788,N_5760,N_5481);
nand U6789 (N_6789,N_4959,N_5604);
xnor U6790 (N_6790,N_5964,N_4565);
nand U6791 (N_6791,N_4567,N_5568);
nor U6792 (N_6792,N_5433,N_4985);
and U6793 (N_6793,N_4750,N_5567);
nor U6794 (N_6794,N_4619,N_5398);
or U6795 (N_6795,N_4886,N_5602);
or U6796 (N_6796,N_5998,N_4737);
or U6797 (N_6797,N_5772,N_5810);
nand U6798 (N_6798,N_4582,N_5556);
xnor U6799 (N_6799,N_4666,N_5666);
xnor U6800 (N_6800,N_5932,N_5816);
nand U6801 (N_6801,N_5267,N_5487);
nand U6802 (N_6802,N_5875,N_4558);
or U6803 (N_6803,N_5693,N_5980);
nor U6804 (N_6804,N_4891,N_4938);
nor U6805 (N_6805,N_5387,N_4853);
or U6806 (N_6806,N_5377,N_5665);
xnor U6807 (N_6807,N_4762,N_5337);
nor U6808 (N_6808,N_5521,N_5638);
xor U6809 (N_6809,N_4844,N_4749);
xnor U6810 (N_6810,N_4822,N_5335);
or U6811 (N_6811,N_4642,N_4864);
xor U6812 (N_6812,N_5425,N_4851);
or U6813 (N_6813,N_5127,N_5499);
xnor U6814 (N_6814,N_4678,N_4503);
nand U6815 (N_6815,N_5297,N_4566);
and U6816 (N_6816,N_5604,N_4854);
and U6817 (N_6817,N_5741,N_5452);
xor U6818 (N_6818,N_4701,N_5707);
xnor U6819 (N_6819,N_5818,N_5000);
xor U6820 (N_6820,N_5858,N_5492);
nand U6821 (N_6821,N_4817,N_4889);
and U6822 (N_6822,N_5191,N_5517);
nand U6823 (N_6823,N_5124,N_5377);
or U6824 (N_6824,N_5601,N_4683);
nor U6825 (N_6825,N_4783,N_4755);
and U6826 (N_6826,N_4552,N_5716);
xnor U6827 (N_6827,N_5926,N_4827);
nor U6828 (N_6828,N_4775,N_5658);
and U6829 (N_6829,N_5184,N_5514);
nand U6830 (N_6830,N_4678,N_5342);
xnor U6831 (N_6831,N_5882,N_5036);
nor U6832 (N_6832,N_4875,N_4954);
or U6833 (N_6833,N_4683,N_4702);
nand U6834 (N_6834,N_5399,N_5383);
xnor U6835 (N_6835,N_4985,N_5030);
nor U6836 (N_6836,N_5375,N_5656);
or U6837 (N_6837,N_5181,N_5964);
or U6838 (N_6838,N_4592,N_5179);
nand U6839 (N_6839,N_4844,N_5574);
and U6840 (N_6840,N_4615,N_5143);
or U6841 (N_6841,N_5458,N_4691);
and U6842 (N_6842,N_5620,N_5106);
or U6843 (N_6843,N_5323,N_5461);
xor U6844 (N_6844,N_5624,N_5587);
xnor U6845 (N_6845,N_4612,N_4833);
and U6846 (N_6846,N_5272,N_4848);
or U6847 (N_6847,N_5433,N_5220);
or U6848 (N_6848,N_4717,N_4698);
or U6849 (N_6849,N_4634,N_5090);
and U6850 (N_6850,N_5661,N_5149);
nor U6851 (N_6851,N_4633,N_4575);
nand U6852 (N_6852,N_5602,N_5692);
or U6853 (N_6853,N_5141,N_5924);
nor U6854 (N_6854,N_5232,N_4997);
nand U6855 (N_6855,N_5394,N_4559);
and U6856 (N_6856,N_5205,N_4606);
nand U6857 (N_6857,N_5903,N_5068);
nand U6858 (N_6858,N_5018,N_5583);
nand U6859 (N_6859,N_4661,N_5293);
xnor U6860 (N_6860,N_5051,N_5219);
xor U6861 (N_6861,N_4629,N_5191);
or U6862 (N_6862,N_5914,N_4502);
or U6863 (N_6863,N_5957,N_5611);
nand U6864 (N_6864,N_4579,N_5007);
nand U6865 (N_6865,N_5064,N_5052);
xor U6866 (N_6866,N_5395,N_5205);
xor U6867 (N_6867,N_5111,N_5626);
nand U6868 (N_6868,N_5530,N_4781);
and U6869 (N_6869,N_4986,N_4946);
and U6870 (N_6870,N_5299,N_4666);
xor U6871 (N_6871,N_5107,N_5938);
xor U6872 (N_6872,N_5918,N_4589);
and U6873 (N_6873,N_5732,N_5340);
nor U6874 (N_6874,N_5834,N_5344);
nand U6875 (N_6875,N_4726,N_5478);
nor U6876 (N_6876,N_5290,N_5789);
and U6877 (N_6877,N_5992,N_5550);
nor U6878 (N_6878,N_5866,N_5955);
nor U6879 (N_6879,N_5345,N_5405);
and U6880 (N_6880,N_5898,N_5576);
xor U6881 (N_6881,N_4902,N_4539);
nor U6882 (N_6882,N_5628,N_5309);
xor U6883 (N_6883,N_5044,N_5220);
or U6884 (N_6884,N_4957,N_5914);
xnor U6885 (N_6885,N_5274,N_4988);
and U6886 (N_6886,N_5313,N_4738);
nor U6887 (N_6887,N_5204,N_5742);
nand U6888 (N_6888,N_5009,N_4726);
nand U6889 (N_6889,N_4535,N_4664);
and U6890 (N_6890,N_5149,N_5850);
nand U6891 (N_6891,N_4766,N_4969);
nand U6892 (N_6892,N_5795,N_5562);
or U6893 (N_6893,N_5274,N_4516);
nand U6894 (N_6894,N_5664,N_5397);
xnor U6895 (N_6895,N_5248,N_5940);
xor U6896 (N_6896,N_5879,N_4732);
nor U6897 (N_6897,N_4587,N_5331);
nor U6898 (N_6898,N_4933,N_4904);
and U6899 (N_6899,N_4949,N_5646);
nor U6900 (N_6900,N_5620,N_5121);
xor U6901 (N_6901,N_5546,N_4793);
or U6902 (N_6902,N_5710,N_5065);
nand U6903 (N_6903,N_4758,N_5477);
nor U6904 (N_6904,N_5655,N_4556);
and U6905 (N_6905,N_5210,N_4896);
nor U6906 (N_6906,N_5635,N_4941);
and U6907 (N_6907,N_5603,N_5581);
or U6908 (N_6908,N_4857,N_4961);
nand U6909 (N_6909,N_5052,N_5697);
nand U6910 (N_6910,N_4571,N_5434);
or U6911 (N_6911,N_5619,N_5472);
nand U6912 (N_6912,N_5726,N_4534);
xor U6913 (N_6913,N_4719,N_5995);
or U6914 (N_6914,N_4631,N_5709);
nor U6915 (N_6915,N_5546,N_5200);
and U6916 (N_6916,N_5128,N_5022);
and U6917 (N_6917,N_5176,N_4967);
and U6918 (N_6918,N_5903,N_5753);
or U6919 (N_6919,N_5188,N_4871);
xor U6920 (N_6920,N_4769,N_5096);
and U6921 (N_6921,N_4578,N_5667);
xnor U6922 (N_6922,N_5307,N_5346);
nand U6923 (N_6923,N_5561,N_4626);
and U6924 (N_6924,N_4659,N_4709);
xor U6925 (N_6925,N_4784,N_5812);
nor U6926 (N_6926,N_5870,N_5257);
nand U6927 (N_6927,N_4580,N_4908);
and U6928 (N_6928,N_4642,N_5302);
xor U6929 (N_6929,N_4689,N_4717);
xnor U6930 (N_6930,N_4633,N_5664);
xnor U6931 (N_6931,N_4564,N_5187);
and U6932 (N_6932,N_4519,N_5129);
or U6933 (N_6933,N_5952,N_5245);
and U6934 (N_6934,N_5252,N_5042);
xnor U6935 (N_6935,N_4823,N_5720);
or U6936 (N_6936,N_4781,N_4893);
and U6937 (N_6937,N_5616,N_5838);
and U6938 (N_6938,N_4559,N_5880);
nor U6939 (N_6939,N_4974,N_5851);
nor U6940 (N_6940,N_4834,N_5310);
and U6941 (N_6941,N_5107,N_5709);
nand U6942 (N_6942,N_4563,N_4752);
or U6943 (N_6943,N_4912,N_5960);
nand U6944 (N_6944,N_5352,N_4651);
nand U6945 (N_6945,N_5572,N_4632);
and U6946 (N_6946,N_5031,N_5725);
nand U6947 (N_6947,N_5641,N_5663);
xor U6948 (N_6948,N_5997,N_5236);
or U6949 (N_6949,N_5616,N_5844);
xnor U6950 (N_6950,N_5995,N_5531);
nor U6951 (N_6951,N_5832,N_5704);
xnor U6952 (N_6952,N_4849,N_4735);
or U6953 (N_6953,N_5432,N_5365);
xnor U6954 (N_6954,N_5313,N_4763);
and U6955 (N_6955,N_5696,N_4842);
nor U6956 (N_6956,N_4737,N_5823);
xnor U6957 (N_6957,N_5067,N_5237);
nand U6958 (N_6958,N_5728,N_5017);
nor U6959 (N_6959,N_5274,N_5278);
or U6960 (N_6960,N_5087,N_5109);
nor U6961 (N_6961,N_5353,N_4927);
nand U6962 (N_6962,N_5573,N_5306);
nand U6963 (N_6963,N_5165,N_5743);
xnor U6964 (N_6964,N_5486,N_5567);
nand U6965 (N_6965,N_5161,N_5164);
xor U6966 (N_6966,N_5346,N_5083);
nor U6967 (N_6967,N_4558,N_5550);
nor U6968 (N_6968,N_5337,N_5332);
xor U6969 (N_6969,N_5262,N_4996);
xor U6970 (N_6970,N_5350,N_5930);
and U6971 (N_6971,N_5315,N_4602);
nand U6972 (N_6972,N_5804,N_5302);
xnor U6973 (N_6973,N_4924,N_4597);
and U6974 (N_6974,N_5490,N_5257);
and U6975 (N_6975,N_4547,N_5234);
nor U6976 (N_6976,N_4601,N_5432);
nand U6977 (N_6977,N_5495,N_5238);
nand U6978 (N_6978,N_5995,N_5802);
nor U6979 (N_6979,N_5745,N_5395);
or U6980 (N_6980,N_5204,N_5503);
nor U6981 (N_6981,N_5253,N_5600);
nor U6982 (N_6982,N_5109,N_5640);
and U6983 (N_6983,N_5038,N_5547);
nor U6984 (N_6984,N_4995,N_5091);
and U6985 (N_6985,N_5561,N_4678);
and U6986 (N_6986,N_5846,N_5640);
or U6987 (N_6987,N_4512,N_5806);
xor U6988 (N_6988,N_4655,N_5258);
nand U6989 (N_6989,N_5393,N_5501);
or U6990 (N_6990,N_4801,N_4974);
nor U6991 (N_6991,N_4731,N_5331);
nand U6992 (N_6992,N_5440,N_4711);
nand U6993 (N_6993,N_4592,N_5343);
and U6994 (N_6994,N_5391,N_4506);
and U6995 (N_6995,N_5476,N_5767);
nand U6996 (N_6996,N_5715,N_5689);
or U6997 (N_6997,N_4523,N_5408);
nand U6998 (N_6998,N_4792,N_5969);
nand U6999 (N_6999,N_4735,N_4966);
and U7000 (N_7000,N_5031,N_5332);
nor U7001 (N_7001,N_5435,N_5507);
nand U7002 (N_7002,N_5543,N_5911);
and U7003 (N_7003,N_5049,N_5054);
nor U7004 (N_7004,N_4504,N_5625);
xor U7005 (N_7005,N_5863,N_5578);
and U7006 (N_7006,N_4861,N_5088);
xnor U7007 (N_7007,N_5376,N_5830);
nand U7008 (N_7008,N_5256,N_5365);
or U7009 (N_7009,N_5565,N_4948);
xor U7010 (N_7010,N_5015,N_5005);
nor U7011 (N_7011,N_4663,N_5761);
nor U7012 (N_7012,N_5517,N_4740);
nand U7013 (N_7013,N_4883,N_4586);
or U7014 (N_7014,N_5011,N_4557);
nor U7015 (N_7015,N_5105,N_5507);
and U7016 (N_7016,N_5272,N_4646);
xor U7017 (N_7017,N_5318,N_5847);
and U7018 (N_7018,N_4640,N_5609);
and U7019 (N_7019,N_5871,N_5318);
and U7020 (N_7020,N_4676,N_4627);
and U7021 (N_7021,N_5006,N_5260);
or U7022 (N_7022,N_5941,N_5575);
xor U7023 (N_7023,N_5317,N_5194);
nor U7024 (N_7024,N_5054,N_4801);
or U7025 (N_7025,N_5493,N_5194);
nand U7026 (N_7026,N_5103,N_4895);
and U7027 (N_7027,N_4811,N_4748);
and U7028 (N_7028,N_5775,N_4501);
xnor U7029 (N_7029,N_5277,N_4738);
and U7030 (N_7030,N_5980,N_4703);
and U7031 (N_7031,N_5225,N_5009);
nand U7032 (N_7032,N_5690,N_5246);
or U7033 (N_7033,N_5580,N_4578);
and U7034 (N_7034,N_5887,N_5310);
nand U7035 (N_7035,N_5291,N_4534);
and U7036 (N_7036,N_5001,N_5800);
nor U7037 (N_7037,N_4999,N_4814);
or U7038 (N_7038,N_5702,N_4502);
nor U7039 (N_7039,N_4651,N_4594);
nor U7040 (N_7040,N_4666,N_5121);
nor U7041 (N_7041,N_4573,N_5304);
nor U7042 (N_7042,N_4623,N_4996);
and U7043 (N_7043,N_5934,N_4845);
xor U7044 (N_7044,N_5061,N_4850);
nor U7045 (N_7045,N_4724,N_5566);
nand U7046 (N_7046,N_5291,N_5838);
xor U7047 (N_7047,N_4842,N_4975);
nand U7048 (N_7048,N_4539,N_5469);
nand U7049 (N_7049,N_5745,N_4821);
and U7050 (N_7050,N_4514,N_5252);
or U7051 (N_7051,N_5268,N_5231);
or U7052 (N_7052,N_5016,N_4943);
nand U7053 (N_7053,N_4955,N_5599);
nand U7054 (N_7054,N_5911,N_4891);
nand U7055 (N_7055,N_4791,N_5059);
or U7056 (N_7056,N_4514,N_5189);
or U7057 (N_7057,N_5608,N_5258);
and U7058 (N_7058,N_4668,N_4625);
and U7059 (N_7059,N_5618,N_5095);
nand U7060 (N_7060,N_5823,N_4569);
and U7061 (N_7061,N_5564,N_4691);
nand U7062 (N_7062,N_5896,N_5003);
xnor U7063 (N_7063,N_4947,N_4568);
nor U7064 (N_7064,N_5802,N_5159);
nor U7065 (N_7065,N_5420,N_4679);
or U7066 (N_7066,N_5271,N_5289);
nand U7067 (N_7067,N_4651,N_5707);
and U7068 (N_7068,N_5526,N_5081);
nor U7069 (N_7069,N_5800,N_5671);
nor U7070 (N_7070,N_5466,N_5750);
nor U7071 (N_7071,N_5192,N_5924);
or U7072 (N_7072,N_4826,N_5847);
nor U7073 (N_7073,N_4774,N_4619);
xor U7074 (N_7074,N_5718,N_5791);
nand U7075 (N_7075,N_5367,N_5759);
xor U7076 (N_7076,N_5761,N_4595);
or U7077 (N_7077,N_5680,N_4826);
nand U7078 (N_7078,N_4903,N_5333);
nand U7079 (N_7079,N_5726,N_4683);
nor U7080 (N_7080,N_5032,N_5991);
nor U7081 (N_7081,N_4610,N_4738);
or U7082 (N_7082,N_4641,N_5908);
nor U7083 (N_7083,N_5277,N_5264);
xnor U7084 (N_7084,N_5610,N_4865);
xor U7085 (N_7085,N_4792,N_4590);
and U7086 (N_7086,N_5546,N_4745);
xnor U7087 (N_7087,N_5536,N_4576);
and U7088 (N_7088,N_5657,N_4910);
xnor U7089 (N_7089,N_5898,N_5878);
nor U7090 (N_7090,N_5086,N_5985);
or U7091 (N_7091,N_5745,N_5998);
nand U7092 (N_7092,N_4730,N_5620);
xor U7093 (N_7093,N_5384,N_4633);
nor U7094 (N_7094,N_4639,N_5030);
nor U7095 (N_7095,N_5327,N_4762);
nand U7096 (N_7096,N_4833,N_5450);
nand U7097 (N_7097,N_5467,N_5542);
nand U7098 (N_7098,N_5706,N_5248);
and U7099 (N_7099,N_5026,N_5374);
xnor U7100 (N_7100,N_4958,N_5721);
xor U7101 (N_7101,N_5389,N_5897);
or U7102 (N_7102,N_5478,N_5743);
and U7103 (N_7103,N_5082,N_4674);
nand U7104 (N_7104,N_4827,N_4999);
or U7105 (N_7105,N_4702,N_5055);
and U7106 (N_7106,N_4993,N_5664);
nand U7107 (N_7107,N_5404,N_5769);
xnor U7108 (N_7108,N_4704,N_4985);
xnor U7109 (N_7109,N_4507,N_5586);
or U7110 (N_7110,N_5481,N_5994);
or U7111 (N_7111,N_4665,N_5011);
xor U7112 (N_7112,N_5749,N_4726);
or U7113 (N_7113,N_5294,N_4794);
and U7114 (N_7114,N_5037,N_5495);
or U7115 (N_7115,N_4812,N_4850);
nor U7116 (N_7116,N_5617,N_4710);
and U7117 (N_7117,N_5822,N_5002);
nor U7118 (N_7118,N_5806,N_5067);
or U7119 (N_7119,N_5078,N_5145);
nand U7120 (N_7120,N_5301,N_5574);
or U7121 (N_7121,N_5005,N_5459);
nor U7122 (N_7122,N_5126,N_4613);
xor U7123 (N_7123,N_5109,N_4943);
xnor U7124 (N_7124,N_4755,N_5676);
and U7125 (N_7125,N_5561,N_5807);
or U7126 (N_7126,N_5887,N_5177);
xor U7127 (N_7127,N_5921,N_4742);
xnor U7128 (N_7128,N_4672,N_5419);
xor U7129 (N_7129,N_5634,N_5093);
nand U7130 (N_7130,N_5740,N_5388);
nand U7131 (N_7131,N_5275,N_4826);
and U7132 (N_7132,N_5490,N_5856);
nand U7133 (N_7133,N_4826,N_5408);
nor U7134 (N_7134,N_4999,N_5612);
and U7135 (N_7135,N_5140,N_4634);
xnor U7136 (N_7136,N_4774,N_5432);
nand U7137 (N_7137,N_5716,N_5748);
nand U7138 (N_7138,N_5481,N_5110);
and U7139 (N_7139,N_5205,N_5257);
or U7140 (N_7140,N_5021,N_4854);
nor U7141 (N_7141,N_5266,N_5725);
nor U7142 (N_7142,N_5680,N_4522);
nor U7143 (N_7143,N_5370,N_5216);
or U7144 (N_7144,N_5806,N_4830);
or U7145 (N_7145,N_4885,N_5714);
or U7146 (N_7146,N_4975,N_5533);
nor U7147 (N_7147,N_4868,N_5896);
or U7148 (N_7148,N_5120,N_4921);
and U7149 (N_7149,N_4856,N_5864);
nand U7150 (N_7150,N_5047,N_5226);
xnor U7151 (N_7151,N_5145,N_5646);
nand U7152 (N_7152,N_5856,N_5315);
nor U7153 (N_7153,N_5669,N_5236);
nor U7154 (N_7154,N_5269,N_5024);
nor U7155 (N_7155,N_5838,N_5223);
or U7156 (N_7156,N_4682,N_5229);
or U7157 (N_7157,N_5283,N_5860);
nand U7158 (N_7158,N_5875,N_5283);
nor U7159 (N_7159,N_5407,N_4702);
nor U7160 (N_7160,N_4856,N_5481);
nand U7161 (N_7161,N_5645,N_4941);
nand U7162 (N_7162,N_5137,N_5066);
and U7163 (N_7163,N_4764,N_5996);
xor U7164 (N_7164,N_5331,N_5466);
and U7165 (N_7165,N_5790,N_5960);
or U7166 (N_7166,N_5876,N_5841);
and U7167 (N_7167,N_5687,N_5216);
nor U7168 (N_7168,N_5457,N_5048);
nand U7169 (N_7169,N_5421,N_5287);
nor U7170 (N_7170,N_5401,N_5962);
or U7171 (N_7171,N_4882,N_5072);
nor U7172 (N_7172,N_5014,N_5677);
or U7173 (N_7173,N_5559,N_5385);
nor U7174 (N_7174,N_5084,N_5209);
nand U7175 (N_7175,N_4972,N_4940);
xor U7176 (N_7176,N_5238,N_4584);
and U7177 (N_7177,N_5597,N_4866);
xor U7178 (N_7178,N_4916,N_5429);
or U7179 (N_7179,N_5534,N_5581);
or U7180 (N_7180,N_5138,N_5823);
nor U7181 (N_7181,N_5213,N_4647);
or U7182 (N_7182,N_5126,N_5669);
nor U7183 (N_7183,N_5034,N_5821);
and U7184 (N_7184,N_5699,N_5320);
nor U7185 (N_7185,N_5443,N_5826);
nor U7186 (N_7186,N_5054,N_4980);
or U7187 (N_7187,N_4669,N_4601);
or U7188 (N_7188,N_4831,N_4765);
nor U7189 (N_7189,N_5015,N_5030);
and U7190 (N_7190,N_4831,N_5044);
and U7191 (N_7191,N_4824,N_5770);
xnor U7192 (N_7192,N_5317,N_5043);
nor U7193 (N_7193,N_5106,N_4660);
nand U7194 (N_7194,N_4730,N_5563);
nand U7195 (N_7195,N_5712,N_5041);
and U7196 (N_7196,N_5053,N_5882);
and U7197 (N_7197,N_5637,N_4977);
and U7198 (N_7198,N_4530,N_5186);
xor U7199 (N_7199,N_5705,N_4936);
nand U7200 (N_7200,N_5324,N_5892);
and U7201 (N_7201,N_5659,N_5188);
and U7202 (N_7202,N_5268,N_4949);
nor U7203 (N_7203,N_4960,N_5657);
nand U7204 (N_7204,N_5030,N_5316);
or U7205 (N_7205,N_5199,N_5154);
xor U7206 (N_7206,N_5331,N_5338);
and U7207 (N_7207,N_5608,N_4656);
nand U7208 (N_7208,N_5424,N_5153);
or U7209 (N_7209,N_4544,N_5942);
nor U7210 (N_7210,N_5943,N_5477);
nor U7211 (N_7211,N_4720,N_5468);
nor U7212 (N_7212,N_5566,N_5767);
xnor U7213 (N_7213,N_5373,N_5345);
xnor U7214 (N_7214,N_5266,N_5509);
nand U7215 (N_7215,N_5110,N_4971);
xor U7216 (N_7216,N_5305,N_5977);
nor U7217 (N_7217,N_4676,N_4500);
or U7218 (N_7218,N_4782,N_4831);
nand U7219 (N_7219,N_5587,N_5402);
nand U7220 (N_7220,N_5369,N_4900);
nor U7221 (N_7221,N_5447,N_5451);
nand U7222 (N_7222,N_5176,N_5912);
nor U7223 (N_7223,N_5514,N_5124);
or U7224 (N_7224,N_5627,N_4952);
or U7225 (N_7225,N_5826,N_4689);
xor U7226 (N_7226,N_4563,N_5744);
or U7227 (N_7227,N_4673,N_5540);
nand U7228 (N_7228,N_4890,N_5061);
nand U7229 (N_7229,N_5499,N_5245);
xor U7230 (N_7230,N_4621,N_5922);
xor U7231 (N_7231,N_5120,N_4584);
or U7232 (N_7232,N_5010,N_5508);
nand U7233 (N_7233,N_5830,N_4984);
xnor U7234 (N_7234,N_5444,N_5733);
nor U7235 (N_7235,N_5199,N_4927);
nand U7236 (N_7236,N_5962,N_5870);
or U7237 (N_7237,N_5454,N_5879);
xor U7238 (N_7238,N_4841,N_5863);
nor U7239 (N_7239,N_5554,N_5678);
or U7240 (N_7240,N_5652,N_5984);
nand U7241 (N_7241,N_5631,N_5809);
nor U7242 (N_7242,N_5978,N_5648);
nand U7243 (N_7243,N_4751,N_5394);
xnor U7244 (N_7244,N_5307,N_5162);
and U7245 (N_7245,N_5256,N_5982);
nand U7246 (N_7246,N_5259,N_5250);
nor U7247 (N_7247,N_4539,N_5812);
and U7248 (N_7248,N_5177,N_5213);
nand U7249 (N_7249,N_4760,N_5970);
and U7250 (N_7250,N_5167,N_4821);
and U7251 (N_7251,N_5379,N_5381);
nor U7252 (N_7252,N_5458,N_5762);
nand U7253 (N_7253,N_5416,N_5938);
xnor U7254 (N_7254,N_4654,N_5747);
and U7255 (N_7255,N_5198,N_5843);
or U7256 (N_7256,N_5932,N_4852);
or U7257 (N_7257,N_5285,N_5066);
or U7258 (N_7258,N_5319,N_4599);
or U7259 (N_7259,N_4695,N_5728);
nor U7260 (N_7260,N_5882,N_4562);
nor U7261 (N_7261,N_4767,N_5284);
nand U7262 (N_7262,N_5459,N_5633);
nor U7263 (N_7263,N_4641,N_5729);
and U7264 (N_7264,N_4687,N_5953);
and U7265 (N_7265,N_5148,N_5961);
nand U7266 (N_7266,N_5922,N_5774);
xor U7267 (N_7267,N_4824,N_5222);
xnor U7268 (N_7268,N_4792,N_5993);
nand U7269 (N_7269,N_5321,N_5158);
nor U7270 (N_7270,N_4541,N_5815);
nor U7271 (N_7271,N_4947,N_5401);
and U7272 (N_7272,N_5910,N_5576);
and U7273 (N_7273,N_4855,N_5976);
nand U7274 (N_7274,N_5027,N_5445);
nor U7275 (N_7275,N_4884,N_4693);
xor U7276 (N_7276,N_4705,N_5476);
or U7277 (N_7277,N_5884,N_5921);
nor U7278 (N_7278,N_4829,N_5999);
or U7279 (N_7279,N_4895,N_4735);
nand U7280 (N_7280,N_5525,N_5677);
nor U7281 (N_7281,N_5883,N_4775);
xor U7282 (N_7282,N_5048,N_5005);
or U7283 (N_7283,N_5151,N_5274);
nor U7284 (N_7284,N_4946,N_4955);
nand U7285 (N_7285,N_5382,N_5875);
and U7286 (N_7286,N_5876,N_5238);
or U7287 (N_7287,N_5730,N_4613);
and U7288 (N_7288,N_5752,N_4737);
and U7289 (N_7289,N_5634,N_5431);
nor U7290 (N_7290,N_4553,N_4666);
xnor U7291 (N_7291,N_4688,N_4904);
nand U7292 (N_7292,N_5025,N_4805);
nor U7293 (N_7293,N_5363,N_5613);
and U7294 (N_7294,N_5443,N_5656);
nand U7295 (N_7295,N_5212,N_5194);
nand U7296 (N_7296,N_5490,N_4930);
xor U7297 (N_7297,N_5765,N_4817);
nand U7298 (N_7298,N_5213,N_5045);
xnor U7299 (N_7299,N_5669,N_5783);
xor U7300 (N_7300,N_5864,N_4690);
xor U7301 (N_7301,N_5788,N_4730);
xnor U7302 (N_7302,N_4659,N_5768);
and U7303 (N_7303,N_4780,N_5722);
nor U7304 (N_7304,N_5568,N_5047);
and U7305 (N_7305,N_5063,N_5153);
nand U7306 (N_7306,N_5749,N_5074);
or U7307 (N_7307,N_5067,N_5025);
or U7308 (N_7308,N_5254,N_5499);
nor U7309 (N_7309,N_5071,N_5228);
xor U7310 (N_7310,N_5789,N_5031);
nor U7311 (N_7311,N_5005,N_5394);
nor U7312 (N_7312,N_5172,N_5569);
or U7313 (N_7313,N_5817,N_5882);
and U7314 (N_7314,N_4660,N_4510);
or U7315 (N_7315,N_5159,N_5091);
and U7316 (N_7316,N_5893,N_5394);
and U7317 (N_7317,N_4966,N_4973);
and U7318 (N_7318,N_5859,N_4749);
or U7319 (N_7319,N_5838,N_5944);
nand U7320 (N_7320,N_5267,N_5447);
xnor U7321 (N_7321,N_5844,N_4941);
nor U7322 (N_7322,N_5208,N_5583);
and U7323 (N_7323,N_4879,N_4882);
nand U7324 (N_7324,N_4968,N_4598);
or U7325 (N_7325,N_5537,N_5391);
nor U7326 (N_7326,N_5535,N_5504);
or U7327 (N_7327,N_5954,N_5461);
nor U7328 (N_7328,N_4827,N_5780);
nand U7329 (N_7329,N_4854,N_5680);
nor U7330 (N_7330,N_5911,N_5924);
and U7331 (N_7331,N_5537,N_5147);
or U7332 (N_7332,N_5716,N_5456);
xnor U7333 (N_7333,N_5107,N_4669);
or U7334 (N_7334,N_5941,N_5159);
or U7335 (N_7335,N_5427,N_5659);
or U7336 (N_7336,N_5235,N_5626);
or U7337 (N_7337,N_4741,N_4933);
nand U7338 (N_7338,N_5397,N_4853);
nor U7339 (N_7339,N_5239,N_5938);
or U7340 (N_7340,N_5583,N_4876);
and U7341 (N_7341,N_4871,N_4698);
xor U7342 (N_7342,N_5273,N_5707);
nor U7343 (N_7343,N_5833,N_4782);
or U7344 (N_7344,N_5630,N_5734);
nor U7345 (N_7345,N_5657,N_4639);
xor U7346 (N_7346,N_5813,N_5984);
xnor U7347 (N_7347,N_5708,N_5315);
nor U7348 (N_7348,N_5215,N_4938);
or U7349 (N_7349,N_5298,N_5161);
or U7350 (N_7350,N_4858,N_4805);
nand U7351 (N_7351,N_4718,N_5941);
or U7352 (N_7352,N_5831,N_5587);
and U7353 (N_7353,N_4865,N_5923);
nor U7354 (N_7354,N_5027,N_5453);
or U7355 (N_7355,N_4641,N_5591);
or U7356 (N_7356,N_4703,N_5478);
or U7357 (N_7357,N_5983,N_4731);
nand U7358 (N_7358,N_5628,N_5235);
or U7359 (N_7359,N_4752,N_4577);
xor U7360 (N_7360,N_5239,N_5381);
and U7361 (N_7361,N_5957,N_4714);
xor U7362 (N_7362,N_5819,N_5758);
nand U7363 (N_7363,N_4607,N_4585);
or U7364 (N_7364,N_4874,N_5963);
or U7365 (N_7365,N_4567,N_5676);
nor U7366 (N_7366,N_4516,N_4742);
xor U7367 (N_7367,N_5649,N_4961);
nand U7368 (N_7368,N_5270,N_4742);
xor U7369 (N_7369,N_5724,N_4827);
and U7370 (N_7370,N_4855,N_5607);
xor U7371 (N_7371,N_5944,N_5431);
and U7372 (N_7372,N_4820,N_5173);
xor U7373 (N_7373,N_4564,N_5651);
and U7374 (N_7374,N_4799,N_5764);
nor U7375 (N_7375,N_4642,N_4635);
xor U7376 (N_7376,N_5692,N_5372);
and U7377 (N_7377,N_5001,N_5909);
nand U7378 (N_7378,N_5602,N_4727);
xor U7379 (N_7379,N_5308,N_5791);
xnor U7380 (N_7380,N_5954,N_5843);
or U7381 (N_7381,N_4931,N_5957);
and U7382 (N_7382,N_5876,N_5297);
nand U7383 (N_7383,N_5882,N_4890);
xnor U7384 (N_7384,N_4792,N_5520);
xnor U7385 (N_7385,N_4787,N_4579);
nand U7386 (N_7386,N_5406,N_5486);
nand U7387 (N_7387,N_4763,N_4730);
xnor U7388 (N_7388,N_5205,N_4748);
and U7389 (N_7389,N_5898,N_5414);
nor U7390 (N_7390,N_5898,N_5148);
nand U7391 (N_7391,N_5949,N_5977);
or U7392 (N_7392,N_5949,N_5150);
and U7393 (N_7393,N_5293,N_4872);
nand U7394 (N_7394,N_4551,N_5271);
or U7395 (N_7395,N_4501,N_4642);
or U7396 (N_7396,N_5960,N_5485);
and U7397 (N_7397,N_4544,N_4757);
xnor U7398 (N_7398,N_5612,N_5187);
or U7399 (N_7399,N_4675,N_5080);
nor U7400 (N_7400,N_5682,N_5914);
nand U7401 (N_7401,N_4800,N_5746);
or U7402 (N_7402,N_4953,N_5776);
nand U7403 (N_7403,N_5709,N_4913);
xor U7404 (N_7404,N_4617,N_5218);
nor U7405 (N_7405,N_5089,N_4588);
nor U7406 (N_7406,N_5387,N_5830);
nor U7407 (N_7407,N_4588,N_4789);
nor U7408 (N_7408,N_5178,N_4639);
nand U7409 (N_7409,N_5175,N_4732);
or U7410 (N_7410,N_5672,N_5264);
xnor U7411 (N_7411,N_5400,N_4932);
xnor U7412 (N_7412,N_4913,N_5157);
or U7413 (N_7413,N_4877,N_5167);
nor U7414 (N_7414,N_5915,N_5492);
nor U7415 (N_7415,N_5427,N_5593);
nor U7416 (N_7416,N_5466,N_5988);
nand U7417 (N_7417,N_5070,N_5219);
or U7418 (N_7418,N_4909,N_5994);
nand U7419 (N_7419,N_4737,N_5533);
xor U7420 (N_7420,N_4922,N_5343);
and U7421 (N_7421,N_4743,N_4961);
xor U7422 (N_7422,N_5215,N_5714);
and U7423 (N_7423,N_5812,N_4794);
nand U7424 (N_7424,N_5968,N_5378);
nor U7425 (N_7425,N_5558,N_4939);
and U7426 (N_7426,N_4742,N_4560);
or U7427 (N_7427,N_5951,N_5187);
xor U7428 (N_7428,N_5415,N_5021);
xnor U7429 (N_7429,N_5244,N_4979);
nand U7430 (N_7430,N_4832,N_5542);
xnor U7431 (N_7431,N_5548,N_4645);
and U7432 (N_7432,N_5900,N_5763);
nor U7433 (N_7433,N_5495,N_5910);
nand U7434 (N_7434,N_5109,N_5339);
nor U7435 (N_7435,N_5830,N_4762);
xnor U7436 (N_7436,N_5161,N_5453);
nand U7437 (N_7437,N_4662,N_5634);
and U7438 (N_7438,N_4710,N_5031);
nor U7439 (N_7439,N_4678,N_4890);
nand U7440 (N_7440,N_5316,N_4753);
xor U7441 (N_7441,N_4629,N_4686);
nand U7442 (N_7442,N_4650,N_4897);
or U7443 (N_7443,N_5964,N_4677);
nand U7444 (N_7444,N_4825,N_5132);
or U7445 (N_7445,N_5219,N_5587);
or U7446 (N_7446,N_5578,N_4638);
or U7447 (N_7447,N_5756,N_5442);
and U7448 (N_7448,N_5497,N_5738);
xnor U7449 (N_7449,N_4550,N_4561);
nor U7450 (N_7450,N_5297,N_4847);
xor U7451 (N_7451,N_5426,N_4784);
nor U7452 (N_7452,N_5916,N_4778);
nand U7453 (N_7453,N_5784,N_4560);
xor U7454 (N_7454,N_5267,N_5530);
xnor U7455 (N_7455,N_4843,N_4940);
nand U7456 (N_7456,N_5283,N_4590);
nor U7457 (N_7457,N_5014,N_5721);
or U7458 (N_7458,N_5226,N_4636);
nand U7459 (N_7459,N_4708,N_4592);
or U7460 (N_7460,N_5389,N_5812);
xor U7461 (N_7461,N_4548,N_5927);
xor U7462 (N_7462,N_5515,N_5081);
nand U7463 (N_7463,N_5375,N_5011);
or U7464 (N_7464,N_5073,N_5122);
xnor U7465 (N_7465,N_5665,N_5042);
or U7466 (N_7466,N_5466,N_5677);
nand U7467 (N_7467,N_4887,N_4915);
and U7468 (N_7468,N_4645,N_5081);
or U7469 (N_7469,N_5726,N_4793);
xnor U7470 (N_7470,N_4829,N_5728);
or U7471 (N_7471,N_5007,N_5176);
or U7472 (N_7472,N_5660,N_4568);
xnor U7473 (N_7473,N_4644,N_5783);
or U7474 (N_7474,N_5223,N_5933);
nand U7475 (N_7475,N_4630,N_4527);
nor U7476 (N_7476,N_5216,N_5679);
or U7477 (N_7477,N_5122,N_4787);
or U7478 (N_7478,N_5585,N_5724);
or U7479 (N_7479,N_5917,N_5687);
xnor U7480 (N_7480,N_5579,N_5284);
nand U7481 (N_7481,N_4816,N_5807);
xor U7482 (N_7482,N_5025,N_4919);
and U7483 (N_7483,N_5354,N_5190);
nand U7484 (N_7484,N_4840,N_4851);
xnor U7485 (N_7485,N_5761,N_5544);
xor U7486 (N_7486,N_5372,N_4753);
xor U7487 (N_7487,N_5302,N_4878);
xor U7488 (N_7488,N_4528,N_5403);
nor U7489 (N_7489,N_5678,N_5426);
xor U7490 (N_7490,N_5248,N_5775);
nand U7491 (N_7491,N_5101,N_5532);
and U7492 (N_7492,N_5820,N_5886);
or U7493 (N_7493,N_5948,N_4700);
xor U7494 (N_7494,N_5273,N_5434);
and U7495 (N_7495,N_5641,N_5285);
nor U7496 (N_7496,N_5150,N_4820);
nand U7497 (N_7497,N_5869,N_4615);
and U7498 (N_7498,N_5508,N_4960);
nor U7499 (N_7499,N_5326,N_5917);
nor U7500 (N_7500,N_6816,N_7297);
xnor U7501 (N_7501,N_7412,N_7379);
xor U7502 (N_7502,N_6485,N_6401);
nand U7503 (N_7503,N_6328,N_6153);
and U7504 (N_7504,N_7021,N_7092);
nor U7505 (N_7505,N_6796,N_6189);
nand U7506 (N_7506,N_6897,N_6354);
xnor U7507 (N_7507,N_6156,N_6681);
xor U7508 (N_7508,N_7415,N_6716);
nand U7509 (N_7509,N_6037,N_7313);
or U7510 (N_7510,N_7263,N_7457);
nor U7511 (N_7511,N_6353,N_6122);
or U7512 (N_7512,N_6415,N_7130);
nor U7513 (N_7513,N_6036,N_6014);
nor U7514 (N_7514,N_7494,N_7119);
xor U7515 (N_7515,N_6024,N_7151);
nand U7516 (N_7516,N_6323,N_7198);
nor U7517 (N_7517,N_6809,N_7411);
xor U7518 (N_7518,N_6017,N_6900);
xnor U7519 (N_7519,N_6868,N_6668);
nor U7520 (N_7520,N_7281,N_7100);
or U7521 (N_7521,N_6850,N_6607);
and U7522 (N_7522,N_6302,N_6553);
and U7523 (N_7523,N_6713,N_6235);
xnor U7524 (N_7524,N_7228,N_6924);
or U7525 (N_7525,N_6314,N_7229);
or U7526 (N_7526,N_7161,N_6107);
nor U7527 (N_7527,N_7186,N_7044);
or U7528 (N_7528,N_6117,N_6594);
nor U7529 (N_7529,N_7256,N_7193);
or U7530 (N_7530,N_6665,N_6957);
xnor U7531 (N_7531,N_7476,N_6199);
or U7532 (N_7532,N_6335,N_6313);
or U7533 (N_7533,N_7454,N_6584);
and U7534 (N_7534,N_7355,N_6774);
nand U7535 (N_7535,N_7472,N_6982);
and U7536 (N_7536,N_7167,N_6987);
xor U7537 (N_7537,N_7022,N_7295);
or U7538 (N_7538,N_7141,N_6345);
nand U7539 (N_7539,N_7413,N_6740);
xor U7540 (N_7540,N_6016,N_6366);
or U7541 (N_7541,N_6089,N_6923);
nand U7542 (N_7542,N_6506,N_6000);
or U7543 (N_7543,N_7145,N_6265);
and U7544 (N_7544,N_6136,N_6085);
or U7545 (N_7545,N_6465,N_7093);
nor U7546 (N_7546,N_6944,N_7393);
or U7547 (N_7547,N_7220,N_7203);
xnor U7548 (N_7548,N_6130,N_6109);
and U7549 (N_7549,N_6775,N_7260);
and U7550 (N_7550,N_6438,N_6564);
nor U7551 (N_7551,N_7002,N_6510);
nand U7552 (N_7552,N_6480,N_6685);
nor U7553 (N_7553,N_6215,N_7210);
nor U7554 (N_7554,N_6046,N_6926);
and U7555 (N_7555,N_6773,N_7230);
xnor U7556 (N_7556,N_6601,N_7479);
or U7557 (N_7557,N_6347,N_6570);
xnor U7558 (N_7558,N_7239,N_6178);
nand U7559 (N_7559,N_6786,N_6116);
nor U7560 (N_7560,N_6249,N_6086);
nor U7561 (N_7561,N_6704,N_6708);
or U7562 (N_7562,N_6534,N_7366);
xor U7563 (N_7563,N_6195,N_6231);
and U7564 (N_7564,N_6884,N_7075);
or U7565 (N_7565,N_7324,N_6625);
nor U7566 (N_7566,N_6543,N_6243);
nand U7567 (N_7567,N_6246,N_6180);
xnor U7568 (N_7568,N_6444,N_6533);
or U7569 (N_7569,N_6292,N_6658);
and U7570 (N_7570,N_6197,N_6812);
nor U7571 (N_7571,N_6646,N_6018);
or U7572 (N_7572,N_6522,N_7270);
nor U7573 (N_7573,N_7316,N_7291);
nor U7574 (N_7574,N_6350,N_6127);
or U7575 (N_7575,N_6204,N_6971);
nor U7576 (N_7576,N_6050,N_6359);
and U7577 (N_7577,N_7327,N_7053);
and U7578 (N_7578,N_6747,N_6078);
or U7579 (N_7579,N_6733,N_6049);
nor U7580 (N_7580,N_6244,N_7041);
and U7581 (N_7581,N_7112,N_6709);
and U7582 (N_7582,N_7120,N_6922);
nor U7583 (N_7583,N_7081,N_6320);
or U7584 (N_7584,N_6279,N_6950);
xor U7585 (N_7585,N_7224,N_7309);
nand U7586 (N_7586,N_7206,N_6009);
xor U7587 (N_7587,N_6141,N_6008);
xnor U7588 (N_7588,N_6710,N_6696);
nor U7589 (N_7589,N_6815,N_6356);
xor U7590 (N_7590,N_7365,N_6660);
or U7591 (N_7591,N_7419,N_7337);
nor U7592 (N_7592,N_6984,N_7356);
or U7593 (N_7593,N_6055,N_7352);
nor U7594 (N_7594,N_6185,N_6737);
or U7595 (N_7595,N_6384,N_6842);
nor U7596 (N_7596,N_7090,N_6479);
or U7597 (N_7597,N_6126,N_6474);
nand U7598 (N_7598,N_7208,N_6834);
xor U7599 (N_7599,N_7487,N_7246);
nor U7600 (N_7600,N_7154,N_6002);
or U7601 (N_7601,N_7249,N_6393);
nor U7602 (N_7602,N_7101,N_6285);
and U7603 (N_7603,N_6011,N_6162);
or U7604 (N_7604,N_7368,N_6993);
and U7605 (N_7605,N_6357,N_6832);
or U7606 (N_7606,N_6382,N_6027);
and U7607 (N_7607,N_6020,N_6829);
nand U7608 (N_7608,N_6132,N_6449);
nor U7609 (N_7609,N_6579,N_6155);
nand U7610 (N_7610,N_6718,N_6568);
nand U7611 (N_7611,N_7212,N_6666);
and U7612 (N_7612,N_6213,N_7456);
and U7613 (N_7613,N_6613,N_6915);
xnor U7614 (N_7614,N_6258,N_6439);
and U7615 (N_7615,N_6380,N_7275);
xor U7616 (N_7616,N_6160,N_7417);
and U7617 (N_7617,N_7284,N_6839);
xnor U7618 (N_7618,N_7358,N_7331);
nor U7619 (N_7619,N_6652,N_7174);
or U7620 (N_7620,N_6170,N_6667);
nor U7621 (N_7621,N_7323,N_7032);
or U7622 (N_7622,N_7498,N_6207);
nor U7623 (N_7623,N_6206,N_6919);
or U7624 (N_7624,N_6073,N_6617);
and U7625 (N_7625,N_6416,N_7162);
and U7626 (N_7626,N_6288,N_6583);
nand U7627 (N_7627,N_6555,N_7084);
xnor U7628 (N_7628,N_6826,N_6720);
and U7629 (N_7629,N_6574,N_6454);
xor U7630 (N_7630,N_6424,N_7332);
nor U7631 (N_7631,N_6503,N_6742);
and U7632 (N_7632,N_6398,N_6598);
nand U7633 (N_7633,N_7303,N_6496);
nand U7634 (N_7634,N_6260,N_7404);
or U7635 (N_7635,N_6348,N_7262);
nand U7636 (N_7636,N_6434,N_6929);
xnor U7637 (N_7637,N_6105,N_6851);
and U7638 (N_7638,N_7395,N_7131);
nor U7639 (N_7639,N_6840,N_7038);
or U7640 (N_7640,N_6032,N_7361);
nand U7641 (N_7641,N_7138,N_6705);
and U7642 (N_7642,N_7216,N_6080);
nand U7643 (N_7643,N_6340,N_6784);
nor U7644 (N_7644,N_6643,N_6837);
or U7645 (N_7645,N_6491,N_7010);
nand U7646 (N_7646,N_6377,N_7460);
and U7647 (N_7647,N_6701,N_6453);
nand U7648 (N_7648,N_6606,N_7347);
nor U7649 (N_7649,N_6163,N_6375);
xnor U7650 (N_7650,N_7423,N_7459);
nand U7651 (N_7651,N_6248,N_6659);
nand U7652 (N_7652,N_7108,N_6931);
xnor U7653 (N_7653,N_7274,N_6270);
nand U7654 (N_7654,N_6626,N_6966);
xor U7655 (N_7655,N_7006,N_7036);
xor U7656 (N_7656,N_7381,N_6226);
xnor U7657 (N_7657,N_7078,N_6630);
and U7658 (N_7658,N_6788,N_6818);
xor U7659 (N_7659,N_6400,N_6410);
and U7660 (N_7660,N_6042,N_6164);
nand U7661 (N_7661,N_7478,N_7047);
or U7662 (N_7662,N_6303,N_6542);
xor U7663 (N_7663,N_7265,N_6167);
nor U7664 (N_7664,N_6239,N_6310);
and U7665 (N_7665,N_6935,N_6979);
xor U7666 (N_7666,N_6822,N_6914);
nand U7667 (N_7667,N_7200,N_6093);
xor U7668 (N_7668,N_6940,N_7083);
xnor U7669 (N_7669,N_6462,N_6906);
nor U7670 (N_7670,N_6166,N_6233);
nand U7671 (N_7671,N_7367,N_6151);
nand U7672 (N_7672,N_6039,N_6111);
nand U7673 (N_7673,N_6925,N_7168);
and U7674 (N_7674,N_6547,N_6804);
xor U7675 (N_7675,N_6365,N_6181);
nand U7676 (N_7676,N_7211,N_7292);
nor U7677 (N_7677,N_6806,N_7434);
and U7678 (N_7678,N_7087,N_7453);
xor U7679 (N_7679,N_6849,N_6290);
and U7680 (N_7680,N_6582,N_7444);
xnor U7681 (N_7681,N_6332,N_7049);
nand U7682 (N_7682,N_6342,N_6566);
or U7683 (N_7683,N_7346,N_6403);
nand U7684 (N_7684,N_6592,N_6487);
xor U7685 (N_7685,N_7004,N_6634);
nand U7686 (N_7686,N_6835,N_6827);
and U7687 (N_7687,N_7402,N_6220);
nor U7688 (N_7688,N_6891,N_7406);
xnor U7689 (N_7689,N_6511,N_6045);
xor U7690 (N_7690,N_7317,N_7429);
nor U7691 (N_7691,N_6425,N_6744);
nand U7692 (N_7692,N_7321,N_6986);
nor U7693 (N_7693,N_7267,N_6945);
or U7694 (N_7694,N_6369,N_7152);
nand U7695 (N_7695,N_6655,N_6072);
or U7696 (N_7696,N_6459,N_7113);
and U7697 (N_7697,N_6799,N_7180);
nand U7698 (N_7698,N_6110,N_6289);
nand U7699 (N_7699,N_6060,N_6992);
xnor U7700 (N_7700,N_7255,N_6322);
nor U7701 (N_7701,N_7136,N_7377);
xor U7702 (N_7702,N_6560,N_6603);
nor U7703 (N_7703,N_6996,N_6174);
and U7704 (N_7704,N_6507,N_6712);
nand U7705 (N_7705,N_7003,N_6108);
and U7706 (N_7706,N_6476,N_6844);
or U7707 (N_7707,N_6255,N_7060);
nand U7708 (N_7708,N_6161,N_6470);
nand U7709 (N_7709,N_6087,N_7050);
xnor U7710 (N_7710,N_6787,N_6767);
nand U7711 (N_7711,N_6682,N_6536);
nand U7712 (N_7712,N_6406,N_6719);
nand U7713 (N_7713,N_6103,N_7240);
xnor U7714 (N_7714,N_6252,N_6885);
nor U7715 (N_7715,N_6308,N_7447);
nand U7716 (N_7716,N_6721,N_7351);
nand U7717 (N_7717,N_6274,N_6730);
nor U7718 (N_7718,N_6590,N_6472);
and U7719 (N_7719,N_6304,N_7371);
xnor U7720 (N_7720,N_6053,N_6192);
and U7721 (N_7721,N_6911,N_7272);
nand U7722 (N_7722,N_6811,N_7149);
nand U7723 (N_7723,N_6693,N_7405);
nand U7724 (N_7724,N_7294,N_6749);
nor U7725 (N_7725,N_6149,N_6988);
or U7726 (N_7726,N_6760,N_7024);
or U7727 (N_7727,N_6673,N_6183);
or U7728 (N_7728,N_6113,N_6545);
and U7729 (N_7729,N_6585,N_6808);
or U7730 (N_7730,N_7349,N_6154);
nor U7731 (N_7731,N_6176,N_6865);
and U7732 (N_7732,N_6970,N_6725);
xnor U7733 (N_7733,N_7278,N_6137);
nor U7734 (N_7734,N_6182,N_7340);
nand U7735 (N_7735,N_7124,N_6841);
nand U7736 (N_7736,N_6650,N_6254);
xor U7737 (N_7737,N_7013,N_7028);
nor U7738 (N_7738,N_7009,N_6781);
or U7739 (N_7739,N_6662,N_6750);
nor U7740 (N_7740,N_6234,N_6836);
xnor U7741 (N_7741,N_6529,N_7362);
nor U7742 (N_7742,N_7132,N_6789);
xor U7743 (N_7743,N_6422,N_6599);
xor U7744 (N_7744,N_7410,N_6862);
xor U7745 (N_7745,N_6229,N_6972);
nand U7746 (N_7746,N_6502,N_6440);
and U7747 (N_7747,N_6724,N_7308);
nand U7748 (N_7748,N_6916,N_6028);
xnor U7749 (N_7749,N_6101,N_6266);
and U7750 (N_7750,N_6441,N_7475);
xnor U7751 (N_7751,N_6663,N_6223);
nor U7752 (N_7752,N_6908,N_7289);
or U7753 (N_7753,N_7178,N_6985);
nand U7754 (N_7754,N_7357,N_7033);
nand U7755 (N_7755,N_7462,N_6031);
nand U7756 (N_7756,N_7104,N_6913);
nand U7757 (N_7757,N_7226,N_6820);
nand U7758 (N_7758,N_6211,N_6515);
and U7759 (N_7759,N_6540,N_6586);
or U7760 (N_7760,N_6346,N_6436);
nand U7761 (N_7761,N_7236,N_6448);
or U7762 (N_7762,N_6427,N_6899);
nor U7763 (N_7763,N_6711,N_6386);
or U7764 (N_7764,N_6561,N_7477);
or U7765 (N_7765,N_6981,N_6129);
nand U7766 (N_7766,N_7116,N_6208);
xnor U7767 (N_7767,N_6272,N_6677);
or U7768 (N_7768,N_7282,N_6146);
nand U7769 (N_7769,N_6418,N_7252);
nor U7770 (N_7770,N_7118,N_7428);
and U7771 (N_7771,N_7209,N_7458);
nor U7772 (N_7772,N_7139,N_7056);
nand U7773 (N_7773,N_6904,N_6281);
nand U7774 (N_7774,N_7133,N_7330);
nor U7775 (N_7775,N_6261,N_6245);
or U7776 (N_7776,N_6135,N_6700);
and U7777 (N_7777,N_6828,N_6473);
nand U7778 (N_7778,N_6959,N_7266);
and U7779 (N_7779,N_7468,N_6397);
and U7780 (N_7780,N_6286,N_6684);
or U7781 (N_7781,N_6691,N_7126);
and U7782 (N_7782,N_6963,N_6445);
and U7783 (N_7783,N_6670,N_6819);
or U7784 (N_7784,N_6637,N_6683);
nor U7785 (N_7785,N_6573,N_6307);
or U7786 (N_7786,N_7205,N_6358);
nor U7787 (N_7787,N_7320,N_6873);
xor U7788 (N_7788,N_6723,N_7189);
nand U7789 (N_7789,N_6692,N_6467);
and U7790 (N_7790,N_6661,N_7285);
nor U7791 (N_7791,N_6977,N_6608);
nor U7792 (N_7792,N_6118,N_6224);
or U7793 (N_7793,N_6589,N_6654);
nor U7794 (N_7794,N_6404,N_6222);
xnor U7795 (N_7795,N_6329,N_7461);
xnor U7796 (N_7796,N_6324,N_6186);
nor U7797 (N_7797,N_6538,N_7353);
nor U7798 (N_7798,N_6896,N_7020);
nand U7799 (N_7799,N_6600,N_6813);
nand U7800 (N_7800,N_7109,N_6757);
and U7801 (N_7801,N_6388,N_6228);
nor U7802 (N_7802,N_6847,N_7467);
xnor U7803 (N_7803,N_7484,N_6690);
xnor U7804 (N_7804,N_6326,N_7440);
or U7805 (N_7805,N_6771,N_6070);
nand U7806 (N_7806,N_7103,N_7250);
nor U7807 (N_7807,N_7076,N_7137);
or U7808 (N_7808,N_7376,N_6785);
and U7809 (N_7809,N_6079,N_7385);
xnor U7810 (N_7810,N_6635,N_6807);
and U7811 (N_7811,N_7300,N_6179);
and U7812 (N_7812,N_6565,N_6952);
or U7813 (N_7813,N_7023,N_7128);
or U7814 (N_7814,N_6707,N_6975);
xnor U7815 (N_7815,N_7296,N_6588);
and U7816 (N_7816,N_6334,N_6864);
xnor U7817 (N_7817,N_6859,N_6408);
or U7818 (N_7818,N_7359,N_6619);
nor U7819 (N_7819,N_6482,N_7435);
nand U7820 (N_7820,N_7223,N_7218);
nand U7821 (N_7821,N_6013,N_6339);
xnor U7822 (N_7822,N_6918,N_6947);
or U7823 (N_7823,N_6509,N_6257);
nand U7824 (N_7824,N_6642,N_6552);
nand U7825 (N_7825,N_7301,N_7222);
or U7826 (N_7826,N_6641,N_6853);
xnor U7827 (N_7827,N_6414,N_6362);
nor U7828 (N_7828,N_7370,N_6483);
xnor U7829 (N_7829,N_6695,N_6190);
nand U7830 (N_7830,N_7311,N_7336);
nor U7831 (N_7831,N_6455,N_6316);
and U7832 (N_7832,N_6953,N_6435);
xnor U7833 (N_7833,N_7052,N_6240);
or U7834 (N_7834,N_7072,N_7019);
and U7835 (N_7835,N_6490,N_6488);
and U7836 (N_7836,N_6044,N_7293);
or U7837 (N_7837,N_7392,N_7325);
xor U7838 (N_7838,N_6604,N_7213);
or U7839 (N_7839,N_6765,N_7172);
xor U7840 (N_7840,N_6012,N_6934);
xor U7841 (N_7841,N_7470,N_7391);
xor U7842 (N_7842,N_6318,N_7463);
and U7843 (N_7843,N_6022,N_6391);
and U7844 (N_7844,N_6264,N_6023);
or U7845 (N_7845,N_7018,N_7062);
nor U7846 (N_7846,N_6120,N_7445);
or U7847 (N_7847,N_6937,N_6201);
nor U7848 (N_7848,N_7054,N_6430);
xnor U7849 (N_7849,N_6015,N_6405);
nand U7850 (N_7850,N_7398,N_6595);
xnor U7851 (N_7851,N_6429,N_6276);
or U7852 (N_7852,N_7110,N_7027);
and U7853 (N_7853,N_6493,N_6351);
nand U7854 (N_7854,N_6743,N_6769);
or U7855 (N_7855,N_6738,N_6399);
xnor U7856 (N_7856,N_6876,N_6040);
nand U7857 (N_7857,N_6291,N_6698);
nand U7858 (N_7858,N_6287,N_6726);
nand U7859 (N_7859,N_6217,N_6768);
nor U7860 (N_7860,N_6620,N_7315);
nor U7861 (N_7861,N_6267,N_6385);
nor U7862 (N_7862,N_6991,N_6390);
nand U7863 (N_7863,N_6212,N_7432);
nor U7864 (N_7864,N_7227,N_6722);
nor U7865 (N_7865,N_6762,N_7102);
nor U7866 (N_7866,N_7369,N_6221);
xor U7867 (N_7867,N_6735,N_6657);
nor U7868 (N_7868,N_7215,N_6958);
xor U7869 (N_7869,N_6144,N_6946);
and U7870 (N_7870,N_6857,N_6063);
and U7871 (N_7871,N_6337,N_7001);
or U7872 (N_7872,N_6321,N_6729);
nand U7873 (N_7873,N_6858,N_6138);
xnor U7874 (N_7874,N_6051,N_6145);
and U7875 (N_7875,N_6360,N_7175);
nor U7876 (N_7876,N_7443,N_6026);
and U7877 (N_7877,N_7146,N_6633);
or U7878 (N_7878,N_6372,N_6428);
nor U7879 (N_7879,N_7287,N_6083);
or U7880 (N_7880,N_6825,N_6352);
nand U7881 (N_7881,N_7283,N_6200);
or U7882 (N_7882,N_6621,N_7214);
and U7883 (N_7883,N_6331,N_7156);
nand U7884 (N_7884,N_7007,N_7058);
nor U7885 (N_7885,N_6336,N_6296);
xor U7886 (N_7886,N_7191,N_6901);
xnor U7887 (N_7887,N_6779,N_6780);
or U7888 (N_7888,N_6715,N_6193);
or U7889 (N_7889,N_6753,N_7492);
xnor U7890 (N_7890,N_6644,N_6466);
nand U7891 (N_7891,N_7196,N_7181);
nand U7892 (N_7892,N_6955,N_6995);
xor U7893 (N_7893,N_6173,N_6525);
or U7894 (N_7894,N_7170,N_6082);
and U7895 (N_7895,N_6202,N_6628);
and U7896 (N_7896,N_6437,N_7111);
nor U7897 (N_7897,N_6803,N_6653);
xnor U7898 (N_7898,N_7234,N_6519);
xor U7899 (N_7899,N_6833,N_6810);
or U7900 (N_7900,N_6047,N_7150);
and U7901 (N_7901,N_6392,N_6319);
nand U7902 (N_7902,N_7177,N_6311);
xor U7903 (N_7903,N_6283,N_6495);
or U7904 (N_7904,N_7436,N_7442);
and U7905 (N_7905,N_6790,N_7166);
nor U7906 (N_7906,N_6315,N_6412);
or U7907 (N_7907,N_7204,N_6535);
and U7908 (N_7908,N_7159,N_6824);
xnor U7909 (N_7909,N_7097,N_7179);
and U7910 (N_7910,N_6327,N_6845);
nor U7911 (N_7911,N_6196,N_6933);
or U7912 (N_7912,N_6305,N_6941);
nand U7913 (N_7913,N_6148,N_7135);
xnor U7914 (N_7914,N_7437,N_6091);
nor U7915 (N_7915,N_6489,N_7448);
nand U7916 (N_7916,N_7094,N_7363);
or U7917 (N_7917,N_6477,N_6782);
nor U7918 (N_7918,N_6299,N_6232);
xnor U7919 (N_7919,N_7482,N_7497);
nand U7920 (N_7920,N_6734,N_6413);
xnor U7921 (N_7921,N_6088,N_6306);
or U7922 (N_7922,N_7399,N_6298);
nand U7923 (N_7923,N_6687,N_7066);
xnor U7924 (N_7924,N_7067,N_7258);
nand U7925 (N_7925,N_7446,N_6094);
xor U7926 (N_7926,N_6843,N_7276);
xnor U7927 (N_7927,N_7396,N_7288);
and U7928 (N_7928,N_7016,N_7305);
or U7929 (N_7929,N_6559,N_6877);
and U7930 (N_7930,N_7207,N_6838);
or U7931 (N_7931,N_7187,N_6805);
nand U7932 (N_7932,N_6949,N_6989);
xor U7933 (N_7933,N_6067,N_6983);
nor U7934 (N_7934,N_6800,N_6184);
and U7935 (N_7935,N_6317,N_6830);
or U7936 (N_7936,N_6333,N_7425);
xnor U7937 (N_7937,N_6518,N_7188);
or U7938 (N_7938,N_6419,N_7106);
xnor U7939 (N_7939,N_6005,N_6624);
or U7940 (N_7940,N_7433,N_6387);
xnor U7941 (N_7941,N_6575,N_6061);
nand U7942 (N_7942,N_7390,N_6759);
xnor U7943 (N_7943,N_7184,N_6098);
nand U7944 (N_7944,N_7025,N_6976);
nand U7945 (N_7945,N_6054,N_6486);
and U7946 (N_7946,N_6764,N_7426);
nand U7947 (N_7947,N_6481,N_6892);
or U7948 (N_7948,N_6100,N_6379);
or U7949 (N_7949,N_6539,N_6587);
nor U7950 (N_7950,N_6821,N_6817);
or U7951 (N_7951,N_6363,N_6175);
nand U7952 (N_7952,N_6562,N_6866);
or U7953 (N_7953,N_7143,N_7345);
nor U7954 (N_7954,N_7235,N_7341);
nor U7955 (N_7955,N_6852,N_6717);
or U7956 (N_7956,N_6938,N_6649);
nand U7957 (N_7957,N_6939,N_6732);
nand U7958 (N_7958,N_6210,N_7354);
nor U7959 (N_7959,N_7098,N_6458);
nand U7960 (N_7960,N_6499,N_6203);
nand U7961 (N_7961,N_6823,N_6112);
or U7962 (N_7962,N_6096,N_6741);
nor U7963 (N_7963,N_6505,N_7247);
and U7964 (N_7964,N_6706,N_7483);
or U7965 (N_7965,N_6898,N_6861);
or U7966 (N_7966,N_6569,N_6227);
nor U7967 (N_7967,N_6038,N_6974);
nand U7968 (N_7968,N_6500,N_7326);
nand U7969 (N_7969,N_6846,N_7190);
nor U7970 (N_7970,N_7243,N_6451);
and U7971 (N_7971,N_6645,N_6128);
or U7972 (N_7972,N_6250,N_7430);
nor U7973 (N_7973,N_6596,N_6389);
xnor U7974 (N_7974,N_6927,N_7299);
or U7975 (N_7975,N_6795,N_6075);
nand U7976 (N_7976,N_6010,N_7029);
xor U7977 (N_7977,N_7400,N_7489);
nand U7978 (N_7978,N_6269,N_7490);
xor U7979 (N_7979,N_6158,N_6463);
nor U7980 (N_7980,N_6033,N_7251);
or U7981 (N_7981,N_6680,N_7232);
nor U7982 (N_7982,N_7464,N_7147);
and U7983 (N_7983,N_6256,N_6278);
or U7984 (N_7984,N_7000,N_6514);
nand U7985 (N_7985,N_6770,N_6763);
xor U7986 (N_7986,N_6421,N_6003);
xnor U7987 (N_7987,N_7343,N_7082);
xnor U7988 (N_7988,N_6802,N_6237);
or U7989 (N_7989,N_6097,N_7407);
and U7990 (N_7990,N_7408,N_6471);
xnor U7991 (N_7991,N_6095,N_6263);
xnor U7992 (N_7992,N_7389,N_6025);
or U7993 (N_7993,N_6065,N_6697);
xor U7994 (N_7994,N_6124,N_6165);
nand U7995 (N_7995,N_6581,N_6867);
and U7996 (N_7996,N_6447,N_7350);
xnor U7997 (N_7997,N_6656,N_6772);
nor U7998 (N_7998,N_6880,N_6856);
nor U7999 (N_7999,N_6411,N_7129);
nand U8000 (N_8000,N_6456,N_6030);
xor U8001 (N_8001,N_6669,N_6119);
nand U8002 (N_8002,N_6280,N_6524);
or U8003 (N_8003,N_6631,N_6139);
nor U8004 (N_8004,N_6544,N_7195);
or U8005 (N_8005,N_7153,N_7261);
and U8006 (N_8006,N_6077,N_6614);
or U8007 (N_8007,N_7171,N_6157);
xor U8008 (N_8008,N_6887,N_7034);
xor U8009 (N_8009,N_6433,N_6567);
nand U8010 (N_8010,N_6373,N_6464);
and U8011 (N_8011,N_6251,N_6344);
or U8012 (N_8012,N_7040,N_6578);
nand U8013 (N_8013,N_7414,N_6370);
nand U8014 (N_8014,N_6301,N_6282);
or U8015 (N_8015,N_6035,N_6968);
and U8016 (N_8016,N_6492,N_7031);
or U8017 (N_8017,N_7388,N_7089);
nand U8018 (N_8018,N_7334,N_6636);
nor U8019 (N_8019,N_7107,N_7014);
or U8020 (N_8020,N_6557,N_7387);
nand U8021 (N_8021,N_6610,N_6494);
or U8022 (N_8022,N_6426,N_7328);
nor U8023 (N_8023,N_6550,N_6879);
xnor U8024 (N_8024,N_7488,N_6874);
and U8025 (N_8025,N_6300,N_7286);
xor U8026 (N_8026,N_6478,N_7302);
and U8027 (N_8027,N_6766,N_7382);
or U8028 (N_8028,N_7048,N_7074);
nor U8029 (N_8029,N_6048,N_6689);
nor U8030 (N_8030,N_6071,N_7485);
or U8031 (N_8031,N_7069,N_6236);
and U8032 (N_8032,N_6532,N_7441);
or U8033 (N_8033,N_6423,N_7314);
xor U8034 (N_8034,N_6576,N_7144);
or U8035 (N_8035,N_6609,N_7493);
or U8036 (N_8036,N_6854,N_7455);
and U8037 (N_8037,N_6672,N_6639);
nand U8038 (N_8038,N_7244,N_6253);
or U8039 (N_8039,N_6034,N_7183);
xnor U8040 (N_8040,N_6973,N_7312);
nor U8041 (N_8041,N_6106,N_7071);
or U8042 (N_8042,N_6062,N_6355);
and U8043 (N_8043,N_6218,N_6541);
nand U8044 (N_8044,N_6870,N_7225);
nand U8045 (N_8045,N_6497,N_6549);
nor U8046 (N_8046,N_6531,N_6443);
or U8047 (N_8047,N_6242,N_7042);
or U8048 (N_8048,N_7045,N_6622);
or U8049 (N_8049,N_6527,N_6394);
nor U8050 (N_8050,N_7115,N_7386);
or U8051 (N_8051,N_6219,N_6104);
nand U8052 (N_8052,N_6041,N_6792);
or U8053 (N_8053,N_6225,N_6194);
or U8054 (N_8054,N_6376,N_7298);
nand U8055 (N_8055,N_6131,N_6558);
nand U8056 (N_8056,N_6090,N_7329);
or U8057 (N_8057,N_6504,N_6883);
or U8058 (N_8058,N_6216,N_7199);
nand U8059 (N_8059,N_7333,N_6990);
nand U8060 (N_8060,N_6123,N_6520);
nor U8061 (N_8061,N_7134,N_6640);
or U8062 (N_8062,N_7397,N_6942);
xor U8063 (N_8063,N_7017,N_6678);
and U8064 (N_8064,N_6930,N_6007);
nor U8065 (N_8065,N_7342,N_6241);
and U8066 (N_8066,N_6508,N_7005);
nor U8067 (N_8067,N_6591,N_7242);
or U8068 (N_8068,N_6848,N_6727);
nand U8069 (N_8069,N_7273,N_6894);
or U8070 (N_8070,N_7063,N_6513);
and U8071 (N_8071,N_7182,N_6728);
or U8072 (N_8072,N_6142,N_7011);
and U8073 (N_8073,N_6450,N_7378);
or U8074 (N_8074,N_6739,N_6675);
nor U8075 (N_8075,N_7030,N_6383);
or U8076 (N_8076,N_6546,N_6756);
nand U8077 (N_8077,N_7086,N_6912);
and U8078 (N_8078,N_6297,N_7248);
xor U8079 (N_8079,N_7192,N_6152);
and U8080 (N_8080,N_6755,N_6115);
or U8081 (N_8081,N_6797,N_7360);
xnor U8082 (N_8082,N_6066,N_6468);
or U8083 (N_8083,N_6702,N_6309);
and U8084 (N_8084,N_6745,N_7280);
nand U8085 (N_8085,N_7123,N_6960);
xnor U8086 (N_8086,N_6021,N_6205);
xor U8087 (N_8087,N_6647,N_6188);
nor U8088 (N_8088,N_7465,N_6731);
or U8089 (N_8089,N_7176,N_6580);
or U8090 (N_8090,N_6168,N_6875);
or U8091 (N_8091,N_6530,N_7114);
and U8092 (N_8092,N_7449,N_6736);
nor U8093 (N_8093,N_6460,N_6863);
or U8094 (N_8094,N_7008,N_6001);
and U8095 (N_8095,N_6407,N_7480);
nor U8096 (N_8096,N_6247,N_7471);
or U8097 (N_8097,N_7438,N_7450);
or U8098 (N_8098,N_6475,N_7080);
nor U8099 (N_8099,N_6159,N_6616);
xnor U8100 (N_8100,N_7418,N_7427);
and U8101 (N_8101,N_6064,N_6629);
nand U8102 (N_8102,N_6209,N_7451);
and U8103 (N_8103,N_6754,N_6259);
nor U8104 (N_8104,N_7015,N_6374);
nor U8105 (N_8105,N_6627,N_6651);
nand U8106 (N_8106,N_6618,N_7486);
nand U8107 (N_8107,N_6501,N_6902);
nor U8108 (N_8108,N_6537,N_7043);
nand U8109 (N_8109,N_7070,N_6994);
or U8110 (N_8110,N_7035,N_7185);
and U8111 (N_8111,N_6230,N_7201);
nand U8112 (N_8112,N_6615,N_7057);
or U8113 (N_8113,N_6978,N_6084);
nand U8114 (N_8114,N_6563,N_7344);
xor U8115 (N_8115,N_6273,N_6431);
or U8116 (N_8116,N_7335,N_6860);
or U8117 (N_8117,N_6703,N_6814);
nand U8118 (N_8118,N_7237,N_6099);
or U8119 (N_8119,N_7233,N_7164);
or U8120 (N_8120,N_6794,N_6150);
or U8121 (N_8121,N_6177,N_7290);
nand U8122 (N_8122,N_7264,N_7257);
nor U8123 (N_8123,N_7155,N_7373);
and U8124 (N_8124,N_7383,N_7452);
or U8125 (N_8125,N_6187,N_7499);
and U8126 (N_8126,N_6056,N_6623);
nand U8127 (N_8127,N_7064,N_6572);
and U8128 (N_8128,N_6452,N_6548);
nand U8129 (N_8129,N_6312,N_7409);
xnor U8130 (N_8130,N_6969,N_7380);
and U8131 (N_8131,N_6277,N_6121);
or U8132 (N_8132,N_6593,N_6381);
nand U8133 (N_8133,N_6004,N_7197);
xor U8134 (N_8134,N_6368,N_6791);
xnor U8135 (N_8135,N_6783,N_6364);
xnor U8136 (N_8136,N_6457,N_7158);
or U8137 (N_8137,N_7421,N_7073);
or U8138 (N_8138,N_6909,N_6903);
nand U8139 (N_8139,N_7061,N_7241);
xnor U8140 (N_8140,N_7142,N_7238);
or U8141 (N_8141,N_6571,N_7403);
nor U8142 (N_8142,N_6612,N_7165);
and U8143 (N_8143,N_7046,N_7374);
or U8144 (N_8144,N_6878,N_6999);
nor U8145 (N_8145,N_6526,N_6058);
and U8146 (N_8146,N_7173,N_6516);
and U8147 (N_8147,N_6461,N_6338);
nor U8148 (N_8148,N_6664,N_7431);
xor U8149 (N_8149,N_6889,N_7169);
or U8150 (N_8150,N_6602,N_6140);
nand U8151 (N_8151,N_6133,N_6556);
and U8152 (N_8152,N_6330,N_6521);
or U8153 (N_8153,N_6855,N_7473);
or U8154 (N_8154,N_7026,N_6831);
xor U8155 (N_8155,N_6632,N_6198);
nor U8156 (N_8156,N_6998,N_7253);
nand U8157 (N_8157,N_6888,N_7091);
xnor U8158 (N_8158,N_6905,N_6962);
and U8159 (N_8159,N_7117,N_6932);
xnor U8160 (N_8160,N_6059,N_7217);
and U8161 (N_8161,N_6967,N_6284);
xnor U8162 (N_8162,N_7481,N_7099);
or U8163 (N_8163,N_6752,N_6961);
nor U8164 (N_8164,N_6928,N_6402);
xor U8165 (N_8165,N_6057,N_7221);
nand U8166 (N_8166,N_6776,N_6638);
nor U8167 (N_8167,N_6361,N_7338);
or U8168 (N_8168,N_7245,N_6758);
nor U8169 (N_8169,N_6214,N_7401);
or U8170 (N_8170,N_7394,N_6798);
nand U8171 (N_8171,N_7306,N_6801);
or U8172 (N_8172,N_7125,N_7348);
nand U8173 (N_8173,N_6262,N_6965);
xnor U8174 (N_8174,N_6686,N_6114);
or U8175 (N_8175,N_7012,N_7088);
and U8176 (N_8176,N_7157,N_6396);
and U8177 (N_8177,N_6295,N_6751);
or U8178 (N_8178,N_6921,N_6793);
nand U8179 (N_8179,N_6019,N_7319);
xnor U8180 (N_8180,N_6920,N_6694);
and U8181 (N_8181,N_7194,N_6688);
and U8182 (N_8182,N_7096,N_6409);
xor U8183 (N_8183,N_7307,N_6577);
nor U8184 (N_8184,N_7105,N_7077);
and U8185 (N_8185,N_6597,N_7163);
nor U8186 (N_8186,N_6052,N_6869);
nand U8187 (N_8187,N_6777,N_7039);
xor U8188 (N_8188,N_7259,N_6882);
xor U8189 (N_8189,N_7364,N_6943);
or U8190 (N_8190,N_6512,N_7122);
nor U8191 (N_8191,N_6917,N_6349);
and U8192 (N_8192,N_6551,N_7304);
nor U8193 (N_8193,N_6076,N_6275);
or U8194 (N_8194,N_7339,N_7279);
and U8195 (N_8195,N_7491,N_7160);
xor U8196 (N_8196,N_7059,N_7420);
or U8197 (N_8197,N_6432,N_6980);
nor U8198 (N_8198,N_6442,N_6092);
or U8199 (N_8199,N_7037,N_6778);
nor U8200 (N_8200,N_7219,N_7496);
or U8201 (N_8201,N_6081,N_6554);
or U8202 (N_8202,N_6143,N_7495);
or U8203 (N_8203,N_6294,N_6029);
nor U8204 (N_8204,N_6068,N_6671);
or U8205 (N_8205,N_6605,N_7051);
nand U8206 (N_8206,N_6893,N_6293);
nand U8207 (N_8207,N_6043,N_7065);
xnor U8208 (N_8208,N_6074,N_6172);
nor U8209 (N_8209,N_6871,N_6956);
nand U8210 (N_8210,N_6367,N_6523);
xor U8211 (N_8211,N_6699,N_6102);
nor U8212 (N_8212,N_7079,N_6069);
nand U8213 (N_8213,N_6517,N_7085);
nand U8214 (N_8214,N_6954,N_6676);
nor U8215 (N_8215,N_7375,N_6936);
xnor U8216 (N_8216,N_6997,N_6948);
and U8217 (N_8217,N_6611,N_6125);
xor U8218 (N_8218,N_6378,N_6498);
or U8219 (N_8219,N_7068,N_6910);
nor U8220 (N_8220,N_6964,N_7148);
and U8221 (N_8221,N_6881,N_6895);
nand U8222 (N_8222,N_6268,N_6484);
or U8223 (N_8223,N_7277,N_6746);
and U8224 (N_8224,N_7231,N_7322);
nand U8225 (N_8225,N_6006,N_6271);
nand U8226 (N_8226,N_7469,N_6674);
xor U8227 (N_8227,N_6134,N_7466);
xor U8228 (N_8228,N_6420,N_7372);
nor U8229 (N_8229,N_6890,N_7121);
or U8230 (N_8230,N_6648,N_6446);
and U8231 (N_8231,N_6679,N_6147);
and U8232 (N_8232,N_7422,N_7095);
or U8233 (N_8233,N_7055,N_7202);
nor U8234 (N_8234,N_6169,N_7127);
or U8235 (N_8235,N_6872,N_6371);
nand U8236 (N_8236,N_7140,N_7384);
xnor U8237 (N_8237,N_6761,N_7416);
or U8238 (N_8238,N_6395,N_7268);
and U8239 (N_8239,N_6171,N_7254);
or U8240 (N_8240,N_6325,N_6238);
or U8241 (N_8241,N_7271,N_7424);
nor U8242 (N_8242,N_6343,N_6191);
and U8243 (N_8243,N_6714,N_6417);
and U8244 (N_8244,N_6886,N_7439);
or U8245 (N_8245,N_6469,N_6341);
and U8246 (N_8246,N_6907,N_7269);
xnor U8247 (N_8247,N_7318,N_6951);
nand U8248 (N_8248,N_7310,N_7474);
xnor U8249 (N_8249,N_6528,N_6748);
and U8250 (N_8250,N_7020,N_6562);
xor U8251 (N_8251,N_6054,N_7235);
nor U8252 (N_8252,N_6325,N_6216);
nor U8253 (N_8253,N_6241,N_6560);
nand U8254 (N_8254,N_6755,N_6020);
nor U8255 (N_8255,N_7071,N_6231);
nor U8256 (N_8256,N_6800,N_6876);
nor U8257 (N_8257,N_7088,N_6852);
nor U8258 (N_8258,N_6408,N_6930);
nor U8259 (N_8259,N_6922,N_7413);
or U8260 (N_8260,N_7028,N_6919);
and U8261 (N_8261,N_6639,N_7480);
nand U8262 (N_8262,N_6316,N_6907);
or U8263 (N_8263,N_6981,N_6496);
or U8264 (N_8264,N_6456,N_6520);
xnor U8265 (N_8265,N_6051,N_7314);
nor U8266 (N_8266,N_6455,N_6896);
xnor U8267 (N_8267,N_6062,N_6403);
nand U8268 (N_8268,N_7435,N_6796);
nor U8269 (N_8269,N_6031,N_6202);
nor U8270 (N_8270,N_7174,N_6955);
nor U8271 (N_8271,N_7464,N_6937);
and U8272 (N_8272,N_6302,N_7113);
nand U8273 (N_8273,N_6597,N_6706);
nand U8274 (N_8274,N_7331,N_7315);
nor U8275 (N_8275,N_6023,N_6385);
nor U8276 (N_8276,N_6502,N_7118);
and U8277 (N_8277,N_6154,N_7042);
nand U8278 (N_8278,N_6357,N_7028);
nand U8279 (N_8279,N_6646,N_6782);
nor U8280 (N_8280,N_6969,N_6712);
xnor U8281 (N_8281,N_6986,N_6067);
nor U8282 (N_8282,N_6300,N_7116);
nand U8283 (N_8283,N_6830,N_6963);
xnor U8284 (N_8284,N_6739,N_6037);
and U8285 (N_8285,N_7003,N_6328);
nand U8286 (N_8286,N_6521,N_7305);
nand U8287 (N_8287,N_6280,N_6099);
nand U8288 (N_8288,N_6449,N_6230);
nand U8289 (N_8289,N_6437,N_7048);
nand U8290 (N_8290,N_6968,N_7458);
and U8291 (N_8291,N_6882,N_7431);
and U8292 (N_8292,N_6218,N_7393);
or U8293 (N_8293,N_7398,N_6124);
xor U8294 (N_8294,N_6842,N_6930);
xnor U8295 (N_8295,N_6998,N_6939);
nand U8296 (N_8296,N_7196,N_7215);
nor U8297 (N_8297,N_7430,N_7272);
and U8298 (N_8298,N_6078,N_7484);
nand U8299 (N_8299,N_6000,N_7120);
nor U8300 (N_8300,N_6190,N_6247);
or U8301 (N_8301,N_6784,N_6102);
or U8302 (N_8302,N_7147,N_6463);
xor U8303 (N_8303,N_6584,N_6216);
or U8304 (N_8304,N_7092,N_7182);
or U8305 (N_8305,N_6820,N_6521);
and U8306 (N_8306,N_6326,N_6445);
and U8307 (N_8307,N_6241,N_6561);
xnor U8308 (N_8308,N_6486,N_6789);
xnor U8309 (N_8309,N_7051,N_6310);
or U8310 (N_8310,N_6375,N_6135);
nand U8311 (N_8311,N_6637,N_7420);
or U8312 (N_8312,N_6876,N_6981);
nor U8313 (N_8313,N_6874,N_7237);
nand U8314 (N_8314,N_6850,N_7439);
nand U8315 (N_8315,N_6112,N_7345);
or U8316 (N_8316,N_6822,N_6845);
xor U8317 (N_8317,N_7299,N_6727);
nor U8318 (N_8318,N_6991,N_6853);
or U8319 (N_8319,N_6850,N_7312);
or U8320 (N_8320,N_6588,N_7430);
nor U8321 (N_8321,N_7453,N_6529);
xnor U8322 (N_8322,N_6079,N_6464);
nand U8323 (N_8323,N_7177,N_7131);
or U8324 (N_8324,N_6340,N_6914);
nand U8325 (N_8325,N_7493,N_6603);
and U8326 (N_8326,N_6363,N_7129);
nor U8327 (N_8327,N_6987,N_6611);
or U8328 (N_8328,N_7128,N_6908);
or U8329 (N_8329,N_7077,N_6462);
nor U8330 (N_8330,N_6977,N_7186);
xor U8331 (N_8331,N_6456,N_6387);
xnor U8332 (N_8332,N_7140,N_6344);
nor U8333 (N_8333,N_7217,N_6387);
and U8334 (N_8334,N_6359,N_7124);
xor U8335 (N_8335,N_6957,N_6173);
nand U8336 (N_8336,N_6502,N_6865);
xor U8337 (N_8337,N_6542,N_7088);
and U8338 (N_8338,N_7340,N_7498);
xnor U8339 (N_8339,N_7363,N_7354);
or U8340 (N_8340,N_6998,N_6778);
or U8341 (N_8341,N_7468,N_6946);
or U8342 (N_8342,N_6746,N_6047);
or U8343 (N_8343,N_7407,N_6551);
or U8344 (N_8344,N_6101,N_7191);
or U8345 (N_8345,N_7021,N_6190);
xor U8346 (N_8346,N_7408,N_6710);
nand U8347 (N_8347,N_6829,N_7424);
or U8348 (N_8348,N_6852,N_7241);
nand U8349 (N_8349,N_6485,N_6598);
nand U8350 (N_8350,N_7387,N_6904);
or U8351 (N_8351,N_6898,N_6206);
nand U8352 (N_8352,N_6440,N_6759);
and U8353 (N_8353,N_6888,N_6127);
nor U8354 (N_8354,N_6205,N_6231);
and U8355 (N_8355,N_6431,N_7262);
and U8356 (N_8356,N_6982,N_7291);
or U8357 (N_8357,N_7380,N_6445);
xnor U8358 (N_8358,N_7427,N_6102);
nand U8359 (N_8359,N_7447,N_6389);
nor U8360 (N_8360,N_6635,N_6420);
or U8361 (N_8361,N_7191,N_6852);
or U8362 (N_8362,N_6766,N_6846);
xnor U8363 (N_8363,N_7234,N_7143);
xor U8364 (N_8364,N_6273,N_7162);
and U8365 (N_8365,N_6993,N_6409);
xnor U8366 (N_8366,N_6341,N_6373);
xor U8367 (N_8367,N_6439,N_7317);
or U8368 (N_8368,N_7123,N_6610);
nand U8369 (N_8369,N_6935,N_6712);
nor U8370 (N_8370,N_6742,N_7029);
and U8371 (N_8371,N_6615,N_6479);
or U8372 (N_8372,N_6435,N_7044);
and U8373 (N_8373,N_6306,N_6246);
nand U8374 (N_8374,N_6693,N_6712);
nand U8375 (N_8375,N_6311,N_7386);
xnor U8376 (N_8376,N_7245,N_7201);
xor U8377 (N_8377,N_6413,N_7201);
or U8378 (N_8378,N_7068,N_7341);
nor U8379 (N_8379,N_7287,N_6811);
and U8380 (N_8380,N_6594,N_6709);
xnor U8381 (N_8381,N_7149,N_6714);
nand U8382 (N_8382,N_6488,N_6985);
nor U8383 (N_8383,N_7439,N_6695);
and U8384 (N_8384,N_7173,N_7164);
nand U8385 (N_8385,N_7045,N_6323);
xor U8386 (N_8386,N_6020,N_6247);
xnor U8387 (N_8387,N_6738,N_6430);
nor U8388 (N_8388,N_7074,N_6173);
and U8389 (N_8389,N_6172,N_6043);
xnor U8390 (N_8390,N_6950,N_6258);
nor U8391 (N_8391,N_7319,N_7443);
or U8392 (N_8392,N_6821,N_6645);
nand U8393 (N_8393,N_7165,N_6156);
or U8394 (N_8394,N_6846,N_6449);
nor U8395 (N_8395,N_6612,N_6270);
nand U8396 (N_8396,N_6725,N_7255);
xnor U8397 (N_8397,N_7083,N_7340);
or U8398 (N_8398,N_7276,N_6950);
xnor U8399 (N_8399,N_6830,N_7060);
xnor U8400 (N_8400,N_7290,N_7175);
nand U8401 (N_8401,N_6311,N_6597);
or U8402 (N_8402,N_6391,N_6292);
xor U8403 (N_8403,N_6826,N_7020);
nor U8404 (N_8404,N_6177,N_6606);
and U8405 (N_8405,N_6391,N_6036);
nand U8406 (N_8406,N_6754,N_7182);
nand U8407 (N_8407,N_7266,N_6493);
nand U8408 (N_8408,N_7380,N_6081);
and U8409 (N_8409,N_6272,N_6956);
or U8410 (N_8410,N_6410,N_6434);
nand U8411 (N_8411,N_6885,N_6732);
xor U8412 (N_8412,N_6417,N_6376);
nor U8413 (N_8413,N_6943,N_6006);
xnor U8414 (N_8414,N_7385,N_6892);
nand U8415 (N_8415,N_6518,N_7468);
nand U8416 (N_8416,N_7099,N_7136);
nand U8417 (N_8417,N_6962,N_7321);
xor U8418 (N_8418,N_6130,N_6936);
or U8419 (N_8419,N_7393,N_6293);
xnor U8420 (N_8420,N_6545,N_6778);
or U8421 (N_8421,N_6410,N_6861);
xnor U8422 (N_8422,N_6390,N_6060);
or U8423 (N_8423,N_6832,N_6379);
nor U8424 (N_8424,N_6994,N_6799);
or U8425 (N_8425,N_6607,N_6881);
nand U8426 (N_8426,N_7170,N_7387);
xor U8427 (N_8427,N_6355,N_6256);
and U8428 (N_8428,N_6327,N_6950);
nand U8429 (N_8429,N_6161,N_7163);
and U8430 (N_8430,N_7265,N_6782);
nand U8431 (N_8431,N_7171,N_6714);
or U8432 (N_8432,N_6868,N_7038);
and U8433 (N_8433,N_6451,N_7363);
xor U8434 (N_8434,N_6119,N_7097);
nand U8435 (N_8435,N_6442,N_6866);
nand U8436 (N_8436,N_7216,N_6614);
xor U8437 (N_8437,N_6805,N_6146);
nand U8438 (N_8438,N_7328,N_6170);
or U8439 (N_8439,N_6873,N_6150);
and U8440 (N_8440,N_6201,N_6332);
or U8441 (N_8441,N_6033,N_6322);
nand U8442 (N_8442,N_6871,N_7416);
xor U8443 (N_8443,N_7355,N_6411);
xor U8444 (N_8444,N_6951,N_6457);
and U8445 (N_8445,N_6179,N_6574);
xor U8446 (N_8446,N_6998,N_7225);
or U8447 (N_8447,N_6205,N_6724);
and U8448 (N_8448,N_7361,N_6830);
xor U8449 (N_8449,N_6425,N_6699);
nand U8450 (N_8450,N_7307,N_7468);
and U8451 (N_8451,N_6507,N_6636);
xnor U8452 (N_8452,N_7035,N_6098);
nor U8453 (N_8453,N_6175,N_7085);
nand U8454 (N_8454,N_7210,N_6666);
or U8455 (N_8455,N_6612,N_6920);
nand U8456 (N_8456,N_7152,N_6082);
nand U8457 (N_8457,N_6744,N_7402);
and U8458 (N_8458,N_6835,N_6912);
and U8459 (N_8459,N_7369,N_6274);
nor U8460 (N_8460,N_6493,N_6963);
or U8461 (N_8461,N_7291,N_6598);
xor U8462 (N_8462,N_6358,N_6806);
xnor U8463 (N_8463,N_7308,N_6980);
xnor U8464 (N_8464,N_6344,N_7116);
nor U8465 (N_8465,N_7339,N_6297);
or U8466 (N_8466,N_7349,N_6940);
or U8467 (N_8467,N_7120,N_6215);
or U8468 (N_8468,N_6482,N_6366);
nand U8469 (N_8469,N_6813,N_7113);
and U8470 (N_8470,N_6415,N_7440);
nor U8471 (N_8471,N_6543,N_7398);
or U8472 (N_8472,N_6376,N_6329);
and U8473 (N_8473,N_6330,N_6078);
or U8474 (N_8474,N_6624,N_6389);
nand U8475 (N_8475,N_7465,N_7170);
nor U8476 (N_8476,N_6283,N_6866);
xor U8477 (N_8477,N_6012,N_7257);
nand U8478 (N_8478,N_7395,N_6711);
or U8479 (N_8479,N_7435,N_6224);
xnor U8480 (N_8480,N_6980,N_6403);
xor U8481 (N_8481,N_7249,N_6754);
and U8482 (N_8482,N_6427,N_6746);
nand U8483 (N_8483,N_6803,N_6120);
xnor U8484 (N_8484,N_6853,N_7248);
and U8485 (N_8485,N_6626,N_6679);
or U8486 (N_8486,N_6434,N_7265);
xor U8487 (N_8487,N_7356,N_7021);
nand U8488 (N_8488,N_7113,N_7491);
and U8489 (N_8489,N_6179,N_6518);
xnor U8490 (N_8490,N_7253,N_6377);
xor U8491 (N_8491,N_6416,N_7117);
and U8492 (N_8492,N_7404,N_6512);
or U8493 (N_8493,N_7133,N_7251);
nand U8494 (N_8494,N_6191,N_6622);
nor U8495 (N_8495,N_6576,N_6583);
nor U8496 (N_8496,N_7212,N_6447);
nand U8497 (N_8497,N_7287,N_6593);
nand U8498 (N_8498,N_6002,N_6705);
or U8499 (N_8499,N_6797,N_6669);
nor U8500 (N_8500,N_6482,N_7213);
or U8501 (N_8501,N_7480,N_6330);
xor U8502 (N_8502,N_6284,N_6153);
or U8503 (N_8503,N_6895,N_7093);
nor U8504 (N_8504,N_6670,N_7267);
or U8505 (N_8505,N_6483,N_6603);
nor U8506 (N_8506,N_6467,N_6136);
and U8507 (N_8507,N_6205,N_6621);
xor U8508 (N_8508,N_7133,N_6855);
or U8509 (N_8509,N_7397,N_7277);
or U8510 (N_8510,N_6647,N_7180);
or U8511 (N_8511,N_6330,N_7041);
and U8512 (N_8512,N_6037,N_7434);
and U8513 (N_8513,N_7256,N_6880);
xnor U8514 (N_8514,N_6829,N_6426);
or U8515 (N_8515,N_6030,N_6074);
nor U8516 (N_8516,N_6469,N_6500);
nand U8517 (N_8517,N_6426,N_7494);
and U8518 (N_8518,N_6802,N_6720);
nor U8519 (N_8519,N_6045,N_6619);
or U8520 (N_8520,N_6844,N_6538);
xor U8521 (N_8521,N_6940,N_6562);
and U8522 (N_8522,N_7212,N_7077);
and U8523 (N_8523,N_7129,N_6413);
nand U8524 (N_8524,N_6950,N_6012);
nand U8525 (N_8525,N_6753,N_7357);
and U8526 (N_8526,N_6129,N_6327);
and U8527 (N_8527,N_7382,N_6749);
nand U8528 (N_8528,N_6034,N_6691);
xor U8529 (N_8529,N_6138,N_6977);
nand U8530 (N_8530,N_6728,N_6644);
xor U8531 (N_8531,N_7215,N_6828);
xnor U8532 (N_8532,N_6133,N_6255);
nor U8533 (N_8533,N_7489,N_7279);
nand U8534 (N_8534,N_6275,N_6933);
nor U8535 (N_8535,N_6505,N_6341);
nand U8536 (N_8536,N_6656,N_6607);
nand U8537 (N_8537,N_6845,N_6912);
and U8538 (N_8538,N_7410,N_6446);
and U8539 (N_8539,N_6976,N_6255);
nor U8540 (N_8540,N_7076,N_6106);
nand U8541 (N_8541,N_6170,N_7279);
nor U8542 (N_8542,N_6343,N_6960);
nand U8543 (N_8543,N_6227,N_7153);
and U8544 (N_8544,N_6712,N_6157);
nand U8545 (N_8545,N_7131,N_7031);
nand U8546 (N_8546,N_7198,N_6729);
or U8547 (N_8547,N_6982,N_7422);
nand U8548 (N_8548,N_6939,N_6226);
or U8549 (N_8549,N_6036,N_7141);
nand U8550 (N_8550,N_6611,N_7285);
and U8551 (N_8551,N_7111,N_6140);
nor U8552 (N_8552,N_6392,N_6068);
nor U8553 (N_8553,N_7096,N_6406);
nor U8554 (N_8554,N_6628,N_6573);
nand U8555 (N_8555,N_6663,N_6717);
nor U8556 (N_8556,N_6638,N_6020);
and U8557 (N_8557,N_6970,N_6546);
and U8558 (N_8558,N_6668,N_6835);
xnor U8559 (N_8559,N_6456,N_6557);
xnor U8560 (N_8560,N_6668,N_6145);
xnor U8561 (N_8561,N_6648,N_6451);
xnor U8562 (N_8562,N_6242,N_7258);
nor U8563 (N_8563,N_7070,N_6881);
nand U8564 (N_8564,N_6542,N_6580);
nor U8565 (N_8565,N_6069,N_7418);
nand U8566 (N_8566,N_7390,N_6193);
and U8567 (N_8567,N_7436,N_7001);
nand U8568 (N_8568,N_6370,N_7154);
xnor U8569 (N_8569,N_6262,N_6718);
nor U8570 (N_8570,N_7221,N_7039);
nand U8571 (N_8571,N_6277,N_6775);
nor U8572 (N_8572,N_7253,N_7040);
nand U8573 (N_8573,N_6191,N_7020);
xnor U8574 (N_8574,N_6512,N_6241);
xnor U8575 (N_8575,N_7156,N_6386);
nor U8576 (N_8576,N_7200,N_6715);
and U8577 (N_8577,N_6255,N_6449);
xnor U8578 (N_8578,N_6748,N_7254);
nand U8579 (N_8579,N_6003,N_6702);
and U8580 (N_8580,N_7246,N_6904);
and U8581 (N_8581,N_7432,N_6486);
or U8582 (N_8582,N_7043,N_6961);
and U8583 (N_8583,N_6307,N_7027);
nor U8584 (N_8584,N_6383,N_7486);
or U8585 (N_8585,N_7484,N_6848);
or U8586 (N_8586,N_6137,N_6544);
nand U8587 (N_8587,N_6084,N_7235);
nand U8588 (N_8588,N_7065,N_6660);
or U8589 (N_8589,N_6751,N_6335);
xor U8590 (N_8590,N_6934,N_7311);
nor U8591 (N_8591,N_7040,N_6945);
nor U8592 (N_8592,N_6011,N_7099);
nand U8593 (N_8593,N_6087,N_6717);
nor U8594 (N_8594,N_6089,N_6251);
and U8595 (N_8595,N_6074,N_6972);
or U8596 (N_8596,N_6659,N_6025);
xnor U8597 (N_8597,N_6530,N_6818);
or U8598 (N_8598,N_6927,N_6945);
or U8599 (N_8599,N_6092,N_7429);
or U8600 (N_8600,N_7221,N_7193);
nor U8601 (N_8601,N_6529,N_6638);
and U8602 (N_8602,N_6583,N_6178);
nor U8603 (N_8603,N_6897,N_7222);
or U8604 (N_8604,N_7034,N_7242);
or U8605 (N_8605,N_6015,N_6842);
and U8606 (N_8606,N_6260,N_6153);
nand U8607 (N_8607,N_6096,N_6209);
nand U8608 (N_8608,N_6552,N_7480);
and U8609 (N_8609,N_6555,N_6492);
and U8610 (N_8610,N_6523,N_7337);
nor U8611 (N_8611,N_6103,N_6832);
nand U8612 (N_8612,N_6008,N_6917);
and U8613 (N_8613,N_6700,N_6226);
nor U8614 (N_8614,N_7221,N_6031);
or U8615 (N_8615,N_6719,N_6933);
nand U8616 (N_8616,N_6832,N_6615);
xor U8617 (N_8617,N_6286,N_6002);
or U8618 (N_8618,N_7497,N_6543);
or U8619 (N_8619,N_6810,N_6859);
xor U8620 (N_8620,N_6768,N_7020);
xnor U8621 (N_8621,N_7270,N_7392);
or U8622 (N_8622,N_6128,N_6928);
and U8623 (N_8623,N_7467,N_6754);
nor U8624 (N_8624,N_7183,N_6551);
and U8625 (N_8625,N_6172,N_6382);
or U8626 (N_8626,N_6971,N_6229);
nand U8627 (N_8627,N_7206,N_6282);
and U8628 (N_8628,N_6391,N_6575);
nand U8629 (N_8629,N_6130,N_7127);
and U8630 (N_8630,N_7269,N_6930);
nand U8631 (N_8631,N_6616,N_6931);
and U8632 (N_8632,N_6446,N_7207);
and U8633 (N_8633,N_7448,N_6067);
nand U8634 (N_8634,N_6439,N_7257);
nor U8635 (N_8635,N_6688,N_6905);
nand U8636 (N_8636,N_6116,N_6751);
nand U8637 (N_8637,N_6627,N_7463);
nor U8638 (N_8638,N_6815,N_6935);
and U8639 (N_8639,N_6834,N_6040);
or U8640 (N_8640,N_7022,N_7113);
or U8641 (N_8641,N_7070,N_6032);
nor U8642 (N_8642,N_6975,N_6855);
nand U8643 (N_8643,N_6799,N_7011);
and U8644 (N_8644,N_7344,N_6863);
nand U8645 (N_8645,N_6003,N_6966);
nand U8646 (N_8646,N_6713,N_6565);
nor U8647 (N_8647,N_6294,N_6207);
nor U8648 (N_8648,N_7277,N_6017);
nand U8649 (N_8649,N_6928,N_6765);
and U8650 (N_8650,N_6063,N_7206);
and U8651 (N_8651,N_7232,N_7265);
and U8652 (N_8652,N_6922,N_7139);
xor U8653 (N_8653,N_7385,N_6152);
nand U8654 (N_8654,N_6567,N_6356);
nor U8655 (N_8655,N_6395,N_6872);
and U8656 (N_8656,N_6306,N_7200);
nand U8657 (N_8657,N_6870,N_6603);
or U8658 (N_8658,N_7285,N_7219);
nand U8659 (N_8659,N_7077,N_7029);
nand U8660 (N_8660,N_7181,N_6043);
xor U8661 (N_8661,N_7141,N_7381);
nand U8662 (N_8662,N_6772,N_7003);
xnor U8663 (N_8663,N_6215,N_6405);
nand U8664 (N_8664,N_7159,N_7049);
and U8665 (N_8665,N_6796,N_6715);
or U8666 (N_8666,N_6221,N_6561);
nor U8667 (N_8667,N_7128,N_6566);
nor U8668 (N_8668,N_6140,N_6118);
and U8669 (N_8669,N_7067,N_6884);
nand U8670 (N_8670,N_6578,N_7208);
and U8671 (N_8671,N_7037,N_7286);
nor U8672 (N_8672,N_6881,N_7088);
or U8673 (N_8673,N_6366,N_6941);
nor U8674 (N_8674,N_6883,N_6232);
and U8675 (N_8675,N_6529,N_6659);
or U8676 (N_8676,N_6204,N_6807);
nand U8677 (N_8677,N_7055,N_6152);
and U8678 (N_8678,N_7385,N_6161);
and U8679 (N_8679,N_7410,N_6825);
nand U8680 (N_8680,N_6931,N_6078);
xnor U8681 (N_8681,N_6712,N_6748);
or U8682 (N_8682,N_6732,N_7431);
nand U8683 (N_8683,N_6760,N_6715);
and U8684 (N_8684,N_6077,N_6369);
and U8685 (N_8685,N_7318,N_6443);
and U8686 (N_8686,N_7193,N_7249);
nor U8687 (N_8687,N_6650,N_7381);
nand U8688 (N_8688,N_6868,N_7264);
xor U8689 (N_8689,N_7320,N_6748);
or U8690 (N_8690,N_6501,N_7253);
xnor U8691 (N_8691,N_6236,N_6168);
or U8692 (N_8692,N_7393,N_7114);
and U8693 (N_8693,N_7143,N_7024);
nor U8694 (N_8694,N_7034,N_6113);
or U8695 (N_8695,N_6001,N_7352);
xor U8696 (N_8696,N_6215,N_6518);
and U8697 (N_8697,N_6037,N_6270);
nand U8698 (N_8698,N_7135,N_6902);
and U8699 (N_8699,N_6011,N_6184);
and U8700 (N_8700,N_7200,N_6871);
nand U8701 (N_8701,N_6046,N_6126);
xor U8702 (N_8702,N_7328,N_7293);
nand U8703 (N_8703,N_7474,N_6056);
xnor U8704 (N_8704,N_6934,N_7205);
xnor U8705 (N_8705,N_7180,N_6168);
xnor U8706 (N_8706,N_6124,N_7129);
or U8707 (N_8707,N_6475,N_7101);
nor U8708 (N_8708,N_6066,N_6982);
and U8709 (N_8709,N_6043,N_7394);
xnor U8710 (N_8710,N_7439,N_6037);
nand U8711 (N_8711,N_6700,N_6746);
nand U8712 (N_8712,N_7301,N_7420);
and U8713 (N_8713,N_7424,N_6149);
nand U8714 (N_8714,N_6477,N_6888);
or U8715 (N_8715,N_6585,N_6881);
or U8716 (N_8716,N_6157,N_7419);
and U8717 (N_8717,N_6244,N_7465);
or U8718 (N_8718,N_6402,N_6631);
nor U8719 (N_8719,N_6335,N_6843);
nand U8720 (N_8720,N_6097,N_7320);
xnor U8721 (N_8721,N_6349,N_7185);
or U8722 (N_8722,N_6266,N_7467);
nor U8723 (N_8723,N_7425,N_6805);
nand U8724 (N_8724,N_7313,N_7022);
nand U8725 (N_8725,N_7028,N_7415);
nor U8726 (N_8726,N_6643,N_7128);
xor U8727 (N_8727,N_6541,N_7239);
xor U8728 (N_8728,N_7066,N_6408);
xor U8729 (N_8729,N_6634,N_6902);
nand U8730 (N_8730,N_7068,N_7272);
or U8731 (N_8731,N_6762,N_7361);
nor U8732 (N_8732,N_6727,N_6127);
nor U8733 (N_8733,N_6447,N_6353);
nand U8734 (N_8734,N_6393,N_6246);
nor U8735 (N_8735,N_6005,N_6619);
xnor U8736 (N_8736,N_6151,N_6233);
xnor U8737 (N_8737,N_6644,N_7423);
nor U8738 (N_8738,N_6358,N_7324);
xor U8739 (N_8739,N_6477,N_7042);
and U8740 (N_8740,N_7017,N_6009);
nor U8741 (N_8741,N_7443,N_6802);
xnor U8742 (N_8742,N_6713,N_7156);
or U8743 (N_8743,N_6695,N_6003);
xor U8744 (N_8744,N_6109,N_7163);
and U8745 (N_8745,N_7009,N_6856);
or U8746 (N_8746,N_6801,N_6517);
xor U8747 (N_8747,N_6637,N_6320);
or U8748 (N_8748,N_6887,N_7318);
or U8749 (N_8749,N_7113,N_7325);
xor U8750 (N_8750,N_6171,N_6073);
nor U8751 (N_8751,N_6289,N_6966);
xor U8752 (N_8752,N_6789,N_6889);
xor U8753 (N_8753,N_6336,N_7105);
nor U8754 (N_8754,N_6591,N_6483);
and U8755 (N_8755,N_6179,N_7208);
and U8756 (N_8756,N_6463,N_6813);
xor U8757 (N_8757,N_6829,N_6357);
xnor U8758 (N_8758,N_6137,N_7212);
and U8759 (N_8759,N_6661,N_7433);
or U8760 (N_8760,N_6206,N_6134);
or U8761 (N_8761,N_6507,N_6887);
or U8762 (N_8762,N_6591,N_6127);
nand U8763 (N_8763,N_6171,N_7187);
nand U8764 (N_8764,N_6521,N_7224);
xnor U8765 (N_8765,N_6695,N_6700);
or U8766 (N_8766,N_6946,N_6020);
nand U8767 (N_8767,N_6534,N_6854);
nand U8768 (N_8768,N_6433,N_6404);
and U8769 (N_8769,N_7328,N_7179);
and U8770 (N_8770,N_7245,N_7069);
xnor U8771 (N_8771,N_6950,N_7011);
xnor U8772 (N_8772,N_7153,N_7105);
xnor U8773 (N_8773,N_6951,N_7102);
or U8774 (N_8774,N_7123,N_6820);
or U8775 (N_8775,N_6020,N_6276);
and U8776 (N_8776,N_6101,N_6232);
and U8777 (N_8777,N_7436,N_6619);
nand U8778 (N_8778,N_7081,N_6397);
nand U8779 (N_8779,N_7218,N_7052);
and U8780 (N_8780,N_6422,N_7164);
or U8781 (N_8781,N_7195,N_7434);
xnor U8782 (N_8782,N_7435,N_6034);
xnor U8783 (N_8783,N_7073,N_7008);
xnor U8784 (N_8784,N_6962,N_6658);
nor U8785 (N_8785,N_7216,N_7424);
nor U8786 (N_8786,N_6009,N_7425);
and U8787 (N_8787,N_7162,N_7155);
xor U8788 (N_8788,N_7359,N_7295);
nor U8789 (N_8789,N_7069,N_7441);
nor U8790 (N_8790,N_6735,N_6255);
xor U8791 (N_8791,N_6270,N_7430);
nand U8792 (N_8792,N_6047,N_6672);
xor U8793 (N_8793,N_6343,N_6356);
nor U8794 (N_8794,N_6193,N_6100);
nand U8795 (N_8795,N_6734,N_6892);
and U8796 (N_8796,N_6310,N_6814);
nor U8797 (N_8797,N_7139,N_7238);
and U8798 (N_8798,N_7283,N_6956);
nor U8799 (N_8799,N_7130,N_7406);
nor U8800 (N_8800,N_6530,N_6654);
nor U8801 (N_8801,N_6057,N_6469);
or U8802 (N_8802,N_7151,N_7402);
xnor U8803 (N_8803,N_7483,N_6233);
and U8804 (N_8804,N_7468,N_6908);
nor U8805 (N_8805,N_7286,N_7495);
and U8806 (N_8806,N_6407,N_6541);
or U8807 (N_8807,N_6035,N_6046);
nand U8808 (N_8808,N_7400,N_6186);
nor U8809 (N_8809,N_6927,N_6503);
and U8810 (N_8810,N_6236,N_6994);
nor U8811 (N_8811,N_6878,N_6843);
xor U8812 (N_8812,N_6751,N_6538);
nor U8813 (N_8813,N_6108,N_7496);
or U8814 (N_8814,N_6810,N_6337);
xnor U8815 (N_8815,N_6671,N_6434);
or U8816 (N_8816,N_6495,N_6684);
xor U8817 (N_8817,N_6113,N_7043);
nor U8818 (N_8818,N_6559,N_6516);
or U8819 (N_8819,N_6116,N_6309);
xor U8820 (N_8820,N_6327,N_7343);
xor U8821 (N_8821,N_6625,N_7091);
nor U8822 (N_8822,N_6064,N_6084);
and U8823 (N_8823,N_6621,N_6352);
or U8824 (N_8824,N_6591,N_7394);
xor U8825 (N_8825,N_7377,N_6872);
nand U8826 (N_8826,N_7161,N_7272);
or U8827 (N_8827,N_6429,N_7274);
nor U8828 (N_8828,N_6235,N_7495);
nor U8829 (N_8829,N_6213,N_6687);
nand U8830 (N_8830,N_6900,N_6742);
and U8831 (N_8831,N_6237,N_7486);
or U8832 (N_8832,N_7319,N_7217);
nand U8833 (N_8833,N_6480,N_6073);
and U8834 (N_8834,N_6568,N_6629);
or U8835 (N_8835,N_6596,N_7031);
or U8836 (N_8836,N_6137,N_6577);
nor U8837 (N_8837,N_6129,N_7341);
xnor U8838 (N_8838,N_6458,N_7491);
and U8839 (N_8839,N_7281,N_7428);
nand U8840 (N_8840,N_6930,N_6428);
and U8841 (N_8841,N_6750,N_6733);
or U8842 (N_8842,N_7354,N_6453);
and U8843 (N_8843,N_7402,N_6862);
and U8844 (N_8844,N_6645,N_7150);
nand U8845 (N_8845,N_6068,N_7050);
nand U8846 (N_8846,N_6047,N_6397);
or U8847 (N_8847,N_6895,N_6528);
and U8848 (N_8848,N_6435,N_6531);
xor U8849 (N_8849,N_6083,N_6115);
nand U8850 (N_8850,N_6992,N_7127);
and U8851 (N_8851,N_6178,N_6134);
nor U8852 (N_8852,N_6617,N_6086);
and U8853 (N_8853,N_7332,N_6818);
nand U8854 (N_8854,N_7085,N_7397);
nor U8855 (N_8855,N_7352,N_7495);
and U8856 (N_8856,N_6590,N_7130);
or U8857 (N_8857,N_6850,N_7277);
nand U8858 (N_8858,N_7463,N_6122);
nand U8859 (N_8859,N_7445,N_7202);
nor U8860 (N_8860,N_7387,N_7414);
or U8861 (N_8861,N_6693,N_7022);
nand U8862 (N_8862,N_7392,N_6054);
and U8863 (N_8863,N_6010,N_6154);
nor U8864 (N_8864,N_6169,N_6404);
nand U8865 (N_8865,N_7320,N_7072);
or U8866 (N_8866,N_6194,N_6061);
nand U8867 (N_8867,N_6871,N_6635);
nor U8868 (N_8868,N_7169,N_7453);
nor U8869 (N_8869,N_6613,N_6991);
or U8870 (N_8870,N_6354,N_6802);
nor U8871 (N_8871,N_6892,N_6351);
or U8872 (N_8872,N_6619,N_6087);
or U8873 (N_8873,N_6346,N_7033);
and U8874 (N_8874,N_6652,N_6327);
nand U8875 (N_8875,N_7206,N_7171);
or U8876 (N_8876,N_7103,N_6717);
or U8877 (N_8877,N_6133,N_6617);
or U8878 (N_8878,N_6355,N_6715);
nand U8879 (N_8879,N_6969,N_7150);
or U8880 (N_8880,N_6333,N_6315);
nor U8881 (N_8881,N_7105,N_6345);
or U8882 (N_8882,N_7266,N_6297);
and U8883 (N_8883,N_7390,N_7252);
nand U8884 (N_8884,N_6792,N_6039);
nor U8885 (N_8885,N_7092,N_6785);
or U8886 (N_8886,N_6726,N_7176);
nand U8887 (N_8887,N_6402,N_6901);
nor U8888 (N_8888,N_6316,N_6662);
or U8889 (N_8889,N_6565,N_7427);
or U8890 (N_8890,N_7391,N_6803);
and U8891 (N_8891,N_7023,N_7163);
or U8892 (N_8892,N_6663,N_6218);
nand U8893 (N_8893,N_6210,N_7249);
nor U8894 (N_8894,N_7134,N_6444);
nor U8895 (N_8895,N_6503,N_7065);
nor U8896 (N_8896,N_6717,N_7153);
and U8897 (N_8897,N_7139,N_6326);
xor U8898 (N_8898,N_7353,N_6589);
xnor U8899 (N_8899,N_7487,N_7051);
nor U8900 (N_8900,N_6986,N_7283);
or U8901 (N_8901,N_6775,N_6969);
xor U8902 (N_8902,N_6107,N_6909);
nor U8903 (N_8903,N_6696,N_6047);
xor U8904 (N_8904,N_6351,N_7116);
and U8905 (N_8905,N_6759,N_7374);
nand U8906 (N_8906,N_6725,N_6077);
nand U8907 (N_8907,N_6629,N_6550);
nor U8908 (N_8908,N_7033,N_6257);
xnor U8909 (N_8909,N_6458,N_6064);
nand U8910 (N_8910,N_6065,N_6607);
or U8911 (N_8911,N_6003,N_6197);
and U8912 (N_8912,N_6903,N_7341);
nor U8913 (N_8913,N_6799,N_6331);
nor U8914 (N_8914,N_7419,N_6234);
nor U8915 (N_8915,N_6586,N_7236);
and U8916 (N_8916,N_7225,N_6517);
nor U8917 (N_8917,N_6657,N_6471);
xor U8918 (N_8918,N_7355,N_6867);
and U8919 (N_8919,N_6075,N_6990);
and U8920 (N_8920,N_6779,N_7047);
or U8921 (N_8921,N_7251,N_6417);
and U8922 (N_8922,N_6451,N_7254);
xnor U8923 (N_8923,N_6621,N_7494);
nand U8924 (N_8924,N_6794,N_6304);
nand U8925 (N_8925,N_7110,N_6662);
xor U8926 (N_8926,N_6241,N_7114);
or U8927 (N_8927,N_6143,N_6342);
xnor U8928 (N_8928,N_6652,N_7388);
nor U8929 (N_8929,N_7342,N_6873);
nor U8930 (N_8930,N_6098,N_6041);
nand U8931 (N_8931,N_6477,N_6572);
or U8932 (N_8932,N_6345,N_6480);
nor U8933 (N_8933,N_7135,N_6227);
xnor U8934 (N_8934,N_7397,N_6533);
or U8935 (N_8935,N_6873,N_7099);
nor U8936 (N_8936,N_6869,N_7441);
or U8937 (N_8937,N_6102,N_7397);
xor U8938 (N_8938,N_6034,N_7145);
and U8939 (N_8939,N_7118,N_6799);
xnor U8940 (N_8940,N_6752,N_6062);
and U8941 (N_8941,N_6223,N_7493);
and U8942 (N_8942,N_6433,N_6170);
xnor U8943 (N_8943,N_7018,N_7487);
or U8944 (N_8944,N_7332,N_7211);
nand U8945 (N_8945,N_6252,N_6950);
nand U8946 (N_8946,N_6564,N_6936);
xnor U8947 (N_8947,N_6059,N_6817);
and U8948 (N_8948,N_7213,N_7297);
or U8949 (N_8949,N_6726,N_6894);
nor U8950 (N_8950,N_6595,N_6954);
or U8951 (N_8951,N_7201,N_6119);
or U8952 (N_8952,N_6814,N_7063);
nand U8953 (N_8953,N_6254,N_6069);
and U8954 (N_8954,N_6460,N_6088);
and U8955 (N_8955,N_6626,N_6640);
or U8956 (N_8956,N_6767,N_7384);
and U8957 (N_8957,N_6521,N_7201);
nand U8958 (N_8958,N_7082,N_7196);
or U8959 (N_8959,N_6486,N_7009);
and U8960 (N_8960,N_6017,N_7450);
nand U8961 (N_8961,N_6770,N_7387);
nor U8962 (N_8962,N_7491,N_6363);
and U8963 (N_8963,N_7245,N_7255);
or U8964 (N_8964,N_6486,N_7435);
nor U8965 (N_8965,N_7042,N_6957);
nor U8966 (N_8966,N_6099,N_6863);
nor U8967 (N_8967,N_6242,N_6332);
nand U8968 (N_8968,N_7044,N_6131);
nand U8969 (N_8969,N_6041,N_6880);
and U8970 (N_8970,N_6657,N_7161);
xnor U8971 (N_8971,N_6075,N_6093);
nor U8972 (N_8972,N_6280,N_6943);
nand U8973 (N_8973,N_6047,N_6396);
and U8974 (N_8974,N_6835,N_7176);
xnor U8975 (N_8975,N_6451,N_6733);
and U8976 (N_8976,N_6508,N_6380);
and U8977 (N_8977,N_6231,N_6182);
and U8978 (N_8978,N_6664,N_6127);
or U8979 (N_8979,N_6420,N_7075);
and U8980 (N_8980,N_6466,N_6561);
nor U8981 (N_8981,N_6264,N_7485);
nor U8982 (N_8982,N_6786,N_7259);
xor U8983 (N_8983,N_7314,N_6238);
xnor U8984 (N_8984,N_6334,N_6301);
or U8985 (N_8985,N_6029,N_7119);
nand U8986 (N_8986,N_7355,N_6200);
or U8987 (N_8987,N_6644,N_6957);
xor U8988 (N_8988,N_6124,N_6724);
and U8989 (N_8989,N_7227,N_6126);
and U8990 (N_8990,N_6907,N_7474);
nor U8991 (N_8991,N_6580,N_6060);
and U8992 (N_8992,N_7403,N_7168);
nor U8993 (N_8993,N_6828,N_6936);
and U8994 (N_8994,N_6866,N_6255);
xor U8995 (N_8995,N_6598,N_6113);
nor U8996 (N_8996,N_7365,N_6498);
and U8997 (N_8997,N_7279,N_6142);
or U8998 (N_8998,N_6615,N_7187);
or U8999 (N_8999,N_7003,N_7019);
xnor U9000 (N_9000,N_8619,N_8047);
nand U9001 (N_9001,N_8379,N_7559);
nand U9002 (N_9002,N_8974,N_8804);
nor U9003 (N_9003,N_8787,N_7526);
or U9004 (N_9004,N_8874,N_7724);
nand U9005 (N_9005,N_8881,N_7728);
and U9006 (N_9006,N_8142,N_8733);
nor U9007 (N_9007,N_8094,N_8178);
and U9008 (N_9008,N_8423,N_8409);
and U9009 (N_9009,N_8986,N_7732);
and U9010 (N_9010,N_8954,N_7830);
xnor U9011 (N_9011,N_7772,N_8742);
nand U9012 (N_9012,N_7590,N_8893);
nor U9013 (N_9013,N_7966,N_8554);
xnor U9014 (N_9014,N_8041,N_7869);
and U9015 (N_9015,N_8244,N_7517);
xor U9016 (N_9016,N_7843,N_7537);
and U9017 (N_9017,N_7828,N_7620);
xnor U9018 (N_9018,N_8664,N_8495);
or U9019 (N_9019,N_8991,N_8795);
xnor U9020 (N_9020,N_8958,N_7706);
or U9021 (N_9021,N_8578,N_8362);
nand U9022 (N_9022,N_7592,N_8239);
nor U9023 (N_9023,N_7886,N_8929);
xor U9024 (N_9024,N_8382,N_8318);
nand U9025 (N_9025,N_8747,N_8214);
nor U9026 (N_9026,N_7527,N_8316);
nor U9027 (N_9027,N_8345,N_7961);
nand U9028 (N_9028,N_7556,N_8801);
or U9029 (N_9029,N_8241,N_8538);
and U9030 (N_9030,N_8890,N_7532);
and U9031 (N_9031,N_7599,N_8820);
and U9032 (N_9032,N_8509,N_8055);
and U9033 (N_9033,N_7936,N_8254);
nor U9034 (N_9034,N_8541,N_8788);
and U9035 (N_9035,N_8597,N_8267);
or U9036 (N_9036,N_8397,N_7916);
nand U9037 (N_9037,N_8411,N_7500);
or U9038 (N_9038,N_7914,N_8628);
or U9039 (N_9039,N_8205,N_7817);
nor U9040 (N_9040,N_7920,N_8764);
xnor U9041 (N_9041,N_7861,N_7725);
nand U9042 (N_9042,N_8573,N_8425);
xnor U9043 (N_9043,N_7822,N_8338);
nand U9044 (N_9044,N_7638,N_8662);
nor U9045 (N_9045,N_7855,N_8852);
nor U9046 (N_9046,N_8160,N_8593);
nor U9047 (N_9047,N_8072,N_8806);
and U9048 (N_9048,N_8431,N_7867);
xnor U9049 (N_9049,N_8661,N_7697);
or U9050 (N_9050,N_8962,N_7747);
nand U9051 (N_9051,N_8175,N_7510);
nor U9052 (N_9052,N_7710,N_8729);
xnor U9053 (N_9053,N_8930,N_8885);
xnor U9054 (N_9054,N_8670,N_8896);
and U9055 (N_9055,N_7603,N_8070);
nor U9056 (N_9056,N_8627,N_8704);
xor U9057 (N_9057,N_7654,N_8319);
nor U9058 (N_9058,N_8665,N_8513);
and U9059 (N_9059,N_7671,N_8129);
xor U9060 (N_9060,N_7678,N_8759);
xnor U9061 (N_9061,N_7972,N_7960);
and U9062 (N_9062,N_8009,N_7845);
and U9063 (N_9063,N_8892,N_8689);
or U9064 (N_9064,N_8410,N_8613);
nand U9065 (N_9065,N_7655,N_8500);
or U9066 (N_9066,N_8184,N_8924);
or U9067 (N_9067,N_8297,N_7739);
or U9068 (N_9068,N_7880,N_8543);
xnor U9069 (N_9069,N_7698,N_7502);
and U9070 (N_9070,N_8906,N_8420);
nor U9071 (N_9071,N_8678,N_8865);
or U9072 (N_9072,N_7505,N_8427);
nand U9073 (N_9073,N_8153,N_7695);
and U9074 (N_9074,N_7594,N_8652);
nor U9075 (N_9075,N_8829,N_8726);
nor U9076 (N_9076,N_7777,N_8372);
and U9077 (N_9077,N_7516,N_7995);
nor U9078 (N_9078,N_7956,N_7874);
or U9079 (N_9079,N_8909,N_8468);
nand U9080 (N_9080,N_8780,N_8832);
and U9081 (N_9081,N_8931,N_8115);
or U9082 (N_9082,N_8353,N_8077);
xnor U9083 (N_9083,N_8220,N_8386);
nor U9084 (N_9084,N_8162,N_7955);
and U9085 (N_9085,N_8935,N_7998);
or U9086 (N_9086,N_8789,N_8794);
and U9087 (N_9087,N_8008,N_8060);
nand U9088 (N_9088,N_8143,N_7737);
nand U9089 (N_9089,N_8128,N_7969);
or U9090 (N_9090,N_8484,N_8154);
or U9091 (N_9091,N_8713,N_8089);
and U9092 (N_9092,N_8540,N_8566);
xor U9093 (N_9093,N_7858,N_7607);
nor U9094 (N_9094,N_8574,N_7799);
or U9095 (N_9095,N_7949,N_8163);
nor U9096 (N_9096,N_7823,N_7504);
xnor U9097 (N_9097,N_7711,N_8100);
nor U9098 (N_9098,N_8586,N_8768);
xnor U9099 (N_9099,N_8398,N_8630);
and U9100 (N_9100,N_8260,N_8440);
xor U9101 (N_9101,N_8135,N_8772);
nor U9102 (N_9102,N_7693,N_8465);
xor U9103 (N_9103,N_8549,N_8149);
or U9104 (N_9104,N_8479,N_7853);
xnor U9105 (N_9105,N_7876,N_7641);
or U9106 (N_9106,N_8104,N_8951);
nor U9107 (N_9107,N_8512,N_7703);
nor U9108 (N_9108,N_7791,N_7952);
and U9109 (N_9109,N_8918,N_8373);
and U9110 (N_9110,N_8034,N_8570);
and U9111 (N_9111,N_8348,N_8843);
nor U9112 (N_9112,N_8022,N_7596);
nor U9113 (N_9113,N_8108,N_8114);
nand U9114 (N_9114,N_7834,N_7913);
xnor U9115 (N_9115,N_8807,N_8288);
and U9116 (N_9116,N_8731,N_7629);
and U9117 (N_9117,N_8914,N_7776);
nand U9118 (N_9118,N_8050,N_8840);
nor U9119 (N_9119,N_7701,N_8413);
and U9120 (N_9120,N_8537,N_7887);
nor U9121 (N_9121,N_7912,N_7587);
and U9122 (N_9122,N_8252,N_8990);
xnor U9123 (N_9123,N_7536,N_7752);
and U9124 (N_9124,N_8478,N_7968);
nor U9125 (N_9125,N_8247,N_8854);
xnor U9126 (N_9126,N_8053,N_7902);
nor U9127 (N_9127,N_8476,N_8728);
or U9128 (N_9128,N_7657,N_8591);
nand U9129 (N_9129,N_7790,N_7636);
xor U9130 (N_9130,N_8816,N_8296);
and U9131 (N_9131,N_8092,N_8195);
and U9132 (N_9132,N_8185,N_8341);
or U9133 (N_9133,N_8922,N_8000);
nand U9134 (N_9134,N_7651,N_7846);
or U9135 (N_9135,N_8636,N_7940);
or U9136 (N_9136,N_8993,N_8227);
xnor U9137 (N_9137,N_8883,N_7922);
xor U9138 (N_9138,N_8818,N_8278);
or U9139 (N_9139,N_8091,N_7925);
nor U9140 (N_9140,N_8847,N_8947);
nand U9141 (N_9141,N_7882,N_8708);
nand U9142 (N_9142,N_8192,N_7770);
xnor U9143 (N_9143,N_8350,N_8324);
nor U9144 (N_9144,N_7754,N_8119);
xnor U9145 (N_9145,N_8793,N_8110);
nand U9146 (N_9146,N_8394,N_8033);
xnor U9147 (N_9147,N_8926,N_8606);
or U9148 (N_9148,N_8601,N_8248);
nor U9149 (N_9149,N_7679,N_8087);
nor U9150 (N_9150,N_7999,N_8402);
and U9151 (N_9151,N_7900,N_7988);
nor U9152 (N_9152,N_8404,N_8377);
xor U9153 (N_9153,N_8870,N_8891);
xnor U9154 (N_9154,N_8528,N_7917);
nor U9155 (N_9155,N_8975,N_7808);
and U9156 (N_9156,N_8849,N_8778);
nor U9157 (N_9157,N_8718,N_8766);
xnor U9158 (N_9158,N_7552,N_8539);
nor U9159 (N_9159,N_8668,N_8457);
and U9160 (N_9160,N_8805,N_8786);
and U9161 (N_9161,N_7633,N_7781);
or U9162 (N_9162,N_7722,N_8577);
nor U9163 (N_9163,N_8051,N_7555);
nand U9164 (N_9164,N_8561,N_8030);
and U9165 (N_9165,N_7899,N_8069);
nand U9166 (N_9166,N_8273,N_7692);
nand U9167 (N_9167,N_7896,N_8463);
and U9168 (N_9168,N_8756,N_7875);
and U9169 (N_9169,N_8658,N_8682);
xnor U9170 (N_9170,N_7736,N_8466);
and U9171 (N_9171,N_8871,N_8284);
or U9172 (N_9172,N_7780,N_7741);
or U9173 (N_9173,N_7616,N_7818);
nand U9174 (N_9174,N_8572,N_8948);
nor U9175 (N_9175,N_8634,N_7745);
or U9176 (N_9176,N_8085,N_7582);
or U9177 (N_9177,N_8904,N_7637);
nand U9178 (N_9178,N_8120,N_7585);
or U9179 (N_9179,N_8810,N_8779);
xor U9180 (N_9180,N_8301,N_8797);
or U9181 (N_9181,N_8639,N_7782);
nand U9182 (N_9182,N_8309,N_8333);
xnor U9183 (N_9183,N_8331,N_8304);
or U9184 (N_9184,N_8898,N_8710);
and U9185 (N_9185,N_8270,N_8356);
xnor U9186 (N_9186,N_7802,N_7801);
nand U9187 (N_9187,N_7986,N_7953);
or U9188 (N_9188,N_8439,N_8702);
nand U9189 (N_9189,N_7542,N_8231);
and U9190 (N_9190,N_8723,N_7577);
and U9191 (N_9191,N_8815,N_8167);
and U9192 (N_9192,N_8230,N_8863);
nand U9193 (N_9193,N_8103,N_8755);
nand U9194 (N_9194,N_8955,N_8113);
nand U9195 (N_9195,N_8151,N_7560);
nand U9196 (N_9196,N_8590,N_8327);
and U9197 (N_9197,N_8204,N_8878);
or U9198 (N_9198,N_8453,N_8263);
and U9199 (N_9199,N_7888,N_8999);
nor U9200 (N_9200,N_8071,N_7879);
and U9201 (N_9201,N_7826,N_8711);
or U9202 (N_9202,N_8531,N_7612);
nor U9203 (N_9203,N_7809,N_8827);
or U9204 (N_9204,N_8587,N_8169);
nand U9205 (N_9205,N_8364,N_7562);
xor U9206 (N_9206,N_8366,N_8322);
and U9207 (N_9207,N_8491,N_7709);
and U9208 (N_9208,N_8242,N_8623);
and U9209 (N_9209,N_8800,N_8443);
nor U9210 (N_9210,N_8503,N_8378);
xnor U9211 (N_9211,N_7981,N_7756);
nor U9212 (N_9212,N_7571,N_8717);
nor U9213 (N_9213,N_8703,N_8403);
nand U9214 (N_9214,N_7575,N_7815);
and U9215 (N_9215,N_8346,N_7719);
or U9216 (N_9216,N_8433,N_8486);
or U9217 (N_9217,N_8166,N_8106);
and U9218 (N_9218,N_7531,N_8837);
xor U9219 (N_9219,N_8551,N_8046);
nand U9220 (N_9220,N_8140,N_8620);
and U9221 (N_9221,N_8920,N_8560);
nor U9222 (N_9222,N_8208,N_8734);
or U9223 (N_9223,N_7622,N_7570);
and U9224 (N_9224,N_8611,N_8158);
nor U9225 (N_9225,N_8957,N_7519);
and U9226 (N_9226,N_7591,N_8029);
or U9227 (N_9227,N_8858,N_8588);
xor U9228 (N_9228,N_8760,N_8553);
nor U9229 (N_9229,N_8493,N_7712);
nand U9230 (N_9230,N_8112,N_7840);
nor U9231 (N_9231,N_7755,N_8349);
nor U9232 (N_9232,N_8375,N_7634);
xor U9233 (N_9233,N_8361,N_8363);
and U9234 (N_9234,N_7850,N_8889);
xor U9235 (N_9235,N_8902,N_8171);
xnor U9236 (N_9236,N_8277,N_8721);
and U9237 (N_9237,N_7690,N_8732);
xor U9238 (N_9238,N_7783,N_7950);
or U9239 (N_9239,N_8025,N_7515);
nand U9240 (N_9240,N_8438,N_8381);
or U9241 (N_9241,N_8691,N_8698);
or U9242 (N_9242,N_7849,N_8651);
or U9243 (N_9243,N_7716,N_8367);
nand U9244 (N_9244,N_8524,N_7918);
xnor U9245 (N_9245,N_7564,N_8095);
xor U9246 (N_9246,N_8763,N_8547);
xnor U9247 (N_9247,N_8196,N_8434);
xor U9248 (N_9248,N_8099,N_8474);
and U9249 (N_9249,N_8645,N_8281);
and U9250 (N_9250,N_8222,N_8170);
or U9251 (N_9251,N_7765,N_8888);
xor U9252 (N_9252,N_7676,N_7885);
or U9253 (N_9253,N_8855,N_7557);
nand U9254 (N_9254,N_8680,N_8499);
xor U9255 (N_9255,N_8532,N_8761);
nand U9256 (N_9256,N_7535,N_8328);
and U9257 (N_9257,N_7865,N_8943);
xnor U9258 (N_9258,N_8335,N_7584);
xor U9259 (N_9259,N_7685,N_8203);
xnor U9260 (N_9260,N_7806,N_8688);
xnor U9261 (N_9261,N_8285,N_7743);
and U9262 (N_9262,N_8769,N_8546);
xnor U9263 (N_9263,N_8102,N_8831);
and U9264 (N_9264,N_8641,N_7829);
or U9265 (N_9265,N_8938,N_8496);
nor U9266 (N_9266,N_8841,N_8988);
nor U9267 (N_9267,N_8121,N_8494);
nand U9268 (N_9268,N_7859,N_8743);
or U9269 (N_9269,N_8441,N_8264);
and U9270 (N_9270,N_7750,N_8207);
xor U9271 (N_9271,N_8152,N_7501);
and U9272 (N_9272,N_8576,N_8730);
xor U9273 (N_9273,N_7661,N_8482);
nor U9274 (N_9274,N_8687,N_8706);
nand U9275 (N_9275,N_8308,N_7904);
and U9276 (N_9276,N_7522,N_8908);
and U9277 (N_9277,N_7694,N_7565);
nor U9278 (N_9278,N_8498,N_8255);
nand U9279 (N_9279,N_8236,N_8635);
nor U9280 (N_9280,N_8995,N_7814);
nor U9281 (N_9281,N_7863,N_8905);
or U9282 (N_9282,N_8853,N_8953);
nor U9283 (N_9283,N_7820,N_8727);
nand U9284 (N_9284,N_8798,N_7740);
and U9285 (N_9285,N_8799,N_8844);
nor U9286 (N_9286,N_7675,N_7906);
nand U9287 (N_9287,N_8568,N_7851);
nand U9288 (N_9288,N_7568,N_8980);
xor U9289 (N_9289,N_8490,N_8666);
nand U9290 (N_9290,N_7841,N_7523);
nand U9291 (N_9291,N_8740,N_8336);
nand U9292 (N_9292,N_7757,N_7976);
nand U9293 (N_9293,N_8998,N_8867);
nand U9294 (N_9294,N_8830,N_8256);
nand U9295 (N_9295,N_8396,N_8834);
or U9296 (N_9296,N_8295,N_8021);
and U9297 (N_9297,N_8464,N_8719);
nor U9298 (N_9298,N_7589,N_8963);
nand U9299 (N_9299,N_8996,N_8006);
nand U9300 (N_9300,N_8667,N_8552);
nor U9301 (N_9301,N_8392,N_8646);
nor U9302 (N_9302,N_8505,N_7554);
xor U9303 (N_9303,N_7816,N_8451);
nor U9304 (N_9304,N_8456,N_8064);
nand U9305 (N_9305,N_8828,N_8020);
nand U9306 (N_9306,N_8605,N_7832);
xnor U9307 (N_9307,N_8294,N_7759);
or U9308 (N_9308,N_8073,N_7611);
nand U9309 (N_9309,N_7549,N_8442);
xnor U9310 (N_9310,N_8251,N_7856);
or U9311 (N_9311,N_8271,N_8229);
or U9312 (N_9312,N_7576,N_8038);
nand U9313 (N_9313,N_7923,N_8040);
and U9314 (N_9314,N_7528,N_8417);
or U9315 (N_9315,N_8298,N_8416);
and U9316 (N_9316,N_7786,N_7550);
or U9317 (N_9317,N_8812,N_8510);
or U9318 (N_9318,N_8369,N_8681);
nand U9319 (N_9319,N_8487,N_7521);
or U9320 (N_9320,N_8556,N_8014);
nand U9321 (N_9321,N_7650,N_7720);
xnor U9322 (N_9322,N_8011,N_7793);
xnor U9323 (N_9323,N_8389,N_8508);
xnor U9324 (N_9324,N_8399,N_8131);
and U9325 (N_9325,N_7928,N_8686);
or U9326 (N_9326,N_8084,N_7768);
xnor U9327 (N_9327,N_8065,N_8714);
nor U9328 (N_9328,N_7677,N_7563);
and U9329 (N_9329,N_8387,N_7803);
nand U9330 (N_9330,N_7919,N_8895);
xnor U9331 (N_9331,N_8982,N_8330);
xor U9332 (N_9332,N_8137,N_8567);
or U9333 (N_9333,N_8638,N_8992);
or U9334 (N_9334,N_7566,N_7893);
or U9335 (N_9335,N_8019,N_8059);
nor U9336 (N_9336,N_7957,N_8783);
or U9337 (N_9337,N_7561,N_8529);
or U9338 (N_9338,N_8901,N_7789);
xnor U9339 (N_9339,N_8640,N_8074);
and U9340 (N_9340,N_8984,N_8481);
nand U9341 (N_9341,N_8024,N_8985);
or U9342 (N_9342,N_8912,N_7942);
nor U9343 (N_9343,N_7715,N_8649);
nand U9344 (N_9344,N_8633,N_7993);
nor U9345 (N_9345,N_7738,N_8432);
and U9346 (N_9346,N_8283,N_8079);
or U9347 (N_9347,N_7898,N_8408);
or U9348 (N_9348,N_7586,N_8693);
nor U9349 (N_9349,N_8968,N_8961);
nor U9350 (N_9350,N_8326,N_7558);
xor U9351 (N_9351,N_8048,N_7658);
nor U9352 (N_9352,N_8249,N_7509);
or U9353 (N_9353,N_8565,N_8562);
nor U9354 (N_9354,N_7862,N_8595);
or U9355 (N_9355,N_8514,N_8967);
nor U9356 (N_9356,N_8809,N_8765);
nor U9357 (N_9357,N_7771,N_7775);
nand U9358 (N_9358,N_8965,N_7503);
and U9359 (N_9359,N_8679,N_7614);
xor U9360 (N_9360,N_8146,N_8360);
nor U9361 (N_9361,N_8545,N_8226);
xnor U9362 (N_9362,N_8879,N_7742);
xor U9363 (N_9363,N_7908,N_8604);
or U9364 (N_9364,N_7933,N_7967);
and U9365 (N_9365,N_8467,N_8268);
nor U9366 (N_9366,N_8861,N_7991);
nor U9367 (N_9367,N_8873,N_7630);
and U9368 (N_9368,N_7890,N_8511);
and U9369 (N_9369,N_8004,N_8186);
nor U9370 (N_9370,N_8157,N_8132);
nand U9371 (N_9371,N_8976,N_8240);
and U9372 (N_9372,N_8107,N_7717);
nand U9373 (N_9373,N_8803,N_7718);
nand U9374 (N_9374,N_8390,N_8564);
nor U9375 (N_9375,N_8882,N_8615);
nand U9376 (N_9376,N_8542,N_7761);
nand U9377 (N_9377,N_8603,N_8007);
or U9378 (N_9378,N_7621,N_8872);
xor U9379 (N_9379,N_7699,N_7787);
and U9380 (N_9380,N_7686,N_8981);
or U9381 (N_9381,N_8944,N_8238);
and U9382 (N_9382,N_7812,N_7663);
nor U9383 (N_9383,N_8475,N_8994);
xor U9384 (N_9384,N_8825,N_8148);
nand U9385 (N_9385,N_8215,N_7970);
and U9386 (N_9386,N_7769,N_7892);
nor U9387 (N_9387,N_8272,N_8483);
xnor U9388 (N_9388,N_8637,N_8090);
nor U9389 (N_9389,N_7926,N_8032);
or U9390 (N_9390,N_7702,N_8673);
and U9391 (N_9391,N_8875,N_7931);
or U9392 (N_9392,N_8307,N_8428);
or U9393 (N_9393,N_8470,N_7895);
xnor U9394 (N_9394,N_8598,N_8447);
nor U9395 (N_9395,N_7696,N_7682);
and U9396 (N_9396,N_8237,N_7911);
xor U9397 (N_9397,N_8013,N_8650);
nor U9398 (N_9398,N_8826,N_8842);
or U9399 (N_9399,N_7598,N_7626);
or U9400 (N_9400,N_7935,N_8973);
xor U9401 (N_9401,N_8243,N_8705);
and U9402 (N_9402,N_8492,N_8683);
nand U9403 (N_9403,N_8675,N_7929);
xor U9404 (N_9404,N_7871,N_8315);
and U9405 (N_9405,N_8534,N_8536);
or U9406 (N_9406,N_8559,N_8471);
or U9407 (N_9407,N_8219,N_8023);
and U9408 (N_9408,N_7656,N_8370);
or U9409 (N_9409,N_8753,N_8429);
xnor U9410 (N_9410,N_8989,N_7792);
and U9411 (N_9411,N_8602,N_8374);
or U9412 (N_9412,N_8934,N_8173);
and U9413 (N_9413,N_7667,N_8201);
nand U9414 (N_9414,N_7878,N_8395);
nand U9415 (N_9415,N_8045,N_7714);
xnor U9416 (N_9416,N_8446,N_7881);
nand U9417 (N_9417,N_8211,N_8579);
nand U9418 (N_9418,N_8111,N_8677);
xnor U9419 (N_9419,N_8280,N_8354);
and U9420 (N_9420,N_8520,N_8876);
xor U9421 (N_9421,N_8857,N_8067);
nand U9422 (N_9422,N_8629,N_7947);
xor U9423 (N_9423,N_8488,N_7649);
and U9424 (N_9424,N_8663,N_7784);
or U9425 (N_9425,N_7653,N_7540);
and U9426 (N_9426,N_7617,N_8838);
xor U9427 (N_9427,N_8003,N_8616);
or U9428 (N_9428,N_7860,N_8784);
xor U9429 (N_9429,N_8262,N_8738);
nand U9430 (N_9430,N_7962,N_7797);
nor U9431 (N_9431,N_8504,N_7681);
xnor U9432 (N_9432,N_8156,N_8548);
or U9433 (N_9433,N_7864,N_8480);
and U9434 (N_9434,N_7837,N_7838);
xor U9435 (N_9435,N_8206,N_8592);
nand U9436 (N_9436,N_8697,N_8235);
nand U9437 (N_9437,N_8122,N_8310);
nand U9438 (N_9438,N_8412,N_7635);
xor U9439 (N_9439,N_7602,N_8596);
or U9440 (N_9440,N_7551,N_8860);
nand U9441 (N_9441,N_8317,N_8359);
or U9442 (N_9442,N_8558,N_8458);
or U9443 (N_9443,N_8342,N_8609);
and U9444 (N_9444,N_8233,N_7762);
and U9445 (N_9445,N_7990,N_7889);
xor U9446 (N_9446,N_8773,N_8979);
xnor U9447 (N_9447,N_7723,N_8462);
and U9448 (N_9448,N_8737,N_8058);
or U9449 (N_9449,N_7733,N_7945);
nand U9450 (N_9450,N_7645,N_8671);
xor U9451 (N_9451,N_8744,N_7615);
nor U9452 (N_9452,N_8161,N_8501);
and U9453 (N_9453,N_8191,N_7613);
xor U9454 (N_9454,N_8197,N_7627);
nand U9455 (N_9455,N_8179,N_8919);
or U9456 (N_9456,N_8581,N_8213);
or U9457 (N_9457,N_8117,N_8915);
xor U9458 (N_9458,N_7533,N_8139);
xnor U9459 (N_9459,N_8771,N_7744);
xor U9460 (N_9460,N_8325,N_7642);
xnor U9461 (N_9461,N_7569,N_7848);
nand U9462 (N_9462,N_8608,N_7643);
nand U9463 (N_9463,N_8405,N_8720);
nor U9464 (N_9464,N_8424,N_8518);
nor U9465 (N_9465,N_7839,N_8282);
nand U9466 (N_9466,N_8631,N_7921);
xor U9467 (N_9467,N_7907,N_7601);
or U9468 (N_9468,N_8725,N_7567);
or U9469 (N_9469,N_8583,N_8724);
or U9470 (N_9470,N_8292,N_8750);
nor U9471 (N_9471,N_8083,N_8625);
xnor U9472 (N_9472,N_8707,N_7796);
nor U9473 (N_9473,N_8515,N_8987);
xor U9474 (N_9474,N_8956,N_8460);
or U9475 (N_9475,N_7763,N_8430);
and U9476 (N_9476,N_8884,N_8887);
nor U9477 (N_9477,N_8617,N_8676);
and U9478 (N_9478,N_7513,N_7779);
and U9479 (N_9479,N_7758,N_8684);
nand U9480 (N_9480,N_8544,N_7707);
xor U9481 (N_9481,N_8563,N_8517);
nor U9482 (N_9482,N_8406,N_8669);
and U9483 (N_9483,N_8632,N_7985);
xor U9484 (N_9484,N_7539,N_7946);
nor U9485 (N_9485,N_8624,N_7688);
xnor U9486 (N_9486,N_8180,N_8530);
xnor U9487 (N_9487,N_8685,N_7943);
and U9488 (N_9488,N_7927,N_8933);
and U9489 (N_9489,N_8368,N_8945);
or U9490 (N_9490,N_8932,N_8224);
xnor U9491 (N_9491,N_7647,N_8393);
nor U9492 (N_9492,N_8977,N_8221);
xor U9493 (N_9493,N_7891,N_7963);
and U9494 (N_9494,N_8334,N_8699);
nor U9495 (N_9495,N_8018,N_8791);
nor U9496 (N_9496,N_8081,N_8261);
nand U9497 (N_9497,N_8253,N_8814);
nor U9498 (N_9498,N_8329,N_8937);
or U9499 (N_9499,N_7821,N_8928);
nor U9500 (N_9500,N_8200,N_8802);
and U9501 (N_9501,N_8066,N_8886);
nand U9502 (N_9502,N_8621,N_8716);
and U9503 (N_9503,N_7573,N_7932);
nand U9504 (N_9504,N_7588,N_8371);
or U9505 (N_9505,N_8134,N_8782);
xor U9506 (N_9506,N_8343,N_8622);
nand U9507 (N_9507,N_7974,N_7646);
and U9508 (N_9508,N_8555,N_8182);
and U9509 (N_9509,N_8299,N_8525);
nor U9510 (N_9510,N_7930,N_8751);
and U9511 (N_9511,N_8654,N_8052);
xor U9512 (N_9512,N_8469,N_7524);
nor U9513 (N_9513,N_8903,N_8250);
or U9514 (N_9514,N_8017,N_7687);
and U9515 (N_9515,N_8913,N_7794);
or U9516 (N_9516,N_7992,N_8997);
and U9517 (N_9517,N_8194,N_8824);
xor U9518 (N_9518,N_8209,N_8557);
or U9519 (N_9519,N_8746,N_7628);
and U9520 (N_9520,N_8502,N_7909);
and U9521 (N_9521,N_7606,N_7619);
nand U9522 (N_9522,N_8489,N_8384);
nand U9523 (N_9523,N_7842,N_8234);
and U9524 (N_9524,N_8454,N_8477);
or U9525 (N_9525,N_7883,N_8694);
nor U9526 (N_9526,N_7625,N_7959);
xor U9527 (N_9527,N_8848,N_8302);
nor U9528 (N_9528,N_8808,N_8877);
or U9529 (N_9529,N_7894,N_8145);
and U9530 (N_9530,N_8712,N_7574);
or U9531 (N_9531,N_8414,N_8337);
and U9532 (N_9532,N_8096,N_8618);
and U9533 (N_9533,N_7753,N_8388);
nand U9534 (N_9534,N_8695,N_8010);
xor U9535 (N_9535,N_8168,N_8228);
and U9536 (N_9536,N_8690,N_8739);
and U9537 (N_9537,N_8426,N_7978);
xnor U9538 (N_9538,N_7954,N_8049);
nand U9539 (N_9539,N_8823,N_8080);
nand U9540 (N_9540,N_8056,N_7600);
or U9541 (N_9541,N_8293,N_8864);
and U9542 (N_9542,N_8497,N_8357);
or U9543 (N_9543,N_7520,N_8358);
nor U9544 (N_9544,N_8418,N_7996);
nand U9545 (N_9545,N_7773,N_7578);
nand U9546 (N_9546,N_8286,N_8550);
and U9547 (N_9547,N_8900,N_7727);
nand U9548 (N_9548,N_8485,N_7746);
and U9549 (N_9549,N_7937,N_8016);
nand U9550 (N_9550,N_8123,N_8391);
xor U9551 (N_9551,N_7729,N_7915);
and U9552 (N_9552,N_8063,N_8754);
or U9553 (N_9553,N_8839,N_8642);
and U9554 (N_9554,N_8340,N_7508);
xor U9555 (N_9555,N_7518,N_8925);
nand U9556 (N_9556,N_8332,N_8612);
or U9557 (N_9557,N_8833,N_8124);
or U9558 (N_9558,N_8819,N_7948);
nand U9559 (N_9559,N_7983,N_7665);
xnor U9560 (N_9560,N_7529,N_8044);
xor U9561 (N_9561,N_8449,N_7831);
or U9562 (N_9562,N_8647,N_8105);
or U9563 (N_9563,N_8057,N_7609);
xor U9564 (N_9564,N_8767,N_7897);
nand U9565 (N_9565,N_8061,N_7735);
and U9566 (N_9566,N_8741,N_8571);
and U9567 (N_9567,N_8585,N_8321);
nand U9568 (N_9568,N_8519,N_8193);
xor U9569 (N_9569,N_8969,N_8098);
nand U9570 (N_9570,N_8450,N_7810);
xor U9571 (N_9571,N_8822,N_8846);
or U9572 (N_9572,N_8949,N_7639);
and U9573 (N_9573,N_8199,N_7704);
xor U9574 (N_9574,N_7873,N_8039);
xnor U9575 (N_9575,N_8522,N_8076);
and U9576 (N_9576,N_7748,N_8126);
xnor U9577 (N_9577,N_8978,N_7721);
nand U9578 (N_9578,N_7593,N_8811);
xnor U9579 (N_9579,N_7659,N_7507);
or U9580 (N_9580,N_7545,N_8435);
nand U9581 (N_9581,N_8164,N_8339);
nand U9582 (N_9582,N_8655,N_8130);
nand U9583 (N_9583,N_7708,N_7766);
or U9584 (N_9584,N_8218,N_8941);
or U9585 (N_9585,N_7547,N_7538);
and U9586 (N_9586,N_8821,N_7610);
xnor U9587 (N_9587,N_8599,N_8835);
xor U9588 (N_9588,N_8736,N_8177);
nand U9589 (N_9589,N_7713,N_8589);
and U9590 (N_9590,N_8792,N_8813);
nor U9591 (N_9591,N_8385,N_8352);
nand U9592 (N_9592,N_8300,N_8850);
nand U9593 (N_9593,N_8289,N_8189);
and U9594 (N_9594,N_8174,N_8657);
or U9595 (N_9595,N_8722,N_8715);
nor U9596 (N_9596,N_8781,N_8674);
and U9597 (N_9597,N_7666,N_8523);
and U9598 (N_9598,N_7534,N_7977);
nand U9599 (N_9599,N_7800,N_7660);
nand U9600 (N_9600,N_8043,N_7700);
xnor U9601 (N_9601,N_8380,N_8700);
and U9602 (N_9602,N_8421,N_8245);
and U9603 (N_9603,N_8959,N_8125);
or U9604 (N_9604,N_8966,N_7785);
nor U9605 (N_9605,N_7975,N_7835);
or U9606 (N_9606,N_8851,N_8983);
or U9607 (N_9607,N_8533,N_8584);
nor U9608 (N_9608,N_8972,N_8594);
nor U9609 (N_9609,N_7512,N_8461);
nor U9610 (N_9610,N_8097,N_8862);
nor U9611 (N_9611,N_8894,N_8917);
nor U9612 (N_9612,N_7905,N_7691);
nor U9613 (N_9613,N_7994,N_8257);
xnor U9614 (N_9614,N_8422,N_7813);
nand U9615 (N_9615,N_8757,N_7795);
xnor U9616 (N_9616,N_7964,N_7984);
xor U9617 (N_9617,N_8656,N_8141);
xor U9618 (N_9618,N_8190,N_8376);
or U9619 (N_9619,N_8181,N_7788);
nor U9620 (N_9620,N_7597,N_7730);
or U9621 (N_9621,N_7673,N_8002);
or U9622 (N_9622,N_8303,N_8188);
nand U9623 (N_9623,N_8709,N_7546);
xnor U9624 (N_9624,N_8653,N_8521);
nor U9625 (N_9625,N_8776,N_8287);
nand U9626 (N_9626,N_7530,N_8775);
or U9627 (N_9627,N_8015,N_7805);
nor U9628 (N_9628,N_8225,N_8323);
and U9629 (N_9629,N_8276,N_7825);
or U9630 (N_9630,N_8068,N_8940);
nand U9631 (N_9631,N_7844,N_8210);
nor U9632 (N_9632,N_7544,N_8939);
or U9633 (N_9633,N_7543,N_8644);
or U9634 (N_9634,N_8312,N_7939);
nor U9635 (N_9635,N_7624,N_8223);
nor U9636 (N_9636,N_8936,N_8749);
nor U9637 (N_9637,N_8659,N_7726);
or U9638 (N_9638,N_8660,N_8859);
nand U9639 (N_9639,N_7847,N_8155);
nor U9640 (N_9640,N_8172,N_8054);
and U9641 (N_9641,N_8028,N_8037);
and U9642 (N_9642,N_8246,N_7605);
nor U9643 (N_9643,N_7971,N_7973);
or U9644 (N_9644,N_8445,N_7689);
xnor U9645 (N_9645,N_7632,N_8614);
nor U9646 (N_9646,N_7857,N_8758);
and U9647 (N_9647,N_8745,N_8165);
or U9648 (N_9648,N_8086,N_7506);
nand U9649 (N_9649,N_8320,N_8897);
xnor U9650 (N_9650,N_8217,N_7595);
nor U9651 (N_9651,N_8610,N_7989);
nor U9652 (N_9652,N_8355,N_8845);
and U9653 (N_9653,N_7553,N_7980);
xnor U9654 (N_9654,N_7872,N_8419);
xnor U9655 (N_9655,N_7669,N_7833);
nor U9656 (N_9656,N_8516,N_7664);
xor U9657 (N_9657,N_8144,N_8198);
nand U9658 (N_9658,N_8347,N_8950);
or U9659 (N_9659,N_8527,N_7877);
nor U9660 (N_9660,N_8866,N_8176);
nor U9661 (N_9661,N_8692,N_8643);
nor U9662 (N_9662,N_8026,N_8774);
xnor U9663 (N_9663,N_8436,N_7618);
and U9664 (N_9664,N_8868,N_7934);
or U9665 (N_9665,N_8952,N_8626);
or U9666 (N_9666,N_8762,N_8042);
and U9667 (N_9667,N_7760,N_7944);
nor U9668 (N_9668,N_8305,N_8314);
and U9669 (N_9669,N_8473,N_7982);
nor U9670 (N_9670,N_8415,N_7668);
nand U9671 (N_9671,N_8290,N_7824);
nand U9672 (N_9672,N_7778,N_8078);
nor U9673 (N_9673,N_7854,N_8005);
or U9674 (N_9674,N_8400,N_7827);
xnor U9675 (N_9675,N_8817,N_8187);
nor U9676 (N_9676,N_8960,N_7979);
or U9677 (N_9677,N_7683,N_7672);
or U9678 (N_9678,N_8101,N_8970);
and U9679 (N_9679,N_8880,N_8472);
xor U9680 (N_9680,N_8790,N_8266);
xor U9681 (N_9681,N_7987,N_8075);
nand U9682 (N_9682,N_8696,N_8964);
or U9683 (N_9683,N_8232,N_7608);
and U9684 (N_9684,N_8942,N_8344);
and U9685 (N_9685,N_8093,N_7819);
nor U9686 (N_9686,N_8946,N_8401);
and U9687 (N_9687,N_8012,N_7548);
xor U9688 (N_9688,N_8265,N_7910);
xnor U9689 (N_9689,N_8600,N_8437);
and U9690 (N_9690,N_8752,N_8748);
and U9691 (N_9691,N_8569,N_8448);
or U9692 (N_9692,N_8202,N_7631);
and U9693 (N_9693,N_8082,N_7648);
nor U9694 (N_9694,N_8001,N_8607);
nand U9695 (N_9695,N_8031,N_8306);
nor U9696 (N_9696,N_7604,N_8907);
nand U9697 (N_9697,N_7525,N_7924);
and U9698 (N_9698,N_7680,N_7811);
or U9699 (N_9699,N_7965,N_8911);
nand U9700 (N_9700,N_8027,N_8147);
and U9701 (N_9701,N_7958,N_8506);
nor U9702 (N_9702,N_8927,N_8582);
nand U9703 (N_9703,N_8183,N_8735);
nor U9704 (N_9704,N_7901,N_8150);
nand U9705 (N_9705,N_7644,N_7511);
nand U9706 (N_9706,N_8455,N_8291);
or U9707 (N_9707,N_8109,N_8036);
and U9708 (N_9708,N_7684,N_8279);
and U9709 (N_9709,N_7581,N_7868);
xor U9710 (N_9710,N_8452,N_7623);
nor U9711 (N_9711,N_8274,N_8444);
nand U9712 (N_9712,N_8770,N_7572);
and U9713 (N_9713,N_8459,N_7804);
xor U9714 (N_9714,N_7705,N_8159);
or U9715 (N_9715,N_8212,N_8580);
nand U9716 (N_9716,N_7583,N_7541);
nor U9717 (N_9717,N_7662,N_8916);
or U9718 (N_9718,N_7807,N_7941);
or U9719 (N_9719,N_8258,N_7579);
nor U9720 (N_9720,N_8796,N_8118);
or U9721 (N_9721,N_8701,N_8575);
nor U9722 (N_9722,N_7751,N_8269);
xnor U9723 (N_9723,N_8971,N_7580);
or U9724 (N_9724,N_7903,N_7731);
xnor U9725 (N_9725,N_8672,N_7674);
or U9726 (N_9726,N_8313,N_8138);
xor U9727 (N_9727,N_8526,N_8910);
or U9728 (N_9728,N_8383,N_8216);
xnor U9729 (N_9729,N_8777,N_8869);
and U9730 (N_9730,N_7938,N_7951);
and U9731 (N_9731,N_7866,N_8836);
and U9732 (N_9732,N_7870,N_8365);
nor U9733 (N_9733,N_8921,N_8856);
nand U9734 (N_9734,N_8133,N_7798);
or U9735 (N_9735,N_7640,N_7734);
or U9736 (N_9736,N_7997,N_8311);
xnor U9737 (N_9737,N_8351,N_7514);
nand U9738 (N_9738,N_8899,N_8923);
nor U9739 (N_9739,N_8275,N_7764);
nor U9740 (N_9740,N_8507,N_7852);
and U9741 (N_9741,N_7884,N_8116);
or U9742 (N_9742,N_8407,N_8035);
or U9743 (N_9743,N_7767,N_8127);
nand U9744 (N_9744,N_7749,N_7652);
xor U9745 (N_9745,N_7836,N_8062);
or U9746 (N_9746,N_8136,N_8535);
and U9747 (N_9747,N_8785,N_8648);
and U9748 (N_9748,N_7670,N_8259);
and U9749 (N_9749,N_8088,N_7774);
nand U9750 (N_9750,N_8783,N_8461);
and U9751 (N_9751,N_7635,N_8278);
or U9752 (N_9752,N_8435,N_8893);
and U9753 (N_9753,N_8022,N_7973);
xnor U9754 (N_9754,N_8749,N_8268);
nand U9755 (N_9755,N_8162,N_8250);
nor U9756 (N_9756,N_8683,N_7508);
or U9757 (N_9757,N_8206,N_7586);
xor U9758 (N_9758,N_8124,N_8646);
nand U9759 (N_9759,N_8723,N_8629);
and U9760 (N_9760,N_8908,N_8587);
and U9761 (N_9761,N_8339,N_7514);
or U9762 (N_9762,N_8476,N_8506);
nor U9763 (N_9763,N_7947,N_8541);
nor U9764 (N_9764,N_8274,N_7742);
nand U9765 (N_9765,N_8232,N_8629);
nand U9766 (N_9766,N_8614,N_8893);
nand U9767 (N_9767,N_7704,N_8513);
nand U9768 (N_9768,N_8306,N_8447);
xor U9769 (N_9769,N_8620,N_8711);
xnor U9770 (N_9770,N_8095,N_7728);
nand U9771 (N_9771,N_8372,N_7936);
nor U9772 (N_9772,N_8568,N_8478);
nand U9773 (N_9773,N_8152,N_7746);
and U9774 (N_9774,N_7994,N_8981);
xnor U9775 (N_9775,N_8589,N_8643);
xor U9776 (N_9776,N_7992,N_7781);
nor U9777 (N_9777,N_8590,N_8867);
nor U9778 (N_9778,N_7717,N_8548);
xnor U9779 (N_9779,N_8229,N_8800);
nor U9780 (N_9780,N_8609,N_8469);
xor U9781 (N_9781,N_7717,N_8397);
or U9782 (N_9782,N_8505,N_8673);
nand U9783 (N_9783,N_8147,N_7725);
xnor U9784 (N_9784,N_8046,N_8730);
nor U9785 (N_9785,N_8032,N_7703);
nor U9786 (N_9786,N_8385,N_8126);
and U9787 (N_9787,N_7630,N_8730);
or U9788 (N_9788,N_8441,N_7510);
and U9789 (N_9789,N_7951,N_8655);
and U9790 (N_9790,N_8907,N_7930);
nor U9791 (N_9791,N_8553,N_7874);
or U9792 (N_9792,N_8112,N_8437);
and U9793 (N_9793,N_8107,N_7730);
xnor U9794 (N_9794,N_8980,N_7630);
and U9795 (N_9795,N_8017,N_8862);
and U9796 (N_9796,N_8316,N_8850);
and U9797 (N_9797,N_8695,N_7696);
nand U9798 (N_9798,N_8618,N_8663);
nor U9799 (N_9799,N_8460,N_7901);
and U9800 (N_9800,N_8907,N_8272);
or U9801 (N_9801,N_7530,N_8547);
or U9802 (N_9802,N_8552,N_8123);
xnor U9803 (N_9803,N_8494,N_7782);
and U9804 (N_9804,N_8633,N_8968);
nand U9805 (N_9805,N_8782,N_7595);
xor U9806 (N_9806,N_7858,N_8656);
nand U9807 (N_9807,N_8586,N_8007);
or U9808 (N_9808,N_8897,N_7761);
and U9809 (N_9809,N_7704,N_8767);
nand U9810 (N_9810,N_8316,N_7701);
nor U9811 (N_9811,N_8098,N_7908);
and U9812 (N_9812,N_8285,N_7952);
or U9813 (N_9813,N_8034,N_8717);
nand U9814 (N_9814,N_7879,N_8575);
and U9815 (N_9815,N_8433,N_7547);
and U9816 (N_9816,N_7532,N_8075);
xnor U9817 (N_9817,N_8370,N_8407);
or U9818 (N_9818,N_8237,N_7685);
and U9819 (N_9819,N_8415,N_7743);
nand U9820 (N_9820,N_8676,N_7929);
xnor U9821 (N_9821,N_8386,N_8879);
xor U9822 (N_9822,N_7879,N_8890);
xnor U9823 (N_9823,N_8358,N_8605);
xnor U9824 (N_9824,N_7641,N_8909);
nand U9825 (N_9825,N_7678,N_8623);
nor U9826 (N_9826,N_7548,N_7822);
nor U9827 (N_9827,N_8719,N_8174);
xnor U9828 (N_9828,N_7723,N_8131);
nor U9829 (N_9829,N_8043,N_7895);
and U9830 (N_9830,N_8556,N_7802);
and U9831 (N_9831,N_8335,N_8457);
and U9832 (N_9832,N_8487,N_8462);
nand U9833 (N_9833,N_7905,N_8586);
and U9834 (N_9834,N_8956,N_8464);
or U9835 (N_9835,N_8692,N_8741);
nand U9836 (N_9836,N_8235,N_7886);
xor U9837 (N_9837,N_8831,N_8423);
and U9838 (N_9838,N_7716,N_8337);
nand U9839 (N_9839,N_7938,N_7581);
nand U9840 (N_9840,N_8153,N_7647);
nor U9841 (N_9841,N_7877,N_8968);
nand U9842 (N_9842,N_7745,N_8905);
and U9843 (N_9843,N_7517,N_8885);
and U9844 (N_9844,N_8090,N_8917);
xnor U9845 (N_9845,N_8618,N_7842);
xor U9846 (N_9846,N_8457,N_8522);
and U9847 (N_9847,N_8969,N_7976);
nand U9848 (N_9848,N_8010,N_8740);
nor U9849 (N_9849,N_8533,N_7857);
and U9850 (N_9850,N_8714,N_8868);
nand U9851 (N_9851,N_8492,N_8312);
and U9852 (N_9852,N_7938,N_8878);
xor U9853 (N_9853,N_8783,N_8445);
xor U9854 (N_9854,N_8851,N_8284);
or U9855 (N_9855,N_8647,N_8818);
nand U9856 (N_9856,N_8623,N_7548);
nand U9857 (N_9857,N_8588,N_8643);
and U9858 (N_9858,N_8334,N_8976);
nand U9859 (N_9859,N_7707,N_8039);
xor U9860 (N_9860,N_8494,N_8486);
or U9861 (N_9861,N_7981,N_7865);
xnor U9862 (N_9862,N_8496,N_8858);
nor U9863 (N_9863,N_7925,N_8385);
nor U9864 (N_9864,N_8740,N_8153);
or U9865 (N_9865,N_8954,N_8828);
and U9866 (N_9866,N_7798,N_7813);
and U9867 (N_9867,N_7820,N_7746);
nand U9868 (N_9868,N_8099,N_8129);
xnor U9869 (N_9869,N_8758,N_8295);
nand U9870 (N_9870,N_8403,N_7633);
and U9871 (N_9871,N_7962,N_7690);
nand U9872 (N_9872,N_8259,N_8486);
or U9873 (N_9873,N_8783,N_7794);
xnor U9874 (N_9874,N_8014,N_7931);
nor U9875 (N_9875,N_8802,N_8208);
and U9876 (N_9876,N_8585,N_8193);
and U9877 (N_9877,N_7717,N_7503);
xnor U9878 (N_9878,N_7711,N_7836);
xor U9879 (N_9879,N_8747,N_8542);
and U9880 (N_9880,N_8417,N_7743);
or U9881 (N_9881,N_8200,N_7978);
xnor U9882 (N_9882,N_8357,N_7714);
and U9883 (N_9883,N_7930,N_8472);
nand U9884 (N_9884,N_8344,N_8046);
nor U9885 (N_9885,N_8149,N_8185);
nor U9886 (N_9886,N_8128,N_7565);
and U9887 (N_9887,N_8802,N_8720);
nand U9888 (N_9888,N_8955,N_8862);
xor U9889 (N_9889,N_8502,N_7898);
nand U9890 (N_9890,N_8929,N_8723);
nand U9891 (N_9891,N_8130,N_8412);
or U9892 (N_9892,N_7851,N_8458);
xor U9893 (N_9893,N_8619,N_7605);
nand U9894 (N_9894,N_8110,N_7927);
nand U9895 (N_9895,N_8783,N_7887);
nor U9896 (N_9896,N_7797,N_8062);
or U9897 (N_9897,N_8745,N_8140);
nor U9898 (N_9898,N_8969,N_7580);
nor U9899 (N_9899,N_8464,N_8582);
xor U9900 (N_9900,N_8110,N_7712);
xnor U9901 (N_9901,N_7986,N_8184);
or U9902 (N_9902,N_7849,N_8483);
nor U9903 (N_9903,N_8871,N_7928);
xnor U9904 (N_9904,N_8156,N_8841);
xor U9905 (N_9905,N_8018,N_7985);
nand U9906 (N_9906,N_8557,N_8969);
or U9907 (N_9907,N_8994,N_8406);
nor U9908 (N_9908,N_8523,N_8275);
or U9909 (N_9909,N_8308,N_8007);
xnor U9910 (N_9910,N_8633,N_8096);
nand U9911 (N_9911,N_8978,N_8750);
xnor U9912 (N_9912,N_7535,N_8539);
nor U9913 (N_9913,N_8648,N_7934);
xor U9914 (N_9914,N_8309,N_8877);
nor U9915 (N_9915,N_8447,N_8008);
and U9916 (N_9916,N_8295,N_8275);
or U9917 (N_9917,N_8923,N_7599);
nand U9918 (N_9918,N_8039,N_7511);
xnor U9919 (N_9919,N_7915,N_7511);
or U9920 (N_9920,N_8683,N_8718);
and U9921 (N_9921,N_8081,N_8243);
nor U9922 (N_9922,N_8861,N_7595);
xor U9923 (N_9923,N_8399,N_8165);
xnor U9924 (N_9924,N_7891,N_8278);
or U9925 (N_9925,N_8620,N_8603);
and U9926 (N_9926,N_8207,N_8924);
xnor U9927 (N_9927,N_8515,N_7533);
or U9928 (N_9928,N_8527,N_7874);
nor U9929 (N_9929,N_8951,N_8263);
xnor U9930 (N_9930,N_8389,N_8991);
nor U9931 (N_9931,N_7907,N_8846);
nor U9932 (N_9932,N_8318,N_7709);
nand U9933 (N_9933,N_8676,N_8713);
or U9934 (N_9934,N_8745,N_7900);
nand U9935 (N_9935,N_8691,N_8797);
nor U9936 (N_9936,N_8153,N_8766);
nor U9937 (N_9937,N_7680,N_7570);
and U9938 (N_9938,N_8744,N_8738);
and U9939 (N_9939,N_7975,N_7934);
xor U9940 (N_9940,N_7936,N_8573);
and U9941 (N_9941,N_8888,N_8856);
nand U9942 (N_9942,N_8661,N_7694);
nand U9943 (N_9943,N_8930,N_7693);
and U9944 (N_9944,N_8162,N_7598);
or U9945 (N_9945,N_8821,N_7527);
and U9946 (N_9946,N_8590,N_8103);
xnor U9947 (N_9947,N_8626,N_7650);
nor U9948 (N_9948,N_8111,N_8308);
or U9949 (N_9949,N_7594,N_8916);
xnor U9950 (N_9950,N_8295,N_8671);
or U9951 (N_9951,N_8054,N_7923);
and U9952 (N_9952,N_8633,N_8811);
nand U9953 (N_9953,N_7978,N_8944);
or U9954 (N_9954,N_8751,N_8401);
nand U9955 (N_9955,N_8363,N_8016);
and U9956 (N_9956,N_8364,N_8747);
xnor U9957 (N_9957,N_8969,N_7658);
nor U9958 (N_9958,N_8531,N_8166);
nand U9959 (N_9959,N_8901,N_8719);
nor U9960 (N_9960,N_8588,N_8711);
nor U9961 (N_9961,N_8594,N_8427);
nand U9962 (N_9962,N_8976,N_8217);
xor U9963 (N_9963,N_7999,N_8865);
and U9964 (N_9964,N_8762,N_8023);
or U9965 (N_9965,N_7842,N_8123);
and U9966 (N_9966,N_8470,N_8005);
or U9967 (N_9967,N_7771,N_8674);
xnor U9968 (N_9968,N_7590,N_8790);
nor U9969 (N_9969,N_7661,N_8186);
nand U9970 (N_9970,N_7840,N_8138);
nor U9971 (N_9971,N_7542,N_8904);
nand U9972 (N_9972,N_8824,N_8718);
xor U9973 (N_9973,N_8078,N_8299);
nor U9974 (N_9974,N_8816,N_8273);
and U9975 (N_9975,N_7662,N_8255);
nor U9976 (N_9976,N_8388,N_8437);
or U9977 (N_9977,N_8009,N_8818);
nand U9978 (N_9978,N_8233,N_7717);
xnor U9979 (N_9979,N_8058,N_8313);
or U9980 (N_9980,N_7906,N_7536);
or U9981 (N_9981,N_7996,N_8925);
nand U9982 (N_9982,N_8352,N_8108);
nand U9983 (N_9983,N_8823,N_7719);
nor U9984 (N_9984,N_7836,N_8230);
nand U9985 (N_9985,N_8158,N_7766);
and U9986 (N_9986,N_7747,N_8368);
and U9987 (N_9987,N_8595,N_8451);
or U9988 (N_9988,N_8159,N_8056);
nand U9989 (N_9989,N_8181,N_8627);
and U9990 (N_9990,N_7952,N_8621);
nor U9991 (N_9991,N_7796,N_7651);
and U9992 (N_9992,N_7818,N_7811);
xnor U9993 (N_9993,N_7930,N_8599);
nand U9994 (N_9994,N_7891,N_8834);
nand U9995 (N_9995,N_7880,N_8631);
xor U9996 (N_9996,N_7754,N_8927);
xor U9997 (N_9997,N_8193,N_8714);
xor U9998 (N_9998,N_8112,N_8855);
xnor U9999 (N_9999,N_8627,N_8210);
nor U10000 (N_10000,N_7838,N_8837);
xnor U10001 (N_10001,N_7786,N_7522);
xnor U10002 (N_10002,N_7850,N_8571);
nand U10003 (N_10003,N_8748,N_8686);
and U10004 (N_10004,N_8199,N_8668);
xnor U10005 (N_10005,N_7544,N_7704);
and U10006 (N_10006,N_8596,N_8290);
nand U10007 (N_10007,N_8047,N_8374);
or U10008 (N_10008,N_7844,N_8241);
nand U10009 (N_10009,N_8657,N_8658);
or U10010 (N_10010,N_7763,N_8778);
nand U10011 (N_10011,N_8722,N_7872);
or U10012 (N_10012,N_8433,N_7997);
and U10013 (N_10013,N_7795,N_8491);
nor U10014 (N_10014,N_8416,N_7657);
nor U10015 (N_10015,N_8567,N_8519);
and U10016 (N_10016,N_7797,N_7865);
or U10017 (N_10017,N_8153,N_8026);
or U10018 (N_10018,N_8586,N_8504);
and U10019 (N_10019,N_8518,N_7963);
and U10020 (N_10020,N_8662,N_8500);
xor U10021 (N_10021,N_8782,N_8738);
or U10022 (N_10022,N_8431,N_7661);
or U10023 (N_10023,N_8401,N_7526);
nor U10024 (N_10024,N_8930,N_8351);
xor U10025 (N_10025,N_8579,N_8348);
nor U10026 (N_10026,N_8548,N_8171);
and U10027 (N_10027,N_7677,N_7892);
xnor U10028 (N_10028,N_8642,N_8556);
or U10029 (N_10029,N_8769,N_7851);
xnor U10030 (N_10030,N_8370,N_8004);
and U10031 (N_10031,N_8916,N_8380);
or U10032 (N_10032,N_7517,N_8072);
nand U10033 (N_10033,N_8228,N_8585);
nor U10034 (N_10034,N_7928,N_8961);
or U10035 (N_10035,N_8169,N_8244);
and U10036 (N_10036,N_8037,N_7698);
and U10037 (N_10037,N_8146,N_8079);
xor U10038 (N_10038,N_8310,N_8369);
nor U10039 (N_10039,N_8526,N_8218);
and U10040 (N_10040,N_8109,N_8021);
nor U10041 (N_10041,N_8817,N_8604);
nor U10042 (N_10042,N_7624,N_8134);
nor U10043 (N_10043,N_8547,N_7884);
or U10044 (N_10044,N_8232,N_8827);
nor U10045 (N_10045,N_7634,N_7595);
nor U10046 (N_10046,N_8031,N_8180);
xnor U10047 (N_10047,N_8106,N_8767);
nor U10048 (N_10048,N_8658,N_8244);
or U10049 (N_10049,N_8413,N_8162);
nor U10050 (N_10050,N_8975,N_7746);
or U10051 (N_10051,N_8734,N_7961);
nor U10052 (N_10052,N_8754,N_8610);
and U10053 (N_10053,N_8391,N_7791);
and U10054 (N_10054,N_7723,N_8015);
xor U10055 (N_10055,N_8191,N_7589);
or U10056 (N_10056,N_8101,N_8777);
or U10057 (N_10057,N_8949,N_8600);
xor U10058 (N_10058,N_8970,N_8963);
nand U10059 (N_10059,N_8390,N_8637);
nor U10060 (N_10060,N_8376,N_7947);
nor U10061 (N_10061,N_7788,N_8655);
nand U10062 (N_10062,N_8828,N_7505);
xnor U10063 (N_10063,N_8556,N_8492);
and U10064 (N_10064,N_7894,N_8081);
and U10065 (N_10065,N_8605,N_8969);
and U10066 (N_10066,N_8124,N_8033);
nand U10067 (N_10067,N_7768,N_8353);
and U10068 (N_10068,N_8787,N_8204);
and U10069 (N_10069,N_7898,N_8945);
nor U10070 (N_10070,N_8561,N_8517);
and U10071 (N_10071,N_8030,N_8992);
nand U10072 (N_10072,N_8445,N_8324);
and U10073 (N_10073,N_8722,N_7965);
and U10074 (N_10074,N_8621,N_7637);
nor U10075 (N_10075,N_8668,N_8791);
xnor U10076 (N_10076,N_8556,N_8003);
xor U10077 (N_10077,N_8625,N_8710);
and U10078 (N_10078,N_8870,N_7767);
or U10079 (N_10079,N_8792,N_7666);
or U10080 (N_10080,N_8444,N_8358);
nand U10081 (N_10081,N_8763,N_8678);
nand U10082 (N_10082,N_7887,N_7741);
nor U10083 (N_10083,N_8911,N_7750);
and U10084 (N_10084,N_7926,N_8098);
nand U10085 (N_10085,N_8791,N_7866);
nand U10086 (N_10086,N_8680,N_8990);
or U10087 (N_10087,N_8582,N_8919);
nand U10088 (N_10088,N_8506,N_8867);
nor U10089 (N_10089,N_8429,N_7969);
xor U10090 (N_10090,N_8390,N_7931);
xor U10091 (N_10091,N_7538,N_7753);
and U10092 (N_10092,N_8650,N_8613);
or U10093 (N_10093,N_7598,N_7854);
and U10094 (N_10094,N_8362,N_8333);
or U10095 (N_10095,N_7821,N_8945);
nand U10096 (N_10096,N_8509,N_8975);
nand U10097 (N_10097,N_8308,N_8181);
and U10098 (N_10098,N_7868,N_8920);
nor U10099 (N_10099,N_8694,N_8063);
xor U10100 (N_10100,N_7569,N_8635);
and U10101 (N_10101,N_8501,N_8209);
nand U10102 (N_10102,N_8385,N_8920);
or U10103 (N_10103,N_8428,N_7798);
or U10104 (N_10104,N_8333,N_8668);
or U10105 (N_10105,N_8829,N_8818);
xnor U10106 (N_10106,N_8530,N_8105);
nor U10107 (N_10107,N_8509,N_7688);
xnor U10108 (N_10108,N_7609,N_7984);
or U10109 (N_10109,N_7608,N_8934);
nand U10110 (N_10110,N_7734,N_8248);
and U10111 (N_10111,N_7779,N_8924);
and U10112 (N_10112,N_7817,N_8915);
nor U10113 (N_10113,N_8636,N_8613);
xnor U10114 (N_10114,N_7648,N_8814);
or U10115 (N_10115,N_8524,N_7784);
xor U10116 (N_10116,N_7648,N_8410);
nor U10117 (N_10117,N_8315,N_7530);
xnor U10118 (N_10118,N_8597,N_8931);
or U10119 (N_10119,N_8169,N_8771);
nor U10120 (N_10120,N_7510,N_7918);
and U10121 (N_10121,N_8287,N_8934);
and U10122 (N_10122,N_8325,N_8783);
or U10123 (N_10123,N_7987,N_8028);
and U10124 (N_10124,N_8652,N_8615);
nor U10125 (N_10125,N_7984,N_7696);
or U10126 (N_10126,N_8257,N_8416);
nand U10127 (N_10127,N_8974,N_8509);
nand U10128 (N_10128,N_8747,N_8731);
xor U10129 (N_10129,N_7517,N_8146);
nand U10130 (N_10130,N_8456,N_7945);
xor U10131 (N_10131,N_8487,N_8345);
or U10132 (N_10132,N_8997,N_8912);
nor U10133 (N_10133,N_7594,N_7855);
and U10134 (N_10134,N_8337,N_8697);
nor U10135 (N_10135,N_8862,N_8727);
xor U10136 (N_10136,N_7886,N_8992);
and U10137 (N_10137,N_8979,N_7936);
nand U10138 (N_10138,N_8005,N_8746);
nor U10139 (N_10139,N_7951,N_7627);
xnor U10140 (N_10140,N_7812,N_8379);
xnor U10141 (N_10141,N_8929,N_8488);
xor U10142 (N_10142,N_8937,N_8256);
xnor U10143 (N_10143,N_8833,N_7782);
xor U10144 (N_10144,N_8964,N_8056);
xor U10145 (N_10145,N_8088,N_8054);
or U10146 (N_10146,N_7829,N_8228);
nor U10147 (N_10147,N_8906,N_8261);
and U10148 (N_10148,N_7829,N_8032);
and U10149 (N_10149,N_8173,N_8692);
or U10150 (N_10150,N_8296,N_7872);
xor U10151 (N_10151,N_7666,N_7788);
and U10152 (N_10152,N_8196,N_7708);
xor U10153 (N_10153,N_8734,N_7689);
nand U10154 (N_10154,N_8008,N_8963);
and U10155 (N_10155,N_7946,N_8080);
nand U10156 (N_10156,N_8082,N_8839);
or U10157 (N_10157,N_8987,N_8225);
or U10158 (N_10158,N_8650,N_8489);
nor U10159 (N_10159,N_8593,N_7664);
and U10160 (N_10160,N_8832,N_8167);
or U10161 (N_10161,N_8588,N_8450);
or U10162 (N_10162,N_8450,N_7554);
nor U10163 (N_10163,N_7675,N_8453);
nand U10164 (N_10164,N_8373,N_8866);
nor U10165 (N_10165,N_7824,N_8904);
nand U10166 (N_10166,N_8544,N_8675);
xor U10167 (N_10167,N_8321,N_7961);
nand U10168 (N_10168,N_8451,N_7875);
nor U10169 (N_10169,N_8813,N_8017);
or U10170 (N_10170,N_7540,N_8603);
xor U10171 (N_10171,N_7619,N_8964);
or U10172 (N_10172,N_8510,N_8192);
xor U10173 (N_10173,N_7828,N_7577);
nand U10174 (N_10174,N_7616,N_8102);
xnor U10175 (N_10175,N_7799,N_7569);
xnor U10176 (N_10176,N_8851,N_7731);
nand U10177 (N_10177,N_8555,N_8158);
or U10178 (N_10178,N_8000,N_8624);
nand U10179 (N_10179,N_7740,N_8309);
nor U10180 (N_10180,N_8975,N_8564);
nand U10181 (N_10181,N_8885,N_8105);
and U10182 (N_10182,N_8643,N_8055);
and U10183 (N_10183,N_8962,N_7876);
nand U10184 (N_10184,N_7863,N_8014);
nor U10185 (N_10185,N_8205,N_7679);
and U10186 (N_10186,N_8940,N_8559);
and U10187 (N_10187,N_7646,N_7825);
xor U10188 (N_10188,N_8347,N_8524);
nor U10189 (N_10189,N_8158,N_8315);
nand U10190 (N_10190,N_7564,N_8517);
nand U10191 (N_10191,N_8394,N_8190);
or U10192 (N_10192,N_8749,N_7528);
xnor U10193 (N_10193,N_8999,N_8143);
nand U10194 (N_10194,N_7580,N_8314);
or U10195 (N_10195,N_8440,N_8003);
nor U10196 (N_10196,N_8085,N_8016);
nand U10197 (N_10197,N_8338,N_8723);
nand U10198 (N_10198,N_8047,N_7639);
nor U10199 (N_10199,N_7525,N_8861);
or U10200 (N_10200,N_8510,N_7926);
and U10201 (N_10201,N_7965,N_8101);
and U10202 (N_10202,N_7998,N_7684);
and U10203 (N_10203,N_8387,N_8877);
and U10204 (N_10204,N_7691,N_8928);
or U10205 (N_10205,N_7657,N_7648);
or U10206 (N_10206,N_7835,N_7607);
xnor U10207 (N_10207,N_8549,N_7945);
xnor U10208 (N_10208,N_8050,N_8004);
or U10209 (N_10209,N_8451,N_8250);
nand U10210 (N_10210,N_8308,N_8971);
xor U10211 (N_10211,N_8881,N_8523);
and U10212 (N_10212,N_8506,N_7928);
and U10213 (N_10213,N_8918,N_8277);
nor U10214 (N_10214,N_8670,N_8513);
nand U10215 (N_10215,N_7618,N_7772);
or U10216 (N_10216,N_8474,N_8279);
xor U10217 (N_10217,N_7537,N_8775);
or U10218 (N_10218,N_8008,N_7789);
nor U10219 (N_10219,N_8029,N_7906);
and U10220 (N_10220,N_8255,N_8213);
nand U10221 (N_10221,N_7888,N_8153);
or U10222 (N_10222,N_8876,N_8741);
and U10223 (N_10223,N_8082,N_7602);
or U10224 (N_10224,N_7745,N_8324);
xor U10225 (N_10225,N_7902,N_8074);
and U10226 (N_10226,N_7820,N_8137);
nor U10227 (N_10227,N_8201,N_8588);
or U10228 (N_10228,N_7547,N_7614);
or U10229 (N_10229,N_7921,N_8739);
and U10230 (N_10230,N_7557,N_7889);
or U10231 (N_10231,N_8473,N_8982);
nor U10232 (N_10232,N_7988,N_8892);
nor U10233 (N_10233,N_8434,N_7893);
xnor U10234 (N_10234,N_7628,N_8305);
and U10235 (N_10235,N_8191,N_8307);
or U10236 (N_10236,N_8484,N_7763);
or U10237 (N_10237,N_8456,N_7726);
xnor U10238 (N_10238,N_8390,N_8698);
nand U10239 (N_10239,N_8040,N_8706);
and U10240 (N_10240,N_8831,N_8351);
nand U10241 (N_10241,N_7547,N_8052);
xnor U10242 (N_10242,N_8198,N_8227);
nand U10243 (N_10243,N_7815,N_8078);
nand U10244 (N_10244,N_8503,N_8430);
nand U10245 (N_10245,N_8441,N_8013);
nand U10246 (N_10246,N_8786,N_8002);
or U10247 (N_10247,N_8838,N_7815);
xor U10248 (N_10248,N_8386,N_8979);
or U10249 (N_10249,N_8624,N_7798);
xor U10250 (N_10250,N_8138,N_8917);
or U10251 (N_10251,N_8876,N_7983);
or U10252 (N_10252,N_7777,N_7798);
nand U10253 (N_10253,N_7525,N_7896);
nand U10254 (N_10254,N_8669,N_7944);
nand U10255 (N_10255,N_8757,N_7842);
and U10256 (N_10256,N_8260,N_7848);
xor U10257 (N_10257,N_8900,N_8702);
nor U10258 (N_10258,N_8495,N_8093);
nor U10259 (N_10259,N_7582,N_8003);
nand U10260 (N_10260,N_8752,N_8819);
or U10261 (N_10261,N_8491,N_8179);
nor U10262 (N_10262,N_7641,N_8605);
nor U10263 (N_10263,N_8871,N_7759);
xnor U10264 (N_10264,N_8853,N_8329);
nand U10265 (N_10265,N_7519,N_7581);
and U10266 (N_10266,N_8258,N_7903);
and U10267 (N_10267,N_7990,N_8787);
or U10268 (N_10268,N_8396,N_7526);
and U10269 (N_10269,N_8041,N_8709);
or U10270 (N_10270,N_8127,N_8565);
xor U10271 (N_10271,N_8798,N_7820);
nor U10272 (N_10272,N_8052,N_8010);
and U10273 (N_10273,N_7616,N_8897);
nand U10274 (N_10274,N_8849,N_8915);
xor U10275 (N_10275,N_8110,N_8078);
or U10276 (N_10276,N_8519,N_8314);
xnor U10277 (N_10277,N_8310,N_7761);
and U10278 (N_10278,N_7670,N_8912);
and U10279 (N_10279,N_7833,N_7630);
and U10280 (N_10280,N_8624,N_7870);
xnor U10281 (N_10281,N_8565,N_8658);
xor U10282 (N_10282,N_7743,N_7576);
and U10283 (N_10283,N_7869,N_8888);
xor U10284 (N_10284,N_7744,N_8323);
xor U10285 (N_10285,N_7939,N_8701);
nand U10286 (N_10286,N_7536,N_7878);
nor U10287 (N_10287,N_7925,N_7740);
xnor U10288 (N_10288,N_8019,N_8560);
or U10289 (N_10289,N_7617,N_8755);
xnor U10290 (N_10290,N_7500,N_7962);
and U10291 (N_10291,N_8120,N_8278);
nand U10292 (N_10292,N_7717,N_8542);
or U10293 (N_10293,N_8909,N_8287);
xor U10294 (N_10294,N_7678,N_7629);
nand U10295 (N_10295,N_7743,N_8346);
nand U10296 (N_10296,N_8578,N_7784);
and U10297 (N_10297,N_8143,N_8509);
nand U10298 (N_10298,N_7790,N_8331);
nor U10299 (N_10299,N_8687,N_7792);
nand U10300 (N_10300,N_7805,N_8194);
and U10301 (N_10301,N_7738,N_8012);
or U10302 (N_10302,N_8632,N_8873);
or U10303 (N_10303,N_8124,N_8353);
nor U10304 (N_10304,N_7767,N_8254);
nand U10305 (N_10305,N_7712,N_7803);
nand U10306 (N_10306,N_8625,N_7606);
or U10307 (N_10307,N_8798,N_8710);
nor U10308 (N_10308,N_8150,N_8272);
and U10309 (N_10309,N_8854,N_8837);
and U10310 (N_10310,N_7759,N_8367);
nor U10311 (N_10311,N_8573,N_8533);
and U10312 (N_10312,N_8997,N_8824);
xor U10313 (N_10313,N_8423,N_8811);
nor U10314 (N_10314,N_8250,N_8198);
xnor U10315 (N_10315,N_8434,N_8418);
or U10316 (N_10316,N_8318,N_8241);
xor U10317 (N_10317,N_8764,N_8847);
nor U10318 (N_10318,N_8322,N_8119);
and U10319 (N_10319,N_8434,N_8445);
xnor U10320 (N_10320,N_8135,N_7906);
or U10321 (N_10321,N_8547,N_8357);
nand U10322 (N_10322,N_8472,N_8943);
nor U10323 (N_10323,N_7593,N_8448);
and U10324 (N_10324,N_7742,N_8668);
or U10325 (N_10325,N_8072,N_7506);
xor U10326 (N_10326,N_8424,N_7522);
nor U10327 (N_10327,N_8376,N_8920);
and U10328 (N_10328,N_8336,N_8816);
xnor U10329 (N_10329,N_8769,N_7882);
nand U10330 (N_10330,N_7612,N_8784);
nand U10331 (N_10331,N_7503,N_8112);
nand U10332 (N_10332,N_8352,N_7822);
xor U10333 (N_10333,N_7548,N_8599);
nand U10334 (N_10334,N_8202,N_8549);
nand U10335 (N_10335,N_7585,N_8374);
nand U10336 (N_10336,N_8574,N_8114);
xnor U10337 (N_10337,N_7665,N_7966);
nand U10338 (N_10338,N_8263,N_8075);
xnor U10339 (N_10339,N_8909,N_7559);
xnor U10340 (N_10340,N_8706,N_8733);
and U10341 (N_10341,N_7600,N_8503);
nand U10342 (N_10342,N_8337,N_7967);
nor U10343 (N_10343,N_8634,N_8701);
xor U10344 (N_10344,N_7786,N_8336);
and U10345 (N_10345,N_7831,N_8985);
nor U10346 (N_10346,N_8859,N_7894);
nor U10347 (N_10347,N_8696,N_8187);
xor U10348 (N_10348,N_8083,N_8399);
or U10349 (N_10349,N_7926,N_8544);
nand U10350 (N_10350,N_8932,N_7955);
nand U10351 (N_10351,N_7994,N_8483);
nor U10352 (N_10352,N_7645,N_7879);
and U10353 (N_10353,N_8067,N_8083);
nand U10354 (N_10354,N_8925,N_7924);
xor U10355 (N_10355,N_8220,N_8955);
or U10356 (N_10356,N_7577,N_8853);
xnor U10357 (N_10357,N_7540,N_8709);
or U10358 (N_10358,N_8492,N_8463);
nor U10359 (N_10359,N_8463,N_7608);
nand U10360 (N_10360,N_8124,N_8160);
and U10361 (N_10361,N_8694,N_7723);
and U10362 (N_10362,N_8961,N_8327);
or U10363 (N_10363,N_7514,N_8273);
or U10364 (N_10364,N_8482,N_8873);
nand U10365 (N_10365,N_7589,N_8237);
and U10366 (N_10366,N_7797,N_8331);
nand U10367 (N_10367,N_8556,N_8929);
or U10368 (N_10368,N_8729,N_7902);
and U10369 (N_10369,N_8076,N_8534);
and U10370 (N_10370,N_8414,N_7500);
xnor U10371 (N_10371,N_8573,N_8681);
nand U10372 (N_10372,N_8821,N_8047);
and U10373 (N_10373,N_8244,N_8905);
and U10374 (N_10374,N_8123,N_7657);
xnor U10375 (N_10375,N_8605,N_8222);
xnor U10376 (N_10376,N_8519,N_7556);
nor U10377 (N_10377,N_7695,N_7787);
or U10378 (N_10378,N_8288,N_7963);
xor U10379 (N_10379,N_8331,N_8389);
xnor U10380 (N_10380,N_8118,N_7804);
nand U10381 (N_10381,N_7845,N_7544);
or U10382 (N_10382,N_8357,N_7535);
and U10383 (N_10383,N_8431,N_8761);
nand U10384 (N_10384,N_7668,N_8367);
nor U10385 (N_10385,N_8970,N_8147);
nand U10386 (N_10386,N_8127,N_7844);
nand U10387 (N_10387,N_8833,N_7552);
or U10388 (N_10388,N_8606,N_8521);
or U10389 (N_10389,N_7889,N_8142);
xor U10390 (N_10390,N_8442,N_8350);
nand U10391 (N_10391,N_8451,N_8740);
xnor U10392 (N_10392,N_8419,N_8973);
nand U10393 (N_10393,N_8995,N_8900);
and U10394 (N_10394,N_8190,N_8721);
nor U10395 (N_10395,N_8832,N_8105);
nor U10396 (N_10396,N_8243,N_8072);
and U10397 (N_10397,N_7606,N_7612);
nand U10398 (N_10398,N_7801,N_7933);
or U10399 (N_10399,N_8518,N_7516);
or U10400 (N_10400,N_8167,N_7707);
nand U10401 (N_10401,N_8706,N_7761);
or U10402 (N_10402,N_7596,N_7746);
and U10403 (N_10403,N_7664,N_8776);
and U10404 (N_10404,N_8811,N_8048);
and U10405 (N_10405,N_7624,N_7788);
or U10406 (N_10406,N_8127,N_7876);
or U10407 (N_10407,N_8052,N_7733);
xnor U10408 (N_10408,N_8765,N_8906);
nor U10409 (N_10409,N_8871,N_8452);
xor U10410 (N_10410,N_7708,N_8849);
and U10411 (N_10411,N_7552,N_8002);
and U10412 (N_10412,N_8215,N_8391);
nor U10413 (N_10413,N_7841,N_8046);
and U10414 (N_10414,N_8735,N_8712);
nand U10415 (N_10415,N_8065,N_8906);
nor U10416 (N_10416,N_7605,N_7609);
nand U10417 (N_10417,N_7782,N_8384);
nor U10418 (N_10418,N_8381,N_8396);
xor U10419 (N_10419,N_8680,N_8512);
nand U10420 (N_10420,N_7962,N_8419);
nor U10421 (N_10421,N_7977,N_8201);
and U10422 (N_10422,N_8656,N_8666);
nor U10423 (N_10423,N_8362,N_8135);
and U10424 (N_10424,N_8916,N_8997);
or U10425 (N_10425,N_8051,N_7562);
and U10426 (N_10426,N_8177,N_8290);
and U10427 (N_10427,N_7680,N_8328);
nand U10428 (N_10428,N_8670,N_7508);
xnor U10429 (N_10429,N_8974,N_8259);
and U10430 (N_10430,N_7556,N_8184);
xor U10431 (N_10431,N_8934,N_7745);
or U10432 (N_10432,N_8913,N_7512);
xor U10433 (N_10433,N_8896,N_8228);
and U10434 (N_10434,N_8480,N_8847);
xnor U10435 (N_10435,N_8608,N_8127);
or U10436 (N_10436,N_7909,N_8788);
nor U10437 (N_10437,N_8478,N_8567);
or U10438 (N_10438,N_8240,N_8102);
xnor U10439 (N_10439,N_8329,N_8379);
nand U10440 (N_10440,N_8838,N_8005);
and U10441 (N_10441,N_7572,N_8350);
and U10442 (N_10442,N_8830,N_8194);
xnor U10443 (N_10443,N_8929,N_8564);
nand U10444 (N_10444,N_8024,N_7655);
or U10445 (N_10445,N_8686,N_8115);
or U10446 (N_10446,N_7697,N_7515);
or U10447 (N_10447,N_8085,N_8817);
nand U10448 (N_10448,N_8170,N_8339);
or U10449 (N_10449,N_8244,N_8678);
and U10450 (N_10450,N_7535,N_8974);
and U10451 (N_10451,N_8131,N_8412);
or U10452 (N_10452,N_7816,N_7758);
nor U10453 (N_10453,N_8963,N_7757);
nand U10454 (N_10454,N_8029,N_8712);
nand U10455 (N_10455,N_8913,N_8186);
or U10456 (N_10456,N_8658,N_8394);
and U10457 (N_10457,N_7527,N_8993);
and U10458 (N_10458,N_8469,N_7999);
and U10459 (N_10459,N_7916,N_8798);
and U10460 (N_10460,N_8985,N_7805);
xnor U10461 (N_10461,N_7718,N_8185);
nand U10462 (N_10462,N_8522,N_8341);
or U10463 (N_10463,N_8466,N_8577);
or U10464 (N_10464,N_7580,N_8484);
nand U10465 (N_10465,N_7731,N_8515);
xor U10466 (N_10466,N_7829,N_8803);
xor U10467 (N_10467,N_8481,N_7746);
xnor U10468 (N_10468,N_8562,N_8837);
xor U10469 (N_10469,N_8818,N_8175);
and U10470 (N_10470,N_8438,N_8878);
nand U10471 (N_10471,N_8470,N_8761);
nor U10472 (N_10472,N_8775,N_7971);
nor U10473 (N_10473,N_8913,N_7612);
or U10474 (N_10474,N_8273,N_8663);
or U10475 (N_10475,N_8253,N_7797);
or U10476 (N_10476,N_7943,N_8860);
nand U10477 (N_10477,N_7618,N_7646);
or U10478 (N_10478,N_7883,N_8699);
xor U10479 (N_10479,N_8133,N_8953);
or U10480 (N_10480,N_8319,N_8372);
nor U10481 (N_10481,N_8763,N_8277);
nor U10482 (N_10482,N_8250,N_8094);
and U10483 (N_10483,N_8213,N_7598);
nor U10484 (N_10484,N_8849,N_8223);
nor U10485 (N_10485,N_8026,N_7721);
nor U10486 (N_10486,N_8219,N_8099);
xor U10487 (N_10487,N_7648,N_8009);
or U10488 (N_10488,N_8232,N_7886);
xor U10489 (N_10489,N_7757,N_8442);
nor U10490 (N_10490,N_8577,N_8337);
and U10491 (N_10491,N_7600,N_7553);
and U10492 (N_10492,N_8811,N_8993);
and U10493 (N_10493,N_8639,N_8467);
xor U10494 (N_10494,N_8967,N_8004);
xor U10495 (N_10495,N_8338,N_7532);
nor U10496 (N_10496,N_7624,N_8466);
nor U10497 (N_10497,N_8100,N_8226);
nor U10498 (N_10498,N_8730,N_8204);
nor U10499 (N_10499,N_8300,N_8921);
or U10500 (N_10500,N_10254,N_9556);
and U10501 (N_10501,N_9107,N_9430);
nand U10502 (N_10502,N_10037,N_9787);
and U10503 (N_10503,N_10096,N_10235);
or U10504 (N_10504,N_10329,N_10109);
and U10505 (N_10505,N_9499,N_9889);
and U10506 (N_10506,N_9192,N_9117);
and U10507 (N_10507,N_9252,N_9687);
nor U10508 (N_10508,N_9401,N_9280);
xor U10509 (N_10509,N_9615,N_9756);
xor U10510 (N_10510,N_10131,N_9495);
xnor U10511 (N_10511,N_10028,N_10186);
or U10512 (N_10512,N_9002,N_9007);
nor U10513 (N_10513,N_10206,N_9932);
nand U10514 (N_10514,N_10091,N_9619);
nor U10515 (N_10515,N_9010,N_10279);
or U10516 (N_10516,N_9504,N_10266);
or U10517 (N_10517,N_10040,N_10288);
nor U10518 (N_10518,N_9954,N_10454);
nand U10519 (N_10519,N_9643,N_9649);
and U10520 (N_10520,N_9744,N_10209);
and U10521 (N_10521,N_9303,N_10274);
nand U10522 (N_10522,N_10436,N_10259);
xnor U10523 (N_10523,N_9282,N_9272);
and U10524 (N_10524,N_10108,N_9371);
xor U10525 (N_10525,N_9682,N_9948);
or U10526 (N_10526,N_9470,N_10126);
nor U10527 (N_10527,N_9033,N_10469);
nor U10528 (N_10528,N_9632,N_9028);
or U10529 (N_10529,N_10075,N_9096);
nor U10530 (N_10530,N_9307,N_9109);
and U10531 (N_10531,N_10322,N_10422);
nand U10532 (N_10532,N_9925,N_9129);
nand U10533 (N_10533,N_9251,N_9613);
nor U10534 (N_10534,N_9661,N_9073);
nand U10535 (N_10535,N_9937,N_9668);
and U10536 (N_10536,N_10294,N_10253);
xnor U10537 (N_10537,N_9999,N_9929);
or U10538 (N_10538,N_9903,N_9350);
xnor U10539 (N_10539,N_9158,N_9098);
xor U10540 (N_10540,N_9531,N_9311);
xor U10541 (N_10541,N_9232,N_9335);
or U10542 (N_10542,N_10029,N_10448);
nor U10543 (N_10543,N_10204,N_9960);
or U10544 (N_10544,N_9398,N_9574);
nor U10545 (N_10545,N_9612,N_9178);
xnor U10546 (N_10546,N_10391,N_10413);
xor U10547 (N_10547,N_10173,N_9936);
nor U10548 (N_10548,N_9213,N_9508);
nand U10549 (N_10549,N_9955,N_9195);
nand U10550 (N_10550,N_9344,N_10210);
nor U10551 (N_10551,N_9587,N_9841);
nand U10552 (N_10552,N_9440,N_10490);
nand U10553 (N_10553,N_10216,N_9655);
nor U10554 (N_10554,N_10095,N_9116);
and U10555 (N_10555,N_9677,N_10372);
or U10556 (N_10556,N_9286,N_10181);
and U10557 (N_10557,N_10359,N_10382);
xnor U10558 (N_10558,N_9309,N_10007);
nand U10559 (N_10559,N_9358,N_9415);
or U10560 (N_10560,N_9281,N_9701);
or U10561 (N_10561,N_9152,N_9961);
or U10562 (N_10562,N_9076,N_9603);
xor U10563 (N_10563,N_9911,N_10057);
and U10564 (N_10564,N_10114,N_10127);
xor U10565 (N_10565,N_9595,N_9862);
and U10566 (N_10566,N_9478,N_9345);
and U10567 (N_10567,N_9568,N_9635);
nand U10568 (N_10568,N_9435,N_10321);
nand U10569 (N_10569,N_9732,N_9299);
nand U10570 (N_10570,N_10384,N_9644);
and U10571 (N_10571,N_9141,N_9446);
xnor U10572 (N_10572,N_10447,N_9260);
xor U10573 (N_10573,N_9815,N_9728);
or U10574 (N_10574,N_9327,N_10174);
or U10575 (N_10575,N_9283,N_9532);
xor U10576 (N_10576,N_9498,N_9293);
xor U10577 (N_10577,N_10213,N_9512);
nand U10578 (N_10578,N_9044,N_9305);
or U10579 (N_10579,N_9792,N_9892);
nand U10580 (N_10580,N_9878,N_10123);
nor U10581 (N_10581,N_9865,N_9411);
xnor U10582 (N_10582,N_9678,N_10357);
and U10583 (N_10583,N_10129,N_9988);
or U10584 (N_10584,N_10412,N_9322);
xnor U10585 (N_10585,N_9434,N_10307);
nor U10586 (N_10586,N_9212,N_9342);
nand U10587 (N_10587,N_9514,N_9108);
and U10588 (N_10588,N_9449,N_9933);
nand U10589 (N_10589,N_10050,N_9118);
nor U10590 (N_10590,N_9242,N_9828);
or U10591 (N_10591,N_10005,N_9263);
nand U10592 (N_10592,N_10199,N_9683);
nand U10593 (N_10593,N_9692,N_9482);
and U10594 (N_10594,N_10032,N_10272);
nor U10595 (N_10595,N_10052,N_9274);
and U10596 (N_10596,N_9253,N_9579);
and U10597 (N_10597,N_9167,N_10257);
or U10598 (N_10598,N_9639,N_10161);
nand U10599 (N_10599,N_9340,N_9196);
and U10600 (N_10600,N_9941,N_9811);
and U10601 (N_10601,N_10136,N_9533);
or U10602 (N_10602,N_10484,N_9699);
or U10603 (N_10603,N_10079,N_10041);
xnor U10604 (N_10604,N_9729,N_9694);
nor U10605 (N_10605,N_9864,N_9777);
nand U10606 (N_10606,N_10227,N_9456);
or U10607 (N_10607,N_9273,N_10067);
and U10608 (N_10608,N_10232,N_9006);
nand U10609 (N_10609,N_9594,N_9951);
or U10610 (N_10610,N_9942,N_9825);
or U10611 (N_10611,N_9588,N_9234);
nand U10612 (N_10612,N_9204,N_10159);
and U10613 (N_10613,N_10142,N_9927);
and U10614 (N_10614,N_9994,N_10330);
and U10615 (N_10615,N_10332,N_9189);
xor U10616 (N_10616,N_10225,N_9236);
nand U10617 (N_10617,N_9604,N_10423);
or U10618 (N_10618,N_9645,N_10107);
xor U10619 (N_10619,N_9857,N_10256);
or U10620 (N_10620,N_10141,N_9974);
nand U10621 (N_10621,N_9560,N_9300);
or U10622 (N_10622,N_9355,N_9339);
nor U10623 (N_10623,N_9187,N_9564);
xor U10624 (N_10624,N_9170,N_9922);
nor U10625 (N_10625,N_9555,N_10416);
and U10626 (N_10626,N_10002,N_9266);
and U10627 (N_10627,N_9490,N_9057);
xor U10628 (N_10628,N_10218,N_9826);
nand U10629 (N_10629,N_9965,N_9205);
nor U10630 (N_10630,N_9709,N_9295);
nand U10631 (N_10631,N_9347,N_9392);
and U10632 (N_10632,N_10405,N_9061);
nor U10633 (N_10633,N_9944,N_9150);
or U10634 (N_10634,N_9558,N_9695);
xor U10635 (N_10635,N_9571,N_9245);
or U10636 (N_10636,N_9886,N_10264);
nand U10637 (N_10637,N_10465,N_9843);
nor U10638 (N_10638,N_9991,N_10287);
and U10639 (N_10639,N_9583,N_9627);
nor U10640 (N_10640,N_9675,N_10429);
nor U10641 (N_10641,N_9853,N_9020);
and U10642 (N_10642,N_9977,N_10080);
xnor U10643 (N_10643,N_10231,N_9525);
nand U10644 (N_10644,N_9641,N_9975);
nand U10645 (N_10645,N_9132,N_10039);
nor U10646 (N_10646,N_10027,N_9492);
or U10647 (N_10647,N_9704,N_9813);
and U10648 (N_10648,N_9503,N_10234);
or U10649 (N_10649,N_9844,N_10115);
nor U10650 (N_10650,N_10143,N_9063);
or U10651 (N_10651,N_9271,N_9467);
and U10652 (N_10652,N_9037,N_9803);
and U10653 (N_10653,N_10166,N_10017);
xor U10654 (N_10654,N_10378,N_9998);
nor U10655 (N_10655,N_10308,N_9084);
or U10656 (N_10656,N_9783,N_10432);
nand U10657 (N_10657,N_10183,N_10111);
and U10658 (N_10658,N_10138,N_9292);
and U10659 (N_10659,N_10201,N_9362);
nor U10660 (N_10660,N_9479,N_9584);
nor U10661 (N_10661,N_10192,N_9773);
and U10662 (N_10662,N_9368,N_10128);
xnor U10663 (N_10663,N_10373,N_9887);
and U10664 (N_10664,N_9209,N_10102);
xnor U10665 (N_10665,N_9698,N_9460);
and U10666 (N_10666,N_10147,N_10315);
xnor U10667 (N_10667,N_9013,N_10393);
xnor U10668 (N_10668,N_9265,N_10046);
nor U10669 (N_10669,N_9461,N_9191);
xor U10670 (N_10670,N_10311,N_9669);
or U10671 (N_10671,N_9774,N_9924);
or U10672 (N_10672,N_10471,N_10386);
nand U10673 (N_10673,N_10325,N_9876);
nor U10674 (N_10674,N_9367,N_10203);
nor U10675 (N_10675,N_10258,N_10358);
nor U10676 (N_10676,N_9953,N_10353);
xnor U10677 (N_10677,N_10292,N_9038);
nand U10678 (N_10678,N_9816,N_10160);
and U10679 (N_10679,N_10006,N_9945);
nor U10680 (N_10680,N_9314,N_9177);
xnor U10681 (N_10681,N_9992,N_9180);
xor U10682 (N_10682,N_10101,N_10026);
xor U10683 (N_10683,N_9854,N_10082);
and U10684 (N_10684,N_10056,N_9294);
and U10685 (N_10685,N_9124,N_10093);
nor U10686 (N_10686,N_9226,N_9278);
nand U10687 (N_10687,N_9050,N_10483);
nand U10688 (N_10688,N_9389,N_9384);
and U10689 (N_10689,N_9329,N_9053);
xor U10690 (N_10690,N_10389,N_9165);
and U10691 (N_10691,N_9671,N_10421);
nor U10692 (N_10692,N_10493,N_10284);
and U10693 (N_10693,N_9468,N_10276);
or U10694 (N_10694,N_9199,N_9420);
xnor U10695 (N_10695,N_9849,N_9730);
or U10696 (N_10696,N_9524,N_9220);
or U10697 (N_10697,N_10494,N_9904);
or U10698 (N_10698,N_10135,N_9636);
xnor U10699 (N_10699,N_9106,N_9254);
or U10700 (N_10700,N_9963,N_10424);
nor U10701 (N_10701,N_10461,N_9772);
xor U10702 (N_10702,N_9239,N_10238);
nor U10703 (N_10703,N_9928,N_9184);
or U10704 (N_10704,N_9032,N_9088);
and U10705 (N_10705,N_9331,N_9312);
xnor U10706 (N_10706,N_9858,N_9664);
and U10707 (N_10707,N_9802,N_10406);
xor U10708 (N_10708,N_9761,N_9867);
and U10709 (N_10709,N_9462,N_9011);
nor U10710 (N_10710,N_10489,N_9978);
xor U10711 (N_10711,N_10347,N_9735);
nor U10712 (N_10712,N_9648,N_10051);
nor U10713 (N_10713,N_9182,N_10148);
xnor U10714 (N_10714,N_10176,N_9838);
nand U10715 (N_10715,N_10185,N_10110);
and U10716 (N_10716,N_9946,N_10223);
or U10717 (N_10717,N_10118,N_9267);
or U10718 (N_10718,N_9754,N_10306);
or U10719 (N_10719,N_9001,N_10468);
xnor U10720 (N_10720,N_9959,N_10170);
nor U10721 (N_10721,N_9289,N_9334);
or U10722 (N_10722,N_9034,N_10088);
and U10723 (N_10723,N_9737,N_9706);
nand U10724 (N_10724,N_9804,N_9256);
nand U10725 (N_10725,N_9386,N_9285);
nor U10726 (N_10726,N_10177,N_9750);
nor U10727 (N_10727,N_9338,N_9169);
and U10728 (N_10728,N_10220,N_10427);
xor U10729 (N_10729,N_9776,N_10298);
nor U10730 (N_10730,N_9755,N_9638);
nand U10731 (N_10731,N_10331,N_9616);
nor U10732 (N_10732,N_9364,N_10450);
and U10733 (N_10733,N_9080,N_9696);
and U10734 (N_10734,N_9353,N_10200);
nand U10735 (N_10735,N_10197,N_9593);
nand U10736 (N_10736,N_9996,N_10409);
nand U10737 (N_10737,N_10379,N_9634);
nand U10738 (N_10738,N_9130,N_9070);
nand U10739 (N_10739,N_9238,N_10191);
and U10740 (N_10740,N_9316,N_10342);
nand U10741 (N_10741,N_9065,N_10163);
xor U10742 (N_10742,N_9374,N_9105);
or U10743 (N_10743,N_9370,N_9484);
nor U10744 (N_10744,N_9214,N_9365);
or U10745 (N_10745,N_10164,N_10252);
nor U10746 (N_10746,N_9341,N_9164);
xnor U10747 (N_10747,N_9569,N_9554);
and U10748 (N_10748,N_10215,N_9599);
nor U10749 (N_10749,N_9685,N_9247);
or U10750 (N_10750,N_9657,N_10383);
nand U10751 (N_10751,N_9742,N_10134);
or U10752 (N_10752,N_9676,N_9015);
nand U10753 (N_10753,N_9526,N_9480);
xor U10754 (N_10754,N_10282,N_9122);
nor U10755 (N_10755,N_9947,N_9137);
nand U10756 (N_10756,N_9651,N_9336);
nor U10757 (N_10757,N_10354,N_10025);
nand U10758 (N_10758,N_9969,N_9784);
or U10759 (N_10759,N_9077,N_9827);
xnor U10760 (N_10760,N_10116,N_10335);
xnor U10761 (N_10761,N_10456,N_9563);
and U10762 (N_10762,N_9097,N_10369);
xnor U10763 (N_10763,N_10497,N_9354);
and U10764 (N_10764,N_9040,N_10376);
and U10765 (N_10765,N_9127,N_9901);
or U10766 (N_10766,N_9487,N_10402);
nand U10767 (N_10767,N_9021,N_10070);
and U10768 (N_10768,N_9663,N_9085);
and U10769 (N_10769,N_9855,N_9059);
and U10770 (N_10770,N_10068,N_10410);
nor U10771 (N_10771,N_10099,N_10281);
nand U10772 (N_10772,N_10303,N_9469);
xnor U10773 (N_10773,N_10009,N_10350);
nand U10774 (N_10774,N_10226,N_9997);
or U10775 (N_10775,N_9869,N_9410);
and U10776 (N_10776,N_9348,N_9790);
nor U10777 (N_10777,N_10351,N_10316);
nand U10778 (N_10778,N_9597,N_9702);
xor U10779 (N_10779,N_9852,N_10364);
xor U10780 (N_10780,N_9891,N_9318);
xor U10781 (N_10781,N_10105,N_9351);
and U10782 (N_10782,N_10289,N_10243);
and U10783 (N_10783,N_9243,N_9095);
and U10784 (N_10784,N_9861,N_10314);
nor U10785 (N_10785,N_9403,N_9993);
xnor U10786 (N_10786,N_9731,N_9986);
or U10787 (N_10787,N_10144,N_9715);
xnor U10788 (N_10788,N_9585,N_10457);
and U10789 (N_10789,N_10362,N_9794);
or U10790 (N_10790,N_10355,N_10090);
xor U10791 (N_10791,N_10229,N_9598);
nor U10792 (N_10792,N_9596,N_9605);
xnor U10793 (N_10793,N_10348,N_9883);
or U10794 (N_10794,N_10149,N_9713);
nor U10795 (N_10795,N_10195,N_9793);
and U10796 (N_10796,N_9897,N_9019);
xnor U10797 (N_10797,N_10334,N_10375);
or U10798 (N_10798,N_9425,N_10444);
xnor U10799 (N_10799,N_9048,N_10319);
nand U10800 (N_10800,N_10438,N_9768);
nand U10801 (N_10801,N_9049,N_9407);
xnor U10802 (N_10802,N_10182,N_9464);
and U10803 (N_10803,N_9818,N_9241);
nand U10804 (N_10804,N_10363,N_9458);
or U10805 (N_10805,N_9438,N_9573);
nor U10806 (N_10806,N_9745,N_9614);
nand U10807 (N_10807,N_10133,N_9580);
xnor U10808 (N_10808,N_10341,N_10491);
or U10809 (N_10809,N_10398,N_9738);
nand U10810 (N_10810,N_9624,N_10187);
or U10811 (N_10811,N_10012,N_10420);
nor U10812 (N_10812,N_9589,N_9427);
nor U10813 (N_10813,N_9653,N_10337);
nor U10814 (N_10814,N_9778,N_10302);
or U10815 (N_10815,N_10260,N_9907);
and U10816 (N_10816,N_9136,N_9016);
and U10817 (N_10817,N_9874,N_9914);
and U10818 (N_10818,N_9210,N_10394);
xor U10819 (N_10819,N_10377,N_9629);
nand U10820 (N_10820,N_9746,N_9194);
or U10821 (N_10821,N_10062,N_10323);
and U10822 (N_10822,N_9443,N_9900);
and U10823 (N_10823,N_9140,N_10124);
and U10824 (N_10824,N_9739,N_9197);
nor U10825 (N_10825,N_9302,N_10300);
nor U10826 (N_10826,N_9457,N_10458);
xor U10827 (N_10827,N_9317,N_10049);
nor U10828 (N_10828,N_9439,N_9349);
nor U10829 (N_10829,N_9513,N_10452);
or U10830 (N_10830,N_9161,N_9646);
or U10831 (N_10831,N_10196,N_9258);
nor U10832 (N_10832,N_10132,N_9511);
nand U10833 (N_10833,N_10167,N_9452);
and U10834 (N_10834,N_9250,N_9602);
nor U10835 (N_10835,N_10250,N_10251);
and U10836 (N_10836,N_9757,N_9722);
or U10837 (N_10837,N_9186,N_10249);
or U10838 (N_10838,N_9003,N_9121);
or U10839 (N_10839,N_10048,N_9246);
nand U10840 (N_10840,N_9544,N_10076);
and U10841 (N_10841,N_9113,N_10061);
and U10842 (N_10842,N_10172,N_9115);
or U10843 (N_10843,N_9175,N_9814);
or U10844 (N_10844,N_9697,N_9832);
xnor U10845 (N_10845,N_9388,N_9801);
xnor U10846 (N_10846,N_10150,N_10273);
or U10847 (N_10847,N_9244,N_9829);
nor U10848 (N_10848,N_9291,N_9575);
nand U10849 (N_10849,N_9369,N_10151);
and U10850 (N_10850,N_9227,N_9767);
and U10851 (N_10851,N_9987,N_9412);
xor U10852 (N_10852,N_10098,N_9419);
and U10853 (N_10853,N_9989,N_9262);
or U10854 (N_10854,N_9740,N_9751);
xor U10855 (N_10855,N_9086,N_10360);
and U10856 (N_10856,N_9270,N_9990);
or U10857 (N_10857,N_10411,N_9147);
nor U10858 (N_10858,N_9375,N_10328);
and U10859 (N_10859,N_10270,N_9939);
nand U10860 (N_10860,N_10368,N_9660);
and U10861 (N_10861,N_9623,N_10313);
and U10862 (N_10862,N_9758,N_9879);
nor U10863 (N_10863,N_10230,N_10474);
nand U10864 (N_10864,N_9310,N_9505);
and U10865 (N_10865,N_9559,N_10092);
or U10866 (N_10866,N_10004,N_10084);
nor U10867 (N_10867,N_9842,N_9224);
xor U10868 (N_10868,N_9895,N_10414);
xnor U10869 (N_10869,N_9798,N_9000);
and U10870 (N_10870,N_9547,N_9770);
nand U10871 (N_10871,N_10214,N_10408);
nor U10872 (N_10872,N_9797,N_10189);
or U10873 (N_10873,N_9700,N_9094);
and U10874 (N_10874,N_10246,N_9519);
or U10875 (N_10875,N_9486,N_9201);
nor U10876 (N_10876,N_10467,N_10459);
and U10877 (N_10877,N_9206,N_10188);
nand U10878 (N_10878,N_9031,N_10024);
nor U10879 (N_10879,N_10295,N_9910);
and U10880 (N_10880,N_10156,N_9819);
xnor U10881 (N_10881,N_9837,N_10441);
nor U10882 (N_10882,N_9507,N_9640);
nor U10883 (N_10883,N_9207,N_9432);
nand U10884 (N_10884,N_9548,N_9385);
nor U10885 (N_10885,N_9567,N_9380);
nor U10886 (N_10886,N_10087,N_9659);
xnor U10887 (N_10887,N_9705,N_9846);
nor U10888 (N_10888,N_9845,N_9215);
and U10889 (N_10889,N_9228,N_10433);
and U10890 (N_10890,N_10291,N_9679);
and U10891 (N_10891,N_9276,N_9926);
nor U10892 (N_10892,N_9870,N_9812);
and U10893 (N_10893,N_9123,N_10395);
and U10894 (N_10894,N_9202,N_9083);
or U10895 (N_10895,N_9930,N_10261);
or U10896 (N_10896,N_9537,N_9022);
or U10897 (N_10897,N_9119,N_9551);
nor U10898 (N_10898,N_9356,N_10366);
and U10899 (N_10899,N_10312,N_9138);
xor U10900 (N_10900,N_10283,N_9885);
nor U10901 (N_10901,N_9120,N_9055);
nand U10902 (N_10902,N_10071,N_9972);
xor U10903 (N_10903,N_9753,N_9459);
nand U10904 (N_10904,N_10194,N_9264);
or U10905 (N_10905,N_9230,N_9967);
nor U10906 (N_10906,N_9691,N_9173);
nor U10907 (N_10907,N_9763,N_9009);
xnor U10908 (N_10908,N_10168,N_9054);
and U10909 (N_10909,N_10304,N_9463);
nand U10910 (N_10910,N_9726,N_9881);
nor U10911 (N_10911,N_9796,N_10404);
or U10912 (N_10912,N_10430,N_9821);
or U10913 (N_10913,N_9851,N_10031);
nand U10914 (N_10914,N_10387,N_9578);
and U10915 (N_10915,N_9808,N_9785);
xnor U10916 (N_10916,N_10333,N_9203);
nor U10917 (N_10917,N_9760,N_10445);
nand U10918 (N_10918,N_10381,N_9647);
nand U10919 (N_10919,N_9717,N_9688);
and U10920 (N_10920,N_9036,N_10171);
nand U10921 (N_10921,N_9982,N_10237);
xnor U10922 (N_10922,N_9060,N_9328);
or U10923 (N_10923,N_10180,N_9520);
nor U10924 (N_10924,N_9741,N_10021);
xnor U10925 (N_10925,N_10339,N_9863);
nand U10926 (N_10926,N_10073,N_9711);
or U10927 (N_10927,N_9154,N_9223);
xor U10928 (N_10928,N_10023,N_9472);
xor U10929 (N_10929,N_9240,N_10106);
or U10930 (N_10930,N_10453,N_9931);
or U10931 (N_10931,N_9500,N_9072);
nor U10932 (N_10932,N_10219,N_10205);
nand U10933 (N_10933,N_9071,N_9572);
nand U10934 (N_10934,N_9454,N_10482);
xor U10935 (N_10935,N_10184,N_9333);
and U10936 (N_10936,N_9915,N_9198);
xnor U10937 (N_10937,N_10297,N_9128);
and U10938 (N_10938,N_9833,N_9943);
nand U10939 (N_10939,N_9540,N_10271);
nand U10940 (N_10940,N_9718,N_9321);
or U10941 (N_10941,N_10078,N_9394);
nor U10942 (N_10942,N_10417,N_9082);
nand U10943 (N_10943,N_9523,N_10486);
or U10944 (N_10944,N_10352,N_10443);
and U10945 (N_10945,N_9748,N_9719);
or U10946 (N_10946,N_10320,N_10003);
and U10947 (N_10947,N_10462,N_10286);
xor U10948 (N_10948,N_10058,N_9237);
and U10949 (N_10949,N_9877,N_9667);
or U10950 (N_10950,N_9235,N_9800);
and U10951 (N_10951,N_9453,N_9543);
xor U10952 (N_10952,N_9284,N_9952);
nand U10953 (N_10953,N_9103,N_9836);
and U10954 (N_10954,N_10152,N_9880);
nand U10955 (N_10955,N_9749,N_9976);
nor U10956 (N_10956,N_9805,N_9672);
nand U10957 (N_10957,N_9830,N_9769);
nand U10958 (N_10958,N_10499,N_10470);
and U10959 (N_10959,N_9233,N_9859);
nor U10960 (N_10960,N_10066,N_10390);
and U10961 (N_10961,N_9581,N_9591);
xor U10962 (N_10962,N_9820,N_10178);
and U10963 (N_10963,N_9346,N_9628);
nand U10964 (N_10964,N_10255,N_10434);
nand U10965 (N_10965,N_9762,N_9143);
nor U10966 (N_10966,N_9890,N_10263);
and U10967 (N_10967,N_9788,N_9373);
xnor U10968 (N_10968,N_10309,N_10428);
nand U10969 (N_10969,N_9423,N_9840);
and U10970 (N_10970,N_9408,N_10435);
xor U10971 (N_10971,N_10439,N_9326);
nand U10972 (N_10972,N_10498,N_10190);
nor U10973 (N_10973,N_10086,N_9087);
nand U10974 (N_10974,N_10097,N_9686);
and U10975 (N_10975,N_10157,N_9488);
xnor U10976 (N_10976,N_9269,N_10162);
xor U10977 (N_10977,N_9509,N_9539);
nand U10978 (N_10978,N_9983,N_9390);
nor U10979 (N_10979,N_10425,N_9476);
or U10980 (N_10980,N_10397,N_9171);
nor U10981 (N_10981,N_10212,N_9066);
nor U10982 (N_10982,N_9973,N_10403);
nor U10983 (N_10983,N_10034,N_9074);
nor U10984 (N_10984,N_9018,N_10392);
xnor U10985 (N_10985,N_9216,N_9079);
and U10986 (N_10986,N_10301,N_9466);
or U10987 (N_10987,N_9069,N_9155);
and U10988 (N_10988,N_10356,N_9279);
xor U10989 (N_10989,N_9257,N_10293);
nand U10990 (N_10990,N_10202,N_9565);
nand U10991 (N_10991,N_10479,N_9436);
nand U10992 (N_10992,N_9723,N_9710);
or U10993 (N_10993,N_9381,N_9261);
nor U10994 (N_10994,N_10047,N_9025);
nor U10995 (N_10995,N_10169,N_9416);
xor U10996 (N_10996,N_9275,N_10008);
nor U10997 (N_10997,N_10247,N_10044);
and U10998 (N_10998,N_10285,N_9550);
or U10999 (N_10999,N_9906,N_9301);
nor U11000 (N_11000,N_10343,N_9610);
and U11001 (N_11001,N_10022,N_9620);
xnor U11002 (N_11002,N_9522,N_9950);
and U11003 (N_11003,N_10094,N_9601);
or U11004 (N_11004,N_9306,N_9397);
xor U11005 (N_11005,N_9743,N_9608);
nor U11006 (N_11006,N_10072,N_9402);
or U11007 (N_11007,N_9027,N_9313);
or U11008 (N_11008,N_9810,N_9125);
xor U11009 (N_11009,N_9428,N_9290);
or U11010 (N_11010,N_10043,N_9824);
nor U11011 (N_11011,N_10437,N_9391);
nand U11012 (N_11012,N_9557,N_9966);
nand U11013 (N_11013,N_9516,N_9985);
nand U11014 (N_11014,N_9866,N_9964);
xor U11015 (N_11015,N_9716,N_10265);
or U11016 (N_11016,N_9689,N_9387);
and U11017 (N_11017,N_9332,N_9008);
or U11018 (N_11018,N_10349,N_9062);
nor U11019 (N_11019,N_9477,N_9934);
or U11020 (N_11020,N_9485,N_10487);
nand U11021 (N_11021,N_9917,N_9043);
xor U11022 (N_11022,N_9727,N_10240);
or U11023 (N_11023,N_9606,N_9287);
and U11024 (N_11024,N_9465,N_9111);
and U11025 (N_11025,N_9888,N_9481);
or U11026 (N_11026,N_10121,N_10492);
nor U11027 (N_11027,N_9782,N_9970);
nor U11028 (N_11028,N_9148,N_9092);
nand U11029 (N_11029,N_9296,N_9089);
and U11030 (N_11030,N_10495,N_10018);
nor U11031 (N_11031,N_9724,N_9856);
and U11032 (N_11032,N_9850,N_9217);
nor U11033 (N_11033,N_10278,N_9670);
xor U11034 (N_11034,N_9592,N_9139);
nor U11035 (N_11035,N_9780,N_9536);
nor U11036 (N_11036,N_9447,N_9030);
and U11037 (N_11037,N_9834,N_9971);
nand U11038 (N_11038,N_9360,N_9156);
or U11039 (N_11039,N_9146,N_9393);
and U11040 (N_11040,N_9357,N_10446);
or U11041 (N_11041,N_10305,N_9100);
nor U11042 (N_11042,N_10154,N_9174);
or U11043 (N_11043,N_9133,N_9546);
xor U11044 (N_11044,N_10399,N_9024);
xor U11045 (N_11045,N_9553,N_9382);
xor U11046 (N_11046,N_10211,N_9791);
nor U11047 (N_11047,N_9145,N_9047);
or U11048 (N_11048,N_9429,N_10125);
or U11049 (N_11049,N_10472,N_9396);
or U11050 (N_11050,N_10036,N_9473);
nor U11051 (N_11051,N_9378,N_10400);
nor U11052 (N_11052,N_9211,N_9494);
nand U11053 (N_11053,N_9268,N_10155);
or U11054 (N_11054,N_9004,N_9673);
nand U11055 (N_11055,N_10222,N_9496);
nor U11056 (N_11056,N_9455,N_10477);
and U11057 (N_11057,N_9570,N_10371);
nand U11058 (N_11058,N_9621,N_9775);
nor U11059 (N_11059,N_9104,N_9534);
and U11060 (N_11060,N_9039,N_9483);
nor U11061 (N_11061,N_10158,N_9297);
or U11062 (N_11062,N_9444,N_9981);
xnor U11063 (N_11063,N_9399,N_9765);
nor U11064 (N_11064,N_9839,N_9527);
and U11065 (N_11065,N_10296,N_9153);
and U11066 (N_11066,N_9075,N_9566);
xor U11067 (N_11067,N_9179,N_10179);
or U11068 (N_11068,N_9530,N_9029);
and U11069 (N_11069,N_9734,N_9134);
or U11070 (N_11070,N_10317,N_9707);
xnor U11071 (N_11071,N_10233,N_9896);
nand U11072 (N_11072,N_9868,N_10065);
and U11073 (N_11073,N_9093,N_9324);
or U11074 (N_11074,N_10290,N_9042);
nor U11075 (N_11075,N_9611,N_10388);
and U11076 (N_11076,N_9909,N_10054);
and U11077 (N_11077,N_9600,N_10103);
nand U11078 (N_11078,N_9014,N_9159);
nand U11079 (N_11079,N_9157,N_10326);
xor U11080 (N_11080,N_9835,N_9376);
nand U11081 (N_11081,N_9144,N_10385);
or U11082 (N_11082,N_9656,N_10476);
and U11083 (N_11083,N_9561,N_9450);
or U11084 (N_11084,N_9681,N_9949);
nand U11085 (N_11085,N_9923,N_9102);
or U11086 (N_11086,N_10146,N_10119);
nand U11087 (N_11087,N_10269,N_9935);
nand U11088 (N_11088,N_9421,N_9956);
nand U11089 (N_11089,N_9642,N_9090);
and U11090 (N_11090,N_9662,N_10139);
nor U11091 (N_11091,N_9166,N_10318);
xor U11092 (N_11092,N_9918,N_10104);
or U11093 (N_11093,N_9799,N_10208);
or U11094 (N_11094,N_9315,N_9860);
nor U11095 (N_11095,N_10033,N_9200);
xor U11096 (N_11096,N_9882,N_10175);
xnor U11097 (N_11097,N_9916,N_9759);
or U11098 (N_11098,N_9160,N_9099);
nand U11099 (N_11099,N_10193,N_9940);
xor U11100 (N_11100,N_9051,N_10346);
nor U11101 (N_11101,N_10480,N_9847);
nand U11102 (N_11102,N_10030,N_9406);
xor U11103 (N_11103,N_9417,N_9383);
or U11104 (N_11104,N_9582,N_10245);
or U11105 (N_11105,N_10165,N_9823);
nor U11106 (N_11106,N_9995,N_10019);
and U11107 (N_11107,N_9521,N_10275);
and U11108 (N_11108,N_9542,N_10431);
nand U11109 (N_11109,N_9919,N_10081);
nor U11110 (N_11110,N_9441,N_9502);
xor U11111 (N_11111,N_10059,N_10451);
nand U11112 (N_11112,N_10241,N_9442);
nor U11113 (N_11113,N_9248,N_9162);
and U11114 (N_11114,N_9831,N_9529);
or U11115 (N_11115,N_9545,N_9135);
xor U11116 (N_11116,N_9422,N_9395);
or U11117 (N_11117,N_9320,N_10077);
nor U11118 (N_11118,N_9437,N_9126);
or U11119 (N_11119,N_9163,N_9781);
or U11120 (N_11120,N_10407,N_9650);
nor U11121 (N_11121,N_9771,N_10120);
and U11122 (N_11122,N_10370,N_9626);
or U11123 (N_11123,N_10455,N_10488);
or U11124 (N_11124,N_9786,N_10464);
nand U11125 (N_11125,N_10137,N_9414);
and U11126 (N_11126,N_9064,N_9622);
xnor U11127 (N_11127,N_9984,N_9779);
or U11128 (N_11128,N_9493,N_10310);
or U11129 (N_11129,N_9552,N_10063);
nor U11130 (N_11130,N_9012,N_9631);
nand U11131 (N_11131,N_10327,N_10463);
or U11132 (N_11132,N_9221,N_10248);
and U11133 (N_11133,N_10473,N_9980);
nor U11134 (N_11134,N_9308,N_10268);
and U11135 (N_11135,N_9026,N_9898);
nand U11136 (N_11136,N_10236,N_9708);
and U11137 (N_11137,N_10198,N_9474);
or U11138 (N_11138,N_10085,N_9506);
nand U11139 (N_11139,N_9809,N_9690);
nand U11140 (N_11140,N_10367,N_9225);
or U11141 (N_11141,N_9445,N_9168);
nor U11142 (N_11142,N_9489,N_9041);
xor U11143 (N_11143,N_9703,N_9298);
nand U11144 (N_11144,N_10153,N_9404);
nor U11145 (N_11145,N_10130,N_10374);
nand U11146 (N_11146,N_9873,N_10396);
and U11147 (N_11147,N_10418,N_10001);
nor U11148 (N_11148,N_10267,N_9894);
or U11149 (N_11149,N_9714,N_10100);
xnor U11150 (N_11150,N_10440,N_9962);
or U11151 (N_11151,N_10242,N_9957);
and U11152 (N_11152,N_9208,N_9372);
nor U11153 (N_11153,N_10401,N_9409);
or U11154 (N_11154,N_10442,N_9617);
or U11155 (N_11155,N_9501,N_9577);
or U11156 (N_11156,N_9288,N_9752);
and U11157 (N_11157,N_9979,N_10485);
nand U11158 (N_11158,N_9451,N_9181);
nand U11159 (N_11159,N_10113,N_10112);
xnor U11160 (N_11160,N_9231,N_10380);
and U11161 (N_11161,N_10340,N_10475);
or U11162 (N_11162,N_9101,N_9848);
or U11163 (N_11163,N_9359,N_9475);
xor U11164 (N_11164,N_9413,N_9058);
nand U11165 (N_11165,N_9325,N_9497);
xor U11166 (N_11166,N_9229,N_9304);
nor U11167 (N_11167,N_10038,N_9193);
or U11168 (N_11168,N_10324,N_9366);
xnor U11169 (N_11169,N_9538,N_9081);
or U11170 (N_11170,N_10035,N_10074);
xor U11171 (N_11171,N_10365,N_9764);
nor U11172 (N_11172,N_9185,N_10045);
nand U11173 (N_11173,N_9068,N_9637);
xnor U11174 (N_11174,N_10064,N_9400);
xnor U11175 (N_11175,N_9872,N_9535);
xnor U11176 (N_11176,N_9078,N_9190);
xnor U11177 (N_11177,N_9343,N_10221);
and U11178 (N_11178,N_10089,N_9795);
xnor U11179 (N_11179,N_9218,N_9255);
or U11180 (N_11180,N_9005,N_10013);
or U11181 (N_11181,N_9219,N_9222);
xor U11182 (N_11182,N_9131,N_10014);
or U11183 (N_11183,N_9352,N_9712);
nor U11184 (N_11184,N_9433,N_9902);
nor U11185 (N_11185,N_10244,N_9517);
or U11186 (N_11186,N_9259,N_9377);
nor U11187 (N_11187,N_10060,N_9045);
xnor U11188 (N_11188,N_9725,N_9736);
xnor U11189 (N_11189,N_9747,N_9337);
or U11190 (N_11190,N_10262,N_9807);
or U11191 (N_11191,N_10010,N_9426);
nor U11192 (N_11192,N_10228,N_9448);
nor U11193 (N_11193,N_9912,N_9142);
nand U11194 (N_11194,N_9920,N_9905);
nor U11195 (N_11195,N_9789,N_9806);
nand U11196 (N_11196,N_10345,N_10015);
nand U11197 (N_11197,N_10011,N_9674);
and U11198 (N_11198,N_10217,N_10140);
nand U11199 (N_11199,N_10481,N_10053);
and U11200 (N_11200,N_9549,N_10299);
nor U11201 (N_11201,N_9323,N_9151);
or U11202 (N_11202,N_10336,N_9528);
nand U11203 (N_11203,N_9363,N_9418);
and U11204 (N_11204,N_10449,N_9379);
nand U11205 (N_11205,N_10117,N_9720);
nand U11206 (N_11206,N_9766,N_9618);
xor U11207 (N_11207,N_10415,N_9515);
xor U11208 (N_11208,N_9424,N_9361);
and U11209 (N_11209,N_9968,N_9319);
nor U11210 (N_11210,N_9625,N_9091);
nor U11211 (N_11211,N_9183,N_9471);
xor U11212 (N_11212,N_10478,N_9590);
nand U11213 (N_11213,N_10419,N_9893);
and U11214 (N_11214,N_9822,N_9035);
nand U11215 (N_11215,N_9908,N_9652);
and U11216 (N_11216,N_9110,N_10069);
and U11217 (N_11217,N_9817,N_10042);
and U11218 (N_11218,N_9017,N_10344);
nor U11219 (N_11219,N_9188,N_9562);
and U11220 (N_11220,N_9607,N_9046);
xnor U11221 (N_11221,N_9277,N_10145);
or U11222 (N_11222,N_9633,N_10426);
nand U11223 (N_11223,N_9067,N_9586);
xnor U11224 (N_11224,N_9149,N_9884);
xor U11225 (N_11225,N_9630,N_9665);
or U11226 (N_11226,N_9733,N_10496);
nor U11227 (N_11227,N_10207,N_9609);
and U11228 (N_11228,N_10280,N_9875);
nor U11229 (N_11229,N_9405,N_9680);
or U11230 (N_11230,N_9721,N_10466);
xnor U11231 (N_11231,N_9114,N_10277);
nor U11232 (N_11232,N_9056,N_9518);
nor U11233 (N_11233,N_9023,N_9330);
nand U11234 (N_11234,N_9958,N_10000);
nand U11235 (N_11235,N_10122,N_9921);
xnor U11236 (N_11236,N_9491,N_9654);
xor U11237 (N_11237,N_9693,N_9052);
and U11238 (N_11238,N_9666,N_10338);
nor U11239 (N_11239,N_10020,N_9576);
nand U11240 (N_11240,N_9684,N_9899);
xor U11241 (N_11241,N_10016,N_9938);
and U11242 (N_11242,N_9913,N_9658);
and U11243 (N_11243,N_9176,N_9871);
nor U11244 (N_11244,N_10361,N_9112);
nor U11245 (N_11245,N_9172,N_9431);
and U11246 (N_11246,N_9510,N_10055);
nor U11247 (N_11247,N_9249,N_10224);
or U11248 (N_11248,N_9541,N_10239);
nand U11249 (N_11249,N_10460,N_10083);
or U11250 (N_11250,N_9496,N_9514);
xor U11251 (N_11251,N_9626,N_10447);
or U11252 (N_11252,N_9846,N_10057);
nand U11253 (N_11253,N_10124,N_10087);
nand U11254 (N_11254,N_9274,N_10462);
and U11255 (N_11255,N_10274,N_9049);
xor U11256 (N_11256,N_9423,N_9999);
or U11257 (N_11257,N_10234,N_10253);
nor U11258 (N_11258,N_9755,N_10232);
nand U11259 (N_11259,N_10266,N_10074);
xnor U11260 (N_11260,N_10467,N_10077);
xnor U11261 (N_11261,N_10030,N_9573);
nor U11262 (N_11262,N_9871,N_10463);
nor U11263 (N_11263,N_9521,N_10435);
xnor U11264 (N_11264,N_9286,N_9642);
xnor U11265 (N_11265,N_9234,N_9187);
and U11266 (N_11266,N_9399,N_9214);
and U11267 (N_11267,N_9798,N_9369);
nand U11268 (N_11268,N_9685,N_10154);
and U11269 (N_11269,N_10454,N_10199);
or U11270 (N_11270,N_9854,N_10134);
or U11271 (N_11271,N_9679,N_9193);
or U11272 (N_11272,N_10316,N_10355);
xnor U11273 (N_11273,N_9955,N_9232);
xnor U11274 (N_11274,N_10069,N_9273);
or U11275 (N_11275,N_9848,N_9595);
nor U11276 (N_11276,N_9900,N_9359);
or U11277 (N_11277,N_9012,N_9883);
nand U11278 (N_11278,N_9706,N_9393);
or U11279 (N_11279,N_9574,N_9828);
nand U11280 (N_11280,N_9223,N_9066);
xor U11281 (N_11281,N_9438,N_9627);
xnor U11282 (N_11282,N_9511,N_10302);
or U11283 (N_11283,N_10050,N_10206);
or U11284 (N_11284,N_9455,N_9418);
or U11285 (N_11285,N_10428,N_9428);
xnor U11286 (N_11286,N_9697,N_9790);
xnor U11287 (N_11287,N_9773,N_9124);
or U11288 (N_11288,N_9005,N_9058);
xnor U11289 (N_11289,N_10498,N_9825);
and U11290 (N_11290,N_10124,N_10237);
and U11291 (N_11291,N_9586,N_9661);
nand U11292 (N_11292,N_9293,N_10379);
or U11293 (N_11293,N_9554,N_9168);
or U11294 (N_11294,N_9067,N_10136);
nor U11295 (N_11295,N_9913,N_9084);
nand U11296 (N_11296,N_10227,N_9006);
nor U11297 (N_11297,N_10466,N_10292);
or U11298 (N_11298,N_10365,N_10467);
nand U11299 (N_11299,N_9108,N_10422);
and U11300 (N_11300,N_9877,N_9494);
nand U11301 (N_11301,N_9805,N_9391);
nor U11302 (N_11302,N_9408,N_9393);
or U11303 (N_11303,N_9521,N_9934);
nand U11304 (N_11304,N_10115,N_9067);
nand U11305 (N_11305,N_10167,N_10370);
nand U11306 (N_11306,N_10466,N_9830);
and U11307 (N_11307,N_9225,N_10271);
and U11308 (N_11308,N_9841,N_9463);
xor U11309 (N_11309,N_10464,N_9375);
nand U11310 (N_11310,N_9184,N_9316);
or U11311 (N_11311,N_9438,N_9954);
xnor U11312 (N_11312,N_9441,N_9397);
nor U11313 (N_11313,N_9474,N_10206);
or U11314 (N_11314,N_9611,N_9452);
nand U11315 (N_11315,N_9494,N_10026);
or U11316 (N_11316,N_10488,N_10471);
xnor U11317 (N_11317,N_10120,N_10348);
nand U11318 (N_11318,N_9299,N_9597);
or U11319 (N_11319,N_9399,N_9960);
or U11320 (N_11320,N_9615,N_9738);
and U11321 (N_11321,N_10187,N_10001);
nor U11322 (N_11322,N_9561,N_9891);
nand U11323 (N_11323,N_9468,N_9372);
xnor U11324 (N_11324,N_9207,N_9239);
xnor U11325 (N_11325,N_10340,N_9204);
xor U11326 (N_11326,N_10420,N_9439);
and U11327 (N_11327,N_9197,N_9935);
nand U11328 (N_11328,N_9278,N_10011);
nor U11329 (N_11329,N_10045,N_9918);
and U11330 (N_11330,N_9590,N_9506);
and U11331 (N_11331,N_10343,N_9694);
nand U11332 (N_11332,N_9540,N_9601);
xor U11333 (N_11333,N_9461,N_10053);
nand U11334 (N_11334,N_9856,N_9616);
xnor U11335 (N_11335,N_10256,N_9390);
xnor U11336 (N_11336,N_10121,N_10405);
and U11337 (N_11337,N_9397,N_9094);
xor U11338 (N_11338,N_9806,N_10420);
and U11339 (N_11339,N_10183,N_9612);
and U11340 (N_11340,N_10218,N_9052);
and U11341 (N_11341,N_9702,N_9022);
nand U11342 (N_11342,N_9923,N_9116);
nand U11343 (N_11343,N_9439,N_10220);
and U11344 (N_11344,N_9817,N_10038);
or U11345 (N_11345,N_9058,N_9040);
or U11346 (N_11346,N_9925,N_9946);
xnor U11347 (N_11347,N_9886,N_9373);
xor U11348 (N_11348,N_9800,N_10033);
nor U11349 (N_11349,N_9638,N_9363);
and U11350 (N_11350,N_10248,N_9069);
or U11351 (N_11351,N_10445,N_9197);
nand U11352 (N_11352,N_9137,N_9505);
nor U11353 (N_11353,N_9892,N_10286);
and U11354 (N_11354,N_9263,N_9202);
nand U11355 (N_11355,N_10390,N_9842);
xnor U11356 (N_11356,N_9922,N_9762);
nor U11357 (N_11357,N_10443,N_9031);
nand U11358 (N_11358,N_9296,N_9377);
nor U11359 (N_11359,N_10441,N_10278);
nand U11360 (N_11360,N_10202,N_9077);
nand U11361 (N_11361,N_10340,N_10047);
and U11362 (N_11362,N_9803,N_9002);
nand U11363 (N_11363,N_9041,N_10168);
and U11364 (N_11364,N_10499,N_9745);
xor U11365 (N_11365,N_9095,N_9521);
or U11366 (N_11366,N_10471,N_10469);
nor U11367 (N_11367,N_10430,N_10490);
and U11368 (N_11368,N_10453,N_10434);
nand U11369 (N_11369,N_10164,N_9682);
nor U11370 (N_11370,N_10426,N_10447);
xor U11371 (N_11371,N_10150,N_9271);
or U11372 (N_11372,N_10156,N_10444);
or U11373 (N_11373,N_9343,N_9912);
nand U11374 (N_11374,N_10360,N_9739);
xnor U11375 (N_11375,N_9746,N_9201);
and U11376 (N_11376,N_9014,N_9440);
xnor U11377 (N_11377,N_9035,N_9282);
nand U11378 (N_11378,N_10214,N_9340);
xor U11379 (N_11379,N_9854,N_9857);
xnor U11380 (N_11380,N_10037,N_9902);
or U11381 (N_11381,N_9888,N_9103);
and U11382 (N_11382,N_9325,N_10243);
nor U11383 (N_11383,N_10168,N_10440);
xnor U11384 (N_11384,N_9330,N_9509);
nand U11385 (N_11385,N_10260,N_9180);
nand U11386 (N_11386,N_9874,N_10245);
xnor U11387 (N_11387,N_9140,N_9130);
and U11388 (N_11388,N_9292,N_9472);
nand U11389 (N_11389,N_9186,N_9767);
nand U11390 (N_11390,N_10390,N_9221);
or U11391 (N_11391,N_9003,N_9715);
or U11392 (N_11392,N_9746,N_9984);
nand U11393 (N_11393,N_9837,N_10475);
or U11394 (N_11394,N_10364,N_9128);
xnor U11395 (N_11395,N_9263,N_9660);
and U11396 (N_11396,N_10006,N_9504);
and U11397 (N_11397,N_10154,N_10398);
and U11398 (N_11398,N_9825,N_9846);
and U11399 (N_11399,N_10242,N_10141);
nand U11400 (N_11400,N_9822,N_9469);
xor U11401 (N_11401,N_9068,N_9766);
nor U11402 (N_11402,N_9070,N_9163);
and U11403 (N_11403,N_9758,N_9190);
xor U11404 (N_11404,N_10346,N_9471);
and U11405 (N_11405,N_10247,N_10167);
nor U11406 (N_11406,N_9832,N_9853);
xnor U11407 (N_11407,N_9839,N_9075);
nand U11408 (N_11408,N_9407,N_10035);
or U11409 (N_11409,N_9352,N_9750);
and U11410 (N_11410,N_9829,N_9691);
xnor U11411 (N_11411,N_9746,N_10259);
nand U11412 (N_11412,N_10495,N_10388);
nand U11413 (N_11413,N_9636,N_10345);
xnor U11414 (N_11414,N_9428,N_9493);
and U11415 (N_11415,N_9537,N_10297);
or U11416 (N_11416,N_9974,N_9565);
nand U11417 (N_11417,N_10143,N_9649);
nand U11418 (N_11418,N_9928,N_9023);
and U11419 (N_11419,N_9576,N_10182);
or U11420 (N_11420,N_9432,N_10455);
nand U11421 (N_11421,N_9991,N_9854);
nor U11422 (N_11422,N_9759,N_9145);
or U11423 (N_11423,N_9770,N_9247);
xor U11424 (N_11424,N_9635,N_10476);
or U11425 (N_11425,N_9957,N_10183);
xor U11426 (N_11426,N_9048,N_10026);
nand U11427 (N_11427,N_9786,N_10253);
xnor U11428 (N_11428,N_10483,N_10184);
or U11429 (N_11429,N_10278,N_10199);
and U11430 (N_11430,N_9338,N_9935);
nor U11431 (N_11431,N_9863,N_10183);
or U11432 (N_11432,N_10458,N_10034);
or U11433 (N_11433,N_9406,N_10138);
nor U11434 (N_11434,N_9948,N_10339);
or U11435 (N_11435,N_10344,N_10351);
nand U11436 (N_11436,N_10144,N_9935);
or U11437 (N_11437,N_10326,N_10232);
or U11438 (N_11438,N_9102,N_10075);
or U11439 (N_11439,N_10163,N_9561);
or U11440 (N_11440,N_10337,N_9715);
or U11441 (N_11441,N_10044,N_9650);
and U11442 (N_11442,N_9256,N_10464);
nor U11443 (N_11443,N_10431,N_9027);
and U11444 (N_11444,N_10188,N_9685);
xnor U11445 (N_11445,N_9284,N_9827);
nand U11446 (N_11446,N_9563,N_10033);
and U11447 (N_11447,N_9331,N_9561);
and U11448 (N_11448,N_9371,N_9614);
and U11449 (N_11449,N_9624,N_10376);
and U11450 (N_11450,N_10045,N_10054);
nand U11451 (N_11451,N_9942,N_9556);
and U11452 (N_11452,N_10416,N_9278);
and U11453 (N_11453,N_10247,N_9849);
nor U11454 (N_11454,N_9396,N_9802);
nor U11455 (N_11455,N_10382,N_9472);
xnor U11456 (N_11456,N_9232,N_9627);
nor U11457 (N_11457,N_10050,N_9772);
and U11458 (N_11458,N_9231,N_9540);
and U11459 (N_11459,N_9625,N_9444);
nor U11460 (N_11460,N_10365,N_10344);
and U11461 (N_11461,N_10408,N_9507);
and U11462 (N_11462,N_9747,N_9505);
and U11463 (N_11463,N_10161,N_9263);
nand U11464 (N_11464,N_10213,N_9439);
or U11465 (N_11465,N_9740,N_9585);
or U11466 (N_11466,N_9268,N_9581);
nor U11467 (N_11467,N_9836,N_10138);
nor U11468 (N_11468,N_9587,N_9289);
nor U11469 (N_11469,N_9753,N_9108);
nor U11470 (N_11470,N_9421,N_9012);
nor U11471 (N_11471,N_9594,N_9712);
nand U11472 (N_11472,N_9162,N_9056);
and U11473 (N_11473,N_9615,N_9271);
nand U11474 (N_11474,N_10247,N_9114);
and U11475 (N_11475,N_9100,N_9979);
nand U11476 (N_11476,N_10215,N_9461);
or U11477 (N_11477,N_9308,N_9078);
nor U11478 (N_11478,N_10007,N_9761);
xnor U11479 (N_11479,N_9171,N_10144);
or U11480 (N_11480,N_9505,N_10118);
xor U11481 (N_11481,N_9633,N_10450);
nor U11482 (N_11482,N_9824,N_9287);
and U11483 (N_11483,N_9422,N_9881);
and U11484 (N_11484,N_9722,N_9549);
nor U11485 (N_11485,N_9014,N_9221);
xor U11486 (N_11486,N_9086,N_9673);
xor U11487 (N_11487,N_10439,N_9238);
or U11488 (N_11488,N_9403,N_10491);
nand U11489 (N_11489,N_9418,N_10171);
nand U11490 (N_11490,N_9981,N_9050);
nand U11491 (N_11491,N_10436,N_9996);
or U11492 (N_11492,N_9494,N_9638);
and U11493 (N_11493,N_10404,N_9268);
and U11494 (N_11494,N_9393,N_10408);
or U11495 (N_11495,N_10208,N_10414);
nand U11496 (N_11496,N_10245,N_9919);
nand U11497 (N_11497,N_9941,N_10388);
xor U11498 (N_11498,N_10149,N_9750);
xor U11499 (N_11499,N_9664,N_9140);
nor U11500 (N_11500,N_10452,N_9519);
and U11501 (N_11501,N_9001,N_9168);
xnor U11502 (N_11502,N_10484,N_9506);
nor U11503 (N_11503,N_10102,N_10060);
nor U11504 (N_11504,N_9032,N_10001);
xor U11505 (N_11505,N_9888,N_9736);
nor U11506 (N_11506,N_9128,N_10397);
or U11507 (N_11507,N_9969,N_9925);
or U11508 (N_11508,N_10136,N_10311);
and U11509 (N_11509,N_10105,N_9314);
and U11510 (N_11510,N_10261,N_10465);
nand U11511 (N_11511,N_10149,N_9555);
nor U11512 (N_11512,N_10002,N_10401);
nor U11513 (N_11513,N_10219,N_10427);
xor U11514 (N_11514,N_9147,N_9318);
nor U11515 (N_11515,N_9591,N_9419);
or U11516 (N_11516,N_10242,N_9438);
and U11517 (N_11517,N_9845,N_10254);
xor U11518 (N_11518,N_9257,N_10371);
nor U11519 (N_11519,N_9901,N_9200);
and U11520 (N_11520,N_10353,N_10080);
nor U11521 (N_11521,N_10153,N_9545);
nor U11522 (N_11522,N_9803,N_9449);
and U11523 (N_11523,N_9027,N_9172);
nor U11524 (N_11524,N_10145,N_9816);
xnor U11525 (N_11525,N_10247,N_9139);
xnor U11526 (N_11526,N_10193,N_9529);
nand U11527 (N_11527,N_9543,N_10009);
xnor U11528 (N_11528,N_10454,N_9081);
nand U11529 (N_11529,N_10302,N_10338);
xnor U11530 (N_11530,N_9588,N_9358);
or U11531 (N_11531,N_10435,N_10138);
and U11532 (N_11532,N_10090,N_9051);
xor U11533 (N_11533,N_9386,N_10340);
nand U11534 (N_11534,N_9756,N_9211);
nand U11535 (N_11535,N_10447,N_10146);
and U11536 (N_11536,N_9352,N_9435);
nor U11537 (N_11537,N_9278,N_10031);
and U11538 (N_11538,N_9089,N_9070);
or U11539 (N_11539,N_9815,N_9473);
nand U11540 (N_11540,N_10104,N_9638);
or U11541 (N_11541,N_10450,N_10186);
and U11542 (N_11542,N_9957,N_10406);
nand U11543 (N_11543,N_10164,N_9452);
or U11544 (N_11544,N_9696,N_9265);
xor U11545 (N_11545,N_10018,N_9884);
nor U11546 (N_11546,N_9487,N_10133);
or U11547 (N_11547,N_9612,N_10148);
or U11548 (N_11548,N_9919,N_9508);
or U11549 (N_11549,N_9390,N_9972);
xor U11550 (N_11550,N_9774,N_10418);
nand U11551 (N_11551,N_9142,N_9144);
and U11552 (N_11552,N_9181,N_10221);
xor U11553 (N_11553,N_10015,N_9062);
and U11554 (N_11554,N_9239,N_10375);
xnor U11555 (N_11555,N_9505,N_9937);
nor U11556 (N_11556,N_9533,N_9114);
xnor U11557 (N_11557,N_9363,N_9663);
xnor U11558 (N_11558,N_9799,N_9892);
or U11559 (N_11559,N_10484,N_10034);
or U11560 (N_11560,N_9123,N_9425);
nor U11561 (N_11561,N_9242,N_10032);
nor U11562 (N_11562,N_9310,N_9532);
nand U11563 (N_11563,N_9926,N_9709);
xnor U11564 (N_11564,N_10274,N_10198);
and U11565 (N_11565,N_9269,N_9349);
nand U11566 (N_11566,N_10103,N_9049);
or U11567 (N_11567,N_9103,N_9253);
nor U11568 (N_11568,N_9229,N_10143);
xnor U11569 (N_11569,N_9176,N_9205);
or U11570 (N_11570,N_10322,N_9755);
and U11571 (N_11571,N_9517,N_10364);
nor U11572 (N_11572,N_9205,N_9669);
or U11573 (N_11573,N_9092,N_9130);
or U11574 (N_11574,N_9436,N_9358);
and U11575 (N_11575,N_9407,N_9871);
nor U11576 (N_11576,N_9361,N_9266);
or U11577 (N_11577,N_9620,N_9242);
nor U11578 (N_11578,N_10229,N_9580);
xnor U11579 (N_11579,N_10116,N_9967);
or U11580 (N_11580,N_9903,N_9158);
xnor U11581 (N_11581,N_9512,N_9510);
or U11582 (N_11582,N_10338,N_9401);
nor U11583 (N_11583,N_10169,N_10470);
and U11584 (N_11584,N_9721,N_9241);
nor U11585 (N_11585,N_10325,N_9816);
and U11586 (N_11586,N_10068,N_10483);
or U11587 (N_11587,N_10164,N_9576);
xor U11588 (N_11588,N_10106,N_9990);
nor U11589 (N_11589,N_9742,N_9495);
nand U11590 (N_11590,N_10483,N_10288);
xor U11591 (N_11591,N_10224,N_10382);
or U11592 (N_11592,N_10338,N_9361);
nor U11593 (N_11593,N_9872,N_9990);
nor U11594 (N_11594,N_10473,N_10121);
and U11595 (N_11595,N_10498,N_9452);
and U11596 (N_11596,N_10198,N_10152);
or U11597 (N_11597,N_10366,N_9660);
and U11598 (N_11598,N_9542,N_10019);
or U11599 (N_11599,N_10374,N_9412);
nor U11600 (N_11600,N_9873,N_9227);
or U11601 (N_11601,N_9077,N_10050);
and U11602 (N_11602,N_10348,N_10164);
nor U11603 (N_11603,N_9438,N_9469);
and U11604 (N_11604,N_9797,N_10245);
nor U11605 (N_11605,N_9723,N_9352);
and U11606 (N_11606,N_9140,N_9193);
and U11607 (N_11607,N_9427,N_9578);
nand U11608 (N_11608,N_10059,N_9683);
xnor U11609 (N_11609,N_9090,N_10483);
or U11610 (N_11610,N_9572,N_9662);
nor U11611 (N_11611,N_9062,N_10403);
nand U11612 (N_11612,N_9471,N_9024);
or U11613 (N_11613,N_10318,N_9302);
and U11614 (N_11614,N_9501,N_10229);
nand U11615 (N_11615,N_10466,N_10108);
or U11616 (N_11616,N_10324,N_9665);
or U11617 (N_11617,N_9950,N_10024);
nand U11618 (N_11618,N_9098,N_9864);
or U11619 (N_11619,N_9116,N_9630);
xor U11620 (N_11620,N_9362,N_10165);
and U11621 (N_11621,N_10438,N_9858);
nor U11622 (N_11622,N_9947,N_10126);
and U11623 (N_11623,N_9413,N_9934);
nor U11624 (N_11624,N_10480,N_10088);
nand U11625 (N_11625,N_9973,N_9821);
xnor U11626 (N_11626,N_9978,N_9482);
xor U11627 (N_11627,N_9554,N_9832);
nor U11628 (N_11628,N_9265,N_9667);
nand U11629 (N_11629,N_10236,N_9072);
or U11630 (N_11630,N_9736,N_9636);
nor U11631 (N_11631,N_10476,N_9650);
or U11632 (N_11632,N_9662,N_10144);
nand U11633 (N_11633,N_10089,N_10023);
nand U11634 (N_11634,N_9942,N_9605);
nor U11635 (N_11635,N_10328,N_9340);
or U11636 (N_11636,N_10142,N_9902);
or U11637 (N_11637,N_9657,N_9540);
or U11638 (N_11638,N_9767,N_9626);
and U11639 (N_11639,N_9896,N_9839);
or U11640 (N_11640,N_9855,N_9945);
and U11641 (N_11641,N_10253,N_9177);
nand U11642 (N_11642,N_9502,N_9733);
xor U11643 (N_11643,N_9638,N_10379);
xor U11644 (N_11644,N_10356,N_9287);
nand U11645 (N_11645,N_9097,N_9577);
nand U11646 (N_11646,N_9609,N_10418);
or U11647 (N_11647,N_9477,N_9849);
xor U11648 (N_11648,N_9974,N_9343);
nand U11649 (N_11649,N_9265,N_9025);
and U11650 (N_11650,N_9211,N_9736);
or U11651 (N_11651,N_10014,N_9741);
or U11652 (N_11652,N_10305,N_10212);
xnor U11653 (N_11653,N_9487,N_9909);
xnor U11654 (N_11654,N_9223,N_10199);
and U11655 (N_11655,N_9351,N_10367);
and U11656 (N_11656,N_9752,N_10217);
and U11657 (N_11657,N_9815,N_9585);
and U11658 (N_11658,N_9449,N_9091);
nor U11659 (N_11659,N_9929,N_9396);
nand U11660 (N_11660,N_9771,N_9471);
nor U11661 (N_11661,N_9330,N_9941);
xnor U11662 (N_11662,N_9633,N_9084);
and U11663 (N_11663,N_9529,N_10483);
nand U11664 (N_11664,N_9852,N_9296);
nand U11665 (N_11665,N_10047,N_9296);
nand U11666 (N_11666,N_10358,N_9412);
or U11667 (N_11667,N_10431,N_9682);
nor U11668 (N_11668,N_9021,N_9881);
xnor U11669 (N_11669,N_9663,N_10048);
and U11670 (N_11670,N_10165,N_10068);
nand U11671 (N_11671,N_9762,N_9035);
and U11672 (N_11672,N_10304,N_10301);
and U11673 (N_11673,N_9411,N_9679);
and U11674 (N_11674,N_10207,N_9418);
xnor U11675 (N_11675,N_9244,N_10019);
or U11676 (N_11676,N_9491,N_9250);
nor U11677 (N_11677,N_9726,N_9929);
and U11678 (N_11678,N_9096,N_9157);
nand U11679 (N_11679,N_10401,N_9405);
nand U11680 (N_11680,N_10327,N_9354);
xor U11681 (N_11681,N_9541,N_9300);
or U11682 (N_11682,N_9079,N_9362);
and U11683 (N_11683,N_10101,N_10163);
xnor U11684 (N_11684,N_9198,N_10443);
nand U11685 (N_11685,N_9742,N_9207);
or U11686 (N_11686,N_9105,N_9560);
nor U11687 (N_11687,N_9202,N_9859);
or U11688 (N_11688,N_10492,N_9664);
and U11689 (N_11689,N_9353,N_10281);
or U11690 (N_11690,N_10172,N_9359);
nand U11691 (N_11691,N_9576,N_10106);
nand U11692 (N_11692,N_10303,N_9200);
xor U11693 (N_11693,N_10011,N_9337);
nand U11694 (N_11694,N_9690,N_9273);
and U11695 (N_11695,N_9907,N_9501);
xor U11696 (N_11696,N_9678,N_9079);
nand U11697 (N_11697,N_9144,N_10206);
and U11698 (N_11698,N_9993,N_9803);
nand U11699 (N_11699,N_9778,N_10440);
nand U11700 (N_11700,N_9789,N_10029);
or U11701 (N_11701,N_10240,N_9428);
nand U11702 (N_11702,N_9796,N_9205);
and U11703 (N_11703,N_9816,N_9782);
or U11704 (N_11704,N_9975,N_10161);
and U11705 (N_11705,N_9819,N_9611);
nor U11706 (N_11706,N_9218,N_10359);
or U11707 (N_11707,N_10451,N_10411);
nand U11708 (N_11708,N_9814,N_10012);
xnor U11709 (N_11709,N_9021,N_9383);
xor U11710 (N_11710,N_9941,N_9317);
nand U11711 (N_11711,N_10068,N_10210);
or U11712 (N_11712,N_9146,N_9945);
or U11713 (N_11713,N_9466,N_9742);
or U11714 (N_11714,N_10326,N_9878);
and U11715 (N_11715,N_10067,N_9661);
nor U11716 (N_11716,N_9955,N_9304);
nand U11717 (N_11717,N_9178,N_9165);
nor U11718 (N_11718,N_9607,N_9071);
or U11719 (N_11719,N_9386,N_9807);
or U11720 (N_11720,N_9603,N_10491);
nand U11721 (N_11721,N_10381,N_9433);
xnor U11722 (N_11722,N_9857,N_10072);
nor U11723 (N_11723,N_10203,N_9379);
and U11724 (N_11724,N_10298,N_9586);
and U11725 (N_11725,N_9495,N_10338);
nor U11726 (N_11726,N_9781,N_10047);
nand U11727 (N_11727,N_10408,N_9814);
nor U11728 (N_11728,N_9233,N_9201);
nor U11729 (N_11729,N_10018,N_10052);
and U11730 (N_11730,N_9298,N_9137);
and U11731 (N_11731,N_10225,N_10350);
xor U11732 (N_11732,N_10285,N_9487);
nor U11733 (N_11733,N_10213,N_9696);
or U11734 (N_11734,N_9519,N_9870);
nor U11735 (N_11735,N_10337,N_9060);
xor U11736 (N_11736,N_10172,N_9209);
xnor U11737 (N_11737,N_9810,N_10326);
or U11738 (N_11738,N_9474,N_9790);
nor U11739 (N_11739,N_10302,N_9067);
xor U11740 (N_11740,N_9345,N_9761);
or U11741 (N_11741,N_9812,N_10310);
or U11742 (N_11742,N_9379,N_10017);
nor U11743 (N_11743,N_9851,N_9451);
xnor U11744 (N_11744,N_9872,N_9095);
or U11745 (N_11745,N_10061,N_9886);
nand U11746 (N_11746,N_10192,N_9025);
or U11747 (N_11747,N_9260,N_9418);
nor U11748 (N_11748,N_9561,N_9382);
or U11749 (N_11749,N_9417,N_10173);
xnor U11750 (N_11750,N_10414,N_9631);
or U11751 (N_11751,N_10492,N_9607);
nand U11752 (N_11752,N_10268,N_9581);
nor U11753 (N_11753,N_10465,N_10375);
or U11754 (N_11754,N_9292,N_9591);
or U11755 (N_11755,N_10399,N_9892);
nor U11756 (N_11756,N_9266,N_9512);
nand U11757 (N_11757,N_9846,N_9860);
and U11758 (N_11758,N_9400,N_9229);
or U11759 (N_11759,N_10449,N_9963);
or U11760 (N_11760,N_10319,N_9967);
or U11761 (N_11761,N_9048,N_9946);
nand U11762 (N_11762,N_9767,N_9013);
and U11763 (N_11763,N_9242,N_9633);
nand U11764 (N_11764,N_10372,N_10259);
xor U11765 (N_11765,N_10447,N_9618);
and U11766 (N_11766,N_9523,N_9599);
or U11767 (N_11767,N_9053,N_9981);
xor U11768 (N_11768,N_10397,N_10262);
nand U11769 (N_11769,N_9989,N_10458);
or U11770 (N_11770,N_9169,N_9450);
xor U11771 (N_11771,N_9772,N_10286);
xnor U11772 (N_11772,N_10109,N_10344);
or U11773 (N_11773,N_9458,N_10216);
nor U11774 (N_11774,N_9725,N_9628);
or U11775 (N_11775,N_10401,N_9151);
and U11776 (N_11776,N_9165,N_9886);
or U11777 (N_11777,N_9440,N_9149);
nand U11778 (N_11778,N_9972,N_9368);
nor U11779 (N_11779,N_9519,N_10055);
xor U11780 (N_11780,N_10435,N_9581);
nand U11781 (N_11781,N_10115,N_9669);
nand U11782 (N_11782,N_10023,N_10038);
or U11783 (N_11783,N_9565,N_9173);
nand U11784 (N_11784,N_9173,N_10314);
and U11785 (N_11785,N_10290,N_10094);
nand U11786 (N_11786,N_9132,N_9757);
or U11787 (N_11787,N_10209,N_9275);
nor U11788 (N_11788,N_9000,N_9538);
and U11789 (N_11789,N_9218,N_9719);
or U11790 (N_11790,N_10013,N_9831);
nand U11791 (N_11791,N_9680,N_9403);
or U11792 (N_11792,N_9689,N_9985);
nand U11793 (N_11793,N_10289,N_9158);
and U11794 (N_11794,N_9373,N_10416);
xnor U11795 (N_11795,N_9917,N_10167);
xor U11796 (N_11796,N_9135,N_10338);
and U11797 (N_11797,N_9301,N_10085);
xor U11798 (N_11798,N_10144,N_9674);
nor U11799 (N_11799,N_10154,N_9057);
nand U11800 (N_11800,N_9881,N_9729);
xor U11801 (N_11801,N_9961,N_9065);
xor U11802 (N_11802,N_9770,N_9045);
or U11803 (N_11803,N_9632,N_9249);
nor U11804 (N_11804,N_9605,N_9558);
nand U11805 (N_11805,N_10036,N_9644);
nand U11806 (N_11806,N_10205,N_9696);
nor U11807 (N_11807,N_9864,N_9442);
or U11808 (N_11808,N_9276,N_10143);
and U11809 (N_11809,N_9417,N_9109);
or U11810 (N_11810,N_10323,N_9580);
nor U11811 (N_11811,N_9764,N_9729);
xor U11812 (N_11812,N_9731,N_9930);
nand U11813 (N_11813,N_9491,N_9178);
or U11814 (N_11814,N_9988,N_10317);
nand U11815 (N_11815,N_9823,N_9092);
nand U11816 (N_11816,N_10198,N_10308);
nor U11817 (N_11817,N_10006,N_9514);
or U11818 (N_11818,N_10154,N_9532);
xnor U11819 (N_11819,N_9354,N_9743);
or U11820 (N_11820,N_10233,N_10433);
and U11821 (N_11821,N_9450,N_9843);
xor U11822 (N_11822,N_10383,N_9943);
or U11823 (N_11823,N_9721,N_10107);
nor U11824 (N_11824,N_9106,N_9662);
xnor U11825 (N_11825,N_9383,N_9892);
nor U11826 (N_11826,N_9809,N_10182);
nor U11827 (N_11827,N_9845,N_10071);
xor U11828 (N_11828,N_10419,N_9218);
nor U11829 (N_11829,N_9858,N_9475);
and U11830 (N_11830,N_9435,N_9316);
nand U11831 (N_11831,N_9509,N_9698);
and U11832 (N_11832,N_9384,N_10182);
or U11833 (N_11833,N_9444,N_9809);
nand U11834 (N_11834,N_9984,N_9629);
nand U11835 (N_11835,N_9814,N_9051);
or U11836 (N_11836,N_9247,N_9203);
nor U11837 (N_11837,N_9886,N_10424);
nand U11838 (N_11838,N_9049,N_9781);
xor U11839 (N_11839,N_9714,N_9642);
and U11840 (N_11840,N_10124,N_9817);
xnor U11841 (N_11841,N_10151,N_9448);
nor U11842 (N_11842,N_9225,N_9075);
or U11843 (N_11843,N_9607,N_10330);
nand U11844 (N_11844,N_9500,N_9682);
nor U11845 (N_11845,N_9754,N_9307);
nor U11846 (N_11846,N_9866,N_9965);
nand U11847 (N_11847,N_10381,N_10418);
nand U11848 (N_11848,N_9222,N_9156);
nand U11849 (N_11849,N_9267,N_10242);
and U11850 (N_11850,N_10093,N_9761);
nand U11851 (N_11851,N_10199,N_9790);
and U11852 (N_11852,N_9436,N_9893);
xor U11853 (N_11853,N_9301,N_9764);
and U11854 (N_11854,N_10423,N_9421);
or U11855 (N_11855,N_9692,N_9015);
nand U11856 (N_11856,N_9653,N_10430);
nor U11857 (N_11857,N_9102,N_9906);
and U11858 (N_11858,N_10423,N_10389);
or U11859 (N_11859,N_10146,N_9225);
and U11860 (N_11860,N_9280,N_9145);
or U11861 (N_11861,N_9342,N_9409);
nand U11862 (N_11862,N_9557,N_9262);
nor U11863 (N_11863,N_9160,N_9316);
nor U11864 (N_11864,N_10375,N_9453);
nand U11865 (N_11865,N_9845,N_9955);
xor U11866 (N_11866,N_9563,N_10206);
or U11867 (N_11867,N_9909,N_10377);
nand U11868 (N_11868,N_9746,N_9394);
nor U11869 (N_11869,N_9588,N_9844);
and U11870 (N_11870,N_10267,N_9370);
nor U11871 (N_11871,N_9660,N_9291);
nor U11872 (N_11872,N_9247,N_10264);
nand U11873 (N_11873,N_10088,N_10142);
or U11874 (N_11874,N_9406,N_10369);
nor U11875 (N_11875,N_10484,N_10021);
or U11876 (N_11876,N_10402,N_10156);
nand U11877 (N_11877,N_9235,N_9134);
nand U11878 (N_11878,N_9568,N_9084);
and U11879 (N_11879,N_10406,N_9687);
and U11880 (N_11880,N_9412,N_9299);
and U11881 (N_11881,N_9124,N_9832);
xnor U11882 (N_11882,N_9645,N_9091);
nor U11883 (N_11883,N_9178,N_10293);
nor U11884 (N_11884,N_9444,N_10123);
or U11885 (N_11885,N_10081,N_9139);
nor U11886 (N_11886,N_10453,N_10126);
or U11887 (N_11887,N_9437,N_10113);
and U11888 (N_11888,N_9147,N_10357);
or U11889 (N_11889,N_9552,N_9918);
and U11890 (N_11890,N_9216,N_9864);
xnor U11891 (N_11891,N_9130,N_9804);
or U11892 (N_11892,N_9990,N_9311);
nor U11893 (N_11893,N_10057,N_9320);
nor U11894 (N_11894,N_10484,N_9731);
or U11895 (N_11895,N_9162,N_9806);
xnor U11896 (N_11896,N_10030,N_9381);
nand U11897 (N_11897,N_9742,N_9261);
nor U11898 (N_11898,N_9275,N_9935);
and U11899 (N_11899,N_9337,N_9119);
xnor U11900 (N_11900,N_10335,N_9612);
nor U11901 (N_11901,N_9594,N_9506);
or U11902 (N_11902,N_9294,N_9821);
or U11903 (N_11903,N_9341,N_9872);
or U11904 (N_11904,N_9441,N_9378);
or U11905 (N_11905,N_9989,N_10184);
nand U11906 (N_11906,N_9559,N_9745);
nand U11907 (N_11907,N_9394,N_9971);
and U11908 (N_11908,N_9987,N_9504);
and U11909 (N_11909,N_9288,N_10002);
and U11910 (N_11910,N_9868,N_9880);
nor U11911 (N_11911,N_10011,N_10103);
and U11912 (N_11912,N_9907,N_10061);
or U11913 (N_11913,N_9860,N_10001);
nand U11914 (N_11914,N_10128,N_9708);
nor U11915 (N_11915,N_9977,N_9577);
and U11916 (N_11916,N_9106,N_9740);
or U11917 (N_11917,N_10483,N_9360);
xnor U11918 (N_11918,N_9722,N_9986);
xor U11919 (N_11919,N_9414,N_10073);
nor U11920 (N_11920,N_9684,N_9325);
and U11921 (N_11921,N_10386,N_9517);
xnor U11922 (N_11922,N_9628,N_9793);
xor U11923 (N_11923,N_9271,N_9546);
nor U11924 (N_11924,N_9344,N_9648);
xor U11925 (N_11925,N_10459,N_9672);
xnor U11926 (N_11926,N_9205,N_9624);
or U11927 (N_11927,N_10491,N_9234);
or U11928 (N_11928,N_10118,N_10129);
or U11929 (N_11929,N_9554,N_9520);
nand U11930 (N_11930,N_10202,N_10372);
nor U11931 (N_11931,N_9812,N_9479);
nand U11932 (N_11932,N_10369,N_10015);
nor U11933 (N_11933,N_10102,N_10011);
nand U11934 (N_11934,N_10149,N_9604);
nor U11935 (N_11935,N_9256,N_9733);
nand U11936 (N_11936,N_9987,N_10314);
xnor U11937 (N_11937,N_10006,N_9885);
nor U11938 (N_11938,N_9693,N_10296);
nand U11939 (N_11939,N_9057,N_10092);
or U11940 (N_11940,N_9289,N_9156);
nor U11941 (N_11941,N_9632,N_9129);
nor U11942 (N_11942,N_10450,N_10197);
or U11943 (N_11943,N_9939,N_9113);
or U11944 (N_11944,N_9208,N_9765);
nand U11945 (N_11945,N_9841,N_9100);
xnor U11946 (N_11946,N_10304,N_9413);
xnor U11947 (N_11947,N_9323,N_10287);
xnor U11948 (N_11948,N_9408,N_9057);
xor U11949 (N_11949,N_9958,N_9112);
and U11950 (N_11950,N_9439,N_10365);
and U11951 (N_11951,N_10311,N_9472);
or U11952 (N_11952,N_10354,N_10017);
or U11953 (N_11953,N_9459,N_10281);
or U11954 (N_11954,N_9393,N_10051);
xnor U11955 (N_11955,N_9080,N_10179);
nand U11956 (N_11956,N_9018,N_9566);
nand U11957 (N_11957,N_9552,N_10310);
or U11958 (N_11958,N_9162,N_9654);
and U11959 (N_11959,N_10438,N_9228);
and U11960 (N_11960,N_9715,N_9266);
nand U11961 (N_11961,N_9504,N_9233);
and U11962 (N_11962,N_10138,N_10067);
xnor U11963 (N_11963,N_10159,N_9869);
xnor U11964 (N_11964,N_9570,N_9721);
xor U11965 (N_11965,N_9478,N_9975);
nor U11966 (N_11966,N_9541,N_9292);
nor U11967 (N_11967,N_10061,N_9533);
nand U11968 (N_11968,N_9261,N_9055);
or U11969 (N_11969,N_10130,N_10319);
or U11970 (N_11970,N_9892,N_9698);
and U11971 (N_11971,N_9402,N_9640);
xnor U11972 (N_11972,N_9706,N_9236);
nand U11973 (N_11973,N_9149,N_9193);
and U11974 (N_11974,N_10248,N_10477);
or U11975 (N_11975,N_9681,N_9552);
or U11976 (N_11976,N_9800,N_10349);
nand U11977 (N_11977,N_10320,N_9922);
and U11978 (N_11978,N_9403,N_9831);
or U11979 (N_11979,N_9247,N_10094);
nand U11980 (N_11980,N_9396,N_9194);
nor U11981 (N_11981,N_9755,N_9436);
xor U11982 (N_11982,N_9566,N_9822);
or U11983 (N_11983,N_9561,N_10279);
or U11984 (N_11984,N_10232,N_9218);
xnor U11985 (N_11985,N_10347,N_10012);
or U11986 (N_11986,N_9813,N_9733);
nand U11987 (N_11987,N_10238,N_9351);
and U11988 (N_11988,N_9535,N_10286);
or U11989 (N_11989,N_9071,N_9540);
and U11990 (N_11990,N_9670,N_10242);
nand U11991 (N_11991,N_9291,N_10044);
or U11992 (N_11992,N_10111,N_10353);
xnor U11993 (N_11993,N_9485,N_10013);
or U11994 (N_11994,N_9689,N_9323);
nor U11995 (N_11995,N_9057,N_9065);
or U11996 (N_11996,N_9888,N_10361);
nand U11997 (N_11997,N_9895,N_9482);
and U11998 (N_11998,N_10253,N_9768);
and U11999 (N_11999,N_9109,N_9865);
xor U12000 (N_12000,N_10607,N_11747);
nor U12001 (N_12001,N_11628,N_10946);
nand U12002 (N_12002,N_11231,N_11339);
nor U12003 (N_12003,N_11674,N_11417);
nand U12004 (N_12004,N_10529,N_11586);
and U12005 (N_12005,N_10907,N_11750);
and U12006 (N_12006,N_11185,N_11596);
or U12007 (N_12007,N_11435,N_11825);
and U12008 (N_12008,N_11313,N_10848);
or U12009 (N_12009,N_11388,N_11241);
nor U12010 (N_12010,N_10780,N_11732);
nor U12011 (N_12011,N_11605,N_11005);
or U12012 (N_12012,N_11360,N_11955);
or U12013 (N_12013,N_11852,N_11340);
xor U12014 (N_12014,N_10899,N_11936);
nand U12015 (N_12015,N_11515,N_11050);
or U12016 (N_12016,N_11723,N_10557);
or U12017 (N_12017,N_11544,N_11549);
or U12018 (N_12018,N_11531,N_10764);
xor U12019 (N_12019,N_11020,N_11572);
or U12020 (N_12020,N_11455,N_11080);
nand U12021 (N_12021,N_10827,N_11437);
nand U12022 (N_12022,N_10865,N_11902);
nand U12023 (N_12023,N_11416,N_11062);
nor U12024 (N_12024,N_10853,N_11726);
nor U12025 (N_12025,N_11295,N_11940);
nor U12026 (N_12026,N_11274,N_10575);
and U12027 (N_12027,N_11139,N_11903);
or U12028 (N_12028,N_11190,N_11907);
xor U12029 (N_12029,N_11662,N_10763);
and U12030 (N_12030,N_11436,N_11075);
nand U12031 (N_12031,N_11973,N_11057);
nor U12032 (N_12032,N_10699,N_10672);
xor U12033 (N_12033,N_10549,N_11843);
xor U12034 (N_12034,N_10733,N_11968);
xnor U12035 (N_12035,N_11823,N_11908);
nor U12036 (N_12036,N_10998,N_11087);
and U12037 (N_12037,N_10519,N_11117);
xor U12038 (N_12038,N_10734,N_11780);
nand U12039 (N_12039,N_11249,N_10837);
nor U12040 (N_12040,N_11119,N_11439);
and U12041 (N_12041,N_10874,N_10993);
or U12042 (N_12042,N_11028,N_11768);
nand U12043 (N_12043,N_10700,N_11795);
nand U12044 (N_12044,N_11332,N_11290);
xor U12045 (N_12045,N_11576,N_11895);
nor U12046 (N_12046,N_11552,N_11326);
or U12047 (N_12047,N_11582,N_11227);
or U12048 (N_12048,N_11483,N_10921);
xor U12049 (N_12049,N_10904,N_10801);
nor U12050 (N_12050,N_10924,N_11857);
and U12051 (N_12051,N_10635,N_10824);
nand U12052 (N_12052,N_10881,N_11868);
and U12053 (N_12053,N_11336,N_11865);
xnor U12054 (N_12054,N_11045,N_11320);
or U12055 (N_12055,N_11162,N_11129);
nor U12056 (N_12056,N_11869,N_11900);
and U12057 (N_12057,N_11137,N_10523);
nand U12058 (N_12058,N_11767,N_11248);
and U12059 (N_12059,N_10631,N_11055);
or U12060 (N_12060,N_10761,N_11929);
xnor U12061 (N_12061,N_11366,N_11074);
nor U12062 (N_12062,N_11545,N_11703);
xor U12063 (N_12063,N_11676,N_11820);
or U12064 (N_12064,N_11851,N_10928);
nand U12065 (N_12065,N_11670,N_11383);
or U12066 (N_12066,N_11950,N_11121);
nand U12067 (N_12067,N_11397,N_10933);
nor U12068 (N_12068,N_11251,N_11101);
nor U12069 (N_12069,N_11229,N_11407);
and U12070 (N_12070,N_11991,N_10569);
nor U12071 (N_12071,N_11447,N_11764);
xor U12072 (N_12072,N_10554,N_11655);
nand U12073 (N_12073,N_10915,N_11223);
xor U12074 (N_12074,N_11584,N_11150);
or U12075 (N_12075,N_11245,N_11860);
nor U12076 (N_12076,N_10883,N_10606);
nor U12077 (N_12077,N_11424,N_11076);
nand U12078 (N_12078,N_11202,N_11499);
xnor U12079 (N_12079,N_10997,N_11328);
nor U12080 (N_12080,N_10566,N_10867);
or U12081 (N_12081,N_11078,N_11421);
xnor U12082 (N_12082,N_11469,N_11719);
and U12083 (N_12083,N_11053,N_10769);
nor U12084 (N_12084,N_10593,N_10846);
nor U12085 (N_12085,N_11694,N_11266);
nor U12086 (N_12086,N_11634,N_11384);
nor U12087 (N_12087,N_11198,N_11714);
and U12088 (N_12088,N_11598,N_10659);
nor U12089 (N_12089,N_10679,N_11555);
or U12090 (N_12090,N_11304,N_11432);
and U12091 (N_12091,N_11650,N_11707);
or U12092 (N_12092,N_11587,N_11562);
nand U12093 (N_12093,N_10614,N_11255);
nand U12094 (N_12094,N_11633,N_11947);
xnor U12095 (N_12095,N_11931,N_10712);
xor U12096 (N_12096,N_11052,N_10947);
nand U12097 (N_12097,N_11367,N_11638);
nor U12098 (N_12098,N_10917,N_10859);
or U12099 (N_12099,N_11413,N_11524);
nor U12100 (N_12100,N_10615,N_10884);
nand U12101 (N_12101,N_11839,N_11099);
and U12102 (N_12102,N_11058,N_10738);
and U12103 (N_12103,N_11807,N_10953);
nor U12104 (N_12104,N_11254,N_10806);
or U12105 (N_12105,N_10804,N_11639);
or U12106 (N_12106,N_11359,N_10788);
and U12107 (N_12107,N_10526,N_11663);
xor U12108 (N_12108,N_10987,N_11517);
xnor U12109 (N_12109,N_10822,N_10646);
nand U12110 (N_12110,N_10617,N_10849);
xor U12111 (N_12111,N_11205,N_11479);
xnor U12112 (N_12112,N_10879,N_11035);
xor U12113 (N_12113,N_11637,N_11946);
nand U12114 (N_12114,N_11140,N_11874);
nand U12115 (N_12115,N_10852,N_11398);
and U12116 (N_12116,N_11525,N_11866);
nand U12117 (N_12117,N_11490,N_10532);
and U12118 (N_12118,N_10990,N_10901);
nor U12119 (N_12119,N_10638,N_11235);
nand U12120 (N_12120,N_11652,N_10817);
and U12121 (N_12121,N_10926,N_11267);
nand U12122 (N_12122,N_10748,N_10759);
nor U12123 (N_12123,N_11518,N_11678);
nand U12124 (N_12124,N_10825,N_10520);
and U12125 (N_12125,N_10751,N_10686);
or U12126 (N_12126,N_10728,N_11867);
nand U12127 (N_12127,N_10685,N_10775);
xnor U12128 (N_12128,N_10755,N_11506);
nor U12129 (N_12129,N_10839,N_10571);
or U12130 (N_12130,N_11463,N_11174);
nor U12131 (N_12131,N_11211,N_10911);
nand U12132 (N_12132,N_11813,N_11399);
nand U12133 (N_12133,N_11563,N_11878);
nand U12134 (N_12134,N_10739,N_11575);
nor U12135 (N_12135,N_10609,N_10522);
and U12136 (N_12136,N_11096,N_11011);
nor U12137 (N_12137,N_10931,N_10586);
xor U12138 (N_12138,N_11998,N_11762);
or U12139 (N_12139,N_11256,N_11146);
and U12140 (N_12140,N_11748,N_10649);
nor U12141 (N_12141,N_10560,N_10666);
nand U12142 (N_12142,N_11606,N_11411);
nand U12143 (N_12143,N_11550,N_11318);
and U12144 (N_12144,N_11126,N_11079);
and U12145 (N_12145,N_11305,N_11220);
nor U12146 (N_12146,N_11039,N_11574);
xnor U12147 (N_12147,N_11932,N_10534);
or U12148 (N_12148,N_11926,N_11412);
and U12149 (N_12149,N_10925,N_11888);
and U12150 (N_12150,N_11391,N_11100);
xor U12151 (N_12151,N_11071,N_11175);
xnor U12152 (N_12152,N_11543,N_11418);
or U12153 (N_12153,N_10886,N_11170);
xnor U12154 (N_12154,N_11191,N_11018);
nand U12155 (N_12155,N_10979,N_10627);
nand U12156 (N_12156,N_11830,N_11493);
and U12157 (N_12157,N_11380,N_10891);
xor U12158 (N_12158,N_11920,N_11921);
or U12159 (N_12159,N_11597,N_10644);
and U12160 (N_12160,N_10779,N_11130);
or U12161 (N_12161,N_11457,N_10744);
nor U12162 (N_12162,N_10982,N_11840);
or U12163 (N_12163,N_11118,N_11183);
and U12164 (N_12164,N_11265,N_11648);
and U12165 (N_12165,N_11937,N_10511);
nand U12166 (N_12166,N_11884,N_11063);
and U12167 (N_12167,N_11453,N_11094);
or U12168 (N_12168,N_11386,N_11646);
and U12169 (N_12169,N_10720,N_11466);
or U12170 (N_12170,N_10625,N_10999);
and U12171 (N_12171,N_11164,N_10658);
or U12172 (N_12172,N_10992,N_11793);
nor U12173 (N_12173,N_11573,N_11643);
or U12174 (N_12174,N_10823,N_11627);
xor U12175 (N_12175,N_11798,N_11307);
xor U12176 (N_12176,N_11914,N_11487);
nand U12177 (N_12177,N_11565,N_11504);
xor U12178 (N_12178,N_11855,N_10515);
nor U12179 (N_12179,N_10785,N_11385);
or U12180 (N_12180,N_10944,N_11116);
xor U12181 (N_12181,N_10912,N_11833);
xnor U12182 (N_12182,N_11355,N_11713);
nor U12183 (N_12183,N_11426,N_11217);
or U12184 (N_12184,N_11242,N_10880);
and U12185 (N_12185,N_11854,N_11072);
or U12186 (N_12186,N_11401,N_10969);
nor U12187 (N_12187,N_11478,N_11836);
nand U12188 (N_12188,N_11083,N_11753);
or U12189 (N_12189,N_11610,N_10657);
and U12190 (N_12190,N_11514,N_11738);
and U12191 (N_12191,N_11147,N_11017);
nor U12192 (N_12192,N_10678,N_10930);
xor U12193 (N_12193,N_11029,N_11067);
xor U12194 (N_12194,N_10637,N_11702);
xnor U12195 (N_12195,N_11476,N_11530);
or U12196 (N_12196,N_10608,N_11448);
or U12197 (N_12197,N_10758,N_11454);
nor U12198 (N_12198,N_11972,N_10596);
xor U12199 (N_12199,N_10564,N_10861);
nor U12200 (N_12200,N_11458,N_11015);
or U12201 (N_12201,N_11601,N_10828);
and U12202 (N_12202,N_11828,N_10976);
nand U12203 (N_12203,N_11644,N_10746);
xor U12204 (N_12204,N_11700,N_11561);
nand U12205 (N_12205,N_11805,N_11960);
nand U12206 (N_12206,N_10762,N_10754);
nand U12207 (N_12207,N_11526,N_11272);
nand U12208 (N_12208,N_11776,N_11289);
and U12209 (N_12209,N_10684,N_11294);
nand U12210 (N_12210,N_11176,N_10794);
nand U12211 (N_12211,N_10991,N_11814);
nor U12212 (N_12212,N_11312,N_11647);
xnor U12213 (N_12213,N_11023,N_11724);
or U12214 (N_12214,N_11465,N_11887);
or U12215 (N_12215,N_11957,N_10690);
nor U12216 (N_12216,N_11329,N_11635);
and U12217 (N_12217,N_11533,N_11761);
nand U12218 (N_12218,N_10851,N_11405);
nor U12219 (N_12219,N_11409,N_10932);
and U12220 (N_12220,N_11989,N_11037);
nor U12221 (N_12221,N_11675,N_10835);
nor U12222 (N_12222,N_10581,N_11066);
xnor U12223 (N_12223,N_11396,N_10524);
and U12224 (N_12224,N_11686,N_10948);
and U12225 (N_12225,N_11194,N_11711);
nand U12226 (N_12226,N_10701,N_10521);
or U12227 (N_12227,N_10961,N_10622);
nand U12228 (N_12228,N_10562,N_11788);
xnor U12229 (N_12229,N_11141,N_10974);
and U12230 (N_12230,N_11240,N_10818);
nand U12231 (N_12231,N_11997,N_11941);
and U12232 (N_12232,N_10798,N_11781);
nor U12233 (N_12233,N_11297,N_11065);
or U12234 (N_12234,N_11155,N_11302);
and U12235 (N_12235,N_11014,N_11911);
or U12236 (N_12236,N_11456,N_11611);
nor U12237 (N_12237,N_11161,N_11371);
xnor U12238 (N_12238,N_11779,N_11898);
xnor U12239 (N_12239,N_11310,N_10945);
nor U12240 (N_12240,N_11275,N_11348);
and U12241 (N_12241,N_11200,N_10927);
nand U12242 (N_12242,N_11209,N_10641);
xor U12243 (N_12243,N_11850,N_11342);
or U12244 (N_12244,N_11812,N_11691);
nor U12245 (N_12245,N_11353,N_10730);
nand U12246 (N_12246,N_11571,N_10873);
xnor U12247 (N_12247,N_11236,N_10781);
xnor U12248 (N_12248,N_11153,N_11016);
and U12249 (N_12249,N_11132,N_11891);
nor U12250 (N_12250,N_11151,N_11566);
xnor U12251 (N_12251,N_11376,N_11001);
and U12252 (N_12252,N_11108,N_10651);
xnor U12253 (N_12253,N_10753,N_11803);
nand U12254 (N_12254,N_11494,N_10624);
xor U12255 (N_12255,N_11237,N_10682);
nand U12256 (N_12256,N_10791,N_11987);
nand U12257 (N_12257,N_11886,N_10501);
xor U12258 (N_12258,N_11002,N_10725);
nand U12259 (N_12259,N_11541,N_11327);
and U12260 (N_12260,N_11690,N_11996);
or U12261 (N_12261,N_10630,N_11934);
or U12262 (N_12262,N_10680,N_11356);
xor U12263 (N_12263,N_10671,N_11640);
nand U12264 (N_12264,N_11428,N_11171);
nor U12265 (N_12265,N_10950,N_11293);
or U12266 (N_12266,N_11979,N_11809);
or U12267 (N_12267,N_10616,N_10592);
or U12268 (N_12268,N_11540,N_10715);
and U12269 (N_12269,N_11993,N_11128);
nor U12270 (N_12270,N_11963,N_11591);
nand U12271 (N_12271,N_11508,N_10600);
xor U12272 (N_12272,N_11300,N_10995);
and U12273 (N_12273,N_11532,N_10536);
or U12274 (N_12274,N_10902,N_11551);
xnor U12275 (N_12275,N_11984,N_11077);
nor U12276 (N_12276,N_11789,N_11093);
nor U12277 (N_12277,N_11896,N_10653);
and U12278 (N_12278,N_11306,N_11815);
nand U12279 (N_12279,N_10517,N_11943);
nor U12280 (N_12280,N_10623,N_11430);
nand U12281 (N_12281,N_10978,N_11226);
and U12282 (N_12282,N_10796,N_11145);
nor U12283 (N_12283,N_11292,N_11033);
xnor U12284 (N_12284,N_11983,N_10655);
xor U12285 (N_12285,N_10578,N_10507);
and U12286 (N_12286,N_11782,N_11459);
nand U12287 (N_12287,N_11743,N_11621);
or U12288 (N_12288,N_11158,N_11600);
or U12289 (N_12289,N_10660,N_11910);
or U12290 (N_12290,N_10537,N_10602);
nor U12291 (N_12291,N_10939,N_11986);
nand U12292 (N_12292,N_11013,N_11107);
and U12293 (N_12293,N_11285,N_10832);
nor U12294 (N_12294,N_10756,N_11480);
nand U12295 (N_12295,N_11475,N_10640);
or U12296 (N_12296,N_11154,N_11064);
nor U12297 (N_12297,N_10777,N_10726);
or U12298 (N_12298,N_11933,N_11239);
or U12299 (N_12299,N_10790,N_11070);
and U12300 (N_12300,N_10888,N_10810);
nand U12301 (N_12301,N_11889,N_11389);
xor U12302 (N_12302,N_11025,N_10548);
or U12303 (N_12303,N_11163,N_11470);
xnor U12304 (N_12304,N_11197,N_10960);
nand U12305 (N_12305,N_10724,N_11927);
nor U12306 (N_12306,N_11420,N_11402);
xnor U12307 (N_12307,N_10567,N_11935);
nand U12308 (N_12308,N_10705,N_10923);
nor U12309 (N_12309,N_11831,N_10603);
or U12310 (N_12310,N_11821,N_11822);
or U12311 (N_12311,N_10513,N_10866);
nand U12312 (N_12312,N_10745,N_11010);
nand U12313 (N_12313,N_10563,N_11721);
nor U12314 (N_12314,N_10709,N_11156);
or U12315 (N_12315,N_10989,N_10750);
nand U12316 (N_12316,N_11451,N_11885);
and U12317 (N_12317,N_11400,N_11007);
nand U12318 (N_12318,N_11992,N_11192);
xor U12319 (N_12319,N_11953,N_10661);
xor U12320 (N_12320,N_11507,N_10510);
or U12321 (N_12321,N_11649,N_10914);
xor U12322 (N_12322,N_11207,N_11682);
and U12323 (N_12323,N_11134,N_11665);
or U12324 (N_12324,N_10772,N_11994);
xor U12325 (N_12325,N_11681,N_10949);
nand U12326 (N_12326,N_11378,N_10882);
xnor U12327 (N_12327,N_11219,N_11602);
nand U12328 (N_12328,N_11036,N_11995);
nand U12329 (N_12329,N_10918,N_11826);
nand U12330 (N_12330,N_11500,N_10943);
and U12331 (N_12331,N_11195,N_11725);
and U12332 (N_12332,N_11485,N_11556);
nor U12333 (N_12333,N_10757,N_11364);
xor U12334 (N_12334,N_10703,N_11568);
nor U12335 (N_12335,N_10539,N_11434);
and U12336 (N_12336,N_10833,N_11497);
xor U12337 (N_12337,N_10552,N_11804);
or U12338 (N_12338,N_10533,N_11614);
or U12339 (N_12339,N_10906,N_11031);
and U12340 (N_12340,N_11212,N_10765);
nor U12341 (N_12341,N_11751,N_10729);
and U12342 (N_12342,N_11509,N_10820);
nand U12343 (N_12343,N_11189,N_11250);
nor U12344 (N_12344,N_11810,N_10692);
nand U12345 (N_12345,N_11742,N_11969);
nor U12346 (N_12346,N_11443,N_10735);
nor U12347 (N_12347,N_11184,N_10908);
or U12348 (N_12348,N_11387,N_11752);
nor U12349 (N_12349,N_10951,N_11999);
xnor U12350 (N_12350,N_10895,N_11109);
nor U12351 (N_12351,N_11299,N_11612);
nand U12352 (N_12352,N_10722,N_11787);
nand U12353 (N_12353,N_11785,N_10583);
nand U12354 (N_12354,N_11930,N_10530);
xor U12355 (N_12355,N_11734,N_10589);
xor U12356 (N_12356,N_11577,N_11971);
and U12357 (N_12357,N_11948,N_10809);
and U12358 (N_12358,N_11693,N_11321);
xor U12359 (N_12359,N_11680,N_11547);
or U12360 (N_12360,N_10694,N_11722);
and U12361 (N_12361,N_11381,N_11361);
nor U12362 (N_12362,N_10704,N_11912);
xnor U12363 (N_12363,N_10965,N_11102);
nor U12364 (N_12364,N_11203,N_11232);
nand U12365 (N_12365,N_10527,N_10736);
nand U12366 (N_12366,N_11131,N_11474);
and U12367 (N_12367,N_11089,N_11863);
and U12368 (N_12368,N_11004,N_11570);
xor U12369 (N_12369,N_11923,N_11090);
nand U12370 (N_12370,N_10547,N_11350);
and U12371 (N_12371,N_11201,N_11791);
nand U12372 (N_12372,N_11442,N_11672);
and U12373 (N_12373,N_11988,N_10508);
and U12374 (N_12374,N_11777,N_11542);
or U12375 (N_12375,N_11775,N_11169);
xnor U12376 (N_12376,N_11578,N_11641);
nand U12377 (N_12377,N_11808,N_10541);
nand U12378 (N_12378,N_11778,N_11939);
or U12379 (N_12379,N_11486,N_11419);
and U12380 (N_12380,N_11666,N_10598);
xor U12381 (N_12381,N_10803,N_11127);
nand U12382 (N_12382,N_11754,N_11848);
nand U12383 (N_12383,N_11861,N_10558);
nand U12384 (N_12384,N_10693,N_11111);
and U12385 (N_12385,N_10771,N_11842);
nor U12386 (N_12386,N_11425,N_11363);
nor U12387 (N_12387,N_11879,N_11873);
xor U12388 (N_12388,N_10985,N_10860);
nand U12389 (N_12389,N_11247,N_10813);
nand U12390 (N_12390,N_11583,N_11214);
or U12391 (N_12391,N_11728,N_11303);
nand U12392 (N_12392,N_11838,N_11182);
nand U12393 (N_12393,N_11379,N_11604);
nand U12394 (N_12394,N_10887,N_10941);
nand U12395 (N_12395,N_10662,N_11603);
nand U12396 (N_12396,N_11133,N_10862);
and U12397 (N_12397,N_11962,N_11097);
or U12398 (N_12398,N_10977,N_10707);
xor U12399 (N_12399,N_10514,N_11315);
and U12400 (N_12400,N_10877,N_10996);
nor U12401 (N_12401,N_11745,N_11216);
and U12402 (N_12402,N_11658,N_10505);
and U12403 (N_12403,N_11343,N_10585);
nor U12404 (N_12404,N_11122,N_11990);
and U12405 (N_12405,N_11187,N_11951);
xor U12406 (N_12406,N_10831,N_10611);
nor U12407 (N_12407,N_10870,N_10970);
nor U12408 (N_12408,N_11165,N_10845);
nor U12409 (N_12409,N_11668,N_11222);
nor U12410 (N_12410,N_11441,N_11283);
nor U12411 (N_12411,N_11279,N_10621);
nand U12412 (N_12412,N_11392,N_10811);
or U12413 (N_12413,N_11982,N_11354);
or U12414 (N_12414,N_10760,N_11268);
or U12415 (N_12415,N_11701,N_10500);
or U12416 (N_12416,N_11536,N_10634);
nor U12417 (N_12417,N_11177,N_11797);
nand U12418 (N_12418,N_10595,N_10687);
and U12419 (N_12419,N_11349,N_10767);
nor U12420 (N_12420,N_11280,N_11692);
nand U12421 (N_12421,N_11160,N_11844);
or U12422 (N_12422,N_10857,N_10584);
xor U12423 (N_12423,N_11624,N_10983);
xnor U12424 (N_12424,N_11204,N_10620);
nor U12425 (N_12425,N_10916,N_11949);
nor U12426 (N_12426,N_11763,N_11422);
nand U12427 (N_12427,N_10905,N_10934);
nand U12428 (N_12428,N_11046,N_11904);
xnor U12429 (N_12429,N_11717,N_11309);
nor U12430 (N_12430,N_11178,N_11414);
nor U12431 (N_12431,N_10876,N_11925);
xnor U12432 (N_12432,N_10697,N_11964);
nor U12433 (N_12433,N_10714,N_10639);
xor U12434 (N_12434,N_11073,N_11370);
nor U12435 (N_12435,N_11038,N_10587);
or U12436 (N_12436,N_11006,N_11186);
xor U12437 (N_12437,N_11375,N_11429);
nand U12438 (N_12438,N_11718,N_10669);
nand U12439 (N_12439,N_11460,N_11684);
nand U12440 (N_12440,N_11330,N_10668);
xnor U12441 (N_12441,N_11569,N_11959);
nor U12442 (N_12442,N_11757,N_11837);
xnor U12443 (N_12443,N_11166,N_10674);
nand U12444 (N_12444,N_11944,N_11756);
xnor U12445 (N_12445,N_11985,N_10717);
and U12446 (N_12446,N_11270,N_11149);
nor U12447 (N_12447,N_10786,N_11511);
and U12448 (N_12448,N_11317,N_11765);
or U12449 (N_12449,N_11730,N_10975);
or U12450 (N_12450,N_11609,N_11243);
nor U12451 (N_12451,N_11567,N_11629);
nand U12452 (N_12452,N_11799,N_10792);
nor U12453 (N_12453,N_11449,N_10604);
xnor U12454 (N_12454,N_11471,N_11528);
nand U12455 (N_12455,N_11081,N_11225);
xor U12456 (N_12456,N_10793,N_11739);
xnor U12457 (N_12457,N_11345,N_11346);
or U12458 (N_12458,N_11301,N_11467);
xnor U12459 (N_12459,N_11636,N_10894);
or U12460 (N_12460,N_11660,N_10841);
xor U12461 (N_12461,N_11196,N_10783);
and U12462 (N_12462,N_11916,N_11382);
and U12463 (N_12463,N_10663,N_11917);
and U12464 (N_12464,N_10675,N_11771);
nand U12465 (N_12465,N_11019,N_10922);
or U12466 (N_12466,N_11864,N_10885);
nor U12467 (N_12467,N_10968,N_11922);
nor U12468 (N_12468,N_10706,N_10789);
nand U12469 (N_12469,N_11088,N_11496);
or U12470 (N_12470,N_10599,N_11769);
xor U12471 (N_12471,N_11905,N_10544);
nor U12472 (N_12472,N_10872,N_11731);
xnor U12473 (N_12473,N_11774,N_11143);
nand U12474 (N_12474,N_11564,N_11811);
xnor U12475 (N_12475,N_11915,N_10506);
xnor U12476 (N_12476,N_11816,N_11026);
and U12477 (N_12477,N_10807,N_11406);
xor U12478 (N_12478,N_10731,N_11427);
or U12479 (N_12479,N_11687,N_11252);
or U12480 (N_12480,N_11817,N_11589);
nand U12481 (N_12481,N_11003,N_11618);
nand U12482 (N_12482,N_11372,N_11462);
and U12483 (N_12483,N_10821,N_11218);
and U12484 (N_12484,N_11112,N_10956);
nand U12485 (N_12485,N_10816,N_11086);
xnor U12486 (N_12486,N_10542,N_10708);
or U12487 (N_12487,N_11193,N_11115);
and U12488 (N_12488,N_11706,N_10568);
or U12489 (N_12489,N_11630,N_11709);
xor U12490 (N_12490,N_11792,N_10619);
nor U12491 (N_12491,N_11325,N_10875);
xor U12492 (N_12492,N_11595,N_11735);
nand U12493 (N_12493,N_11452,N_11032);
nor U12494 (N_12494,N_11488,N_11492);
or U12495 (N_12495,N_10980,N_10696);
nor U12496 (N_12496,N_10525,N_11790);
xnor U12497 (N_12497,N_10778,N_11311);
nand U12498 (N_12498,N_11651,N_10898);
and U12499 (N_12499,N_11834,N_10555);
xor U12500 (N_12500,N_11827,N_10850);
and U12501 (N_12501,N_11978,N_10509);
or U12502 (N_12502,N_11059,N_10721);
nand U12503 (N_12503,N_10826,N_11308);
nand U12504 (N_12504,N_10727,N_10543);
xnor U12505 (N_12505,N_10652,N_10732);
or U12506 (N_12506,N_11148,N_11410);
xnor U12507 (N_12507,N_11590,N_11558);
or U12508 (N_12508,N_11892,N_10890);
xnor U12509 (N_12509,N_11450,N_10768);
nand U12510 (N_12510,N_10590,N_11259);
xor U12511 (N_12511,N_11374,N_11581);
nor U12512 (N_12512,N_11736,N_10551);
nor U12513 (N_12513,N_10787,N_10643);
nor U12514 (N_12514,N_11468,N_11626);
nand U12515 (N_12515,N_11104,N_10795);
nor U12516 (N_12516,N_11503,N_11796);
xnor U12517 (N_12517,N_11390,N_10574);
nand U12518 (N_12518,N_11806,N_10957);
and U12519 (N_12519,N_10576,N_11890);
nand U12520 (N_12520,N_10829,N_11210);
and U12521 (N_12521,N_11699,N_11871);
or U12522 (N_12522,N_10910,N_10691);
or U12523 (N_12523,N_11337,N_10695);
xor U12524 (N_12524,N_11049,N_11673);
and U12525 (N_12525,N_10830,N_10972);
nor U12526 (N_12526,N_11472,N_10920);
nand U12527 (N_12527,N_11091,N_11846);
xor U12528 (N_12528,N_11051,N_11705);
or U12529 (N_12529,N_11829,N_11755);
xor U12530 (N_12530,N_10940,N_11491);
nand U12531 (N_12531,N_10665,N_11897);
and U12532 (N_12532,N_11619,N_10858);
or U12533 (N_12533,N_11246,N_11446);
xnor U12534 (N_12534,N_11188,N_10952);
xor U12535 (N_12535,N_11585,N_10909);
or U12536 (N_12536,N_11977,N_11473);
or U12537 (N_12537,N_10868,N_10504);
nand U12538 (N_12538,N_10676,N_11284);
or U12539 (N_12539,N_10591,N_10994);
or U12540 (N_12540,N_11882,N_11976);
and U12541 (N_12541,N_10889,N_11881);
or U12542 (N_12542,N_11872,N_11261);
and U12543 (N_12543,N_11281,N_10565);
nand U12544 (N_12544,N_10844,N_11082);
xnor U12545 (N_12545,N_10766,N_11909);
nand U12546 (N_12546,N_11440,N_11928);
nand U12547 (N_12547,N_11659,N_11331);
and U12548 (N_12548,N_11616,N_10935);
nand U12549 (N_12549,N_11234,N_11230);
or U12550 (N_12550,N_11818,N_10834);
and U12551 (N_12551,N_11906,N_10561);
nand U12552 (N_12552,N_11720,N_11362);
nor U12553 (N_12553,N_11710,N_11546);
nor U12554 (N_12554,N_11858,N_11669);
nor U12555 (N_12555,N_10962,N_11352);
nor U12556 (N_12556,N_10774,N_10688);
nor U12557 (N_12557,N_11027,N_11919);
xnor U12558 (N_12558,N_11257,N_10752);
nand U12559 (N_12559,N_11445,N_11124);
or U12560 (N_12560,N_11980,N_11945);
nand U12561 (N_12561,N_11548,N_11138);
xor U12562 (N_12562,N_10737,N_11291);
xor U12563 (N_12563,N_11593,N_11512);
nor U12564 (N_12564,N_10698,N_11438);
xor U12565 (N_12565,N_11654,N_11880);
nand U12566 (N_12566,N_11802,N_10656);
nor U12567 (N_12567,N_10605,N_11704);
nand U12568 (N_12568,N_11484,N_11685);
nand U12569 (N_12569,N_10986,N_11110);
or U12570 (N_12570,N_10538,N_10838);
xor U12571 (N_12571,N_10799,N_11369);
xor U12572 (N_12572,N_11883,N_11258);
and U12573 (N_12573,N_11009,N_10776);
or U12574 (N_12574,N_10749,N_11824);
xnor U12575 (N_12575,N_11608,N_11553);
nor U12576 (N_12576,N_11733,N_11617);
xnor U12577 (N_12577,N_11084,N_11277);
and U12578 (N_12578,N_11727,N_10546);
nor U12579 (N_12579,N_11206,N_11952);
xnor U12580 (N_12580,N_10647,N_11224);
nor U12581 (N_12581,N_11853,N_11180);
or U12582 (N_12582,N_11415,N_10723);
nor U12583 (N_12583,N_10664,N_11334);
nand U12584 (N_12584,N_11683,N_10800);
or U12585 (N_12585,N_11238,N_11773);
or U12586 (N_12586,N_10570,N_11688);
or U12587 (N_12587,N_11594,N_11632);
and U12588 (N_12588,N_10988,N_11368);
xnor U12589 (N_12589,N_11276,N_11894);
nand U12590 (N_12590,N_11631,N_11938);
nor U12591 (N_12591,N_11539,N_11966);
or U12592 (N_12592,N_11365,N_11282);
nor U12593 (N_12593,N_10670,N_11461);
or U12594 (N_12594,N_10955,N_11695);
or U12595 (N_12595,N_11136,N_10959);
and U12596 (N_12596,N_10629,N_10577);
nor U12597 (N_12597,N_11758,N_11870);
or U12598 (N_12598,N_11579,N_11625);
nand U12599 (N_12599,N_11319,N_10681);
or U12600 (N_12600,N_10582,N_11677);
nand U12601 (N_12601,N_10812,N_10601);
nand U12602 (N_12602,N_10503,N_11744);
and U12603 (N_12603,N_11377,N_11269);
nor U12604 (N_12604,N_10903,N_11120);
or U12605 (N_12605,N_11847,N_11296);
xnor U12606 (N_12606,N_11698,N_10878);
and U12607 (N_12607,N_11008,N_11314);
and U12608 (N_12608,N_11288,N_10840);
nand U12609 (N_12609,N_11729,N_10718);
or U12610 (N_12610,N_11061,N_11974);
or U12611 (N_12611,N_11835,N_11716);
nor U12612 (N_12612,N_11298,N_10645);
and U12613 (N_12613,N_11954,N_11689);
nand U12614 (N_12614,N_10540,N_11607);
or U12615 (N_12615,N_11521,N_11273);
or U12616 (N_12616,N_10632,N_11642);
nor U12617 (N_12617,N_10642,N_10747);
or U12618 (N_12618,N_11351,N_10936);
or U12619 (N_12619,N_10966,N_10773);
xor U12620 (N_12620,N_11233,N_11105);
nor U12621 (N_12621,N_10559,N_11263);
and U12622 (N_12622,N_11021,N_11482);
nand U12623 (N_12623,N_11505,N_11519);
nand U12624 (N_12624,N_11357,N_10929);
nor U12625 (N_12625,N_11286,N_11172);
nand U12626 (N_12626,N_11522,N_10814);
nor U12627 (N_12627,N_11030,N_11667);
or U12628 (N_12628,N_10597,N_10636);
nor U12629 (N_12629,N_11877,N_11253);
and U12630 (N_12630,N_11221,N_11322);
nand U12631 (N_12631,N_11664,N_10856);
and U12632 (N_12632,N_11875,N_11024);
xor U12633 (N_12633,N_11344,N_11144);
or U12634 (N_12634,N_10667,N_11958);
and U12635 (N_12635,N_10770,N_10618);
nor U12636 (N_12636,N_10843,N_10854);
xor U12637 (N_12637,N_11069,N_10984);
or U12638 (N_12638,N_11358,N_10710);
and U12639 (N_12639,N_10797,N_10892);
or U12640 (N_12640,N_11431,N_11179);
or U12641 (N_12641,N_11554,N_11040);
and U12642 (N_12642,N_11845,N_11749);
nand U12643 (N_12643,N_11098,N_10550);
or U12644 (N_12644,N_11048,N_11740);
or U12645 (N_12645,N_11901,N_11022);
nor U12646 (N_12646,N_10689,N_11042);
xor U12647 (N_12647,N_10784,N_10743);
and U12648 (N_12648,N_11712,N_11786);
nand U12649 (N_12649,N_10528,N_11622);
xor U12650 (N_12650,N_11056,N_11746);
xor U12651 (N_12651,N_11085,N_10633);
or U12652 (N_12652,N_10863,N_11856);
nor U12653 (N_12653,N_10553,N_11168);
nor U12654 (N_12654,N_10819,N_11501);
or U12655 (N_12655,N_11696,N_11395);
nand U12656 (N_12656,N_10855,N_11152);
or U12657 (N_12657,N_10626,N_11034);
and U12658 (N_12658,N_11333,N_11956);
or U12659 (N_12659,N_11656,N_10971);
nor U12660 (N_12660,N_11516,N_11862);
xor U12661 (N_12661,N_11819,N_10967);
and U12662 (N_12662,N_11043,N_10805);
xnor U12663 (N_12663,N_11341,N_11615);
xnor U12664 (N_12664,N_10871,N_11167);
nor U12665 (N_12665,N_11125,N_11679);
nor U12666 (N_12666,N_10802,N_10628);
nand U12667 (N_12667,N_11433,N_10580);
xor U12668 (N_12668,N_11783,N_11535);
nor U12669 (N_12669,N_11913,N_10613);
and U12670 (N_12670,N_11278,N_10815);
nand U12671 (N_12671,N_11520,N_11671);
or U12672 (N_12672,N_10650,N_11213);
and U12673 (N_12673,N_11068,N_11975);
or U12674 (N_12674,N_11114,N_10893);
nand U12675 (N_12675,N_11095,N_10896);
nor U12676 (N_12676,N_10897,N_10502);
or U12677 (N_12677,N_11899,N_11538);
xor U12678 (N_12678,N_10677,N_11741);
and U12679 (N_12679,N_11316,N_10864);
nand U12680 (N_12680,N_10973,N_11159);
nor U12681 (N_12681,N_11092,N_11961);
and U12682 (N_12682,N_10648,N_11408);
or U12683 (N_12683,N_11697,N_11181);
xnor U12684 (N_12684,N_11645,N_11106);
nand U12685 (N_12685,N_10842,N_10958);
nor U12686 (N_12686,N_10919,N_10808);
nand U12687 (N_12687,N_10573,N_11859);
and U12688 (N_12688,N_11477,N_11444);
and U12689 (N_12689,N_11849,N_10512);
xnor U12690 (N_12690,N_10711,N_11794);
nor U12691 (N_12691,N_11715,N_10847);
nand U12692 (N_12692,N_10963,N_10719);
or U12693 (N_12693,N_10942,N_11580);
and U12694 (N_12694,N_11784,N_11404);
nor U12695 (N_12695,N_11557,N_11534);
and U12696 (N_12696,N_10900,N_11592);
nor U12697 (N_12697,N_10610,N_11766);
or U12698 (N_12698,N_11832,N_11489);
or U12699 (N_12699,N_11942,N_11394);
or U12700 (N_12700,N_11228,N_11708);
xor U12701 (N_12701,N_11103,N_11041);
or U12702 (N_12702,N_11620,N_11737);
xor U12703 (N_12703,N_11523,N_11653);
and U12704 (N_12704,N_10869,N_11924);
xor U12705 (N_12705,N_11481,N_10612);
nor U12706 (N_12706,N_11772,N_11970);
or U12707 (N_12707,N_11760,N_11324);
and U12708 (N_12708,N_10518,N_11613);
xnor U12709 (N_12709,N_11770,N_11323);
and U12710 (N_12710,N_10702,N_11559);
nor U12711 (N_12711,N_11199,N_11403);
and U12712 (N_12712,N_11510,N_11335);
or U12713 (N_12713,N_10937,N_11588);
and U12714 (N_12714,N_11157,N_11893);
xnor U12715 (N_12715,N_11800,N_10594);
or U12716 (N_12716,N_11244,N_10588);
and U12717 (N_12717,N_11965,N_11423);
nand U12718 (N_12718,N_11560,N_10531);
xor U12719 (N_12719,N_10713,N_11123);
nor U12720 (N_12720,N_11502,N_11967);
and U12721 (N_12721,N_11271,N_10654);
nor U12722 (N_12722,N_11918,N_10535);
nor U12723 (N_12723,N_11262,N_10673);
nand U12724 (N_12724,N_11047,N_10683);
or U12725 (N_12725,N_11135,N_10556);
or U12726 (N_12726,N_11599,N_11264);
xnor U12727 (N_12727,N_11623,N_10741);
or U12728 (N_12728,N_10742,N_11529);
xnor U12729 (N_12729,N_10938,N_10572);
nand U12730 (N_12730,N_11373,N_11537);
nand U12731 (N_12731,N_11215,N_11393);
nand U12732 (N_12732,N_11498,N_11012);
nand U12733 (N_12733,N_11044,N_10981);
xnor U12734 (N_12734,N_11338,N_11054);
nand U12735 (N_12735,N_10913,N_10716);
and U12736 (N_12736,N_11981,N_10782);
nand U12737 (N_12737,N_11759,N_11208);
or U12738 (N_12738,N_10740,N_11173);
xor U12739 (N_12739,N_11113,N_11260);
or U12740 (N_12740,N_10516,N_11801);
or U12741 (N_12741,N_11527,N_10836);
and U12742 (N_12742,N_10579,N_10954);
or U12743 (N_12743,N_10545,N_11841);
or U12744 (N_12744,N_11347,N_11060);
nand U12745 (N_12745,N_11000,N_11513);
nor U12746 (N_12746,N_10964,N_11287);
xnor U12747 (N_12747,N_11142,N_11495);
xor U12748 (N_12748,N_11657,N_11464);
and U12749 (N_12749,N_11876,N_11661);
nor U12750 (N_12750,N_11131,N_10708);
xor U12751 (N_12751,N_10911,N_11574);
nor U12752 (N_12752,N_10851,N_10763);
nor U12753 (N_12753,N_11835,N_11482);
and U12754 (N_12754,N_11632,N_10628);
nor U12755 (N_12755,N_11330,N_10728);
nand U12756 (N_12756,N_11762,N_11234);
xor U12757 (N_12757,N_11377,N_11450);
nand U12758 (N_12758,N_11408,N_11478);
nor U12759 (N_12759,N_10541,N_11140);
nand U12760 (N_12760,N_11415,N_11452);
xnor U12761 (N_12761,N_11978,N_11414);
and U12762 (N_12762,N_10870,N_10780);
nand U12763 (N_12763,N_10880,N_10562);
and U12764 (N_12764,N_11223,N_11180);
nor U12765 (N_12765,N_11781,N_11691);
or U12766 (N_12766,N_10708,N_10537);
or U12767 (N_12767,N_10760,N_10563);
nor U12768 (N_12768,N_11002,N_11869);
and U12769 (N_12769,N_11985,N_10610);
nor U12770 (N_12770,N_11398,N_10950);
and U12771 (N_12771,N_11215,N_10914);
or U12772 (N_12772,N_10681,N_11886);
and U12773 (N_12773,N_11739,N_11450);
xor U12774 (N_12774,N_11131,N_11371);
nand U12775 (N_12775,N_11687,N_11469);
nand U12776 (N_12776,N_11078,N_11372);
nor U12777 (N_12777,N_11966,N_11615);
xor U12778 (N_12778,N_11950,N_11600);
nor U12779 (N_12779,N_11960,N_11110);
xor U12780 (N_12780,N_11373,N_10925);
nand U12781 (N_12781,N_10960,N_11536);
nand U12782 (N_12782,N_11736,N_10869);
and U12783 (N_12783,N_11647,N_11600);
and U12784 (N_12784,N_11280,N_10972);
and U12785 (N_12785,N_11904,N_11327);
nor U12786 (N_12786,N_11807,N_11462);
and U12787 (N_12787,N_10508,N_10938);
nand U12788 (N_12788,N_11983,N_11523);
and U12789 (N_12789,N_11989,N_11623);
or U12790 (N_12790,N_11049,N_10863);
and U12791 (N_12791,N_10946,N_10960);
xnor U12792 (N_12792,N_10550,N_11110);
nand U12793 (N_12793,N_10731,N_11036);
xor U12794 (N_12794,N_11263,N_11688);
xor U12795 (N_12795,N_11567,N_11189);
or U12796 (N_12796,N_11633,N_10907);
xor U12797 (N_12797,N_10669,N_11860);
or U12798 (N_12798,N_10790,N_11113);
nor U12799 (N_12799,N_11954,N_11070);
nand U12800 (N_12800,N_10903,N_11816);
nand U12801 (N_12801,N_10968,N_10524);
nor U12802 (N_12802,N_10666,N_11640);
and U12803 (N_12803,N_11416,N_11312);
nor U12804 (N_12804,N_10589,N_11412);
or U12805 (N_12805,N_11861,N_10765);
nand U12806 (N_12806,N_10778,N_11862);
or U12807 (N_12807,N_10729,N_10798);
or U12808 (N_12808,N_11149,N_11935);
or U12809 (N_12809,N_11234,N_11254);
or U12810 (N_12810,N_11088,N_11344);
nand U12811 (N_12811,N_11662,N_11183);
nand U12812 (N_12812,N_11216,N_10915);
and U12813 (N_12813,N_11979,N_10719);
and U12814 (N_12814,N_11010,N_11153);
nand U12815 (N_12815,N_11776,N_10670);
and U12816 (N_12816,N_11606,N_11802);
xor U12817 (N_12817,N_10767,N_11196);
or U12818 (N_12818,N_11778,N_11810);
or U12819 (N_12819,N_11303,N_11978);
nor U12820 (N_12820,N_11654,N_11856);
nand U12821 (N_12821,N_11854,N_11827);
or U12822 (N_12822,N_11004,N_10953);
or U12823 (N_12823,N_11729,N_11325);
nor U12824 (N_12824,N_11906,N_11921);
nor U12825 (N_12825,N_11224,N_10525);
nor U12826 (N_12826,N_10549,N_10901);
nor U12827 (N_12827,N_11533,N_10634);
and U12828 (N_12828,N_11124,N_11611);
xor U12829 (N_12829,N_10773,N_11392);
nand U12830 (N_12830,N_11816,N_11564);
nand U12831 (N_12831,N_11200,N_10544);
nor U12832 (N_12832,N_11419,N_11783);
and U12833 (N_12833,N_10921,N_11008);
nand U12834 (N_12834,N_10860,N_11987);
xnor U12835 (N_12835,N_11875,N_11662);
or U12836 (N_12836,N_10772,N_10598);
or U12837 (N_12837,N_10761,N_10863);
nand U12838 (N_12838,N_10503,N_11797);
or U12839 (N_12839,N_10824,N_11098);
xor U12840 (N_12840,N_11765,N_10832);
nor U12841 (N_12841,N_11242,N_11879);
nor U12842 (N_12842,N_11530,N_11144);
nor U12843 (N_12843,N_11718,N_11451);
or U12844 (N_12844,N_11664,N_11712);
nand U12845 (N_12845,N_10626,N_10619);
nor U12846 (N_12846,N_11457,N_10520);
nand U12847 (N_12847,N_11327,N_11482);
xnor U12848 (N_12848,N_11213,N_10759);
nand U12849 (N_12849,N_11286,N_10970);
nand U12850 (N_12850,N_10690,N_11513);
nor U12851 (N_12851,N_11062,N_11055);
nand U12852 (N_12852,N_11036,N_11615);
nor U12853 (N_12853,N_10509,N_11750);
nand U12854 (N_12854,N_11356,N_11910);
nor U12855 (N_12855,N_11786,N_10915);
or U12856 (N_12856,N_11441,N_10679);
nor U12857 (N_12857,N_11482,N_11909);
and U12858 (N_12858,N_11486,N_11006);
or U12859 (N_12859,N_10501,N_10869);
and U12860 (N_12860,N_11203,N_11486);
or U12861 (N_12861,N_11860,N_11390);
and U12862 (N_12862,N_11837,N_11836);
or U12863 (N_12863,N_11518,N_11104);
xnor U12864 (N_12864,N_11813,N_11688);
xnor U12865 (N_12865,N_10909,N_11640);
nor U12866 (N_12866,N_10523,N_10997);
and U12867 (N_12867,N_11781,N_11180);
nor U12868 (N_12868,N_11756,N_11395);
nand U12869 (N_12869,N_10992,N_10999);
xor U12870 (N_12870,N_11277,N_11099);
nand U12871 (N_12871,N_11730,N_11883);
and U12872 (N_12872,N_10722,N_10940);
and U12873 (N_12873,N_11515,N_10570);
nand U12874 (N_12874,N_11656,N_11998);
and U12875 (N_12875,N_11361,N_11754);
xnor U12876 (N_12876,N_10790,N_11871);
or U12877 (N_12877,N_11856,N_11718);
xor U12878 (N_12878,N_10813,N_10645);
or U12879 (N_12879,N_11486,N_10973);
nor U12880 (N_12880,N_10760,N_11550);
xnor U12881 (N_12881,N_11557,N_10939);
xor U12882 (N_12882,N_11669,N_11821);
nand U12883 (N_12883,N_11147,N_11884);
nor U12884 (N_12884,N_11791,N_11826);
xor U12885 (N_12885,N_10627,N_11992);
nor U12886 (N_12886,N_11819,N_10961);
or U12887 (N_12887,N_10943,N_11730);
nand U12888 (N_12888,N_10822,N_11586);
and U12889 (N_12889,N_11951,N_11302);
or U12890 (N_12890,N_11665,N_11131);
nand U12891 (N_12891,N_11622,N_10725);
xnor U12892 (N_12892,N_11541,N_11565);
nand U12893 (N_12893,N_11530,N_11113);
nor U12894 (N_12894,N_11704,N_10820);
and U12895 (N_12895,N_11383,N_11396);
nor U12896 (N_12896,N_11260,N_11064);
xor U12897 (N_12897,N_10667,N_11686);
xor U12898 (N_12898,N_10983,N_11737);
xor U12899 (N_12899,N_10597,N_10738);
nand U12900 (N_12900,N_11120,N_11681);
xor U12901 (N_12901,N_11123,N_11700);
nor U12902 (N_12902,N_11162,N_11708);
nor U12903 (N_12903,N_11605,N_11627);
nand U12904 (N_12904,N_10815,N_11239);
and U12905 (N_12905,N_11981,N_10874);
xor U12906 (N_12906,N_10886,N_11528);
xnor U12907 (N_12907,N_11980,N_11612);
nor U12908 (N_12908,N_10640,N_11866);
nand U12909 (N_12909,N_10561,N_11639);
and U12910 (N_12910,N_11313,N_11647);
xor U12911 (N_12911,N_11983,N_11126);
xnor U12912 (N_12912,N_10790,N_11037);
nor U12913 (N_12913,N_10864,N_11263);
and U12914 (N_12914,N_11464,N_11659);
nor U12915 (N_12915,N_10900,N_11923);
and U12916 (N_12916,N_11839,N_11417);
xnor U12917 (N_12917,N_11004,N_11288);
nor U12918 (N_12918,N_11200,N_11509);
nand U12919 (N_12919,N_11658,N_11210);
xor U12920 (N_12920,N_10811,N_11805);
or U12921 (N_12921,N_11600,N_10872);
xor U12922 (N_12922,N_11527,N_11239);
nand U12923 (N_12923,N_11150,N_11421);
and U12924 (N_12924,N_11110,N_11477);
xnor U12925 (N_12925,N_11058,N_11407);
and U12926 (N_12926,N_10677,N_11337);
nor U12927 (N_12927,N_11921,N_11405);
nor U12928 (N_12928,N_10967,N_10805);
or U12929 (N_12929,N_10690,N_11281);
or U12930 (N_12930,N_10716,N_11430);
nor U12931 (N_12931,N_11486,N_11818);
nor U12932 (N_12932,N_11691,N_10685);
nand U12933 (N_12933,N_11655,N_10585);
xnor U12934 (N_12934,N_11226,N_11726);
and U12935 (N_12935,N_10622,N_11140);
xnor U12936 (N_12936,N_11712,N_11709);
nor U12937 (N_12937,N_11843,N_11398);
and U12938 (N_12938,N_10670,N_10824);
nand U12939 (N_12939,N_10548,N_11559);
xor U12940 (N_12940,N_10618,N_10599);
xnor U12941 (N_12941,N_11322,N_11808);
xnor U12942 (N_12942,N_11666,N_10713);
xor U12943 (N_12943,N_10807,N_11067);
or U12944 (N_12944,N_11327,N_10520);
xor U12945 (N_12945,N_10775,N_11040);
nand U12946 (N_12946,N_10669,N_11989);
xnor U12947 (N_12947,N_11513,N_11578);
nor U12948 (N_12948,N_11844,N_10833);
and U12949 (N_12949,N_10795,N_11076);
nand U12950 (N_12950,N_10825,N_11547);
and U12951 (N_12951,N_11399,N_11501);
xnor U12952 (N_12952,N_11000,N_10763);
xor U12953 (N_12953,N_11543,N_11561);
or U12954 (N_12954,N_10875,N_10817);
and U12955 (N_12955,N_10927,N_10559);
or U12956 (N_12956,N_10517,N_11688);
or U12957 (N_12957,N_10526,N_11885);
xnor U12958 (N_12958,N_11555,N_11543);
and U12959 (N_12959,N_11676,N_11172);
nor U12960 (N_12960,N_11958,N_10713);
nor U12961 (N_12961,N_10969,N_10824);
nand U12962 (N_12962,N_11018,N_10611);
nor U12963 (N_12963,N_11656,N_10502);
and U12964 (N_12964,N_10758,N_11401);
or U12965 (N_12965,N_11380,N_10614);
nor U12966 (N_12966,N_11946,N_10729);
xnor U12967 (N_12967,N_11717,N_11288);
nor U12968 (N_12968,N_11926,N_10995);
nor U12969 (N_12969,N_11955,N_11542);
nand U12970 (N_12970,N_11965,N_10708);
nand U12971 (N_12971,N_10892,N_11352);
and U12972 (N_12972,N_10723,N_10551);
xnor U12973 (N_12973,N_10619,N_11085);
nor U12974 (N_12974,N_11757,N_11297);
nor U12975 (N_12975,N_11969,N_11007);
or U12976 (N_12976,N_11122,N_10635);
nor U12977 (N_12977,N_10556,N_11848);
or U12978 (N_12978,N_10571,N_11023);
nand U12979 (N_12979,N_11592,N_10582);
and U12980 (N_12980,N_11098,N_10874);
nor U12981 (N_12981,N_11364,N_11365);
nand U12982 (N_12982,N_11934,N_11849);
nor U12983 (N_12983,N_10571,N_10553);
nor U12984 (N_12984,N_11729,N_10748);
and U12985 (N_12985,N_10953,N_10543);
nand U12986 (N_12986,N_11059,N_10573);
and U12987 (N_12987,N_10582,N_10564);
or U12988 (N_12988,N_10732,N_10740);
and U12989 (N_12989,N_11240,N_11027);
and U12990 (N_12990,N_11015,N_11814);
nor U12991 (N_12991,N_10506,N_11682);
xnor U12992 (N_12992,N_11180,N_11862);
or U12993 (N_12993,N_11259,N_10567);
nand U12994 (N_12994,N_11251,N_10895);
nor U12995 (N_12995,N_10676,N_11224);
nand U12996 (N_12996,N_11149,N_11835);
nand U12997 (N_12997,N_11673,N_10994);
or U12998 (N_12998,N_11673,N_10750);
xor U12999 (N_12999,N_11746,N_10989);
nor U13000 (N_13000,N_11436,N_11920);
nor U13001 (N_13001,N_11292,N_11859);
nor U13002 (N_13002,N_11587,N_11355);
or U13003 (N_13003,N_11409,N_10979);
or U13004 (N_13004,N_10755,N_11172);
nor U13005 (N_13005,N_10840,N_10708);
xor U13006 (N_13006,N_11167,N_10752);
nor U13007 (N_13007,N_10616,N_11244);
nor U13008 (N_13008,N_10728,N_11103);
xnor U13009 (N_13009,N_11852,N_11273);
and U13010 (N_13010,N_10715,N_10663);
xor U13011 (N_13011,N_11312,N_10933);
nor U13012 (N_13012,N_10861,N_10985);
nand U13013 (N_13013,N_11827,N_11831);
nand U13014 (N_13014,N_10629,N_10568);
or U13015 (N_13015,N_10802,N_11629);
nand U13016 (N_13016,N_11304,N_11055);
and U13017 (N_13017,N_10816,N_11968);
nand U13018 (N_13018,N_11670,N_10790);
xnor U13019 (N_13019,N_10997,N_11506);
nor U13020 (N_13020,N_10606,N_10684);
xor U13021 (N_13021,N_11192,N_11680);
xnor U13022 (N_13022,N_11240,N_10780);
or U13023 (N_13023,N_11385,N_10906);
xor U13024 (N_13024,N_11327,N_11116);
xnor U13025 (N_13025,N_10556,N_11551);
or U13026 (N_13026,N_10643,N_11209);
and U13027 (N_13027,N_11720,N_10683);
or U13028 (N_13028,N_11215,N_11137);
nor U13029 (N_13029,N_10518,N_11891);
nor U13030 (N_13030,N_11136,N_10929);
nand U13031 (N_13031,N_11347,N_10742);
xor U13032 (N_13032,N_11412,N_11197);
nor U13033 (N_13033,N_10845,N_11731);
and U13034 (N_13034,N_11735,N_10838);
and U13035 (N_13035,N_10866,N_11957);
and U13036 (N_13036,N_10575,N_11209);
or U13037 (N_13037,N_11631,N_11446);
nand U13038 (N_13038,N_11896,N_11578);
and U13039 (N_13039,N_11848,N_11907);
or U13040 (N_13040,N_11798,N_11958);
xor U13041 (N_13041,N_11517,N_10780);
and U13042 (N_13042,N_10980,N_10834);
nor U13043 (N_13043,N_10721,N_10651);
nor U13044 (N_13044,N_11042,N_11294);
nor U13045 (N_13045,N_10999,N_10584);
and U13046 (N_13046,N_11296,N_10526);
nor U13047 (N_13047,N_11265,N_11341);
nand U13048 (N_13048,N_11495,N_10979);
or U13049 (N_13049,N_11844,N_11871);
nand U13050 (N_13050,N_11729,N_11285);
nand U13051 (N_13051,N_11915,N_11015);
xor U13052 (N_13052,N_11822,N_11057);
xnor U13053 (N_13053,N_10537,N_11092);
xnor U13054 (N_13054,N_10542,N_10963);
or U13055 (N_13055,N_11394,N_11476);
and U13056 (N_13056,N_11497,N_11536);
or U13057 (N_13057,N_11949,N_10767);
nand U13058 (N_13058,N_10641,N_11559);
nor U13059 (N_13059,N_11949,N_10964);
nand U13060 (N_13060,N_10591,N_10946);
nand U13061 (N_13061,N_11593,N_11418);
and U13062 (N_13062,N_11616,N_11347);
and U13063 (N_13063,N_10867,N_11055);
nor U13064 (N_13064,N_11486,N_11998);
nor U13065 (N_13065,N_11154,N_11239);
xnor U13066 (N_13066,N_10718,N_11781);
nand U13067 (N_13067,N_10919,N_11806);
nor U13068 (N_13068,N_10856,N_11532);
and U13069 (N_13069,N_10623,N_10797);
or U13070 (N_13070,N_10978,N_11174);
or U13071 (N_13071,N_11022,N_11321);
and U13072 (N_13072,N_11225,N_11684);
xor U13073 (N_13073,N_11180,N_10544);
nor U13074 (N_13074,N_10595,N_11211);
xnor U13075 (N_13075,N_10817,N_10879);
xor U13076 (N_13076,N_10984,N_10940);
and U13077 (N_13077,N_11863,N_10621);
and U13078 (N_13078,N_11408,N_11804);
nand U13079 (N_13079,N_10710,N_11539);
and U13080 (N_13080,N_11947,N_10839);
nand U13081 (N_13081,N_10843,N_10602);
nand U13082 (N_13082,N_10849,N_10971);
nor U13083 (N_13083,N_10726,N_11094);
nor U13084 (N_13084,N_11857,N_10945);
nor U13085 (N_13085,N_11631,N_10821);
nand U13086 (N_13086,N_11848,N_10632);
nand U13087 (N_13087,N_11596,N_11600);
or U13088 (N_13088,N_10582,N_10541);
and U13089 (N_13089,N_11199,N_10684);
xor U13090 (N_13090,N_11171,N_11259);
nor U13091 (N_13091,N_11730,N_11890);
nor U13092 (N_13092,N_11129,N_11946);
nor U13093 (N_13093,N_11454,N_11753);
or U13094 (N_13094,N_11837,N_10877);
nor U13095 (N_13095,N_11581,N_11804);
xnor U13096 (N_13096,N_10936,N_10603);
and U13097 (N_13097,N_11861,N_11341);
and U13098 (N_13098,N_11536,N_10701);
nor U13099 (N_13099,N_11331,N_11111);
nor U13100 (N_13100,N_10944,N_11423);
or U13101 (N_13101,N_11395,N_11494);
nor U13102 (N_13102,N_11563,N_11701);
nor U13103 (N_13103,N_11908,N_10681);
nand U13104 (N_13104,N_11618,N_11712);
nor U13105 (N_13105,N_11197,N_11856);
or U13106 (N_13106,N_10793,N_11448);
and U13107 (N_13107,N_10800,N_11867);
nand U13108 (N_13108,N_11211,N_11754);
xnor U13109 (N_13109,N_10974,N_11528);
nand U13110 (N_13110,N_10567,N_11558);
or U13111 (N_13111,N_11410,N_11752);
and U13112 (N_13112,N_11524,N_10537);
or U13113 (N_13113,N_11172,N_11725);
xor U13114 (N_13114,N_11530,N_10633);
xor U13115 (N_13115,N_11981,N_11376);
nor U13116 (N_13116,N_10925,N_10798);
nand U13117 (N_13117,N_11084,N_10533);
and U13118 (N_13118,N_10839,N_11051);
nand U13119 (N_13119,N_11358,N_11846);
or U13120 (N_13120,N_11483,N_11985);
nor U13121 (N_13121,N_11925,N_10542);
xor U13122 (N_13122,N_10946,N_10991);
nand U13123 (N_13123,N_11330,N_11226);
and U13124 (N_13124,N_11089,N_11378);
xor U13125 (N_13125,N_11022,N_11260);
nor U13126 (N_13126,N_10793,N_10873);
xor U13127 (N_13127,N_11259,N_11580);
nor U13128 (N_13128,N_10519,N_11193);
or U13129 (N_13129,N_11869,N_11329);
nor U13130 (N_13130,N_11104,N_11849);
xnor U13131 (N_13131,N_11622,N_11535);
nor U13132 (N_13132,N_11593,N_10681);
nor U13133 (N_13133,N_10601,N_11653);
nor U13134 (N_13134,N_11457,N_11120);
nor U13135 (N_13135,N_10847,N_10898);
or U13136 (N_13136,N_10999,N_11257);
or U13137 (N_13137,N_10829,N_10976);
and U13138 (N_13138,N_11493,N_10782);
xor U13139 (N_13139,N_11907,N_11043);
and U13140 (N_13140,N_10565,N_10596);
or U13141 (N_13141,N_11272,N_11748);
nand U13142 (N_13142,N_11788,N_11036);
or U13143 (N_13143,N_11326,N_11525);
nand U13144 (N_13144,N_11979,N_11419);
xor U13145 (N_13145,N_10928,N_10644);
and U13146 (N_13146,N_11318,N_11262);
and U13147 (N_13147,N_11203,N_11265);
nor U13148 (N_13148,N_11406,N_11804);
nand U13149 (N_13149,N_10711,N_11495);
nor U13150 (N_13150,N_11231,N_11198);
nor U13151 (N_13151,N_10951,N_11499);
or U13152 (N_13152,N_11812,N_10999);
or U13153 (N_13153,N_11098,N_11315);
and U13154 (N_13154,N_10608,N_10652);
or U13155 (N_13155,N_11601,N_11719);
nand U13156 (N_13156,N_11573,N_10727);
and U13157 (N_13157,N_11232,N_10710);
nand U13158 (N_13158,N_11464,N_11801);
or U13159 (N_13159,N_11649,N_11698);
nor U13160 (N_13160,N_11508,N_11967);
or U13161 (N_13161,N_10500,N_11706);
nand U13162 (N_13162,N_10846,N_11002);
xnor U13163 (N_13163,N_11883,N_10595);
or U13164 (N_13164,N_10525,N_10914);
nand U13165 (N_13165,N_11029,N_10572);
xor U13166 (N_13166,N_10988,N_10619);
xnor U13167 (N_13167,N_11201,N_11593);
and U13168 (N_13168,N_11805,N_11571);
nand U13169 (N_13169,N_11300,N_11352);
and U13170 (N_13170,N_11579,N_11390);
or U13171 (N_13171,N_11838,N_11244);
xor U13172 (N_13172,N_11081,N_11053);
xor U13173 (N_13173,N_11407,N_11796);
and U13174 (N_13174,N_11925,N_11381);
nand U13175 (N_13175,N_11800,N_11216);
xnor U13176 (N_13176,N_10823,N_11213);
nand U13177 (N_13177,N_11041,N_11913);
xor U13178 (N_13178,N_11648,N_10636);
nor U13179 (N_13179,N_11732,N_11752);
xor U13180 (N_13180,N_11225,N_10981);
xnor U13181 (N_13181,N_11732,N_11000);
or U13182 (N_13182,N_10684,N_10616);
and U13183 (N_13183,N_11836,N_11486);
or U13184 (N_13184,N_11674,N_11458);
and U13185 (N_13185,N_11167,N_11937);
or U13186 (N_13186,N_11642,N_10546);
nor U13187 (N_13187,N_10656,N_10744);
xnor U13188 (N_13188,N_11904,N_10820);
and U13189 (N_13189,N_11723,N_11935);
nor U13190 (N_13190,N_10603,N_10567);
nor U13191 (N_13191,N_11442,N_11618);
nor U13192 (N_13192,N_10948,N_11035);
and U13193 (N_13193,N_10671,N_10516);
or U13194 (N_13194,N_11697,N_11251);
nor U13195 (N_13195,N_11353,N_10621);
nand U13196 (N_13196,N_10886,N_10617);
nor U13197 (N_13197,N_11020,N_11206);
or U13198 (N_13198,N_11070,N_11330);
or U13199 (N_13199,N_11875,N_11265);
and U13200 (N_13200,N_11773,N_10912);
and U13201 (N_13201,N_11704,N_10615);
or U13202 (N_13202,N_10848,N_11877);
and U13203 (N_13203,N_10922,N_11602);
or U13204 (N_13204,N_11515,N_11886);
or U13205 (N_13205,N_11402,N_11562);
or U13206 (N_13206,N_11688,N_10507);
xnor U13207 (N_13207,N_11186,N_11944);
and U13208 (N_13208,N_11722,N_10568);
nand U13209 (N_13209,N_10853,N_11789);
nor U13210 (N_13210,N_11818,N_10706);
xnor U13211 (N_13211,N_11610,N_11640);
nand U13212 (N_13212,N_11368,N_11915);
nand U13213 (N_13213,N_10655,N_10604);
and U13214 (N_13214,N_11929,N_10881);
or U13215 (N_13215,N_11667,N_11982);
nor U13216 (N_13216,N_11669,N_11677);
xor U13217 (N_13217,N_11271,N_10750);
xnor U13218 (N_13218,N_11259,N_11600);
and U13219 (N_13219,N_11448,N_10734);
nand U13220 (N_13220,N_10688,N_11858);
nor U13221 (N_13221,N_11502,N_10973);
and U13222 (N_13222,N_11798,N_11801);
nand U13223 (N_13223,N_10704,N_10733);
nor U13224 (N_13224,N_11641,N_11027);
and U13225 (N_13225,N_10723,N_11414);
xor U13226 (N_13226,N_10857,N_11519);
or U13227 (N_13227,N_10727,N_11214);
nand U13228 (N_13228,N_10689,N_10641);
xor U13229 (N_13229,N_11506,N_11790);
xnor U13230 (N_13230,N_11506,N_11277);
xnor U13231 (N_13231,N_10545,N_11385);
nand U13232 (N_13232,N_11389,N_10584);
nand U13233 (N_13233,N_11841,N_11925);
or U13234 (N_13234,N_11240,N_11888);
nand U13235 (N_13235,N_10901,N_11537);
nand U13236 (N_13236,N_10523,N_11927);
or U13237 (N_13237,N_10628,N_11337);
or U13238 (N_13238,N_10730,N_11123);
and U13239 (N_13239,N_11142,N_10586);
xnor U13240 (N_13240,N_10630,N_11879);
xor U13241 (N_13241,N_10586,N_11446);
or U13242 (N_13242,N_11872,N_10561);
xor U13243 (N_13243,N_10835,N_11295);
and U13244 (N_13244,N_11911,N_11395);
and U13245 (N_13245,N_11551,N_11835);
and U13246 (N_13246,N_10965,N_11071);
and U13247 (N_13247,N_10953,N_11611);
or U13248 (N_13248,N_11409,N_10640);
nand U13249 (N_13249,N_11147,N_10991);
nor U13250 (N_13250,N_11194,N_11801);
or U13251 (N_13251,N_11317,N_10831);
nor U13252 (N_13252,N_10638,N_11208);
or U13253 (N_13253,N_11734,N_11190);
and U13254 (N_13254,N_11618,N_10648);
xor U13255 (N_13255,N_11612,N_11138);
and U13256 (N_13256,N_11977,N_10987);
and U13257 (N_13257,N_11038,N_11980);
xnor U13258 (N_13258,N_10920,N_11811);
and U13259 (N_13259,N_11284,N_11497);
and U13260 (N_13260,N_11848,N_11780);
nand U13261 (N_13261,N_11328,N_11964);
and U13262 (N_13262,N_11438,N_11237);
nor U13263 (N_13263,N_11271,N_11798);
nor U13264 (N_13264,N_11482,N_11433);
nand U13265 (N_13265,N_10557,N_11898);
nor U13266 (N_13266,N_10791,N_10958);
xnor U13267 (N_13267,N_10617,N_11249);
and U13268 (N_13268,N_10749,N_11640);
nor U13269 (N_13269,N_10674,N_10994);
nor U13270 (N_13270,N_11653,N_10967);
or U13271 (N_13271,N_10537,N_11905);
xor U13272 (N_13272,N_10633,N_10577);
xor U13273 (N_13273,N_11369,N_11523);
nor U13274 (N_13274,N_11536,N_11842);
or U13275 (N_13275,N_11384,N_10703);
or U13276 (N_13276,N_11572,N_10833);
and U13277 (N_13277,N_10944,N_10874);
and U13278 (N_13278,N_11456,N_11609);
or U13279 (N_13279,N_10634,N_11689);
nand U13280 (N_13280,N_11979,N_11289);
xnor U13281 (N_13281,N_11460,N_10791);
nor U13282 (N_13282,N_11375,N_11568);
and U13283 (N_13283,N_10993,N_10808);
nor U13284 (N_13284,N_11158,N_11721);
nor U13285 (N_13285,N_11347,N_10987);
xnor U13286 (N_13286,N_11523,N_10985);
nand U13287 (N_13287,N_11646,N_11510);
nand U13288 (N_13288,N_11325,N_11680);
xor U13289 (N_13289,N_11219,N_11325);
xor U13290 (N_13290,N_11246,N_10873);
or U13291 (N_13291,N_11289,N_11903);
nor U13292 (N_13292,N_10565,N_10708);
and U13293 (N_13293,N_10962,N_10698);
xnor U13294 (N_13294,N_11055,N_10566);
nor U13295 (N_13295,N_10915,N_10674);
xnor U13296 (N_13296,N_10886,N_11353);
nand U13297 (N_13297,N_11287,N_11687);
nand U13298 (N_13298,N_11070,N_10762);
xor U13299 (N_13299,N_10665,N_10592);
nor U13300 (N_13300,N_11280,N_11847);
or U13301 (N_13301,N_11680,N_10857);
nor U13302 (N_13302,N_11307,N_10690);
or U13303 (N_13303,N_10964,N_11573);
xor U13304 (N_13304,N_11675,N_10849);
xor U13305 (N_13305,N_11920,N_11599);
or U13306 (N_13306,N_10813,N_11263);
xor U13307 (N_13307,N_11355,N_10646);
nand U13308 (N_13308,N_11241,N_11514);
nand U13309 (N_13309,N_11165,N_10591);
or U13310 (N_13310,N_11211,N_11177);
xnor U13311 (N_13311,N_11420,N_11298);
and U13312 (N_13312,N_11097,N_10907);
xnor U13313 (N_13313,N_11088,N_11398);
nor U13314 (N_13314,N_11098,N_11831);
nand U13315 (N_13315,N_11904,N_11367);
nand U13316 (N_13316,N_10560,N_11441);
or U13317 (N_13317,N_10863,N_11339);
or U13318 (N_13318,N_11762,N_11386);
xor U13319 (N_13319,N_11210,N_11675);
nor U13320 (N_13320,N_11067,N_11308);
nor U13321 (N_13321,N_11874,N_11187);
nand U13322 (N_13322,N_10573,N_10553);
and U13323 (N_13323,N_10908,N_10974);
nand U13324 (N_13324,N_11616,N_11709);
xnor U13325 (N_13325,N_11803,N_11309);
and U13326 (N_13326,N_10666,N_11150);
nor U13327 (N_13327,N_10688,N_11054);
or U13328 (N_13328,N_10847,N_11647);
or U13329 (N_13329,N_11984,N_11316);
nand U13330 (N_13330,N_11011,N_11868);
and U13331 (N_13331,N_11599,N_10756);
xor U13332 (N_13332,N_11641,N_10704);
nand U13333 (N_13333,N_11134,N_10580);
nor U13334 (N_13334,N_11175,N_11677);
xnor U13335 (N_13335,N_10723,N_11673);
xnor U13336 (N_13336,N_11316,N_10860);
or U13337 (N_13337,N_11817,N_11003);
xor U13338 (N_13338,N_10705,N_11212);
and U13339 (N_13339,N_11413,N_11675);
or U13340 (N_13340,N_11963,N_10959);
nand U13341 (N_13341,N_11220,N_11936);
nor U13342 (N_13342,N_10877,N_11065);
or U13343 (N_13343,N_11069,N_10549);
nand U13344 (N_13344,N_11221,N_11668);
nand U13345 (N_13345,N_10906,N_11370);
nand U13346 (N_13346,N_11103,N_11505);
nand U13347 (N_13347,N_11596,N_10989);
nor U13348 (N_13348,N_11331,N_10958);
and U13349 (N_13349,N_11313,N_11087);
and U13350 (N_13350,N_11707,N_11400);
or U13351 (N_13351,N_11587,N_11230);
nand U13352 (N_13352,N_10540,N_11559);
xor U13353 (N_13353,N_11997,N_11864);
xor U13354 (N_13354,N_11796,N_10872);
or U13355 (N_13355,N_11007,N_11559);
nor U13356 (N_13356,N_10632,N_11850);
nor U13357 (N_13357,N_11204,N_11287);
and U13358 (N_13358,N_11551,N_11641);
or U13359 (N_13359,N_11635,N_11570);
xnor U13360 (N_13360,N_11524,N_11779);
nor U13361 (N_13361,N_11177,N_10556);
and U13362 (N_13362,N_11366,N_10858);
nand U13363 (N_13363,N_11597,N_11892);
nand U13364 (N_13364,N_10821,N_11113);
nor U13365 (N_13365,N_11020,N_10878);
xor U13366 (N_13366,N_11644,N_11823);
nor U13367 (N_13367,N_11431,N_11218);
and U13368 (N_13368,N_11218,N_11162);
and U13369 (N_13369,N_11645,N_11560);
nand U13370 (N_13370,N_10739,N_11623);
nand U13371 (N_13371,N_10601,N_10767);
and U13372 (N_13372,N_10507,N_10723);
xor U13373 (N_13373,N_10670,N_10564);
nor U13374 (N_13374,N_11654,N_11778);
xor U13375 (N_13375,N_10507,N_11384);
xor U13376 (N_13376,N_10723,N_10739);
xnor U13377 (N_13377,N_11274,N_11051);
or U13378 (N_13378,N_11044,N_10974);
xnor U13379 (N_13379,N_11544,N_10520);
or U13380 (N_13380,N_11753,N_11793);
xor U13381 (N_13381,N_11850,N_11422);
xor U13382 (N_13382,N_11016,N_11616);
or U13383 (N_13383,N_10757,N_10981);
xor U13384 (N_13384,N_11991,N_11976);
nor U13385 (N_13385,N_10624,N_11087);
xnor U13386 (N_13386,N_10859,N_10821);
and U13387 (N_13387,N_10906,N_11026);
xor U13388 (N_13388,N_11913,N_11187);
nor U13389 (N_13389,N_11617,N_10697);
nand U13390 (N_13390,N_10980,N_11380);
nand U13391 (N_13391,N_11631,N_10961);
and U13392 (N_13392,N_11290,N_10600);
and U13393 (N_13393,N_11717,N_11125);
or U13394 (N_13394,N_10586,N_10697);
or U13395 (N_13395,N_11609,N_10778);
or U13396 (N_13396,N_11745,N_10507);
and U13397 (N_13397,N_11408,N_11787);
xnor U13398 (N_13398,N_11317,N_11050);
nor U13399 (N_13399,N_11948,N_11975);
or U13400 (N_13400,N_11132,N_10550);
nand U13401 (N_13401,N_11450,N_10598);
nand U13402 (N_13402,N_11129,N_11392);
xnor U13403 (N_13403,N_11093,N_11306);
and U13404 (N_13404,N_10541,N_11401);
nor U13405 (N_13405,N_10765,N_10659);
nor U13406 (N_13406,N_10758,N_11281);
nor U13407 (N_13407,N_10896,N_10538);
or U13408 (N_13408,N_11791,N_11286);
and U13409 (N_13409,N_10706,N_11024);
nor U13410 (N_13410,N_11407,N_10977);
xnor U13411 (N_13411,N_10577,N_10742);
nand U13412 (N_13412,N_11962,N_11091);
nand U13413 (N_13413,N_11541,N_11501);
nor U13414 (N_13414,N_10994,N_11140);
or U13415 (N_13415,N_10596,N_11286);
xnor U13416 (N_13416,N_11838,N_11164);
nor U13417 (N_13417,N_11033,N_11330);
nand U13418 (N_13418,N_11792,N_10993);
nor U13419 (N_13419,N_10543,N_11768);
nor U13420 (N_13420,N_11838,N_11219);
and U13421 (N_13421,N_11335,N_11781);
nor U13422 (N_13422,N_11874,N_11809);
nor U13423 (N_13423,N_10922,N_11865);
nor U13424 (N_13424,N_10862,N_11427);
nor U13425 (N_13425,N_11148,N_11414);
nand U13426 (N_13426,N_11014,N_10829);
and U13427 (N_13427,N_11172,N_11217);
nand U13428 (N_13428,N_10629,N_10635);
or U13429 (N_13429,N_10515,N_11588);
xor U13430 (N_13430,N_11576,N_11846);
nor U13431 (N_13431,N_11780,N_11592);
nand U13432 (N_13432,N_11332,N_10751);
xnor U13433 (N_13433,N_10517,N_10839);
and U13434 (N_13434,N_11877,N_11021);
or U13435 (N_13435,N_10692,N_11094);
xor U13436 (N_13436,N_11316,N_11978);
or U13437 (N_13437,N_11272,N_10774);
and U13438 (N_13438,N_11139,N_11461);
and U13439 (N_13439,N_11225,N_10644);
and U13440 (N_13440,N_10779,N_11298);
nor U13441 (N_13441,N_11742,N_10618);
and U13442 (N_13442,N_10660,N_10977);
or U13443 (N_13443,N_11733,N_11332);
xor U13444 (N_13444,N_10790,N_10880);
xor U13445 (N_13445,N_10937,N_10540);
xor U13446 (N_13446,N_11447,N_11389);
xor U13447 (N_13447,N_11076,N_10995);
nor U13448 (N_13448,N_10842,N_10722);
or U13449 (N_13449,N_11157,N_11251);
nand U13450 (N_13450,N_11178,N_10707);
xor U13451 (N_13451,N_10597,N_11589);
xnor U13452 (N_13452,N_10550,N_10506);
or U13453 (N_13453,N_11822,N_11985);
nor U13454 (N_13454,N_10897,N_10559);
and U13455 (N_13455,N_11162,N_11696);
or U13456 (N_13456,N_10906,N_11960);
and U13457 (N_13457,N_11746,N_10726);
nand U13458 (N_13458,N_10940,N_10806);
or U13459 (N_13459,N_11701,N_11735);
nand U13460 (N_13460,N_10696,N_10784);
and U13461 (N_13461,N_11383,N_11516);
nor U13462 (N_13462,N_10852,N_11299);
and U13463 (N_13463,N_10904,N_11221);
and U13464 (N_13464,N_11730,N_11559);
nand U13465 (N_13465,N_11662,N_10570);
and U13466 (N_13466,N_10656,N_11013);
or U13467 (N_13467,N_10798,N_10792);
nand U13468 (N_13468,N_11252,N_11201);
or U13469 (N_13469,N_10742,N_10877);
nor U13470 (N_13470,N_11394,N_11670);
xor U13471 (N_13471,N_10658,N_10852);
and U13472 (N_13472,N_11090,N_10581);
and U13473 (N_13473,N_10723,N_11007);
nand U13474 (N_13474,N_10959,N_10846);
nor U13475 (N_13475,N_11307,N_11917);
nand U13476 (N_13476,N_11824,N_11500);
and U13477 (N_13477,N_10591,N_11172);
nand U13478 (N_13478,N_11055,N_10945);
nor U13479 (N_13479,N_11646,N_10709);
xnor U13480 (N_13480,N_11424,N_10828);
or U13481 (N_13481,N_11213,N_11469);
nand U13482 (N_13482,N_10542,N_10933);
xor U13483 (N_13483,N_11356,N_11433);
nor U13484 (N_13484,N_10806,N_11921);
nand U13485 (N_13485,N_11196,N_11022);
nand U13486 (N_13486,N_10715,N_10598);
and U13487 (N_13487,N_10694,N_11014);
or U13488 (N_13488,N_11858,N_10843);
xor U13489 (N_13489,N_11892,N_11064);
nor U13490 (N_13490,N_11086,N_10893);
xnor U13491 (N_13491,N_10753,N_11829);
nand U13492 (N_13492,N_11317,N_11239);
nor U13493 (N_13493,N_10922,N_11205);
nand U13494 (N_13494,N_10819,N_11018);
or U13495 (N_13495,N_10990,N_11685);
nand U13496 (N_13496,N_11774,N_11805);
or U13497 (N_13497,N_10817,N_11651);
nand U13498 (N_13498,N_11637,N_10869);
nand U13499 (N_13499,N_11602,N_11448);
nor U13500 (N_13500,N_12388,N_13211);
or U13501 (N_13501,N_12023,N_13010);
or U13502 (N_13502,N_12424,N_12116);
xor U13503 (N_13503,N_12902,N_12532);
nor U13504 (N_13504,N_13460,N_12262);
xnor U13505 (N_13505,N_12406,N_12491);
nor U13506 (N_13506,N_12544,N_13375);
nand U13507 (N_13507,N_12346,N_12697);
and U13508 (N_13508,N_12257,N_12530);
or U13509 (N_13509,N_12175,N_13086);
nor U13510 (N_13510,N_12502,N_12205);
and U13511 (N_13511,N_12075,N_13120);
nand U13512 (N_13512,N_12467,N_13224);
nor U13513 (N_13513,N_13112,N_13268);
xnor U13514 (N_13514,N_12417,N_13118);
and U13515 (N_13515,N_12165,N_12831);
nand U13516 (N_13516,N_12947,N_13472);
and U13517 (N_13517,N_13279,N_12071);
and U13518 (N_13518,N_12107,N_12315);
nor U13519 (N_13519,N_12999,N_12508);
and U13520 (N_13520,N_12885,N_12275);
nor U13521 (N_13521,N_12726,N_12207);
nor U13522 (N_13522,N_12084,N_12110);
or U13523 (N_13523,N_13180,N_12523);
nor U13524 (N_13524,N_12933,N_12171);
nand U13525 (N_13525,N_12358,N_12874);
and U13526 (N_13526,N_12799,N_12036);
or U13527 (N_13527,N_13035,N_12626);
and U13528 (N_13528,N_12568,N_12056);
nand U13529 (N_13529,N_12479,N_13148);
or U13530 (N_13530,N_13184,N_12377);
nand U13531 (N_13531,N_13384,N_12890);
nand U13532 (N_13532,N_13027,N_13365);
nor U13533 (N_13533,N_12781,N_12640);
nand U13534 (N_13534,N_12436,N_13030);
nor U13535 (N_13535,N_12836,N_12181);
nand U13536 (N_13536,N_12382,N_12334);
or U13537 (N_13537,N_12385,N_12952);
xnor U13538 (N_13538,N_13139,N_12266);
nand U13539 (N_13539,N_12279,N_13473);
nand U13540 (N_13540,N_13409,N_13443);
nand U13541 (N_13541,N_12895,N_12119);
nand U13542 (N_13542,N_12337,N_13267);
nand U13543 (N_13543,N_13069,N_12345);
and U13544 (N_13544,N_13194,N_12540);
xnor U13545 (N_13545,N_12583,N_12151);
nor U13546 (N_13546,N_12734,N_13039);
xnor U13547 (N_13547,N_13372,N_13026);
and U13548 (N_13548,N_12797,N_12559);
and U13549 (N_13549,N_13437,N_12187);
nand U13550 (N_13550,N_12839,N_12659);
and U13551 (N_13551,N_12919,N_12511);
nand U13552 (N_13552,N_12130,N_12251);
xor U13553 (N_13553,N_12231,N_12085);
nand U13554 (N_13554,N_12962,N_12249);
nand U13555 (N_13555,N_12029,N_12955);
or U13556 (N_13556,N_12133,N_12915);
or U13557 (N_13557,N_12732,N_12022);
or U13558 (N_13558,N_12795,N_12191);
nand U13559 (N_13559,N_12609,N_12440);
nor U13560 (N_13560,N_12330,N_12764);
nor U13561 (N_13561,N_12225,N_12679);
nand U13562 (N_13562,N_13178,N_12988);
nor U13563 (N_13563,N_12213,N_13444);
nor U13564 (N_13564,N_12921,N_13367);
nand U13565 (N_13565,N_13442,N_13309);
nand U13566 (N_13566,N_12473,N_12967);
and U13567 (N_13567,N_12433,N_12001);
nor U13568 (N_13568,N_12801,N_13411);
or U13569 (N_13569,N_13018,N_12215);
nor U13570 (N_13570,N_12632,N_13161);
nor U13571 (N_13571,N_12796,N_13420);
nor U13572 (N_13572,N_12405,N_12013);
xor U13573 (N_13573,N_12716,N_13360);
nor U13574 (N_13574,N_12966,N_12254);
nor U13575 (N_13575,N_12835,N_12193);
xor U13576 (N_13576,N_13247,N_12709);
and U13577 (N_13577,N_12222,N_12192);
xnor U13578 (N_13578,N_13374,N_12256);
xor U13579 (N_13579,N_12286,N_13031);
nand U13580 (N_13580,N_12490,N_12513);
and U13581 (N_13581,N_12354,N_12157);
and U13582 (N_13582,N_12940,N_12746);
nor U13583 (N_13583,N_12139,N_12653);
nor U13584 (N_13584,N_12147,N_12025);
or U13585 (N_13585,N_13412,N_12333);
nor U13586 (N_13586,N_12169,N_12236);
nand U13587 (N_13587,N_13257,N_12360);
nand U13588 (N_13588,N_12815,N_13157);
and U13589 (N_13589,N_12898,N_12365);
and U13590 (N_13590,N_12123,N_12682);
and U13591 (N_13591,N_12783,N_13377);
xnor U13592 (N_13592,N_12366,N_12515);
or U13593 (N_13593,N_13017,N_13048);
xnor U13594 (N_13594,N_13400,N_12888);
xnor U13595 (N_13595,N_12153,N_13325);
nor U13596 (N_13596,N_12401,N_12549);
and U13597 (N_13597,N_12922,N_12299);
xor U13598 (N_13598,N_12847,N_12418);
xor U13599 (N_13599,N_12828,N_12787);
nand U13600 (N_13600,N_12229,N_12772);
xnor U13601 (N_13601,N_12011,N_12793);
and U13602 (N_13602,N_13353,N_13106);
nor U13603 (N_13603,N_12259,N_12826);
and U13604 (N_13604,N_12317,N_13192);
and U13605 (N_13605,N_13088,N_12364);
nor U13606 (N_13606,N_12925,N_12019);
nor U13607 (N_13607,N_12372,N_12611);
nor U13608 (N_13608,N_12060,N_13153);
nand U13609 (N_13609,N_12688,N_12356);
and U13610 (N_13610,N_12670,N_12900);
xnor U13611 (N_13611,N_12809,N_12042);
nor U13612 (N_13612,N_12224,N_12076);
nand U13613 (N_13613,N_13401,N_12498);
or U13614 (N_13614,N_13083,N_12751);
or U13615 (N_13615,N_12520,N_12630);
and U13616 (N_13616,N_12590,N_12661);
and U13617 (N_13617,N_12371,N_12004);
nand U13618 (N_13618,N_12641,N_12455);
or U13619 (N_13619,N_12182,N_12876);
xnor U13620 (N_13620,N_13102,N_13396);
or U13621 (N_13621,N_12297,N_12748);
xnor U13622 (N_13622,N_12743,N_12505);
nand U13623 (N_13623,N_13172,N_12577);
xor U13624 (N_13624,N_12383,N_12072);
or U13625 (N_13625,N_13117,N_12015);
and U13626 (N_13626,N_12629,N_13285);
and U13627 (N_13627,N_12063,N_12573);
nor U13628 (N_13628,N_12179,N_12930);
nand U13629 (N_13629,N_13466,N_13149);
nand U13630 (N_13630,N_13040,N_12046);
xor U13631 (N_13631,N_12950,N_12690);
nand U13632 (N_13632,N_13449,N_13008);
nor U13633 (N_13633,N_13345,N_12802);
nor U13634 (N_13634,N_12488,N_13022);
xnor U13635 (N_13635,N_13494,N_12677);
or U13636 (N_13636,N_12817,N_13168);
xor U13637 (N_13637,N_13091,N_12840);
xor U13638 (N_13638,N_13060,N_12627);
and U13639 (N_13639,N_12094,N_12850);
nor U13640 (N_13640,N_12204,N_12245);
nor U13641 (N_13641,N_12453,N_13395);
xnor U13642 (N_13642,N_12662,N_12020);
nor U13643 (N_13643,N_12270,N_12282);
and U13644 (N_13644,N_13333,N_13230);
and U13645 (N_13645,N_12176,N_12706);
and U13646 (N_13646,N_12136,N_12048);
or U13647 (N_13647,N_13484,N_13128);
nand U13648 (N_13648,N_12811,N_12931);
or U13649 (N_13649,N_12854,N_12792);
or U13650 (N_13650,N_13202,N_12212);
xor U13651 (N_13651,N_12412,N_13366);
or U13652 (N_13652,N_13436,N_12477);
and U13653 (N_13653,N_12353,N_12963);
and U13654 (N_13654,N_13093,N_13435);
or U13655 (N_13655,N_12397,N_13077);
or U13656 (N_13656,N_12342,N_12914);
nand U13657 (N_13657,N_13323,N_13020);
xnor U13658 (N_13658,N_12824,N_12102);
nor U13659 (N_13659,N_13355,N_12946);
or U13660 (N_13660,N_13273,N_13417);
or U13661 (N_13661,N_12129,N_12504);
nor U13662 (N_13662,N_12314,N_13201);
nand U13663 (N_13663,N_13012,N_13144);
nand U13664 (N_13664,N_13110,N_12126);
nor U13665 (N_13665,N_12769,N_12866);
or U13666 (N_13666,N_12565,N_12984);
or U13667 (N_13667,N_13124,N_12343);
and U13668 (N_13668,N_12545,N_12118);
or U13669 (N_13669,N_13085,N_12782);
nand U13670 (N_13670,N_12059,N_12460);
or U13671 (N_13671,N_13237,N_12427);
nor U13672 (N_13672,N_13481,N_12429);
nor U13673 (N_13673,N_13164,N_13403);
nor U13674 (N_13674,N_12923,N_12276);
or U13675 (N_13675,N_12444,N_12725);
nor U13676 (N_13676,N_13463,N_13082);
nand U13677 (N_13677,N_12132,N_12587);
nand U13678 (N_13678,N_13131,N_12209);
or U13679 (N_13679,N_12750,N_12869);
and U13680 (N_13680,N_12492,N_12198);
or U13681 (N_13681,N_12537,N_12271);
nor U13682 (N_13682,N_12434,N_12887);
xnor U13683 (N_13683,N_12618,N_12759);
nand U13684 (N_13684,N_13245,N_12973);
nor U13685 (N_13685,N_12516,N_12543);
nor U13686 (N_13686,N_12621,N_12298);
or U13687 (N_13687,N_12935,N_12762);
nor U13688 (N_13688,N_12990,N_13146);
nand U13689 (N_13689,N_12367,N_12425);
nand U13690 (N_13690,N_12886,N_13258);
xor U13691 (N_13691,N_12808,N_12435);
or U13692 (N_13692,N_13475,N_12472);
nor U13693 (N_13693,N_12610,N_12218);
xor U13694 (N_13694,N_13482,N_13072);
nand U13695 (N_13695,N_13014,N_12936);
or U13696 (N_13696,N_12422,N_13147);
xor U13697 (N_13697,N_12622,N_13121);
xnor U13698 (N_13698,N_12100,N_12143);
or U13699 (N_13699,N_12379,N_12997);
nand U13700 (N_13700,N_12985,N_13260);
or U13701 (N_13701,N_13446,N_12834);
nor U13702 (N_13702,N_13169,N_13136);
and U13703 (N_13703,N_12313,N_13308);
nor U13704 (N_13704,N_12778,N_12723);
nor U13705 (N_13705,N_13174,N_13423);
and U13706 (N_13706,N_13339,N_12645);
nand U13707 (N_13707,N_12387,N_12538);
nor U13708 (N_13708,N_13291,N_12838);
xnor U13709 (N_13709,N_12863,N_12323);
and U13710 (N_13710,N_13495,N_13092);
or U13711 (N_13711,N_13456,N_12979);
xor U13712 (N_13712,N_13370,N_12395);
nor U13713 (N_13713,N_12786,N_12572);
nor U13714 (N_13714,N_13324,N_13327);
and U13715 (N_13715,N_12052,N_13050);
and U13716 (N_13716,N_13392,N_12080);
and U13717 (N_13717,N_13068,N_12867);
nand U13718 (N_13718,N_12833,N_12135);
and U13719 (N_13719,N_12109,N_12780);
xor U13720 (N_13720,N_13154,N_13498);
xor U13721 (N_13721,N_12669,N_12305);
nor U13722 (N_13722,N_12026,N_12005);
xor U13723 (N_13723,N_12686,N_12771);
nor U13724 (N_13724,N_12785,N_12602);
xnor U13725 (N_13725,N_12055,N_12635);
and U13726 (N_13726,N_13455,N_13253);
xor U13727 (N_13727,N_12068,N_13344);
or U13728 (N_13728,N_12580,N_13028);
or U13729 (N_13729,N_13242,N_12457);
nor U13730 (N_13730,N_12039,N_12054);
or U13731 (N_13731,N_13490,N_13262);
nor U13732 (N_13732,N_12090,N_12829);
xnor U13733 (N_13733,N_13087,N_13364);
nand U13734 (N_13734,N_12357,N_12494);
nand U13735 (N_13735,N_13239,N_13496);
and U13736 (N_13736,N_12864,N_13122);
nand U13737 (N_13737,N_12875,N_12774);
nor U13738 (N_13738,N_12616,N_12093);
nor U13739 (N_13739,N_12570,N_12252);
nor U13740 (N_13740,N_13249,N_12956);
xnor U13741 (N_13741,N_13470,N_12376);
nand U13742 (N_13742,N_13450,N_12658);
and U13743 (N_13743,N_12167,N_12291);
and U13744 (N_13744,N_13135,N_12766);
xor U13745 (N_13745,N_12197,N_12837);
and U13746 (N_13746,N_13464,N_12668);
nand U13747 (N_13747,N_12431,N_12302);
or U13748 (N_13748,N_12428,N_12241);
or U13749 (N_13749,N_12637,N_13143);
nand U13750 (N_13750,N_12553,N_12937);
and U13751 (N_13751,N_13424,N_12507);
nand U13752 (N_13752,N_13270,N_13447);
nor U13753 (N_13753,N_12087,N_12698);
nor U13754 (N_13754,N_13371,N_13233);
nor U13755 (N_13755,N_12702,N_12972);
or U13756 (N_13756,N_12159,N_13288);
xor U13757 (N_13757,N_12542,N_12033);
nor U13758 (N_13758,N_12959,N_12451);
xnor U13759 (N_13759,N_12908,N_12576);
or U13760 (N_13760,N_12721,N_13032);
nor U13761 (N_13761,N_12238,N_12288);
nand U13762 (N_13762,N_13218,N_12715);
nand U13763 (N_13763,N_12692,N_13338);
nand U13764 (N_13764,N_13362,N_12893);
nor U13765 (N_13765,N_12442,N_12014);
or U13766 (N_13766,N_13382,N_12807);
xor U13767 (N_13767,N_13177,N_13066);
nor U13768 (N_13768,N_12407,N_13497);
nand U13769 (N_13769,N_12430,N_13431);
or U13770 (N_13770,N_13369,N_12034);
xnor U13771 (N_13771,N_12594,N_13408);
nand U13772 (N_13772,N_13105,N_13254);
nor U13773 (N_13773,N_13234,N_12037);
xor U13774 (N_13774,N_13256,N_12518);
nand U13775 (N_13775,N_12882,N_12339);
and U13776 (N_13776,N_13151,N_13196);
or U13777 (N_13777,N_12703,N_12131);
or U13778 (N_13778,N_12281,N_13381);
nor U13779 (N_13779,N_12862,N_13299);
or U13780 (N_13780,N_12304,N_13071);
xor U13781 (N_13781,N_13138,N_12633);
nor U13782 (N_13782,N_13397,N_13252);
nand U13783 (N_13783,N_13264,N_13007);
nor U13784 (N_13784,N_12981,N_12446);
or U13785 (N_13785,N_13289,N_13385);
nor U13786 (N_13786,N_12269,N_12514);
or U13787 (N_13787,N_13329,N_13387);
and U13788 (N_13788,N_12533,N_13489);
nor U13789 (N_13789,N_12903,N_12199);
xor U13790 (N_13790,N_12138,N_12873);
nand U13791 (N_13791,N_13038,N_12227);
or U13792 (N_13792,N_13115,N_12678);
nand U13793 (N_13793,N_12685,N_12894);
nand U13794 (N_13794,N_13021,N_12680);
nor U13795 (N_13795,N_12535,N_12273);
nand U13796 (N_13796,N_13130,N_12600);
and U13797 (N_13797,N_12718,N_13142);
and U13798 (N_13798,N_12813,N_12951);
xnor U13799 (N_13799,N_12308,N_13337);
nand U13800 (N_13800,N_13223,N_12582);
xor U13801 (N_13801,N_12907,N_13140);
nor U13802 (N_13802,N_12789,N_12486);
nand U13803 (N_13803,N_12880,N_12163);
xnor U13804 (N_13804,N_12998,N_12328);
or U13805 (N_13805,N_13134,N_12283);
and U13806 (N_13806,N_12841,N_13046);
xor U13807 (N_13807,N_12221,N_13214);
xor U13808 (N_13808,N_13053,N_12805);
nor U13809 (N_13809,N_12311,N_13426);
nand U13810 (N_13810,N_12158,N_12174);
nand U13811 (N_13811,N_13363,N_12247);
xor U13812 (N_13812,N_12699,N_13292);
nand U13813 (N_13813,N_12563,N_12591);
and U13814 (N_13814,N_12468,N_12745);
nor U13815 (N_13815,N_12768,N_13492);
xnor U13816 (N_13816,N_12681,N_12760);
nand U13817 (N_13817,N_12326,N_12183);
xor U13818 (N_13818,N_12905,N_13210);
and U13819 (N_13819,N_12369,N_12050);
and U13820 (N_13820,N_12825,N_12539);
nand U13821 (N_13821,N_12024,N_12932);
nand U13822 (N_13822,N_12464,N_12177);
xnor U13823 (N_13823,N_13283,N_12082);
xnor U13824 (N_13824,N_13199,N_12079);
and U13825 (N_13825,N_12917,N_13306);
xnor U13826 (N_13826,N_12219,N_13343);
xor U13827 (N_13827,N_13269,N_13261);
or U13828 (N_13828,N_12250,N_13491);
nor U13829 (N_13829,N_12557,N_13359);
nand U13830 (N_13830,N_12858,N_12099);
or U13831 (N_13831,N_12375,N_12307);
xnor U13832 (N_13832,N_12711,N_12470);
xnor U13833 (N_13833,N_12237,N_12896);
or U13834 (N_13834,N_13413,N_12977);
xor U13835 (N_13835,N_12414,N_12673);
or U13836 (N_13836,N_12607,N_13259);
xnor U13837 (N_13837,N_12415,N_12560);
and U13838 (N_13838,N_12010,N_12426);
nand U13839 (N_13839,N_13373,N_13055);
and U13840 (N_13840,N_13155,N_12744);
or U13841 (N_13841,N_12340,N_12089);
nand U13842 (N_13842,N_12027,N_12722);
and U13843 (N_13843,N_12978,N_12909);
and U13844 (N_13844,N_12810,N_12848);
or U13845 (N_13845,N_12644,N_12649);
nor U13846 (N_13846,N_12740,N_13265);
nand U13847 (N_13847,N_12230,N_12704);
or U13848 (N_13848,N_12280,N_13064);
nor U13849 (N_13849,N_12113,N_12755);
or U13850 (N_13850,N_13282,N_12599);
nand U13851 (N_13851,N_12551,N_12466);
and U13852 (N_13852,N_13439,N_13175);
xor U13853 (N_13853,N_12713,N_12140);
xnor U13854 (N_13854,N_13297,N_12620);
xor U13855 (N_13855,N_12053,N_12788);
nand U13856 (N_13856,N_12106,N_12916);
nor U13857 (N_13857,N_12884,N_13099);
xor U13858 (N_13858,N_12613,N_12812);
nor U13859 (N_13859,N_13109,N_13181);
or U13860 (N_13860,N_12295,N_12974);
xor U13861 (N_13861,N_12203,N_12399);
xnor U13862 (N_13862,N_12593,N_13216);
nand U13863 (N_13863,N_12729,N_12986);
nand U13864 (N_13864,N_13347,N_12449);
and U13865 (N_13865,N_12261,N_13284);
and U13866 (N_13866,N_12021,N_13281);
or U13867 (N_13867,N_12581,N_12156);
xnor U13868 (N_13868,N_13469,N_13335);
nand U13869 (N_13869,N_12349,N_13378);
or U13870 (N_13870,N_12853,N_12400);
nand U13871 (N_13871,N_12168,N_12861);
and U13872 (N_13872,N_13386,N_13326);
or U13873 (N_13873,N_12043,N_13019);
nor U13874 (N_13874,N_12693,N_12883);
and U13875 (N_13875,N_12064,N_13126);
nand U13876 (N_13876,N_13402,N_13244);
xnor U13877 (N_13877,N_12953,N_13079);
nand U13878 (N_13878,N_12394,N_12592);
and U13879 (N_13879,N_12125,N_13388);
and U13880 (N_13880,N_12120,N_12517);
xor U13881 (N_13881,N_13485,N_12881);
nor U13882 (N_13882,N_13451,N_12246);
and U13883 (N_13883,N_12651,N_12028);
or U13884 (N_13884,N_13133,N_12614);
nor U13885 (N_13885,N_12569,N_12934);
and U13886 (N_13886,N_12958,N_12499);
or U13887 (N_13887,N_12008,N_13465);
or U13888 (N_13888,N_13272,N_12512);
and U13889 (N_13889,N_12728,N_12501);
and U13890 (N_13890,N_12278,N_13176);
or U13891 (N_13891,N_12827,N_12944);
or U13892 (N_13892,N_13204,N_13024);
or U13893 (N_13893,N_13225,N_12776);
nor U13894 (N_13894,N_12660,N_12552);
or U13895 (N_13895,N_12724,N_13390);
nor U13896 (N_13896,N_13453,N_12370);
and U13897 (N_13897,N_13129,N_12982);
nand U13898 (N_13898,N_12194,N_12992);
nand U13899 (N_13899,N_13215,N_12717);
nor U13900 (N_13900,N_12154,N_12462);
and U13901 (N_13901,N_12814,N_13432);
xor U13902 (N_13902,N_13051,N_12579);
and U13903 (N_13903,N_12567,N_12180);
xor U13904 (N_13904,N_12189,N_12104);
and U13905 (N_13905,N_12761,N_13059);
nor U13906 (N_13906,N_12105,N_12701);
xnor U13907 (N_13907,N_12939,N_13222);
nor U13908 (N_13908,N_12228,N_13452);
xor U13909 (N_13909,N_13278,N_13219);
and U13910 (N_13910,N_12438,N_12571);
xor U13911 (N_13911,N_12240,N_13195);
and U13912 (N_13912,N_12901,N_13054);
nor U13913 (N_13913,N_13389,N_13043);
nand U13914 (N_13914,N_12737,N_12361);
nand U13915 (N_13915,N_12519,N_12957);
and U13916 (N_13916,N_12469,N_12478);
or U13917 (N_13917,N_12976,N_12122);
xnor U13918 (N_13918,N_13352,N_13468);
nor U13919 (N_13919,N_13312,N_13049);
xnor U13920 (N_13920,N_12964,N_12081);
nor U13921 (N_13921,N_12720,N_12355);
nand U13922 (N_13922,N_12458,N_12320);
nor U13923 (N_13923,N_12484,N_13226);
nand U13924 (N_13924,N_13041,N_12487);
and U13925 (N_13925,N_12534,N_12821);
and U13926 (N_13926,N_12244,N_13015);
xor U13927 (N_13927,N_12991,N_12057);
and U13928 (N_13928,N_12146,N_12736);
nor U13929 (N_13929,N_13428,N_12851);
nor U13930 (N_13930,N_12712,N_13029);
and U13931 (N_13931,N_13074,N_12095);
nor U13932 (N_13932,N_13203,N_12258);
xor U13933 (N_13933,N_13346,N_12348);
xor U13934 (N_13934,N_13348,N_12172);
and U13935 (N_13935,N_12860,N_13217);
nor U13936 (N_13936,N_12753,N_12767);
nand U13937 (N_13937,N_13034,N_13189);
xor U13938 (N_13938,N_13073,N_13094);
and U13939 (N_13939,N_12798,N_12648);
nand U13940 (N_13940,N_12344,N_12619);
and U13941 (N_13941,N_12904,N_12527);
or U13942 (N_13942,N_13350,N_13440);
nand U13943 (N_13943,N_12012,N_12846);
and U13944 (N_13944,N_12758,N_12474);
and U13945 (N_13945,N_13294,N_13045);
and U13946 (N_13946,N_12960,N_12877);
xor U13947 (N_13947,N_12735,N_12918);
nor U13948 (N_13948,N_13036,N_13295);
xor U13949 (N_13949,N_12970,N_12954);
xnor U13950 (N_13950,N_13044,N_12016);
nor U13951 (N_13951,N_13016,N_13243);
nand U13952 (N_13952,N_12248,N_12303);
nor U13953 (N_13953,N_13187,N_13061);
and U13954 (N_13954,N_12352,N_12708);
nor U13955 (N_13955,N_12938,N_13137);
xnor U13956 (N_13956,N_12719,N_12994);
nor U13957 (N_13957,N_12754,N_13321);
and U13958 (N_13958,N_12503,N_12657);
and U13959 (N_13959,N_13477,N_13070);
or U13960 (N_13960,N_12656,N_12843);
xor U13961 (N_13961,N_12253,N_13290);
or U13962 (N_13962,N_12942,N_12409);
nand U13963 (N_13963,N_12987,N_12301);
and U13964 (N_13964,N_13221,N_12526);
and U13965 (N_13965,N_12742,N_12707);
or U13966 (N_13966,N_13002,N_12277);
or U13967 (N_13967,N_12456,N_12684);
and U13968 (N_13968,N_13065,N_12077);
and U13969 (N_13969,N_13351,N_12439);
xor U13970 (N_13970,N_12561,N_12111);
and U13971 (N_13971,N_13445,N_12003);
nand U13972 (N_13972,N_13057,N_12115);
xnor U13973 (N_13973,N_13042,N_12624);
nand U13974 (N_13974,N_12522,N_13058);
nand U13975 (N_13975,N_13004,N_12265);
and U13976 (N_13976,N_12927,N_13000);
nand U13977 (N_13977,N_12804,N_12009);
nor U13978 (N_13978,N_12906,N_12752);
or U13979 (N_13979,N_12373,N_13319);
xnor U13980 (N_13980,N_12214,N_12264);
or U13981 (N_13981,N_13441,N_12683);
xnor U13982 (N_13982,N_12341,N_13037);
xnor U13983 (N_13983,N_12351,N_12818);
and U13984 (N_13984,N_12235,N_13255);
or U13985 (N_13985,N_13100,N_13185);
nand U13986 (N_13986,N_13098,N_12675);
and U13987 (N_13987,N_12643,N_12445);
nand U13988 (N_13988,N_13274,N_12312);
or U13989 (N_13989,N_13227,N_12849);
and U13990 (N_13990,N_12646,N_12070);
xnor U13991 (N_13991,N_12413,N_12450);
nand U13992 (N_13992,N_12741,N_12625);
or U13993 (N_13993,N_12574,N_12223);
nor U13994 (N_13994,N_12318,N_12398);
xor U13995 (N_13995,N_12233,N_12447);
xor U13996 (N_13996,N_13033,N_13145);
xnor U13997 (N_13997,N_12206,N_12667);
nor U13998 (N_13998,N_13429,N_12443);
or U13999 (N_13999,N_12747,N_12995);
xnor U14000 (N_14000,N_12047,N_13302);
and U14001 (N_14001,N_13368,N_12292);
or U14002 (N_14002,N_13123,N_13310);
and U14003 (N_14003,N_13166,N_12949);
and U14004 (N_14004,N_12733,N_12870);
xnor U14005 (N_14005,N_12506,N_12289);
xnor U14006 (N_14006,N_13159,N_12666);
or U14007 (N_14007,N_12128,N_12272);
and U14008 (N_14008,N_12556,N_12731);
xnor U14009 (N_14009,N_12359,N_12671);
and U14010 (N_14010,N_12336,N_12996);
nor U14011 (N_14011,N_12842,N_12293);
nor U14012 (N_14012,N_12380,N_12097);
or U14013 (N_14013,N_12421,N_12411);
and U14014 (N_14014,N_13127,N_13427);
and U14015 (N_14015,N_13084,N_12239);
and U14016 (N_14016,N_12393,N_12152);
or U14017 (N_14017,N_12309,N_13454);
and U14018 (N_14018,N_12528,N_12142);
nor U14019 (N_14019,N_12926,N_13416);
nand U14020 (N_14020,N_12555,N_13006);
nor U14021 (N_14021,N_12083,N_13275);
and U14022 (N_14022,N_13235,N_13191);
nor U14023 (N_14023,N_13407,N_12695);
nor U14024 (N_14024,N_12773,N_12051);
and U14025 (N_14025,N_12166,N_12822);
or U14026 (N_14026,N_13173,N_13391);
or U14027 (N_14027,N_13206,N_12529);
nor U14028 (N_14028,N_12067,N_12605);
nand U14029 (N_14029,N_12200,N_12103);
nand U14030 (N_14030,N_12615,N_12868);
nor U14031 (N_14031,N_12017,N_13476);
xnor U14032 (N_14032,N_13023,N_13479);
xor U14033 (N_14033,N_13287,N_13314);
or U14034 (N_14034,N_12612,N_13125);
nor U14035 (N_14035,N_13080,N_12588);
and U14036 (N_14036,N_12536,N_13213);
or U14037 (N_14037,N_12710,N_12639);
xnor U14038 (N_14038,N_12820,N_13304);
nor U14039 (N_14039,N_13459,N_12274);
or U14040 (N_14040,N_13116,N_12403);
or U14041 (N_14041,N_12608,N_12124);
or U14042 (N_14042,N_13220,N_13076);
or U14043 (N_14043,N_12816,N_12041);
xnor U14044 (N_14044,N_13340,N_13114);
nand U14045 (N_14045,N_12601,N_13334);
nand U14046 (N_14046,N_12830,N_12208);
or U14047 (N_14047,N_12654,N_13251);
nand U14048 (N_14048,N_12329,N_12475);
nand U14049 (N_14049,N_12859,N_13316);
nor U14050 (N_14050,N_12562,N_13003);
and U14051 (N_14051,N_12623,N_13376);
or U14052 (N_14052,N_13160,N_12040);
nor U14053 (N_14053,N_12584,N_12030);
xor U14054 (N_14054,N_12416,N_12546);
and U14055 (N_14055,N_12112,N_12390);
nand U14056 (N_14056,N_12471,N_13461);
nand U14057 (N_14057,N_12929,N_12170);
xnor U14058 (N_14058,N_13167,N_13328);
xnor U14059 (N_14059,N_12652,N_12943);
or U14060 (N_14060,N_12290,N_12459);
xor U14061 (N_14061,N_12948,N_12756);
or U14062 (N_14062,N_13349,N_13322);
xor U14063 (N_14063,N_13425,N_12777);
xnor U14064 (N_14064,N_13163,N_12993);
or U14065 (N_14065,N_12910,N_12216);
and U14066 (N_14066,N_12049,N_13394);
and U14067 (N_14067,N_12631,N_13471);
or U14068 (N_14068,N_12201,N_12144);
nand U14069 (N_14069,N_13358,N_13434);
xor U14070 (N_14070,N_12547,N_12700);
xnor U14071 (N_14071,N_13342,N_12396);
nand U14072 (N_14072,N_13212,N_13300);
nand U14073 (N_14073,N_13303,N_12696);
nand U14074 (N_14074,N_12554,N_13296);
xor U14075 (N_14075,N_12879,N_13081);
nor U14076 (N_14076,N_12186,N_12098);
or U14077 (N_14077,N_13414,N_12091);
nor U14078 (N_14078,N_12674,N_12483);
or U14079 (N_14079,N_13380,N_12044);
or U14080 (N_14080,N_12368,N_12550);
xnor U14081 (N_14081,N_12045,N_13119);
or U14082 (N_14082,N_13276,N_12331);
xnor U14083 (N_14083,N_12730,N_13238);
nand U14084 (N_14084,N_12548,N_12074);
and U14085 (N_14085,N_12790,N_12603);
nor U14086 (N_14086,N_13067,N_12928);
or U14087 (N_14087,N_12595,N_13165);
nand U14088 (N_14088,N_12763,N_12589);
or U14089 (N_14089,N_12965,N_12891);
nor U14090 (N_14090,N_12392,N_12073);
xnor U14091 (N_14091,N_12007,N_12689);
nor U14092 (N_14092,N_13205,N_12636);
xor U14093 (N_14093,N_12687,N_12497);
and U14094 (N_14094,N_13062,N_12220);
and U14095 (N_14095,N_12691,N_12521);
nand U14096 (N_14096,N_12101,N_13467);
nand U14097 (N_14097,N_12389,N_13356);
nand U14098 (N_14098,N_13132,N_13493);
and U14099 (N_14099,N_13487,N_13075);
xor U14100 (N_14100,N_13186,N_12606);
nand U14101 (N_14101,N_12749,N_13419);
nor U14102 (N_14102,N_13486,N_13182);
and U14103 (N_14103,N_12694,N_12316);
or U14104 (N_14104,N_12941,N_12374);
xnor U14105 (N_14105,N_12108,N_12217);
nor U14106 (N_14106,N_12437,N_12496);
xnor U14107 (N_14107,N_13383,N_13478);
nand U14108 (N_14108,N_12770,N_12482);
nand U14109 (N_14109,N_13311,N_12127);
xnor U14110 (N_14110,N_13107,N_12481);
and U14111 (N_14111,N_13250,N_13280);
xnor U14112 (N_14112,N_12500,N_12531);
or U14113 (N_14113,N_13170,N_13404);
xor U14114 (N_14114,N_12969,N_13228);
nand U14115 (N_14115,N_12121,N_12448);
nand U14116 (N_14116,N_12260,N_12794);
xnor U14117 (N_14117,N_12114,N_12347);
and U14118 (N_14118,N_13318,N_12844);
or U14119 (N_14119,N_13150,N_13001);
or U14120 (N_14120,N_13399,N_12285);
xnor U14121 (N_14121,N_12294,N_12058);
nor U14122 (N_14122,N_13005,N_13266);
and U14123 (N_14123,N_13056,N_12065);
nand U14124 (N_14124,N_12173,N_12461);
and U14125 (N_14125,N_12319,N_13305);
xor U14126 (N_14126,N_12596,N_12018);
or U14127 (N_14127,N_13232,N_12465);
nor U14128 (N_14128,N_12210,N_12775);
nand U14129 (N_14129,N_12647,N_13448);
and U14130 (N_14130,N_12855,N_12306);
and U14131 (N_14131,N_12911,N_12268);
xnor U14132 (N_14132,N_12150,N_13171);
nor U14133 (N_14133,N_12791,N_12897);
xnor U14134 (N_14134,N_12493,N_12441);
or U14135 (N_14135,N_12338,N_12634);
nand U14136 (N_14136,N_12525,N_13156);
nand U14137 (N_14137,N_12524,N_13047);
nand U14138 (N_14138,N_13457,N_13483);
nand U14139 (N_14139,N_12006,N_12463);
or U14140 (N_14140,N_13111,N_12586);
nor U14141 (N_14141,N_12162,N_13330);
nor U14142 (N_14142,N_12000,N_12384);
or U14143 (N_14143,N_12296,N_13301);
and U14144 (N_14144,N_12161,N_12510);
or U14145 (N_14145,N_12196,N_13458);
xnor U14146 (N_14146,N_12664,N_13097);
and U14147 (N_14147,N_12381,N_13438);
nor U14148 (N_14148,N_13013,N_13179);
or U14149 (N_14149,N_12137,N_13263);
nor U14150 (N_14150,N_13277,N_13499);
or U14151 (N_14151,N_12149,N_12485);
xnor U14152 (N_14152,N_12857,N_12575);
or U14153 (N_14153,N_13190,N_12727);
and U14154 (N_14154,N_12784,N_12989);
xnor U14155 (N_14155,N_12432,N_13025);
xor U14156 (N_14156,N_13271,N_12920);
or U14157 (N_14157,N_12061,N_12420);
xor U14158 (N_14158,N_12913,N_12738);
xor U14159 (N_14159,N_12714,N_12509);
or U14160 (N_14160,N_12062,N_13207);
and U14161 (N_14161,N_13320,N_12148);
nor U14162 (N_14162,N_12035,N_12335);
and U14163 (N_14163,N_12803,N_12327);
or U14164 (N_14164,N_13011,N_13354);
xor U14165 (N_14165,N_13248,N_13193);
xor U14166 (N_14166,N_13240,N_12300);
xnor U14167 (N_14167,N_12878,N_12267);
nor U14168 (N_14168,N_12185,N_12806);
nand U14169 (N_14169,N_12454,N_12779);
xnor U14170 (N_14170,N_12362,N_12160);
nor U14171 (N_14171,N_12410,N_12889);
nor U14172 (N_14172,N_12066,N_13361);
nand U14173 (N_14173,N_12096,N_13293);
and U14174 (N_14174,N_13113,N_12408);
or U14175 (N_14175,N_12284,N_12255);
or U14176 (N_14176,N_13197,N_12739);
and U14177 (N_14177,N_13162,N_12665);
nand U14178 (N_14178,N_12597,N_12852);
nand U14179 (N_14179,N_12190,N_12476);
nand U14180 (N_14180,N_12924,N_12819);
nor U14181 (N_14181,N_12404,N_12195);
or U14182 (N_14182,N_12032,N_13009);
nand U14183 (N_14183,N_12765,N_12971);
nor U14184 (N_14184,N_13317,N_12086);
and U14185 (N_14185,N_12391,N_13241);
xor U14186 (N_14186,N_12350,N_13188);
nand U14187 (N_14187,N_12263,N_12202);
nand U14188 (N_14188,N_12541,N_13357);
nor U14189 (N_14189,N_12856,N_13198);
and U14190 (N_14190,N_12155,N_12480);
and U14191 (N_14191,N_12961,N_13103);
nor U14192 (N_14192,N_12402,N_12178);
and U14193 (N_14193,N_13052,N_12558);
nand U14194 (N_14194,N_12363,N_12628);
nand U14195 (N_14195,N_13315,N_12031);
nor U14196 (N_14196,N_13313,N_12945);
nand U14197 (N_14197,N_12865,N_13152);
xnor U14198 (N_14198,N_12287,N_13421);
nor U14199 (N_14199,N_12663,N_13231);
or U14200 (N_14200,N_12578,N_13336);
and U14201 (N_14201,N_12386,N_12705);
nand U14202 (N_14202,N_12232,N_13108);
and U14203 (N_14203,N_13341,N_12321);
or U14204 (N_14204,N_12234,N_13379);
and U14205 (N_14205,N_12243,N_12325);
nor U14206 (N_14206,N_13331,N_12188);
xor U14207 (N_14207,N_12598,N_12655);
nand U14208 (N_14208,N_13090,N_12566);
xnor U14209 (N_14209,N_12069,N_13398);
nand U14210 (N_14210,N_13236,N_12638);
nor U14211 (N_14211,N_13200,N_12650);
nor U14212 (N_14212,N_13141,N_13430);
nand U14213 (N_14213,N_12419,N_12164);
and U14214 (N_14214,N_12088,N_12980);
or U14215 (N_14215,N_13078,N_12832);
xor U14216 (N_14216,N_12823,N_12672);
and U14217 (N_14217,N_12184,N_12968);
and U14218 (N_14218,N_12322,N_12892);
xor U14219 (N_14219,N_13298,N_12899);
nand U14220 (N_14220,N_13246,N_12452);
nor U14221 (N_14221,N_13183,N_13418);
nand U14222 (N_14222,N_12092,N_13462);
nand U14223 (N_14223,N_12038,N_13158);
nor U14224 (N_14224,N_13480,N_13410);
xor U14225 (N_14225,N_12676,N_12983);
and U14226 (N_14226,N_12604,N_12871);
nand U14227 (N_14227,N_12495,N_12564);
nor U14228 (N_14228,N_12002,N_12617);
nor U14229 (N_14229,N_13474,N_13332);
and U14230 (N_14230,N_13406,N_13422);
xor U14231 (N_14231,N_13229,N_13488);
xor U14232 (N_14232,N_12117,N_13209);
or U14233 (N_14233,N_12872,N_12423);
nand U14234 (N_14234,N_12226,N_13063);
xor U14235 (N_14235,N_13433,N_12642);
nor U14236 (N_14236,N_12324,N_12141);
xor U14237 (N_14237,N_13095,N_12585);
nor U14238 (N_14238,N_13101,N_12332);
and U14239 (N_14239,N_12800,N_13286);
nor U14240 (N_14240,N_13089,N_13096);
or U14241 (N_14241,N_13393,N_12145);
xor U14242 (N_14242,N_13208,N_12378);
and U14243 (N_14243,N_12912,N_12242);
nand U14244 (N_14244,N_13405,N_12134);
xnor U14245 (N_14245,N_12489,N_12757);
or U14246 (N_14246,N_13307,N_12211);
nor U14247 (N_14247,N_13415,N_12975);
xor U14248 (N_14248,N_12845,N_12310);
nand U14249 (N_14249,N_12078,N_13104);
and U14250 (N_14250,N_12844,N_13443);
xor U14251 (N_14251,N_13213,N_13487);
nand U14252 (N_14252,N_12608,N_13327);
nor U14253 (N_14253,N_13190,N_13079);
xnor U14254 (N_14254,N_12033,N_12050);
xnor U14255 (N_14255,N_12912,N_12829);
nor U14256 (N_14256,N_13483,N_12683);
and U14257 (N_14257,N_13230,N_12370);
nand U14258 (N_14258,N_12166,N_12177);
xnor U14259 (N_14259,N_12172,N_12263);
nand U14260 (N_14260,N_13209,N_12833);
nand U14261 (N_14261,N_13235,N_13117);
and U14262 (N_14262,N_12793,N_13030);
and U14263 (N_14263,N_12575,N_12033);
xnor U14264 (N_14264,N_13297,N_13115);
or U14265 (N_14265,N_12039,N_12204);
nand U14266 (N_14266,N_12948,N_12408);
xor U14267 (N_14267,N_12163,N_12806);
xnor U14268 (N_14268,N_13488,N_12679);
or U14269 (N_14269,N_12887,N_12839);
nand U14270 (N_14270,N_13405,N_13359);
or U14271 (N_14271,N_13089,N_12748);
nand U14272 (N_14272,N_13057,N_12417);
nor U14273 (N_14273,N_12736,N_12009);
xor U14274 (N_14274,N_12175,N_12341);
xor U14275 (N_14275,N_12868,N_13076);
nor U14276 (N_14276,N_13316,N_12323);
and U14277 (N_14277,N_12230,N_12574);
or U14278 (N_14278,N_12738,N_12718);
nand U14279 (N_14279,N_12309,N_13458);
nand U14280 (N_14280,N_13498,N_12327);
nand U14281 (N_14281,N_13391,N_13365);
nor U14282 (N_14282,N_13303,N_12880);
or U14283 (N_14283,N_13100,N_12127);
nor U14284 (N_14284,N_13389,N_13206);
or U14285 (N_14285,N_13187,N_12678);
nand U14286 (N_14286,N_12246,N_12855);
nor U14287 (N_14287,N_12091,N_12126);
nor U14288 (N_14288,N_13130,N_13021);
nor U14289 (N_14289,N_12276,N_13390);
and U14290 (N_14290,N_12265,N_12741);
xnor U14291 (N_14291,N_13366,N_12301);
and U14292 (N_14292,N_12243,N_12641);
nor U14293 (N_14293,N_12146,N_13019);
nand U14294 (N_14294,N_13112,N_12976);
or U14295 (N_14295,N_13091,N_12682);
and U14296 (N_14296,N_12162,N_12210);
nand U14297 (N_14297,N_13376,N_12344);
and U14298 (N_14298,N_12349,N_12269);
and U14299 (N_14299,N_12642,N_12517);
and U14300 (N_14300,N_12868,N_13186);
or U14301 (N_14301,N_13309,N_12479);
or U14302 (N_14302,N_12488,N_13364);
or U14303 (N_14303,N_13296,N_13171);
xor U14304 (N_14304,N_13296,N_13238);
or U14305 (N_14305,N_12627,N_12992);
nand U14306 (N_14306,N_12545,N_12616);
or U14307 (N_14307,N_12717,N_13470);
nand U14308 (N_14308,N_12920,N_12333);
or U14309 (N_14309,N_12178,N_12691);
nor U14310 (N_14310,N_12500,N_12968);
or U14311 (N_14311,N_13207,N_13270);
and U14312 (N_14312,N_12753,N_12171);
and U14313 (N_14313,N_12180,N_12321);
xor U14314 (N_14314,N_12230,N_12886);
and U14315 (N_14315,N_12865,N_13240);
or U14316 (N_14316,N_12448,N_13447);
and U14317 (N_14317,N_12098,N_12390);
nor U14318 (N_14318,N_12709,N_12167);
nor U14319 (N_14319,N_12784,N_12469);
or U14320 (N_14320,N_13057,N_12913);
or U14321 (N_14321,N_12865,N_12509);
xor U14322 (N_14322,N_13044,N_12422);
xor U14323 (N_14323,N_12325,N_13168);
nand U14324 (N_14324,N_13482,N_13472);
nor U14325 (N_14325,N_12282,N_12604);
nor U14326 (N_14326,N_13333,N_12922);
and U14327 (N_14327,N_12433,N_13369);
or U14328 (N_14328,N_13269,N_12338);
nand U14329 (N_14329,N_12014,N_12060);
xor U14330 (N_14330,N_12161,N_13087);
nor U14331 (N_14331,N_13450,N_13347);
nor U14332 (N_14332,N_12898,N_12124);
and U14333 (N_14333,N_13392,N_12848);
xnor U14334 (N_14334,N_13459,N_13303);
xor U14335 (N_14335,N_12312,N_12691);
or U14336 (N_14336,N_12131,N_12925);
nor U14337 (N_14337,N_12758,N_12204);
or U14338 (N_14338,N_12195,N_13131);
nand U14339 (N_14339,N_12677,N_12804);
xnor U14340 (N_14340,N_12953,N_12725);
and U14341 (N_14341,N_13386,N_13044);
or U14342 (N_14342,N_13039,N_13116);
and U14343 (N_14343,N_12824,N_12410);
or U14344 (N_14344,N_12333,N_12991);
or U14345 (N_14345,N_12229,N_12405);
xnor U14346 (N_14346,N_12551,N_12896);
or U14347 (N_14347,N_13238,N_12234);
nor U14348 (N_14348,N_12556,N_13384);
or U14349 (N_14349,N_13462,N_13278);
xnor U14350 (N_14350,N_13250,N_13482);
or U14351 (N_14351,N_13313,N_13149);
xor U14352 (N_14352,N_12151,N_12747);
and U14353 (N_14353,N_13166,N_12048);
or U14354 (N_14354,N_12341,N_13073);
xnor U14355 (N_14355,N_12889,N_12624);
nor U14356 (N_14356,N_13114,N_13283);
or U14357 (N_14357,N_12424,N_12236);
nor U14358 (N_14358,N_13422,N_13211);
or U14359 (N_14359,N_12065,N_12897);
xnor U14360 (N_14360,N_12582,N_12090);
and U14361 (N_14361,N_12880,N_12775);
xnor U14362 (N_14362,N_13148,N_13111);
or U14363 (N_14363,N_12003,N_12622);
nand U14364 (N_14364,N_12212,N_12438);
nand U14365 (N_14365,N_12021,N_13309);
nor U14366 (N_14366,N_13361,N_12783);
nand U14367 (N_14367,N_13472,N_12349);
nor U14368 (N_14368,N_13405,N_12669);
xor U14369 (N_14369,N_12663,N_13091);
xor U14370 (N_14370,N_13256,N_12447);
nor U14371 (N_14371,N_12782,N_12294);
nand U14372 (N_14372,N_12634,N_13333);
nor U14373 (N_14373,N_12432,N_12999);
and U14374 (N_14374,N_12803,N_12308);
xnor U14375 (N_14375,N_13025,N_12122);
xor U14376 (N_14376,N_12127,N_12473);
nor U14377 (N_14377,N_13072,N_13480);
or U14378 (N_14378,N_12749,N_13069);
nor U14379 (N_14379,N_12908,N_13191);
and U14380 (N_14380,N_13299,N_12665);
nor U14381 (N_14381,N_12635,N_12228);
and U14382 (N_14382,N_12691,N_12260);
nand U14383 (N_14383,N_12480,N_13211);
nor U14384 (N_14384,N_12064,N_12929);
or U14385 (N_14385,N_13058,N_12864);
or U14386 (N_14386,N_13265,N_12298);
and U14387 (N_14387,N_12887,N_12038);
xor U14388 (N_14388,N_12905,N_13274);
nor U14389 (N_14389,N_13286,N_12908);
nand U14390 (N_14390,N_12816,N_13237);
nor U14391 (N_14391,N_12407,N_12303);
nor U14392 (N_14392,N_12620,N_12481);
and U14393 (N_14393,N_12002,N_13067);
nand U14394 (N_14394,N_13345,N_12748);
xor U14395 (N_14395,N_12825,N_12531);
xnor U14396 (N_14396,N_13100,N_12955);
and U14397 (N_14397,N_13473,N_12966);
or U14398 (N_14398,N_12777,N_13288);
or U14399 (N_14399,N_12377,N_12801);
nor U14400 (N_14400,N_13298,N_13056);
nand U14401 (N_14401,N_12399,N_12278);
nor U14402 (N_14402,N_13302,N_13069);
or U14403 (N_14403,N_12276,N_12955);
or U14404 (N_14404,N_12393,N_12253);
and U14405 (N_14405,N_12786,N_12215);
and U14406 (N_14406,N_12927,N_13125);
nand U14407 (N_14407,N_13031,N_12745);
and U14408 (N_14408,N_13210,N_12006);
nor U14409 (N_14409,N_12553,N_13380);
nand U14410 (N_14410,N_13163,N_12076);
and U14411 (N_14411,N_13049,N_13134);
nor U14412 (N_14412,N_13222,N_12285);
or U14413 (N_14413,N_12111,N_12566);
nand U14414 (N_14414,N_12749,N_13291);
and U14415 (N_14415,N_13481,N_12974);
or U14416 (N_14416,N_12431,N_12264);
nor U14417 (N_14417,N_12087,N_12393);
xor U14418 (N_14418,N_12876,N_12729);
or U14419 (N_14419,N_13005,N_13295);
and U14420 (N_14420,N_13286,N_12368);
nor U14421 (N_14421,N_12873,N_12143);
nor U14422 (N_14422,N_12814,N_12956);
nor U14423 (N_14423,N_12296,N_12324);
and U14424 (N_14424,N_12790,N_13384);
or U14425 (N_14425,N_13221,N_12860);
and U14426 (N_14426,N_12145,N_13107);
nand U14427 (N_14427,N_13245,N_12540);
or U14428 (N_14428,N_12815,N_13395);
or U14429 (N_14429,N_13123,N_12458);
and U14430 (N_14430,N_12608,N_12598);
nand U14431 (N_14431,N_13228,N_12423);
and U14432 (N_14432,N_13302,N_12061);
nand U14433 (N_14433,N_12960,N_12242);
nor U14434 (N_14434,N_12165,N_12308);
nor U14435 (N_14435,N_13420,N_13447);
nor U14436 (N_14436,N_12195,N_12935);
xor U14437 (N_14437,N_12918,N_12269);
or U14438 (N_14438,N_12199,N_12052);
nor U14439 (N_14439,N_13018,N_13334);
nand U14440 (N_14440,N_13062,N_12903);
nand U14441 (N_14441,N_13499,N_13236);
nand U14442 (N_14442,N_12479,N_12663);
nand U14443 (N_14443,N_12934,N_12410);
nor U14444 (N_14444,N_12235,N_13072);
or U14445 (N_14445,N_12760,N_13480);
or U14446 (N_14446,N_13127,N_12121);
nand U14447 (N_14447,N_13444,N_13479);
or U14448 (N_14448,N_12255,N_12105);
nor U14449 (N_14449,N_12004,N_12892);
or U14450 (N_14450,N_12640,N_12052);
or U14451 (N_14451,N_12591,N_12704);
nor U14452 (N_14452,N_12458,N_12346);
nor U14453 (N_14453,N_12030,N_12573);
and U14454 (N_14454,N_13343,N_12785);
xor U14455 (N_14455,N_13365,N_12675);
nor U14456 (N_14456,N_12581,N_12764);
nor U14457 (N_14457,N_13125,N_13486);
and U14458 (N_14458,N_12918,N_13156);
or U14459 (N_14459,N_12365,N_12433);
nand U14460 (N_14460,N_12525,N_12622);
xor U14461 (N_14461,N_12598,N_12922);
nand U14462 (N_14462,N_13480,N_13323);
xnor U14463 (N_14463,N_12210,N_12788);
xor U14464 (N_14464,N_12348,N_12644);
or U14465 (N_14465,N_13382,N_12626);
nor U14466 (N_14466,N_12677,N_12052);
nand U14467 (N_14467,N_12005,N_12441);
nand U14468 (N_14468,N_12183,N_12232);
nand U14469 (N_14469,N_12751,N_13306);
nor U14470 (N_14470,N_12120,N_13196);
and U14471 (N_14471,N_13078,N_12490);
and U14472 (N_14472,N_12002,N_12748);
and U14473 (N_14473,N_13395,N_13398);
nor U14474 (N_14474,N_12787,N_12437);
nand U14475 (N_14475,N_13115,N_12168);
xor U14476 (N_14476,N_13309,N_13003);
nand U14477 (N_14477,N_13498,N_12329);
and U14478 (N_14478,N_12376,N_12375);
and U14479 (N_14479,N_12487,N_13410);
nor U14480 (N_14480,N_13367,N_13138);
nor U14481 (N_14481,N_12927,N_12949);
nor U14482 (N_14482,N_12768,N_12532);
nor U14483 (N_14483,N_12147,N_12894);
nand U14484 (N_14484,N_12568,N_12130);
xor U14485 (N_14485,N_13476,N_12078);
nor U14486 (N_14486,N_13177,N_13362);
xnor U14487 (N_14487,N_12358,N_13138);
or U14488 (N_14488,N_13452,N_13180);
nand U14489 (N_14489,N_12006,N_12627);
xnor U14490 (N_14490,N_12582,N_13136);
nor U14491 (N_14491,N_12915,N_13058);
and U14492 (N_14492,N_13141,N_13182);
or U14493 (N_14493,N_13060,N_13007);
or U14494 (N_14494,N_12748,N_13059);
xnor U14495 (N_14495,N_12648,N_12654);
nor U14496 (N_14496,N_12338,N_12343);
nor U14497 (N_14497,N_12165,N_13459);
and U14498 (N_14498,N_13461,N_12370);
nor U14499 (N_14499,N_13300,N_12117);
nand U14500 (N_14500,N_12074,N_12153);
xnor U14501 (N_14501,N_12581,N_12191);
and U14502 (N_14502,N_12114,N_12060);
nor U14503 (N_14503,N_13436,N_13031);
nor U14504 (N_14504,N_13327,N_12763);
nand U14505 (N_14505,N_12859,N_12473);
nor U14506 (N_14506,N_13222,N_13071);
xnor U14507 (N_14507,N_12430,N_12585);
nand U14508 (N_14508,N_12900,N_13295);
nor U14509 (N_14509,N_12202,N_12888);
nand U14510 (N_14510,N_12967,N_12002);
xor U14511 (N_14511,N_13160,N_13182);
nor U14512 (N_14512,N_12357,N_12903);
or U14513 (N_14513,N_12944,N_13155);
xnor U14514 (N_14514,N_12864,N_12323);
nor U14515 (N_14515,N_12381,N_13399);
nor U14516 (N_14516,N_12710,N_13481);
and U14517 (N_14517,N_12830,N_12250);
nand U14518 (N_14518,N_12764,N_13277);
nand U14519 (N_14519,N_12841,N_12675);
or U14520 (N_14520,N_12342,N_12297);
xnor U14521 (N_14521,N_13256,N_12834);
nor U14522 (N_14522,N_12597,N_12553);
nor U14523 (N_14523,N_12342,N_13319);
or U14524 (N_14524,N_12727,N_12658);
or U14525 (N_14525,N_12668,N_12446);
nor U14526 (N_14526,N_13405,N_13368);
xnor U14527 (N_14527,N_12244,N_12907);
or U14528 (N_14528,N_12657,N_12828);
nand U14529 (N_14529,N_13054,N_13212);
and U14530 (N_14530,N_12566,N_12554);
xnor U14531 (N_14531,N_13037,N_13010);
or U14532 (N_14532,N_12059,N_12266);
or U14533 (N_14533,N_12209,N_13243);
and U14534 (N_14534,N_12887,N_12464);
nand U14535 (N_14535,N_13099,N_12400);
or U14536 (N_14536,N_12469,N_13322);
and U14537 (N_14537,N_13216,N_12799);
nand U14538 (N_14538,N_12291,N_12078);
xor U14539 (N_14539,N_12902,N_13082);
nor U14540 (N_14540,N_13120,N_12286);
and U14541 (N_14541,N_12175,N_12336);
nand U14542 (N_14542,N_12092,N_12762);
nor U14543 (N_14543,N_13246,N_12954);
and U14544 (N_14544,N_13237,N_13306);
and U14545 (N_14545,N_13486,N_12330);
nor U14546 (N_14546,N_12590,N_13341);
and U14547 (N_14547,N_12569,N_12470);
xnor U14548 (N_14548,N_12913,N_12310);
and U14549 (N_14549,N_12364,N_13153);
nor U14550 (N_14550,N_12290,N_13293);
nand U14551 (N_14551,N_12493,N_12068);
or U14552 (N_14552,N_13225,N_12519);
or U14553 (N_14553,N_12227,N_12300);
or U14554 (N_14554,N_13105,N_13405);
xnor U14555 (N_14555,N_12265,N_13383);
and U14556 (N_14556,N_13334,N_13307);
nand U14557 (N_14557,N_12647,N_12745);
and U14558 (N_14558,N_12999,N_12899);
nor U14559 (N_14559,N_12832,N_12905);
or U14560 (N_14560,N_12166,N_12524);
xnor U14561 (N_14561,N_12811,N_12038);
xnor U14562 (N_14562,N_12306,N_12164);
or U14563 (N_14563,N_12179,N_13052);
xnor U14564 (N_14564,N_12773,N_13033);
or U14565 (N_14565,N_12070,N_13254);
or U14566 (N_14566,N_13168,N_13343);
xor U14567 (N_14567,N_12255,N_12276);
nand U14568 (N_14568,N_12423,N_13287);
and U14569 (N_14569,N_13499,N_12731);
and U14570 (N_14570,N_13167,N_12922);
nand U14571 (N_14571,N_12459,N_13292);
xor U14572 (N_14572,N_13319,N_13473);
xnor U14573 (N_14573,N_13096,N_12147);
nor U14574 (N_14574,N_12611,N_13362);
nor U14575 (N_14575,N_12479,N_12907);
nor U14576 (N_14576,N_12700,N_13134);
nand U14577 (N_14577,N_12930,N_13430);
nor U14578 (N_14578,N_13018,N_12802);
or U14579 (N_14579,N_12960,N_13200);
xor U14580 (N_14580,N_13464,N_12432);
xor U14581 (N_14581,N_12899,N_12509);
and U14582 (N_14582,N_12830,N_12171);
and U14583 (N_14583,N_12052,N_12821);
and U14584 (N_14584,N_12736,N_12248);
or U14585 (N_14585,N_13439,N_12168);
or U14586 (N_14586,N_12380,N_12521);
nand U14587 (N_14587,N_12798,N_13209);
nor U14588 (N_14588,N_12219,N_13130);
or U14589 (N_14589,N_13438,N_12620);
or U14590 (N_14590,N_12885,N_12841);
and U14591 (N_14591,N_12141,N_13394);
nor U14592 (N_14592,N_12294,N_12308);
xor U14593 (N_14593,N_12169,N_12701);
and U14594 (N_14594,N_12563,N_12212);
or U14595 (N_14595,N_12687,N_12623);
and U14596 (N_14596,N_12678,N_12037);
and U14597 (N_14597,N_12857,N_13196);
and U14598 (N_14598,N_13005,N_12690);
nor U14599 (N_14599,N_12744,N_13217);
or U14600 (N_14600,N_13075,N_12687);
or U14601 (N_14601,N_12083,N_13313);
nor U14602 (N_14602,N_12202,N_12106);
nand U14603 (N_14603,N_12084,N_13012);
or U14604 (N_14604,N_12133,N_12928);
or U14605 (N_14605,N_12813,N_12408);
nand U14606 (N_14606,N_13158,N_12080);
nor U14607 (N_14607,N_13283,N_12283);
and U14608 (N_14608,N_13012,N_12995);
nor U14609 (N_14609,N_12777,N_12183);
or U14610 (N_14610,N_12597,N_13426);
xor U14611 (N_14611,N_12593,N_12220);
xor U14612 (N_14612,N_12920,N_13495);
nand U14613 (N_14613,N_13432,N_12160);
and U14614 (N_14614,N_12344,N_12601);
xnor U14615 (N_14615,N_13046,N_12338);
nor U14616 (N_14616,N_12455,N_12606);
or U14617 (N_14617,N_12863,N_13099);
nand U14618 (N_14618,N_12559,N_12829);
nand U14619 (N_14619,N_13139,N_13002);
nor U14620 (N_14620,N_13133,N_12015);
and U14621 (N_14621,N_12004,N_13122);
nand U14622 (N_14622,N_12973,N_12570);
nor U14623 (N_14623,N_13159,N_12209);
or U14624 (N_14624,N_12458,N_12782);
xnor U14625 (N_14625,N_12190,N_12481);
and U14626 (N_14626,N_13208,N_13045);
nand U14627 (N_14627,N_13268,N_12489);
xnor U14628 (N_14628,N_12162,N_12919);
xor U14629 (N_14629,N_13248,N_13345);
xor U14630 (N_14630,N_13118,N_12955);
or U14631 (N_14631,N_12110,N_12739);
xor U14632 (N_14632,N_12443,N_13412);
nand U14633 (N_14633,N_12654,N_12992);
and U14634 (N_14634,N_12594,N_12232);
and U14635 (N_14635,N_13409,N_12616);
and U14636 (N_14636,N_13360,N_12966);
nor U14637 (N_14637,N_12880,N_13095);
or U14638 (N_14638,N_12830,N_12946);
nand U14639 (N_14639,N_13363,N_12329);
xnor U14640 (N_14640,N_12733,N_12274);
and U14641 (N_14641,N_12450,N_12251);
or U14642 (N_14642,N_13381,N_12767);
and U14643 (N_14643,N_12897,N_12012);
and U14644 (N_14644,N_12883,N_13264);
nand U14645 (N_14645,N_13314,N_13135);
and U14646 (N_14646,N_13349,N_12382);
xor U14647 (N_14647,N_12626,N_12888);
or U14648 (N_14648,N_13260,N_12468);
nand U14649 (N_14649,N_12495,N_12674);
and U14650 (N_14650,N_13059,N_12516);
or U14651 (N_14651,N_12309,N_13388);
nand U14652 (N_14652,N_12779,N_13457);
or U14653 (N_14653,N_12150,N_13132);
nand U14654 (N_14654,N_13334,N_12492);
nand U14655 (N_14655,N_12734,N_12215);
and U14656 (N_14656,N_12027,N_12090);
or U14657 (N_14657,N_12974,N_12697);
or U14658 (N_14658,N_12604,N_12129);
and U14659 (N_14659,N_12924,N_13215);
and U14660 (N_14660,N_12673,N_13303);
nand U14661 (N_14661,N_12590,N_12613);
nand U14662 (N_14662,N_13048,N_13029);
or U14663 (N_14663,N_12492,N_13467);
or U14664 (N_14664,N_13160,N_13218);
xnor U14665 (N_14665,N_12718,N_13248);
and U14666 (N_14666,N_13444,N_12810);
xnor U14667 (N_14667,N_12568,N_12233);
nor U14668 (N_14668,N_13280,N_13001);
or U14669 (N_14669,N_12198,N_12853);
nand U14670 (N_14670,N_12787,N_12518);
or U14671 (N_14671,N_12410,N_12791);
or U14672 (N_14672,N_12524,N_12755);
and U14673 (N_14673,N_12634,N_12381);
nand U14674 (N_14674,N_13224,N_12680);
and U14675 (N_14675,N_12623,N_12796);
nor U14676 (N_14676,N_13295,N_12394);
nor U14677 (N_14677,N_12301,N_12930);
xnor U14678 (N_14678,N_13362,N_12945);
xnor U14679 (N_14679,N_12892,N_12541);
nor U14680 (N_14680,N_12599,N_12687);
nor U14681 (N_14681,N_12307,N_12692);
or U14682 (N_14682,N_13461,N_12897);
nand U14683 (N_14683,N_12949,N_12760);
nor U14684 (N_14684,N_12289,N_12829);
nor U14685 (N_14685,N_12840,N_12100);
or U14686 (N_14686,N_12694,N_13110);
or U14687 (N_14687,N_12978,N_12586);
or U14688 (N_14688,N_12549,N_13482);
nor U14689 (N_14689,N_13228,N_12862);
and U14690 (N_14690,N_13446,N_13459);
nand U14691 (N_14691,N_12627,N_12265);
nor U14692 (N_14692,N_13267,N_13244);
xor U14693 (N_14693,N_12704,N_13048);
nor U14694 (N_14694,N_12187,N_12672);
and U14695 (N_14695,N_12497,N_12388);
nor U14696 (N_14696,N_13399,N_13474);
xnor U14697 (N_14697,N_13467,N_13369);
and U14698 (N_14698,N_13322,N_12540);
and U14699 (N_14699,N_13235,N_12284);
nand U14700 (N_14700,N_13480,N_13062);
and U14701 (N_14701,N_12188,N_12307);
and U14702 (N_14702,N_12538,N_12603);
xor U14703 (N_14703,N_13081,N_13276);
or U14704 (N_14704,N_13327,N_12459);
and U14705 (N_14705,N_12552,N_12284);
and U14706 (N_14706,N_12098,N_12778);
nand U14707 (N_14707,N_13298,N_12742);
nand U14708 (N_14708,N_12919,N_12781);
and U14709 (N_14709,N_12439,N_13404);
or U14710 (N_14710,N_12270,N_12827);
and U14711 (N_14711,N_12077,N_13427);
and U14712 (N_14712,N_12123,N_12917);
nand U14713 (N_14713,N_12674,N_13441);
nand U14714 (N_14714,N_13299,N_12687);
nand U14715 (N_14715,N_13268,N_12292);
and U14716 (N_14716,N_12772,N_13288);
xnor U14717 (N_14717,N_13276,N_12130);
xnor U14718 (N_14718,N_12018,N_12213);
or U14719 (N_14719,N_12652,N_12268);
or U14720 (N_14720,N_13293,N_12667);
xor U14721 (N_14721,N_12001,N_12855);
xnor U14722 (N_14722,N_12962,N_12879);
nand U14723 (N_14723,N_12153,N_12469);
nor U14724 (N_14724,N_13395,N_13163);
xor U14725 (N_14725,N_13434,N_12615);
nor U14726 (N_14726,N_12649,N_13477);
or U14727 (N_14727,N_12833,N_13174);
nand U14728 (N_14728,N_13010,N_12438);
nand U14729 (N_14729,N_12086,N_13299);
xor U14730 (N_14730,N_12648,N_13354);
and U14731 (N_14731,N_13391,N_12874);
xnor U14732 (N_14732,N_13480,N_12236);
nand U14733 (N_14733,N_13271,N_13056);
or U14734 (N_14734,N_12500,N_12959);
nor U14735 (N_14735,N_13436,N_12745);
nand U14736 (N_14736,N_13304,N_12899);
and U14737 (N_14737,N_13262,N_12120);
and U14738 (N_14738,N_12613,N_12902);
nand U14739 (N_14739,N_13143,N_12514);
xnor U14740 (N_14740,N_12731,N_12258);
nor U14741 (N_14741,N_12354,N_12777);
nor U14742 (N_14742,N_12966,N_13145);
nand U14743 (N_14743,N_13144,N_13236);
and U14744 (N_14744,N_13458,N_12737);
nor U14745 (N_14745,N_12289,N_12226);
nand U14746 (N_14746,N_12648,N_12065);
nand U14747 (N_14747,N_12060,N_12147);
nand U14748 (N_14748,N_12921,N_12845);
or U14749 (N_14749,N_12614,N_13007);
and U14750 (N_14750,N_12058,N_13281);
xnor U14751 (N_14751,N_12886,N_12408);
nand U14752 (N_14752,N_12907,N_12261);
xor U14753 (N_14753,N_12117,N_12590);
or U14754 (N_14754,N_13058,N_12617);
or U14755 (N_14755,N_13360,N_12407);
nor U14756 (N_14756,N_13261,N_13488);
nand U14757 (N_14757,N_13255,N_12647);
xnor U14758 (N_14758,N_12334,N_12314);
or U14759 (N_14759,N_13438,N_12487);
or U14760 (N_14760,N_13359,N_13261);
or U14761 (N_14761,N_12185,N_12009);
and U14762 (N_14762,N_13476,N_12938);
nor U14763 (N_14763,N_13369,N_12452);
or U14764 (N_14764,N_13060,N_12457);
nor U14765 (N_14765,N_12677,N_12543);
nand U14766 (N_14766,N_12727,N_12183);
or U14767 (N_14767,N_12812,N_12753);
nor U14768 (N_14768,N_12306,N_12348);
nand U14769 (N_14769,N_12089,N_13088);
or U14770 (N_14770,N_12545,N_13492);
xnor U14771 (N_14771,N_12185,N_12557);
or U14772 (N_14772,N_12838,N_12891);
nand U14773 (N_14773,N_13427,N_12763);
and U14774 (N_14774,N_13397,N_12792);
or U14775 (N_14775,N_12352,N_12624);
nor U14776 (N_14776,N_13299,N_13271);
and U14777 (N_14777,N_12435,N_13076);
and U14778 (N_14778,N_13153,N_12072);
and U14779 (N_14779,N_13470,N_12034);
and U14780 (N_14780,N_13010,N_12944);
or U14781 (N_14781,N_12902,N_13064);
and U14782 (N_14782,N_13128,N_12918);
or U14783 (N_14783,N_13074,N_12273);
nor U14784 (N_14784,N_13303,N_12850);
nor U14785 (N_14785,N_12742,N_12827);
or U14786 (N_14786,N_12718,N_12916);
or U14787 (N_14787,N_13208,N_12854);
nand U14788 (N_14788,N_12197,N_12975);
nor U14789 (N_14789,N_12869,N_12213);
nand U14790 (N_14790,N_13301,N_13070);
nor U14791 (N_14791,N_12887,N_12653);
or U14792 (N_14792,N_12964,N_13196);
nand U14793 (N_14793,N_12465,N_13238);
or U14794 (N_14794,N_13314,N_12408);
nand U14795 (N_14795,N_13245,N_12972);
nor U14796 (N_14796,N_12711,N_13233);
or U14797 (N_14797,N_13475,N_12113);
and U14798 (N_14798,N_12392,N_13466);
nand U14799 (N_14799,N_12165,N_13215);
or U14800 (N_14800,N_12373,N_12026);
nand U14801 (N_14801,N_12321,N_12393);
or U14802 (N_14802,N_12044,N_12725);
nor U14803 (N_14803,N_13478,N_13487);
and U14804 (N_14804,N_13140,N_13170);
nor U14805 (N_14805,N_12853,N_12628);
nand U14806 (N_14806,N_12138,N_12216);
nor U14807 (N_14807,N_13318,N_12738);
and U14808 (N_14808,N_12894,N_12457);
or U14809 (N_14809,N_13366,N_12734);
xor U14810 (N_14810,N_13399,N_13491);
nor U14811 (N_14811,N_13313,N_12489);
nand U14812 (N_14812,N_13034,N_12102);
xor U14813 (N_14813,N_12638,N_13241);
or U14814 (N_14814,N_13304,N_13397);
and U14815 (N_14815,N_12718,N_12683);
and U14816 (N_14816,N_12275,N_12759);
or U14817 (N_14817,N_13117,N_13106);
xnor U14818 (N_14818,N_12165,N_13151);
nand U14819 (N_14819,N_12105,N_12264);
and U14820 (N_14820,N_13044,N_12136);
or U14821 (N_14821,N_12093,N_12917);
and U14822 (N_14822,N_12794,N_12086);
nor U14823 (N_14823,N_12694,N_13140);
xnor U14824 (N_14824,N_13142,N_12963);
nand U14825 (N_14825,N_12847,N_12989);
xnor U14826 (N_14826,N_12158,N_12926);
or U14827 (N_14827,N_12049,N_13301);
xor U14828 (N_14828,N_12884,N_13076);
xnor U14829 (N_14829,N_12703,N_12704);
nor U14830 (N_14830,N_12191,N_13169);
and U14831 (N_14831,N_13096,N_12961);
nand U14832 (N_14832,N_13287,N_12449);
or U14833 (N_14833,N_13443,N_12318);
nand U14834 (N_14834,N_12930,N_13033);
nand U14835 (N_14835,N_12543,N_12603);
nor U14836 (N_14836,N_13174,N_13245);
and U14837 (N_14837,N_12653,N_13119);
and U14838 (N_14838,N_13194,N_12588);
or U14839 (N_14839,N_13226,N_13043);
and U14840 (N_14840,N_13143,N_12968);
or U14841 (N_14841,N_13414,N_12978);
or U14842 (N_14842,N_12885,N_13483);
xor U14843 (N_14843,N_12649,N_12977);
nor U14844 (N_14844,N_12005,N_13320);
xor U14845 (N_14845,N_13216,N_13240);
nand U14846 (N_14846,N_12564,N_12911);
and U14847 (N_14847,N_12488,N_12684);
and U14848 (N_14848,N_12817,N_13321);
or U14849 (N_14849,N_13058,N_12653);
or U14850 (N_14850,N_13200,N_12227);
nand U14851 (N_14851,N_13416,N_12639);
nand U14852 (N_14852,N_13256,N_12638);
nor U14853 (N_14853,N_13486,N_12837);
nand U14854 (N_14854,N_13379,N_12311);
and U14855 (N_14855,N_13313,N_13385);
nand U14856 (N_14856,N_12254,N_12429);
and U14857 (N_14857,N_12514,N_12657);
nand U14858 (N_14858,N_13242,N_12698);
and U14859 (N_14859,N_12832,N_12111);
xnor U14860 (N_14860,N_13456,N_13015);
nor U14861 (N_14861,N_12403,N_12043);
nand U14862 (N_14862,N_12411,N_13133);
and U14863 (N_14863,N_12310,N_12036);
xnor U14864 (N_14864,N_12661,N_12009);
or U14865 (N_14865,N_13023,N_13346);
nor U14866 (N_14866,N_13194,N_12360);
nand U14867 (N_14867,N_13148,N_12098);
nand U14868 (N_14868,N_12035,N_12357);
and U14869 (N_14869,N_12519,N_12698);
xor U14870 (N_14870,N_12319,N_12470);
nor U14871 (N_14871,N_12097,N_13048);
or U14872 (N_14872,N_12054,N_12064);
nand U14873 (N_14873,N_12609,N_12826);
xnor U14874 (N_14874,N_12844,N_13310);
xnor U14875 (N_14875,N_12634,N_13289);
nand U14876 (N_14876,N_12213,N_12231);
xnor U14877 (N_14877,N_12571,N_12875);
and U14878 (N_14878,N_12581,N_13237);
nor U14879 (N_14879,N_12628,N_12754);
nor U14880 (N_14880,N_13347,N_13277);
xor U14881 (N_14881,N_12764,N_12020);
or U14882 (N_14882,N_13104,N_12473);
nor U14883 (N_14883,N_12561,N_12312);
or U14884 (N_14884,N_12631,N_13240);
and U14885 (N_14885,N_13117,N_13466);
nor U14886 (N_14886,N_13431,N_12256);
nor U14887 (N_14887,N_12961,N_13084);
and U14888 (N_14888,N_13169,N_13378);
and U14889 (N_14889,N_13448,N_12258);
or U14890 (N_14890,N_13315,N_12037);
xor U14891 (N_14891,N_12197,N_13342);
nand U14892 (N_14892,N_13210,N_12536);
nor U14893 (N_14893,N_12057,N_12341);
nor U14894 (N_14894,N_13217,N_12747);
xor U14895 (N_14895,N_12564,N_12287);
nand U14896 (N_14896,N_12085,N_12489);
and U14897 (N_14897,N_12358,N_12936);
and U14898 (N_14898,N_13306,N_12279);
xnor U14899 (N_14899,N_12778,N_12864);
nand U14900 (N_14900,N_12209,N_12137);
nor U14901 (N_14901,N_13164,N_12347);
or U14902 (N_14902,N_12655,N_12878);
nand U14903 (N_14903,N_12067,N_13024);
nand U14904 (N_14904,N_12622,N_12826);
xnor U14905 (N_14905,N_13201,N_13350);
or U14906 (N_14906,N_12062,N_12736);
or U14907 (N_14907,N_13238,N_12538);
and U14908 (N_14908,N_13357,N_12507);
nor U14909 (N_14909,N_13208,N_13220);
nor U14910 (N_14910,N_13304,N_12829);
and U14911 (N_14911,N_12599,N_13453);
and U14912 (N_14912,N_12068,N_13139);
xor U14913 (N_14913,N_12375,N_12226);
and U14914 (N_14914,N_12925,N_12829);
nor U14915 (N_14915,N_12674,N_13262);
nand U14916 (N_14916,N_12435,N_12312);
or U14917 (N_14917,N_13150,N_13328);
nand U14918 (N_14918,N_12082,N_12389);
and U14919 (N_14919,N_13415,N_13265);
nand U14920 (N_14920,N_12936,N_13492);
or U14921 (N_14921,N_13350,N_12068);
or U14922 (N_14922,N_13034,N_12106);
nand U14923 (N_14923,N_12378,N_12130);
or U14924 (N_14924,N_12307,N_13182);
nand U14925 (N_14925,N_12098,N_13339);
nor U14926 (N_14926,N_12943,N_12746);
nand U14927 (N_14927,N_12652,N_12807);
nor U14928 (N_14928,N_12896,N_13408);
nand U14929 (N_14929,N_12377,N_13380);
and U14930 (N_14930,N_12973,N_13179);
nand U14931 (N_14931,N_12520,N_12483);
and U14932 (N_14932,N_12113,N_12814);
or U14933 (N_14933,N_12303,N_13363);
or U14934 (N_14934,N_12289,N_12221);
nand U14935 (N_14935,N_12471,N_12944);
nand U14936 (N_14936,N_12156,N_12630);
nand U14937 (N_14937,N_12666,N_12833);
nand U14938 (N_14938,N_12994,N_12116);
xor U14939 (N_14939,N_12263,N_12497);
xor U14940 (N_14940,N_12861,N_12840);
and U14941 (N_14941,N_13179,N_12391);
nor U14942 (N_14942,N_12595,N_12310);
and U14943 (N_14943,N_13212,N_13124);
and U14944 (N_14944,N_12014,N_12617);
and U14945 (N_14945,N_12222,N_12226);
and U14946 (N_14946,N_13058,N_12642);
and U14947 (N_14947,N_12782,N_12425);
or U14948 (N_14948,N_13348,N_12777);
xnor U14949 (N_14949,N_12857,N_12400);
and U14950 (N_14950,N_12966,N_12813);
nand U14951 (N_14951,N_13142,N_12262);
and U14952 (N_14952,N_12424,N_13295);
nand U14953 (N_14953,N_12340,N_12626);
nor U14954 (N_14954,N_12254,N_12045);
or U14955 (N_14955,N_12458,N_12695);
nand U14956 (N_14956,N_12702,N_13327);
and U14957 (N_14957,N_13091,N_13070);
or U14958 (N_14958,N_13317,N_12589);
and U14959 (N_14959,N_12307,N_13049);
nor U14960 (N_14960,N_12736,N_12956);
nor U14961 (N_14961,N_13297,N_12599);
nand U14962 (N_14962,N_13234,N_13137);
or U14963 (N_14963,N_12762,N_12699);
or U14964 (N_14964,N_12763,N_12019);
nand U14965 (N_14965,N_13336,N_12321);
nand U14966 (N_14966,N_13089,N_13445);
nor U14967 (N_14967,N_12765,N_13392);
or U14968 (N_14968,N_12508,N_12764);
nor U14969 (N_14969,N_12942,N_12138);
xnor U14970 (N_14970,N_12458,N_12187);
and U14971 (N_14971,N_13269,N_13307);
or U14972 (N_14972,N_12591,N_13173);
nor U14973 (N_14973,N_12043,N_12837);
nor U14974 (N_14974,N_12553,N_13476);
or U14975 (N_14975,N_12541,N_12739);
nand U14976 (N_14976,N_12371,N_13246);
nand U14977 (N_14977,N_12213,N_12039);
or U14978 (N_14978,N_12305,N_12074);
or U14979 (N_14979,N_12483,N_12463);
xnor U14980 (N_14980,N_13147,N_13158);
or U14981 (N_14981,N_13495,N_12003);
nor U14982 (N_14982,N_12897,N_12215);
xnor U14983 (N_14983,N_12028,N_12887);
or U14984 (N_14984,N_12753,N_13435);
nand U14985 (N_14985,N_12485,N_13239);
xnor U14986 (N_14986,N_13333,N_12294);
nor U14987 (N_14987,N_12407,N_13414);
and U14988 (N_14988,N_13375,N_12198);
nand U14989 (N_14989,N_13373,N_13022);
nor U14990 (N_14990,N_12535,N_12609);
nor U14991 (N_14991,N_12786,N_12779);
and U14992 (N_14992,N_13305,N_13119);
xor U14993 (N_14993,N_13305,N_12945);
or U14994 (N_14994,N_13410,N_12920);
and U14995 (N_14995,N_12046,N_12205);
xor U14996 (N_14996,N_13344,N_13136);
nand U14997 (N_14997,N_12285,N_12365);
and U14998 (N_14998,N_13035,N_13274);
nor U14999 (N_14999,N_13414,N_13271);
or UO_0 (O_0,N_13916,N_13769);
and UO_1 (O_1,N_13654,N_14387);
xnor UO_2 (O_2,N_13625,N_14336);
or UO_3 (O_3,N_14505,N_14028);
nand UO_4 (O_4,N_14339,N_13729);
nor UO_5 (O_5,N_14244,N_14018);
nor UO_6 (O_6,N_14254,N_14702);
and UO_7 (O_7,N_13567,N_13737);
nor UO_8 (O_8,N_14301,N_14984);
xor UO_9 (O_9,N_14682,N_14791);
or UO_10 (O_10,N_13576,N_14823);
or UO_11 (O_11,N_14590,N_14826);
nor UO_12 (O_12,N_13589,N_14478);
and UO_13 (O_13,N_14316,N_14989);
and UO_14 (O_14,N_13698,N_14651);
or UO_15 (O_15,N_14183,N_14382);
or UO_16 (O_16,N_14976,N_14374);
or UO_17 (O_17,N_14899,N_14740);
or UO_18 (O_18,N_14249,N_13914);
nor UO_19 (O_19,N_14125,N_13547);
xor UO_20 (O_20,N_14345,N_14334);
nand UO_21 (O_21,N_14430,N_13629);
or UO_22 (O_22,N_14748,N_13688);
nor UO_23 (O_23,N_14852,N_14104);
or UO_24 (O_24,N_14425,N_14137);
xor UO_25 (O_25,N_14695,N_13682);
and UO_26 (O_26,N_13930,N_13995);
nand UO_27 (O_27,N_14147,N_14156);
nand UO_28 (O_28,N_13848,N_14206);
or UO_29 (O_29,N_14732,N_14413);
xor UO_30 (O_30,N_14835,N_14502);
xor UO_31 (O_31,N_13996,N_14615);
and UO_32 (O_32,N_14436,N_14893);
and UO_33 (O_33,N_14781,N_14068);
nand UO_34 (O_34,N_13728,N_14986);
xnor UO_35 (O_35,N_13550,N_13814);
nor UO_36 (O_36,N_14884,N_13934);
nand UO_37 (O_37,N_13545,N_13689);
nand UO_38 (O_38,N_13568,N_13620);
or UO_39 (O_39,N_14012,N_14882);
nor UO_40 (O_40,N_14067,N_13598);
xnor UO_41 (O_41,N_13932,N_14433);
or UO_42 (O_42,N_14353,N_14631);
and UO_43 (O_43,N_14900,N_14971);
and UO_44 (O_44,N_14721,N_13999);
xnor UO_45 (O_45,N_14140,N_14600);
xor UO_46 (O_46,N_13865,N_14924);
and UO_47 (O_47,N_14308,N_13884);
nand UO_48 (O_48,N_14321,N_13572);
nand UO_49 (O_49,N_13778,N_13871);
nor UO_50 (O_50,N_13773,N_14077);
or UO_51 (O_51,N_14807,N_13549);
and UO_52 (O_52,N_14785,N_13507);
xor UO_53 (O_53,N_14449,N_14609);
and UO_54 (O_54,N_14938,N_14383);
or UO_55 (O_55,N_14720,N_13882);
or UO_56 (O_56,N_14729,N_14337);
nor UO_57 (O_57,N_13684,N_14146);
nor UO_58 (O_58,N_14714,N_13763);
xnor UO_59 (O_59,N_13789,N_13734);
and UO_60 (O_60,N_14375,N_14874);
or UO_61 (O_61,N_14945,N_13588);
nor UO_62 (O_62,N_13532,N_14639);
nand UO_63 (O_63,N_14532,N_13851);
nand UO_64 (O_64,N_13829,N_14351);
nor UO_65 (O_65,N_14038,N_14839);
xor UO_66 (O_66,N_14859,N_14010);
or UO_67 (O_67,N_14107,N_13958);
nand UO_68 (O_68,N_13849,N_14955);
nor UO_69 (O_69,N_14736,N_14849);
nor UO_70 (O_70,N_13745,N_13577);
or UO_71 (O_71,N_13675,N_14484);
xnor UO_72 (O_72,N_14084,N_14547);
nor UO_73 (O_73,N_14559,N_13879);
and UO_74 (O_74,N_14006,N_13883);
nand UO_75 (O_75,N_14522,N_13539);
or UO_76 (O_76,N_14396,N_14024);
nor UO_77 (O_77,N_14920,N_13847);
nand UO_78 (O_78,N_14355,N_14833);
or UO_79 (O_79,N_13519,N_14090);
nor UO_80 (O_80,N_13944,N_13509);
nand UO_81 (O_81,N_14551,N_14057);
and UO_82 (O_82,N_14412,N_13513);
xnor UO_83 (O_83,N_14579,N_14369);
xor UO_84 (O_84,N_14969,N_14359);
nand UO_85 (O_85,N_14535,N_14469);
or UO_86 (O_86,N_14529,N_13708);
xor UO_87 (O_87,N_14769,N_14799);
xnor UO_88 (O_88,N_13786,N_13881);
or UO_89 (O_89,N_13810,N_13861);
nor UO_90 (O_90,N_14890,N_13942);
or UO_91 (O_91,N_13659,N_13713);
or UO_92 (O_92,N_14891,N_13854);
nor UO_93 (O_93,N_14466,N_13523);
or UO_94 (O_94,N_14297,N_14222);
nand UO_95 (O_95,N_13959,N_14592);
xor UO_96 (O_96,N_13649,N_14101);
or UO_97 (O_97,N_14232,N_13735);
and UO_98 (O_98,N_14442,N_14652);
or UO_99 (O_99,N_14565,N_13771);
or UO_100 (O_100,N_14069,N_14628);
and UO_101 (O_101,N_14817,N_14541);
and UO_102 (O_102,N_14908,N_13543);
and UO_103 (O_103,N_14548,N_14256);
xnor UO_104 (O_104,N_14824,N_13945);
and UO_105 (O_105,N_14406,N_14014);
and UO_106 (O_106,N_14919,N_14685);
or UO_107 (O_107,N_14634,N_13899);
or UO_108 (O_108,N_14870,N_14867);
nand UO_109 (O_109,N_13901,N_14755);
xor UO_110 (O_110,N_14260,N_14997);
or UO_111 (O_111,N_14191,N_14462);
nor UO_112 (O_112,N_13823,N_14693);
nand UO_113 (O_113,N_14161,N_13950);
or UO_114 (O_114,N_14831,N_14468);
xor UO_115 (O_115,N_13955,N_14519);
and UO_116 (O_116,N_14197,N_14338);
nor UO_117 (O_117,N_13667,N_14362);
xor UO_118 (O_118,N_13716,N_13749);
nor UO_119 (O_119,N_13746,N_14784);
and UO_120 (O_120,N_13650,N_14610);
nand UO_121 (O_121,N_14931,N_14832);
nor UO_122 (O_122,N_14860,N_14019);
nand UO_123 (O_123,N_14388,N_13967);
xnor UO_124 (O_124,N_14918,N_13681);
nand UO_125 (O_125,N_14758,N_14072);
and UO_126 (O_126,N_14681,N_14789);
nand UO_127 (O_127,N_14738,N_14991);
and UO_128 (O_128,N_14779,N_14135);
nor UO_129 (O_129,N_14778,N_14295);
xor UO_130 (O_130,N_13866,N_13564);
nor UO_131 (O_131,N_13834,N_14795);
nor UO_132 (O_132,N_14536,N_14042);
and UO_133 (O_133,N_14542,N_13727);
or UO_134 (O_134,N_14453,N_14507);
or UO_135 (O_135,N_14647,N_14401);
and UO_136 (O_136,N_13836,N_14952);
and UO_137 (O_137,N_14193,N_14127);
or UO_138 (O_138,N_14648,N_13972);
or UO_139 (O_139,N_13556,N_14927);
nor UO_140 (O_140,N_14731,N_14698);
xor UO_141 (O_141,N_13977,N_13919);
nand UO_142 (O_142,N_14950,N_14240);
and UO_143 (O_143,N_14854,N_13685);
nand UO_144 (O_144,N_14129,N_14613);
nor UO_145 (O_145,N_13692,N_13726);
nand UO_146 (O_146,N_14805,N_14379);
nor UO_147 (O_147,N_14344,N_14747);
and UO_148 (O_148,N_13691,N_14110);
or UO_149 (O_149,N_14076,N_13824);
nor UO_150 (O_150,N_14490,N_13792);
xnor UO_151 (O_151,N_14864,N_13574);
xnor UO_152 (O_152,N_13639,N_14100);
xor UO_153 (O_153,N_14585,N_14460);
and UO_154 (O_154,N_14207,N_13788);
and UO_155 (O_155,N_13898,N_14112);
nor UO_156 (O_156,N_14116,N_13571);
and UO_157 (O_157,N_14684,N_14058);
and UO_158 (O_158,N_13638,N_14134);
nor UO_159 (O_159,N_14538,N_13918);
and UO_160 (O_160,N_14939,N_13806);
nor UO_161 (O_161,N_14461,N_13538);
and UO_162 (O_162,N_14080,N_13864);
xor UO_163 (O_163,N_14537,N_14558);
xor UO_164 (O_164,N_13961,N_14996);
nor UO_165 (O_165,N_13604,N_14054);
xnor UO_166 (O_166,N_14403,N_14262);
and UO_167 (O_167,N_14782,N_14837);
or UO_168 (O_168,N_13935,N_14828);
or UO_169 (O_169,N_14840,N_13828);
and UO_170 (O_170,N_14964,N_14053);
nor UO_171 (O_171,N_13926,N_14347);
nor UO_172 (O_172,N_14153,N_14342);
and UO_173 (O_173,N_14354,N_14661);
or UO_174 (O_174,N_14581,N_13785);
and UO_175 (O_175,N_13776,N_13596);
xnor UO_176 (O_176,N_14987,N_14437);
nand UO_177 (O_177,N_14357,N_14489);
and UO_178 (O_178,N_14589,N_14117);
xor UO_179 (O_179,N_13674,N_14052);
nand UO_180 (O_180,N_14944,N_13570);
or UO_181 (O_181,N_13744,N_14757);
or UO_182 (O_182,N_14570,N_13575);
nor UO_183 (O_183,N_13796,N_13906);
nand UO_184 (O_184,N_14421,N_14340);
or UO_185 (O_185,N_13634,N_13801);
and UO_186 (O_186,N_14448,N_14348);
nor UO_187 (O_187,N_13578,N_14119);
xor UO_188 (O_188,N_13712,N_14377);
or UO_189 (O_189,N_14764,N_13584);
nor UO_190 (O_190,N_14584,N_14177);
xnor UO_191 (O_191,N_13647,N_13764);
and UO_192 (O_192,N_14213,N_14994);
nand UO_193 (O_193,N_14236,N_14349);
and UO_194 (O_194,N_14158,N_14754);
xnor UO_195 (O_195,N_14319,N_14903);
xor UO_196 (O_196,N_14620,N_14500);
xnor UO_197 (O_197,N_14335,N_14166);
nand UO_198 (O_198,N_13582,N_14850);
nor UO_199 (O_199,N_14465,N_13943);
or UO_200 (O_200,N_14103,N_13740);
xor UO_201 (O_201,N_14091,N_14482);
nand UO_202 (O_202,N_14414,N_14325);
nand UO_203 (O_203,N_14056,N_14573);
nor UO_204 (O_204,N_14801,N_14051);
and UO_205 (O_205,N_13895,N_13803);
xnor UO_206 (O_206,N_14270,N_14133);
and UO_207 (O_207,N_13984,N_14762);
xnor UO_208 (O_208,N_14668,N_14591);
nor UO_209 (O_209,N_14739,N_14305);
or UO_210 (O_210,N_13911,N_13892);
nand UO_211 (O_211,N_13599,N_13817);
or UO_212 (O_212,N_13887,N_14595);
nor UO_213 (O_213,N_14564,N_13794);
and UO_214 (O_214,N_13795,N_13753);
nor UO_215 (O_215,N_13970,N_14128);
nand UO_216 (O_216,N_14518,N_14247);
and UO_217 (O_217,N_13951,N_14873);
xnor UO_218 (O_218,N_14201,N_14367);
and UO_219 (O_219,N_13700,N_14567);
xnor UO_220 (O_220,N_14641,N_14350);
xnor UO_221 (O_221,N_14456,N_14094);
xor UO_222 (O_222,N_13630,N_13525);
or UO_223 (O_223,N_13891,N_14632);
or UO_224 (O_224,N_14095,N_13956);
and UO_225 (O_225,N_14243,N_14679);
or UO_226 (O_226,N_14196,N_14717);
or UO_227 (O_227,N_13907,N_14642);
xnor UO_228 (O_228,N_13989,N_14200);
nand UO_229 (O_229,N_14809,N_14926);
and UO_230 (O_230,N_13548,N_14176);
or UO_231 (O_231,N_14307,N_13842);
and UO_232 (O_232,N_14138,N_14497);
nor UO_233 (O_233,N_14626,N_14189);
nand UO_234 (O_234,N_14370,N_14814);
and UO_235 (O_235,N_14263,N_13998);
or UO_236 (O_236,N_14376,N_14261);
nand UO_237 (O_237,N_13645,N_14552);
or UO_238 (O_238,N_14672,N_14399);
and UO_239 (O_239,N_14509,N_14568);
and UO_240 (O_240,N_13720,N_13888);
and UO_241 (O_241,N_14363,N_14982);
or UO_242 (O_242,N_14735,N_14188);
nor UO_243 (O_243,N_13867,N_14190);
nor UO_244 (O_244,N_14390,N_14673);
and UO_245 (O_245,N_14088,N_14861);
and UO_246 (O_246,N_14312,N_13562);
or UO_247 (O_247,N_14961,N_14296);
or UO_248 (O_248,N_14265,N_14149);
and UO_249 (O_249,N_13660,N_14278);
or UO_250 (O_250,N_13535,N_14773);
or UO_251 (O_251,N_13731,N_14358);
nor UO_252 (O_252,N_14109,N_14474);
nor UO_253 (O_253,N_14148,N_14599);
xnor UO_254 (O_254,N_14637,N_14032);
or UO_255 (O_255,N_13939,N_14667);
and UO_256 (O_256,N_14875,N_14210);
and UO_257 (O_257,N_13678,N_14666);
xor UO_258 (O_258,N_14633,N_13949);
and UO_259 (O_259,N_13971,N_13591);
nor UO_260 (O_260,N_13511,N_14513);
nand UO_261 (O_261,N_14934,N_14970);
or UO_262 (O_262,N_13710,N_14528);
nand UO_263 (O_263,N_14527,N_14040);
xnor UO_264 (O_264,N_14441,N_13602);
xor UO_265 (O_265,N_14612,N_14315);
xnor UO_266 (O_266,N_13858,N_14005);
or UO_267 (O_267,N_14768,N_13832);
or UO_268 (O_268,N_14851,N_14677);
and UO_269 (O_269,N_14108,N_13644);
and UO_270 (O_270,N_13723,N_13504);
xnor UO_271 (O_271,N_14417,N_13669);
nand UO_272 (O_272,N_14230,N_14343);
xor UO_273 (O_273,N_14689,N_13921);
nor UO_274 (O_274,N_13515,N_14749);
and UO_275 (O_275,N_13615,N_14877);
xor UO_276 (O_276,N_14604,N_13623);
and UO_277 (O_277,N_13752,N_14907);
xor UO_278 (O_278,N_13982,N_14487);
and UO_279 (O_279,N_13846,N_13718);
nand UO_280 (O_280,N_14871,N_13985);
xor UO_281 (O_281,N_14726,N_13812);
nand UO_282 (O_282,N_14578,N_14766);
nor UO_283 (O_283,N_14120,N_13987);
and UO_284 (O_284,N_14182,N_13553);
or UO_285 (O_285,N_14957,N_14404);
and UO_286 (O_286,N_14479,N_14838);
or UO_287 (O_287,N_14777,N_14154);
xor UO_288 (O_288,N_14495,N_14415);
xnor UO_289 (O_289,N_14221,N_13819);
nand UO_290 (O_290,N_13910,N_14883);
or UO_291 (O_291,N_14025,N_14715);
or UO_292 (O_292,N_14352,N_13501);
xor UO_293 (O_293,N_14744,N_13637);
and UO_294 (O_294,N_13830,N_13920);
and UO_295 (O_295,N_14205,N_13527);
or UO_296 (O_296,N_14886,N_13671);
xnor UO_297 (O_297,N_14725,N_13791);
xor UO_298 (O_298,N_14092,N_13779);
nor UO_299 (O_299,N_14765,N_14400);
and UO_300 (O_300,N_14458,N_14501);
nand UO_301 (O_301,N_14075,N_14793);
or UO_302 (O_302,N_13973,N_14029);
xnor UO_303 (O_303,N_14391,N_14163);
nor UO_304 (O_304,N_14627,N_14802);
and UO_305 (O_305,N_13612,N_14439);
and UO_306 (O_306,N_13631,N_14365);
nor UO_307 (O_307,N_14252,N_14728);
nand UO_308 (O_308,N_14311,N_13923);
xnor UO_309 (O_309,N_14921,N_14447);
nand UO_310 (O_310,N_13711,N_14402);
or UO_311 (O_311,N_14905,N_14130);
xnor UO_312 (O_312,N_14422,N_13948);
nand UO_313 (O_313,N_14911,N_13757);
xnor UO_314 (O_314,N_14533,N_13811);
or UO_315 (O_315,N_14942,N_14514);
or UO_316 (O_316,N_13903,N_14630);
nor UO_317 (O_317,N_13521,N_14203);
or UO_318 (O_318,N_14373,N_14653);
nor UO_319 (O_319,N_13859,N_13632);
or UO_320 (O_320,N_13761,N_14023);
or UO_321 (O_321,N_13839,N_13536);
or UO_322 (O_322,N_14954,N_13852);
nor UO_323 (O_323,N_14546,N_14385);
or UO_324 (O_324,N_13544,N_13636);
or UO_325 (O_325,N_14033,N_13936);
xnor UO_326 (O_326,N_14803,N_14678);
nand UO_327 (O_327,N_14277,N_13904);
and UO_328 (O_328,N_14691,N_13651);
xor UO_329 (O_329,N_13551,N_14115);
nor UO_330 (O_330,N_13826,N_14360);
and UO_331 (O_331,N_14635,N_14515);
or UO_332 (O_332,N_13520,N_14499);
xnor UO_333 (O_333,N_14186,N_14164);
or UO_334 (O_334,N_14872,N_14792);
nor UO_335 (O_335,N_14951,N_13704);
or UO_336 (O_336,N_13941,N_14445);
nand UO_337 (O_337,N_14978,N_14046);
and UO_338 (O_338,N_14111,N_14159);
nor UO_339 (O_339,N_13868,N_13503);
or UO_340 (O_340,N_14371,N_14572);
nand UO_341 (O_341,N_14250,N_13673);
nand UO_342 (O_342,N_13502,N_14842);
xor UO_343 (O_343,N_13743,N_13793);
and UO_344 (O_344,N_13980,N_14910);
and UO_345 (O_345,N_13896,N_14577);
xnor UO_346 (O_346,N_14272,N_14550);
or UO_347 (O_347,N_13686,N_13872);
nand UO_348 (O_348,N_14096,N_13557);
xor UO_349 (O_349,N_14259,N_14155);
nand UO_350 (O_350,N_13885,N_14786);
nand UO_351 (O_351,N_14880,N_14914);
nand UO_352 (O_352,N_14988,N_13862);
nand UO_353 (O_353,N_13831,N_14061);
and UO_354 (O_354,N_14083,N_13991);
nand UO_355 (O_355,N_14424,N_13770);
xor UO_356 (O_356,N_14574,N_14366);
nand UO_357 (O_357,N_14995,N_13546);
xnor UO_358 (O_358,N_14645,N_14411);
nand UO_359 (O_359,N_14796,N_14322);
and UO_360 (O_360,N_14772,N_14444);
xnor UO_361 (O_361,N_13593,N_14692);
xor UO_362 (O_362,N_14560,N_14037);
or UO_363 (O_363,N_14055,N_13755);
nor UO_364 (O_364,N_13601,N_14967);
nor UO_365 (O_365,N_14790,N_14407);
xor UO_366 (O_366,N_14993,N_14361);
and UO_367 (O_367,N_14394,N_14708);
xor UO_368 (O_368,N_13821,N_14030);
nand UO_369 (O_369,N_14936,N_14162);
or UO_370 (O_370,N_14284,N_14865);
nand UO_371 (O_371,N_14718,N_14670);
xor UO_372 (O_372,N_14271,N_14794);
nor UO_373 (O_373,N_14226,N_14602);
nand UO_374 (O_374,N_14016,N_14733);
nor UO_375 (O_375,N_14869,N_13643);
xor UO_376 (O_376,N_14257,N_13924);
or UO_377 (O_377,N_13869,N_14300);
nand UO_378 (O_378,N_14812,N_13626);
nor UO_379 (O_379,N_14743,N_14123);
nor UO_380 (O_380,N_14876,N_14434);
nor UO_381 (O_381,N_14330,N_14687);
nand UO_382 (O_382,N_14273,N_14477);
or UO_383 (O_383,N_14915,N_14082);
or UO_384 (O_384,N_14834,N_14846);
or UO_385 (O_385,N_13687,N_14575);
and UO_386 (O_386,N_14225,N_14195);
or UO_387 (O_387,N_14897,N_13751);
and UO_388 (O_388,N_13677,N_14118);
or UO_389 (O_389,N_14956,N_14486);
and UO_390 (O_390,N_13838,N_13528);
and UO_391 (O_391,N_13610,N_14549);
nand UO_392 (O_392,N_14804,N_14664);
xor UO_393 (O_393,N_14853,N_14429);
or UO_394 (O_394,N_14064,N_13510);
nand UO_395 (O_395,N_14291,N_14675);
nor UO_396 (O_396,N_13974,N_14021);
and UO_397 (O_397,N_14496,N_14488);
nand UO_398 (O_398,N_14346,N_14822);
nor UO_399 (O_399,N_13760,N_14912);
nand UO_400 (O_400,N_13542,N_13714);
or UO_401 (O_401,N_13621,N_13524);
xnor UO_402 (O_402,N_13709,N_14294);
nor UO_403 (O_403,N_14821,N_13701);
and UO_404 (O_404,N_13850,N_13878);
nor UO_405 (O_405,N_14650,N_14686);
or UO_406 (O_406,N_13693,N_14255);
nand UO_407 (O_407,N_14211,N_13706);
nor UO_408 (O_408,N_14829,N_13683);
and UO_409 (O_409,N_14504,N_14212);
nor UO_410 (O_410,N_14654,N_13635);
nor UO_411 (O_411,N_13840,N_14697);
xor UO_412 (O_412,N_14034,N_14144);
or UO_413 (O_413,N_14087,N_13915);
or UO_414 (O_414,N_13799,N_14566);
nor UO_415 (O_415,N_13890,N_13870);
or UO_416 (O_416,N_13863,N_14827);
or UO_417 (O_417,N_14384,N_14719);
or UO_418 (O_418,N_14776,N_14198);
or UO_419 (O_419,N_13561,N_13512);
nand UO_420 (O_420,N_14694,N_13900);
or UO_421 (O_421,N_14623,N_14426);
nand UO_422 (O_422,N_14480,N_14596);
or UO_423 (O_423,N_13954,N_13783);
nand UO_424 (O_424,N_14676,N_13702);
xor UO_425 (O_425,N_14431,N_13952);
xor UO_426 (O_426,N_14446,N_13889);
xnor UO_427 (O_427,N_14202,N_14493);
nor UO_428 (O_428,N_14081,N_14601);
xor UO_429 (O_429,N_13500,N_14381);
nand UO_430 (O_430,N_14690,N_14026);
nor UO_431 (O_431,N_14862,N_14761);
nand UO_432 (O_432,N_14475,N_14467);
nor UO_433 (O_433,N_13975,N_14539);
or UO_434 (O_434,N_14009,N_14928);
xnor UO_435 (O_435,N_14949,N_13762);
xor UO_436 (O_436,N_14665,N_14015);
and UO_437 (O_437,N_14086,N_13559);
nor UO_438 (O_438,N_14659,N_14309);
or UO_439 (O_439,N_14783,N_14975);
or UO_440 (O_440,N_14410,N_13725);
or UO_441 (O_441,N_14750,N_14711);
nand UO_442 (O_442,N_13707,N_14450);
nor UO_443 (O_443,N_13913,N_14065);
xor UO_444 (O_444,N_14131,N_14660);
xor UO_445 (O_445,N_13624,N_14231);
or UO_446 (O_446,N_14341,N_14368);
nand UO_447 (O_447,N_13517,N_14455);
nand UO_448 (O_448,N_14048,N_14220);
xor UO_449 (O_449,N_14810,N_13573);
or UO_450 (O_450,N_14745,N_14516);
xnor UO_451 (O_451,N_13979,N_14098);
nand UO_452 (O_452,N_14953,N_14658);
or UO_453 (O_453,N_13595,N_14848);
xnor UO_454 (O_454,N_14844,N_14280);
and UO_455 (O_455,N_14160,N_14264);
or UO_456 (O_456,N_14638,N_14451);
or UO_457 (O_457,N_13617,N_14286);
and UO_458 (O_458,N_14171,N_14473);
xor UO_459 (O_459,N_13505,N_13940);
and UO_460 (O_460,N_14287,N_13628);
and UO_461 (O_461,N_14644,N_14963);
nor UO_462 (O_462,N_13988,N_14616);
or UO_463 (O_463,N_13614,N_14857);
nand UO_464 (O_464,N_14699,N_13668);
xnor UO_465 (O_465,N_14770,N_14895);
or UO_466 (O_466,N_14730,N_14845);
nor UO_467 (O_467,N_14419,N_14132);
xor UO_468 (O_468,N_14930,N_14248);
nand UO_469 (O_469,N_13963,N_14204);
nor UO_470 (O_470,N_14416,N_13648);
nor UO_471 (O_471,N_14947,N_14798);
or UO_472 (O_472,N_14471,N_13531);
xor UO_473 (O_473,N_13606,N_13530);
xnor UO_474 (O_474,N_14904,N_14598);
or UO_475 (O_475,N_14003,N_14901);
nor UO_476 (O_476,N_13603,N_13790);
and UO_477 (O_477,N_14737,N_14289);
or UO_478 (O_478,N_14960,N_13736);
nor UO_479 (O_479,N_13680,N_14935);
and UO_480 (O_480,N_14011,N_13966);
xnor UO_481 (O_481,N_13797,N_13581);
xor UO_482 (O_482,N_14605,N_13880);
nand UO_483 (O_483,N_14680,N_13784);
xnor UO_484 (O_484,N_14013,N_14288);
nand UO_485 (O_485,N_14215,N_14071);
nand UO_486 (O_486,N_13537,N_14275);
and UO_487 (O_487,N_13613,N_13741);
and UO_488 (O_488,N_13640,N_13694);
and UO_489 (O_489,N_13611,N_14246);
or UO_490 (O_490,N_13937,N_13666);
or UO_491 (O_491,N_13526,N_14483);
nor UO_492 (O_492,N_14258,N_14093);
or UO_493 (O_493,N_14304,N_14800);
nor UO_494 (O_494,N_13855,N_14517);
or UO_495 (O_495,N_14524,N_14998);
nor UO_496 (O_496,N_13809,N_14655);
and UO_497 (O_497,N_14126,N_14896);
or UO_498 (O_498,N_14656,N_14887);
nor UO_499 (O_499,N_14356,N_14556);
xor UO_500 (O_500,N_13750,N_14888);
nand UO_501 (O_501,N_13893,N_13815);
nand UO_502 (O_502,N_14121,N_14775);
xor UO_503 (O_503,N_14588,N_13585);
or UO_504 (O_504,N_13927,N_14863);
and UO_505 (O_505,N_14741,N_13697);
nor UO_506 (O_506,N_13627,N_14723);
and UO_507 (O_507,N_13619,N_14443);
nand UO_508 (O_508,N_14165,N_14925);
or UO_509 (O_509,N_14705,N_14932);
and UO_510 (O_510,N_13800,N_14281);
nand UO_511 (O_511,N_14561,N_14303);
nand UO_512 (O_512,N_13747,N_14510);
or UO_513 (O_513,N_13925,N_14788);
xnor UO_514 (O_514,N_13820,N_14700);
nor UO_515 (O_515,N_14031,N_14079);
or UO_516 (O_516,N_14405,N_14485);
and UO_517 (O_517,N_14526,N_13845);
nor UO_518 (O_518,N_14181,N_14320);
or UO_519 (O_519,N_14228,N_14587);
nor UO_520 (O_520,N_14855,N_14313);
nor UO_521 (O_521,N_14820,N_14622);
xnor UO_522 (O_522,N_14923,N_14216);
and UO_523 (O_523,N_14688,N_13873);
xor UO_524 (O_524,N_14318,N_14576);
and UO_525 (O_525,N_14624,N_14734);
and UO_526 (O_526,N_14968,N_13960);
xnor UO_527 (O_527,N_13665,N_13518);
and UO_528 (O_528,N_13554,N_14269);
or UO_529 (O_529,N_14427,N_14227);
nand UO_530 (O_530,N_13768,N_13739);
or UO_531 (O_531,N_14251,N_14941);
and UO_532 (O_532,N_14224,N_14386);
nor UO_533 (O_533,N_14085,N_13670);
and UO_534 (O_534,N_13983,N_13529);
nor UO_535 (O_535,N_14326,N_13695);
nor UO_536 (O_536,N_14078,N_14751);
xor UO_537 (O_537,N_13997,N_14290);
xor UO_538 (O_538,N_14563,N_14314);
or UO_539 (O_539,N_14174,N_14122);
or UO_540 (O_540,N_14981,N_13875);
nand UO_541 (O_541,N_14797,N_14192);
nand UO_542 (O_542,N_14457,N_13837);
nand UO_543 (O_543,N_14506,N_14742);
nor UO_544 (O_544,N_14136,N_14555);
nor UO_545 (O_545,N_14380,N_13733);
xor UO_546 (O_546,N_13835,N_13633);
xnor UO_547 (O_547,N_14724,N_14008);
xor UO_548 (O_548,N_13579,N_13690);
nor UO_549 (O_549,N_14614,N_14073);
xor UO_550 (O_550,N_14293,N_13597);
xnor UO_551 (O_551,N_13586,N_14238);
nor UO_552 (O_552,N_13679,N_13876);
or UO_553 (O_553,N_13798,N_14836);
and UO_554 (O_554,N_13986,N_13843);
nand UO_555 (O_555,N_13732,N_13874);
nor UO_556 (O_556,N_14266,N_14825);
nand UO_557 (O_557,N_14571,N_14707);
or UO_558 (O_558,N_14841,N_13565);
nor UO_559 (O_559,N_14916,N_14102);
or UO_560 (O_560,N_14492,N_14617);
xor UO_561 (O_561,N_14063,N_14027);
or UO_562 (O_562,N_13922,N_14557);
nand UO_563 (O_563,N_14167,N_13860);
xnor UO_564 (O_564,N_14965,N_14173);
or UO_565 (O_565,N_14180,N_14440);
nand UO_566 (O_566,N_13516,N_14819);
or UO_567 (O_567,N_13580,N_13993);
and UO_568 (O_568,N_14141,N_14806);
and UO_569 (O_569,N_14621,N_14049);
or UO_570 (O_570,N_14607,N_14113);
nor UO_571 (O_571,N_14157,N_13827);
and UO_572 (O_572,N_14323,N_14521);
nor UO_573 (O_573,N_14234,N_14597);
xor UO_574 (O_574,N_14889,N_14992);
and UO_575 (O_575,N_14178,N_14554);
nor UO_576 (O_576,N_13990,N_14716);
nand UO_577 (O_577,N_13802,N_13600);
nand UO_578 (O_578,N_14674,N_13777);
xor UO_579 (O_579,N_13969,N_14712);
nor UO_580 (O_580,N_14372,N_14324);
xnor UO_581 (O_581,N_14759,N_14233);
or UO_582 (O_582,N_13912,N_14858);
or UO_583 (O_583,N_13641,N_14432);
nor UO_584 (O_584,N_13658,N_14124);
and UO_585 (O_585,N_13722,N_13938);
and UO_586 (O_586,N_14771,N_14237);
nand UO_587 (O_587,N_14285,N_14544);
nand UO_588 (O_588,N_14209,N_13653);
nor UO_589 (O_589,N_14868,N_14847);
nor UO_590 (O_590,N_14472,N_13533);
xor UO_591 (O_591,N_13696,N_14937);
or UO_592 (O_592,N_14948,N_13608);
nor UO_593 (O_593,N_14097,N_14044);
nor UO_594 (O_594,N_14606,N_14306);
nor UO_595 (O_595,N_14640,N_14946);
nand UO_596 (O_596,N_14331,N_13902);
nand UO_597 (O_597,N_14618,N_14922);
nor UO_598 (O_598,N_14459,N_14977);
or UO_599 (O_599,N_14636,N_14105);
xnor UO_600 (O_600,N_14047,N_13774);
or UO_601 (O_601,N_14017,N_14787);
and UO_602 (O_602,N_14512,N_14282);
nor UO_603 (O_603,N_14170,N_14036);
xor UO_604 (O_604,N_13818,N_14435);
or UO_605 (O_605,N_14780,N_14959);
xor UO_606 (O_606,N_14543,N_14274);
xor UO_607 (O_607,N_14218,N_13705);
xnor UO_608 (O_608,N_13767,N_13908);
nand UO_609 (O_609,N_14333,N_13555);
xnor UO_610 (O_610,N_13699,N_14898);
nand UO_611 (O_611,N_14746,N_13759);
and UO_612 (O_612,N_14267,N_14169);
nand UO_613 (O_613,N_14917,N_14974);
nand UO_614 (O_614,N_13994,N_13622);
nand UO_615 (O_615,N_14856,N_13844);
nand UO_616 (O_616,N_13721,N_14973);
or UO_617 (O_617,N_14398,N_13962);
and UO_618 (O_618,N_13816,N_13780);
or UO_619 (O_619,N_14508,N_14902);
nand UO_620 (O_620,N_14913,N_13583);
nor UO_621 (O_621,N_13657,N_14043);
xor UO_622 (O_622,N_14683,N_13964);
xor UO_623 (O_623,N_14470,N_14143);
and UO_624 (O_624,N_13756,N_13616);
or UO_625 (O_625,N_14878,N_14525);
nor UO_626 (O_626,N_13618,N_13877);
nor UO_627 (O_627,N_13663,N_14393);
and UO_628 (O_628,N_14420,N_13672);
or UO_629 (O_629,N_14106,N_14151);
nand UO_630 (O_630,N_13506,N_14022);
nand UO_631 (O_631,N_14843,N_13931);
or UO_632 (O_632,N_14007,N_14696);
and UO_633 (O_633,N_13929,N_14979);
nand UO_634 (O_634,N_13782,N_13953);
or UO_635 (O_635,N_14586,N_14179);
nand UO_636 (O_636,N_14906,N_14881);
xnor UO_637 (O_637,N_14142,N_14753);
nand UO_638 (O_638,N_13947,N_14752);
or UO_639 (O_639,N_14214,N_14958);
nor UO_640 (O_640,N_14299,N_14438);
and UO_641 (O_641,N_14643,N_14229);
xor UO_642 (O_642,N_14452,N_14463);
nand UO_643 (O_643,N_14663,N_14980);
nand UO_644 (O_644,N_14545,N_14763);
nand UO_645 (O_645,N_14966,N_14185);
or UO_646 (O_646,N_13933,N_13592);
nor UO_647 (O_647,N_13772,N_14039);
and UO_648 (O_648,N_13738,N_13661);
nand UO_649 (O_649,N_14530,N_14253);
nor UO_650 (O_650,N_14990,N_14378);
nand UO_651 (O_651,N_13730,N_14152);
nand UO_652 (O_652,N_13552,N_14657);
xor UO_653 (O_653,N_13758,N_14020);
nand UO_654 (O_654,N_14818,N_14608);
xnor UO_655 (O_655,N_14327,N_14235);
xor UO_656 (O_656,N_14710,N_14423);
or UO_657 (O_657,N_13569,N_14611);
xnor UO_658 (O_658,N_14511,N_14476);
nand UO_659 (O_659,N_14866,N_14328);
or UO_660 (O_660,N_14619,N_13587);
nor UO_661 (O_661,N_14662,N_14139);
or UO_662 (O_662,N_14364,N_14830);
nand UO_663 (O_663,N_14114,N_14208);
and UO_664 (O_664,N_14649,N_13787);
xor UO_665 (O_665,N_13897,N_13703);
nand UO_666 (O_666,N_13781,N_14892);
nor UO_667 (O_667,N_14706,N_14756);
xor UO_668 (O_668,N_14060,N_13917);
nand UO_669 (O_669,N_14494,N_13646);
and UO_670 (O_670,N_13825,N_13590);
xnor UO_671 (O_671,N_14418,N_13664);
and UO_672 (O_672,N_14503,N_14150);
and UO_673 (O_673,N_14002,N_13856);
nand UO_674 (O_674,N_13717,N_13905);
and UO_675 (O_675,N_14534,N_14972);
nand UO_676 (O_676,N_14242,N_13642);
nor UO_677 (O_677,N_14671,N_14879);
nand UO_678 (O_678,N_13968,N_14940);
nor UO_679 (O_679,N_13594,N_14722);
nor UO_680 (O_680,N_13560,N_14603);
xor UO_681 (O_681,N_13853,N_14241);
nor UO_682 (O_682,N_13766,N_13909);
and UO_683 (O_683,N_14999,N_14145);
xnor UO_684 (O_684,N_14219,N_14194);
xor UO_685 (O_685,N_14045,N_14059);
nor UO_686 (O_686,N_14815,N_14704);
xor UO_687 (O_687,N_14245,N_14050);
and UO_688 (O_688,N_14491,N_14943);
xor UO_689 (O_689,N_13656,N_14816);
and UO_690 (O_690,N_13609,N_14464);
xor UO_691 (O_691,N_13719,N_14962);
nor UO_692 (O_692,N_13508,N_14000);
nand UO_693 (O_693,N_14041,N_14070);
nand UO_694 (O_694,N_14292,N_13558);
or UO_695 (O_695,N_13981,N_14540);
and UO_696 (O_696,N_14727,N_13805);
or UO_697 (O_697,N_13992,N_14397);
or UO_698 (O_698,N_13662,N_14239);
xor UO_699 (O_699,N_14099,N_14268);
xor UO_700 (O_700,N_14553,N_14593);
or UO_701 (O_701,N_14074,N_14184);
or UO_702 (O_702,N_14709,N_13976);
or UO_703 (O_703,N_14066,N_14669);
nor UO_704 (O_704,N_14454,N_14713);
nor UO_705 (O_705,N_13514,N_13724);
xnor UO_706 (O_706,N_14004,N_14172);
and UO_707 (O_707,N_14302,N_13841);
nand UO_708 (O_708,N_13715,N_14583);
nor UO_709 (O_709,N_13808,N_13754);
and UO_710 (O_710,N_13652,N_14392);
and UO_711 (O_711,N_13886,N_14569);
and UO_712 (O_712,N_14283,N_14625);
nand UO_713 (O_713,N_14562,N_14035);
nand UO_714 (O_714,N_13563,N_14531);
xor UO_715 (O_715,N_14217,N_14885);
or UO_716 (O_716,N_14813,N_14811);
or UO_717 (O_717,N_14894,N_14332);
nand UO_718 (O_718,N_14199,N_13607);
nor UO_719 (O_719,N_14909,N_14062);
xor UO_720 (O_720,N_13978,N_13540);
nor UO_721 (O_721,N_13894,N_13566);
nand UO_722 (O_722,N_14223,N_14395);
nor UO_723 (O_723,N_14594,N_14409);
or UO_724 (O_724,N_13946,N_14520);
nor UO_725 (O_725,N_14523,N_14279);
nand UO_726 (O_726,N_13676,N_14310);
xnor UO_727 (O_727,N_13833,N_13748);
nor UO_728 (O_728,N_14317,N_13807);
nor UO_729 (O_729,N_14168,N_13857);
xor UO_730 (O_730,N_13775,N_14646);
and UO_731 (O_731,N_14329,N_13605);
xnor UO_732 (O_732,N_14187,N_14408);
and UO_733 (O_733,N_14985,N_14580);
or UO_734 (O_734,N_14298,N_14428);
nand UO_735 (O_735,N_13957,N_13522);
and UO_736 (O_736,N_14001,N_14774);
nand UO_737 (O_737,N_14276,N_14701);
and UO_738 (O_738,N_13534,N_14175);
xnor UO_739 (O_739,N_14703,N_14498);
xor UO_740 (O_740,N_13965,N_14760);
and UO_741 (O_741,N_13928,N_13813);
xor UO_742 (O_742,N_13541,N_13804);
xor UO_743 (O_743,N_14481,N_14933);
xnor UO_744 (O_744,N_13822,N_14629);
nand UO_745 (O_745,N_13742,N_14929);
and UO_746 (O_746,N_14808,N_13765);
or UO_747 (O_747,N_14767,N_14983);
nor UO_748 (O_748,N_13655,N_14582);
nand UO_749 (O_749,N_14089,N_14389);
nor UO_750 (O_750,N_14225,N_13579);
nor UO_751 (O_751,N_14190,N_13549);
nand UO_752 (O_752,N_14541,N_13674);
nor UO_753 (O_753,N_14962,N_14714);
nand UO_754 (O_754,N_13734,N_14727);
xnor UO_755 (O_755,N_13695,N_14709);
nand UO_756 (O_756,N_14490,N_14531);
xor UO_757 (O_757,N_13880,N_14158);
nand UO_758 (O_758,N_14012,N_14786);
nor UO_759 (O_759,N_14965,N_13764);
nand UO_760 (O_760,N_14709,N_14944);
nand UO_761 (O_761,N_13926,N_13521);
nor UO_762 (O_762,N_14190,N_14187);
and UO_763 (O_763,N_14209,N_14309);
nand UO_764 (O_764,N_13777,N_14513);
or UO_765 (O_765,N_14863,N_13770);
or UO_766 (O_766,N_14660,N_13974);
xor UO_767 (O_767,N_13718,N_14046);
nand UO_768 (O_768,N_14712,N_14203);
nor UO_769 (O_769,N_14938,N_14004);
or UO_770 (O_770,N_14700,N_13954);
and UO_771 (O_771,N_13820,N_13955);
xor UO_772 (O_772,N_13885,N_14713);
xor UO_773 (O_773,N_14077,N_14894);
xnor UO_774 (O_774,N_14404,N_14193);
nand UO_775 (O_775,N_14507,N_14535);
nor UO_776 (O_776,N_14387,N_14196);
or UO_777 (O_777,N_14104,N_14475);
nor UO_778 (O_778,N_14936,N_13811);
nand UO_779 (O_779,N_14425,N_14977);
nand UO_780 (O_780,N_14772,N_13639);
nor UO_781 (O_781,N_14243,N_13708);
or UO_782 (O_782,N_13549,N_13898);
or UO_783 (O_783,N_14400,N_14717);
or UO_784 (O_784,N_14371,N_13521);
xnor UO_785 (O_785,N_13626,N_14480);
nand UO_786 (O_786,N_14964,N_13660);
xnor UO_787 (O_787,N_14367,N_14245);
nand UO_788 (O_788,N_13773,N_13605);
nor UO_789 (O_789,N_14949,N_13666);
nor UO_790 (O_790,N_14825,N_13945);
nand UO_791 (O_791,N_13685,N_13910);
nand UO_792 (O_792,N_14798,N_14801);
and UO_793 (O_793,N_13955,N_14900);
nand UO_794 (O_794,N_14845,N_13712);
nand UO_795 (O_795,N_14927,N_13525);
nor UO_796 (O_796,N_14550,N_14325);
and UO_797 (O_797,N_14759,N_14424);
and UO_798 (O_798,N_13608,N_14578);
or UO_799 (O_799,N_14038,N_13590);
nor UO_800 (O_800,N_14207,N_13822);
nor UO_801 (O_801,N_14163,N_13642);
and UO_802 (O_802,N_13701,N_14201);
and UO_803 (O_803,N_14835,N_13952);
nor UO_804 (O_804,N_14963,N_13914);
nand UO_805 (O_805,N_14320,N_14971);
nor UO_806 (O_806,N_13874,N_14491);
and UO_807 (O_807,N_14002,N_13544);
nor UO_808 (O_808,N_14738,N_14814);
xnor UO_809 (O_809,N_14892,N_14017);
xor UO_810 (O_810,N_14954,N_13831);
nand UO_811 (O_811,N_14499,N_13527);
xnor UO_812 (O_812,N_14723,N_13561);
xor UO_813 (O_813,N_13721,N_13514);
nor UO_814 (O_814,N_13521,N_13860);
nand UO_815 (O_815,N_14032,N_13784);
xnor UO_816 (O_816,N_13929,N_13743);
or UO_817 (O_817,N_14454,N_14433);
nand UO_818 (O_818,N_13637,N_13605);
and UO_819 (O_819,N_14251,N_13964);
and UO_820 (O_820,N_14594,N_14926);
and UO_821 (O_821,N_14913,N_14019);
xor UO_822 (O_822,N_13908,N_14233);
xnor UO_823 (O_823,N_14364,N_13947);
nor UO_824 (O_824,N_13964,N_14963);
or UO_825 (O_825,N_14950,N_14951);
xnor UO_826 (O_826,N_13816,N_13807);
nand UO_827 (O_827,N_13979,N_14977);
nand UO_828 (O_828,N_13551,N_14567);
nor UO_829 (O_829,N_14648,N_13656);
or UO_830 (O_830,N_14302,N_14160);
nand UO_831 (O_831,N_13873,N_14595);
nor UO_832 (O_832,N_14095,N_14163);
nand UO_833 (O_833,N_14988,N_13660);
and UO_834 (O_834,N_14997,N_14749);
nand UO_835 (O_835,N_14978,N_13749);
nand UO_836 (O_836,N_14315,N_14855);
and UO_837 (O_837,N_13910,N_14901);
nand UO_838 (O_838,N_14263,N_14736);
nor UO_839 (O_839,N_13689,N_14498);
and UO_840 (O_840,N_14594,N_14374);
and UO_841 (O_841,N_14682,N_13693);
nor UO_842 (O_842,N_14461,N_13587);
or UO_843 (O_843,N_13882,N_13683);
and UO_844 (O_844,N_13896,N_13670);
or UO_845 (O_845,N_14384,N_13759);
nor UO_846 (O_846,N_14201,N_13933);
or UO_847 (O_847,N_14474,N_14047);
and UO_848 (O_848,N_14615,N_14372);
or UO_849 (O_849,N_14027,N_14149);
and UO_850 (O_850,N_14199,N_14782);
and UO_851 (O_851,N_14054,N_13912);
or UO_852 (O_852,N_14533,N_14225);
or UO_853 (O_853,N_13549,N_14001);
xor UO_854 (O_854,N_14053,N_14572);
xnor UO_855 (O_855,N_14928,N_14182);
or UO_856 (O_856,N_13803,N_14083);
nor UO_857 (O_857,N_13955,N_14071);
and UO_858 (O_858,N_13578,N_14747);
nand UO_859 (O_859,N_14186,N_13936);
nand UO_860 (O_860,N_14855,N_14348);
xnor UO_861 (O_861,N_13878,N_14868);
nand UO_862 (O_862,N_13696,N_14580);
and UO_863 (O_863,N_14991,N_14802);
nor UO_864 (O_864,N_14816,N_14927);
nor UO_865 (O_865,N_14287,N_13651);
nor UO_866 (O_866,N_14616,N_13946);
nor UO_867 (O_867,N_14449,N_14387);
or UO_868 (O_868,N_14598,N_14994);
nand UO_869 (O_869,N_14073,N_14891);
xor UO_870 (O_870,N_14843,N_14455);
nor UO_871 (O_871,N_13600,N_14157);
or UO_872 (O_872,N_13934,N_13962);
nand UO_873 (O_873,N_13732,N_14420);
nor UO_874 (O_874,N_14977,N_14165);
nor UO_875 (O_875,N_14711,N_14251);
xnor UO_876 (O_876,N_14759,N_14605);
xnor UO_877 (O_877,N_13719,N_14331);
or UO_878 (O_878,N_14548,N_14615);
nand UO_879 (O_879,N_14384,N_14066);
and UO_880 (O_880,N_13638,N_13865);
nand UO_881 (O_881,N_14015,N_13958);
and UO_882 (O_882,N_14907,N_14530);
nand UO_883 (O_883,N_14913,N_14125);
nor UO_884 (O_884,N_13677,N_14634);
xnor UO_885 (O_885,N_14189,N_14325);
and UO_886 (O_886,N_14891,N_13804);
nand UO_887 (O_887,N_14780,N_14638);
nor UO_888 (O_888,N_13769,N_13906);
nor UO_889 (O_889,N_13681,N_14741);
xnor UO_890 (O_890,N_14111,N_14569);
and UO_891 (O_891,N_13724,N_14971);
nor UO_892 (O_892,N_14211,N_13656);
nor UO_893 (O_893,N_14156,N_14039);
or UO_894 (O_894,N_13804,N_13572);
and UO_895 (O_895,N_13507,N_14316);
or UO_896 (O_896,N_14525,N_13586);
xnor UO_897 (O_897,N_14030,N_13556);
nand UO_898 (O_898,N_13786,N_13811);
or UO_899 (O_899,N_14886,N_13862);
and UO_900 (O_900,N_14692,N_14809);
or UO_901 (O_901,N_13845,N_14632);
and UO_902 (O_902,N_14968,N_14331);
or UO_903 (O_903,N_14967,N_13590);
and UO_904 (O_904,N_14365,N_14594);
or UO_905 (O_905,N_13530,N_14702);
nand UO_906 (O_906,N_14512,N_14399);
nand UO_907 (O_907,N_14546,N_14941);
or UO_908 (O_908,N_13918,N_14481);
nor UO_909 (O_909,N_13635,N_13813);
nand UO_910 (O_910,N_14642,N_14896);
nand UO_911 (O_911,N_13922,N_14985);
or UO_912 (O_912,N_14706,N_13920);
or UO_913 (O_913,N_14254,N_14597);
nand UO_914 (O_914,N_13824,N_13506);
or UO_915 (O_915,N_14319,N_13908);
nand UO_916 (O_916,N_14744,N_14069);
or UO_917 (O_917,N_13622,N_14805);
xor UO_918 (O_918,N_14151,N_14095);
nor UO_919 (O_919,N_14468,N_14541);
and UO_920 (O_920,N_14312,N_14549);
nand UO_921 (O_921,N_13838,N_14843);
or UO_922 (O_922,N_14318,N_14025);
and UO_923 (O_923,N_13757,N_14395);
and UO_924 (O_924,N_13827,N_14706);
nand UO_925 (O_925,N_14563,N_14227);
nand UO_926 (O_926,N_14600,N_13844);
xnor UO_927 (O_927,N_14408,N_14863);
nor UO_928 (O_928,N_14176,N_13674);
xor UO_929 (O_929,N_14772,N_13868);
nand UO_930 (O_930,N_14664,N_14506);
or UO_931 (O_931,N_13914,N_14405);
xnor UO_932 (O_932,N_14949,N_13501);
nor UO_933 (O_933,N_13828,N_14552);
xnor UO_934 (O_934,N_14915,N_14260);
nor UO_935 (O_935,N_14904,N_13767);
and UO_936 (O_936,N_14184,N_14388);
xnor UO_937 (O_937,N_14179,N_14801);
xor UO_938 (O_938,N_14099,N_14461);
and UO_939 (O_939,N_13557,N_14049);
nand UO_940 (O_940,N_13710,N_14052);
and UO_941 (O_941,N_13793,N_14809);
nor UO_942 (O_942,N_13955,N_13554);
nor UO_943 (O_943,N_13932,N_14180);
or UO_944 (O_944,N_13705,N_14736);
nand UO_945 (O_945,N_14092,N_14731);
xnor UO_946 (O_946,N_13528,N_13851);
nand UO_947 (O_947,N_14790,N_14546);
and UO_948 (O_948,N_14420,N_14462);
xor UO_949 (O_949,N_14204,N_13523);
or UO_950 (O_950,N_13731,N_13894);
nor UO_951 (O_951,N_13572,N_13705);
and UO_952 (O_952,N_14252,N_14612);
nand UO_953 (O_953,N_13934,N_13615);
and UO_954 (O_954,N_13721,N_13572);
xnor UO_955 (O_955,N_13690,N_14652);
nor UO_956 (O_956,N_14433,N_14412);
nor UO_957 (O_957,N_13624,N_14060);
nor UO_958 (O_958,N_13641,N_13735);
nor UO_959 (O_959,N_14552,N_14879);
and UO_960 (O_960,N_14864,N_14828);
xor UO_961 (O_961,N_13793,N_14986);
and UO_962 (O_962,N_14501,N_13559);
xnor UO_963 (O_963,N_14807,N_14610);
nor UO_964 (O_964,N_14801,N_13539);
and UO_965 (O_965,N_13721,N_14248);
nor UO_966 (O_966,N_14471,N_14419);
nor UO_967 (O_967,N_14986,N_14513);
or UO_968 (O_968,N_13985,N_13626);
nand UO_969 (O_969,N_14249,N_14148);
nor UO_970 (O_970,N_13723,N_13600);
or UO_971 (O_971,N_13985,N_13769);
xor UO_972 (O_972,N_14504,N_13701);
xnor UO_973 (O_973,N_13813,N_13839);
nand UO_974 (O_974,N_14569,N_14604);
and UO_975 (O_975,N_14478,N_13569);
nor UO_976 (O_976,N_13855,N_14334);
nand UO_977 (O_977,N_14463,N_14963);
xor UO_978 (O_978,N_14332,N_13624);
and UO_979 (O_979,N_13743,N_14073);
nand UO_980 (O_980,N_14660,N_14393);
xor UO_981 (O_981,N_13690,N_13718);
nand UO_982 (O_982,N_13711,N_14942);
and UO_983 (O_983,N_14447,N_14415);
or UO_984 (O_984,N_14456,N_14885);
or UO_985 (O_985,N_13613,N_14340);
nand UO_986 (O_986,N_14071,N_13837);
nand UO_987 (O_987,N_14467,N_13872);
or UO_988 (O_988,N_14766,N_13946);
or UO_989 (O_989,N_14828,N_14208);
nor UO_990 (O_990,N_13774,N_13819);
nand UO_991 (O_991,N_13729,N_14884);
nor UO_992 (O_992,N_14750,N_14965);
nand UO_993 (O_993,N_14983,N_14804);
and UO_994 (O_994,N_14866,N_14659);
xor UO_995 (O_995,N_13654,N_14140);
or UO_996 (O_996,N_13965,N_14889);
xnor UO_997 (O_997,N_14686,N_14866);
nand UO_998 (O_998,N_14947,N_13502);
and UO_999 (O_999,N_14708,N_13674);
or UO_1000 (O_1000,N_14025,N_14498);
xor UO_1001 (O_1001,N_14568,N_14533);
or UO_1002 (O_1002,N_14012,N_13941);
or UO_1003 (O_1003,N_14443,N_14163);
or UO_1004 (O_1004,N_13555,N_14326);
nor UO_1005 (O_1005,N_14056,N_13934);
nand UO_1006 (O_1006,N_14223,N_14255);
xor UO_1007 (O_1007,N_14273,N_14061);
nand UO_1008 (O_1008,N_14078,N_13539);
or UO_1009 (O_1009,N_14519,N_13537);
nand UO_1010 (O_1010,N_14670,N_14520);
nor UO_1011 (O_1011,N_14086,N_14349);
or UO_1012 (O_1012,N_14058,N_14283);
xor UO_1013 (O_1013,N_14567,N_13936);
or UO_1014 (O_1014,N_14541,N_14214);
xnor UO_1015 (O_1015,N_13865,N_13693);
xor UO_1016 (O_1016,N_14985,N_14241);
xor UO_1017 (O_1017,N_14299,N_14567);
nor UO_1018 (O_1018,N_14362,N_14012);
or UO_1019 (O_1019,N_14286,N_14670);
and UO_1020 (O_1020,N_14973,N_14168);
nor UO_1021 (O_1021,N_14710,N_13880);
and UO_1022 (O_1022,N_13914,N_14020);
nor UO_1023 (O_1023,N_13576,N_14769);
xnor UO_1024 (O_1024,N_14154,N_14621);
xor UO_1025 (O_1025,N_14887,N_14868);
xnor UO_1026 (O_1026,N_14962,N_14641);
and UO_1027 (O_1027,N_14655,N_13763);
xor UO_1028 (O_1028,N_14945,N_14540);
nor UO_1029 (O_1029,N_14320,N_14983);
xnor UO_1030 (O_1030,N_13752,N_13820);
and UO_1031 (O_1031,N_13685,N_14510);
nor UO_1032 (O_1032,N_14091,N_13619);
nand UO_1033 (O_1033,N_14982,N_13777);
nand UO_1034 (O_1034,N_14143,N_13949);
and UO_1035 (O_1035,N_13665,N_14273);
nor UO_1036 (O_1036,N_13804,N_13995);
nand UO_1037 (O_1037,N_14049,N_14587);
xor UO_1038 (O_1038,N_13754,N_14915);
nand UO_1039 (O_1039,N_13866,N_13618);
or UO_1040 (O_1040,N_14799,N_14037);
or UO_1041 (O_1041,N_14359,N_14136);
nor UO_1042 (O_1042,N_13705,N_14201);
nor UO_1043 (O_1043,N_14231,N_14087);
or UO_1044 (O_1044,N_14160,N_14244);
xor UO_1045 (O_1045,N_14555,N_14663);
or UO_1046 (O_1046,N_13965,N_14932);
and UO_1047 (O_1047,N_13970,N_14452);
and UO_1048 (O_1048,N_13762,N_14276);
nor UO_1049 (O_1049,N_14937,N_14940);
nor UO_1050 (O_1050,N_14827,N_14398);
xnor UO_1051 (O_1051,N_14175,N_14262);
or UO_1052 (O_1052,N_14402,N_13897);
xor UO_1053 (O_1053,N_13546,N_14943);
or UO_1054 (O_1054,N_14593,N_14564);
xor UO_1055 (O_1055,N_13585,N_14139);
nand UO_1056 (O_1056,N_13608,N_14756);
or UO_1057 (O_1057,N_13554,N_13537);
nand UO_1058 (O_1058,N_14137,N_13572);
nand UO_1059 (O_1059,N_14961,N_14791);
and UO_1060 (O_1060,N_14684,N_13734);
nand UO_1061 (O_1061,N_14349,N_14747);
nand UO_1062 (O_1062,N_13843,N_13568);
nor UO_1063 (O_1063,N_13571,N_13964);
nor UO_1064 (O_1064,N_14287,N_14046);
xor UO_1065 (O_1065,N_13837,N_14823);
xnor UO_1066 (O_1066,N_14266,N_14374);
nor UO_1067 (O_1067,N_14215,N_13751);
xnor UO_1068 (O_1068,N_13642,N_13722);
nand UO_1069 (O_1069,N_13509,N_14714);
and UO_1070 (O_1070,N_14731,N_13897);
or UO_1071 (O_1071,N_14142,N_14806);
nor UO_1072 (O_1072,N_14626,N_14347);
nand UO_1073 (O_1073,N_13893,N_14175);
or UO_1074 (O_1074,N_13829,N_14470);
and UO_1075 (O_1075,N_13907,N_13506);
xor UO_1076 (O_1076,N_14525,N_13850);
xor UO_1077 (O_1077,N_13986,N_14055);
or UO_1078 (O_1078,N_14284,N_13951);
or UO_1079 (O_1079,N_14792,N_14259);
nor UO_1080 (O_1080,N_13742,N_13603);
or UO_1081 (O_1081,N_13751,N_13889);
nor UO_1082 (O_1082,N_13916,N_13806);
or UO_1083 (O_1083,N_13977,N_13622);
nor UO_1084 (O_1084,N_14065,N_14313);
nor UO_1085 (O_1085,N_13827,N_14540);
or UO_1086 (O_1086,N_13740,N_14938);
nand UO_1087 (O_1087,N_14482,N_14684);
nor UO_1088 (O_1088,N_14759,N_14918);
nand UO_1089 (O_1089,N_14621,N_14490);
or UO_1090 (O_1090,N_13641,N_14878);
nand UO_1091 (O_1091,N_14525,N_14790);
xnor UO_1092 (O_1092,N_13551,N_14751);
xor UO_1093 (O_1093,N_14539,N_13787);
nand UO_1094 (O_1094,N_14533,N_14646);
nor UO_1095 (O_1095,N_14669,N_14537);
nor UO_1096 (O_1096,N_13712,N_14691);
nand UO_1097 (O_1097,N_13683,N_14419);
nor UO_1098 (O_1098,N_13751,N_14612);
or UO_1099 (O_1099,N_14584,N_13694);
and UO_1100 (O_1100,N_13501,N_14069);
xor UO_1101 (O_1101,N_14769,N_14586);
xnor UO_1102 (O_1102,N_14237,N_13573);
nor UO_1103 (O_1103,N_13601,N_13874);
nor UO_1104 (O_1104,N_13521,N_14566);
and UO_1105 (O_1105,N_14285,N_14012);
or UO_1106 (O_1106,N_14734,N_14451);
xor UO_1107 (O_1107,N_13669,N_14769);
nand UO_1108 (O_1108,N_13578,N_14144);
nor UO_1109 (O_1109,N_13974,N_14038);
nor UO_1110 (O_1110,N_13808,N_14899);
nand UO_1111 (O_1111,N_13960,N_14329);
and UO_1112 (O_1112,N_13995,N_13706);
or UO_1113 (O_1113,N_13977,N_13940);
and UO_1114 (O_1114,N_14491,N_14929);
xnor UO_1115 (O_1115,N_14105,N_14632);
nor UO_1116 (O_1116,N_14106,N_13974);
nor UO_1117 (O_1117,N_13901,N_14458);
or UO_1118 (O_1118,N_14719,N_14705);
xor UO_1119 (O_1119,N_14430,N_13627);
or UO_1120 (O_1120,N_14584,N_14907);
or UO_1121 (O_1121,N_14833,N_14071);
nand UO_1122 (O_1122,N_14531,N_13670);
and UO_1123 (O_1123,N_14957,N_14454);
or UO_1124 (O_1124,N_13843,N_13545);
nor UO_1125 (O_1125,N_14208,N_14574);
nor UO_1126 (O_1126,N_14219,N_14952);
or UO_1127 (O_1127,N_14782,N_13814);
and UO_1128 (O_1128,N_14334,N_13795);
xnor UO_1129 (O_1129,N_14246,N_14444);
xnor UO_1130 (O_1130,N_14162,N_13848);
and UO_1131 (O_1131,N_14530,N_14702);
nor UO_1132 (O_1132,N_14647,N_14184);
and UO_1133 (O_1133,N_14030,N_14503);
or UO_1134 (O_1134,N_13587,N_14675);
or UO_1135 (O_1135,N_14758,N_14553);
xnor UO_1136 (O_1136,N_14862,N_13844);
nand UO_1137 (O_1137,N_14597,N_14615);
nor UO_1138 (O_1138,N_13604,N_14551);
nand UO_1139 (O_1139,N_13522,N_13749);
nor UO_1140 (O_1140,N_14255,N_14163);
and UO_1141 (O_1141,N_13721,N_14953);
nand UO_1142 (O_1142,N_13565,N_14220);
or UO_1143 (O_1143,N_14808,N_14019);
nor UO_1144 (O_1144,N_14106,N_13808);
or UO_1145 (O_1145,N_13968,N_14864);
xor UO_1146 (O_1146,N_13594,N_14085);
xor UO_1147 (O_1147,N_13736,N_13770);
xnor UO_1148 (O_1148,N_13607,N_13983);
nand UO_1149 (O_1149,N_14574,N_14775);
xor UO_1150 (O_1150,N_13955,N_14808);
or UO_1151 (O_1151,N_14576,N_14230);
and UO_1152 (O_1152,N_14774,N_13919);
xnor UO_1153 (O_1153,N_14966,N_14311);
xor UO_1154 (O_1154,N_14960,N_13642);
nor UO_1155 (O_1155,N_13995,N_14142);
nand UO_1156 (O_1156,N_13611,N_14430);
nor UO_1157 (O_1157,N_13887,N_13832);
xnor UO_1158 (O_1158,N_14702,N_14050);
and UO_1159 (O_1159,N_14821,N_13741);
and UO_1160 (O_1160,N_13806,N_14120);
and UO_1161 (O_1161,N_14889,N_13996);
or UO_1162 (O_1162,N_14530,N_14022);
xnor UO_1163 (O_1163,N_13812,N_13700);
and UO_1164 (O_1164,N_14788,N_14443);
nor UO_1165 (O_1165,N_13503,N_14514);
and UO_1166 (O_1166,N_13588,N_14157);
xnor UO_1167 (O_1167,N_14522,N_14402);
or UO_1168 (O_1168,N_13627,N_14131);
or UO_1169 (O_1169,N_13626,N_14446);
or UO_1170 (O_1170,N_13904,N_14325);
xnor UO_1171 (O_1171,N_13934,N_14246);
or UO_1172 (O_1172,N_14557,N_14872);
or UO_1173 (O_1173,N_13834,N_14399);
xor UO_1174 (O_1174,N_14433,N_14051);
nand UO_1175 (O_1175,N_14269,N_14826);
or UO_1176 (O_1176,N_13702,N_14851);
or UO_1177 (O_1177,N_13807,N_14294);
xor UO_1178 (O_1178,N_13960,N_14263);
nand UO_1179 (O_1179,N_14966,N_13983);
xor UO_1180 (O_1180,N_14773,N_14769);
xnor UO_1181 (O_1181,N_14233,N_13909);
xnor UO_1182 (O_1182,N_13878,N_14168);
and UO_1183 (O_1183,N_14003,N_13721);
nand UO_1184 (O_1184,N_14222,N_14034);
nand UO_1185 (O_1185,N_14429,N_13628);
xor UO_1186 (O_1186,N_13708,N_14194);
nand UO_1187 (O_1187,N_14927,N_14480);
and UO_1188 (O_1188,N_14705,N_14400);
nor UO_1189 (O_1189,N_14425,N_13969);
nand UO_1190 (O_1190,N_13811,N_14257);
nor UO_1191 (O_1191,N_14313,N_14363);
or UO_1192 (O_1192,N_14729,N_14624);
or UO_1193 (O_1193,N_14263,N_14004);
or UO_1194 (O_1194,N_13910,N_13586);
nand UO_1195 (O_1195,N_13567,N_14862);
xnor UO_1196 (O_1196,N_14918,N_14846);
nor UO_1197 (O_1197,N_13888,N_13892);
or UO_1198 (O_1198,N_14033,N_14023);
and UO_1199 (O_1199,N_14671,N_14517);
nor UO_1200 (O_1200,N_14108,N_14713);
and UO_1201 (O_1201,N_14113,N_14910);
nor UO_1202 (O_1202,N_14670,N_14220);
and UO_1203 (O_1203,N_14841,N_14017);
nor UO_1204 (O_1204,N_13641,N_13890);
xnor UO_1205 (O_1205,N_13807,N_13744);
nand UO_1206 (O_1206,N_13839,N_14755);
xnor UO_1207 (O_1207,N_13889,N_13958);
and UO_1208 (O_1208,N_14155,N_13937);
and UO_1209 (O_1209,N_14220,N_14210);
or UO_1210 (O_1210,N_14976,N_13836);
xnor UO_1211 (O_1211,N_13751,N_13575);
nor UO_1212 (O_1212,N_14384,N_14065);
xor UO_1213 (O_1213,N_14729,N_13519);
nand UO_1214 (O_1214,N_13717,N_14448);
nor UO_1215 (O_1215,N_14442,N_14223);
xnor UO_1216 (O_1216,N_14440,N_13878);
xnor UO_1217 (O_1217,N_13957,N_14022);
nor UO_1218 (O_1218,N_14478,N_13635);
and UO_1219 (O_1219,N_14081,N_14061);
or UO_1220 (O_1220,N_14142,N_14391);
nand UO_1221 (O_1221,N_13662,N_14634);
or UO_1222 (O_1222,N_14022,N_13819);
nand UO_1223 (O_1223,N_14191,N_13681);
xor UO_1224 (O_1224,N_14100,N_13857);
and UO_1225 (O_1225,N_13857,N_14049);
or UO_1226 (O_1226,N_14093,N_14370);
and UO_1227 (O_1227,N_14175,N_14868);
nand UO_1228 (O_1228,N_13536,N_14212);
or UO_1229 (O_1229,N_14226,N_14663);
nor UO_1230 (O_1230,N_14331,N_14565);
nor UO_1231 (O_1231,N_14017,N_14521);
nor UO_1232 (O_1232,N_14576,N_14850);
nand UO_1233 (O_1233,N_14339,N_14177);
xor UO_1234 (O_1234,N_14280,N_14854);
or UO_1235 (O_1235,N_13721,N_13752);
and UO_1236 (O_1236,N_14591,N_13598);
and UO_1237 (O_1237,N_14448,N_13584);
or UO_1238 (O_1238,N_14820,N_14770);
nor UO_1239 (O_1239,N_14744,N_14908);
nand UO_1240 (O_1240,N_14774,N_14869);
nand UO_1241 (O_1241,N_13899,N_14161);
nor UO_1242 (O_1242,N_13772,N_13978);
and UO_1243 (O_1243,N_13776,N_13522);
and UO_1244 (O_1244,N_14853,N_14904);
and UO_1245 (O_1245,N_14909,N_14223);
and UO_1246 (O_1246,N_13630,N_13928);
and UO_1247 (O_1247,N_14083,N_13820);
nor UO_1248 (O_1248,N_14368,N_14125);
or UO_1249 (O_1249,N_13614,N_14387);
and UO_1250 (O_1250,N_14679,N_14265);
nand UO_1251 (O_1251,N_14604,N_14201);
and UO_1252 (O_1252,N_13985,N_13679);
and UO_1253 (O_1253,N_14799,N_14984);
nand UO_1254 (O_1254,N_14088,N_14111);
or UO_1255 (O_1255,N_14845,N_14906);
and UO_1256 (O_1256,N_14182,N_13666);
and UO_1257 (O_1257,N_14241,N_13789);
nand UO_1258 (O_1258,N_14603,N_14480);
xnor UO_1259 (O_1259,N_13689,N_14586);
or UO_1260 (O_1260,N_14344,N_14718);
xnor UO_1261 (O_1261,N_14276,N_13993);
xnor UO_1262 (O_1262,N_13971,N_14632);
or UO_1263 (O_1263,N_14669,N_14116);
xor UO_1264 (O_1264,N_14896,N_14581);
xor UO_1265 (O_1265,N_14582,N_13765);
and UO_1266 (O_1266,N_14164,N_14967);
or UO_1267 (O_1267,N_13841,N_14544);
nor UO_1268 (O_1268,N_14729,N_14798);
xnor UO_1269 (O_1269,N_13554,N_14451);
nor UO_1270 (O_1270,N_14201,N_13668);
xor UO_1271 (O_1271,N_14713,N_13712);
nor UO_1272 (O_1272,N_13597,N_14594);
xor UO_1273 (O_1273,N_14140,N_13945);
xor UO_1274 (O_1274,N_14969,N_14237);
and UO_1275 (O_1275,N_13625,N_14488);
nor UO_1276 (O_1276,N_14826,N_14589);
and UO_1277 (O_1277,N_14074,N_14786);
and UO_1278 (O_1278,N_14781,N_13627);
and UO_1279 (O_1279,N_14015,N_14472);
or UO_1280 (O_1280,N_14774,N_13530);
xor UO_1281 (O_1281,N_14939,N_13936);
and UO_1282 (O_1282,N_14349,N_14843);
or UO_1283 (O_1283,N_14030,N_14501);
and UO_1284 (O_1284,N_14046,N_13706);
or UO_1285 (O_1285,N_14745,N_14525);
nor UO_1286 (O_1286,N_14635,N_14404);
and UO_1287 (O_1287,N_13732,N_14038);
nor UO_1288 (O_1288,N_14105,N_13943);
nand UO_1289 (O_1289,N_14576,N_14740);
and UO_1290 (O_1290,N_13731,N_14464);
nand UO_1291 (O_1291,N_14562,N_14781);
xnor UO_1292 (O_1292,N_14007,N_14196);
and UO_1293 (O_1293,N_14633,N_14541);
nand UO_1294 (O_1294,N_14754,N_14321);
and UO_1295 (O_1295,N_13868,N_13796);
xor UO_1296 (O_1296,N_13594,N_14043);
and UO_1297 (O_1297,N_13875,N_14340);
xnor UO_1298 (O_1298,N_13817,N_14469);
and UO_1299 (O_1299,N_14340,N_14216);
and UO_1300 (O_1300,N_13648,N_14004);
or UO_1301 (O_1301,N_14725,N_13606);
or UO_1302 (O_1302,N_14776,N_13895);
nor UO_1303 (O_1303,N_14431,N_14470);
nand UO_1304 (O_1304,N_14219,N_14190);
and UO_1305 (O_1305,N_13603,N_13761);
nand UO_1306 (O_1306,N_14572,N_14379);
and UO_1307 (O_1307,N_14185,N_14152);
xor UO_1308 (O_1308,N_13596,N_14960);
xor UO_1309 (O_1309,N_13675,N_13803);
xnor UO_1310 (O_1310,N_13878,N_13549);
or UO_1311 (O_1311,N_14122,N_14774);
nand UO_1312 (O_1312,N_14576,N_14296);
and UO_1313 (O_1313,N_14978,N_14533);
nor UO_1314 (O_1314,N_13642,N_14178);
nor UO_1315 (O_1315,N_14022,N_13697);
and UO_1316 (O_1316,N_14305,N_13977);
and UO_1317 (O_1317,N_14336,N_13731);
xnor UO_1318 (O_1318,N_13979,N_14914);
xnor UO_1319 (O_1319,N_14792,N_14838);
nand UO_1320 (O_1320,N_14611,N_14201);
nor UO_1321 (O_1321,N_14531,N_13552);
xor UO_1322 (O_1322,N_14074,N_14741);
xnor UO_1323 (O_1323,N_14139,N_13557);
nor UO_1324 (O_1324,N_14479,N_14580);
nor UO_1325 (O_1325,N_14053,N_13591);
nand UO_1326 (O_1326,N_14069,N_14987);
nand UO_1327 (O_1327,N_14603,N_14103);
nand UO_1328 (O_1328,N_13723,N_14197);
or UO_1329 (O_1329,N_13791,N_13784);
nand UO_1330 (O_1330,N_14986,N_14630);
xor UO_1331 (O_1331,N_14714,N_13826);
nand UO_1332 (O_1332,N_14200,N_14284);
nor UO_1333 (O_1333,N_14375,N_14349);
and UO_1334 (O_1334,N_14863,N_13656);
and UO_1335 (O_1335,N_14580,N_14926);
or UO_1336 (O_1336,N_14303,N_14776);
or UO_1337 (O_1337,N_13812,N_13982);
xor UO_1338 (O_1338,N_13505,N_14090);
nor UO_1339 (O_1339,N_14560,N_14410);
nand UO_1340 (O_1340,N_14096,N_14076);
and UO_1341 (O_1341,N_14556,N_13975);
xor UO_1342 (O_1342,N_14093,N_14660);
nand UO_1343 (O_1343,N_14675,N_13772);
or UO_1344 (O_1344,N_14221,N_14813);
xnor UO_1345 (O_1345,N_13677,N_14919);
xnor UO_1346 (O_1346,N_13907,N_14306);
nor UO_1347 (O_1347,N_14223,N_14080);
nor UO_1348 (O_1348,N_14581,N_13673);
and UO_1349 (O_1349,N_14661,N_14849);
nand UO_1350 (O_1350,N_14693,N_14558);
or UO_1351 (O_1351,N_14198,N_14149);
xnor UO_1352 (O_1352,N_14891,N_13649);
nand UO_1353 (O_1353,N_13943,N_14249);
nand UO_1354 (O_1354,N_13932,N_13704);
nand UO_1355 (O_1355,N_14677,N_13910);
and UO_1356 (O_1356,N_13690,N_13549);
or UO_1357 (O_1357,N_14836,N_14366);
nand UO_1358 (O_1358,N_14681,N_14574);
or UO_1359 (O_1359,N_14992,N_14441);
nor UO_1360 (O_1360,N_14289,N_13629);
nor UO_1361 (O_1361,N_14459,N_14225);
and UO_1362 (O_1362,N_14073,N_13903);
and UO_1363 (O_1363,N_13801,N_14062);
nand UO_1364 (O_1364,N_14936,N_13842);
nor UO_1365 (O_1365,N_14028,N_14811);
xnor UO_1366 (O_1366,N_14019,N_14633);
or UO_1367 (O_1367,N_14848,N_14539);
and UO_1368 (O_1368,N_13970,N_14932);
xnor UO_1369 (O_1369,N_14808,N_14332);
nand UO_1370 (O_1370,N_14257,N_14099);
nor UO_1371 (O_1371,N_14183,N_14334);
or UO_1372 (O_1372,N_14870,N_14726);
nand UO_1373 (O_1373,N_14888,N_13824);
nor UO_1374 (O_1374,N_14529,N_14177);
or UO_1375 (O_1375,N_14466,N_13643);
nor UO_1376 (O_1376,N_13959,N_14906);
xnor UO_1377 (O_1377,N_14308,N_14185);
nand UO_1378 (O_1378,N_14240,N_14380);
nor UO_1379 (O_1379,N_14546,N_14931);
nor UO_1380 (O_1380,N_14810,N_14705);
nor UO_1381 (O_1381,N_13820,N_14816);
or UO_1382 (O_1382,N_14425,N_14835);
xnor UO_1383 (O_1383,N_14583,N_14489);
nand UO_1384 (O_1384,N_14728,N_13984);
nand UO_1385 (O_1385,N_14260,N_14612);
nand UO_1386 (O_1386,N_14955,N_13853);
xor UO_1387 (O_1387,N_13982,N_14921);
or UO_1388 (O_1388,N_14944,N_14224);
xnor UO_1389 (O_1389,N_14033,N_13903);
nor UO_1390 (O_1390,N_14295,N_13586);
xnor UO_1391 (O_1391,N_14707,N_14156);
nand UO_1392 (O_1392,N_13956,N_14080);
and UO_1393 (O_1393,N_13715,N_14329);
xnor UO_1394 (O_1394,N_14010,N_13797);
nor UO_1395 (O_1395,N_14529,N_14094);
xnor UO_1396 (O_1396,N_13630,N_14826);
xnor UO_1397 (O_1397,N_13666,N_13932);
and UO_1398 (O_1398,N_13553,N_14387);
xor UO_1399 (O_1399,N_14416,N_13608);
and UO_1400 (O_1400,N_14315,N_14767);
xnor UO_1401 (O_1401,N_14408,N_13624);
or UO_1402 (O_1402,N_13934,N_14583);
xor UO_1403 (O_1403,N_13878,N_14930);
nand UO_1404 (O_1404,N_13649,N_14402);
nand UO_1405 (O_1405,N_14888,N_13918);
and UO_1406 (O_1406,N_13506,N_14057);
or UO_1407 (O_1407,N_13622,N_14345);
nor UO_1408 (O_1408,N_14336,N_14941);
and UO_1409 (O_1409,N_14511,N_14418);
xnor UO_1410 (O_1410,N_14880,N_14423);
nand UO_1411 (O_1411,N_14661,N_14552);
nor UO_1412 (O_1412,N_14446,N_14941);
xnor UO_1413 (O_1413,N_14161,N_13781);
or UO_1414 (O_1414,N_14166,N_14422);
nand UO_1415 (O_1415,N_14543,N_14715);
or UO_1416 (O_1416,N_14511,N_14225);
or UO_1417 (O_1417,N_14061,N_14229);
nor UO_1418 (O_1418,N_13581,N_14559);
nand UO_1419 (O_1419,N_14183,N_13821);
nor UO_1420 (O_1420,N_14478,N_14610);
and UO_1421 (O_1421,N_13943,N_13935);
xnor UO_1422 (O_1422,N_14471,N_14325);
xnor UO_1423 (O_1423,N_13724,N_14562);
or UO_1424 (O_1424,N_14886,N_13568);
xor UO_1425 (O_1425,N_14029,N_13622);
nand UO_1426 (O_1426,N_13815,N_13949);
xor UO_1427 (O_1427,N_13601,N_13604);
and UO_1428 (O_1428,N_14036,N_14765);
or UO_1429 (O_1429,N_13767,N_14064);
nand UO_1430 (O_1430,N_14129,N_14844);
xnor UO_1431 (O_1431,N_13699,N_14346);
nand UO_1432 (O_1432,N_13771,N_13819);
and UO_1433 (O_1433,N_14504,N_14506);
and UO_1434 (O_1434,N_14096,N_13818);
nor UO_1435 (O_1435,N_14608,N_13699);
and UO_1436 (O_1436,N_14736,N_13622);
or UO_1437 (O_1437,N_14455,N_13826);
xnor UO_1438 (O_1438,N_14130,N_13941);
or UO_1439 (O_1439,N_14049,N_14668);
nand UO_1440 (O_1440,N_14907,N_14688);
and UO_1441 (O_1441,N_14346,N_13980);
nor UO_1442 (O_1442,N_14275,N_14954);
xor UO_1443 (O_1443,N_14220,N_14437);
xor UO_1444 (O_1444,N_14997,N_14398);
nand UO_1445 (O_1445,N_13962,N_14183);
nand UO_1446 (O_1446,N_14590,N_14655);
nor UO_1447 (O_1447,N_14502,N_14433);
nand UO_1448 (O_1448,N_14166,N_14698);
and UO_1449 (O_1449,N_13893,N_13517);
nand UO_1450 (O_1450,N_14215,N_13875);
nor UO_1451 (O_1451,N_14236,N_14258);
xor UO_1452 (O_1452,N_14532,N_13784);
or UO_1453 (O_1453,N_14089,N_13545);
or UO_1454 (O_1454,N_14393,N_14740);
nand UO_1455 (O_1455,N_13908,N_13829);
xnor UO_1456 (O_1456,N_13679,N_13916);
xnor UO_1457 (O_1457,N_14700,N_14932);
or UO_1458 (O_1458,N_13771,N_14135);
and UO_1459 (O_1459,N_14201,N_13501);
or UO_1460 (O_1460,N_13973,N_14148);
or UO_1461 (O_1461,N_14809,N_13711);
nor UO_1462 (O_1462,N_14683,N_13974);
or UO_1463 (O_1463,N_14244,N_13856);
and UO_1464 (O_1464,N_14055,N_13647);
nor UO_1465 (O_1465,N_13729,N_14273);
xor UO_1466 (O_1466,N_14978,N_14259);
xor UO_1467 (O_1467,N_14278,N_13780);
and UO_1468 (O_1468,N_14247,N_14708);
xnor UO_1469 (O_1469,N_13783,N_14391);
and UO_1470 (O_1470,N_14889,N_14170);
nand UO_1471 (O_1471,N_14280,N_13821);
nand UO_1472 (O_1472,N_14069,N_14696);
xor UO_1473 (O_1473,N_13706,N_14306);
nand UO_1474 (O_1474,N_14538,N_14009);
nor UO_1475 (O_1475,N_14895,N_14579);
nor UO_1476 (O_1476,N_14054,N_14731);
and UO_1477 (O_1477,N_14428,N_14296);
or UO_1478 (O_1478,N_14731,N_14057);
nand UO_1479 (O_1479,N_14956,N_14391);
nand UO_1480 (O_1480,N_14388,N_13972);
and UO_1481 (O_1481,N_14557,N_14354);
xnor UO_1482 (O_1482,N_14498,N_14628);
nand UO_1483 (O_1483,N_14492,N_13858);
or UO_1484 (O_1484,N_14887,N_14541);
or UO_1485 (O_1485,N_14875,N_14320);
nand UO_1486 (O_1486,N_14533,N_14157);
nor UO_1487 (O_1487,N_13627,N_14188);
and UO_1488 (O_1488,N_14054,N_14962);
and UO_1489 (O_1489,N_14965,N_14271);
nor UO_1490 (O_1490,N_14765,N_13884);
and UO_1491 (O_1491,N_13884,N_13785);
or UO_1492 (O_1492,N_14674,N_14773);
nor UO_1493 (O_1493,N_14360,N_13671);
nor UO_1494 (O_1494,N_13935,N_13714);
or UO_1495 (O_1495,N_13845,N_13836);
xnor UO_1496 (O_1496,N_14995,N_13505);
and UO_1497 (O_1497,N_14324,N_13889);
xnor UO_1498 (O_1498,N_14873,N_14453);
xor UO_1499 (O_1499,N_14350,N_13757);
nor UO_1500 (O_1500,N_14984,N_14913);
and UO_1501 (O_1501,N_14539,N_13584);
nor UO_1502 (O_1502,N_13925,N_14818);
nand UO_1503 (O_1503,N_14865,N_14736);
nand UO_1504 (O_1504,N_14618,N_13714);
nor UO_1505 (O_1505,N_14069,N_14476);
xor UO_1506 (O_1506,N_13721,N_14347);
nand UO_1507 (O_1507,N_14167,N_14530);
nand UO_1508 (O_1508,N_14548,N_13762);
nor UO_1509 (O_1509,N_14123,N_14944);
or UO_1510 (O_1510,N_14211,N_14034);
xnor UO_1511 (O_1511,N_13555,N_13884);
or UO_1512 (O_1512,N_14868,N_13781);
nand UO_1513 (O_1513,N_14481,N_14769);
or UO_1514 (O_1514,N_14149,N_13972);
and UO_1515 (O_1515,N_14502,N_14033);
xnor UO_1516 (O_1516,N_14588,N_14490);
nor UO_1517 (O_1517,N_14549,N_14114);
nand UO_1518 (O_1518,N_14035,N_14262);
and UO_1519 (O_1519,N_14261,N_14826);
nor UO_1520 (O_1520,N_14464,N_14721);
and UO_1521 (O_1521,N_14241,N_13646);
and UO_1522 (O_1522,N_14658,N_14464);
or UO_1523 (O_1523,N_13803,N_13962);
or UO_1524 (O_1524,N_14008,N_14529);
nand UO_1525 (O_1525,N_14187,N_14873);
nor UO_1526 (O_1526,N_14016,N_14359);
or UO_1527 (O_1527,N_14100,N_14952);
nor UO_1528 (O_1528,N_13615,N_14185);
nor UO_1529 (O_1529,N_14848,N_14732);
nand UO_1530 (O_1530,N_14371,N_13821);
and UO_1531 (O_1531,N_13919,N_13788);
nand UO_1532 (O_1532,N_13640,N_13845);
nand UO_1533 (O_1533,N_14214,N_14412);
or UO_1534 (O_1534,N_14968,N_14812);
xor UO_1535 (O_1535,N_14985,N_13690);
nand UO_1536 (O_1536,N_14735,N_14465);
nor UO_1537 (O_1537,N_14176,N_14692);
and UO_1538 (O_1538,N_14511,N_14966);
nand UO_1539 (O_1539,N_14711,N_14787);
nor UO_1540 (O_1540,N_13604,N_14540);
and UO_1541 (O_1541,N_14019,N_13792);
nor UO_1542 (O_1542,N_13791,N_13792);
xor UO_1543 (O_1543,N_13990,N_14434);
xor UO_1544 (O_1544,N_14814,N_14030);
nand UO_1545 (O_1545,N_14912,N_14943);
nor UO_1546 (O_1546,N_13738,N_13731);
xnor UO_1547 (O_1547,N_13679,N_14856);
and UO_1548 (O_1548,N_14917,N_13632);
or UO_1549 (O_1549,N_14963,N_14603);
and UO_1550 (O_1550,N_13634,N_14995);
and UO_1551 (O_1551,N_13959,N_14703);
xnor UO_1552 (O_1552,N_14000,N_14683);
or UO_1553 (O_1553,N_14284,N_13686);
xor UO_1554 (O_1554,N_13993,N_14452);
and UO_1555 (O_1555,N_13553,N_14312);
and UO_1556 (O_1556,N_13672,N_14175);
and UO_1557 (O_1557,N_14982,N_14098);
nor UO_1558 (O_1558,N_14510,N_14186);
xnor UO_1559 (O_1559,N_13843,N_14796);
or UO_1560 (O_1560,N_13987,N_14286);
or UO_1561 (O_1561,N_14563,N_13997);
nor UO_1562 (O_1562,N_14927,N_13859);
or UO_1563 (O_1563,N_14247,N_14774);
nor UO_1564 (O_1564,N_14040,N_13996);
nor UO_1565 (O_1565,N_13686,N_14227);
nand UO_1566 (O_1566,N_14974,N_13951);
nand UO_1567 (O_1567,N_14958,N_14135);
nand UO_1568 (O_1568,N_14461,N_13790);
and UO_1569 (O_1569,N_13571,N_14228);
xnor UO_1570 (O_1570,N_14942,N_13795);
or UO_1571 (O_1571,N_14156,N_14851);
nand UO_1572 (O_1572,N_14902,N_13811);
xor UO_1573 (O_1573,N_13613,N_13810);
xnor UO_1574 (O_1574,N_13589,N_14021);
nand UO_1575 (O_1575,N_14140,N_14294);
nor UO_1576 (O_1576,N_13535,N_14249);
nand UO_1577 (O_1577,N_14318,N_13559);
and UO_1578 (O_1578,N_14825,N_13703);
xor UO_1579 (O_1579,N_14209,N_13645);
nand UO_1580 (O_1580,N_13659,N_14222);
xnor UO_1581 (O_1581,N_13517,N_14170);
or UO_1582 (O_1582,N_13829,N_13740);
xor UO_1583 (O_1583,N_14510,N_14151);
xor UO_1584 (O_1584,N_13877,N_13928);
and UO_1585 (O_1585,N_13663,N_14870);
nor UO_1586 (O_1586,N_14112,N_13893);
or UO_1587 (O_1587,N_13751,N_13527);
or UO_1588 (O_1588,N_13772,N_13960);
or UO_1589 (O_1589,N_13908,N_14564);
nand UO_1590 (O_1590,N_14202,N_14950);
xor UO_1591 (O_1591,N_14576,N_14535);
nor UO_1592 (O_1592,N_14001,N_14557);
nor UO_1593 (O_1593,N_13959,N_14983);
xor UO_1594 (O_1594,N_13881,N_13743);
xor UO_1595 (O_1595,N_14828,N_14292);
and UO_1596 (O_1596,N_14592,N_14236);
and UO_1597 (O_1597,N_14994,N_14613);
xnor UO_1598 (O_1598,N_14581,N_14068);
xor UO_1599 (O_1599,N_14733,N_14017);
nor UO_1600 (O_1600,N_14621,N_14897);
nand UO_1601 (O_1601,N_14224,N_14990);
nor UO_1602 (O_1602,N_14095,N_14585);
xor UO_1603 (O_1603,N_13897,N_14464);
xnor UO_1604 (O_1604,N_14042,N_14328);
or UO_1605 (O_1605,N_14387,N_14751);
or UO_1606 (O_1606,N_13915,N_14116);
nand UO_1607 (O_1607,N_13685,N_14613);
xor UO_1608 (O_1608,N_13719,N_13999);
or UO_1609 (O_1609,N_14186,N_14948);
nor UO_1610 (O_1610,N_14448,N_14510);
or UO_1611 (O_1611,N_13598,N_14533);
or UO_1612 (O_1612,N_13930,N_14617);
or UO_1613 (O_1613,N_13982,N_14981);
or UO_1614 (O_1614,N_14784,N_13685);
nand UO_1615 (O_1615,N_14775,N_13886);
xnor UO_1616 (O_1616,N_14831,N_14614);
nand UO_1617 (O_1617,N_14732,N_13654);
nand UO_1618 (O_1618,N_13986,N_14672);
nor UO_1619 (O_1619,N_13709,N_13802);
xnor UO_1620 (O_1620,N_14163,N_13540);
nor UO_1621 (O_1621,N_14673,N_14033);
and UO_1622 (O_1622,N_14037,N_14947);
or UO_1623 (O_1623,N_13755,N_14791);
xor UO_1624 (O_1624,N_14374,N_13520);
or UO_1625 (O_1625,N_14711,N_14272);
or UO_1626 (O_1626,N_14118,N_13676);
and UO_1627 (O_1627,N_14230,N_14582);
nand UO_1628 (O_1628,N_14815,N_14791);
xor UO_1629 (O_1629,N_14131,N_14383);
nor UO_1630 (O_1630,N_14505,N_14401);
or UO_1631 (O_1631,N_14226,N_13882);
or UO_1632 (O_1632,N_14236,N_14983);
or UO_1633 (O_1633,N_14087,N_13739);
nand UO_1634 (O_1634,N_13820,N_14301);
nand UO_1635 (O_1635,N_14842,N_14691);
xnor UO_1636 (O_1636,N_14573,N_14702);
nand UO_1637 (O_1637,N_13594,N_14370);
and UO_1638 (O_1638,N_14611,N_14592);
and UO_1639 (O_1639,N_13829,N_13638);
xor UO_1640 (O_1640,N_13895,N_13506);
and UO_1641 (O_1641,N_13532,N_14859);
nand UO_1642 (O_1642,N_13794,N_14134);
or UO_1643 (O_1643,N_14720,N_13836);
nor UO_1644 (O_1644,N_14716,N_14196);
nor UO_1645 (O_1645,N_14781,N_14097);
xor UO_1646 (O_1646,N_14405,N_13823);
or UO_1647 (O_1647,N_13842,N_14925);
or UO_1648 (O_1648,N_13601,N_14753);
or UO_1649 (O_1649,N_14196,N_13973);
nor UO_1650 (O_1650,N_14885,N_14982);
and UO_1651 (O_1651,N_13952,N_14486);
xor UO_1652 (O_1652,N_14651,N_14856);
nor UO_1653 (O_1653,N_14783,N_14399);
or UO_1654 (O_1654,N_14373,N_14426);
nor UO_1655 (O_1655,N_14721,N_14920);
xnor UO_1656 (O_1656,N_14103,N_14763);
or UO_1657 (O_1657,N_14838,N_13838);
or UO_1658 (O_1658,N_13853,N_14453);
or UO_1659 (O_1659,N_13969,N_14678);
nand UO_1660 (O_1660,N_14582,N_14791);
nor UO_1661 (O_1661,N_14327,N_13925);
and UO_1662 (O_1662,N_14284,N_14655);
or UO_1663 (O_1663,N_14124,N_13898);
xor UO_1664 (O_1664,N_13558,N_14183);
or UO_1665 (O_1665,N_13795,N_14466);
nand UO_1666 (O_1666,N_13582,N_14176);
nand UO_1667 (O_1667,N_13975,N_13928);
xnor UO_1668 (O_1668,N_13974,N_14051);
nor UO_1669 (O_1669,N_14622,N_14684);
nor UO_1670 (O_1670,N_13762,N_13945);
nor UO_1671 (O_1671,N_13702,N_13597);
nand UO_1672 (O_1672,N_14413,N_13546);
nand UO_1673 (O_1673,N_13684,N_14237);
nor UO_1674 (O_1674,N_14470,N_13702);
xor UO_1675 (O_1675,N_14122,N_14181);
and UO_1676 (O_1676,N_14208,N_13780);
nor UO_1677 (O_1677,N_14198,N_14217);
xnor UO_1678 (O_1678,N_13921,N_14794);
and UO_1679 (O_1679,N_14292,N_14701);
and UO_1680 (O_1680,N_14687,N_14161);
or UO_1681 (O_1681,N_14907,N_13889);
or UO_1682 (O_1682,N_13670,N_14048);
and UO_1683 (O_1683,N_14356,N_14589);
xor UO_1684 (O_1684,N_14465,N_14518);
or UO_1685 (O_1685,N_13594,N_13951);
nand UO_1686 (O_1686,N_14264,N_14013);
nand UO_1687 (O_1687,N_14980,N_14905);
xor UO_1688 (O_1688,N_13973,N_13650);
nand UO_1689 (O_1689,N_13951,N_14166);
nand UO_1690 (O_1690,N_14948,N_13901);
xor UO_1691 (O_1691,N_14627,N_14089);
xor UO_1692 (O_1692,N_14694,N_14288);
xor UO_1693 (O_1693,N_13725,N_14259);
and UO_1694 (O_1694,N_13517,N_13717);
and UO_1695 (O_1695,N_13717,N_13666);
and UO_1696 (O_1696,N_14920,N_14694);
and UO_1697 (O_1697,N_14995,N_14231);
nand UO_1698 (O_1698,N_14058,N_13606);
or UO_1699 (O_1699,N_13760,N_13642);
and UO_1700 (O_1700,N_14231,N_14331);
nand UO_1701 (O_1701,N_14122,N_14580);
nor UO_1702 (O_1702,N_14911,N_13908);
or UO_1703 (O_1703,N_13998,N_13773);
nand UO_1704 (O_1704,N_14875,N_13503);
nand UO_1705 (O_1705,N_14955,N_13673);
nand UO_1706 (O_1706,N_13559,N_14368);
and UO_1707 (O_1707,N_14838,N_14459);
and UO_1708 (O_1708,N_13860,N_14064);
and UO_1709 (O_1709,N_13866,N_13544);
nand UO_1710 (O_1710,N_14110,N_13527);
or UO_1711 (O_1711,N_14026,N_14328);
or UO_1712 (O_1712,N_14161,N_14107);
xor UO_1713 (O_1713,N_14023,N_14989);
xor UO_1714 (O_1714,N_14408,N_13731);
or UO_1715 (O_1715,N_13834,N_14523);
nand UO_1716 (O_1716,N_13511,N_14681);
or UO_1717 (O_1717,N_13578,N_13853);
or UO_1718 (O_1718,N_14794,N_13504);
or UO_1719 (O_1719,N_13684,N_13738);
and UO_1720 (O_1720,N_14442,N_14834);
nand UO_1721 (O_1721,N_13542,N_14294);
xnor UO_1722 (O_1722,N_14401,N_14356);
or UO_1723 (O_1723,N_14564,N_13892);
and UO_1724 (O_1724,N_14297,N_14936);
and UO_1725 (O_1725,N_14373,N_13563);
xor UO_1726 (O_1726,N_14052,N_13545);
or UO_1727 (O_1727,N_14713,N_14577);
nand UO_1728 (O_1728,N_14189,N_14251);
or UO_1729 (O_1729,N_13988,N_14703);
and UO_1730 (O_1730,N_14194,N_13776);
and UO_1731 (O_1731,N_13897,N_14743);
and UO_1732 (O_1732,N_13802,N_13944);
and UO_1733 (O_1733,N_13704,N_14198);
and UO_1734 (O_1734,N_14770,N_14725);
and UO_1735 (O_1735,N_13910,N_13565);
xnor UO_1736 (O_1736,N_14937,N_14645);
nand UO_1737 (O_1737,N_13788,N_14544);
nand UO_1738 (O_1738,N_14867,N_14685);
nor UO_1739 (O_1739,N_14184,N_13856);
nand UO_1740 (O_1740,N_13751,N_14767);
xor UO_1741 (O_1741,N_14212,N_14161);
xnor UO_1742 (O_1742,N_14453,N_14771);
and UO_1743 (O_1743,N_14066,N_13646);
nor UO_1744 (O_1744,N_13576,N_14073);
and UO_1745 (O_1745,N_14936,N_14695);
nand UO_1746 (O_1746,N_14367,N_13684);
nor UO_1747 (O_1747,N_14659,N_14330);
nand UO_1748 (O_1748,N_13920,N_14834);
xnor UO_1749 (O_1749,N_14565,N_14672);
nand UO_1750 (O_1750,N_14390,N_14534);
nor UO_1751 (O_1751,N_14229,N_13653);
nand UO_1752 (O_1752,N_14217,N_13831);
nand UO_1753 (O_1753,N_13772,N_14604);
and UO_1754 (O_1754,N_14468,N_14107);
nor UO_1755 (O_1755,N_14237,N_14105);
nand UO_1756 (O_1756,N_14612,N_14150);
nand UO_1757 (O_1757,N_14505,N_14574);
nand UO_1758 (O_1758,N_14347,N_14878);
xor UO_1759 (O_1759,N_13892,N_14712);
or UO_1760 (O_1760,N_14868,N_14233);
nand UO_1761 (O_1761,N_13503,N_14176);
or UO_1762 (O_1762,N_14513,N_14977);
nor UO_1763 (O_1763,N_14335,N_13869);
or UO_1764 (O_1764,N_14261,N_14186);
nor UO_1765 (O_1765,N_14694,N_14240);
xor UO_1766 (O_1766,N_14316,N_13785);
nand UO_1767 (O_1767,N_14968,N_14280);
and UO_1768 (O_1768,N_14224,N_14049);
xnor UO_1769 (O_1769,N_13519,N_14130);
and UO_1770 (O_1770,N_14992,N_14672);
nor UO_1771 (O_1771,N_14189,N_14869);
or UO_1772 (O_1772,N_14510,N_13904);
nand UO_1773 (O_1773,N_14146,N_14690);
nor UO_1774 (O_1774,N_13959,N_14267);
or UO_1775 (O_1775,N_14433,N_13525);
nand UO_1776 (O_1776,N_13584,N_14227);
and UO_1777 (O_1777,N_14689,N_13657);
and UO_1778 (O_1778,N_13865,N_13878);
or UO_1779 (O_1779,N_14265,N_14320);
and UO_1780 (O_1780,N_14444,N_13717);
or UO_1781 (O_1781,N_14638,N_13802);
or UO_1782 (O_1782,N_13902,N_14841);
nor UO_1783 (O_1783,N_14687,N_13503);
nand UO_1784 (O_1784,N_14568,N_13888);
or UO_1785 (O_1785,N_13955,N_14174);
nand UO_1786 (O_1786,N_14356,N_14343);
and UO_1787 (O_1787,N_13656,N_14813);
nand UO_1788 (O_1788,N_14443,N_14533);
and UO_1789 (O_1789,N_14488,N_14130);
nor UO_1790 (O_1790,N_14622,N_13736);
xor UO_1791 (O_1791,N_14509,N_14930);
and UO_1792 (O_1792,N_14170,N_13913);
or UO_1793 (O_1793,N_13915,N_14752);
or UO_1794 (O_1794,N_14666,N_14338);
xor UO_1795 (O_1795,N_14494,N_13779);
nand UO_1796 (O_1796,N_14735,N_13532);
xor UO_1797 (O_1797,N_14628,N_14080);
nand UO_1798 (O_1798,N_14810,N_13605);
or UO_1799 (O_1799,N_14554,N_13826);
or UO_1800 (O_1800,N_14137,N_13500);
nand UO_1801 (O_1801,N_14584,N_14816);
or UO_1802 (O_1802,N_14075,N_14727);
and UO_1803 (O_1803,N_14817,N_13548);
xnor UO_1804 (O_1804,N_14566,N_14545);
and UO_1805 (O_1805,N_14980,N_13995);
nand UO_1806 (O_1806,N_13588,N_13667);
nand UO_1807 (O_1807,N_14439,N_14943);
xnor UO_1808 (O_1808,N_14542,N_14616);
nand UO_1809 (O_1809,N_14531,N_14032);
and UO_1810 (O_1810,N_14073,N_13796);
and UO_1811 (O_1811,N_14896,N_14829);
xnor UO_1812 (O_1812,N_14826,N_14395);
nor UO_1813 (O_1813,N_14890,N_13609);
nor UO_1814 (O_1814,N_14859,N_14086);
or UO_1815 (O_1815,N_14421,N_13940);
nand UO_1816 (O_1816,N_13677,N_14760);
or UO_1817 (O_1817,N_14392,N_14076);
xnor UO_1818 (O_1818,N_13515,N_14841);
nand UO_1819 (O_1819,N_13904,N_14580);
or UO_1820 (O_1820,N_14469,N_13884);
xor UO_1821 (O_1821,N_13594,N_14834);
and UO_1822 (O_1822,N_13734,N_13854);
nor UO_1823 (O_1823,N_14989,N_14004);
nand UO_1824 (O_1824,N_13636,N_13749);
and UO_1825 (O_1825,N_14645,N_14884);
nor UO_1826 (O_1826,N_14595,N_14647);
nand UO_1827 (O_1827,N_14157,N_14662);
nor UO_1828 (O_1828,N_14631,N_14620);
xor UO_1829 (O_1829,N_13658,N_14566);
nand UO_1830 (O_1830,N_14055,N_14623);
nand UO_1831 (O_1831,N_14974,N_14828);
and UO_1832 (O_1832,N_14157,N_13592);
xor UO_1833 (O_1833,N_14735,N_13938);
or UO_1834 (O_1834,N_14721,N_14876);
or UO_1835 (O_1835,N_13972,N_14454);
xor UO_1836 (O_1836,N_14741,N_14432);
nand UO_1837 (O_1837,N_14662,N_13559);
and UO_1838 (O_1838,N_14149,N_13546);
or UO_1839 (O_1839,N_14058,N_13875);
or UO_1840 (O_1840,N_14790,N_14540);
and UO_1841 (O_1841,N_14188,N_14064);
and UO_1842 (O_1842,N_14126,N_13736);
nor UO_1843 (O_1843,N_13817,N_13629);
xor UO_1844 (O_1844,N_13533,N_14778);
nand UO_1845 (O_1845,N_13810,N_14428);
xnor UO_1846 (O_1846,N_14684,N_14637);
and UO_1847 (O_1847,N_13866,N_14057);
or UO_1848 (O_1848,N_14381,N_13928);
or UO_1849 (O_1849,N_13928,N_13915);
xor UO_1850 (O_1850,N_14628,N_13573);
or UO_1851 (O_1851,N_13609,N_13560);
xnor UO_1852 (O_1852,N_14929,N_14972);
and UO_1853 (O_1853,N_13645,N_14188);
xnor UO_1854 (O_1854,N_13585,N_14232);
xor UO_1855 (O_1855,N_13600,N_14358);
nand UO_1856 (O_1856,N_13802,N_13727);
or UO_1857 (O_1857,N_14496,N_13644);
or UO_1858 (O_1858,N_14319,N_13720);
or UO_1859 (O_1859,N_14623,N_14484);
xnor UO_1860 (O_1860,N_13790,N_14721);
xnor UO_1861 (O_1861,N_14307,N_14094);
nor UO_1862 (O_1862,N_14219,N_13786);
xor UO_1863 (O_1863,N_14224,N_13512);
nand UO_1864 (O_1864,N_14998,N_14532);
xnor UO_1865 (O_1865,N_14434,N_14752);
and UO_1866 (O_1866,N_14008,N_14497);
nor UO_1867 (O_1867,N_14191,N_14578);
or UO_1868 (O_1868,N_14557,N_14260);
xnor UO_1869 (O_1869,N_14391,N_13667);
or UO_1870 (O_1870,N_14958,N_13569);
nand UO_1871 (O_1871,N_14554,N_14294);
xnor UO_1872 (O_1872,N_13716,N_14881);
nor UO_1873 (O_1873,N_13542,N_13813);
xnor UO_1874 (O_1874,N_14773,N_14487);
xor UO_1875 (O_1875,N_14729,N_14949);
and UO_1876 (O_1876,N_13506,N_14776);
or UO_1877 (O_1877,N_14354,N_13883);
or UO_1878 (O_1878,N_14670,N_13801);
nand UO_1879 (O_1879,N_13595,N_14689);
xor UO_1880 (O_1880,N_14287,N_14984);
or UO_1881 (O_1881,N_14718,N_14714);
and UO_1882 (O_1882,N_14667,N_13501);
xnor UO_1883 (O_1883,N_13632,N_14576);
nor UO_1884 (O_1884,N_13782,N_13797);
nand UO_1885 (O_1885,N_14988,N_14081);
nor UO_1886 (O_1886,N_14533,N_14053);
or UO_1887 (O_1887,N_13573,N_14721);
xor UO_1888 (O_1888,N_14236,N_13880);
nor UO_1889 (O_1889,N_13709,N_14351);
and UO_1890 (O_1890,N_14113,N_14896);
xor UO_1891 (O_1891,N_14511,N_14182);
and UO_1892 (O_1892,N_14483,N_13522);
nor UO_1893 (O_1893,N_13749,N_14904);
or UO_1894 (O_1894,N_14860,N_13941);
and UO_1895 (O_1895,N_13921,N_14869);
or UO_1896 (O_1896,N_14843,N_13705);
nand UO_1897 (O_1897,N_13870,N_13899);
or UO_1898 (O_1898,N_13798,N_14734);
xnor UO_1899 (O_1899,N_13582,N_14990);
nor UO_1900 (O_1900,N_13631,N_14494);
and UO_1901 (O_1901,N_14302,N_14396);
and UO_1902 (O_1902,N_13609,N_14811);
nor UO_1903 (O_1903,N_14344,N_13605);
or UO_1904 (O_1904,N_14911,N_14702);
or UO_1905 (O_1905,N_14166,N_13792);
nor UO_1906 (O_1906,N_13807,N_14969);
or UO_1907 (O_1907,N_14061,N_13573);
nand UO_1908 (O_1908,N_13789,N_14334);
and UO_1909 (O_1909,N_13763,N_14376);
and UO_1910 (O_1910,N_14376,N_13714);
xnor UO_1911 (O_1911,N_13974,N_14209);
nor UO_1912 (O_1912,N_14855,N_14982);
or UO_1913 (O_1913,N_13605,N_14955);
and UO_1914 (O_1914,N_14671,N_14264);
nor UO_1915 (O_1915,N_13980,N_14995);
and UO_1916 (O_1916,N_14514,N_14649);
xor UO_1917 (O_1917,N_14857,N_14919);
nand UO_1918 (O_1918,N_14532,N_13983);
xor UO_1919 (O_1919,N_14176,N_13664);
xor UO_1920 (O_1920,N_14592,N_14011);
nor UO_1921 (O_1921,N_14364,N_14508);
nor UO_1922 (O_1922,N_14228,N_14452);
nand UO_1923 (O_1923,N_13591,N_14365);
nor UO_1924 (O_1924,N_13524,N_13563);
and UO_1925 (O_1925,N_13569,N_14104);
and UO_1926 (O_1926,N_13896,N_14288);
and UO_1927 (O_1927,N_14361,N_13563);
nor UO_1928 (O_1928,N_13626,N_14545);
nor UO_1929 (O_1929,N_14457,N_13800);
or UO_1930 (O_1930,N_14526,N_14884);
nor UO_1931 (O_1931,N_14571,N_13885);
or UO_1932 (O_1932,N_14918,N_14077);
nand UO_1933 (O_1933,N_14061,N_14367);
xnor UO_1934 (O_1934,N_14778,N_14464);
nor UO_1935 (O_1935,N_13775,N_14307);
nand UO_1936 (O_1936,N_13747,N_14013);
nor UO_1937 (O_1937,N_14245,N_14237);
and UO_1938 (O_1938,N_13696,N_14460);
nor UO_1939 (O_1939,N_13699,N_14131);
xnor UO_1940 (O_1940,N_14913,N_14507);
or UO_1941 (O_1941,N_14704,N_13533);
nand UO_1942 (O_1942,N_13799,N_14634);
nor UO_1943 (O_1943,N_13964,N_13611);
nand UO_1944 (O_1944,N_14444,N_14373);
or UO_1945 (O_1945,N_14990,N_13966);
nand UO_1946 (O_1946,N_14214,N_14574);
and UO_1947 (O_1947,N_14198,N_13711);
and UO_1948 (O_1948,N_14971,N_14021);
xnor UO_1949 (O_1949,N_14514,N_14226);
nand UO_1950 (O_1950,N_14960,N_14124);
xnor UO_1951 (O_1951,N_13995,N_14377);
or UO_1952 (O_1952,N_13641,N_14507);
nor UO_1953 (O_1953,N_14877,N_14727);
nor UO_1954 (O_1954,N_14597,N_14460);
nor UO_1955 (O_1955,N_13572,N_14334);
or UO_1956 (O_1956,N_13880,N_14564);
and UO_1957 (O_1957,N_14147,N_14538);
and UO_1958 (O_1958,N_14829,N_14238);
nor UO_1959 (O_1959,N_14221,N_14657);
and UO_1960 (O_1960,N_14942,N_13518);
and UO_1961 (O_1961,N_14317,N_14052);
nor UO_1962 (O_1962,N_14232,N_14910);
xor UO_1963 (O_1963,N_14252,N_14033);
or UO_1964 (O_1964,N_14351,N_14700);
xnor UO_1965 (O_1965,N_13591,N_14681);
nand UO_1966 (O_1966,N_14208,N_13681);
and UO_1967 (O_1967,N_13910,N_14054);
xnor UO_1968 (O_1968,N_14084,N_14790);
or UO_1969 (O_1969,N_14429,N_14966);
or UO_1970 (O_1970,N_14566,N_14382);
or UO_1971 (O_1971,N_14405,N_14787);
xnor UO_1972 (O_1972,N_13967,N_14497);
nor UO_1973 (O_1973,N_13631,N_13933);
nand UO_1974 (O_1974,N_14222,N_13807);
nor UO_1975 (O_1975,N_14812,N_14616);
nand UO_1976 (O_1976,N_14943,N_14764);
nand UO_1977 (O_1977,N_14482,N_14624);
nand UO_1978 (O_1978,N_13830,N_14659);
xor UO_1979 (O_1979,N_14838,N_13721);
and UO_1980 (O_1980,N_14460,N_14252);
nand UO_1981 (O_1981,N_14110,N_14029);
or UO_1982 (O_1982,N_13788,N_14355);
nand UO_1983 (O_1983,N_14169,N_14297);
nand UO_1984 (O_1984,N_13859,N_14883);
or UO_1985 (O_1985,N_13726,N_14146);
or UO_1986 (O_1986,N_14441,N_14128);
xnor UO_1987 (O_1987,N_13505,N_14533);
or UO_1988 (O_1988,N_14783,N_13794);
or UO_1989 (O_1989,N_14080,N_14806);
and UO_1990 (O_1990,N_13655,N_14476);
nor UO_1991 (O_1991,N_14961,N_14550);
nor UO_1992 (O_1992,N_14391,N_14011);
and UO_1993 (O_1993,N_14429,N_14543);
and UO_1994 (O_1994,N_14872,N_14990);
nor UO_1995 (O_1995,N_14181,N_13859);
and UO_1996 (O_1996,N_14882,N_14760);
nor UO_1997 (O_1997,N_14908,N_14103);
xnor UO_1998 (O_1998,N_14791,N_14668);
nor UO_1999 (O_1999,N_14953,N_13546);
endmodule