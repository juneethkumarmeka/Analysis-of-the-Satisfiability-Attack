module basic_500_3000_500_4_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_488,In_105);
nor U1 (N_1,In_9,In_101);
or U2 (N_2,In_108,In_75);
or U3 (N_3,In_282,In_409);
nand U4 (N_4,In_181,In_286);
xnor U5 (N_5,In_98,In_112);
nand U6 (N_6,In_257,In_198);
and U7 (N_7,In_53,In_344);
nand U8 (N_8,In_363,In_396);
nor U9 (N_9,In_325,In_425);
nand U10 (N_10,In_432,In_273);
nor U11 (N_11,In_251,In_35);
or U12 (N_12,In_403,In_377);
or U13 (N_13,In_66,In_358);
and U14 (N_14,In_335,In_236);
or U15 (N_15,In_65,In_24);
nand U16 (N_16,In_380,In_364);
nor U17 (N_17,In_139,In_362);
or U18 (N_18,In_287,In_427);
nor U19 (N_19,In_39,In_88);
and U20 (N_20,In_72,In_448);
or U21 (N_21,In_111,In_367);
or U22 (N_22,In_136,In_152);
nand U23 (N_23,In_373,In_302);
nor U24 (N_24,In_34,In_308);
and U25 (N_25,In_319,In_383);
nand U26 (N_26,In_232,In_482);
and U27 (N_27,In_324,In_200);
xor U28 (N_28,In_390,In_94);
or U29 (N_29,In_384,In_244);
and U30 (N_30,In_155,In_180);
and U31 (N_31,In_276,In_428);
xor U32 (N_32,In_320,In_197);
or U33 (N_33,In_394,In_32);
or U34 (N_34,In_168,In_116);
nand U35 (N_35,In_30,In_387);
nand U36 (N_36,In_243,In_379);
and U37 (N_37,In_43,In_103);
xor U38 (N_38,In_256,In_222);
nand U39 (N_39,In_199,In_290);
or U40 (N_40,In_16,In_188);
nor U41 (N_41,In_331,In_63);
nor U42 (N_42,In_350,In_418);
or U43 (N_43,In_146,In_453);
nor U44 (N_44,In_374,In_494);
nand U45 (N_45,In_420,In_399);
nor U46 (N_46,In_104,In_144);
xnor U47 (N_47,In_359,In_346);
and U48 (N_48,In_372,In_398);
xor U49 (N_49,In_449,In_412);
xnor U50 (N_50,In_122,In_347);
xnor U51 (N_51,In_392,In_393);
nor U52 (N_52,In_457,In_334);
xor U53 (N_53,In_441,In_460);
or U54 (N_54,In_71,In_247);
or U55 (N_55,In_433,In_120);
and U56 (N_56,In_81,In_215);
xnor U57 (N_57,In_493,In_458);
or U58 (N_58,In_311,In_134);
and U59 (N_59,In_326,In_14);
or U60 (N_60,In_430,In_321);
and U61 (N_61,In_316,In_401);
or U62 (N_62,In_22,In_499);
or U63 (N_63,In_61,In_317);
and U64 (N_64,In_107,In_205);
or U65 (N_65,In_456,In_267);
nor U66 (N_66,In_312,In_291);
or U67 (N_67,In_391,In_218);
and U68 (N_68,In_2,In_224);
and U69 (N_69,In_130,In_261);
xnor U70 (N_70,In_309,In_85);
nand U71 (N_71,In_477,In_31);
and U72 (N_72,In_327,In_459);
xor U73 (N_73,In_231,In_495);
xor U74 (N_74,In_249,In_12);
and U75 (N_75,In_361,In_365);
and U76 (N_76,In_44,In_370);
nand U77 (N_77,In_260,In_138);
or U78 (N_78,In_410,In_92);
or U79 (N_79,In_20,In_162);
nand U80 (N_80,In_382,In_330);
or U81 (N_81,In_190,In_141);
nand U82 (N_82,In_27,In_51);
nor U83 (N_83,In_313,In_296);
nand U84 (N_84,In_113,In_167);
xnor U85 (N_85,In_164,In_354);
xnor U86 (N_86,In_288,In_69);
xor U87 (N_87,In_413,In_151);
and U88 (N_88,In_442,In_351);
xnor U89 (N_89,In_10,In_315);
or U90 (N_90,In_411,In_233);
nand U91 (N_91,In_169,In_343);
xor U92 (N_92,In_73,In_87);
nor U93 (N_93,In_258,In_234);
nor U94 (N_94,In_323,In_26);
xor U95 (N_95,In_227,In_270);
xnor U96 (N_96,In_48,In_481);
and U97 (N_97,In_280,In_297);
and U98 (N_98,In_110,In_452);
nand U99 (N_99,In_40,In_90);
xnor U100 (N_100,In_473,In_158);
nand U101 (N_101,In_443,In_17);
or U102 (N_102,In_194,In_255);
xnor U103 (N_103,In_230,In_49);
xor U104 (N_104,In_269,In_414);
or U105 (N_105,In_422,In_89);
nor U106 (N_106,In_467,In_471);
xnor U107 (N_107,In_118,In_23);
nor U108 (N_108,In_239,In_114);
nand U109 (N_109,In_496,In_100);
and U110 (N_110,In_42,In_153);
nor U111 (N_111,In_15,In_419);
or U112 (N_112,In_429,In_307);
nor U113 (N_113,In_339,In_212);
nor U114 (N_114,In_62,In_440);
or U115 (N_115,In_45,In_491);
nor U116 (N_116,In_83,In_191);
or U117 (N_117,In_463,In_192);
nand U118 (N_118,In_126,In_333);
xor U119 (N_119,In_208,In_479);
nor U120 (N_120,In_464,In_68);
nor U121 (N_121,In_274,In_163);
or U122 (N_122,In_283,In_226);
and U123 (N_123,In_140,In_210);
nand U124 (N_124,In_397,In_462);
or U125 (N_125,In_59,In_97);
nor U126 (N_126,In_264,In_439);
xor U127 (N_127,In_124,In_156);
nor U128 (N_128,In_400,In_252);
nand U129 (N_129,In_119,In_29);
nor U130 (N_130,In_366,In_298);
nor U131 (N_131,In_182,In_193);
nand U132 (N_132,In_360,In_117);
xnor U133 (N_133,In_240,In_489);
or U134 (N_134,In_203,In_421);
or U135 (N_135,In_50,In_294);
nand U136 (N_136,In_173,In_11);
nor U137 (N_137,In_478,In_121);
xnor U138 (N_138,In_480,In_357);
nor U139 (N_139,In_201,In_238);
nor U140 (N_140,In_468,In_160);
nand U141 (N_141,In_484,In_213);
xnor U142 (N_142,In_127,In_466);
nor U143 (N_143,In_214,In_241);
nand U144 (N_144,In_349,In_295);
xor U145 (N_145,In_5,In_474);
or U146 (N_146,In_143,In_259);
xnor U147 (N_147,In_148,In_6);
and U148 (N_148,In_470,In_303);
nor U149 (N_149,In_46,In_487);
or U150 (N_150,In_483,In_99);
or U151 (N_151,In_245,In_41);
or U152 (N_152,In_301,In_137);
xnor U153 (N_153,In_490,In_228);
xnor U154 (N_154,In_171,In_246);
or U155 (N_155,In_207,In_314);
or U156 (N_156,In_211,In_328);
and U157 (N_157,In_202,In_128);
xnor U158 (N_158,In_38,In_125);
nand U159 (N_159,In_216,In_60);
nand U160 (N_160,In_78,In_389);
xnor U161 (N_161,In_345,In_284);
or U162 (N_162,In_135,In_271);
nor U163 (N_163,In_96,In_436);
xnor U164 (N_164,In_278,In_242);
nor U165 (N_165,In_109,In_332);
nor U166 (N_166,In_166,In_381);
nand U167 (N_167,In_0,In_434);
nand U168 (N_168,In_447,In_454);
and U169 (N_169,In_170,In_80);
xnor U170 (N_170,In_322,In_444);
or U171 (N_171,In_266,In_165);
and U172 (N_172,In_341,In_476);
and U173 (N_173,In_93,In_424);
and U174 (N_174,In_318,In_378);
and U175 (N_175,In_475,In_348);
nand U176 (N_176,In_189,In_426);
xor U177 (N_177,In_55,In_187);
and U178 (N_178,In_250,In_337);
nand U179 (N_179,In_157,In_54);
or U180 (N_180,In_265,In_272);
and U181 (N_181,In_465,In_289);
nor U182 (N_182,In_179,In_195);
nor U183 (N_183,In_47,In_18);
nand U184 (N_184,In_147,In_498);
and U185 (N_185,In_371,In_281);
and U186 (N_186,In_340,In_115);
and U187 (N_187,In_219,In_76);
xnor U188 (N_188,In_175,In_395);
nand U189 (N_189,In_21,In_279);
or U190 (N_190,In_445,In_417);
nor U191 (N_191,In_497,In_235);
xor U192 (N_192,In_416,In_84);
or U193 (N_193,In_106,In_229);
nor U194 (N_194,In_408,In_74);
or U195 (N_195,In_102,In_329);
and U196 (N_196,In_196,In_406);
nand U197 (N_197,In_293,In_91);
nand U198 (N_198,In_338,In_28);
xnor U199 (N_199,In_145,In_300);
nand U200 (N_200,In_19,In_217);
or U201 (N_201,In_369,In_52);
and U202 (N_202,In_25,In_355);
and U203 (N_203,In_172,In_402);
xnor U204 (N_204,In_178,In_469);
nand U205 (N_205,In_388,In_451);
nor U206 (N_206,In_64,In_186);
nand U207 (N_207,In_33,In_237);
nand U208 (N_208,In_386,In_123);
nand U209 (N_209,In_310,In_56);
xnor U210 (N_210,In_268,In_133);
or U211 (N_211,In_176,In_306);
and U212 (N_212,In_285,In_7);
nand U213 (N_213,In_305,In_86);
and U214 (N_214,In_431,In_485);
nor U215 (N_215,In_13,In_446);
xnor U216 (N_216,In_154,In_37);
nor U217 (N_217,In_1,In_159);
nor U218 (N_218,In_336,In_375);
nor U219 (N_219,In_437,In_263);
nand U220 (N_220,In_415,In_4);
nor U221 (N_221,In_184,In_342);
nor U222 (N_222,In_435,In_299);
nor U223 (N_223,In_58,In_220);
xor U224 (N_224,In_275,In_353);
or U225 (N_225,In_423,In_262);
or U226 (N_226,In_221,In_450);
nand U227 (N_227,In_209,In_149);
and U228 (N_228,In_407,In_82);
nand U229 (N_229,In_95,In_461);
nor U230 (N_230,In_248,In_150);
and U231 (N_231,In_472,In_292);
nor U232 (N_232,In_492,In_36);
nand U233 (N_233,In_254,In_277);
or U234 (N_234,In_3,In_376);
xnor U235 (N_235,In_352,In_304);
nand U236 (N_236,In_131,In_455);
or U237 (N_237,In_253,In_129);
xor U238 (N_238,In_57,In_385);
xnor U239 (N_239,In_486,In_404);
nand U240 (N_240,In_204,In_368);
nand U241 (N_241,In_132,In_438);
xor U242 (N_242,In_183,In_225);
or U243 (N_243,In_67,In_79);
xor U244 (N_244,In_206,In_185);
or U245 (N_245,In_142,In_77);
and U246 (N_246,In_174,In_223);
or U247 (N_247,In_161,In_405);
xnor U248 (N_248,In_356,In_70);
or U249 (N_249,In_177,In_8);
xnor U250 (N_250,In_27,In_301);
and U251 (N_251,In_441,In_172);
nor U252 (N_252,In_480,In_383);
or U253 (N_253,In_347,In_118);
nor U254 (N_254,In_62,In_327);
nand U255 (N_255,In_222,In_102);
or U256 (N_256,In_444,In_468);
and U257 (N_257,In_227,In_210);
nand U258 (N_258,In_338,In_130);
or U259 (N_259,In_450,In_466);
and U260 (N_260,In_358,In_159);
nand U261 (N_261,In_307,In_11);
and U262 (N_262,In_478,In_309);
and U263 (N_263,In_251,In_458);
nand U264 (N_264,In_4,In_83);
or U265 (N_265,In_370,In_433);
and U266 (N_266,In_166,In_404);
and U267 (N_267,In_237,In_386);
and U268 (N_268,In_347,In_2);
and U269 (N_269,In_280,In_14);
and U270 (N_270,In_207,In_277);
nor U271 (N_271,In_282,In_38);
or U272 (N_272,In_475,In_322);
xnor U273 (N_273,In_466,In_118);
or U274 (N_274,In_136,In_347);
or U275 (N_275,In_392,In_348);
nor U276 (N_276,In_435,In_43);
nand U277 (N_277,In_94,In_445);
and U278 (N_278,In_50,In_425);
xor U279 (N_279,In_144,In_11);
and U280 (N_280,In_467,In_165);
nor U281 (N_281,In_482,In_98);
xnor U282 (N_282,In_15,In_90);
xnor U283 (N_283,In_243,In_369);
nand U284 (N_284,In_404,In_461);
and U285 (N_285,In_330,In_157);
nor U286 (N_286,In_141,In_278);
or U287 (N_287,In_208,In_339);
nor U288 (N_288,In_426,In_440);
nand U289 (N_289,In_10,In_208);
and U290 (N_290,In_70,In_11);
and U291 (N_291,In_201,In_51);
or U292 (N_292,In_72,In_79);
or U293 (N_293,In_444,In_75);
nor U294 (N_294,In_397,In_290);
nor U295 (N_295,In_337,In_490);
and U296 (N_296,In_221,In_157);
nor U297 (N_297,In_195,In_347);
nand U298 (N_298,In_120,In_101);
nor U299 (N_299,In_126,In_169);
or U300 (N_300,In_410,In_196);
nor U301 (N_301,In_475,In_228);
nor U302 (N_302,In_358,In_188);
nand U303 (N_303,In_435,In_296);
nor U304 (N_304,In_452,In_400);
and U305 (N_305,In_37,In_104);
xor U306 (N_306,In_91,In_121);
nand U307 (N_307,In_162,In_7);
or U308 (N_308,In_7,In_39);
or U309 (N_309,In_439,In_177);
and U310 (N_310,In_123,In_418);
nor U311 (N_311,In_469,In_385);
or U312 (N_312,In_9,In_63);
and U313 (N_313,In_76,In_366);
and U314 (N_314,In_65,In_354);
xor U315 (N_315,In_314,In_324);
nor U316 (N_316,In_93,In_77);
or U317 (N_317,In_316,In_306);
nor U318 (N_318,In_170,In_421);
nand U319 (N_319,In_238,In_25);
xnor U320 (N_320,In_2,In_106);
xor U321 (N_321,In_308,In_149);
or U322 (N_322,In_326,In_126);
xor U323 (N_323,In_192,In_86);
xor U324 (N_324,In_182,In_171);
or U325 (N_325,In_298,In_181);
nand U326 (N_326,In_150,In_437);
and U327 (N_327,In_52,In_407);
nand U328 (N_328,In_208,In_151);
nor U329 (N_329,In_416,In_417);
and U330 (N_330,In_170,In_333);
nor U331 (N_331,In_77,In_410);
or U332 (N_332,In_283,In_471);
or U333 (N_333,In_222,In_479);
nand U334 (N_334,In_67,In_139);
nand U335 (N_335,In_277,In_184);
or U336 (N_336,In_124,In_231);
nor U337 (N_337,In_467,In_144);
nand U338 (N_338,In_410,In_120);
xnor U339 (N_339,In_115,In_469);
nor U340 (N_340,In_133,In_116);
nand U341 (N_341,In_97,In_389);
xnor U342 (N_342,In_137,In_241);
nor U343 (N_343,In_439,In_495);
nor U344 (N_344,In_437,In_471);
nor U345 (N_345,In_66,In_4);
and U346 (N_346,In_408,In_453);
xnor U347 (N_347,In_469,In_18);
nand U348 (N_348,In_347,In_134);
and U349 (N_349,In_222,In_489);
or U350 (N_350,In_354,In_30);
and U351 (N_351,In_95,In_363);
nand U352 (N_352,In_489,In_343);
and U353 (N_353,In_460,In_358);
or U354 (N_354,In_213,In_199);
and U355 (N_355,In_122,In_305);
nor U356 (N_356,In_143,In_91);
nand U357 (N_357,In_190,In_20);
and U358 (N_358,In_184,In_477);
xor U359 (N_359,In_497,In_228);
xnor U360 (N_360,In_271,In_116);
nand U361 (N_361,In_331,In_336);
nand U362 (N_362,In_444,In_166);
nand U363 (N_363,In_173,In_378);
and U364 (N_364,In_2,In_237);
or U365 (N_365,In_364,In_387);
nor U366 (N_366,In_2,In_391);
and U367 (N_367,In_344,In_121);
xnor U368 (N_368,In_339,In_241);
nor U369 (N_369,In_422,In_3);
xnor U370 (N_370,In_102,In_364);
nand U371 (N_371,In_243,In_120);
nand U372 (N_372,In_477,In_66);
nor U373 (N_373,In_260,In_112);
nor U374 (N_374,In_56,In_398);
and U375 (N_375,In_307,In_289);
nor U376 (N_376,In_435,In_159);
or U377 (N_377,In_199,In_391);
or U378 (N_378,In_10,In_470);
nand U379 (N_379,In_312,In_409);
xor U380 (N_380,In_140,In_264);
xor U381 (N_381,In_312,In_215);
nand U382 (N_382,In_13,In_358);
nand U383 (N_383,In_410,In_488);
nor U384 (N_384,In_413,In_259);
nor U385 (N_385,In_411,In_303);
nand U386 (N_386,In_443,In_465);
nor U387 (N_387,In_407,In_349);
and U388 (N_388,In_435,In_379);
xnor U389 (N_389,In_493,In_150);
nor U390 (N_390,In_148,In_135);
or U391 (N_391,In_210,In_131);
xnor U392 (N_392,In_145,In_285);
xor U393 (N_393,In_177,In_446);
xnor U394 (N_394,In_485,In_89);
nor U395 (N_395,In_183,In_281);
nor U396 (N_396,In_491,In_420);
xor U397 (N_397,In_274,In_32);
xor U398 (N_398,In_329,In_330);
or U399 (N_399,In_393,In_290);
nor U400 (N_400,In_19,In_82);
xor U401 (N_401,In_61,In_59);
nor U402 (N_402,In_415,In_201);
xor U403 (N_403,In_293,In_27);
and U404 (N_404,In_471,In_380);
nand U405 (N_405,In_436,In_419);
and U406 (N_406,In_116,In_288);
nand U407 (N_407,In_8,In_45);
and U408 (N_408,In_308,In_310);
and U409 (N_409,In_447,In_245);
or U410 (N_410,In_8,In_486);
xor U411 (N_411,In_332,In_144);
nor U412 (N_412,In_116,In_314);
nand U413 (N_413,In_301,In_341);
xor U414 (N_414,In_414,In_50);
xor U415 (N_415,In_337,In_128);
nand U416 (N_416,In_183,In_300);
xnor U417 (N_417,In_430,In_66);
or U418 (N_418,In_351,In_493);
or U419 (N_419,In_220,In_216);
or U420 (N_420,In_318,In_137);
and U421 (N_421,In_365,In_374);
or U422 (N_422,In_454,In_194);
or U423 (N_423,In_251,In_125);
and U424 (N_424,In_367,In_44);
or U425 (N_425,In_218,In_396);
or U426 (N_426,In_306,In_385);
nor U427 (N_427,In_491,In_300);
xnor U428 (N_428,In_407,In_15);
or U429 (N_429,In_370,In_88);
nor U430 (N_430,In_175,In_223);
xor U431 (N_431,In_242,In_167);
nand U432 (N_432,In_51,In_470);
nand U433 (N_433,In_189,In_177);
xor U434 (N_434,In_372,In_4);
and U435 (N_435,In_208,In_73);
nor U436 (N_436,In_315,In_443);
or U437 (N_437,In_375,In_79);
or U438 (N_438,In_282,In_442);
and U439 (N_439,In_380,In_188);
nor U440 (N_440,In_118,In_159);
nand U441 (N_441,In_20,In_397);
and U442 (N_442,In_186,In_275);
nor U443 (N_443,In_455,In_237);
and U444 (N_444,In_380,In_397);
or U445 (N_445,In_305,In_209);
xnor U446 (N_446,In_80,In_180);
nor U447 (N_447,In_496,In_194);
and U448 (N_448,In_90,In_53);
or U449 (N_449,In_215,In_117);
and U450 (N_450,In_277,In_490);
xnor U451 (N_451,In_35,In_21);
xor U452 (N_452,In_255,In_167);
and U453 (N_453,In_422,In_14);
nand U454 (N_454,In_341,In_52);
nand U455 (N_455,In_7,In_29);
nand U456 (N_456,In_329,In_192);
or U457 (N_457,In_254,In_262);
or U458 (N_458,In_494,In_212);
or U459 (N_459,In_170,In_427);
nor U460 (N_460,In_476,In_206);
nand U461 (N_461,In_386,In_286);
xor U462 (N_462,In_250,In_242);
or U463 (N_463,In_449,In_19);
xnor U464 (N_464,In_350,In_274);
and U465 (N_465,In_169,In_395);
or U466 (N_466,In_177,In_64);
xor U467 (N_467,In_444,In_170);
or U468 (N_468,In_24,In_497);
or U469 (N_469,In_364,In_133);
nand U470 (N_470,In_340,In_403);
or U471 (N_471,In_323,In_183);
nor U472 (N_472,In_365,In_140);
or U473 (N_473,In_123,In_364);
nand U474 (N_474,In_13,In_304);
or U475 (N_475,In_83,In_144);
and U476 (N_476,In_339,In_49);
xnor U477 (N_477,In_458,In_322);
xor U478 (N_478,In_304,In_465);
or U479 (N_479,In_215,In_342);
and U480 (N_480,In_305,In_107);
or U481 (N_481,In_65,In_342);
nand U482 (N_482,In_324,In_105);
nand U483 (N_483,In_34,In_107);
nor U484 (N_484,In_193,In_289);
xnor U485 (N_485,In_388,In_474);
nor U486 (N_486,In_469,In_380);
xor U487 (N_487,In_315,In_440);
and U488 (N_488,In_162,In_22);
or U489 (N_489,In_460,In_171);
xor U490 (N_490,In_106,In_89);
and U491 (N_491,In_261,In_450);
nor U492 (N_492,In_131,In_346);
or U493 (N_493,In_34,In_100);
and U494 (N_494,In_305,In_363);
xor U495 (N_495,In_303,In_203);
nor U496 (N_496,In_52,In_402);
and U497 (N_497,In_388,In_458);
or U498 (N_498,In_488,In_450);
and U499 (N_499,In_285,In_476);
xor U500 (N_500,In_147,In_314);
nand U501 (N_501,In_148,In_157);
or U502 (N_502,In_450,In_265);
nand U503 (N_503,In_452,In_335);
xor U504 (N_504,In_73,In_82);
nor U505 (N_505,In_92,In_204);
or U506 (N_506,In_55,In_485);
or U507 (N_507,In_410,In_306);
or U508 (N_508,In_390,In_442);
nor U509 (N_509,In_390,In_166);
xor U510 (N_510,In_457,In_33);
xnor U511 (N_511,In_127,In_176);
xor U512 (N_512,In_400,In_381);
nand U513 (N_513,In_123,In_266);
xor U514 (N_514,In_12,In_141);
xnor U515 (N_515,In_426,In_187);
nor U516 (N_516,In_422,In_28);
xor U517 (N_517,In_320,In_308);
or U518 (N_518,In_59,In_485);
or U519 (N_519,In_151,In_224);
or U520 (N_520,In_16,In_480);
xor U521 (N_521,In_299,In_420);
xor U522 (N_522,In_240,In_229);
and U523 (N_523,In_69,In_86);
nor U524 (N_524,In_39,In_52);
nand U525 (N_525,In_219,In_480);
nand U526 (N_526,In_154,In_70);
or U527 (N_527,In_255,In_254);
or U528 (N_528,In_42,In_82);
xnor U529 (N_529,In_74,In_325);
or U530 (N_530,In_382,In_198);
or U531 (N_531,In_446,In_421);
nor U532 (N_532,In_77,In_268);
nand U533 (N_533,In_247,In_278);
nand U534 (N_534,In_397,In_475);
nand U535 (N_535,In_422,In_431);
nand U536 (N_536,In_221,In_81);
nand U537 (N_537,In_141,In_210);
and U538 (N_538,In_443,In_279);
nor U539 (N_539,In_65,In_222);
nand U540 (N_540,In_30,In_5);
nor U541 (N_541,In_345,In_455);
or U542 (N_542,In_406,In_271);
nor U543 (N_543,In_329,In_195);
nor U544 (N_544,In_346,In_371);
and U545 (N_545,In_95,In_107);
nand U546 (N_546,In_40,In_246);
or U547 (N_547,In_80,In_298);
or U548 (N_548,In_398,In_442);
nor U549 (N_549,In_23,In_41);
xnor U550 (N_550,In_120,In_489);
nand U551 (N_551,In_317,In_92);
nand U552 (N_552,In_341,In_298);
xor U553 (N_553,In_388,In_375);
nor U554 (N_554,In_152,In_455);
nor U555 (N_555,In_246,In_9);
nand U556 (N_556,In_346,In_115);
nand U557 (N_557,In_144,In_425);
nor U558 (N_558,In_123,In_46);
nand U559 (N_559,In_38,In_414);
and U560 (N_560,In_151,In_227);
and U561 (N_561,In_414,In_219);
or U562 (N_562,In_478,In_496);
and U563 (N_563,In_42,In_426);
xnor U564 (N_564,In_301,In_232);
xnor U565 (N_565,In_417,In_3);
xor U566 (N_566,In_92,In_36);
or U567 (N_567,In_421,In_134);
nand U568 (N_568,In_264,In_336);
nand U569 (N_569,In_355,In_464);
and U570 (N_570,In_411,In_56);
or U571 (N_571,In_202,In_302);
nor U572 (N_572,In_213,In_165);
xnor U573 (N_573,In_373,In_18);
nand U574 (N_574,In_424,In_470);
and U575 (N_575,In_379,In_28);
nor U576 (N_576,In_99,In_485);
nand U577 (N_577,In_361,In_484);
nand U578 (N_578,In_468,In_261);
nor U579 (N_579,In_469,In_330);
xor U580 (N_580,In_33,In_135);
or U581 (N_581,In_136,In_403);
or U582 (N_582,In_89,In_200);
and U583 (N_583,In_62,In_102);
and U584 (N_584,In_231,In_25);
and U585 (N_585,In_345,In_51);
nor U586 (N_586,In_447,In_119);
xnor U587 (N_587,In_401,In_398);
or U588 (N_588,In_141,In_204);
or U589 (N_589,In_396,In_183);
nor U590 (N_590,In_200,In_20);
or U591 (N_591,In_119,In_474);
and U592 (N_592,In_282,In_90);
nand U593 (N_593,In_401,In_149);
nand U594 (N_594,In_86,In_107);
nand U595 (N_595,In_455,In_65);
or U596 (N_596,In_184,In_254);
and U597 (N_597,In_235,In_456);
xnor U598 (N_598,In_159,In_137);
nor U599 (N_599,In_354,In_297);
or U600 (N_600,In_345,In_246);
and U601 (N_601,In_60,In_245);
or U602 (N_602,In_322,In_163);
nor U603 (N_603,In_488,In_407);
xnor U604 (N_604,In_449,In_363);
and U605 (N_605,In_314,In_220);
nor U606 (N_606,In_206,In_463);
or U607 (N_607,In_132,In_36);
or U608 (N_608,In_248,In_424);
and U609 (N_609,In_279,In_405);
or U610 (N_610,In_351,In_108);
or U611 (N_611,In_313,In_486);
nand U612 (N_612,In_407,In_90);
nand U613 (N_613,In_24,In_233);
xor U614 (N_614,In_10,In_441);
xor U615 (N_615,In_442,In_267);
and U616 (N_616,In_6,In_91);
or U617 (N_617,In_318,In_99);
nor U618 (N_618,In_383,In_20);
xnor U619 (N_619,In_380,In_214);
xor U620 (N_620,In_318,In_478);
nor U621 (N_621,In_260,In_235);
xnor U622 (N_622,In_389,In_178);
and U623 (N_623,In_178,In_381);
nor U624 (N_624,In_17,In_162);
and U625 (N_625,In_58,In_12);
and U626 (N_626,In_140,In_152);
nand U627 (N_627,In_261,In_197);
nor U628 (N_628,In_5,In_430);
nor U629 (N_629,In_382,In_43);
nand U630 (N_630,In_20,In_336);
xor U631 (N_631,In_60,In_2);
or U632 (N_632,In_130,In_438);
xnor U633 (N_633,In_481,In_234);
or U634 (N_634,In_127,In_413);
and U635 (N_635,In_279,In_43);
or U636 (N_636,In_55,In_435);
and U637 (N_637,In_111,In_473);
and U638 (N_638,In_459,In_265);
nand U639 (N_639,In_97,In_236);
nand U640 (N_640,In_302,In_307);
nor U641 (N_641,In_251,In_16);
or U642 (N_642,In_395,In_42);
or U643 (N_643,In_403,In_184);
and U644 (N_644,In_487,In_205);
or U645 (N_645,In_90,In_334);
or U646 (N_646,In_488,In_177);
nand U647 (N_647,In_151,In_306);
nand U648 (N_648,In_91,In_303);
and U649 (N_649,In_449,In_299);
nand U650 (N_650,In_14,In_21);
and U651 (N_651,In_331,In_108);
xnor U652 (N_652,In_472,In_236);
nor U653 (N_653,In_81,In_350);
or U654 (N_654,In_499,In_25);
nor U655 (N_655,In_331,In_160);
or U656 (N_656,In_268,In_390);
nand U657 (N_657,In_405,In_344);
nand U658 (N_658,In_329,In_427);
nor U659 (N_659,In_492,In_391);
nor U660 (N_660,In_271,In_106);
nor U661 (N_661,In_338,In_107);
xnor U662 (N_662,In_373,In_71);
or U663 (N_663,In_299,In_296);
xnor U664 (N_664,In_199,In_339);
and U665 (N_665,In_185,In_36);
xnor U666 (N_666,In_278,In_269);
or U667 (N_667,In_301,In_20);
or U668 (N_668,In_492,In_62);
or U669 (N_669,In_52,In_82);
or U670 (N_670,In_22,In_471);
nand U671 (N_671,In_489,In_200);
nand U672 (N_672,In_298,In_31);
or U673 (N_673,In_263,In_139);
xnor U674 (N_674,In_486,In_153);
nand U675 (N_675,In_462,In_224);
or U676 (N_676,In_175,In_97);
and U677 (N_677,In_414,In_280);
and U678 (N_678,In_58,In_336);
nor U679 (N_679,In_444,In_381);
or U680 (N_680,In_238,In_72);
nor U681 (N_681,In_4,In_84);
nor U682 (N_682,In_201,In_95);
nor U683 (N_683,In_102,In_488);
and U684 (N_684,In_75,In_236);
or U685 (N_685,In_410,In_143);
nand U686 (N_686,In_414,In_0);
or U687 (N_687,In_109,In_491);
xnor U688 (N_688,In_52,In_126);
and U689 (N_689,In_473,In_291);
nor U690 (N_690,In_12,In_69);
or U691 (N_691,In_449,In_326);
nor U692 (N_692,In_366,In_36);
nor U693 (N_693,In_231,In_367);
nor U694 (N_694,In_129,In_64);
nand U695 (N_695,In_407,In_350);
nor U696 (N_696,In_399,In_191);
nand U697 (N_697,In_102,In_400);
nor U698 (N_698,In_409,In_34);
xnor U699 (N_699,In_426,In_481);
and U700 (N_700,In_62,In_7);
xnor U701 (N_701,In_260,In_277);
nand U702 (N_702,In_455,In_445);
xor U703 (N_703,In_392,In_207);
or U704 (N_704,In_204,In_410);
nor U705 (N_705,In_134,In_310);
xnor U706 (N_706,In_121,In_295);
nor U707 (N_707,In_221,In_251);
nor U708 (N_708,In_441,In_304);
nor U709 (N_709,In_307,In_248);
nand U710 (N_710,In_139,In_191);
xnor U711 (N_711,In_202,In_458);
and U712 (N_712,In_403,In_392);
nand U713 (N_713,In_96,In_45);
or U714 (N_714,In_494,In_129);
or U715 (N_715,In_185,In_144);
xnor U716 (N_716,In_448,In_495);
nor U717 (N_717,In_475,In_380);
nor U718 (N_718,In_284,In_185);
nor U719 (N_719,In_490,In_442);
or U720 (N_720,In_256,In_326);
nand U721 (N_721,In_327,In_147);
nand U722 (N_722,In_233,In_464);
nand U723 (N_723,In_325,In_207);
xnor U724 (N_724,In_82,In_430);
and U725 (N_725,In_379,In_311);
nor U726 (N_726,In_25,In_78);
and U727 (N_727,In_399,In_169);
nor U728 (N_728,In_406,In_318);
and U729 (N_729,In_236,In_321);
and U730 (N_730,In_419,In_288);
or U731 (N_731,In_241,In_429);
xor U732 (N_732,In_386,In_296);
nand U733 (N_733,In_297,In_39);
and U734 (N_734,In_88,In_60);
or U735 (N_735,In_205,In_349);
nor U736 (N_736,In_483,In_463);
and U737 (N_737,In_376,In_104);
xnor U738 (N_738,In_470,In_269);
and U739 (N_739,In_312,In_98);
xor U740 (N_740,In_227,In_14);
or U741 (N_741,In_202,In_416);
xnor U742 (N_742,In_297,In_138);
xor U743 (N_743,In_343,In_267);
nor U744 (N_744,In_438,In_452);
or U745 (N_745,In_257,In_231);
nor U746 (N_746,In_474,In_142);
nor U747 (N_747,In_20,In_207);
xnor U748 (N_748,In_9,In_451);
and U749 (N_749,In_178,In_407);
nand U750 (N_750,N_362,N_732);
nor U751 (N_751,N_639,N_156);
nor U752 (N_752,N_204,N_637);
nor U753 (N_753,N_647,N_16);
or U754 (N_754,N_66,N_277);
and U755 (N_755,N_583,N_106);
nor U756 (N_756,N_36,N_683);
xnor U757 (N_757,N_88,N_128);
xnor U758 (N_758,N_234,N_314);
xnor U759 (N_759,N_311,N_219);
xnor U760 (N_760,N_181,N_169);
nor U761 (N_761,N_472,N_555);
or U762 (N_762,N_64,N_720);
xor U763 (N_763,N_225,N_25);
or U764 (N_764,N_684,N_587);
nor U765 (N_765,N_40,N_523);
and U766 (N_766,N_86,N_265);
xnor U767 (N_767,N_586,N_350);
xnor U768 (N_768,N_680,N_561);
nor U769 (N_769,N_655,N_742);
and U770 (N_770,N_13,N_443);
xor U771 (N_771,N_255,N_266);
xnor U772 (N_772,N_308,N_30);
and U773 (N_773,N_323,N_295);
nand U774 (N_774,N_540,N_629);
nand U775 (N_775,N_528,N_662);
xnor U776 (N_776,N_221,N_107);
xor U777 (N_777,N_290,N_663);
nor U778 (N_778,N_320,N_457);
xor U779 (N_779,N_356,N_313);
nor U780 (N_780,N_82,N_746);
xor U781 (N_781,N_393,N_409);
xor U782 (N_782,N_612,N_432);
nand U783 (N_783,N_8,N_212);
or U784 (N_784,N_116,N_450);
or U785 (N_785,N_653,N_304);
xor U786 (N_786,N_672,N_344);
and U787 (N_787,N_147,N_203);
or U788 (N_788,N_208,N_584);
or U789 (N_789,N_187,N_456);
or U790 (N_790,N_389,N_363);
nand U791 (N_791,N_482,N_231);
nor U792 (N_792,N_97,N_724);
xnor U793 (N_793,N_309,N_26);
or U794 (N_794,N_137,N_278);
xor U795 (N_795,N_486,N_174);
or U796 (N_796,N_142,N_595);
xnor U797 (N_797,N_455,N_74);
and U798 (N_798,N_711,N_339);
nor U799 (N_799,N_469,N_287);
and U800 (N_800,N_183,N_39);
xor U801 (N_801,N_448,N_84);
nand U802 (N_802,N_246,N_638);
and U803 (N_803,N_570,N_236);
and U804 (N_804,N_240,N_360);
or U805 (N_805,N_155,N_85);
xor U806 (N_806,N_307,N_370);
nor U807 (N_807,N_330,N_485);
xnor U808 (N_808,N_607,N_238);
nor U809 (N_809,N_585,N_623);
xnor U810 (N_810,N_121,N_705);
nand U811 (N_811,N_703,N_37);
or U812 (N_812,N_110,N_618);
nor U813 (N_813,N_163,N_524);
xnor U814 (N_814,N_94,N_251);
and U815 (N_815,N_60,N_691);
nand U816 (N_816,N_220,N_275);
nand U817 (N_817,N_127,N_197);
or U818 (N_818,N_264,N_748);
nor U819 (N_819,N_382,N_145);
or U820 (N_820,N_466,N_699);
nor U821 (N_821,N_20,N_256);
nor U822 (N_822,N_267,N_398);
or U823 (N_823,N_616,N_345);
and U824 (N_824,N_546,N_374);
or U825 (N_825,N_130,N_42);
nor U826 (N_826,N_46,N_723);
and U827 (N_827,N_564,N_715);
or U828 (N_828,N_736,N_118);
or U829 (N_829,N_5,N_424);
nand U830 (N_830,N_475,N_654);
and U831 (N_831,N_114,N_452);
nor U832 (N_832,N_373,N_708);
nor U833 (N_833,N_138,N_376);
or U834 (N_834,N_451,N_721);
nor U835 (N_835,N_168,N_605);
or U836 (N_836,N_553,N_505);
nand U837 (N_837,N_429,N_415);
nor U838 (N_838,N_681,N_159);
xor U839 (N_839,N_157,N_425);
nor U840 (N_840,N_481,N_29);
nand U841 (N_841,N_588,N_222);
nand U842 (N_842,N_24,N_704);
and U843 (N_843,N_65,N_151);
or U844 (N_844,N_508,N_354);
or U845 (N_845,N_454,N_213);
xnor U846 (N_846,N_148,N_227);
nand U847 (N_847,N_651,N_743);
nor U848 (N_848,N_559,N_375);
nand U849 (N_849,N_658,N_202);
or U850 (N_850,N_75,N_2);
and U851 (N_851,N_657,N_58);
nand U852 (N_852,N_368,N_115);
nor U853 (N_853,N_606,N_310);
xor U854 (N_854,N_334,N_596);
or U855 (N_855,N_648,N_284);
or U856 (N_856,N_512,N_92);
and U857 (N_857,N_641,N_158);
and U858 (N_858,N_93,N_661);
or U859 (N_859,N_534,N_297);
nand U860 (N_860,N_462,N_133);
xor U861 (N_861,N_513,N_150);
or U862 (N_862,N_269,N_132);
xor U863 (N_863,N_601,N_511);
nand U864 (N_864,N_614,N_427);
nand U865 (N_865,N_192,N_49);
or U866 (N_866,N_631,N_119);
nor U867 (N_867,N_140,N_332);
and U868 (N_868,N_272,N_161);
and U869 (N_869,N_281,N_500);
and U870 (N_870,N_81,N_733);
xnor U871 (N_871,N_687,N_293);
and U872 (N_872,N_399,N_531);
and U873 (N_873,N_70,N_18);
nand U874 (N_874,N_739,N_396);
nand U875 (N_875,N_378,N_179);
xor U876 (N_876,N_62,N_645);
nor U877 (N_877,N_390,N_660);
nor U878 (N_878,N_242,N_303);
nor U879 (N_879,N_198,N_357);
nand U880 (N_880,N_701,N_490);
nor U881 (N_881,N_397,N_34);
nand U882 (N_882,N_327,N_685);
nand U883 (N_883,N_263,N_283);
and U884 (N_884,N_604,N_194);
xnor U885 (N_885,N_228,N_417);
or U886 (N_886,N_31,N_441);
or U887 (N_887,N_253,N_359);
and U888 (N_888,N_117,N_483);
xnor U889 (N_889,N_135,N_669);
and U890 (N_890,N_442,N_697);
nand U891 (N_891,N_589,N_254);
nand U892 (N_892,N_223,N_366);
nand U893 (N_893,N_494,N_257);
and U894 (N_894,N_395,N_279);
and U895 (N_895,N_745,N_319);
and U896 (N_896,N_173,N_394);
nand U897 (N_897,N_385,N_575);
nor U898 (N_898,N_69,N_568);
nand U899 (N_899,N_577,N_111);
and U900 (N_900,N_671,N_643);
nor U901 (N_901,N_302,N_690);
nor U902 (N_902,N_152,N_175);
or U903 (N_903,N_608,N_247);
or U904 (N_904,N_516,N_633);
or U905 (N_905,N_4,N_248);
or U906 (N_906,N_15,N_317);
nor U907 (N_907,N_549,N_90);
nor U908 (N_908,N_68,N_96);
or U909 (N_909,N_502,N_722);
xor U910 (N_910,N_83,N_299);
nor U911 (N_911,N_649,N_526);
or U912 (N_912,N_108,N_41);
or U913 (N_913,N_560,N_414);
or U914 (N_914,N_519,N_95);
nor U915 (N_915,N_177,N_706);
nor U916 (N_916,N_474,N_740);
and U917 (N_917,N_689,N_55);
xor U918 (N_918,N_698,N_459);
and U919 (N_919,N_453,N_205);
or U920 (N_920,N_400,N_333);
nand U921 (N_921,N_478,N_261);
nor U922 (N_922,N_479,N_436);
nor U923 (N_923,N_141,N_592);
and U924 (N_924,N_321,N_244);
nand U925 (N_925,N_507,N_113);
nor U926 (N_926,N_445,N_692);
xor U927 (N_927,N_727,N_518);
and U928 (N_928,N_229,N_749);
nor U929 (N_929,N_408,N_422);
nor U930 (N_930,N_217,N_471);
nor U931 (N_931,N_11,N_433);
xnor U932 (N_932,N_741,N_285);
or U933 (N_933,N_123,N_144);
or U934 (N_934,N_610,N_291);
and U935 (N_935,N_252,N_384);
xnor U936 (N_936,N_465,N_707);
xor U937 (N_937,N_460,N_573);
and U938 (N_938,N_590,N_340);
or U939 (N_939,N_547,N_714);
nand U940 (N_940,N_712,N_403);
xnor U941 (N_941,N_582,N_668);
xnor U942 (N_942,N_501,N_172);
and U943 (N_943,N_218,N_383);
nand U944 (N_944,N_176,N_391);
nor U945 (N_945,N_365,N_622);
or U946 (N_946,N_125,N_324);
xnor U947 (N_947,N_377,N_656);
xor U948 (N_948,N_301,N_210);
xnor U949 (N_949,N_530,N_315);
and U950 (N_950,N_579,N_129);
and U951 (N_951,N_726,N_473);
xnor U952 (N_952,N_634,N_325);
xor U953 (N_953,N_61,N_28);
and U954 (N_954,N_139,N_189);
or U955 (N_955,N_619,N_670);
and U956 (N_956,N_47,N_613);
nor U957 (N_957,N_27,N_666);
nor U958 (N_958,N_50,N_734);
xor U959 (N_959,N_421,N_620);
or U960 (N_960,N_617,N_153);
nand U961 (N_961,N_353,N_686);
nor U962 (N_962,N_7,N_67);
xnor U963 (N_963,N_89,N_273);
nor U964 (N_964,N_259,N_274);
or U965 (N_965,N_480,N_630);
and U966 (N_966,N_43,N_444);
xor U967 (N_967,N_430,N_372);
nor U968 (N_968,N_493,N_600);
nand U969 (N_969,N_54,N_413);
or U970 (N_970,N_53,N_160);
xnor U971 (N_971,N_611,N_17);
xor U972 (N_972,N_336,N_463);
and U973 (N_973,N_541,N_659);
and U974 (N_974,N_149,N_386);
nor U975 (N_975,N_642,N_22);
xnor U976 (N_976,N_535,N_419);
xnor U977 (N_977,N_352,N_529);
nor U978 (N_978,N_38,N_286);
and U979 (N_979,N_348,N_744);
nand U980 (N_980,N_401,N_675);
nand U981 (N_981,N_499,N_558);
and U982 (N_982,N_23,N_688);
and U983 (N_983,N_381,N_180);
or U984 (N_984,N_418,N_567);
or U985 (N_985,N_525,N_367);
and U986 (N_986,N_628,N_468);
nand U987 (N_987,N_306,N_615);
xor U988 (N_988,N_335,N_548);
nor U989 (N_989,N_329,N_536);
and U990 (N_990,N_371,N_358);
nand U991 (N_991,N_624,N_102);
xnor U992 (N_992,N_59,N_713);
nand U993 (N_993,N_646,N_435);
or U994 (N_994,N_44,N_79);
nor U995 (N_995,N_166,N_195);
nand U996 (N_996,N_45,N_718);
nor U997 (N_997,N_674,N_98);
xor U998 (N_998,N_167,N_209);
nand U999 (N_999,N_215,N_241);
nor U1000 (N_1000,N_292,N_364);
nand U1001 (N_1001,N_747,N_537);
nand U1002 (N_1002,N_504,N_316);
or U1003 (N_1003,N_124,N_693);
nand U1004 (N_1004,N_48,N_388);
nor U1005 (N_1005,N_201,N_503);
nand U1006 (N_1006,N_598,N_122);
nand U1007 (N_1007,N_556,N_562);
or U1008 (N_1008,N_57,N_294);
xor U1009 (N_1009,N_185,N_488);
nand U1010 (N_1010,N_10,N_346);
or U1011 (N_1011,N_679,N_262);
nand U1012 (N_1012,N_276,N_162);
nor U1013 (N_1013,N_514,N_32);
xor U1014 (N_1014,N_412,N_143);
and U1015 (N_1015,N_337,N_565);
and U1016 (N_1016,N_591,N_542);
nor U1017 (N_1017,N_164,N_627);
xor U1018 (N_1018,N_545,N_270);
xor U1019 (N_1019,N_322,N_380);
nor U1020 (N_1020,N_571,N_12);
or U1021 (N_1021,N_496,N_282);
nand U1022 (N_1022,N_467,N_477);
nor U1023 (N_1023,N_0,N_458);
or U1024 (N_1024,N_437,N_578);
nand U1025 (N_1025,N_343,N_361);
and U1026 (N_1026,N_35,N_461);
nor U1027 (N_1027,N_677,N_440);
or U1028 (N_1028,N_126,N_328);
or U1029 (N_1029,N_603,N_543);
nand U1030 (N_1030,N_19,N_387);
nor U1031 (N_1031,N_199,N_100);
and U1032 (N_1032,N_51,N_532);
nand U1033 (N_1033,N_678,N_21);
nand U1034 (N_1034,N_644,N_190);
and U1035 (N_1035,N_527,N_33);
or U1036 (N_1036,N_416,N_318);
or U1037 (N_1037,N_136,N_245);
or U1038 (N_1038,N_312,N_235);
nand U1039 (N_1039,N_574,N_551);
xnor U1040 (N_1040,N_517,N_552);
xor U1041 (N_1041,N_676,N_226);
xnor U1042 (N_1042,N_580,N_331);
nor U1043 (N_1043,N_298,N_206);
nand U1044 (N_1044,N_599,N_520);
nand U1045 (N_1045,N_91,N_56);
and U1046 (N_1046,N_484,N_550);
xor U1047 (N_1047,N_700,N_426);
nand U1048 (N_1048,N_725,N_439);
or U1049 (N_1049,N_243,N_506);
nor U1050 (N_1050,N_428,N_154);
xnor U1051 (N_1051,N_544,N_510);
or U1052 (N_1052,N_76,N_233);
nor U1053 (N_1053,N_635,N_216);
xor U1054 (N_1054,N_80,N_184);
xnor U1055 (N_1055,N_392,N_131);
and U1056 (N_1056,N_404,N_449);
nand U1057 (N_1057,N_112,N_63);
nor U1058 (N_1058,N_341,N_77);
nand U1059 (N_1059,N_492,N_563);
nor U1060 (N_1060,N_188,N_104);
nor U1061 (N_1061,N_719,N_182);
or U1062 (N_1062,N_729,N_230);
and U1063 (N_1063,N_196,N_521);
and U1064 (N_1064,N_557,N_280);
or U1065 (N_1065,N_355,N_737);
or U1066 (N_1066,N_305,N_509);
nand U1067 (N_1067,N_597,N_52);
nand U1068 (N_1068,N_326,N_476);
and U1069 (N_1069,N_423,N_487);
and U1070 (N_1070,N_271,N_178);
nor U1071 (N_1071,N_411,N_710);
xnor U1072 (N_1072,N_410,N_625);
and U1073 (N_1073,N_640,N_268);
and U1074 (N_1074,N_105,N_6);
nand U1075 (N_1075,N_193,N_171);
or U1076 (N_1076,N_664,N_438);
and U1077 (N_1077,N_101,N_609);
and U1078 (N_1078,N_515,N_351);
or U1079 (N_1079,N_14,N_447);
nor U1080 (N_1080,N_214,N_9);
and U1081 (N_1081,N_191,N_338);
or U1082 (N_1082,N_402,N_288);
xnor U1083 (N_1083,N_200,N_497);
xor U1084 (N_1084,N_71,N_146);
nor U1085 (N_1085,N_522,N_728);
or U1086 (N_1086,N_731,N_491);
or U1087 (N_1087,N_300,N_554);
or U1088 (N_1088,N_258,N_420);
xor U1089 (N_1089,N_626,N_538);
nor U1090 (N_1090,N_717,N_566);
xnor U1091 (N_1091,N_602,N_431);
or U1092 (N_1092,N_572,N_709);
and U1093 (N_1093,N_652,N_694);
nor U1094 (N_1094,N_673,N_1);
nor U1095 (N_1095,N_237,N_87);
xnor U1096 (N_1096,N_738,N_239);
nor U1097 (N_1097,N_78,N_120);
and U1098 (N_1098,N_621,N_186);
nand U1099 (N_1099,N_581,N_695);
nor U1100 (N_1100,N_716,N_593);
nand U1101 (N_1101,N_211,N_379);
nand U1102 (N_1102,N_498,N_735);
nor U1103 (N_1103,N_165,N_730);
and U1104 (N_1104,N_405,N_170);
nand U1105 (N_1105,N_224,N_73);
nand U1106 (N_1106,N_207,N_296);
nand U1107 (N_1107,N_103,N_569);
and U1108 (N_1108,N_576,N_594);
nor U1109 (N_1109,N_667,N_342);
nand U1110 (N_1110,N_495,N_347);
nand U1111 (N_1111,N_636,N_407);
nor U1112 (N_1112,N_533,N_289);
or U1113 (N_1113,N_702,N_406);
nor U1114 (N_1114,N_539,N_696);
or U1115 (N_1115,N_434,N_489);
xnor U1116 (N_1116,N_470,N_260);
xnor U1117 (N_1117,N_232,N_650);
nand U1118 (N_1118,N_134,N_369);
or U1119 (N_1119,N_3,N_446);
nor U1120 (N_1120,N_72,N_349);
or U1121 (N_1121,N_250,N_249);
nand U1122 (N_1122,N_464,N_665);
nand U1123 (N_1123,N_682,N_109);
or U1124 (N_1124,N_99,N_632);
and U1125 (N_1125,N_104,N_219);
nor U1126 (N_1126,N_717,N_318);
nor U1127 (N_1127,N_423,N_507);
or U1128 (N_1128,N_617,N_274);
xor U1129 (N_1129,N_699,N_452);
and U1130 (N_1130,N_480,N_598);
and U1131 (N_1131,N_284,N_214);
nand U1132 (N_1132,N_135,N_723);
and U1133 (N_1133,N_336,N_167);
nor U1134 (N_1134,N_422,N_31);
and U1135 (N_1135,N_357,N_516);
and U1136 (N_1136,N_460,N_142);
and U1137 (N_1137,N_602,N_492);
and U1138 (N_1138,N_455,N_564);
xor U1139 (N_1139,N_594,N_729);
nand U1140 (N_1140,N_156,N_147);
and U1141 (N_1141,N_540,N_200);
nor U1142 (N_1142,N_265,N_746);
nor U1143 (N_1143,N_515,N_658);
nor U1144 (N_1144,N_734,N_66);
nand U1145 (N_1145,N_335,N_84);
nor U1146 (N_1146,N_87,N_100);
nor U1147 (N_1147,N_133,N_568);
or U1148 (N_1148,N_667,N_106);
nand U1149 (N_1149,N_290,N_442);
or U1150 (N_1150,N_669,N_428);
nor U1151 (N_1151,N_77,N_710);
or U1152 (N_1152,N_409,N_176);
and U1153 (N_1153,N_396,N_103);
xnor U1154 (N_1154,N_270,N_133);
and U1155 (N_1155,N_411,N_103);
xor U1156 (N_1156,N_175,N_72);
and U1157 (N_1157,N_10,N_378);
nand U1158 (N_1158,N_342,N_35);
or U1159 (N_1159,N_165,N_621);
nor U1160 (N_1160,N_701,N_225);
nor U1161 (N_1161,N_337,N_14);
nand U1162 (N_1162,N_195,N_202);
and U1163 (N_1163,N_438,N_202);
xor U1164 (N_1164,N_127,N_512);
or U1165 (N_1165,N_424,N_587);
or U1166 (N_1166,N_610,N_59);
or U1167 (N_1167,N_662,N_217);
nand U1168 (N_1168,N_37,N_409);
nor U1169 (N_1169,N_255,N_43);
nand U1170 (N_1170,N_496,N_487);
nand U1171 (N_1171,N_306,N_217);
or U1172 (N_1172,N_186,N_390);
xnor U1173 (N_1173,N_525,N_124);
or U1174 (N_1174,N_649,N_94);
nand U1175 (N_1175,N_687,N_386);
xor U1176 (N_1176,N_386,N_44);
and U1177 (N_1177,N_392,N_166);
nand U1178 (N_1178,N_462,N_453);
or U1179 (N_1179,N_149,N_710);
xor U1180 (N_1180,N_258,N_34);
and U1181 (N_1181,N_705,N_382);
nor U1182 (N_1182,N_598,N_78);
or U1183 (N_1183,N_521,N_480);
and U1184 (N_1184,N_628,N_313);
or U1185 (N_1185,N_526,N_639);
xnor U1186 (N_1186,N_226,N_558);
xnor U1187 (N_1187,N_381,N_653);
and U1188 (N_1188,N_669,N_307);
nor U1189 (N_1189,N_440,N_551);
xor U1190 (N_1190,N_594,N_608);
or U1191 (N_1191,N_22,N_666);
or U1192 (N_1192,N_637,N_80);
and U1193 (N_1193,N_670,N_403);
or U1194 (N_1194,N_362,N_644);
or U1195 (N_1195,N_491,N_377);
or U1196 (N_1196,N_23,N_424);
nand U1197 (N_1197,N_1,N_618);
xnor U1198 (N_1198,N_560,N_586);
and U1199 (N_1199,N_143,N_553);
nor U1200 (N_1200,N_681,N_45);
nand U1201 (N_1201,N_713,N_387);
and U1202 (N_1202,N_406,N_293);
nor U1203 (N_1203,N_714,N_668);
xnor U1204 (N_1204,N_133,N_36);
nor U1205 (N_1205,N_22,N_695);
and U1206 (N_1206,N_595,N_116);
and U1207 (N_1207,N_532,N_246);
and U1208 (N_1208,N_727,N_677);
nor U1209 (N_1209,N_520,N_171);
and U1210 (N_1210,N_179,N_675);
xnor U1211 (N_1211,N_344,N_117);
xnor U1212 (N_1212,N_239,N_500);
nand U1213 (N_1213,N_227,N_386);
xnor U1214 (N_1214,N_250,N_31);
xor U1215 (N_1215,N_518,N_498);
or U1216 (N_1216,N_663,N_84);
and U1217 (N_1217,N_510,N_602);
nand U1218 (N_1218,N_348,N_590);
xnor U1219 (N_1219,N_674,N_357);
and U1220 (N_1220,N_430,N_130);
nor U1221 (N_1221,N_360,N_657);
and U1222 (N_1222,N_139,N_123);
nand U1223 (N_1223,N_69,N_244);
or U1224 (N_1224,N_459,N_63);
nor U1225 (N_1225,N_86,N_207);
and U1226 (N_1226,N_459,N_26);
xor U1227 (N_1227,N_701,N_621);
xnor U1228 (N_1228,N_604,N_504);
nor U1229 (N_1229,N_209,N_623);
xnor U1230 (N_1230,N_549,N_302);
xnor U1231 (N_1231,N_595,N_327);
or U1232 (N_1232,N_459,N_101);
nand U1233 (N_1233,N_146,N_413);
nor U1234 (N_1234,N_51,N_2);
nor U1235 (N_1235,N_732,N_669);
and U1236 (N_1236,N_700,N_27);
nor U1237 (N_1237,N_128,N_564);
nor U1238 (N_1238,N_380,N_622);
and U1239 (N_1239,N_21,N_605);
xnor U1240 (N_1240,N_447,N_99);
xnor U1241 (N_1241,N_1,N_304);
or U1242 (N_1242,N_580,N_462);
and U1243 (N_1243,N_685,N_745);
nand U1244 (N_1244,N_553,N_3);
xnor U1245 (N_1245,N_341,N_558);
or U1246 (N_1246,N_105,N_114);
nor U1247 (N_1247,N_89,N_392);
xnor U1248 (N_1248,N_746,N_209);
nand U1249 (N_1249,N_690,N_277);
nor U1250 (N_1250,N_183,N_518);
nor U1251 (N_1251,N_61,N_176);
nand U1252 (N_1252,N_350,N_740);
or U1253 (N_1253,N_259,N_279);
or U1254 (N_1254,N_621,N_57);
nor U1255 (N_1255,N_363,N_669);
or U1256 (N_1256,N_358,N_179);
xor U1257 (N_1257,N_452,N_355);
xor U1258 (N_1258,N_578,N_538);
nand U1259 (N_1259,N_536,N_413);
xor U1260 (N_1260,N_51,N_519);
xor U1261 (N_1261,N_181,N_582);
or U1262 (N_1262,N_691,N_462);
nand U1263 (N_1263,N_66,N_701);
or U1264 (N_1264,N_344,N_563);
and U1265 (N_1265,N_444,N_743);
or U1266 (N_1266,N_581,N_178);
nor U1267 (N_1267,N_606,N_688);
nor U1268 (N_1268,N_425,N_628);
and U1269 (N_1269,N_26,N_563);
nand U1270 (N_1270,N_24,N_234);
or U1271 (N_1271,N_300,N_494);
nor U1272 (N_1272,N_747,N_287);
or U1273 (N_1273,N_704,N_747);
nand U1274 (N_1274,N_608,N_563);
xnor U1275 (N_1275,N_608,N_616);
nor U1276 (N_1276,N_631,N_601);
nor U1277 (N_1277,N_728,N_290);
nor U1278 (N_1278,N_539,N_353);
nor U1279 (N_1279,N_487,N_377);
nor U1280 (N_1280,N_130,N_725);
and U1281 (N_1281,N_621,N_35);
or U1282 (N_1282,N_217,N_360);
xnor U1283 (N_1283,N_421,N_17);
nand U1284 (N_1284,N_612,N_446);
xor U1285 (N_1285,N_498,N_647);
nand U1286 (N_1286,N_194,N_485);
xnor U1287 (N_1287,N_21,N_363);
xor U1288 (N_1288,N_643,N_91);
nor U1289 (N_1289,N_264,N_413);
nor U1290 (N_1290,N_242,N_572);
xnor U1291 (N_1291,N_333,N_384);
and U1292 (N_1292,N_676,N_186);
xnor U1293 (N_1293,N_403,N_508);
nand U1294 (N_1294,N_481,N_391);
xnor U1295 (N_1295,N_554,N_708);
nand U1296 (N_1296,N_734,N_9);
and U1297 (N_1297,N_587,N_124);
nand U1298 (N_1298,N_35,N_146);
nor U1299 (N_1299,N_165,N_73);
or U1300 (N_1300,N_227,N_501);
and U1301 (N_1301,N_153,N_740);
xnor U1302 (N_1302,N_578,N_499);
and U1303 (N_1303,N_430,N_684);
xnor U1304 (N_1304,N_272,N_120);
nor U1305 (N_1305,N_506,N_342);
and U1306 (N_1306,N_637,N_429);
xnor U1307 (N_1307,N_145,N_402);
and U1308 (N_1308,N_107,N_458);
nor U1309 (N_1309,N_565,N_21);
and U1310 (N_1310,N_150,N_102);
or U1311 (N_1311,N_192,N_437);
nand U1312 (N_1312,N_415,N_341);
nor U1313 (N_1313,N_741,N_178);
and U1314 (N_1314,N_162,N_451);
xnor U1315 (N_1315,N_166,N_500);
and U1316 (N_1316,N_56,N_642);
xor U1317 (N_1317,N_70,N_47);
or U1318 (N_1318,N_474,N_566);
or U1319 (N_1319,N_346,N_624);
nand U1320 (N_1320,N_596,N_74);
nor U1321 (N_1321,N_165,N_525);
nor U1322 (N_1322,N_589,N_311);
xor U1323 (N_1323,N_41,N_525);
nand U1324 (N_1324,N_301,N_9);
or U1325 (N_1325,N_737,N_315);
nand U1326 (N_1326,N_648,N_193);
and U1327 (N_1327,N_627,N_124);
nor U1328 (N_1328,N_404,N_442);
xnor U1329 (N_1329,N_597,N_332);
nand U1330 (N_1330,N_45,N_394);
nor U1331 (N_1331,N_491,N_388);
or U1332 (N_1332,N_77,N_430);
nand U1333 (N_1333,N_296,N_693);
nor U1334 (N_1334,N_11,N_743);
nand U1335 (N_1335,N_13,N_747);
nor U1336 (N_1336,N_248,N_313);
nor U1337 (N_1337,N_458,N_277);
and U1338 (N_1338,N_147,N_353);
and U1339 (N_1339,N_445,N_621);
and U1340 (N_1340,N_9,N_343);
xor U1341 (N_1341,N_529,N_2);
or U1342 (N_1342,N_318,N_142);
nor U1343 (N_1343,N_226,N_361);
or U1344 (N_1344,N_199,N_410);
xnor U1345 (N_1345,N_147,N_455);
and U1346 (N_1346,N_530,N_708);
xor U1347 (N_1347,N_632,N_201);
xor U1348 (N_1348,N_492,N_434);
and U1349 (N_1349,N_465,N_742);
or U1350 (N_1350,N_233,N_178);
or U1351 (N_1351,N_178,N_195);
xor U1352 (N_1352,N_593,N_15);
and U1353 (N_1353,N_47,N_588);
or U1354 (N_1354,N_440,N_402);
nand U1355 (N_1355,N_571,N_27);
nor U1356 (N_1356,N_414,N_234);
xor U1357 (N_1357,N_529,N_477);
or U1358 (N_1358,N_536,N_582);
nand U1359 (N_1359,N_644,N_119);
nor U1360 (N_1360,N_189,N_117);
and U1361 (N_1361,N_732,N_554);
xor U1362 (N_1362,N_749,N_474);
nor U1363 (N_1363,N_32,N_436);
nand U1364 (N_1364,N_463,N_78);
and U1365 (N_1365,N_677,N_378);
nand U1366 (N_1366,N_240,N_727);
nor U1367 (N_1367,N_520,N_376);
nand U1368 (N_1368,N_561,N_68);
or U1369 (N_1369,N_373,N_35);
nand U1370 (N_1370,N_290,N_580);
nor U1371 (N_1371,N_40,N_679);
and U1372 (N_1372,N_358,N_622);
xnor U1373 (N_1373,N_644,N_4);
xor U1374 (N_1374,N_204,N_180);
xor U1375 (N_1375,N_271,N_227);
nor U1376 (N_1376,N_637,N_65);
xor U1377 (N_1377,N_606,N_370);
and U1378 (N_1378,N_175,N_739);
and U1379 (N_1379,N_246,N_23);
or U1380 (N_1380,N_457,N_129);
and U1381 (N_1381,N_547,N_191);
nor U1382 (N_1382,N_485,N_83);
nand U1383 (N_1383,N_607,N_284);
nand U1384 (N_1384,N_160,N_321);
nand U1385 (N_1385,N_250,N_282);
nor U1386 (N_1386,N_543,N_214);
and U1387 (N_1387,N_347,N_309);
nand U1388 (N_1388,N_196,N_32);
nand U1389 (N_1389,N_313,N_239);
xnor U1390 (N_1390,N_418,N_244);
xor U1391 (N_1391,N_621,N_680);
nand U1392 (N_1392,N_499,N_71);
and U1393 (N_1393,N_52,N_236);
and U1394 (N_1394,N_59,N_410);
nor U1395 (N_1395,N_361,N_444);
xor U1396 (N_1396,N_275,N_32);
nor U1397 (N_1397,N_313,N_452);
nor U1398 (N_1398,N_110,N_551);
xor U1399 (N_1399,N_301,N_516);
nand U1400 (N_1400,N_506,N_89);
or U1401 (N_1401,N_263,N_351);
or U1402 (N_1402,N_643,N_291);
nand U1403 (N_1403,N_655,N_146);
nor U1404 (N_1404,N_147,N_529);
nand U1405 (N_1405,N_500,N_477);
nor U1406 (N_1406,N_230,N_301);
or U1407 (N_1407,N_198,N_135);
xor U1408 (N_1408,N_740,N_166);
nor U1409 (N_1409,N_445,N_271);
xnor U1410 (N_1410,N_290,N_570);
nand U1411 (N_1411,N_298,N_170);
nor U1412 (N_1412,N_434,N_215);
nand U1413 (N_1413,N_118,N_227);
and U1414 (N_1414,N_560,N_191);
nand U1415 (N_1415,N_533,N_448);
nor U1416 (N_1416,N_242,N_96);
and U1417 (N_1417,N_340,N_482);
nor U1418 (N_1418,N_178,N_84);
or U1419 (N_1419,N_340,N_76);
nand U1420 (N_1420,N_693,N_13);
nor U1421 (N_1421,N_274,N_526);
nand U1422 (N_1422,N_190,N_267);
or U1423 (N_1423,N_101,N_699);
and U1424 (N_1424,N_122,N_442);
nor U1425 (N_1425,N_215,N_480);
nand U1426 (N_1426,N_623,N_451);
and U1427 (N_1427,N_108,N_425);
nor U1428 (N_1428,N_265,N_116);
nor U1429 (N_1429,N_726,N_199);
xnor U1430 (N_1430,N_6,N_442);
xnor U1431 (N_1431,N_599,N_622);
nand U1432 (N_1432,N_320,N_216);
nand U1433 (N_1433,N_48,N_693);
nand U1434 (N_1434,N_553,N_441);
xor U1435 (N_1435,N_385,N_657);
and U1436 (N_1436,N_55,N_598);
nor U1437 (N_1437,N_384,N_344);
and U1438 (N_1438,N_404,N_266);
nor U1439 (N_1439,N_543,N_296);
xnor U1440 (N_1440,N_213,N_259);
nor U1441 (N_1441,N_29,N_543);
nor U1442 (N_1442,N_637,N_292);
or U1443 (N_1443,N_474,N_155);
and U1444 (N_1444,N_715,N_457);
nand U1445 (N_1445,N_428,N_111);
xor U1446 (N_1446,N_232,N_235);
or U1447 (N_1447,N_236,N_143);
nand U1448 (N_1448,N_424,N_413);
or U1449 (N_1449,N_333,N_203);
nor U1450 (N_1450,N_528,N_278);
nand U1451 (N_1451,N_534,N_426);
nand U1452 (N_1452,N_592,N_454);
or U1453 (N_1453,N_489,N_451);
and U1454 (N_1454,N_485,N_203);
and U1455 (N_1455,N_254,N_356);
nor U1456 (N_1456,N_131,N_736);
nor U1457 (N_1457,N_89,N_125);
or U1458 (N_1458,N_461,N_318);
nor U1459 (N_1459,N_451,N_688);
nand U1460 (N_1460,N_77,N_246);
nand U1461 (N_1461,N_12,N_615);
or U1462 (N_1462,N_100,N_297);
xnor U1463 (N_1463,N_733,N_507);
nand U1464 (N_1464,N_223,N_328);
or U1465 (N_1465,N_609,N_632);
xor U1466 (N_1466,N_82,N_352);
or U1467 (N_1467,N_695,N_508);
and U1468 (N_1468,N_489,N_264);
xor U1469 (N_1469,N_641,N_103);
nand U1470 (N_1470,N_747,N_741);
and U1471 (N_1471,N_697,N_144);
or U1472 (N_1472,N_292,N_466);
and U1473 (N_1473,N_13,N_622);
xnor U1474 (N_1474,N_14,N_267);
or U1475 (N_1475,N_314,N_556);
nand U1476 (N_1476,N_203,N_554);
nor U1477 (N_1477,N_167,N_309);
or U1478 (N_1478,N_353,N_83);
nand U1479 (N_1479,N_547,N_98);
xor U1480 (N_1480,N_519,N_482);
nand U1481 (N_1481,N_736,N_255);
xor U1482 (N_1482,N_550,N_259);
xnor U1483 (N_1483,N_613,N_82);
xnor U1484 (N_1484,N_265,N_402);
xnor U1485 (N_1485,N_451,N_312);
xor U1486 (N_1486,N_173,N_547);
and U1487 (N_1487,N_720,N_87);
nand U1488 (N_1488,N_214,N_712);
nand U1489 (N_1489,N_405,N_198);
nand U1490 (N_1490,N_697,N_298);
and U1491 (N_1491,N_573,N_260);
or U1492 (N_1492,N_739,N_543);
and U1493 (N_1493,N_162,N_563);
nor U1494 (N_1494,N_69,N_137);
or U1495 (N_1495,N_20,N_10);
nor U1496 (N_1496,N_700,N_592);
or U1497 (N_1497,N_309,N_517);
and U1498 (N_1498,N_531,N_21);
xnor U1499 (N_1499,N_703,N_334);
or U1500 (N_1500,N_1379,N_833);
nand U1501 (N_1501,N_992,N_803);
xnor U1502 (N_1502,N_1213,N_1432);
nand U1503 (N_1503,N_891,N_1318);
and U1504 (N_1504,N_1304,N_1003);
nor U1505 (N_1505,N_937,N_948);
nor U1506 (N_1506,N_1498,N_1325);
nor U1507 (N_1507,N_816,N_1152);
xnor U1508 (N_1508,N_962,N_1161);
xnor U1509 (N_1509,N_760,N_1065);
or U1510 (N_1510,N_1445,N_1074);
nand U1511 (N_1511,N_1350,N_1006);
xnor U1512 (N_1512,N_1156,N_1218);
or U1513 (N_1513,N_1020,N_1259);
or U1514 (N_1514,N_961,N_1334);
xor U1515 (N_1515,N_915,N_1396);
xnor U1516 (N_1516,N_936,N_767);
or U1517 (N_1517,N_1419,N_1321);
nand U1518 (N_1518,N_998,N_1060);
nor U1519 (N_1519,N_884,N_947);
nand U1520 (N_1520,N_861,N_1182);
and U1521 (N_1521,N_987,N_1464);
nand U1522 (N_1522,N_1028,N_974);
nand U1523 (N_1523,N_1437,N_1068);
xnor U1524 (N_1524,N_1211,N_1052);
or U1525 (N_1525,N_862,N_1133);
and U1526 (N_1526,N_818,N_864);
nand U1527 (N_1527,N_972,N_1064);
xor U1528 (N_1528,N_1271,N_1104);
nand U1529 (N_1529,N_1367,N_831);
xnor U1530 (N_1530,N_1188,N_1184);
and U1531 (N_1531,N_1115,N_1377);
nand U1532 (N_1532,N_1193,N_1401);
xnor U1533 (N_1533,N_958,N_1103);
xor U1534 (N_1534,N_1476,N_878);
nor U1535 (N_1535,N_868,N_999);
nand U1536 (N_1536,N_970,N_1411);
nand U1537 (N_1537,N_1100,N_805);
nor U1538 (N_1538,N_839,N_1235);
or U1539 (N_1539,N_979,N_777);
xnor U1540 (N_1540,N_1384,N_866);
xor U1541 (N_1541,N_1143,N_1314);
or U1542 (N_1542,N_1004,N_1059);
xor U1543 (N_1543,N_836,N_801);
nor U1544 (N_1544,N_1058,N_1335);
nor U1545 (N_1545,N_1478,N_1409);
nor U1546 (N_1546,N_1310,N_851);
nand U1547 (N_1547,N_847,N_953);
and U1548 (N_1548,N_896,N_1257);
xor U1549 (N_1549,N_1374,N_1390);
or U1550 (N_1550,N_1269,N_822);
or U1551 (N_1551,N_771,N_1410);
and U1552 (N_1552,N_931,N_1383);
or U1553 (N_1553,N_882,N_1078);
or U1554 (N_1554,N_911,N_1460);
and U1555 (N_1555,N_1395,N_1360);
nand U1556 (N_1556,N_770,N_967);
xor U1557 (N_1557,N_1424,N_1239);
or U1558 (N_1558,N_823,N_980);
and U1559 (N_1559,N_1479,N_1405);
nor U1560 (N_1560,N_1482,N_1340);
nand U1561 (N_1561,N_796,N_932);
xor U1562 (N_1562,N_1062,N_933);
nand U1563 (N_1563,N_892,N_1435);
nand U1564 (N_1564,N_905,N_874);
or U1565 (N_1565,N_834,N_1233);
and U1566 (N_1566,N_869,N_893);
xor U1567 (N_1567,N_988,N_842);
and U1568 (N_1568,N_957,N_1163);
or U1569 (N_1569,N_1418,N_1431);
xnor U1570 (N_1570,N_1346,N_1048);
and U1571 (N_1571,N_807,N_1167);
xor U1572 (N_1572,N_912,N_879);
nor U1573 (N_1573,N_1012,N_1180);
nand U1574 (N_1574,N_1046,N_1347);
and U1575 (N_1575,N_1324,N_850);
and U1576 (N_1576,N_759,N_786);
nor U1577 (N_1577,N_1242,N_757);
xor U1578 (N_1578,N_916,N_794);
nor U1579 (N_1579,N_873,N_1177);
or U1580 (N_1580,N_1047,N_806);
and U1581 (N_1581,N_855,N_1077);
or U1582 (N_1582,N_942,N_1311);
xnor U1583 (N_1583,N_1333,N_1372);
nor U1584 (N_1584,N_1034,N_930);
nand U1585 (N_1585,N_1015,N_1249);
and U1586 (N_1586,N_1356,N_1465);
nor U1587 (N_1587,N_1147,N_844);
and U1588 (N_1588,N_766,N_835);
or U1589 (N_1589,N_1237,N_872);
nor U1590 (N_1590,N_1394,N_1404);
and U1591 (N_1591,N_1490,N_1055);
nor U1592 (N_1592,N_1329,N_754);
or U1593 (N_1593,N_1274,N_1024);
nand U1594 (N_1594,N_1099,N_990);
nand U1595 (N_1595,N_1201,N_1290);
xor U1596 (N_1596,N_1270,N_1176);
and U1597 (N_1597,N_1284,N_966);
and U1598 (N_1598,N_1426,N_1328);
nor U1599 (N_1599,N_924,N_1462);
nand U1600 (N_1600,N_1477,N_1199);
and U1601 (N_1601,N_761,N_986);
or U1602 (N_1602,N_1191,N_1470);
nor U1603 (N_1603,N_787,N_824);
or U1604 (N_1604,N_1086,N_1150);
xnor U1605 (N_1605,N_1469,N_1122);
or U1606 (N_1606,N_1456,N_1491);
and U1607 (N_1607,N_1467,N_1054);
xor U1608 (N_1608,N_785,N_1095);
nor U1609 (N_1609,N_938,N_1175);
nor U1610 (N_1610,N_955,N_956);
and U1611 (N_1611,N_1309,N_1025);
and U1612 (N_1612,N_1185,N_1417);
nor U1613 (N_1613,N_1033,N_800);
nand U1614 (N_1614,N_929,N_1234);
nor U1615 (N_1615,N_849,N_1198);
nor U1616 (N_1616,N_1022,N_923);
and U1617 (N_1617,N_1348,N_1073);
nand U1618 (N_1618,N_1056,N_1407);
nor U1619 (N_1619,N_1101,N_1124);
and U1620 (N_1620,N_1219,N_809);
or U1621 (N_1621,N_1458,N_815);
xor U1622 (N_1622,N_1109,N_996);
and U1623 (N_1623,N_1111,N_1220);
nand U1624 (N_1624,N_994,N_1398);
and U1625 (N_1625,N_821,N_1297);
nand U1626 (N_1626,N_1131,N_1369);
nor U1627 (N_1627,N_1412,N_1416);
and U1628 (N_1628,N_1169,N_814);
or U1629 (N_1629,N_1359,N_913);
and U1630 (N_1630,N_1063,N_1238);
and U1631 (N_1631,N_1387,N_1388);
and U1632 (N_1632,N_1119,N_1051);
xor U1633 (N_1633,N_1391,N_969);
and U1634 (N_1634,N_1151,N_1089);
or U1635 (N_1635,N_812,N_925);
nand U1636 (N_1636,N_1082,N_1493);
or U1637 (N_1637,N_1438,N_830);
nor U1638 (N_1638,N_1113,N_1208);
xnor U1639 (N_1639,N_795,N_1475);
xnor U1640 (N_1640,N_858,N_1069);
or U1641 (N_1641,N_1040,N_1107);
xnor U1642 (N_1642,N_1164,N_1382);
or U1643 (N_1643,N_1230,N_837);
and U1644 (N_1644,N_1355,N_1322);
and U1645 (N_1645,N_1140,N_982);
xor U1646 (N_1646,N_1495,N_926);
nor U1647 (N_1647,N_1305,N_1466);
or U1648 (N_1648,N_1041,N_1031);
nand U1649 (N_1649,N_1053,N_776);
nand U1650 (N_1650,N_1275,N_1423);
nor U1651 (N_1651,N_897,N_825);
or U1652 (N_1652,N_1406,N_1102);
xnor U1653 (N_1653,N_1453,N_774);
nand U1654 (N_1654,N_1026,N_1029);
xnor U1655 (N_1655,N_1447,N_1168);
nor U1656 (N_1656,N_1291,N_1446);
xor U1657 (N_1657,N_1190,N_826);
or U1658 (N_1658,N_1017,N_1061);
and U1659 (N_1659,N_1158,N_1245);
xnor U1660 (N_1660,N_1076,N_960);
nand U1661 (N_1661,N_859,N_1299);
and U1662 (N_1662,N_920,N_1427);
nand U1663 (N_1663,N_1197,N_983);
nand U1664 (N_1664,N_1492,N_832);
or U1665 (N_1665,N_1452,N_1090);
nor U1666 (N_1666,N_1215,N_904);
nor U1667 (N_1667,N_1085,N_1016);
xor U1668 (N_1668,N_1186,N_1187);
xnor U1669 (N_1669,N_779,N_1358);
and U1670 (N_1670,N_1376,N_1231);
and U1671 (N_1671,N_944,N_1132);
or U1672 (N_1672,N_1232,N_1489);
nand U1673 (N_1673,N_798,N_921);
or U1674 (N_1674,N_1195,N_883);
nand U1675 (N_1675,N_993,N_1341);
nor U1676 (N_1676,N_1108,N_1472);
or U1677 (N_1677,N_764,N_1096);
nand U1678 (N_1678,N_1092,N_1018);
and U1679 (N_1679,N_1362,N_1281);
and U1680 (N_1680,N_1134,N_1455);
nor U1681 (N_1681,N_1414,N_1084);
nor U1682 (N_1682,N_1021,N_1389);
nor U1683 (N_1683,N_1166,N_1162);
nand U1684 (N_1684,N_1228,N_782);
xor U1685 (N_1685,N_1200,N_881);
and U1686 (N_1686,N_950,N_1212);
or U1687 (N_1687,N_750,N_804);
or U1688 (N_1688,N_1011,N_1287);
nor U1689 (N_1689,N_1364,N_841);
nand U1690 (N_1690,N_1045,N_783);
or U1691 (N_1691,N_1136,N_1146);
nand U1692 (N_1692,N_1392,N_1474);
nor U1693 (N_1693,N_1067,N_1248);
and U1694 (N_1694,N_1153,N_1300);
nor U1695 (N_1695,N_880,N_1128);
xor U1696 (N_1696,N_1327,N_808);
nand U1697 (N_1697,N_1043,N_863);
nor U1698 (N_1698,N_1430,N_1436);
or U1699 (N_1699,N_1293,N_791);
nand U1700 (N_1700,N_1352,N_1203);
nand U1701 (N_1701,N_1080,N_1373);
nor U1702 (N_1702,N_1137,N_1386);
xnor U1703 (N_1703,N_1170,N_829);
nand U1704 (N_1704,N_888,N_1266);
and U1705 (N_1705,N_852,N_810);
or U1706 (N_1706,N_778,N_952);
and U1707 (N_1707,N_1487,N_1339);
nor U1708 (N_1708,N_1255,N_1192);
xnor U1709 (N_1709,N_781,N_1038);
or U1710 (N_1710,N_934,N_1315);
xnor U1711 (N_1711,N_1267,N_1439);
and U1712 (N_1712,N_819,N_840);
xnor U1713 (N_1713,N_1091,N_811);
and U1714 (N_1714,N_1402,N_1443);
nor U1715 (N_1715,N_1178,N_901);
nand U1716 (N_1716,N_1308,N_946);
nand U1717 (N_1717,N_976,N_1292);
nand U1718 (N_1718,N_1205,N_963);
nor U1719 (N_1719,N_753,N_1121);
and U1720 (N_1720,N_789,N_1371);
or U1721 (N_1721,N_1194,N_1296);
xnor U1722 (N_1722,N_1425,N_1361);
or U1723 (N_1723,N_1112,N_1258);
nor U1724 (N_1724,N_1461,N_1349);
or U1725 (N_1725,N_964,N_1036);
nand U1726 (N_1726,N_1105,N_1142);
xnor U1727 (N_1727,N_828,N_1114);
xnor U1728 (N_1728,N_1481,N_1499);
and U1729 (N_1729,N_1283,N_1050);
or U1730 (N_1730,N_1210,N_1440);
and U1731 (N_1731,N_1110,N_954);
or U1732 (N_1732,N_1353,N_1268);
and U1733 (N_1733,N_1375,N_1366);
or U1734 (N_1734,N_894,N_1130);
nor U1735 (N_1735,N_793,N_1400);
or U1736 (N_1736,N_1144,N_752);
or U1737 (N_1737,N_856,N_1206);
or U1738 (N_1738,N_1254,N_1243);
xnor U1739 (N_1739,N_1256,N_1236);
xnor U1740 (N_1740,N_1301,N_1286);
nor U1741 (N_1741,N_1260,N_1485);
nand U1742 (N_1742,N_799,N_1240);
or U1743 (N_1743,N_1253,N_1035);
or U1744 (N_1744,N_941,N_1072);
xnor U1745 (N_1745,N_1363,N_1181);
xor U1746 (N_1746,N_1421,N_940);
nand U1747 (N_1747,N_875,N_1138);
nand U1748 (N_1748,N_1118,N_1368);
and U1749 (N_1749,N_977,N_1480);
and U1750 (N_1750,N_1316,N_1226);
or U1751 (N_1751,N_1032,N_927);
or U1752 (N_1752,N_1330,N_1393);
nand U1753 (N_1753,N_1019,N_939);
xor U1754 (N_1754,N_890,N_1399);
xor U1755 (N_1755,N_984,N_1039);
and U1756 (N_1756,N_1486,N_1223);
nand U1757 (N_1757,N_1380,N_1331);
and U1758 (N_1758,N_775,N_1098);
and U1759 (N_1759,N_1160,N_1488);
nor U1760 (N_1760,N_1428,N_1083);
and U1761 (N_1761,N_1494,N_1442);
nand U1762 (N_1762,N_1204,N_1042);
nor U1763 (N_1763,N_1273,N_1221);
or U1764 (N_1764,N_949,N_1450);
xor U1765 (N_1765,N_788,N_1433);
and U1766 (N_1766,N_1276,N_1277);
xnor U1767 (N_1767,N_889,N_1342);
and U1768 (N_1768,N_1295,N_772);
xnor U1769 (N_1769,N_1326,N_1357);
and U1770 (N_1770,N_1337,N_1454);
nor U1771 (N_1771,N_1149,N_1279);
xor U1772 (N_1772,N_928,N_1217);
xnor U1773 (N_1773,N_813,N_867);
xnor U1774 (N_1774,N_780,N_1189);
nor U1775 (N_1775,N_756,N_1225);
or U1776 (N_1776,N_973,N_1247);
or U1777 (N_1777,N_1145,N_1280);
nand U1778 (N_1778,N_995,N_802);
nor U1779 (N_1779,N_1007,N_1120);
nand U1780 (N_1780,N_945,N_1459);
nand U1781 (N_1781,N_1473,N_1264);
nor U1782 (N_1782,N_1323,N_1457);
or U1783 (N_1783,N_1252,N_1209);
or U1784 (N_1784,N_1282,N_755);
nor U1785 (N_1785,N_899,N_827);
nor U1786 (N_1786,N_975,N_1429);
or U1787 (N_1787,N_1251,N_854);
or U1788 (N_1788,N_1241,N_908);
xnor U1789 (N_1789,N_1449,N_959);
nand U1790 (N_1790,N_784,N_768);
nand U1791 (N_1791,N_1378,N_985);
xnor U1792 (N_1792,N_1227,N_1354);
xnor U1793 (N_1793,N_1001,N_1141);
or U1794 (N_1794,N_1183,N_1159);
nor U1795 (N_1795,N_997,N_1009);
or U1796 (N_1796,N_1312,N_1123);
nand U1797 (N_1797,N_1434,N_1126);
nand U1798 (N_1798,N_1117,N_1037);
nand U1799 (N_1799,N_1079,N_1013);
nor U1800 (N_1800,N_971,N_1154);
nand U1801 (N_1801,N_1484,N_1403);
and U1802 (N_1802,N_1351,N_885);
xor U1803 (N_1803,N_1313,N_838);
nand U1804 (N_1804,N_887,N_1422);
and U1805 (N_1805,N_902,N_871);
xnor U1806 (N_1806,N_1261,N_1246);
nor U1807 (N_1807,N_910,N_1179);
nand U1808 (N_1808,N_1049,N_765);
and U1809 (N_1809,N_758,N_886);
xor U1810 (N_1810,N_1173,N_817);
nor U1811 (N_1811,N_1030,N_876);
or U1812 (N_1812,N_1332,N_1262);
and U1813 (N_1813,N_1397,N_1066);
nor U1814 (N_1814,N_865,N_773);
or U1815 (N_1815,N_1288,N_918);
nand U1816 (N_1816,N_1345,N_1222);
xnor U1817 (N_1817,N_1165,N_1307);
xor U1818 (N_1818,N_1008,N_1289);
and U1819 (N_1819,N_1317,N_1302);
nand U1820 (N_1820,N_820,N_1000);
nor U1821 (N_1821,N_763,N_1448);
xor U1822 (N_1822,N_843,N_1306);
nand U1823 (N_1823,N_877,N_1127);
nand U1824 (N_1824,N_860,N_797);
xor U1825 (N_1825,N_1071,N_1135);
or U1826 (N_1826,N_1097,N_906);
or U1827 (N_1827,N_1497,N_1320);
xnor U1828 (N_1828,N_1172,N_1202);
or U1829 (N_1829,N_857,N_1088);
and U1830 (N_1830,N_968,N_845);
or U1831 (N_1831,N_1415,N_1044);
nor U1832 (N_1832,N_1214,N_1344);
xor U1833 (N_1833,N_1451,N_895);
xnor U1834 (N_1834,N_1370,N_1216);
nand U1835 (N_1835,N_846,N_1148);
or U1836 (N_1836,N_1116,N_909);
or U1837 (N_1837,N_1155,N_1196);
nor U1838 (N_1838,N_792,N_1094);
or U1839 (N_1839,N_870,N_1171);
or U1840 (N_1840,N_989,N_762);
nand U1841 (N_1841,N_1010,N_935);
or U1842 (N_1842,N_1278,N_1298);
xor U1843 (N_1843,N_1285,N_1413);
xnor U1844 (N_1844,N_1294,N_1075);
nand U1845 (N_1845,N_1139,N_790);
nand U1846 (N_1846,N_1157,N_1250);
or U1847 (N_1847,N_917,N_1265);
nor U1848 (N_1848,N_1005,N_1272);
and U1849 (N_1849,N_1023,N_1303);
or U1850 (N_1850,N_1125,N_922);
nand U1851 (N_1851,N_1129,N_1014);
or U1852 (N_1852,N_1463,N_1444);
and U1853 (N_1853,N_1057,N_951);
or U1854 (N_1854,N_1244,N_1093);
xor U1855 (N_1855,N_1381,N_1002);
xnor U1856 (N_1856,N_1319,N_898);
nor U1857 (N_1857,N_848,N_1468);
xor U1858 (N_1858,N_981,N_1385);
nand U1859 (N_1859,N_1420,N_1229);
or U1860 (N_1860,N_1263,N_978);
nand U1861 (N_1861,N_751,N_1070);
or U1862 (N_1862,N_907,N_769);
and U1863 (N_1863,N_1207,N_991);
and U1864 (N_1864,N_943,N_1471);
or U1865 (N_1865,N_903,N_1174);
xor U1866 (N_1866,N_1081,N_1027);
and U1867 (N_1867,N_1483,N_1336);
nor U1868 (N_1868,N_1343,N_1338);
nor U1869 (N_1869,N_965,N_914);
xnor U1870 (N_1870,N_919,N_1496);
nor U1871 (N_1871,N_1365,N_853);
and U1872 (N_1872,N_1224,N_1087);
xnor U1873 (N_1873,N_900,N_1106);
or U1874 (N_1874,N_1441,N_1408);
nor U1875 (N_1875,N_1477,N_754);
or U1876 (N_1876,N_1407,N_846);
or U1877 (N_1877,N_815,N_1210);
or U1878 (N_1878,N_1118,N_1361);
xnor U1879 (N_1879,N_922,N_1016);
nand U1880 (N_1880,N_1447,N_1081);
nand U1881 (N_1881,N_883,N_1366);
nor U1882 (N_1882,N_1312,N_1324);
xor U1883 (N_1883,N_994,N_1417);
nand U1884 (N_1884,N_1424,N_925);
nor U1885 (N_1885,N_1242,N_1175);
nor U1886 (N_1886,N_883,N_1003);
or U1887 (N_1887,N_1498,N_1454);
and U1888 (N_1888,N_885,N_1469);
xnor U1889 (N_1889,N_1028,N_1477);
nand U1890 (N_1890,N_1083,N_992);
or U1891 (N_1891,N_1082,N_1435);
or U1892 (N_1892,N_1327,N_983);
nand U1893 (N_1893,N_1230,N_857);
nand U1894 (N_1894,N_754,N_1443);
nand U1895 (N_1895,N_807,N_1043);
and U1896 (N_1896,N_930,N_1236);
nor U1897 (N_1897,N_1249,N_1152);
nor U1898 (N_1898,N_826,N_1266);
and U1899 (N_1899,N_1180,N_1176);
nor U1900 (N_1900,N_777,N_1196);
and U1901 (N_1901,N_971,N_1487);
xor U1902 (N_1902,N_1253,N_1339);
nand U1903 (N_1903,N_767,N_991);
and U1904 (N_1904,N_1279,N_1453);
nor U1905 (N_1905,N_1422,N_934);
and U1906 (N_1906,N_862,N_782);
xnor U1907 (N_1907,N_908,N_1358);
nor U1908 (N_1908,N_1408,N_1312);
and U1909 (N_1909,N_1087,N_1108);
and U1910 (N_1910,N_856,N_1017);
nor U1911 (N_1911,N_1112,N_1408);
nand U1912 (N_1912,N_993,N_1102);
or U1913 (N_1913,N_1366,N_806);
or U1914 (N_1914,N_1095,N_1236);
nor U1915 (N_1915,N_1252,N_1178);
nand U1916 (N_1916,N_985,N_1055);
and U1917 (N_1917,N_1007,N_832);
xor U1918 (N_1918,N_831,N_858);
xnor U1919 (N_1919,N_888,N_1196);
nand U1920 (N_1920,N_1311,N_762);
and U1921 (N_1921,N_879,N_1212);
nand U1922 (N_1922,N_836,N_1393);
nor U1923 (N_1923,N_936,N_1492);
nand U1924 (N_1924,N_751,N_986);
or U1925 (N_1925,N_800,N_786);
or U1926 (N_1926,N_984,N_1160);
and U1927 (N_1927,N_1361,N_898);
xor U1928 (N_1928,N_931,N_1049);
nand U1929 (N_1929,N_843,N_1189);
nand U1930 (N_1930,N_1361,N_1031);
nand U1931 (N_1931,N_1153,N_1357);
nor U1932 (N_1932,N_1092,N_1391);
and U1933 (N_1933,N_1362,N_1456);
nand U1934 (N_1934,N_834,N_1396);
nand U1935 (N_1935,N_1020,N_1482);
xnor U1936 (N_1936,N_1383,N_1405);
nor U1937 (N_1937,N_1410,N_1315);
and U1938 (N_1938,N_1269,N_1082);
and U1939 (N_1939,N_1477,N_1122);
and U1940 (N_1940,N_987,N_1115);
or U1941 (N_1941,N_884,N_1148);
xor U1942 (N_1942,N_885,N_1061);
nor U1943 (N_1943,N_1112,N_1102);
xnor U1944 (N_1944,N_1302,N_910);
and U1945 (N_1945,N_962,N_975);
and U1946 (N_1946,N_893,N_1035);
nor U1947 (N_1947,N_1416,N_1177);
nor U1948 (N_1948,N_1481,N_1168);
or U1949 (N_1949,N_847,N_799);
xnor U1950 (N_1950,N_1095,N_992);
or U1951 (N_1951,N_1027,N_999);
or U1952 (N_1952,N_1184,N_1221);
and U1953 (N_1953,N_1079,N_887);
nor U1954 (N_1954,N_1408,N_1263);
and U1955 (N_1955,N_1250,N_1432);
nand U1956 (N_1956,N_1284,N_1285);
or U1957 (N_1957,N_845,N_1023);
nand U1958 (N_1958,N_814,N_1471);
nand U1959 (N_1959,N_1384,N_1009);
and U1960 (N_1960,N_1040,N_1190);
xor U1961 (N_1961,N_1389,N_1026);
and U1962 (N_1962,N_1486,N_1073);
xor U1963 (N_1963,N_1027,N_1166);
nand U1964 (N_1964,N_1292,N_1245);
nand U1965 (N_1965,N_759,N_838);
nand U1966 (N_1966,N_1115,N_1367);
and U1967 (N_1967,N_1218,N_959);
and U1968 (N_1968,N_1271,N_941);
nor U1969 (N_1969,N_933,N_1423);
xor U1970 (N_1970,N_1428,N_1187);
nor U1971 (N_1971,N_1217,N_1083);
or U1972 (N_1972,N_896,N_1400);
and U1973 (N_1973,N_874,N_1138);
nand U1974 (N_1974,N_1048,N_1414);
nand U1975 (N_1975,N_1402,N_1195);
or U1976 (N_1976,N_1160,N_1496);
and U1977 (N_1977,N_836,N_756);
nor U1978 (N_1978,N_1064,N_1391);
or U1979 (N_1979,N_872,N_1082);
and U1980 (N_1980,N_1233,N_1121);
or U1981 (N_1981,N_1295,N_1009);
and U1982 (N_1982,N_1456,N_868);
xnor U1983 (N_1983,N_860,N_1063);
and U1984 (N_1984,N_1102,N_779);
and U1985 (N_1985,N_1293,N_933);
nand U1986 (N_1986,N_917,N_1097);
or U1987 (N_1987,N_1063,N_1366);
nor U1988 (N_1988,N_1419,N_999);
or U1989 (N_1989,N_985,N_1475);
nand U1990 (N_1990,N_889,N_1353);
or U1991 (N_1991,N_1143,N_1184);
xor U1992 (N_1992,N_1392,N_1104);
nand U1993 (N_1993,N_997,N_1084);
nor U1994 (N_1994,N_1130,N_1339);
nand U1995 (N_1995,N_1363,N_1037);
or U1996 (N_1996,N_869,N_785);
nand U1997 (N_1997,N_978,N_819);
and U1998 (N_1998,N_876,N_1393);
or U1999 (N_1999,N_1093,N_945);
and U2000 (N_2000,N_787,N_913);
xnor U2001 (N_2001,N_1336,N_1303);
nand U2002 (N_2002,N_1461,N_1251);
xor U2003 (N_2003,N_1253,N_1439);
or U2004 (N_2004,N_918,N_1227);
xnor U2005 (N_2005,N_1231,N_779);
xor U2006 (N_2006,N_975,N_1066);
nor U2007 (N_2007,N_1286,N_1050);
nor U2008 (N_2008,N_1048,N_1083);
or U2009 (N_2009,N_1181,N_1151);
nor U2010 (N_2010,N_1352,N_1028);
xor U2011 (N_2011,N_1197,N_838);
and U2012 (N_2012,N_1462,N_1149);
nor U2013 (N_2013,N_802,N_1364);
or U2014 (N_2014,N_1117,N_862);
xor U2015 (N_2015,N_1220,N_1202);
or U2016 (N_2016,N_1178,N_1147);
nand U2017 (N_2017,N_851,N_955);
xor U2018 (N_2018,N_1076,N_1188);
nand U2019 (N_2019,N_1103,N_890);
xnor U2020 (N_2020,N_1195,N_1047);
or U2021 (N_2021,N_1267,N_1124);
nor U2022 (N_2022,N_1428,N_1126);
and U2023 (N_2023,N_1261,N_841);
or U2024 (N_2024,N_1012,N_944);
or U2025 (N_2025,N_1094,N_1041);
or U2026 (N_2026,N_1050,N_1274);
nand U2027 (N_2027,N_1285,N_1040);
xor U2028 (N_2028,N_1169,N_1296);
xnor U2029 (N_2029,N_1342,N_1189);
and U2030 (N_2030,N_952,N_913);
nor U2031 (N_2031,N_1390,N_757);
and U2032 (N_2032,N_789,N_979);
nand U2033 (N_2033,N_1393,N_1015);
or U2034 (N_2034,N_943,N_1296);
nand U2035 (N_2035,N_1340,N_1176);
xnor U2036 (N_2036,N_1004,N_1107);
and U2037 (N_2037,N_1369,N_751);
xor U2038 (N_2038,N_1028,N_1264);
nand U2039 (N_2039,N_1035,N_1422);
and U2040 (N_2040,N_860,N_1019);
nand U2041 (N_2041,N_1193,N_1104);
and U2042 (N_2042,N_982,N_963);
and U2043 (N_2043,N_1238,N_1486);
xor U2044 (N_2044,N_1300,N_1351);
or U2045 (N_2045,N_1245,N_837);
and U2046 (N_2046,N_872,N_780);
nand U2047 (N_2047,N_1360,N_828);
and U2048 (N_2048,N_1074,N_1497);
and U2049 (N_2049,N_851,N_1315);
and U2050 (N_2050,N_1224,N_1277);
or U2051 (N_2051,N_1127,N_794);
or U2052 (N_2052,N_892,N_969);
nor U2053 (N_2053,N_1432,N_1263);
nand U2054 (N_2054,N_909,N_984);
or U2055 (N_2055,N_815,N_1327);
nand U2056 (N_2056,N_842,N_1224);
nand U2057 (N_2057,N_1057,N_1472);
nand U2058 (N_2058,N_1239,N_785);
nor U2059 (N_2059,N_814,N_994);
and U2060 (N_2060,N_1220,N_1316);
or U2061 (N_2061,N_1011,N_928);
nor U2062 (N_2062,N_770,N_1288);
nor U2063 (N_2063,N_1303,N_1018);
xor U2064 (N_2064,N_1249,N_1365);
xnor U2065 (N_2065,N_893,N_1153);
xor U2066 (N_2066,N_1026,N_1003);
nand U2067 (N_2067,N_1406,N_1291);
and U2068 (N_2068,N_1190,N_770);
nor U2069 (N_2069,N_1393,N_1006);
nor U2070 (N_2070,N_978,N_898);
or U2071 (N_2071,N_1225,N_1308);
and U2072 (N_2072,N_1221,N_1371);
and U2073 (N_2073,N_1404,N_1492);
nor U2074 (N_2074,N_1494,N_1128);
xor U2075 (N_2075,N_1333,N_766);
nor U2076 (N_2076,N_1117,N_1434);
nor U2077 (N_2077,N_1473,N_1249);
nand U2078 (N_2078,N_1431,N_803);
or U2079 (N_2079,N_1359,N_939);
xor U2080 (N_2080,N_1252,N_1421);
or U2081 (N_2081,N_944,N_905);
nor U2082 (N_2082,N_1455,N_909);
nand U2083 (N_2083,N_821,N_1275);
or U2084 (N_2084,N_1146,N_1215);
and U2085 (N_2085,N_832,N_888);
nand U2086 (N_2086,N_1003,N_1050);
xnor U2087 (N_2087,N_1447,N_1448);
and U2088 (N_2088,N_1055,N_822);
xor U2089 (N_2089,N_1216,N_1026);
and U2090 (N_2090,N_1168,N_792);
xnor U2091 (N_2091,N_1106,N_1477);
xnor U2092 (N_2092,N_1493,N_868);
or U2093 (N_2093,N_1185,N_1369);
nor U2094 (N_2094,N_1429,N_846);
nand U2095 (N_2095,N_1017,N_999);
and U2096 (N_2096,N_952,N_1175);
nor U2097 (N_2097,N_1038,N_1444);
or U2098 (N_2098,N_1178,N_985);
and U2099 (N_2099,N_956,N_1360);
or U2100 (N_2100,N_1029,N_887);
nand U2101 (N_2101,N_1229,N_779);
or U2102 (N_2102,N_1080,N_1310);
xor U2103 (N_2103,N_1383,N_1460);
nor U2104 (N_2104,N_1384,N_978);
nand U2105 (N_2105,N_855,N_1319);
and U2106 (N_2106,N_1402,N_1433);
and U2107 (N_2107,N_1406,N_1456);
xor U2108 (N_2108,N_1308,N_1216);
and U2109 (N_2109,N_1340,N_785);
and U2110 (N_2110,N_1298,N_1289);
nand U2111 (N_2111,N_1029,N_1058);
xor U2112 (N_2112,N_1047,N_914);
or U2113 (N_2113,N_1318,N_941);
and U2114 (N_2114,N_1328,N_988);
nor U2115 (N_2115,N_1366,N_824);
and U2116 (N_2116,N_1112,N_1294);
xor U2117 (N_2117,N_987,N_1155);
or U2118 (N_2118,N_1074,N_882);
nor U2119 (N_2119,N_1157,N_1100);
and U2120 (N_2120,N_1087,N_774);
nand U2121 (N_2121,N_1032,N_1205);
xnor U2122 (N_2122,N_1297,N_1180);
nor U2123 (N_2123,N_1257,N_1153);
nor U2124 (N_2124,N_1240,N_772);
nor U2125 (N_2125,N_891,N_1060);
and U2126 (N_2126,N_1292,N_1003);
or U2127 (N_2127,N_1444,N_1230);
xnor U2128 (N_2128,N_859,N_1035);
and U2129 (N_2129,N_1491,N_1137);
and U2130 (N_2130,N_772,N_910);
xnor U2131 (N_2131,N_1115,N_880);
nor U2132 (N_2132,N_1331,N_957);
nand U2133 (N_2133,N_879,N_1452);
or U2134 (N_2134,N_869,N_846);
nand U2135 (N_2135,N_1060,N_759);
or U2136 (N_2136,N_1048,N_1280);
or U2137 (N_2137,N_1219,N_1206);
or U2138 (N_2138,N_891,N_796);
and U2139 (N_2139,N_1305,N_792);
or U2140 (N_2140,N_854,N_1445);
xor U2141 (N_2141,N_1229,N_848);
nor U2142 (N_2142,N_765,N_870);
xor U2143 (N_2143,N_1446,N_1062);
nand U2144 (N_2144,N_1348,N_1462);
and U2145 (N_2145,N_847,N_1493);
nor U2146 (N_2146,N_1226,N_1096);
and U2147 (N_2147,N_1394,N_1106);
nand U2148 (N_2148,N_1319,N_1468);
and U2149 (N_2149,N_1168,N_816);
nor U2150 (N_2150,N_893,N_1374);
and U2151 (N_2151,N_869,N_804);
and U2152 (N_2152,N_846,N_953);
nor U2153 (N_2153,N_1480,N_918);
nand U2154 (N_2154,N_1332,N_754);
nor U2155 (N_2155,N_855,N_1226);
xor U2156 (N_2156,N_1065,N_866);
xor U2157 (N_2157,N_1378,N_1171);
nor U2158 (N_2158,N_880,N_873);
xor U2159 (N_2159,N_835,N_992);
and U2160 (N_2160,N_1284,N_1169);
xnor U2161 (N_2161,N_928,N_1484);
nor U2162 (N_2162,N_1417,N_819);
nand U2163 (N_2163,N_1137,N_866);
or U2164 (N_2164,N_1051,N_1455);
or U2165 (N_2165,N_906,N_1183);
nor U2166 (N_2166,N_1176,N_841);
or U2167 (N_2167,N_798,N_1288);
nor U2168 (N_2168,N_1219,N_1150);
and U2169 (N_2169,N_1407,N_1196);
nor U2170 (N_2170,N_1104,N_1171);
and U2171 (N_2171,N_1432,N_969);
nor U2172 (N_2172,N_751,N_1475);
or U2173 (N_2173,N_1256,N_1301);
nor U2174 (N_2174,N_938,N_1281);
or U2175 (N_2175,N_1348,N_884);
and U2176 (N_2176,N_1403,N_779);
nor U2177 (N_2177,N_904,N_1464);
and U2178 (N_2178,N_1132,N_1330);
and U2179 (N_2179,N_1173,N_882);
nor U2180 (N_2180,N_1117,N_869);
nand U2181 (N_2181,N_1179,N_1120);
xnor U2182 (N_2182,N_1047,N_1378);
or U2183 (N_2183,N_860,N_821);
and U2184 (N_2184,N_870,N_1227);
nand U2185 (N_2185,N_1427,N_1099);
xor U2186 (N_2186,N_1215,N_1148);
nand U2187 (N_2187,N_1271,N_766);
nor U2188 (N_2188,N_1421,N_1115);
xnor U2189 (N_2189,N_1352,N_896);
nor U2190 (N_2190,N_879,N_1105);
nor U2191 (N_2191,N_820,N_1177);
xnor U2192 (N_2192,N_1044,N_1223);
xnor U2193 (N_2193,N_995,N_1443);
nor U2194 (N_2194,N_808,N_945);
nand U2195 (N_2195,N_1292,N_772);
and U2196 (N_2196,N_752,N_1439);
nand U2197 (N_2197,N_1092,N_1241);
nand U2198 (N_2198,N_877,N_1269);
or U2199 (N_2199,N_1345,N_1299);
nor U2200 (N_2200,N_1194,N_1383);
nand U2201 (N_2201,N_1477,N_1446);
nor U2202 (N_2202,N_841,N_876);
nand U2203 (N_2203,N_1421,N_873);
nor U2204 (N_2204,N_947,N_1314);
or U2205 (N_2205,N_820,N_924);
nor U2206 (N_2206,N_1073,N_1431);
or U2207 (N_2207,N_815,N_861);
nand U2208 (N_2208,N_1202,N_1275);
nor U2209 (N_2209,N_918,N_1182);
or U2210 (N_2210,N_819,N_1311);
or U2211 (N_2211,N_964,N_814);
nor U2212 (N_2212,N_1395,N_854);
xor U2213 (N_2213,N_1426,N_1247);
or U2214 (N_2214,N_782,N_1007);
and U2215 (N_2215,N_1184,N_901);
nand U2216 (N_2216,N_769,N_1458);
nand U2217 (N_2217,N_1471,N_1180);
or U2218 (N_2218,N_1021,N_1161);
nand U2219 (N_2219,N_1120,N_1377);
nor U2220 (N_2220,N_1040,N_1348);
nor U2221 (N_2221,N_948,N_969);
and U2222 (N_2222,N_1401,N_919);
nor U2223 (N_2223,N_892,N_759);
xnor U2224 (N_2224,N_1362,N_1498);
nor U2225 (N_2225,N_976,N_983);
nand U2226 (N_2226,N_827,N_872);
xor U2227 (N_2227,N_968,N_1137);
nand U2228 (N_2228,N_997,N_1074);
or U2229 (N_2229,N_1128,N_1253);
nand U2230 (N_2230,N_1284,N_982);
xor U2231 (N_2231,N_1179,N_1080);
xnor U2232 (N_2232,N_1166,N_1481);
and U2233 (N_2233,N_759,N_1130);
or U2234 (N_2234,N_760,N_1210);
and U2235 (N_2235,N_1438,N_828);
nand U2236 (N_2236,N_995,N_885);
xor U2237 (N_2237,N_1472,N_976);
and U2238 (N_2238,N_1347,N_874);
and U2239 (N_2239,N_809,N_1146);
nor U2240 (N_2240,N_1351,N_1085);
or U2241 (N_2241,N_1303,N_829);
nor U2242 (N_2242,N_1439,N_798);
nor U2243 (N_2243,N_1133,N_1481);
or U2244 (N_2244,N_804,N_982);
nor U2245 (N_2245,N_758,N_847);
nand U2246 (N_2246,N_1486,N_833);
nor U2247 (N_2247,N_1133,N_859);
nand U2248 (N_2248,N_952,N_1337);
xnor U2249 (N_2249,N_1374,N_770);
nor U2250 (N_2250,N_2066,N_1557);
nand U2251 (N_2251,N_1649,N_1927);
and U2252 (N_2252,N_1513,N_2085);
xnor U2253 (N_2253,N_1634,N_1975);
xor U2254 (N_2254,N_1815,N_2121);
xor U2255 (N_2255,N_1753,N_2205);
and U2256 (N_2256,N_1705,N_1543);
nand U2257 (N_2257,N_1695,N_1841);
nor U2258 (N_2258,N_1702,N_2213);
and U2259 (N_2259,N_2130,N_1784);
or U2260 (N_2260,N_1908,N_1662);
nand U2261 (N_2261,N_1780,N_1777);
nor U2262 (N_2262,N_1934,N_1997);
and U2263 (N_2263,N_1607,N_1672);
xor U2264 (N_2264,N_1575,N_1597);
nand U2265 (N_2265,N_2062,N_1503);
nand U2266 (N_2266,N_1520,N_2026);
nor U2267 (N_2267,N_1576,N_1535);
nand U2268 (N_2268,N_1623,N_2200);
or U2269 (N_2269,N_2137,N_2091);
or U2270 (N_2270,N_1883,N_2183);
and U2271 (N_2271,N_1787,N_1963);
nor U2272 (N_2272,N_1831,N_2214);
xnor U2273 (N_2273,N_2078,N_1516);
nand U2274 (N_2274,N_1659,N_1585);
and U2275 (N_2275,N_1862,N_2049);
and U2276 (N_2276,N_1731,N_2207);
nand U2277 (N_2277,N_1986,N_1866);
xor U2278 (N_2278,N_1899,N_2015);
or U2279 (N_2279,N_1637,N_1707);
and U2280 (N_2280,N_1763,N_2054);
or U2281 (N_2281,N_1636,N_2225);
nand U2282 (N_2282,N_2055,N_2122);
xor U2283 (N_2283,N_1527,N_1727);
nand U2284 (N_2284,N_1999,N_2124);
nand U2285 (N_2285,N_2249,N_1948);
or U2286 (N_2286,N_1933,N_1626);
nand U2287 (N_2287,N_1788,N_2003);
xnor U2288 (N_2288,N_2136,N_2173);
nand U2289 (N_2289,N_1791,N_2140);
and U2290 (N_2290,N_1526,N_2228);
xnor U2291 (N_2291,N_2059,N_1656);
nand U2292 (N_2292,N_1762,N_1728);
or U2293 (N_2293,N_1589,N_2032);
or U2294 (N_2294,N_2029,N_2013);
xnor U2295 (N_2295,N_1742,N_1868);
nand U2296 (N_2296,N_1559,N_1772);
nand U2297 (N_2297,N_1698,N_1511);
nor U2298 (N_2298,N_1794,N_1587);
nor U2299 (N_2299,N_2219,N_2156);
nand U2300 (N_2300,N_1774,N_2119);
or U2301 (N_2301,N_1766,N_1798);
nand U2302 (N_2302,N_1936,N_1845);
xnor U2303 (N_2303,N_2113,N_1853);
or U2304 (N_2304,N_1850,N_2198);
nor U2305 (N_2305,N_1805,N_1972);
nor U2306 (N_2306,N_1800,N_1771);
xnor U2307 (N_2307,N_1680,N_1856);
or U2308 (N_2308,N_1758,N_1920);
or U2309 (N_2309,N_1951,N_1533);
xor U2310 (N_2310,N_1603,N_2114);
or U2311 (N_2311,N_1564,N_2157);
nand U2312 (N_2312,N_1956,N_1571);
and U2313 (N_2313,N_1631,N_1998);
xor U2314 (N_2314,N_2170,N_1736);
and U2315 (N_2315,N_1923,N_1692);
or U2316 (N_2316,N_1645,N_1994);
nor U2317 (N_2317,N_1669,N_1706);
nor U2318 (N_2318,N_1872,N_1593);
nor U2319 (N_2319,N_2144,N_1852);
nor U2320 (N_2320,N_2218,N_2036);
and U2321 (N_2321,N_1996,N_2152);
and U2322 (N_2322,N_1922,N_1945);
nand U2323 (N_2323,N_1717,N_2115);
nor U2324 (N_2324,N_2216,N_1653);
nand U2325 (N_2325,N_1847,N_2125);
nand U2326 (N_2326,N_1993,N_1870);
xnor U2327 (N_2327,N_2040,N_2084);
nand U2328 (N_2328,N_1688,N_2063);
or U2329 (N_2329,N_1573,N_1884);
nand U2330 (N_2330,N_1961,N_1666);
nor U2331 (N_2331,N_2155,N_1889);
nand U2332 (N_2332,N_2051,N_2068);
xnor U2333 (N_2333,N_2222,N_1854);
or U2334 (N_2334,N_2171,N_2175);
nand U2335 (N_2335,N_2240,N_1801);
nand U2336 (N_2336,N_2018,N_1646);
or U2337 (N_2337,N_1964,N_1861);
and U2338 (N_2338,N_1682,N_1925);
and U2339 (N_2339,N_1867,N_2025);
nor U2340 (N_2340,N_1594,N_1586);
nand U2341 (N_2341,N_1830,N_2165);
or U2342 (N_2342,N_1907,N_2038);
nor U2343 (N_2343,N_2077,N_2012);
and U2344 (N_2344,N_1745,N_1654);
xor U2345 (N_2345,N_2129,N_1882);
nand U2346 (N_2346,N_2166,N_1793);
nand U2347 (N_2347,N_1517,N_2224);
xor U2348 (N_2348,N_1877,N_2027);
nand U2349 (N_2349,N_1921,N_1592);
or U2350 (N_2350,N_1675,N_2209);
nor U2351 (N_2351,N_1690,N_1509);
and U2352 (N_2352,N_1844,N_1799);
and U2353 (N_2353,N_2094,N_1935);
and U2354 (N_2354,N_2072,N_1937);
nand U2355 (N_2355,N_1909,N_1810);
and U2356 (N_2356,N_1544,N_2208);
or U2357 (N_2357,N_1782,N_2231);
xor U2358 (N_2358,N_1931,N_1940);
and U2359 (N_2359,N_2006,N_1540);
or U2360 (N_2360,N_2215,N_2168);
xnor U2361 (N_2361,N_1761,N_2162);
or U2362 (N_2362,N_1942,N_2185);
nor U2363 (N_2363,N_2141,N_1809);
and U2364 (N_2364,N_1673,N_1823);
nor U2365 (N_2365,N_1510,N_2108);
xnor U2366 (N_2366,N_1812,N_2065);
nand U2367 (N_2367,N_2202,N_2096);
nor U2368 (N_2368,N_2004,N_2057);
nand U2369 (N_2369,N_1685,N_1827);
nor U2370 (N_2370,N_1642,N_2154);
xnor U2371 (N_2371,N_2247,N_2052);
and U2372 (N_2372,N_2098,N_2022);
nor U2373 (N_2373,N_1569,N_2246);
or U2374 (N_2374,N_2079,N_2020);
xnor U2375 (N_2375,N_1506,N_1952);
or U2376 (N_2376,N_2071,N_2034);
xnor U2377 (N_2377,N_1657,N_1764);
xnor U2378 (N_2378,N_1613,N_2145);
nor U2379 (N_2379,N_1895,N_1752);
nand U2380 (N_2380,N_1944,N_1878);
nor U2381 (N_2381,N_1542,N_1818);
xnor U2382 (N_2382,N_1532,N_2196);
nand U2383 (N_2383,N_2187,N_1765);
xnor U2384 (N_2384,N_1683,N_2160);
and U2385 (N_2385,N_1817,N_1678);
or U2386 (N_2386,N_1840,N_1596);
nor U2387 (N_2387,N_1658,N_1679);
xnor U2388 (N_2388,N_1518,N_2158);
or U2389 (N_2389,N_2082,N_1523);
nor U2390 (N_2390,N_1838,N_1591);
nand U2391 (N_2391,N_2212,N_1730);
and U2392 (N_2392,N_1624,N_1821);
nand U2393 (N_2393,N_1950,N_1887);
nor U2394 (N_2394,N_1712,N_1767);
and U2395 (N_2395,N_1807,N_1790);
nand U2396 (N_2396,N_2179,N_2153);
nor U2397 (N_2397,N_1713,N_1770);
nor U2398 (N_2398,N_2159,N_2092);
and U2399 (N_2399,N_2244,N_1667);
xnor U2400 (N_2400,N_1684,N_2241);
xnor U2401 (N_2401,N_1606,N_1803);
xnor U2402 (N_2402,N_1579,N_1545);
xnor U2403 (N_2403,N_2042,N_1505);
and U2404 (N_2404,N_1632,N_1917);
xor U2405 (N_2405,N_1595,N_1751);
nand U2406 (N_2406,N_1693,N_1570);
xnor U2407 (N_2407,N_1556,N_1834);
xnor U2408 (N_2408,N_1833,N_1990);
xor U2409 (N_2409,N_1725,N_1514);
nand U2410 (N_2410,N_1608,N_2147);
or U2411 (N_2411,N_1911,N_2227);
or U2412 (N_2412,N_1720,N_1863);
and U2413 (N_2413,N_1939,N_1574);
and U2414 (N_2414,N_1962,N_1677);
xnor U2415 (N_2415,N_2109,N_1808);
and U2416 (N_2416,N_1581,N_1555);
and U2417 (N_2417,N_2024,N_2234);
nor U2418 (N_2418,N_1829,N_1567);
nor U2419 (N_2419,N_1648,N_1835);
or U2420 (N_2420,N_2067,N_1749);
xnor U2421 (N_2421,N_1890,N_1843);
xnor U2422 (N_2422,N_2053,N_2123);
nand U2423 (N_2423,N_1970,N_2019);
and U2424 (N_2424,N_1891,N_1881);
and U2425 (N_2425,N_1709,N_1633);
xnor U2426 (N_2426,N_2070,N_1836);
and U2427 (N_2427,N_1629,N_2100);
nor U2428 (N_2428,N_1610,N_2104);
xnor U2429 (N_2429,N_2169,N_1898);
xor U2430 (N_2430,N_2189,N_1551);
nor U2431 (N_2431,N_1584,N_2112);
nor U2432 (N_2432,N_2086,N_1857);
and U2433 (N_2433,N_1701,N_2076);
and U2434 (N_2434,N_1860,N_2111);
nor U2435 (N_2435,N_2223,N_1548);
xnor U2436 (N_2436,N_1824,N_1865);
nor U2437 (N_2437,N_1876,N_2181);
or U2438 (N_2438,N_1813,N_1786);
and U2439 (N_2439,N_2007,N_2002);
or U2440 (N_2440,N_2177,N_2164);
nor U2441 (N_2441,N_1814,N_2194);
nor U2442 (N_2442,N_1601,N_1738);
nor U2443 (N_2443,N_1987,N_1915);
xnor U2444 (N_2444,N_1902,N_1630);
xor U2445 (N_2445,N_2217,N_1565);
xnor U2446 (N_2446,N_1747,N_2044);
nand U2447 (N_2447,N_1910,N_2232);
or U2448 (N_2448,N_2047,N_1757);
or U2449 (N_2449,N_2033,N_2178);
xor U2450 (N_2450,N_1529,N_2046);
nand U2451 (N_2451,N_1674,N_2116);
and U2452 (N_2452,N_1519,N_1622);
nor U2453 (N_2453,N_1995,N_2041);
or U2454 (N_2454,N_1769,N_1580);
or U2455 (N_2455,N_2117,N_1588);
nand U2456 (N_2456,N_1741,N_1992);
and U2457 (N_2457,N_1792,N_2005);
or U2458 (N_2458,N_2135,N_1954);
and U2459 (N_2459,N_1718,N_1617);
or U2460 (N_2460,N_1811,N_2206);
xnor U2461 (N_2461,N_2193,N_1528);
nor U2462 (N_2462,N_2069,N_1982);
or U2463 (N_2463,N_1716,N_2190);
or U2464 (N_2464,N_1822,N_1750);
nand U2465 (N_2465,N_1979,N_2045);
xnor U2466 (N_2466,N_1566,N_1816);
nand U2467 (N_2467,N_1754,N_2210);
or U2468 (N_2468,N_1896,N_1947);
xor U2469 (N_2469,N_1819,N_2235);
xor U2470 (N_2470,N_1627,N_1930);
and U2471 (N_2471,N_1748,N_1894);
xnor U2472 (N_2472,N_1924,N_1616);
nand U2473 (N_2473,N_2238,N_1913);
or U2474 (N_2474,N_2014,N_2151);
and U2475 (N_2475,N_1957,N_2134);
nor U2476 (N_2476,N_2083,N_1644);
xnor U2477 (N_2477,N_1665,N_2095);
nand U2478 (N_2478,N_1612,N_2127);
or U2479 (N_2479,N_1719,N_2087);
or U2480 (N_2480,N_1694,N_2248);
nor U2481 (N_2481,N_1953,N_1976);
xnor U2482 (N_2482,N_1703,N_1561);
xnor U2483 (N_2483,N_1904,N_1609);
or U2484 (N_2484,N_1806,N_1755);
nor U2485 (N_2485,N_2073,N_1966);
xor U2486 (N_2486,N_1522,N_1660);
nor U2487 (N_2487,N_2102,N_1602);
or U2488 (N_2488,N_1943,N_1611);
and U2489 (N_2489,N_1577,N_1977);
nand U2490 (N_2490,N_1625,N_1710);
nand U2491 (N_2491,N_1547,N_1973);
and U2492 (N_2492,N_1971,N_1796);
and U2493 (N_2493,N_1640,N_2236);
nor U2494 (N_2494,N_1534,N_2090);
nor U2495 (N_2495,N_1989,N_1960);
and U2496 (N_2496,N_1906,N_1980);
nor U2497 (N_2497,N_2037,N_1614);
nand U2498 (N_2498,N_1869,N_1916);
nor U2499 (N_2499,N_2000,N_1691);
or U2500 (N_2500,N_1704,N_2035);
nor U2501 (N_2501,N_1714,N_1858);
nand U2502 (N_2502,N_2161,N_1668);
and U2503 (N_2503,N_1639,N_2074);
xor U2504 (N_2504,N_2009,N_2139);
nor U2505 (N_2505,N_1746,N_1900);
nor U2506 (N_2506,N_1671,N_1897);
xor U2507 (N_2507,N_1721,N_1837);
or U2508 (N_2508,N_2186,N_1500);
nor U2509 (N_2509,N_1783,N_2061);
nor U2510 (N_2510,N_1985,N_2106);
or U2511 (N_2511,N_1958,N_2017);
nor U2512 (N_2512,N_2230,N_1628);
nand U2513 (N_2513,N_1531,N_1991);
nor U2514 (N_2514,N_2008,N_2150);
and U2515 (N_2515,N_1880,N_1619);
or U2516 (N_2516,N_1700,N_2043);
nand U2517 (N_2517,N_1553,N_2203);
or U2518 (N_2518,N_1501,N_1536);
or U2519 (N_2519,N_2064,N_1926);
nor U2520 (N_2520,N_2081,N_1743);
nand U2521 (N_2521,N_1846,N_1549);
nor U2522 (N_2522,N_1789,N_1615);
xor U2523 (N_2523,N_2050,N_2048);
nand U2524 (N_2524,N_1732,N_2099);
xnor U2525 (N_2525,N_2126,N_1515);
and U2526 (N_2526,N_2028,N_2172);
xor U2527 (N_2527,N_1578,N_1650);
nor U2528 (N_2528,N_1946,N_2131);
or U2529 (N_2529,N_1729,N_1696);
and U2530 (N_2530,N_2128,N_1874);
or U2531 (N_2531,N_1525,N_1851);
nand U2532 (N_2532,N_2199,N_1879);
and U2533 (N_2533,N_1885,N_1583);
nor U2534 (N_2534,N_1768,N_1699);
and U2535 (N_2535,N_1621,N_2105);
and U2536 (N_2536,N_2058,N_2132);
nand U2537 (N_2537,N_2101,N_2176);
xnor U2538 (N_2538,N_2204,N_1552);
and U2539 (N_2539,N_1599,N_2030);
nand U2540 (N_2540,N_1598,N_2107);
nor U2541 (N_2541,N_1839,N_1502);
nor U2542 (N_2542,N_1820,N_1504);
or U2543 (N_2543,N_1638,N_1849);
or U2544 (N_2544,N_1600,N_1733);
nor U2545 (N_2545,N_1842,N_2001);
nor U2546 (N_2546,N_1737,N_1670);
xor U2547 (N_2547,N_2010,N_1563);
xor U2548 (N_2548,N_1938,N_1539);
xnor U2549 (N_2549,N_1723,N_1983);
and U2550 (N_2550,N_2011,N_1859);
and U2551 (N_2551,N_1892,N_1965);
or U2552 (N_2552,N_1568,N_1663);
or U2553 (N_2553,N_1550,N_1969);
and U2554 (N_2554,N_2093,N_1572);
xor U2555 (N_2555,N_1740,N_1641);
and U2556 (N_2556,N_1855,N_1744);
xor U2557 (N_2557,N_2023,N_2197);
and U2558 (N_2558,N_1825,N_1886);
or U2559 (N_2559,N_2149,N_2089);
xnor U2560 (N_2560,N_1795,N_1756);
and U2561 (N_2561,N_2220,N_1686);
xor U2562 (N_2562,N_1826,N_1888);
nor U2563 (N_2563,N_1722,N_1676);
xor U2564 (N_2564,N_1652,N_1848);
and U2565 (N_2565,N_1554,N_1618);
nor U2566 (N_2566,N_1919,N_1508);
xor U2567 (N_2567,N_2138,N_1776);
and U2568 (N_2568,N_1785,N_1726);
xnor U2569 (N_2569,N_2133,N_1681);
and U2570 (N_2570,N_1778,N_1984);
and U2571 (N_2571,N_1643,N_2242);
and U2572 (N_2572,N_2182,N_1773);
and U2573 (N_2573,N_1959,N_1912);
nand U2574 (N_2574,N_1932,N_1968);
xnor U2575 (N_2575,N_2146,N_1779);
nor U2576 (N_2576,N_1760,N_1546);
xor U2577 (N_2577,N_2184,N_2201);
nand U2578 (N_2578,N_1651,N_1955);
and U2579 (N_2579,N_1558,N_1655);
or U2580 (N_2580,N_1914,N_1521);
and U2581 (N_2581,N_2174,N_1538);
nor U2582 (N_2582,N_2118,N_1697);
or U2583 (N_2583,N_1775,N_1893);
nand U2584 (N_2584,N_1530,N_1967);
nand U2585 (N_2585,N_2192,N_1918);
nor U2586 (N_2586,N_1524,N_2229);
and U2587 (N_2587,N_2142,N_2239);
xnor U2588 (N_2588,N_2191,N_2188);
and U2589 (N_2589,N_1832,N_1735);
and U2590 (N_2590,N_2195,N_1689);
or U2591 (N_2591,N_1871,N_2016);
and U2592 (N_2592,N_1562,N_2075);
and U2593 (N_2593,N_2021,N_2120);
xnor U2594 (N_2594,N_1804,N_1873);
nor U2595 (N_2595,N_1929,N_1507);
nand U2596 (N_2596,N_2226,N_1781);
nor U2597 (N_2597,N_2243,N_2056);
xor U2598 (N_2598,N_1903,N_2088);
and U2599 (N_2599,N_2031,N_1974);
and U2600 (N_2600,N_1988,N_1724);
xnor U2601 (N_2601,N_2211,N_1620);
xor U2602 (N_2602,N_1759,N_1582);
xnor U2603 (N_2603,N_2163,N_1708);
nor U2604 (N_2604,N_1661,N_2148);
nor U2605 (N_2605,N_1941,N_1687);
nand U2606 (N_2606,N_1739,N_1734);
or U2607 (N_2607,N_1664,N_2110);
nor U2608 (N_2608,N_2237,N_1981);
nand U2609 (N_2609,N_2097,N_2180);
xnor U2610 (N_2610,N_1949,N_2080);
or U2611 (N_2611,N_1828,N_2143);
nand U2612 (N_2612,N_1512,N_1928);
xnor U2613 (N_2613,N_1537,N_1590);
or U2614 (N_2614,N_2039,N_1875);
nand U2615 (N_2615,N_1604,N_1864);
xor U2616 (N_2616,N_1715,N_1978);
or U2617 (N_2617,N_1635,N_2103);
xnor U2618 (N_2618,N_2167,N_2060);
and U2619 (N_2619,N_1541,N_1647);
or U2620 (N_2620,N_1711,N_1797);
or U2621 (N_2621,N_2233,N_1901);
xnor U2622 (N_2622,N_1560,N_1802);
and U2623 (N_2623,N_1905,N_2245);
or U2624 (N_2624,N_2221,N_1605);
or U2625 (N_2625,N_1614,N_2159);
xor U2626 (N_2626,N_1608,N_1906);
nor U2627 (N_2627,N_1997,N_1841);
or U2628 (N_2628,N_1923,N_1877);
nand U2629 (N_2629,N_1560,N_1862);
xnor U2630 (N_2630,N_1735,N_2000);
and U2631 (N_2631,N_2185,N_2053);
and U2632 (N_2632,N_2245,N_1782);
nand U2633 (N_2633,N_2136,N_1520);
nor U2634 (N_2634,N_1861,N_1834);
nand U2635 (N_2635,N_1643,N_2128);
and U2636 (N_2636,N_1964,N_1532);
nor U2637 (N_2637,N_1814,N_2226);
nor U2638 (N_2638,N_2191,N_1625);
nand U2639 (N_2639,N_1612,N_1500);
nand U2640 (N_2640,N_2004,N_1670);
xor U2641 (N_2641,N_1891,N_1788);
xor U2642 (N_2642,N_1766,N_1542);
and U2643 (N_2643,N_1508,N_1850);
nor U2644 (N_2644,N_2017,N_1816);
nand U2645 (N_2645,N_1598,N_1522);
xor U2646 (N_2646,N_1914,N_1724);
xnor U2647 (N_2647,N_2031,N_1878);
and U2648 (N_2648,N_1559,N_2100);
and U2649 (N_2649,N_2018,N_1606);
nand U2650 (N_2650,N_2151,N_2216);
nand U2651 (N_2651,N_2038,N_2022);
and U2652 (N_2652,N_1746,N_1579);
nor U2653 (N_2653,N_1945,N_2197);
nor U2654 (N_2654,N_2180,N_1538);
nand U2655 (N_2655,N_1628,N_1962);
or U2656 (N_2656,N_1533,N_2069);
and U2657 (N_2657,N_2074,N_2000);
nor U2658 (N_2658,N_1840,N_1898);
xor U2659 (N_2659,N_1550,N_2138);
nor U2660 (N_2660,N_1869,N_1788);
and U2661 (N_2661,N_1839,N_1505);
nand U2662 (N_2662,N_2102,N_1810);
and U2663 (N_2663,N_2180,N_1914);
or U2664 (N_2664,N_1753,N_1682);
and U2665 (N_2665,N_2204,N_1764);
nand U2666 (N_2666,N_1873,N_2194);
or U2667 (N_2667,N_2219,N_2222);
or U2668 (N_2668,N_2018,N_1511);
nor U2669 (N_2669,N_1900,N_2034);
nand U2670 (N_2670,N_2168,N_1609);
nor U2671 (N_2671,N_1614,N_2018);
nor U2672 (N_2672,N_1503,N_1847);
nor U2673 (N_2673,N_1563,N_2075);
nand U2674 (N_2674,N_1742,N_1660);
nor U2675 (N_2675,N_1567,N_1766);
nand U2676 (N_2676,N_1629,N_1899);
xnor U2677 (N_2677,N_1799,N_1723);
xnor U2678 (N_2678,N_1612,N_1712);
nor U2679 (N_2679,N_1672,N_1644);
and U2680 (N_2680,N_1709,N_1798);
and U2681 (N_2681,N_1894,N_2238);
nand U2682 (N_2682,N_1713,N_2060);
or U2683 (N_2683,N_1722,N_2114);
xnor U2684 (N_2684,N_1714,N_2167);
nand U2685 (N_2685,N_1895,N_2006);
and U2686 (N_2686,N_2134,N_2219);
xnor U2687 (N_2687,N_1980,N_2182);
nor U2688 (N_2688,N_1806,N_2227);
nor U2689 (N_2689,N_1695,N_1508);
or U2690 (N_2690,N_1778,N_2072);
nand U2691 (N_2691,N_2088,N_1911);
and U2692 (N_2692,N_1544,N_2156);
nor U2693 (N_2693,N_1824,N_2162);
nor U2694 (N_2694,N_1530,N_1618);
nor U2695 (N_2695,N_1711,N_1740);
xnor U2696 (N_2696,N_1515,N_2147);
nand U2697 (N_2697,N_1697,N_2200);
or U2698 (N_2698,N_1564,N_1751);
or U2699 (N_2699,N_2074,N_2029);
nand U2700 (N_2700,N_1510,N_2009);
nor U2701 (N_2701,N_1539,N_1545);
nand U2702 (N_2702,N_2202,N_2209);
xor U2703 (N_2703,N_1663,N_1739);
or U2704 (N_2704,N_1639,N_1583);
or U2705 (N_2705,N_1665,N_1962);
and U2706 (N_2706,N_1643,N_1869);
nor U2707 (N_2707,N_2192,N_2081);
nand U2708 (N_2708,N_2064,N_1883);
xor U2709 (N_2709,N_1641,N_2066);
or U2710 (N_2710,N_1763,N_1966);
nor U2711 (N_2711,N_1854,N_1531);
nand U2712 (N_2712,N_1836,N_2024);
or U2713 (N_2713,N_1681,N_2003);
nand U2714 (N_2714,N_1707,N_1980);
nand U2715 (N_2715,N_2023,N_2052);
and U2716 (N_2716,N_1670,N_2081);
xor U2717 (N_2717,N_2077,N_1650);
nand U2718 (N_2718,N_2068,N_2040);
and U2719 (N_2719,N_1667,N_2078);
or U2720 (N_2720,N_2192,N_2133);
and U2721 (N_2721,N_2073,N_1908);
or U2722 (N_2722,N_1911,N_1734);
nor U2723 (N_2723,N_1877,N_1555);
nor U2724 (N_2724,N_1882,N_1950);
and U2725 (N_2725,N_1974,N_2025);
or U2726 (N_2726,N_1659,N_1536);
or U2727 (N_2727,N_1595,N_2103);
nand U2728 (N_2728,N_1753,N_1623);
nand U2729 (N_2729,N_1654,N_1977);
and U2730 (N_2730,N_2091,N_1513);
xnor U2731 (N_2731,N_2133,N_1500);
nor U2732 (N_2732,N_1616,N_1575);
nor U2733 (N_2733,N_2159,N_1956);
or U2734 (N_2734,N_2011,N_1811);
and U2735 (N_2735,N_1707,N_1705);
nand U2736 (N_2736,N_1613,N_2043);
xnor U2737 (N_2737,N_2232,N_1524);
nor U2738 (N_2738,N_2117,N_1860);
or U2739 (N_2739,N_1870,N_1842);
nor U2740 (N_2740,N_1810,N_1903);
nand U2741 (N_2741,N_1827,N_1906);
or U2742 (N_2742,N_1705,N_1584);
and U2743 (N_2743,N_1512,N_1726);
or U2744 (N_2744,N_1942,N_1782);
and U2745 (N_2745,N_1903,N_1595);
xor U2746 (N_2746,N_1787,N_1982);
nand U2747 (N_2747,N_2242,N_1543);
and U2748 (N_2748,N_1986,N_1918);
and U2749 (N_2749,N_1643,N_1576);
nand U2750 (N_2750,N_1972,N_2140);
xor U2751 (N_2751,N_2061,N_2241);
nand U2752 (N_2752,N_1625,N_1778);
nand U2753 (N_2753,N_2142,N_1832);
and U2754 (N_2754,N_1964,N_1765);
xnor U2755 (N_2755,N_1876,N_1968);
and U2756 (N_2756,N_1699,N_2090);
nor U2757 (N_2757,N_2166,N_1552);
or U2758 (N_2758,N_1908,N_1622);
and U2759 (N_2759,N_2165,N_1567);
xor U2760 (N_2760,N_2103,N_1946);
xnor U2761 (N_2761,N_1690,N_1575);
nand U2762 (N_2762,N_2016,N_1903);
or U2763 (N_2763,N_2051,N_1679);
nor U2764 (N_2764,N_2112,N_2101);
and U2765 (N_2765,N_2249,N_1738);
xnor U2766 (N_2766,N_2022,N_2205);
xor U2767 (N_2767,N_1517,N_2164);
and U2768 (N_2768,N_1966,N_1706);
nor U2769 (N_2769,N_2093,N_2231);
or U2770 (N_2770,N_1546,N_1758);
and U2771 (N_2771,N_1799,N_1891);
xor U2772 (N_2772,N_1616,N_1701);
xor U2773 (N_2773,N_1510,N_1763);
xor U2774 (N_2774,N_2143,N_2084);
and U2775 (N_2775,N_1594,N_1776);
xnor U2776 (N_2776,N_1520,N_2212);
xnor U2777 (N_2777,N_2227,N_2186);
xnor U2778 (N_2778,N_2016,N_2036);
nand U2779 (N_2779,N_2025,N_1621);
nor U2780 (N_2780,N_1889,N_2037);
and U2781 (N_2781,N_1936,N_1716);
xor U2782 (N_2782,N_1579,N_1611);
and U2783 (N_2783,N_1512,N_2106);
nand U2784 (N_2784,N_2217,N_1856);
nor U2785 (N_2785,N_2241,N_2096);
xor U2786 (N_2786,N_1625,N_2246);
and U2787 (N_2787,N_1959,N_1878);
nor U2788 (N_2788,N_1557,N_1743);
or U2789 (N_2789,N_1677,N_1994);
nor U2790 (N_2790,N_1869,N_2166);
and U2791 (N_2791,N_1720,N_2128);
nor U2792 (N_2792,N_2203,N_2159);
or U2793 (N_2793,N_1805,N_2163);
xor U2794 (N_2794,N_2100,N_2012);
nand U2795 (N_2795,N_2118,N_1848);
and U2796 (N_2796,N_1502,N_2002);
and U2797 (N_2797,N_1744,N_1899);
xor U2798 (N_2798,N_2087,N_1755);
or U2799 (N_2799,N_1657,N_2185);
nand U2800 (N_2800,N_1928,N_1827);
nor U2801 (N_2801,N_1900,N_1769);
nor U2802 (N_2802,N_1616,N_2056);
xnor U2803 (N_2803,N_1632,N_1665);
nor U2804 (N_2804,N_1828,N_2125);
nor U2805 (N_2805,N_1652,N_1945);
nor U2806 (N_2806,N_1574,N_2010);
or U2807 (N_2807,N_1977,N_2164);
or U2808 (N_2808,N_1586,N_1990);
xor U2809 (N_2809,N_1686,N_1790);
nand U2810 (N_2810,N_2090,N_2179);
nand U2811 (N_2811,N_1563,N_1736);
or U2812 (N_2812,N_1823,N_1883);
and U2813 (N_2813,N_1855,N_2148);
nor U2814 (N_2814,N_1786,N_2166);
nor U2815 (N_2815,N_2103,N_2133);
and U2816 (N_2816,N_1765,N_1934);
nand U2817 (N_2817,N_1845,N_1786);
nor U2818 (N_2818,N_2093,N_1927);
or U2819 (N_2819,N_1575,N_2202);
or U2820 (N_2820,N_1530,N_2201);
nand U2821 (N_2821,N_1513,N_1632);
nor U2822 (N_2822,N_1980,N_1709);
nor U2823 (N_2823,N_1787,N_1720);
or U2824 (N_2824,N_1715,N_1617);
or U2825 (N_2825,N_1820,N_2113);
xnor U2826 (N_2826,N_1847,N_1537);
nor U2827 (N_2827,N_2053,N_2217);
nand U2828 (N_2828,N_1588,N_2188);
or U2829 (N_2829,N_1778,N_1533);
xnor U2830 (N_2830,N_1857,N_1968);
xnor U2831 (N_2831,N_1860,N_1863);
nor U2832 (N_2832,N_2249,N_1989);
or U2833 (N_2833,N_2089,N_2002);
nand U2834 (N_2834,N_1966,N_2018);
and U2835 (N_2835,N_1699,N_1987);
or U2836 (N_2836,N_1904,N_2015);
nand U2837 (N_2837,N_1667,N_1841);
nor U2838 (N_2838,N_1555,N_2217);
or U2839 (N_2839,N_1666,N_1946);
nand U2840 (N_2840,N_1994,N_1763);
and U2841 (N_2841,N_1919,N_1710);
xor U2842 (N_2842,N_1750,N_1707);
or U2843 (N_2843,N_1919,N_1595);
nand U2844 (N_2844,N_1514,N_2229);
xnor U2845 (N_2845,N_1830,N_1740);
or U2846 (N_2846,N_1751,N_1697);
and U2847 (N_2847,N_1662,N_2059);
and U2848 (N_2848,N_1595,N_1819);
nor U2849 (N_2849,N_1933,N_2051);
nand U2850 (N_2850,N_1932,N_1839);
or U2851 (N_2851,N_1869,N_1690);
and U2852 (N_2852,N_1982,N_1532);
nor U2853 (N_2853,N_1741,N_1967);
or U2854 (N_2854,N_1705,N_1754);
nand U2855 (N_2855,N_2015,N_1967);
or U2856 (N_2856,N_1696,N_1580);
and U2857 (N_2857,N_2196,N_2057);
or U2858 (N_2858,N_2159,N_1556);
xnor U2859 (N_2859,N_1577,N_2171);
and U2860 (N_2860,N_2175,N_1572);
and U2861 (N_2861,N_1892,N_1851);
nor U2862 (N_2862,N_1895,N_1567);
nor U2863 (N_2863,N_1957,N_1781);
nand U2864 (N_2864,N_1802,N_2248);
nand U2865 (N_2865,N_1961,N_2083);
nor U2866 (N_2866,N_1506,N_2032);
nand U2867 (N_2867,N_1592,N_2203);
and U2868 (N_2868,N_1800,N_1989);
and U2869 (N_2869,N_2001,N_1863);
and U2870 (N_2870,N_1673,N_2045);
nor U2871 (N_2871,N_2067,N_2069);
and U2872 (N_2872,N_1589,N_2072);
xor U2873 (N_2873,N_1525,N_1881);
or U2874 (N_2874,N_1783,N_2116);
nor U2875 (N_2875,N_2148,N_1574);
and U2876 (N_2876,N_2227,N_1759);
and U2877 (N_2877,N_1954,N_1826);
and U2878 (N_2878,N_1979,N_1634);
nand U2879 (N_2879,N_1563,N_1756);
xnor U2880 (N_2880,N_1887,N_1589);
or U2881 (N_2881,N_1971,N_2120);
nand U2882 (N_2882,N_1529,N_1735);
and U2883 (N_2883,N_1801,N_2222);
and U2884 (N_2884,N_2234,N_2189);
or U2885 (N_2885,N_2129,N_2210);
or U2886 (N_2886,N_1664,N_1773);
nor U2887 (N_2887,N_1817,N_2217);
xor U2888 (N_2888,N_2082,N_1638);
nor U2889 (N_2889,N_1615,N_1602);
or U2890 (N_2890,N_2092,N_2247);
or U2891 (N_2891,N_1811,N_1921);
xnor U2892 (N_2892,N_1865,N_1527);
or U2893 (N_2893,N_2226,N_1631);
xnor U2894 (N_2894,N_1613,N_2094);
nor U2895 (N_2895,N_1507,N_1965);
nor U2896 (N_2896,N_2239,N_1950);
nand U2897 (N_2897,N_2020,N_2200);
nor U2898 (N_2898,N_1973,N_2079);
xnor U2899 (N_2899,N_1607,N_2119);
and U2900 (N_2900,N_2089,N_1757);
and U2901 (N_2901,N_1742,N_1526);
nor U2902 (N_2902,N_1506,N_2237);
nand U2903 (N_2903,N_1839,N_1930);
xor U2904 (N_2904,N_1760,N_1836);
xnor U2905 (N_2905,N_1808,N_1977);
or U2906 (N_2906,N_1572,N_1660);
xnor U2907 (N_2907,N_2232,N_2140);
or U2908 (N_2908,N_2112,N_2194);
nor U2909 (N_2909,N_1981,N_1838);
and U2910 (N_2910,N_2184,N_2055);
nand U2911 (N_2911,N_1938,N_1826);
or U2912 (N_2912,N_2124,N_2217);
xnor U2913 (N_2913,N_1741,N_1917);
nand U2914 (N_2914,N_2078,N_1658);
nand U2915 (N_2915,N_1565,N_1697);
nor U2916 (N_2916,N_2241,N_2113);
or U2917 (N_2917,N_2094,N_1661);
or U2918 (N_2918,N_1737,N_1769);
or U2919 (N_2919,N_2025,N_2245);
nand U2920 (N_2920,N_1927,N_1579);
xor U2921 (N_2921,N_1701,N_1822);
or U2922 (N_2922,N_1698,N_2190);
or U2923 (N_2923,N_1504,N_2017);
nor U2924 (N_2924,N_2065,N_1569);
xnor U2925 (N_2925,N_1666,N_1998);
nand U2926 (N_2926,N_2107,N_1845);
xnor U2927 (N_2927,N_1670,N_2217);
nor U2928 (N_2928,N_1673,N_1615);
xor U2929 (N_2929,N_1948,N_1501);
and U2930 (N_2930,N_1604,N_1772);
xor U2931 (N_2931,N_1730,N_2227);
and U2932 (N_2932,N_1654,N_1655);
nor U2933 (N_2933,N_1649,N_2195);
nor U2934 (N_2934,N_1761,N_1660);
or U2935 (N_2935,N_1738,N_1787);
nor U2936 (N_2936,N_1644,N_1788);
and U2937 (N_2937,N_1993,N_1704);
or U2938 (N_2938,N_1513,N_2101);
or U2939 (N_2939,N_1957,N_1780);
nor U2940 (N_2940,N_1553,N_1909);
nor U2941 (N_2941,N_1919,N_1930);
nand U2942 (N_2942,N_1824,N_1790);
and U2943 (N_2943,N_1746,N_1895);
xnor U2944 (N_2944,N_1641,N_2050);
and U2945 (N_2945,N_1673,N_1618);
or U2946 (N_2946,N_1892,N_1665);
nor U2947 (N_2947,N_1799,N_2229);
nor U2948 (N_2948,N_1514,N_1950);
or U2949 (N_2949,N_1827,N_1718);
or U2950 (N_2950,N_1640,N_1767);
xnor U2951 (N_2951,N_2224,N_2112);
and U2952 (N_2952,N_1798,N_1976);
nand U2953 (N_2953,N_1524,N_1934);
xnor U2954 (N_2954,N_2029,N_1642);
nand U2955 (N_2955,N_2136,N_1528);
or U2956 (N_2956,N_1727,N_2238);
nor U2957 (N_2957,N_1835,N_2003);
nand U2958 (N_2958,N_2097,N_1845);
nand U2959 (N_2959,N_1517,N_2140);
xnor U2960 (N_2960,N_1814,N_2174);
xnor U2961 (N_2961,N_1864,N_2106);
xnor U2962 (N_2962,N_1691,N_1933);
nor U2963 (N_2963,N_1918,N_1991);
nand U2964 (N_2964,N_2085,N_1654);
nand U2965 (N_2965,N_1620,N_2163);
nor U2966 (N_2966,N_1988,N_1509);
and U2967 (N_2967,N_1828,N_1903);
or U2968 (N_2968,N_2237,N_1521);
xor U2969 (N_2969,N_1988,N_2149);
or U2970 (N_2970,N_1838,N_1574);
nor U2971 (N_2971,N_1706,N_1584);
nor U2972 (N_2972,N_1798,N_1956);
xnor U2973 (N_2973,N_2116,N_1851);
nor U2974 (N_2974,N_1668,N_1831);
nand U2975 (N_2975,N_2103,N_2171);
nor U2976 (N_2976,N_2224,N_2171);
or U2977 (N_2977,N_1916,N_1849);
and U2978 (N_2978,N_1841,N_2109);
and U2979 (N_2979,N_2094,N_2114);
nand U2980 (N_2980,N_1739,N_1591);
xnor U2981 (N_2981,N_2106,N_2136);
xnor U2982 (N_2982,N_1635,N_2172);
xor U2983 (N_2983,N_1760,N_1824);
nor U2984 (N_2984,N_2098,N_1806);
nor U2985 (N_2985,N_1762,N_1994);
or U2986 (N_2986,N_1993,N_1825);
nor U2987 (N_2987,N_1614,N_1977);
and U2988 (N_2988,N_1805,N_1747);
or U2989 (N_2989,N_2187,N_1981);
and U2990 (N_2990,N_1636,N_1590);
nand U2991 (N_2991,N_2242,N_1652);
and U2992 (N_2992,N_1887,N_2051);
and U2993 (N_2993,N_1674,N_2231);
nand U2994 (N_2994,N_1945,N_1800);
nand U2995 (N_2995,N_2167,N_2099);
or U2996 (N_2996,N_1617,N_2077);
nor U2997 (N_2997,N_2164,N_1533);
or U2998 (N_2998,N_1845,N_2086);
xor U2999 (N_2999,N_2161,N_1757);
nand UO_0 (O_0,N_2598,N_2888);
or UO_1 (O_1,N_2409,N_2910);
nor UO_2 (O_2,N_2963,N_2950);
and UO_3 (O_3,N_2810,N_2413);
and UO_4 (O_4,N_2825,N_2412);
nand UO_5 (O_5,N_2821,N_2383);
nor UO_6 (O_6,N_2776,N_2541);
or UO_7 (O_7,N_2555,N_2742);
xor UO_8 (O_8,N_2414,N_2483);
nor UO_9 (O_9,N_2933,N_2619);
nor UO_10 (O_10,N_2283,N_2687);
and UO_11 (O_11,N_2417,N_2840);
or UO_12 (O_12,N_2572,N_2790);
and UO_13 (O_13,N_2864,N_2425);
nor UO_14 (O_14,N_2672,N_2689);
nor UO_15 (O_15,N_2537,N_2889);
and UO_16 (O_16,N_2779,N_2335);
nor UO_17 (O_17,N_2739,N_2977);
nor UO_18 (O_18,N_2624,N_2818);
and UO_19 (O_19,N_2700,N_2749);
or UO_20 (O_20,N_2652,N_2843);
nor UO_21 (O_21,N_2860,N_2964);
or UO_22 (O_22,N_2431,N_2463);
xor UO_23 (O_23,N_2813,N_2307);
nor UO_24 (O_24,N_2556,N_2433);
or UO_25 (O_25,N_2395,N_2728);
nand UO_26 (O_26,N_2927,N_2873);
and UO_27 (O_27,N_2390,N_2774);
or UO_28 (O_28,N_2903,N_2449);
xor UO_29 (O_29,N_2268,N_2877);
and UO_30 (O_30,N_2688,N_2945);
xor UO_31 (O_31,N_2710,N_2550);
nor UO_32 (O_32,N_2302,N_2525);
nor UO_33 (O_33,N_2384,N_2783);
nor UO_34 (O_34,N_2536,N_2967);
nand UO_35 (O_35,N_2394,N_2533);
or UO_36 (O_36,N_2979,N_2276);
nand UO_37 (O_37,N_2909,N_2714);
nand UO_38 (O_38,N_2605,N_2988);
or UO_39 (O_39,N_2786,N_2995);
nor UO_40 (O_40,N_2701,N_2321);
nor UO_41 (O_41,N_2703,N_2416);
and UO_42 (O_42,N_2679,N_2982);
or UO_43 (O_43,N_2581,N_2668);
xor UO_44 (O_44,N_2435,N_2316);
xor UO_45 (O_45,N_2820,N_2626);
and UO_46 (O_46,N_2750,N_2271);
and UO_47 (O_47,N_2415,N_2633);
nand UO_48 (O_48,N_2830,N_2275);
and UO_49 (O_49,N_2486,N_2570);
nand UO_50 (O_50,N_2315,N_2844);
nand UO_51 (O_51,N_2938,N_2369);
xnor UO_52 (O_52,N_2498,N_2490);
nand UO_53 (O_53,N_2992,N_2812);
and UO_54 (O_54,N_2625,N_2420);
and UO_55 (O_55,N_2639,N_2727);
nor UO_56 (O_56,N_2292,N_2939);
nand UO_57 (O_57,N_2968,N_2929);
xnor UO_58 (O_58,N_2874,N_2788);
or UO_59 (O_59,N_2586,N_2677);
and UO_60 (O_60,N_2352,N_2721);
xnor UO_61 (O_61,N_2971,N_2870);
xor UO_62 (O_62,N_2252,N_2583);
xor UO_63 (O_63,N_2985,N_2955);
or UO_64 (O_64,N_2584,N_2530);
or UO_65 (O_65,N_2765,N_2332);
and UO_66 (O_66,N_2656,N_2862);
or UO_67 (O_67,N_2879,N_2998);
nand UO_68 (O_68,N_2607,N_2850);
and UO_69 (O_69,N_2775,N_2565);
xor UO_70 (O_70,N_2694,N_2257);
xnor UO_71 (O_71,N_2311,N_2817);
or UO_72 (O_72,N_2661,N_2443);
or UO_73 (O_73,N_2482,N_2623);
and UO_74 (O_74,N_2338,N_2915);
nand UO_75 (O_75,N_2682,N_2319);
or UO_76 (O_76,N_2685,N_2675);
or UO_77 (O_77,N_2738,N_2616);
nor UO_78 (O_78,N_2488,N_2989);
nor UO_79 (O_79,N_2699,N_2254);
xor UO_80 (O_80,N_2886,N_2378);
xor UO_81 (O_81,N_2917,N_2865);
xor UO_82 (O_82,N_2339,N_2631);
or UO_83 (O_83,N_2962,N_2331);
nand UO_84 (O_84,N_2920,N_2780);
nor UO_85 (O_85,N_2323,N_2853);
or UO_86 (O_86,N_2399,N_2717);
nand UO_87 (O_87,N_2477,N_2871);
nand UO_88 (O_88,N_2396,N_2558);
and UO_89 (O_89,N_2499,N_2940);
nand UO_90 (O_90,N_2599,N_2492);
and UO_91 (O_91,N_2330,N_2262);
or UO_92 (O_92,N_2838,N_2702);
xnor UO_93 (O_93,N_2568,N_2861);
nor UO_94 (O_94,N_2837,N_2856);
nor UO_95 (O_95,N_2997,N_2676);
nand UO_96 (O_96,N_2441,N_2648);
or UO_97 (O_97,N_2697,N_2404);
or UO_98 (O_98,N_2932,N_2961);
xnor UO_99 (O_99,N_2759,N_2552);
or UO_100 (O_100,N_2644,N_2804);
or UO_101 (O_101,N_2345,N_2503);
nor UO_102 (O_102,N_2344,N_2294);
xnor UO_103 (O_103,N_2993,N_2747);
nor UO_104 (O_104,N_2826,N_2424);
xnor UO_105 (O_105,N_2547,N_2312);
xnor UO_106 (O_106,N_2975,N_2400);
nand UO_107 (O_107,N_2410,N_2287);
xor UO_108 (O_108,N_2919,N_2502);
or UO_109 (O_109,N_2811,N_2884);
nor UO_110 (O_110,N_2348,N_2304);
xor UO_111 (O_111,N_2725,N_2373);
and UO_112 (O_112,N_2359,N_2418);
nor UO_113 (O_113,N_2513,N_2461);
nand UO_114 (O_114,N_2892,N_2693);
or UO_115 (O_115,N_2347,N_2912);
nor UO_116 (O_116,N_2479,N_2526);
nand UO_117 (O_117,N_2907,N_2680);
nand UO_118 (O_118,N_2476,N_2613);
or UO_119 (O_119,N_2669,N_2388);
xnor UO_120 (O_120,N_2432,N_2617);
nor UO_121 (O_121,N_2868,N_2391);
nand UO_122 (O_122,N_2723,N_2847);
nor UO_123 (O_123,N_2407,N_2758);
or UO_124 (O_124,N_2953,N_2458);
xor UO_125 (O_125,N_2996,N_2585);
nand UO_126 (O_126,N_2712,N_2554);
and UO_127 (O_127,N_2726,N_2539);
nor UO_128 (O_128,N_2855,N_2258);
nand UO_129 (O_129,N_2670,N_2802);
nand UO_130 (O_130,N_2914,N_2942);
nand UO_131 (O_131,N_2459,N_2447);
nand UO_132 (O_132,N_2289,N_2898);
xor UO_133 (O_133,N_2485,N_2343);
xor UO_134 (O_134,N_2990,N_2282);
nand UO_135 (O_135,N_2535,N_2506);
and UO_136 (O_136,N_2715,N_2380);
nand UO_137 (O_137,N_2666,N_2859);
nor UO_138 (O_138,N_2883,N_2571);
and UO_139 (O_139,N_2590,N_2904);
and UO_140 (O_140,N_2578,N_2722);
and UO_141 (O_141,N_2752,N_2846);
nand UO_142 (O_142,N_2867,N_2521);
xor UO_143 (O_143,N_2274,N_2356);
nor UO_144 (O_144,N_2709,N_2895);
nand UO_145 (O_145,N_2575,N_2615);
or UO_146 (O_146,N_2760,N_2908);
and UO_147 (O_147,N_2819,N_2934);
xor UO_148 (O_148,N_2328,N_2660);
nand UO_149 (O_149,N_2958,N_2926);
xnor UO_150 (O_150,N_2753,N_2828);
and UO_151 (O_151,N_2365,N_2564);
and UO_152 (O_152,N_2496,N_2845);
nor UO_153 (O_153,N_2250,N_2970);
xor UO_154 (O_154,N_2815,N_2785);
xnor UO_155 (O_155,N_2632,N_2469);
and UO_156 (O_156,N_2729,N_2944);
nor UO_157 (O_157,N_2439,N_2473);
or UO_158 (O_158,N_2403,N_2580);
xor UO_159 (O_159,N_2422,N_2382);
and UO_160 (O_160,N_2634,N_2305);
or UO_161 (O_161,N_2540,N_2466);
or UO_162 (O_162,N_2787,N_2470);
and UO_163 (O_163,N_2596,N_2520);
xnor UO_164 (O_164,N_2354,N_2673);
nand UO_165 (O_165,N_2379,N_2800);
nor UO_166 (O_166,N_2293,N_2561);
nand UO_167 (O_167,N_2451,N_2515);
nor UO_168 (O_168,N_2336,N_2579);
nand UO_169 (O_169,N_2935,N_2872);
nor UO_170 (O_170,N_2772,N_2562);
nor UO_171 (O_171,N_2754,N_2662);
and UO_172 (O_172,N_2353,N_2474);
or UO_173 (O_173,N_2740,N_2854);
xor UO_174 (O_174,N_2692,N_2973);
or UO_175 (O_175,N_2265,N_2518);
and UO_176 (O_176,N_2822,N_2716);
and UO_177 (O_177,N_2504,N_2442);
or UO_178 (O_178,N_2548,N_2999);
xnor UO_179 (O_179,N_2374,N_2902);
or UO_180 (O_180,N_2429,N_2719);
nor UO_181 (O_181,N_2767,N_2887);
nor UO_182 (O_182,N_2491,N_2733);
or UO_183 (O_183,N_2455,N_2627);
or UO_184 (O_184,N_2991,N_2894);
or UO_185 (O_185,N_2882,N_2387);
nand UO_186 (O_186,N_2875,N_2600);
nor UO_187 (O_187,N_2505,N_2322);
xor UO_188 (O_188,N_2299,N_2885);
nor UO_189 (O_189,N_2730,N_2534);
and UO_190 (O_190,N_2256,N_2794);
xor UO_191 (O_191,N_2300,N_2796);
nand UO_192 (O_192,N_2454,N_2251);
xnor UO_193 (O_193,N_2402,N_2645);
nand UO_194 (O_194,N_2711,N_2833);
and UO_195 (O_195,N_2360,N_2279);
or UO_196 (O_196,N_2770,N_2511);
or UO_197 (O_197,N_2475,N_2553);
nor UO_198 (O_198,N_2392,N_2930);
and UO_199 (O_199,N_2746,N_2649);
or UO_200 (O_200,N_2705,N_2763);
and UO_201 (O_201,N_2642,N_2465);
nor UO_202 (O_202,N_2543,N_2597);
xnor UO_203 (O_203,N_2984,N_2436);
xnor UO_204 (O_204,N_2974,N_2411);
or UO_205 (O_205,N_2456,N_2588);
xnor UO_206 (O_206,N_2582,N_2936);
and UO_207 (O_207,N_2650,N_2437);
nor UO_208 (O_208,N_2507,N_2948);
nor UO_209 (O_209,N_2266,N_2731);
nand UO_210 (O_210,N_2695,N_2638);
nand UO_211 (O_211,N_2277,N_2255);
nand UO_212 (O_212,N_2514,N_2768);
nand UO_213 (O_213,N_2683,N_2678);
nand UO_214 (O_214,N_2324,N_2516);
and UO_215 (O_215,N_2528,N_2745);
and UO_216 (O_216,N_2314,N_2773);
nand UO_217 (O_217,N_2295,N_2286);
and UO_218 (O_218,N_2921,N_2736);
nor UO_219 (O_219,N_2364,N_2659);
nor UO_220 (O_220,N_2987,N_2611);
and UO_221 (O_221,N_2529,N_2489);
and UO_222 (O_222,N_2947,N_2741);
or UO_223 (O_223,N_2781,N_2327);
xor UO_224 (O_224,N_2836,N_2735);
xor UO_225 (O_225,N_2296,N_2574);
xor UO_226 (O_226,N_2829,N_2366);
nor UO_227 (O_227,N_2737,N_2972);
and UO_228 (O_228,N_2756,N_2743);
nor UO_229 (O_229,N_2983,N_2658);
and UO_230 (O_230,N_2782,N_2309);
xnor UO_231 (O_231,N_2891,N_2284);
xor UO_232 (O_232,N_2959,N_2280);
xnor UO_233 (O_233,N_2832,N_2791);
nand UO_234 (O_234,N_2896,N_2622);
nand UO_235 (O_235,N_2674,N_2361);
or UO_236 (O_236,N_2440,N_2375);
nor UO_237 (O_237,N_2592,N_2544);
or UO_238 (O_238,N_2602,N_2497);
xor UO_239 (O_239,N_2508,N_2748);
nor UO_240 (O_240,N_2281,N_2601);
xor UO_241 (O_241,N_2798,N_2576);
xor UO_242 (O_242,N_2952,N_2724);
and UO_243 (O_243,N_2792,N_2372);
nor UO_244 (O_244,N_2333,N_2799);
nand UO_245 (O_245,N_2367,N_2851);
xnor UO_246 (O_246,N_2519,N_2965);
xor UO_247 (O_247,N_2423,N_2542);
nand UO_248 (O_248,N_2771,N_2777);
nor UO_249 (O_249,N_2567,N_2452);
or UO_250 (O_250,N_2664,N_2494);
nor UO_251 (O_251,N_2522,N_2744);
nand UO_252 (O_252,N_2849,N_2428);
xor UO_253 (O_253,N_2797,N_2897);
nor UO_254 (O_254,N_2591,N_2493);
and UO_255 (O_255,N_2696,N_2831);
and UO_256 (O_256,N_2438,N_2757);
and UO_257 (O_257,N_2708,N_2557);
and UO_258 (O_258,N_2563,N_2858);
xor UO_259 (O_259,N_2839,N_2966);
or UO_260 (O_260,N_2793,N_2462);
xor UO_261 (O_261,N_2318,N_2329);
and UO_262 (O_262,N_2337,N_2573);
nor UO_263 (O_263,N_2317,N_2637);
xnor UO_264 (O_264,N_2606,N_2545);
xnor UO_265 (O_265,N_2981,N_2303);
nor UO_266 (O_266,N_2809,N_2517);
xor UO_267 (O_267,N_2946,N_2900);
xnor UO_268 (O_268,N_2654,N_2646);
xnor UO_269 (O_269,N_2943,N_2698);
nor UO_270 (O_270,N_2263,N_2636);
or UO_271 (O_271,N_2653,N_2937);
or UO_272 (O_272,N_2480,N_2389);
and UO_273 (O_273,N_2595,N_2406);
nor UO_274 (O_274,N_2720,N_2925);
nand UO_275 (O_275,N_2272,N_2986);
and UO_276 (O_276,N_2893,N_2824);
and UO_277 (O_277,N_2467,N_2253);
nor UO_278 (O_278,N_2290,N_2298);
nor UO_279 (O_279,N_2628,N_2341);
and UO_280 (O_280,N_2401,N_2647);
xor UO_281 (O_281,N_2707,N_2559);
or UO_282 (O_282,N_2538,N_2994);
nor UO_283 (O_283,N_2806,N_2620);
and UO_284 (O_284,N_2430,N_2852);
and UO_285 (O_285,N_2495,N_2446);
nor UO_286 (O_286,N_2911,N_2630);
xor UO_287 (O_287,N_2381,N_2450);
or UO_288 (O_288,N_2784,N_2612);
and UO_289 (O_289,N_2594,N_2655);
and UO_290 (O_290,N_2922,N_2878);
and UO_291 (O_291,N_2814,N_2866);
and UO_292 (O_292,N_2549,N_2807);
nor UO_293 (O_293,N_2509,N_2448);
xor UO_294 (O_294,N_2681,N_2808);
and UO_295 (O_295,N_2890,N_2512);
nor UO_296 (O_296,N_2604,N_2484);
nand UO_297 (O_297,N_2566,N_2405);
or UO_298 (O_298,N_2269,N_2453);
nand UO_299 (O_299,N_2635,N_2362);
or UO_300 (O_300,N_2931,N_2609);
xor UO_301 (O_301,N_2827,N_2924);
or UO_302 (O_302,N_2718,N_2941);
nor UO_303 (O_303,N_2641,N_2691);
xnor UO_304 (O_304,N_2928,N_2789);
nand UO_305 (O_305,N_2686,N_2325);
and UO_306 (O_306,N_2834,N_2665);
nor UO_307 (O_307,N_2427,N_2346);
nand UO_308 (O_308,N_2334,N_2426);
and UO_309 (O_309,N_2732,N_2313);
or UO_310 (O_310,N_2444,N_2264);
xnor UO_311 (O_311,N_2532,N_2308);
xnor UO_312 (O_312,N_2464,N_2267);
xor UO_313 (O_313,N_2371,N_2960);
xor UO_314 (O_314,N_2949,N_2671);
xor UO_315 (O_315,N_2761,N_2629);
xor UO_316 (O_316,N_2842,N_2951);
nor UO_317 (O_317,N_2795,N_2385);
and UO_318 (O_318,N_2755,N_2651);
and UO_319 (O_319,N_2876,N_2560);
nor UO_320 (O_320,N_2546,N_2301);
and UO_321 (O_321,N_2523,N_2823);
nand UO_322 (O_322,N_2434,N_2734);
nand UO_323 (O_323,N_2569,N_2481);
and UO_324 (O_324,N_2478,N_2357);
nor UO_325 (O_325,N_2320,N_2587);
or UO_326 (O_326,N_2778,N_2706);
xor UO_327 (O_327,N_2419,N_2270);
nor UO_328 (O_328,N_2589,N_2349);
or UO_329 (O_329,N_2278,N_2913);
and UO_330 (O_330,N_2769,N_2857);
or UO_331 (O_331,N_2969,N_2916);
nor UO_332 (O_332,N_2377,N_2551);
or UO_333 (O_333,N_2285,N_2398);
nand UO_334 (O_334,N_2704,N_2501);
or UO_335 (O_335,N_2863,N_2976);
nand UO_336 (O_336,N_2880,N_2684);
xor UO_337 (O_337,N_2881,N_2762);
nor UO_338 (O_338,N_2835,N_2640);
or UO_339 (O_339,N_2487,N_2531);
nor UO_340 (O_340,N_2841,N_2690);
nor UO_341 (O_341,N_2291,N_2524);
nand UO_342 (O_342,N_2363,N_2351);
xor UO_343 (O_343,N_2350,N_2906);
or UO_344 (O_344,N_2355,N_2500);
nand UO_345 (O_345,N_2764,N_2603);
nor UO_346 (O_346,N_2310,N_2801);
and UO_347 (O_347,N_2621,N_2342);
nand UO_348 (O_348,N_2472,N_2408);
and UO_349 (O_349,N_2899,N_2657);
xor UO_350 (O_350,N_2288,N_2306);
nand UO_351 (O_351,N_2386,N_2805);
xor UO_352 (O_352,N_2376,N_2261);
nand UO_353 (O_353,N_2273,N_2923);
or UO_354 (O_354,N_2978,N_2460);
nor UO_355 (O_355,N_2957,N_2457);
nand UO_356 (O_356,N_2471,N_2618);
xor UO_357 (O_357,N_2260,N_2869);
xor UO_358 (O_358,N_2803,N_2358);
xor UO_359 (O_359,N_2751,N_2643);
nand UO_360 (O_360,N_2608,N_2368);
and UO_361 (O_361,N_2297,N_2816);
nand UO_362 (O_362,N_2614,N_2663);
nor UO_363 (O_363,N_2901,N_2918);
nor UO_364 (O_364,N_2713,N_2577);
or UO_365 (O_365,N_2393,N_2956);
nand UO_366 (O_366,N_2445,N_2340);
nand UO_367 (O_367,N_2980,N_2421);
nor UO_368 (O_368,N_2610,N_2593);
nand UO_369 (O_369,N_2370,N_2397);
nand UO_370 (O_370,N_2527,N_2848);
xnor UO_371 (O_371,N_2259,N_2667);
and UO_372 (O_372,N_2326,N_2905);
and UO_373 (O_373,N_2954,N_2468);
nand UO_374 (O_374,N_2510,N_2766);
nand UO_375 (O_375,N_2680,N_2469);
and UO_376 (O_376,N_2667,N_2534);
xnor UO_377 (O_377,N_2268,N_2972);
or UO_378 (O_378,N_2823,N_2789);
nand UO_379 (O_379,N_2797,N_2873);
and UO_380 (O_380,N_2657,N_2688);
xor UO_381 (O_381,N_2914,N_2949);
nor UO_382 (O_382,N_2476,N_2886);
xor UO_383 (O_383,N_2770,N_2341);
nand UO_384 (O_384,N_2708,N_2662);
and UO_385 (O_385,N_2403,N_2540);
nand UO_386 (O_386,N_2361,N_2896);
and UO_387 (O_387,N_2349,N_2545);
and UO_388 (O_388,N_2647,N_2668);
nor UO_389 (O_389,N_2325,N_2970);
or UO_390 (O_390,N_2823,N_2630);
or UO_391 (O_391,N_2744,N_2397);
and UO_392 (O_392,N_2413,N_2664);
and UO_393 (O_393,N_2455,N_2271);
xor UO_394 (O_394,N_2942,N_2282);
and UO_395 (O_395,N_2598,N_2760);
and UO_396 (O_396,N_2627,N_2321);
or UO_397 (O_397,N_2882,N_2621);
or UO_398 (O_398,N_2257,N_2824);
and UO_399 (O_399,N_2349,N_2283);
xor UO_400 (O_400,N_2519,N_2529);
xnor UO_401 (O_401,N_2922,N_2361);
nand UO_402 (O_402,N_2824,N_2789);
or UO_403 (O_403,N_2323,N_2463);
nor UO_404 (O_404,N_2524,N_2859);
and UO_405 (O_405,N_2354,N_2964);
nor UO_406 (O_406,N_2665,N_2988);
xnor UO_407 (O_407,N_2740,N_2449);
and UO_408 (O_408,N_2958,N_2663);
nor UO_409 (O_409,N_2265,N_2526);
nand UO_410 (O_410,N_2856,N_2943);
nand UO_411 (O_411,N_2579,N_2600);
xnor UO_412 (O_412,N_2533,N_2311);
nor UO_413 (O_413,N_2422,N_2900);
or UO_414 (O_414,N_2455,N_2894);
or UO_415 (O_415,N_2297,N_2719);
nor UO_416 (O_416,N_2298,N_2924);
nand UO_417 (O_417,N_2370,N_2781);
nor UO_418 (O_418,N_2615,N_2743);
nand UO_419 (O_419,N_2979,N_2578);
xnor UO_420 (O_420,N_2816,N_2689);
and UO_421 (O_421,N_2389,N_2957);
xnor UO_422 (O_422,N_2370,N_2403);
nand UO_423 (O_423,N_2523,N_2521);
nor UO_424 (O_424,N_2960,N_2910);
nand UO_425 (O_425,N_2557,N_2394);
or UO_426 (O_426,N_2270,N_2538);
or UO_427 (O_427,N_2946,N_2807);
nor UO_428 (O_428,N_2305,N_2408);
xnor UO_429 (O_429,N_2344,N_2467);
nand UO_430 (O_430,N_2551,N_2411);
or UO_431 (O_431,N_2705,N_2689);
nor UO_432 (O_432,N_2892,N_2384);
nand UO_433 (O_433,N_2789,N_2273);
nor UO_434 (O_434,N_2503,N_2521);
or UO_435 (O_435,N_2835,N_2750);
nand UO_436 (O_436,N_2903,N_2498);
and UO_437 (O_437,N_2916,N_2330);
and UO_438 (O_438,N_2983,N_2320);
nand UO_439 (O_439,N_2482,N_2398);
xor UO_440 (O_440,N_2373,N_2318);
nand UO_441 (O_441,N_2634,N_2694);
xnor UO_442 (O_442,N_2303,N_2557);
or UO_443 (O_443,N_2718,N_2754);
xor UO_444 (O_444,N_2864,N_2378);
xnor UO_445 (O_445,N_2289,N_2721);
nand UO_446 (O_446,N_2262,N_2499);
and UO_447 (O_447,N_2481,N_2490);
or UO_448 (O_448,N_2540,N_2387);
nor UO_449 (O_449,N_2618,N_2950);
nor UO_450 (O_450,N_2695,N_2310);
nor UO_451 (O_451,N_2351,N_2808);
nor UO_452 (O_452,N_2706,N_2940);
nor UO_453 (O_453,N_2676,N_2666);
xor UO_454 (O_454,N_2641,N_2618);
or UO_455 (O_455,N_2582,N_2666);
and UO_456 (O_456,N_2839,N_2741);
nor UO_457 (O_457,N_2761,N_2745);
xor UO_458 (O_458,N_2599,N_2787);
nand UO_459 (O_459,N_2510,N_2611);
nor UO_460 (O_460,N_2670,N_2256);
or UO_461 (O_461,N_2584,N_2501);
xor UO_462 (O_462,N_2364,N_2988);
or UO_463 (O_463,N_2437,N_2893);
and UO_464 (O_464,N_2707,N_2926);
nand UO_465 (O_465,N_2635,N_2906);
and UO_466 (O_466,N_2784,N_2529);
xnor UO_467 (O_467,N_2406,N_2965);
and UO_468 (O_468,N_2988,N_2865);
nor UO_469 (O_469,N_2864,N_2982);
or UO_470 (O_470,N_2489,N_2881);
and UO_471 (O_471,N_2940,N_2757);
or UO_472 (O_472,N_2432,N_2786);
or UO_473 (O_473,N_2526,N_2504);
and UO_474 (O_474,N_2996,N_2602);
nor UO_475 (O_475,N_2391,N_2387);
nor UO_476 (O_476,N_2451,N_2908);
and UO_477 (O_477,N_2615,N_2961);
nor UO_478 (O_478,N_2840,N_2325);
nor UO_479 (O_479,N_2545,N_2506);
or UO_480 (O_480,N_2587,N_2537);
nor UO_481 (O_481,N_2967,N_2866);
xor UO_482 (O_482,N_2917,N_2354);
or UO_483 (O_483,N_2733,N_2848);
xnor UO_484 (O_484,N_2293,N_2360);
and UO_485 (O_485,N_2824,N_2311);
nand UO_486 (O_486,N_2503,N_2413);
nand UO_487 (O_487,N_2815,N_2535);
nand UO_488 (O_488,N_2643,N_2260);
and UO_489 (O_489,N_2405,N_2779);
nand UO_490 (O_490,N_2967,N_2534);
and UO_491 (O_491,N_2913,N_2733);
and UO_492 (O_492,N_2947,N_2983);
and UO_493 (O_493,N_2772,N_2994);
nand UO_494 (O_494,N_2923,N_2800);
xor UO_495 (O_495,N_2644,N_2875);
nor UO_496 (O_496,N_2661,N_2721);
xnor UO_497 (O_497,N_2872,N_2923);
or UO_498 (O_498,N_2274,N_2477);
or UO_499 (O_499,N_2424,N_2466);
endmodule