module basic_1500_15000_2000_5_levels_1xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_794,In_1037);
or U1 (N_1,In_1162,In_44);
nor U2 (N_2,In_379,In_36);
and U3 (N_3,In_1253,In_1146);
nand U4 (N_4,In_82,In_1279);
and U5 (N_5,In_616,In_610);
or U6 (N_6,In_429,In_450);
nor U7 (N_7,In_678,In_1143);
and U8 (N_8,In_157,In_364);
nand U9 (N_9,In_700,In_611);
and U10 (N_10,In_772,In_966);
and U11 (N_11,In_1188,In_400);
and U12 (N_12,In_1415,In_735);
or U13 (N_13,In_107,In_1255);
and U14 (N_14,In_1335,In_1176);
nor U15 (N_15,In_171,In_147);
xor U16 (N_16,In_96,In_25);
nor U17 (N_17,In_211,In_447);
nand U18 (N_18,In_1205,In_949);
nand U19 (N_19,In_487,In_485);
nor U20 (N_20,In_1339,In_191);
nand U21 (N_21,In_560,In_961);
nor U22 (N_22,In_494,In_116);
nand U23 (N_23,In_456,In_838);
nor U24 (N_24,In_329,In_876);
or U25 (N_25,In_344,In_940);
nand U26 (N_26,In_1052,In_213);
nor U27 (N_27,In_1319,In_757);
and U28 (N_28,In_644,In_1252);
and U29 (N_29,In_279,In_1298);
or U30 (N_30,In_189,In_480);
nand U31 (N_31,In_1216,In_1151);
or U32 (N_32,In_597,In_811);
and U33 (N_33,In_1387,In_813);
nor U34 (N_34,In_40,In_1439);
and U35 (N_35,In_73,In_695);
nor U36 (N_36,In_1030,In_1442);
nor U37 (N_37,In_396,In_1425);
nand U38 (N_38,In_1196,In_1066);
nand U39 (N_39,In_579,In_35);
nor U40 (N_40,In_1383,In_412);
nor U41 (N_41,In_862,In_852);
and U42 (N_42,In_820,In_499);
nor U43 (N_43,In_51,In_1284);
and U44 (N_44,In_424,In_796);
nand U45 (N_45,In_657,In_1134);
nor U46 (N_46,In_655,In_42);
or U47 (N_47,In_1226,In_1189);
nand U48 (N_48,In_584,In_566);
nand U49 (N_49,In_1122,In_267);
nand U50 (N_50,In_1085,In_1330);
nor U51 (N_51,In_1103,In_495);
nor U52 (N_52,In_1104,In_615);
or U53 (N_53,In_284,In_679);
and U54 (N_54,In_1471,In_462);
and U55 (N_55,In_767,In_1469);
nor U56 (N_56,In_1013,In_1117);
and U57 (N_57,In_343,In_511);
or U58 (N_58,In_658,In_843);
nand U59 (N_59,In_88,In_1408);
and U60 (N_60,In_346,In_15);
and U61 (N_61,In_1126,In_355);
nor U62 (N_62,In_448,In_316);
nor U63 (N_63,In_633,In_369);
nand U64 (N_64,In_198,In_1435);
and U65 (N_65,In_605,In_713);
or U66 (N_66,In_926,In_1395);
or U67 (N_67,In_1398,In_8);
and U68 (N_68,In_287,In_588);
nand U69 (N_69,In_87,In_421);
or U70 (N_70,In_427,In_1076);
nor U71 (N_71,In_805,In_85);
nor U72 (N_72,In_1078,In_188);
nor U73 (N_73,In_1356,In_1479);
nor U74 (N_74,In_817,In_734);
and U75 (N_75,In_1108,In_259);
xnor U76 (N_76,In_234,In_722);
nand U77 (N_77,In_525,In_1424);
or U78 (N_78,In_760,In_1467);
nand U79 (N_79,In_310,In_620);
nor U80 (N_80,In_115,In_1083);
nor U81 (N_81,In_1263,In_870);
and U82 (N_82,In_11,In_240);
nand U83 (N_83,In_1265,In_306);
nor U84 (N_84,In_361,In_650);
and U85 (N_85,In_840,In_458);
or U86 (N_86,In_235,In_590);
nand U87 (N_87,In_223,In_124);
and U88 (N_88,In_634,In_1324);
nand U89 (N_89,In_1025,In_1266);
and U90 (N_90,In_1481,In_517);
or U91 (N_91,In_304,In_667);
or U92 (N_92,In_52,In_739);
nor U93 (N_93,In_676,In_1486);
nand U94 (N_94,In_842,In_380);
and U95 (N_95,In_163,In_1268);
and U96 (N_96,In_1341,In_309);
nand U97 (N_97,In_442,In_86);
and U98 (N_98,In_26,In_438);
nand U99 (N_99,In_1307,In_1305);
or U100 (N_100,In_604,In_1494);
and U101 (N_101,In_1049,In_652);
nand U102 (N_102,In_1109,In_375);
nor U103 (N_103,In_437,In_472);
and U104 (N_104,In_1296,In_1264);
and U105 (N_105,In_753,In_335);
or U106 (N_106,In_324,In_965);
nand U107 (N_107,In_715,In_801);
nand U108 (N_108,In_1292,In_272);
nor U109 (N_109,In_793,In_413);
or U110 (N_110,In_670,In_1212);
or U111 (N_111,In_166,In_210);
and U112 (N_112,In_420,In_866);
and U113 (N_113,In_768,In_1297);
and U114 (N_114,In_1115,In_270);
nor U115 (N_115,In_879,In_1453);
and U116 (N_116,In_815,In_20);
or U117 (N_117,In_514,In_617);
nor U118 (N_118,In_473,In_135);
or U119 (N_119,In_175,In_299);
nand U120 (N_120,In_798,In_405);
or U121 (N_121,In_1419,In_1051);
or U122 (N_122,In_573,In_901);
and U123 (N_123,In_1325,In_452);
or U124 (N_124,In_905,In_699);
and U125 (N_125,In_902,In_141);
or U126 (N_126,In_504,In_218);
or U127 (N_127,In_137,In_692);
or U128 (N_128,In_476,In_94);
nand U129 (N_129,In_673,In_698);
or U130 (N_130,In_185,In_155);
and U131 (N_131,In_72,In_933);
nor U132 (N_132,In_323,In_449);
nand U133 (N_133,In_580,In_505);
nor U134 (N_134,In_1254,In_880);
or U135 (N_135,In_22,In_1023);
nor U136 (N_136,In_732,In_626);
or U137 (N_137,In_809,In_935);
and U138 (N_138,In_194,In_30);
nor U139 (N_139,In_510,In_91);
and U140 (N_140,In_280,In_221);
and U141 (N_141,In_277,In_59);
nor U142 (N_142,In_4,In_745);
nor U143 (N_143,In_336,In_1300);
nor U144 (N_144,In_981,In_1154);
nor U145 (N_145,In_558,In_453);
nand U146 (N_146,In_1185,In_460);
or U147 (N_147,In_41,In_656);
nor U148 (N_148,In_1231,In_374);
nor U149 (N_149,In_1138,In_1239);
and U150 (N_150,In_998,In_1074);
or U151 (N_151,In_29,In_1369);
or U152 (N_152,In_747,In_50);
xnor U153 (N_153,In_1422,In_500);
and U154 (N_154,In_49,In_1147);
and U155 (N_155,In_1290,In_603);
or U156 (N_156,In_409,In_889);
or U157 (N_157,In_948,In_632);
or U158 (N_158,In_983,In_729);
xnor U159 (N_159,In_660,In_1357);
nor U160 (N_160,In_1396,In_112);
or U161 (N_161,In_868,In_1064);
nand U162 (N_162,In_1321,In_418);
and U163 (N_163,In_119,In_1044);
nand U164 (N_164,In_1179,In_716);
or U165 (N_165,In_482,In_1178);
nand U166 (N_166,In_985,In_627);
nand U167 (N_167,In_647,In_1145);
and U168 (N_168,In_984,In_321);
nor U169 (N_169,In_451,In_195);
nand U170 (N_170,In_1294,In_1441);
and U171 (N_171,In_106,In_992);
nand U172 (N_172,In_1436,In_170);
nand U173 (N_173,In_90,In_370);
nand U174 (N_174,In_1140,In_1372);
nor U175 (N_175,In_822,In_654);
or U176 (N_176,In_600,In_501);
nand U177 (N_177,In_1125,In_54);
and U178 (N_178,In_378,In_980);
nor U179 (N_179,In_704,In_792);
nand U180 (N_180,In_1116,In_1468);
and U181 (N_181,In_376,In_1149);
nor U182 (N_182,In_1423,In_1403);
and U183 (N_183,In_1135,In_239);
and U184 (N_184,In_204,In_1412);
nor U185 (N_185,In_382,In_1275);
nor U186 (N_186,In_152,In_1416);
nand U187 (N_187,In_710,In_964);
nor U188 (N_188,In_963,In_758);
nand U189 (N_189,In_553,In_407);
and U190 (N_190,In_75,In_896);
nand U191 (N_191,In_1080,In_1454);
nor U192 (N_192,In_1086,In_797);
or U193 (N_193,In_83,In_1092);
or U194 (N_194,In_907,In_542);
and U195 (N_195,In_457,In_1225);
or U196 (N_196,In_1096,In_23);
and U197 (N_197,In_489,In_1114);
nor U198 (N_198,In_111,In_1053);
or U199 (N_199,In_443,In_918);
or U200 (N_200,In_562,In_773);
nand U201 (N_201,In_996,In_283);
nand U202 (N_202,In_247,In_62);
and U203 (N_203,In_1337,In_1248);
or U204 (N_204,In_238,In_608);
nor U205 (N_205,In_21,In_1362);
and U206 (N_206,In_415,In_1353);
nor U207 (N_207,In_187,In_97);
and U208 (N_208,In_569,In_180);
nand U209 (N_209,In_1230,In_1458);
or U210 (N_210,In_78,In_268);
or U211 (N_211,In_1497,In_854);
and U212 (N_212,In_894,In_520);
and U213 (N_213,In_1437,In_1077);
nor U214 (N_214,In_289,In_691);
or U215 (N_215,In_1148,In_953);
or U216 (N_216,In_661,In_1198);
and U217 (N_217,In_954,In_850);
or U218 (N_218,In_799,In_1452);
or U219 (N_219,In_340,In_408);
nor U220 (N_220,In_664,In_215);
or U221 (N_221,In_1301,In_395);
or U222 (N_222,In_1048,In_183);
and U223 (N_223,In_790,In_1464);
nand U224 (N_224,In_623,In_1118);
or U225 (N_225,In_1244,In_1462);
nand U226 (N_226,In_737,In_174);
nand U227 (N_227,In_298,In_781);
nand U228 (N_228,In_1169,In_1318);
nand U229 (N_229,In_1182,In_1496);
nor U230 (N_230,In_131,In_242);
nor U231 (N_231,In_1120,In_911);
or U232 (N_232,In_1431,In_1009);
and U233 (N_233,In_76,In_574);
nand U234 (N_234,In_151,In_509);
or U235 (N_235,In_322,In_296);
and U236 (N_236,In_613,In_830);
and U237 (N_237,In_1152,In_977);
and U238 (N_238,In_751,In_554);
and U239 (N_239,In_432,In_292);
or U240 (N_240,In_601,In_1006);
nor U241 (N_241,In_1093,In_856);
nor U242 (N_242,In_269,In_467);
nor U243 (N_243,In_1336,In_461);
or U244 (N_244,In_498,In_341);
and U245 (N_245,In_176,In_784);
and U246 (N_246,In_28,In_1455);
or U247 (N_247,In_1043,In_1283);
nor U248 (N_248,In_1381,In_252);
nand U249 (N_249,In_65,In_317);
nand U250 (N_250,In_944,In_828);
or U251 (N_251,In_1022,In_102);
and U252 (N_252,In_356,In_744);
and U253 (N_253,In_971,In_313);
nor U254 (N_254,In_924,In_1032);
or U255 (N_255,In_548,In_6);
or U256 (N_256,In_728,In_960);
nand U257 (N_257,In_291,In_290);
and U258 (N_258,In_136,In_1012);
or U259 (N_259,In_463,In_1378);
or U260 (N_260,In_973,In_1312);
nand U261 (N_261,In_683,In_1488);
nor U262 (N_262,In_861,In_669);
nand U263 (N_263,In_503,In_1068);
or U264 (N_264,In_1180,In_64);
nand U265 (N_265,In_230,In_668);
xnor U266 (N_266,In_146,In_567);
and U267 (N_267,In_786,In_575);
and U268 (N_268,In_121,In_618);
or U269 (N_269,In_318,In_950);
nand U270 (N_270,In_591,In_783);
and U271 (N_271,In_551,In_161);
nand U272 (N_272,In_1081,In_1495);
nor U273 (N_273,In_1034,In_707);
and U274 (N_274,In_646,In_968);
and U275 (N_275,In_226,In_1172);
nand U276 (N_276,In_196,In_800);
and U277 (N_277,In_1262,In_1338);
or U278 (N_278,In_1465,In_1167);
and U279 (N_279,In_864,In_1367);
or U280 (N_280,In_63,In_513);
and U281 (N_281,In_888,In_771);
or U282 (N_282,In_1130,In_543);
or U283 (N_283,In_1221,In_168);
and U284 (N_284,In_465,In_422);
nor U285 (N_285,In_301,In_1240);
nand U286 (N_286,In_763,In_398);
nor U287 (N_287,In_696,In_975);
or U288 (N_288,In_1476,In_243);
and U289 (N_289,In_1366,In_987);
or U290 (N_290,In_937,In_1380);
nor U291 (N_291,In_74,In_1070);
and U292 (N_292,In_1021,In_1272);
nor U293 (N_293,In_172,In_821);
and U294 (N_294,In_570,In_552);
nor U295 (N_295,In_851,In_390);
or U296 (N_296,In_1327,In_261);
nor U297 (N_297,In_2,In_858);
and U298 (N_298,In_315,In_92);
nor U299 (N_299,In_496,In_571);
nand U300 (N_300,In_848,In_1207);
or U301 (N_301,In_1346,In_10);
or U302 (N_302,In_628,In_621);
nor U303 (N_303,In_526,In_406);
nand U304 (N_304,In_991,In_697);
and U305 (N_305,In_1157,In_913);
nand U306 (N_306,In_780,In_860);
nor U307 (N_307,In_1020,In_774);
xnor U308 (N_308,In_231,In_1177);
nor U309 (N_309,In_997,In_1087);
and U310 (N_310,In_648,In_662);
or U311 (N_311,In_764,In_140);
nor U312 (N_312,In_1133,In_1245);
nand U313 (N_313,In_1038,In_1379);
nand U314 (N_314,In_263,In_994);
nand U315 (N_315,In_1224,In_689);
nor U316 (N_316,In_593,In_743);
or U317 (N_317,In_1102,In_1163);
nand U318 (N_318,In_53,In_37);
nor U319 (N_319,In_769,In_1175);
or U320 (N_320,In_491,In_401);
or U321 (N_321,In_182,In_190);
nor U322 (N_322,In_589,In_557);
nor U323 (N_323,In_307,In_159);
nand U324 (N_324,In_779,In_24);
or U325 (N_325,In_990,In_1075);
and U326 (N_326,In_1128,In_148);
nand U327 (N_327,In_572,In_123);
and U328 (N_328,In_807,In_416);
and U329 (N_329,In_93,In_538);
nor U330 (N_330,In_81,In_1232);
nand U331 (N_331,In_1050,In_1215);
nor U332 (N_332,In_216,In_903);
nand U333 (N_333,In_1399,In_444);
and U334 (N_334,In_833,In_1348);
and U335 (N_335,In_727,In_77);
nor U336 (N_336,In_1098,In_1153);
or U337 (N_337,In_1417,In_459);
and U338 (N_338,In_320,In_167);
xnor U339 (N_339,In_651,In_976);
nand U340 (N_340,In_1235,In_359);
nand U341 (N_341,In_530,In_80);
nor U342 (N_342,In_849,In_712);
nor U343 (N_343,In_912,In_1384);
nor U344 (N_344,In_1474,In_1273);
or U345 (N_345,In_474,In_57);
nand U346 (N_346,In_430,In_1282);
and U347 (N_347,In_1041,In_855);
or U348 (N_348,In_1256,In_1413);
or U349 (N_349,In_865,In_1127);
or U350 (N_350,In_1069,In_731);
or U351 (N_351,In_909,In_431);
nand U352 (N_352,In_711,In_1490);
or U353 (N_353,In_425,In_1472);
nand U354 (N_354,In_599,In_193);
and U355 (N_355,In_1061,In_362);
or U356 (N_356,In_469,In_1187);
nor U357 (N_357,In_587,In_671);
and U358 (N_358,In_1027,In_349);
and U359 (N_359,In_104,In_222);
nand U360 (N_360,In_775,In_1332);
and U361 (N_361,In_47,In_789);
nand U362 (N_362,In_1036,In_1040);
and U363 (N_363,In_1402,In_921);
nand U364 (N_364,In_232,In_470);
and U365 (N_365,In_791,In_411);
nor U366 (N_366,In_1160,In_1042);
or U367 (N_367,In_14,In_1371);
nand U368 (N_368,In_393,In_1161);
and U369 (N_369,In_549,In_1035);
or U370 (N_370,In_1352,In_1101);
nor U371 (N_371,In_1368,In_56);
or U372 (N_372,In_874,In_1234);
or U373 (N_373,In_1004,In_528);
and U374 (N_374,In_1391,In_1063);
and U375 (N_375,In_1440,In_1055);
or U376 (N_376,In_1426,In_675);
nor U377 (N_377,In_1123,In_348);
nand U378 (N_378,In_563,In_1446);
and U379 (N_379,In_122,In_1438);
nor U380 (N_380,In_1241,In_908);
nand U381 (N_381,In_585,In_643);
or U382 (N_382,In_1113,In_607);
or U383 (N_383,In_99,In_512);
nor U384 (N_384,In_682,In_748);
nand U385 (N_385,In_177,In_873);
or U386 (N_386,In_684,In_1156);
nor U387 (N_387,In_598,In_829);
nand U388 (N_388,In_947,In_1447);
and U389 (N_389,In_1173,In_314);
nand U390 (N_390,In_1026,In_265);
nand U391 (N_391,In_885,In_441);
and U392 (N_392,In_943,In_900);
nor U393 (N_393,In_1124,In_1278);
nor U394 (N_394,In_612,In_1267);
nand U395 (N_395,In_67,In_1394);
and U396 (N_396,In_319,In_66);
and U397 (N_397,In_802,In_445);
and U398 (N_398,In_19,In_788);
nor U399 (N_399,In_1045,In_1106);
and U400 (N_400,In_392,In_55);
nand U401 (N_401,In_819,In_1259);
or U402 (N_402,In_1158,In_1445);
or U403 (N_403,In_529,In_1320);
and U404 (N_404,In_98,In_352);
nand U405 (N_405,In_701,In_545);
nand U406 (N_406,In_824,In_875);
nor U407 (N_407,In_931,In_351);
nor U408 (N_408,In_1010,In_1406);
nor U409 (N_409,In_39,In_297);
and U410 (N_410,In_426,In_845);
and U411 (N_411,In_200,In_1223);
xor U412 (N_412,In_1411,In_224);
nand U413 (N_413,In_844,In_1202);
and U414 (N_414,In_1277,In_1095);
nand U415 (N_415,In_7,In_179);
and U416 (N_416,In_1466,In_1191);
nor U417 (N_417,In_1091,In_1463);
or U418 (N_418,In_1112,In_100);
nand U419 (N_419,In_127,In_1386);
nand U420 (N_420,In_1475,In_878);
nor U421 (N_421,In_160,In_659);
or U422 (N_422,In_1480,In_1477);
and U423 (N_423,In_33,In_872);
and U424 (N_424,In_1129,In_1203);
and U425 (N_425,In_154,In_1105);
or U426 (N_426,In_206,In_1190);
or U427 (N_427,In_665,In_1342);
or U428 (N_428,In_726,In_1473);
nand U429 (N_429,In_1005,In_372);
nand U430 (N_430,In_714,In_736);
or U431 (N_431,In_1249,In_433);
nand U432 (N_432,In_423,In_540);
nand U433 (N_433,In_1388,In_978);
nand U434 (N_434,In_752,In_345);
nor U435 (N_435,In_776,In_688);
or U436 (N_436,In_826,In_740);
nand U437 (N_437,In_244,In_150);
and U438 (N_438,In_955,In_446);
and U439 (N_439,In_114,In_1304);
nand U440 (N_440,In_1432,In_165);
nand U441 (N_441,In_32,In_1291);
nand U442 (N_442,In_1355,In_1159);
and U443 (N_443,In_666,In_619);
and U444 (N_444,In_381,In_831);
and U445 (N_445,In_1016,In_302);
or U446 (N_446,In_1186,In_945);
or U447 (N_447,In_582,In_1323);
nor U448 (N_448,In_834,In_1450);
and U449 (N_449,In_142,In_1459);
and U450 (N_450,In_867,In_0);
nand U451 (N_451,In_256,In_761);
and U452 (N_452,In_846,In_233);
and U453 (N_453,In_338,In_1246);
or U454 (N_454,In_818,In_730);
nand U455 (N_455,In_755,In_625);
nand U456 (N_456,In_103,In_1168);
or U457 (N_457,In_1329,In_1420);
nand U458 (N_458,In_832,In_1326);
nand U459 (N_459,In_1349,In_1197);
and U460 (N_460,In_565,In_386);
and U461 (N_461,In_1311,In_1410);
or U462 (N_462,In_910,In_946);
nor U463 (N_463,In_914,In_559);
or U464 (N_464,In_1456,In_1247);
and U465 (N_465,In_31,In_839);
or U466 (N_466,In_254,In_326);
or U467 (N_467,In_1200,In_237);
or U468 (N_468,In_248,In_787);
or U469 (N_469,In_337,In_404);
nand U470 (N_470,In_178,In_389);
and U471 (N_471,In_419,In_785);
nor U472 (N_472,In_506,In_347);
or U473 (N_473,In_533,In_539);
or U474 (N_474,In_576,In_892);
and U475 (N_475,In_1201,In_217);
nand U476 (N_476,In_568,In_1409);
nand U477 (N_477,In_835,In_1316);
and U478 (N_478,In_464,In_920);
or U479 (N_479,In_1288,In_738);
nor U480 (N_480,In_592,In_521);
or U481 (N_481,In_982,In_162);
xor U482 (N_482,In_823,In_1236);
nand U483 (N_483,In_1195,In_1062);
nand U484 (N_484,In_622,In_354);
xnor U485 (N_485,In_479,In_71);
or U486 (N_486,In_756,In_795);
and U487 (N_487,In_1181,In_1213);
or U488 (N_488,In_311,In_1056);
xnor U489 (N_489,In_1390,In_202);
and U490 (N_490,In_132,In_1217);
nand U491 (N_491,In_749,In_1171);
or U492 (N_492,In_645,In_951);
or U493 (N_493,In_1222,In_484);
and U494 (N_494,In_967,In_979);
or U495 (N_495,In_368,In_1132);
nor U496 (N_496,In_929,In_1489);
or U497 (N_497,In_932,In_1270);
or U498 (N_498,In_881,In_1033);
nand U499 (N_499,In_934,In_1347);
nor U500 (N_500,In_1392,In_1242);
nor U501 (N_501,In_1460,In_1059);
or U502 (N_502,In_331,In_899);
nand U503 (N_503,In_1155,In_930);
or U504 (N_504,In_255,In_522);
and U505 (N_505,In_523,In_810);
nand U506 (N_506,In_1429,In_917);
nor U507 (N_507,In_1039,In_928);
and U508 (N_508,In_249,In_1377);
and U509 (N_509,In_923,In_1280);
or U510 (N_510,In_391,In_1094);
nor U511 (N_511,In_471,In_1003);
and U512 (N_512,In_95,In_260);
and U513 (N_513,In_1443,In_271);
or U514 (N_514,In_212,In_1233);
nor U515 (N_515,In_286,In_723);
nand U516 (N_516,In_535,In_1260);
nor U517 (N_517,In_1088,In_890);
nand U518 (N_518,In_101,In_541);
nand U519 (N_519,In_1204,In_640);
or U520 (N_520,In_827,In_435);
nand U521 (N_521,In_1054,In_5);
or U522 (N_522,In_1089,In_718);
nand U523 (N_523,In_962,In_118);
or U524 (N_524,In_759,In_1360);
nor U525 (N_525,In_1449,In_241);
and U526 (N_526,In_897,In_1071);
nand U527 (N_527,In_502,In_1418);
and U528 (N_528,In_886,In_1261);
xor U529 (N_529,In_898,In_332);
nand U530 (N_530,In_493,In_606);
nor U531 (N_531,In_266,In_969);
and U532 (N_532,In_12,In_1018);
nor U533 (N_533,In_139,In_884);
nor U534 (N_534,In_125,In_1276);
and U535 (N_535,In_956,In_1073);
or U536 (N_536,In_1218,In_614);
nand U537 (N_537,In_468,In_79);
or U538 (N_538,In_1219,In_1271);
nor U539 (N_539,In_869,In_1111);
and U540 (N_540,In_806,In_1015);
nand U541 (N_541,In_1002,In_537);
nand U542 (N_542,In_203,In_328);
nand U543 (N_543,In_1482,In_1310);
nand U544 (N_544,In_1199,In_693);
and U545 (N_545,In_1139,In_555);
nor U546 (N_546,In_253,In_719);
and U547 (N_547,In_816,In_782);
or U548 (N_548,In_532,In_721);
nor U549 (N_549,In_350,In_915);
nor U550 (N_550,In_516,In_305);
and U551 (N_551,In_1174,In_518);
nand U552 (N_552,In_108,In_577);
nor U553 (N_553,In_486,In_365);
and U554 (N_554,In_988,In_120);
or U555 (N_555,In_158,In_534);
and U556 (N_556,In_536,In_702);
nor U557 (N_557,In_995,In_906);
nand U558 (N_558,In_629,In_925);
and U559 (N_559,In_293,In_245);
and U560 (N_560,In_274,In_1322);
nand U561 (N_561,In_1451,In_273);
or U562 (N_562,In_209,In_282);
nor U563 (N_563,In_1011,In_1485);
or U564 (N_564,In_48,In_970);
and U565 (N_565,In_109,In_531);
nor U566 (N_566,In_1404,In_1315);
or U567 (N_567,In_746,In_1350);
or U568 (N_568,In_208,In_1499);
nand U569 (N_569,In_1306,In_281);
and U570 (N_570,In_871,In_680);
and U571 (N_571,In_250,In_750);
and U572 (N_572,In_1286,In_1487);
and U573 (N_573,In_1192,In_1028);
and U574 (N_574,In_1328,In_1457);
or U575 (N_575,In_1314,In_825);
nor U576 (N_576,In_681,In_402);
nor U577 (N_577,In_1150,In_1100);
or U578 (N_578,In_1427,In_207);
nand U579 (N_579,In_1082,In_1433);
or U580 (N_580,In_105,In_672);
nor U581 (N_581,In_857,In_229);
and U582 (N_582,In_371,In_578);
nor U583 (N_583,In_45,In_1401);
or U584 (N_584,In_1029,In_1484);
nor U585 (N_585,In_957,In_295);
and U586 (N_586,In_993,In_434);
nor U587 (N_587,In_687,In_1414);
nor U588 (N_588,In_1375,In_1370);
and U589 (N_589,In_1385,In_84);
nand U590 (N_590,In_1001,In_1057);
nor U591 (N_591,In_214,In_360);
nor U592 (N_592,In_1193,In_1046);
or U593 (N_593,In_1165,In_89);
nand U594 (N_594,In_129,In_808);
or U595 (N_595,In_1299,In_936);
nor U596 (N_596,In_725,In_145);
nor U597 (N_597,In_547,In_1345);
or U598 (N_598,In_507,In_853);
or U599 (N_599,In_524,In_1492);
nor U600 (N_600,In_1250,In_804);
or U601 (N_601,In_1359,In_1428);
nand U602 (N_602,In_1214,In_1493);
nand U603 (N_603,In_724,In_1097);
and U604 (N_604,In_262,In_636);
nand U605 (N_605,In_1363,In_134);
nor U606 (N_606,In_778,In_492);
nand U607 (N_607,In_300,In_1206);
nor U608 (N_608,In_1364,In_164);
and U609 (N_609,In_417,In_938);
or U610 (N_610,In_1065,In_397);
nor U611 (N_611,In_1008,In_303);
nor U612 (N_612,In_919,In_126);
nor U613 (N_613,In_596,In_327);
or U614 (N_614,In_916,In_1470);
or U615 (N_615,In_1483,In_227);
nor U616 (N_616,In_1397,In_941);
nor U617 (N_617,In_1024,In_720);
nand U618 (N_618,In_477,In_153);
nand U619 (N_619,In_637,In_1331);
and U620 (N_620,In_490,In_288);
nor U621 (N_621,In_1227,In_564);
or U622 (N_622,In_387,In_863);
and U623 (N_623,In_18,In_481);
or U624 (N_624,In_638,In_766);
nand U625 (N_625,In_246,In_803);
or U626 (N_626,In_594,In_373);
nand U627 (N_627,In_595,In_1274);
or U628 (N_628,In_475,In_1090);
nand U629 (N_629,In_1293,In_1258);
xor U630 (N_630,In_43,In_1211);
nor U631 (N_631,In_184,In_497);
nor U632 (N_632,In_974,In_1137);
and U633 (N_633,In_1170,In_1);
nor U634 (N_634,In_388,In_762);
nor U635 (N_635,In_837,In_1400);
and U636 (N_636,In_770,In_143);
nand U637 (N_637,In_922,In_353);
and U638 (N_638,In_1308,In_1121);
or U639 (N_639,In_61,In_765);
or U640 (N_640,In_1478,In_706);
and U641 (N_641,In_1194,In_228);
nor U642 (N_642,In_841,In_891);
nor U643 (N_643,In_1210,In_1084);
nor U644 (N_644,In_1141,In_3);
nor U645 (N_645,In_893,In_1303);
nand U646 (N_646,In_225,In_34);
or U647 (N_647,In_58,In_410);
or U648 (N_648,In_358,In_1269);
or U649 (N_649,In_1072,In_708);
and U650 (N_650,In_649,In_1334);
and U651 (N_651,In_113,In_1376);
or U652 (N_652,In_653,In_1354);
or U653 (N_653,In_635,In_952);
nand U654 (N_654,In_27,In_414);
and U655 (N_655,In_330,In_385);
nor U656 (N_656,In_236,In_859);
nand U657 (N_657,In_561,In_717);
or U658 (N_658,In_363,In_927);
and U659 (N_659,In_186,In_399);
nor U660 (N_660,In_882,In_1382);
or U661 (N_661,In_1251,In_439);
and U662 (N_662,In_1067,In_1498);
nand U663 (N_663,In_690,In_38);
nand U664 (N_664,In_483,In_192);
or U665 (N_665,In_904,In_1281);
or U666 (N_666,In_958,In_1119);
nor U667 (N_667,In_703,In_1491);
or U668 (N_668,In_1434,In_1344);
or U669 (N_669,In_339,In_285);
nand U670 (N_670,In_677,In_384);
nor U671 (N_671,In_1144,In_939);
nor U672 (N_672,In_199,In_1309);
and U673 (N_673,In_1361,In_488);
nand U674 (N_674,In_1358,In_130);
and U675 (N_675,In_455,In_519);
and U676 (N_676,In_440,In_733);
nor U677 (N_677,In_1351,In_1405);
and U678 (N_678,In_1131,In_1058);
nor U679 (N_679,In_639,In_1365);
or U680 (N_680,In_1238,In_586);
and U681 (N_681,In_686,In_128);
or U682 (N_682,In_334,In_16);
nor U683 (N_683,In_60,In_1430);
and U684 (N_684,In_133,In_877);
nor U685 (N_685,In_972,In_1285);
or U686 (N_686,In_709,In_989);
nor U687 (N_687,In_1184,In_357);
nor U688 (N_688,In_1220,In_1208);
or U689 (N_689,In_144,In_1000);
nand U690 (N_690,In_1079,In_403);
nor U691 (N_691,In_602,In_219);
or U692 (N_692,In_13,In_197);
nor U693 (N_693,In_377,In_69);
nor U694 (N_694,In_1107,In_1209);
nand U695 (N_695,In_1237,In_895);
or U696 (N_696,In_1228,In_325);
and U697 (N_697,In_308,In_220);
and U698 (N_698,In_812,In_1448);
and U699 (N_699,In_333,In_986);
or U700 (N_700,In_436,In_276);
and U701 (N_701,In_1461,In_181);
nor U702 (N_702,In_1289,In_70);
nand U703 (N_703,In_149,In_366);
nand U704 (N_704,In_544,In_546);
nand U705 (N_705,In_9,In_367);
nor U706 (N_706,In_1317,In_883);
and U707 (N_707,In_312,In_1243);
nor U708 (N_708,In_1444,In_631);
and U709 (N_709,In_466,In_454);
or U710 (N_710,In_742,In_556);
or U711 (N_711,In_527,In_624);
nor U712 (N_712,In_741,In_694);
or U713 (N_713,In_847,In_581);
or U714 (N_714,In_17,In_278);
and U715 (N_715,In_138,In_1060);
nor U716 (N_716,In_609,In_1166);
xnor U717 (N_717,In_1019,In_1333);
nand U718 (N_718,In_1183,In_1343);
or U719 (N_719,In_394,In_1257);
or U720 (N_720,In_1099,In_630);
nand U721 (N_721,In_342,In_814);
and U722 (N_722,In_1295,In_836);
or U723 (N_723,In_1302,In_515);
nand U724 (N_724,In_583,In_428);
or U725 (N_725,In_251,In_201);
and U726 (N_726,In_508,In_674);
nand U727 (N_727,In_1110,In_1287);
and U728 (N_728,In_294,In_1031);
nand U729 (N_729,In_173,In_275);
and U730 (N_730,In_999,In_110);
or U731 (N_731,In_887,In_550);
and U732 (N_732,In_959,In_478);
nor U733 (N_733,In_1373,In_1014);
or U734 (N_734,In_1313,In_1017);
or U735 (N_735,In_383,In_1407);
and U736 (N_736,In_169,In_156);
and U737 (N_737,In_663,In_754);
nor U738 (N_738,In_642,In_68);
nand U739 (N_739,In_942,In_1374);
nor U740 (N_740,In_685,In_1164);
and U741 (N_741,In_258,In_641);
nor U742 (N_742,In_1142,In_705);
nand U743 (N_743,In_257,In_1421);
nor U744 (N_744,In_1047,In_777);
nand U745 (N_745,In_264,In_205);
and U746 (N_746,In_1389,In_1136);
nor U747 (N_747,In_1229,In_1340);
and U748 (N_748,In_117,In_46);
and U749 (N_749,In_1393,In_1007);
nand U750 (N_750,In_6,In_1145);
nor U751 (N_751,In_529,In_897);
nand U752 (N_752,In_938,In_697);
or U753 (N_753,In_302,In_688);
and U754 (N_754,In_708,In_1477);
and U755 (N_755,In_1170,In_1099);
and U756 (N_756,In_472,In_896);
nor U757 (N_757,In_1490,In_832);
nand U758 (N_758,In_1148,In_1464);
nand U759 (N_759,In_1211,In_1001);
and U760 (N_760,In_635,In_540);
nor U761 (N_761,In_1307,In_743);
or U762 (N_762,In_1202,In_1129);
and U763 (N_763,In_662,In_1352);
and U764 (N_764,In_806,In_928);
or U765 (N_765,In_251,In_529);
nor U766 (N_766,In_69,In_424);
nand U767 (N_767,In_635,In_859);
nand U768 (N_768,In_78,In_267);
nor U769 (N_769,In_161,In_654);
and U770 (N_770,In_1410,In_1435);
or U771 (N_771,In_235,In_1148);
nor U772 (N_772,In_1396,In_386);
nor U773 (N_773,In_565,In_706);
nand U774 (N_774,In_720,In_1388);
or U775 (N_775,In_584,In_81);
and U776 (N_776,In_448,In_728);
nor U777 (N_777,In_245,In_487);
nand U778 (N_778,In_5,In_929);
or U779 (N_779,In_1438,In_242);
or U780 (N_780,In_671,In_944);
nor U781 (N_781,In_243,In_1462);
nand U782 (N_782,In_1202,In_312);
nand U783 (N_783,In_920,In_59);
nor U784 (N_784,In_1177,In_78);
and U785 (N_785,In_112,In_817);
and U786 (N_786,In_1228,In_1233);
nor U787 (N_787,In_1377,In_1265);
and U788 (N_788,In_648,In_90);
or U789 (N_789,In_128,In_417);
nand U790 (N_790,In_423,In_1102);
and U791 (N_791,In_243,In_484);
and U792 (N_792,In_900,In_235);
nand U793 (N_793,In_539,In_1185);
nand U794 (N_794,In_569,In_121);
or U795 (N_795,In_1243,In_236);
nand U796 (N_796,In_331,In_628);
nor U797 (N_797,In_1392,In_111);
and U798 (N_798,In_1398,In_1054);
nand U799 (N_799,In_510,In_207);
nand U800 (N_800,In_366,In_458);
or U801 (N_801,In_527,In_1046);
nor U802 (N_802,In_643,In_120);
and U803 (N_803,In_1310,In_289);
nand U804 (N_804,In_584,In_985);
nor U805 (N_805,In_711,In_733);
nor U806 (N_806,In_743,In_336);
nand U807 (N_807,In_792,In_1487);
nor U808 (N_808,In_496,In_708);
nand U809 (N_809,In_1005,In_216);
nand U810 (N_810,In_870,In_152);
nand U811 (N_811,In_954,In_1344);
or U812 (N_812,In_729,In_432);
nand U813 (N_813,In_706,In_992);
and U814 (N_814,In_242,In_477);
nand U815 (N_815,In_15,In_12);
and U816 (N_816,In_941,In_73);
nor U817 (N_817,In_778,In_153);
nor U818 (N_818,In_646,In_900);
nor U819 (N_819,In_1325,In_448);
and U820 (N_820,In_964,In_904);
and U821 (N_821,In_1176,In_1194);
nor U822 (N_822,In_601,In_686);
nor U823 (N_823,In_775,In_41);
nor U824 (N_824,In_781,In_1009);
nand U825 (N_825,In_971,In_736);
and U826 (N_826,In_692,In_1030);
and U827 (N_827,In_285,In_304);
or U828 (N_828,In_522,In_1393);
nand U829 (N_829,In_124,In_1477);
or U830 (N_830,In_785,In_543);
and U831 (N_831,In_1451,In_283);
nand U832 (N_832,In_1021,In_253);
and U833 (N_833,In_1368,In_227);
nor U834 (N_834,In_1098,In_1382);
or U835 (N_835,In_591,In_666);
nand U836 (N_836,In_181,In_65);
nand U837 (N_837,In_1461,In_1343);
nor U838 (N_838,In_507,In_646);
and U839 (N_839,In_1049,In_320);
nand U840 (N_840,In_885,In_1327);
or U841 (N_841,In_870,In_802);
or U842 (N_842,In_908,In_214);
nand U843 (N_843,In_972,In_1297);
nand U844 (N_844,In_291,In_1055);
nor U845 (N_845,In_245,In_1406);
nor U846 (N_846,In_1138,In_155);
and U847 (N_847,In_700,In_600);
nand U848 (N_848,In_341,In_1319);
nand U849 (N_849,In_1259,In_516);
nor U850 (N_850,In_1237,In_1494);
or U851 (N_851,In_94,In_943);
or U852 (N_852,In_1461,In_229);
nand U853 (N_853,In_857,In_55);
nor U854 (N_854,In_1093,In_465);
or U855 (N_855,In_575,In_27);
nand U856 (N_856,In_555,In_1064);
or U857 (N_857,In_527,In_999);
and U858 (N_858,In_1244,In_881);
nand U859 (N_859,In_429,In_63);
nand U860 (N_860,In_1265,In_1238);
nor U861 (N_861,In_478,In_509);
and U862 (N_862,In_64,In_226);
or U863 (N_863,In_600,In_822);
xnor U864 (N_864,In_905,In_954);
and U865 (N_865,In_1288,In_122);
and U866 (N_866,In_1440,In_1305);
or U867 (N_867,In_845,In_904);
and U868 (N_868,In_55,In_611);
or U869 (N_869,In_514,In_334);
or U870 (N_870,In_1204,In_909);
nand U871 (N_871,In_982,In_557);
nor U872 (N_872,In_858,In_233);
nor U873 (N_873,In_284,In_868);
nor U874 (N_874,In_1043,In_751);
nand U875 (N_875,In_415,In_1032);
nand U876 (N_876,In_1405,In_124);
xnor U877 (N_877,In_316,In_127);
and U878 (N_878,In_537,In_817);
or U879 (N_879,In_815,In_201);
and U880 (N_880,In_502,In_481);
nor U881 (N_881,In_949,In_554);
and U882 (N_882,In_669,In_794);
or U883 (N_883,In_98,In_641);
nand U884 (N_884,In_186,In_22);
nor U885 (N_885,In_1270,In_252);
and U886 (N_886,In_942,In_71);
nor U887 (N_887,In_1144,In_695);
nand U888 (N_888,In_1311,In_388);
and U889 (N_889,In_613,In_647);
and U890 (N_890,In_27,In_1029);
or U891 (N_891,In_378,In_1215);
or U892 (N_892,In_15,In_1096);
nor U893 (N_893,In_79,In_276);
nand U894 (N_894,In_356,In_949);
nand U895 (N_895,In_1291,In_829);
nor U896 (N_896,In_1285,In_497);
nand U897 (N_897,In_1437,In_724);
and U898 (N_898,In_881,In_68);
or U899 (N_899,In_480,In_1357);
xor U900 (N_900,In_1246,In_1433);
and U901 (N_901,In_1145,In_864);
or U902 (N_902,In_1222,In_1475);
nand U903 (N_903,In_1339,In_1072);
and U904 (N_904,In_68,In_1032);
nor U905 (N_905,In_916,In_861);
or U906 (N_906,In_288,In_947);
nor U907 (N_907,In_1254,In_997);
or U908 (N_908,In_439,In_917);
or U909 (N_909,In_140,In_100);
or U910 (N_910,In_1162,In_1105);
and U911 (N_911,In_679,In_601);
nand U912 (N_912,In_676,In_218);
and U913 (N_913,In_187,In_402);
nor U914 (N_914,In_793,In_629);
or U915 (N_915,In_369,In_266);
and U916 (N_916,In_706,In_923);
nor U917 (N_917,In_1271,In_1147);
nand U918 (N_918,In_293,In_1480);
and U919 (N_919,In_308,In_181);
nor U920 (N_920,In_1130,In_1333);
and U921 (N_921,In_1243,In_878);
nand U922 (N_922,In_1275,In_903);
nor U923 (N_923,In_1464,In_1273);
nor U924 (N_924,In_1097,In_387);
and U925 (N_925,In_264,In_1415);
nor U926 (N_926,In_184,In_398);
nand U927 (N_927,In_1020,In_1141);
nand U928 (N_928,In_463,In_1146);
or U929 (N_929,In_1404,In_873);
nor U930 (N_930,In_1492,In_866);
or U931 (N_931,In_1124,In_798);
nor U932 (N_932,In_395,In_259);
nor U933 (N_933,In_1143,In_295);
nor U934 (N_934,In_1000,In_428);
or U935 (N_935,In_1146,In_93);
nand U936 (N_936,In_704,In_271);
nand U937 (N_937,In_417,In_1094);
or U938 (N_938,In_861,In_239);
or U939 (N_939,In_42,In_30);
nand U940 (N_940,In_25,In_1085);
nand U941 (N_941,In_1235,In_94);
or U942 (N_942,In_1419,In_1135);
nor U943 (N_943,In_746,In_507);
or U944 (N_944,In_1470,In_460);
nor U945 (N_945,In_498,In_146);
or U946 (N_946,In_176,In_298);
or U947 (N_947,In_557,In_710);
and U948 (N_948,In_791,In_559);
nand U949 (N_949,In_1030,In_1265);
nor U950 (N_950,In_249,In_913);
or U951 (N_951,In_1,In_603);
nand U952 (N_952,In_262,In_550);
nor U953 (N_953,In_1086,In_1184);
nor U954 (N_954,In_685,In_618);
nand U955 (N_955,In_238,In_992);
and U956 (N_956,In_1174,In_914);
or U957 (N_957,In_1491,In_675);
or U958 (N_958,In_762,In_1287);
nor U959 (N_959,In_809,In_117);
and U960 (N_960,In_1274,In_1175);
nor U961 (N_961,In_471,In_354);
nand U962 (N_962,In_1319,In_254);
nand U963 (N_963,In_441,In_961);
nand U964 (N_964,In_925,In_1324);
nand U965 (N_965,In_520,In_833);
and U966 (N_966,In_1410,In_925);
and U967 (N_967,In_97,In_1155);
and U968 (N_968,In_6,In_157);
or U969 (N_969,In_849,In_730);
or U970 (N_970,In_649,In_237);
nor U971 (N_971,In_166,In_63);
nand U972 (N_972,In_781,In_414);
and U973 (N_973,In_1101,In_1045);
or U974 (N_974,In_154,In_827);
or U975 (N_975,In_427,In_1281);
nor U976 (N_976,In_740,In_1346);
and U977 (N_977,In_148,In_511);
nand U978 (N_978,In_247,In_1457);
and U979 (N_979,In_1330,In_536);
nand U980 (N_980,In_639,In_151);
nor U981 (N_981,In_1265,In_362);
and U982 (N_982,In_330,In_1382);
nor U983 (N_983,In_32,In_817);
or U984 (N_984,In_531,In_415);
or U985 (N_985,In_570,In_612);
or U986 (N_986,In_122,In_711);
or U987 (N_987,In_1078,In_331);
nor U988 (N_988,In_1471,In_824);
nand U989 (N_989,In_1024,In_576);
and U990 (N_990,In_918,In_1284);
and U991 (N_991,In_878,In_1324);
and U992 (N_992,In_1179,In_417);
nand U993 (N_993,In_955,In_273);
nor U994 (N_994,In_1329,In_12);
nand U995 (N_995,In_6,In_322);
and U996 (N_996,In_1305,In_1483);
nand U997 (N_997,In_20,In_543);
xnor U998 (N_998,In_1032,In_125);
or U999 (N_999,In_338,In_1316);
nor U1000 (N_1000,In_1335,In_194);
and U1001 (N_1001,In_842,In_928);
and U1002 (N_1002,In_289,In_708);
nand U1003 (N_1003,In_50,In_78);
or U1004 (N_1004,In_1050,In_245);
nand U1005 (N_1005,In_620,In_713);
and U1006 (N_1006,In_721,In_496);
or U1007 (N_1007,In_119,In_1264);
and U1008 (N_1008,In_607,In_1205);
or U1009 (N_1009,In_634,In_1229);
nor U1010 (N_1010,In_833,In_626);
nor U1011 (N_1011,In_45,In_1320);
nand U1012 (N_1012,In_1425,In_1137);
nor U1013 (N_1013,In_571,In_460);
or U1014 (N_1014,In_1172,In_417);
and U1015 (N_1015,In_1265,In_151);
nand U1016 (N_1016,In_1017,In_259);
nor U1017 (N_1017,In_473,In_211);
or U1018 (N_1018,In_1324,In_816);
nor U1019 (N_1019,In_1315,In_749);
nor U1020 (N_1020,In_804,In_1471);
and U1021 (N_1021,In_210,In_409);
nand U1022 (N_1022,In_439,In_1195);
nand U1023 (N_1023,In_889,In_267);
and U1024 (N_1024,In_1069,In_1001);
nor U1025 (N_1025,In_1053,In_733);
nor U1026 (N_1026,In_294,In_1120);
nor U1027 (N_1027,In_430,In_1092);
nor U1028 (N_1028,In_1289,In_1136);
and U1029 (N_1029,In_710,In_233);
nand U1030 (N_1030,In_1442,In_1132);
nor U1031 (N_1031,In_580,In_164);
and U1032 (N_1032,In_1064,In_171);
or U1033 (N_1033,In_717,In_869);
nand U1034 (N_1034,In_787,In_948);
and U1035 (N_1035,In_57,In_1148);
nand U1036 (N_1036,In_872,In_1166);
or U1037 (N_1037,In_370,In_1164);
or U1038 (N_1038,In_165,In_351);
nand U1039 (N_1039,In_403,In_392);
and U1040 (N_1040,In_775,In_586);
nor U1041 (N_1041,In_1431,In_559);
nor U1042 (N_1042,In_19,In_1474);
and U1043 (N_1043,In_17,In_561);
nor U1044 (N_1044,In_1490,In_1286);
and U1045 (N_1045,In_159,In_543);
nor U1046 (N_1046,In_440,In_663);
nand U1047 (N_1047,In_395,In_1365);
and U1048 (N_1048,In_461,In_900);
or U1049 (N_1049,In_1466,In_1141);
and U1050 (N_1050,In_207,In_716);
or U1051 (N_1051,In_1321,In_749);
or U1052 (N_1052,In_769,In_931);
nor U1053 (N_1053,In_810,In_825);
nor U1054 (N_1054,In_800,In_1295);
nand U1055 (N_1055,In_622,In_924);
nand U1056 (N_1056,In_1071,In_285);
and U1057 (N_1057,In_1444,In_202);
nor U1058 (N_1058,In_859,In_603);
nand U1059 (N_1059,In_342,In_1181);
and U1060 (N_1060,In_818,In_1493);
nor U1061 (N_1061,In_1000,In_227);
or U1062 (N_1062,In_134,In_262);
or U1063 (N_1063,In_266,In_1499);
nand U1064 (N_1064,In_460,In_702);
nand U1065 (N_1065,In_444,In_447);
nand U1066 (N_1066,In_152,In_532);
and U1067 (N_1067,In_316,In_680);
or U1068 (N_1068,In_942,In_580);
and U1069 (N_1069,In_620,In_1179);
and U1070 (N_1070,In_449,In_879);
and U1071 (N_1071,In_1367,In_550);
nor U1072 (N_1072,In_42,In_1372);
and U1073 (N_1073,In_850,In_175);
and U1074 (N_1074,In_1257,In_121);
or U1075 (N_1075,In_72,In_169);
or U1076 (N_1076,In_1134,In_1440);
and U1077 (N_1077,In_242,In_395);
or U1078 (N_1078,In_1285,In_814);
nor U1079 (N_1079,In_1453,In_146);
nand U1080 (N_1080,In_54,In_517);
or U1081 (N_1081,In_1267,In_637);
or U1082 (N_1082,In_306,In_963);
and U1083 (N_1083,In_155,In_1363);
and U1084 (N_1084,In_1063,In_82);
and U1085 (N_1085,In_854,In_1352);
nor U1086 (N_1086,In_1040,In_1094);
and U1087 (N_1087,In_797,In_776);
nand U1088 (N_1088,In_397,In_566);
nor U1089 (N_1089,In_1002,In_1021);
or U1090 (N_1090,In_1049,In_481);
or U1091 (N_1091,In_717,In_218);
nor U1092 (N_1092,In_832,In_1452);
or U1093 (N_1093,In_1197,In_26);
and U1094 (N_1094,In_146,In_45);
or U1095 (N_1095,In_1479,In_1319);
nand U1096 (N_1096,In_1355,In_397);
nor U1097 (N_1097,In_752,In_841);
nand U1098 (N_1098,In_202,In_735);
nor U1099 (N_1099,In_24,In_254);
nand U1100 (N_1100,In_530,In_508);
or U1101 (N_1101,In_652,In_859);
or U1102 (N_1102,In_509,In_571);
or U1103 (N_1103,In_231,In_566);
and U1104 (N_1104,In_1211,In_220);
nand U1105 (N_1105,In_1136,In_1254);
or U1106 (N_1106,In_1054,In_1043);
or U1107 (N_1107,In_1318,In_439);
nand U1108 (N_1108,In_501,In_1315);
or U1109 (N_1109,In_1457,In_1070);
nand U1110 (N_1110,In_966,In_1140);
nor U1111 (N_1111,In_121,In_1043);
and U1112 (N_1112,In_753,In_26);
nor U1113 (N_1113,In_1222,In_1418);
nor U1114 (N_1114,In_1178,In_792);
and U1115 (N_1115,In_857,In_599);
and U1116 (N_1116,In_1115,In_372);
nor U1117 (N_1117,In_416,In_417);
nor U1118 (N_1118,In_131,In_165);
and U1119 (N_1119,In_1197,In_605);
nor U1120 (N_1120,In_806,In_436);
nand U1121 (N_1121,In_669,In_576);
or U1122 (N_1122,In_1487,In_1465);
nor U1123 (N_1123,In_1002,In_877);
or U1124 (N_1124,In_586,In_1466);
or U1125 (N_1125,In_507,In_1432);
or U1126 (N_1126,In_1311,In_1028);
nor U1127 (N_1127,In_682,In_1107);
or U1128 (N_1128,In_259,In_489);
nor U1129 (N_1129,In_930,In_552);
nor U1130 (N_1130,In_1123,In_337);
and U1131 (N_1131,In_1300,In_811);
nand U1132 (N_1132,In_1234,In_1105);
or U1133 (N_1133,In_1078,In_125);
nand U1134 (N_1134,In_860,In_112);
nor U1135 (N_1135,In_884,In_1044);
xnor U1136 (N_1136,In_1176,In_1417);
nor U1137 (N_1137,In_1216,In_973);
nor U1138 (N_1138,In_1076,In_812);
or U1139 (N_1139,In_1040,In_917);
nor U1140 (N_1140,In_973,In_521);
nor U1141 (N_1141,In_93,In_1254);
nor U1142 (N_1142,In_674,In_450);
nor U1143 (N_1143,In_834,In_1012);
nand U1144 (N_1144,In_62,In_765);
or U1145 (N_1145,In_910,In_261);
nand U1146 (N_1146,In_675,In_274);
and U1147 (N_1147,In_1223,In_346);
and U1148 (N_1148,In_1289,In_1047);
or U1149 (N_1149,In_1159,In_1283);
or U1150 (N_1150,In_1456,In_256);
nand U1151 (N_1151,In_236,In_1184);
nand U1152 (N_1152,In_1268,In_1106);
or U1153 (N_1153,In_424,In_1488);
and U1154 (N_1154,In_463,In_1019);
and U1155 (N_1155,In_1225,In_819);
nor U1156 (N_1156,In_289,In_835);
and U1157 (N_1157,In_152,In_142);
and U1158 (N_1158,In_1274,In_323);
and U1159 (N_1159,In_914,In_39);
nor U1160 (N_1160,In_268,In_83);
or U1161 (N_1161,In_1034,In_1153);
nand U1162 (N_1162,In_960,In_445);
nor U1163 (N_1163,In_1401,In_360);
nor U1164 (N_1164,In_706,In_1237);
nand U1165 (N_1165,In_1306,In_1442);
and U1166 (N_1166,In_749,In_1297);
nand U1167 (N_1167,In_430,In_739);
nor U1168 (N_1168,In_279,In_812);
nand U1169 (N_1169,In_394,In_798);
or U1170 (N_1170,In_362,In_1245);
nand U1171 (N_1171,In_349,In_1304);
or U1172 (N_1172,In_1390,In_1313);
nand U1173 (N_1173,In_343,In_259);
xor U1174 (N_1174,In_993,In_126);
nor U1175 (N_1175,In_63,In_1138);
or U1176 (N_1176,In_46,In_672);
nor U1177 (N_1177,In_681,In_145);
nor U1178 (N_1178,In_1276,In_1126);
nand U1179 (N_1179,In_1161,In_592);
or U1180 (N_1180,In_699,In_442);
nor U1181 (N_1181,In_392,In_283);
and U1182 (N_1182,In_979,In_1260);
and U1183 (N_1183,In_1144,In_1108);
nand U1184 (N_1184,In_850,In_427);
nand U1185 (N_1185,In_540,In_1068);
nor U1186 (N_1186,In_342,In_1082);
nor U1187 (N_1187,In_1244,In_977);
nand U1188 (N_1188,In_390,In_232);
nor U1189 (N_1189,In_700,In_513);
and U1190 (N_1190,In_657,In_348);
xor U1191 (N_1191,In_1191,In_971);
nor U1192 (N_1192,In_22,In_566);
or U1193 (N_1193,In_225,In_527);
or U1194 (N_1194,In_979,In_539);
nand U1195 (N_1195,In_363,In_1283);
and U1196 (N_1196,In_1480,In_842);
or U1197 (N_1197,In_325,In_122);
and U1198 (N_1198,In_586,In_251);
or U1199 (N_1199,In_884,In_1052);
nor U1200 (N_1200,In_930,In_820);
or U1201 (N_1201,In_890,In_863);
nand U1202 (N_1202,In_187,In_1058);
nand U1203 (N_1203,In_705,In_1304);
nor U1204 (N_1204,In_550,In_1323);
nor U1205 (N_1205,In_247,In_162);
nand U1206 (N_1206,In_916,In_852);
nor U1207 (N_1207,In_834,In_804);
nor U1208 (N_1208,In_1323,In_951);
nor U1209 (N_1209,In_748,In_1199);
or U1210 (N_1210,In_1245,In_247);
and U1211 (N_1211,In_469,In_384);
or U1212 (N_1212,In_1381,In_856);
nor U1213 (N_1213,In_1030,In_694);
nor U1214 (N_1214,In_345,In_343);
or U1215 (N_1215,In_447,In_487);
nor U1216 (N_1216,In_427,In_843);
and U1217 (N_1217,In_363,In_1359);
and U1218 (N_1218,In_864,In_1215);
and U1219 (N_1219,In_233,In_662);
nor U1220 (N_1220,In_1045,In_756);
or U1221 (N_1221,In_570,In_257);
or U1222 (N_1222,In_1382,In_293);
nand U1223 (N_1223,In_1393,In_260);
xnor U1224 (N_1224,In_837,In_1306);
or U1225 (N_1225,In_938,In_618);
or U1226 (N_1226,In_832,In_397);
nand U1227 (N_1227,In_853,In_1200);
nor U1228 (N_1228,In_497,In_1479);
nand U1229 (N_1229,In_1400,In_1487);
or U1230 (N_1230,In_184,In_1354);
or U1231 (N_1231,In_908,In_268);
and U1232 (N_1232,In_305,In_1055);
or U1233 (N_1233,In_317,In_265);
or U1234 (N_1234,In_64,In_321);
or U1235 (N_1235,In_905,In_835);
nor U1236 (N_1236,In_225,In_678);
nor U1237 (N_1237,In_892,In_80);
nand U1238 (N_1238,In_831,In_243);
or U1239 (N_1239,In_1222,In_784);
nand U1240 (N_1240,In_93,In_658);
nand U1241 (N_1241,In_589,In_1365);
nor U1242 (N_1242,In_27,In_700);
nand U1243 (N_1243,In_876,In_1061);
nor U1244 (N_1244,In_1227,In_683);
nor U1245 (N_1245,In_451,In_81);
nand U1246 (N_1246,In_74,In_1461);
or U1247 (N_1247,In_1196,In_646);
and U1248 (N_1248,In_468,In_1431);
and U1249 (N_1249,In_1009,In_72);
or U1250 (N_1250,In_699,In_1154);
nand U1251 (N_1251,In_59,In_466);
or U1252 (N_1252,In_913,In_1188);
and U1253 (N_1253,In_1344,In_629);
nand U1254 (N_1254,In_1285,In_417);
or U1255 (N_1255,In_500,In_404);
or U1256 (N_1256,In_997,In_518);
and U1257 (N_1257,In_844,In_1392);
nor U1258 (N_1258,In_192,In_1191);
and U1259 (N_1259,In_718,In_372);
and U1260 (N_1260,In_126,In_253);
nor U1261 (N_1261,In_732,In_1017);
nor U1262 (N_1262,In_1126,In_985);
and U1263 (N_1263,In_367,In_1237);
or U1264 (N_1264,In_306,In_1108);
nand U1265 (N_1265,In_1330,In_926);
nand U1266 (N_1266,In_288,In_1037);
and U1267 (N_1267,In_1253,In_724);
nor U1268 (N_1268,In_1437,In_526);
or U1269 (N_1269,In_690,In_411);
nand U1270 (N_1270,In_43,In_425);
nor U1271 (N_1271,In_446,In_1082);
nand U1272 (N_1272,In_443,In_1080);
nor U1273 (N_1273,In_553,In_1486);
nor U1274 (N_1274,In_774,In_805);
and U1275 (N_1275,In_483,In_723);
or U1276 (N_1276,In_1371,In_161);
and U1277 (N_1277,In_364,In_690);
and U1278 (N_1278,In_232,In_613);
and U1279 (N_1279,In_1280,In_419);
nand U1280 (N_1280,In_132,In_732);
nor U1281 (N_1281,In_492,In_87);
and U1282 (N_1282,In_1377,In_1139);
nand U1283 (N_1283,In_728,In_895);
and U1284 (N_1284,In_51,In_199);
or U1285 (N_1285,In_0,In_614);
nor U1286 (N_1286,In_481,In_1191);
nor U1287 (N_1287,In_720,In_162);
nand U1288 (N_1288,In_903,In_408);
nor U1289 (N_1289,In_626,In_1285);
and U1290 (N_1290,In_979,In_1068);
or U1291 (N_1291,In_482,In_1171);
nor U1292 (N_1292,In_31,In_1033);
xor U1293 (N_1293,In_76,In_51);
nand U1294 (N_1294,In_1233,In_870);
or U1295 (N_1295,In_536,In_901);
or U1296 (N_1296,In_808,In_834);
or U1297 (N_1297,In_1380,In_94);
nand U1298 (N_1298,In_1138,In_337);
nand U1299 (N_1299,In_897,In_1232);
nor U1300 (N_1300,In_1171,In_1424);
xnor U1301 (N_1301,In_1012,In_385);
or U1302 (N_1302,In_346,In_1406);
or U1303 (N_1303,In_1218,In_1450);
and U1304 (N_1304,In_546,In_360);
or U1305 (N_1305,In_1488,In_1059);
nor U1306 (N_1306,In_438,In_828);
nor U1307 (N_1307,In_818,In_1173);
and U1308 (N_1308,In_190,In_900);
and U1309 (N_1309,In_392,In_1066);
and U1310 (N_1310,In_1308,In_1276);
or U1311 (N_1311,In_404,In_379);
or U1312 (N_1312,In_134,In_718);
or U1313 (N_1313,In_71,In_817);
nand U1314 (N_1314,In_1001,In_687);
nor U1315 (N_1315,In_1302,In_1057);
and U1316 (N_1316,In_1439,In_630);
nand U1317 (N_1317,In_72,In_1278);
nand U1318 (N_1318,In_869,In_418);
and U1319 (N_1319,In_833,In_548);
nor U1320 (N_1320,In_405,In_1099);
or U1321 (N_1321,In_995,In_638);
and U1322 (N_1322,In_886,In_1420);
nor U1323 (N_1323,In_154,In_299);
or U1324 (N_1324,In_1126,In_525);
nand U1325 (N_1325,In_1118,In_236);
and U1326 (N_1326,In_708,In_268);
or U1327 (N_1327,In_580,In_1246);
and U1328 (N_1328,In_555,In_8);
or U1329 (N_1329,In_852,In_483);
xor U1330 (N_1330,In_648,In_149);
nor U1331 (N_1331,In_544,In_697);
and U1332 (N_1332,In_780,In_1362);
or U1333 (N_1333,In_836,In_926);
and U1334 (N_1334,In_2,In_842);
or U1335 (N_1335,In_1474,In_1264);
nor U1336 (N_1336,In_882,In_1149);
nor U1337 (N_1337,In_794,In_757);
or U1338 (N_1338,In_1050,In_857);
nor U1339 (N_1339,In_567,In_1401);
or U1340 (N_1340,In_1400,In_359);
nor U1341 (N_1341,In_1082,In_617);
and U1342 (N_1342,In_342,In_1419);
or U1343 (N_1343,In_1435,In_710);
or U1344 (N_1344,In_166,In_1351);
nor U1345 (N_1345,In_1118,In_562);
nand U1346 (N_1346,In_1436,In_329);
and U1347 (N_1347,In_696,In_359);
nand U1348 (N_1348,In_179,In_767);
nor U1349 (N_1349,In_1007,In_999);
or U1350 (N_1350,In_461,In_422);
nand U1351 (N_1351,In_1072,In_1147);
and U1352 (N_1352,In_133,In_773);
nor U1353 (N_1353,In_244,In_1172);
xnor U1354 (N_1354,In_687,In_1420);
nand U1355 (N_1355,In_840,In_834);
nand U1356 (N_1356,In_579,In_1291);
nand U1357 (N_1357,In_1014,In_561);
and U1358 (N_1358,In_1020,In_1308);
nor U1359 (N_1359,In_637,In_678);
or U1360 (N_1360,In_459,In_850);
and U1361 (N_1361,In_310,In_292);
and U1362 (N_1362,In_617,In_1040);
and U1363 (N_1363,In_658,In_486);
or U1364 (N_1364,In_1407,In_1122);
or U1365 (N_1365,In_1105,In_598);
nor U1366 (N_1366,In_1458,In_1289);
nor U1367 (N_1367,In_692,In_637);
nor U1368 (N_1368,In_387,In_317);
nand U1369 (N_1369,In_447,In_636);
nor U1370 (N_1370,In_770,In_445);
nor U1371 (N_1371,In_419,In_352);
and U1372 (N_1372,In_8,In_981);
nand U1373 (N_1373,In_752,In_263);
nand U1374 (N_1374,In_300,In_725);
and U1375 (N_1375,In_353,In_444);
nor U1376 (N_1376,In_137,In_1174);
or U1377 (N_1377,In_122,In_601);
nand U1378 (N_1378,In_762,In_460);
nand U1379 (N_1379,In_143,In_837);
nor U1380 (N_1380,In_779,In_727);
or U1381 (N_1381,In_477,In_971);
nor U1382 (N_1382,In_329,In_14);
and U1383 (N_1383,In_1028,In_549);
nor U1384 (N_1384,In_568,In_75);
or U1385 (N_1385,In_180,In_1386);
nor U1386 (N_1386,In_118,In_687);
xnor U1387 (N_1387,In_961,In_574);
nor U1388 (N_1388,In_335,In_207);
nor U1389 (N_1389,In_1022,In_330);
or U1390 (N_1390,In_1105,In_90);
nand U1391 (N_1391,In_1118,In_1190);
and U1392 (N_1392,In_364,In_839);
nor U1393 (N_1393,In_648,In_1225);
or U1394 (N_1394,In_1474,In_519);
or U1395 (N_1395,In_1465,In_870);
and U1396 (N_1396,In_931,In_814);
or U1397 (N_1397,In_823,In_844);
nand U1398 (N_1398,In_227,In_339);
and U1399 (N_1399,In_1174,In_1403);
or U1400 (N_1400,In_446,In_219);
nand U1401 (N_1401,In_910,In_680);
nor U1402 (N_1402,In_1380,In_111);
and U1403 (N_1403,In_1376,In_1088);
nor U1404 (N_1404,In_1238,In_1152);
or U1405 (N_1405,In_682,In_419);
or U1406 (N_1406,In_25,In_20);
and U1407 (N_1407,In_40,In_1116);
nand U1408 (N_1408,In_1444,In_867);
nand U1409 (N_1409,In_1011,In_501);
nor U1410 (N_1410,In_495,In_249);
nor U1411 (N_1411,In_638,In_409);
nand U1412 (N_1412,In_980,In_257);
or U1413 (N_1413,In_497,In_647);
nor U1414 (N_1414,In_1393,In_198);
or U1415 (N_1415,In_634,In_443);
nand U1416 (N_1416,In_917,In_834);
and U1417 (N_1417,In_737,In_903);
nand U1418 (N_1418,In_1450,In_229);
or U1419 (N_1419,In_10,In_1364);
nand U1420 (N_1420,In_1091,In_772);
or U1421 (N_1421,In_490,In_664);
or U1422 (N_1422,In_1045,In_856);
nor U1423 (N_1423,In_1320,In_544);
nand U1424 (N_1424,In_717,In_1462);
nor U1425 (N_1425,In_901,In_1308);
nor U1426 (N_1426,In_1393,In_399);
or U1427 (N_1427,In_51,In_1484);
and U1428 (N_1428,In_454,In_556);
or U1429 (N_1429,In_1,In_680);
or U1430 (N_1430,In_805,In_856);
or U1431 (N_1431,In_482,In_879);
and U1432 (N_1432,In_406,In_819);
or U1433 (N_1433,In_481,In_1239);
nor U1434 (N_1434,In_1280,In_261);
and U1435 (N_1435,In_998,In_544);
and U1436 (N_1436,In_319,In_378);
and U1437 (N_1437,In_462,In_56);
nor U1438 (N_1438,In_377,In_1019);
nor U1439 (N_1439,In_1440,In_160);
nor U1440 (N_1440,In_1117,In_1399);
or U1441 (N_1441,In_22,In_1381);
and U1442 (N_1442,In_1327,In_1343);
nor U1443 (N_1443,In_1487,In_478);
nor U1444 (N_1444,In_433,In_718);
nand U1445 (N_1445,In_157,In_228);
and U1446 (N_1446,In_1267,In_153);
and U1447 (N_1447,In_1366,In_1131);
nor U1448 (N_1448,In_1048,In_28);
nor U1449 (N_1449,In_124,In_1063);
nor U1450 (N_1450,In_916,In_1358);
xor U1451 (N_1451,In_161,In_1307);
nor U1452 (N_1452,In_1402,In_745);
nor U1453 (N_1453,In_1488,In_615);
nand U1454 (N_1454,In_551,In_1057);
nor U1455 (N_1455,In_363,In_375);
nand U1456 (N_1456,In_1259,In_643);
nor U1457 (N_1457,In_804,In_850);
or U1458 (N_1458,In_11,In_162);
nand U1459 (N_1459,In_1347,In_706);
nand U1460 (N_1460,In_702,In_836);
nand U1461 (N_1461,In_22,In_1461);
or U1462 (N_1462,In_1206,In_962);
or U1463 (N_1463,In_1091,In_45);
and U1464 (N_1464,In_1043,In_1495);
nor U1465 (N_1465,In_694,In_49);
nor U1466 (N_1466,In_1078,In_596);
or U1467 (N_1467,In_1478,In_766);
nand U1468 (N_1468,In_536,In_348);
and U1469 (N_1469,In_1421,In_659);
or U1470 (N_1470,In_83,In_462);
nand U1471 (N_1471,In_1378,In_1308);
nor U1472 (N_1472,In_888,In_234);
and U1473 (N_1473,In_1216,In_1030);
nor U1474 (N_1474,In_851,In_994);
nand U1475 (N_1475,In_799,In_708);
and U1476 (N_1476,In_144,In_995);
nand U1477 (N_1477,In_1272,In_124);
xor U1478 (N_1478,In_957,In_508);
nor U1479 (N_1479,In_900,In_801);
or U1480 (N_1480,In_31,In_607);
nand U1481 (N_1481,In_418,In_38);
nand U1482 (N_1482,In_1410,In_192);
nand U1483 (N_1483,In_69,In_1494);
and U1484 (N_1484,In_959,In_723);
and U1485 (N_1485,In_731,In_647);
nand U1486 (N_1486,In_1306,In_1070);
nand U1487 (N_1487,In_971,In_1477);
nand U1488 (N_1488,In_482,In_991);
and U1489 (N_1489,In_659,In_10);
and U1490 (N_1490,In_1082,In_252);
nor U1491 (N_1491,In_1110,In_93);
and U1492 (N_1492,In_1280,In_1370);
xor U1493 (N_1493,In_813,In_946);
nor U1494 (N_1494,In_576,In_286);
nor U1495 (N_1495,In_412,In_894);
and U1496 (N_1496,In_404,In_1262);
and U1497 (N_1497,In_482,In_113);
nor U1498 (N_1498,In_165,In_867);
or U1499 (N_1499,In_279,In_1116);
and U1500 (N_1500,In_1127,In_1049);
nand U1501 (N_1501,In_1426,In_806);
nand U1502 (N_1502,In_904,In_819);
nor U1503 (N_1503,In_1412,In_961);
nand U1504 (N_1504,In_818,In_202);
nor U1505 (N_1505,In_530,In_481);
and U1506 (N_1506,In_466,In_89);
nor U1507 (N_1507,In_468,In_952);
nor U1508 (N_1508,In_67,In_1210);
xnor U1509 (N_1509,In_716,In_1229);
nand U1510 (N_1510,In_80,In_538);
or U1511 (N_1511,In_578,In_465);
nand U1512 (N_1512,In_667,In_791);
nor U1513 (N_1513,In_1329,In_566);
and U1514 (N_1514,In_305,In_542);
and U1515 (N_1515,In_637,In_665);
nand U1516 (N_1516,In_41,In_261);
or U1517 (N_1517,In_1359,In_711);
or U1518 (N_1518,In_1038,In_517);
nand U1519 (N_1519,In_1449,In_995);
or U1520 (N_1520,In_764,In_335);
and U1521 (N_1521,In_360,In_1040);
nor U1522 (N_1522,In_393,In_1014);
nand U1523 (N_1523,In_1338,In_557);
nor U1524 (N_1524,In_553,In_975);
or U1525 (N_1525,In_1225,In_1328);
nor U1526 (N_1526,In_1085,In_1386);
nand U1527 (N_1527,In_1399,In_585);
nor U1528 (N_1528,In_572,In_449);
nor U1529 (N_1529,In_554,In_889);
or U1530 (N_1530,In_966,In_1113);
and U1531 (N_1531,In_137,In_1439);
nor U1532 (N_1532,In_1183,In_1166);
and U1533 (N_1533,In_1286,In_1096);
nor U1534 (N_1534,In_1349,In_1318);
nor U1535 (N_1535,In_943,In_1333);
and U1536 (N_1536,In_276,In_1337);
nand U1537 (N_1537,In_173,In_491);
nor U1538 (N_1538,In_93,In_1207);
nor U1539 (N_1539,In_1157,In_1235);
nor U1540 (N_1540,In_1329,In_414);
or U1541 (N_1541,In_1419,In_923);
and U1542 (N_1542,In_962,In_237);
or U1543 (N_1543,In_1415,In_1020);
nand U1544 (N_1544,In_292,In_860);
or U1545 (N_1545,In_162,In_1099);
and U1546 (N_1546,In_234,In_1492);
nand U1547 (N_1547,In_1304,In_454);
nand U1548 (N_1548,In_718,In_117);
nor U1549 (N_1549,In_430,In_1136);
nand U1550 (N_1550,In_606,In_1174);
nand U1551 (N_1551,In_1101,In_495);
or U1552 (N_1552,In_164,In_553);
or U1553 (N_1553,In_492,In_524);
or U1554 (N_1554,In_1053,In_804);
or U1555 (N_1555,In_103,In_1384);
nand U1556 (N_1556,In_678,In_56);
nand U1557 (N_1557,In_299,In_313);
and U1558 (N_1558,In_433,In_899);
nor U1559 (N_1559,In_1272,In_704);
nand U1560 (N_1560,In_1013,In_596);
nand U1561 (N_1561,In_109,In_1400);
nand U1562 (N_1562,In_932,In_1147);
nor U1563 (N_1563,In_1427,In_1360);
or U1564 (N_1564,In_465,In_921);
and U1565 (N_1565,In_61,In_1289);
nand U1566 (N_1566,In_1496,In_1195);
nor U1567 (N_1567,In_1161,In_272);
or U1568 (N_1568,In_853,In_159);
nor U1569 (N_1569,In_565,In_978);
or U1570 (N_1570,In_977,In_954);
nor U1571 (N_1571,In_920,In_256);
nor U1572 (N_1572,In_500,In_718);
or U1573 (N_1573,In_189,In_1478);
nor U1574 (N_1574,In_890,In_915);
nor U1575 (N_1575,In_438,In_657);
and U1576 (N_1576,In_1461,In_767);
nand U1577 (N_1577,In_786,In_1484);
nor U1578 (N_1578,In_1050,In_1013);
and U1579 (N_1579,In_1263,In_1227);
xnor U1580 (N_1580,In_102,In_880);
nor U1581 (N_1581,In_1428,In_1216);
and U1582 (N_1582,In_1027,In_84);
and U1583 (N_1583,In_961,In_104);
nor U1584 (N_1584,In_1470,In_935);
nor U1585 (N_1585,In_892,In_1256);
and U1586 (N_1586,In_924,In_316);
nand U1587 (N_1587,In_1499,In_1465);
and U1588 (N_1588,In_771,In_949);
nand U1589 (N_1589,In_25,In_583);
nand U1590 (N_1590,In_928,In_873);
or U1591 (N_1591,In_577,In_592);
nand U1592 (N_1592,In_1295,In_346);
or U1593 (N_1593,In_160,In_372);
or U1594 (N_1594,In_1483,In_48);
or U1595 (N_1595,In_699,In_779);
nor U1596 (N_1596,In_417,In_57);
and U1597 (N_1597,In_1426,In_91);
or U1598 (N_1598,In_343,In_1147);
or U1599 (N_1599,In_570,In_996);
nand U1600 (N_1600,In_1087,In_725);
nor U1601 (N_1601,In_57,In_1156);
nor U1602 (N_1602,In_270,In_1482);
and U1603 (N_1603,In_290,In_528);
and U1604 (N_1604,In_1224,In_1139);
nand U1605 (N_1605,In_1237,In_1232);
or U1606 (N_1606,In_176,In_270);
or U1607 (N_1607,In_1381,In_956);
or U1608 (N_1608,In_882,In_584);
nor U1609 (N_1609,In_47,In_16);
and U1610 (N_1610,In_1247,In_890);
or U1611 (N_1611,In_1453,In_1115);
and U1612 (N_1612,In_284,In_1233);
nor U1613 (N_1613,In_779,In_208);
or U1614 (N_1614,In_552,In_1468);
nand U1615 (N_1615,In_640,In_108);
nand U1616 (N_1616,In_1466,In_1385);
and U1617 (N_1617,In_1027,In_324);
or U1618 (N_1618,In_799,In_1014);
and U1619 (N_1619,In_755,In_933);
nand U1620 (N_1620,In_885,In_127);
nand U1621 (N_1621,In_922,In_1303);
or U1622 (N_1622,In_820,In_585);
and U1623 (N_1623,In_1432,In_589);
or U1624 (N_1624,In_874,In_906);
nor U1625 (N_1625,In_937,In_183);
nor U1626 (N_1626,In_1326,In_1052);
or U1627 (N_1627,In_812,In_1137);
and U1628 (N_1628,In_927,In_250);
nand U1629 (N_1629,In_1414,In_783);
nor U1630 (N_1630,In_221,In_1157);
or U1631 (N_1631,In_882,In_1447);
nor U1632 (N_1632,In_161,In_443);
nand U1633 (N_1633,In_1210,In_283);
nor U1634 (N_1634,In_220,In_1296);
or U1635 (N_1635,In_636,In_237);
or U1636 (N_1636,In_1466,In_629);
or U1637 (N_1637,In_430,In_154);
and U1638 (N_1638,In_270,In_1260);
and U1639 (N_1639,In_297,In_695);
or U1640 (N_1640,In_1271,In_86);
or U1641 (N_1641,In_965,In_1416);
nand U1642 (N_1642,In_1489,In_1122);
nor U1643 (N_1643,In_138,In_624);
or U1644 (N_1644,In_658,In_1193);
nand U1645 (N_1645,In_771,In_446);
and U1646 (N_1646,In_1421,In_393);
nor U1647 (N_1647,In_42,In_513);
or U1648 (N_1648,In_874,In_143);
or U1649 (N_1649,In_18,In_615);
or U1650 (N_1650,In_453,In_522);
or U1651 (N_1651,In_308,In_405);
and U1652 (N_1652,In_1156,In_556);
nor U1653 (N_1653,In_104,In_797);
or U1654 (N_1654,In_580,In_1427);
nand U1655 (N_1655,In_1456,In_648);
nor U1656 (N_1656,In_1232,In_1385);
and U1657 (N_1657,In_506,In_155);
nor U1658 (N_1658,In_1035,In_623);
nor U1659 (N_1659,In_1112,In_1286);
and U1660 (N_1660,In_137,In_919);
or U1661 (N_1661,In_303,In_1398);
or U1662 (N_1662,In_1466,In_513);
nor U1663 (N_1663,In_1177,In_903);
nand U1664 (N_1664,In_1439,In_10);
nor U1665 (N_1665,In_990,In_1147);
nand U1666 (N_1666,In_495,In_714);
or U1667 (N_1667,In_1436,In_186);
nand U1668 (N_1668,In_292,In_1123);
nand U1669 (N_1669,In_337,In_854);
or U1670 (N_1670,In_1306,In_1086);
and U1671 (N_1671,In_1461,In_16);
nand U1672 (N_1672,In_1439,In_434);
nor U1673 (N_1673,In_1480,In_1086);
nor U1674 (N_1674,In_84,In_1013);
or U1675 (N_1675,In_501,In_427);
nor U1676 (N_1676,In_1078,In_1356);
nor U1677 (N_1677,In_1409,In_713);
or U1678 (N_1678,In_1020,In_675);
xnor U1679 (N_1679,In_663,In_1431);
or U1680 (N_1680,In_1086,In_419);
or U1681 (N_1681,In_38,In_455);
and U1682 (N_1682,In_183,In_43);
or U1683 (N_1683,In_248,In_1433);
and U1684 (N_1684,In_604,In_270);
and U1685 (N_1685,In_1297,In_1111);
nand U1686 (N_1686,In_943,In_1130);
nand U1687 (N_1687,In_248,In_660);
nand U1688 (N_1688,In_14,In_1320);
nand U1689 (N_1689,In_312,In_25);
and U1690 (N_1690,In_1062,In_465);
or U1691 (N_1691,In_20,In_807);
and U1692 (N_1692,In_471,In_975);
and U1693 (N_1693,In_1211,In_1021);
and U1694 (N_1694,In_1166,In_1333);
and U1695 (N_1695,In_1239,In_1224);
and U1696 (N_1696,In_881,In_820);
nor U1697 (N_1697,In_102,In_861);
or U1698 (N_1698,In_1398,In_531);
nand U1699 (N_1699,In_606,In_627);
nor U1700 (N_1700,In_742,In_509);
nand U1701 (N_1701,In_854,In_1393);
or U1702 (N_1702,In_1200,In_38);
and U1703 (N_1703,In_1363,In_132);
and U1704 (N_1704,In_221,In_490);
nor U1705 (N_1705,In_636,In_1475);
nand U1706 (N_1706,In_977,In_1006);
and U1707 (N_1707,In_1293,In_526);
or U1708 (N_1708,In_44,In_366);
nand U1709 (N_1709,In_1389,In_6);
and U1710 (N_1710,In_598,In_707);
and U1711 (N_1711,In_716,In_322);
nand U1712 (N_1712,In_518,In_111);
or U1713 (N_1713,In_1333,In_1180);
nor U1714 (N_1714,In_505,In_651);
nand U1715 (N_1715,In_894,In_1069);
nor U1716 (N_1716,In_622,In_453);
nor U1717 (N_1717,In_1174,In_791);
and U1718 (N_1718,In_1219,In_1455);
and U1719 (N_1719,In_1346,In_1317);
and U1720 (N_1720,In_339,In_994);
nand U1721 (N_1721,In_1426,In_255);
and U1722 (N_1722,In_852,In_552);
or U1723 (N_1723,In_689,In_325);
xnor U1724 (N_1724,In_1452,In_213);
or U1725 (N_1725,In_1365,In_974);
or U1726 (N_1726,In_43,In_726);
or U1727 (N_1727,In_950,In_695);
or U1728 (N_1728,In_41,In_462);
nor U1729 (N_1729,In_391,In_676);
nor U1730 (N_1730,In_950,In_1244);
or U1731 (N_1731,In_2,In_1030);
or U1732 (N_1732,In_597,In_1420);
or U1733 (N_1733,In_272,In_636);
and U1734 (N_1734,In_649,In_1490);
nand U1735 (N_1735,In_454,In_1215);
nor U1736 (N_1736,In_1040,In_320);
nor U1737 (N_1737,In_1465,In_997);
or U1738 (N_1738,In_1352,In_43);
nand U1739 (N_1739,In_1186,In_1452);
and U1740 (N_1740,In_127,In_1330);
or U1741 (N_1741,In_1229,In_345);
and U1742 (N_1742,In_1430,In_1105);
or U1743 (N_1743,In_41,In_966);
and U1744 (N_1744,In_678,In_71);
nand U1745 (N_1745,In_1227,In_28);
nand U1746 (N_1746,In_957,In_32);
and U1747 (N_1747,In_1076,In_976);
nor U1748 (N_1748,In_642,In_872);
or U1749 (N_1749,In_433,In_890);
nand U1750 (N_1750,In_162,In_76);
and U1751 (N_1751,In_1182,In_800);
or U1752 (N_1752,In_1095,In_1282);
or U1753 (N_1753,In_747,In_902);
and U1754 (N_1754,In_207,In_1113);
nor U1755 (N_1755,In_86,In_965);
or U1756 (N_1756,In_1106,In_936);
nor U1757 (N_1757,In_177,In_308);
or U1758 (N_1758,In_272,In_389);
or U1759 (N_1759,In_673,In_534);
nor U1760 (N_1760,In_206,In_1015);
or U1761 (N_1761,In_740,In_1236);
or U1762 (N_1762,In_800,In_963);
nand U1763 (N_1763,In_1363,In_1489);
or U1764 (N_1764,In_722,In_1271);
nand U1765 (N_1765,In_394,In_372);
or U1766 (N_1766,In_640,In_476);
nor U1767 (N_1767,In_521,In_305);
nand U1768 (N_1768,In_1379,In_169);
and U1769 (N_1769,In_1414,In_551);
or U1770 (N_1770,In_1053,In_1432);
nor U1771 (N_1771,In_732,In_467);
nor U1772 (N_1772,In_752,In_1077);
nand U1773 (N_1773,In_1052,In_161);
nand U1774 (N_1774,In_135,In_754);
nand U1775 (N_1775,In_292,In_1367);
nor U1776 (N_1776,In_1315,In_955);
nand U1777 (N_1777,In_721,In_1212);
nand U1778 (N_1778,In_340,In_14);
and U1779 (N_1779,In_1379,In_1151);
nand U1780 (N_1780,In_1334,In_1416);
or U1781 (N_1781,In_187,In_508);
or U1782 (N_1782,In_522,In_1048);
nor U1783 (N_1783,In_1203,In_741);
nor U1784 (N_1784,In_1364,In_189);
nor U1785 (N_1785,In_559,In_546);
and U1786 (N_1786,In_1044,In_1138);
or U1787 (N_1787,In_613,In_685);
and U1788 (N_1788,In_750,In_636);
or U1789 (N_1789,In_269,In_661);
or U1790 (N_1790,In_710,In_262);
nor U1791 (N_1791,In_611,In_1285);
nand U1792 (N_1792,In_1019,In_1062);
nand U1793 (N_1793,In_1303,In_1291);
nor U1794 (N_1794,In_1350,In_383);
or U1795 (N_1795,In_1,In_775);
or U1796 (N_1796,In_1393,In_667);
and U1797 (N_1797,In_439,In_844);
or U1798 (N_1798,In_445,In_475);
nor U1799 (N_1799,In_1271,In_1068);
or U1800 (N_1800,In_1348,In_1252);
nand U1801 (N_1801,In_1413,In_177);
nand U1802 (N_1802,In_40,In_134);
nor U1803 (N_1803,In_1094,In_618);
or U1804 (N_1804,In_1499,In_1462);
nand U1805 (N_1805,In_793,In_19);
nand U1806 (N_1806,In_400,In_1451);
nor U1807 (N_1807,In_963,In_510);
xor U1808 (N_1808,In_774,In_1297);
or U1809 (N_1809,In_1291,In_1281);
and U1810 (N_1810,In_423,In_237);
nand U1811 (N_1811,In_478,In_1421);
nand U1812 (N_1812,In_338,In_534);
nor U1813 (N_1813,In_272,In_1331);
nand U1814 (N_1814,In_1219,In_327);
nand U1815 (N_1815,In_703,In_523);
or U1816 (N_1816,In_738,In_823);
nor U1817 (N_1817,In_712,In_1128);
or U1818 (N_1818,In_1192,In_1333);
nand U1819 (N_1819,In_342,In_1281);
nand U1820 (N_1820,In_686,In_996);
or U1821 (N_1821,In_1323,In_1247);
nor U1822 (N_1822,In_315,In_915);
nand U1823 (N_1823,In_472,In_796);
nor U1824 (N_1824,In_625,In_1119);
nor U1825 (N_1825,In_483,In_70);
nor U1826 (N_1826,In_664,In_520);
and U1827 (N_1827,In_764,In_221);
and U1828 (N_1828,In_215,In_604);
nand U1829 (N_1829,In_1306,In_154);
nor U1830 (N_1830,In_508,In_305);
nand U1831 (N_1831,In_752,In_233);
or U1832 (N_1832,In_292,In_637);
or U1833 (N_1833,In_960,In_1457);
and U1834 (N_1834,In_1207,In_228);
nand U1835 (N_1835,In_587,In_543);
nand U1836 (N_1836,In_1039,In_44);
nor U1837 (N_1837,In_1191,In_1078);
nand U1838 (N_1838,In_1260,In_372);
nand U1839 (N_1839,In_1001,In_316);
or U1840 (N_1840,In_1191,In_823);
nor U1841 (N_1841,In_396,In_1098);
nand U1842 (N_1842,In_1022,In_198);
nor U1843 (N_1843,In_849,In_1184);
and U1844 (N_1844,In_939,In_0);
nor U1845 (N_1845,In_733,In_1136);
nor U1846 (N_1846,In_722,In_586);
and U1847 (N_1847,In_43,In_1354);
nor U1848 (N_1848,In_9,In_229);
nor U1849 (N_1849,In_1450,In_945);
and U1850 (N_1850,In_1220,In_1074);
and U1851 (N_1851,In_142,In_50);
and U1852 (N_1852,In_1211,In_721);
nand U1853 (N_1853,In_404,In_1306);
or U1854 (N_1854,In_102,In_269);
nand U1855 (N_1855,In_1371,In_409);
nand U1856 (N_1856,In_1088,In_1320);
and U1857 (N_1857,In_540,In_1263);
and U1858 (N_1858,In_465,In_32);
nor U1859 (N_1859,In_1312,In_1000);
and U1860 (N_1860,In_1261,In_1351);
nor U1861 (N_1861,In_456,In_662);
and U1862 (N_1862,In_92,In_1100);
nor U1863 (N_1863,In_333,In_292);
or U1864 (N_1864,In_548,In_867);
and U1865 (N_1865,In_694,In_1009);
nand U1866 (N_1866,In_1492,In_1077);
or U1867 (N_1867,In_12,In_685);
nand U1868 (N_1868,In_767,In_753);
and U1869 (N_1869,In_371,In_929);
and U1870 (N_1870,In_1306,In_158);
or U1871 (N_1871,In_13,In_953);
or U1872 (N_1872,In_802,In_168);
or U1873 (N_1873,In_704,In_1170);
and U1874 (N_1874,In_1088,In_361);
or U1875 (N_1875,In_359,In_841);
nand U1876 (N_1876,In_695,In_1429);
nand U1877 (N_1877,In_1449,In_997);
nand U1878 (N_1878,In_1467,In_820);
or U1879 (N_1879,In_812,In_876);
nor U1880 (N_1880,In_202,In_1045);
nand U1881 (N_1881,In_867,In_231);
nor U1882 (N_1882,In_1090,In_196);
xor U1883 (N_1883,In_178,In_1023);
nor U1884 (N_1884,In_279,In_1382);
and U1885 (N_1885,In_908,In_66);
or U1886 (N_1886,In_797,In_1289);
or U1887 (N_1887,In_1462,In_955);
or U1888 (N_1888,In_754,In_554);
or U1889 (N_1889,In_825,In_578);
or U1890 (N_1890,In_913,In_1366);
nand U1891 (N_1891,In_937,In_384);
nor U1892 (N_1892,In_1450,In_352);
or U1893 (N_1893,In_958,In_441);
nor U1894 (N_1894,In_426,In_1154);
and U1895 (N_1895,In_1388,In_1287);
nor U1896 (N_1896,In_161,In_60);
nand U1897 (N_1897,In_964,In_1315);
nor U1898 (N_1898,In_1105,In_948);
nor U1899 (N_1899,In_1041,In_648);
nand U1900 (N_1900,In_322,In_482);
nor U1901 (N_1901,In_329,In_1485);
nor U1902 (N_1902,In_470,In_432);
nor U1903 (N_1903,In_358,In_115);
nor U1904 (N_1904,In_84,In_1394);
nor U1905 (N_1905,In_526,In_863);
nor U1906 (N_1906,In_745,In_264);
nand U1907 (N_1907,In_891,In_547);
nand U1908 (N_1908,In_562,In_809);
or U1909 (N_1909,In_835,In_280);
or U1910 (N_1910,In_518,In_1286);
nor U1911 (N_1911,In_401,In_587);
and U1912 (N_1912,In_1152,In_86);
nor U1913 (N_1913,In_125,In_1246);
nand U1914 (N_1914,In_1281,In_996);
nor U1915 (N_1915,In_1153,In_1094);
and U1916 (N_1916,In_900,In_771);
or U1917 (N_1917,In_1295,In_881);
nand U1918 (N_1918,In_1245,In_938);
nor U1919 (N_1919,In_204,In_1188);
nor U1920 (N_1920,In_787,In_1141);
or U1921 (N_1921,In_1225,In_786);
or U1922 (N_1922,In_720,In_296);
nor U1923 (N_1923,In_592,In_1150);
or U1924 (N_1924,In_1110,In_1424);
nand U1925 (N_1925,In_734,In_533);
nand U1926 (N_1926,In_903,In_9);
nor U1927 (N_1927,In_961,In_11);
nor U1928 (N_1928,In_660,In_161);
nor U1929 (N_1929,In_689,In_1143);
nand U1930 (N_1930,In_1151,In_1122);
and U1931 (N_1931,In_1347,In_612);
or U1932 (N_1932,In_1069,In_997);
nor U1933 (N_1933,In_217,In_212);
and U1934 (N_1934,In_250,In_944);
nand U1935 (N_1935,In_163,In_184);
or U1936 (N_1936,In_1321,In_989);
nand U1937 (N_1937,In_1064,In_667);
or U1938 (N_1938,In_1289,In_214);
nand U1939 (N_1939,In_457,In_6);
or U1940 (N_1940,In_335,In_1131);
nand U1941 (N_1941,In_1459,In_729);
and U1942 (N_1942,In_1057,In_1186);
or U1943 (N_1943,In_739,In_1484);
nand U1944 (N_1944,In_498,In_825);
nand U1945 (N_1945,In_232,In_975);
or U1946 (N_1946,In_1221,In_715);
nand U1947 (N_1947,In_200,In_991);
or U1948 (N_1948,In_499,In_685);
nor U1949 (N_1949,In_1186,In_32);
nor U1950 (N_1950,In_1356,In_1358);
nor U1951 (N_1951,In_1027,In_965);
and U1952 (N_1952,In_1371,In_564);
nor U1953 (N_1953,In_102,In_927);
and U1954 (N_1954,In_1198,In_1482);
and U1955 (N_1955,In_433,In_724);
or U1956 (N_1956,In_349,In_131);
nor U1957 (N_1957,In_525,In_1183);
or U1958 (N_1958,In_1402,In_1309);
and U1959 (N_1959,In_356,In_972);
nand U1960 (N_1960,In_519,In_1329);
and U1961 (N_1961,In_1062,In_200);
or U1962 (N_1962,In_694,In_133);
nor U1963 (N_1963,In_567,In_1394);
and U1964 (N_1964,In_1279,In_654);
nand U1965 (N_1965,In_1420,In_1422);
nor U1966 (N_1966,In_906,In_74);
nor U1967 (N_1967,In_1363,In_37);
or U1968 (N_1968,In_485,In_885);
and U1969 (N_1969,In_15,In_315);
nand U1970 (N_1970,In_952,In_165);
nor U1971 (N_1971,In_167,In_225);
nor U1972 (N_1972,In_1250,In_494);
nand U1973 (N_1973,In_845,In_773);
nor U1974 (N_1974,In_573,In_658);
nor U1975 (N_1975,In_830,In_378);
nor U1976 (N_1976,In_1490,In_1101);
or U1977 (N_1977,In_799,In_1147);
nor U1978 (N_1978,In_348,In_1442);
nor U1979 (N_1979,In_19,In_1009);
or U1980 (N_1980,In_1073,In_1286);
nand U1981 (N_1981,In_561,In_950);
nand U1982 (N_1982,In_1146,In_669);
and U1983 (N_1983,In_1079,In_1086);
or U1984 (N_1984,In_109,In_1266);
and U1985 (N_1985,In_934,In_377);
nand U1986 (N_1986,In_1319,In_868);
and U1987 (N_1987,In_1110,In_445);
nand U1988 (N_1988,In_1441,In_1412);
nand U1989 (N_1989,In_1038,In_47);
nand U1990 (N_1990,In_596,In_1225);
nand U1991 (N_1991,In_226,In_1001);
and U1992 (N_1992,In_46,In_135);
or U1993 (N_1993,In_408,In_448);
nor U1994 (N_1994,In_1189,In_1331);
and U1995 (N_1995,In_353,In_1055);
nand U1996 (N_1996,In_1027,In_1359);
and U1997 (N_1997,In_1210,In_790);
nand U1998 (N_1998,In_642,In_773);
xnor U1999 (N_1999,In_1398,In_1120);
and U2000 (N_2000,In_179,In_1399);
nor U2001 (N_2001,In_396,In_627);
or U2002 (N_2002,In_344,In_212);
and U2003 (N_2003,In_118,In_983);
nor U2004 (N_2004,In_1348,In_1116);
nor U2005 (N_2005,In_257,In_100);
nand U2006 (N_2006,In_869,In_811);
or U2007 (N_2007,In_1275,In_1362);
and U2008 (N_2008,In_277,In_168);
nor U2009 (N_2009,In_1334,In_888);
nor U2010 (N_2010,In_423,In_171);
or U2011 (N_2011,In_920,In_880);
nor U2012 (N_2012,In_146,In_1309);
and U2013 (N_2013,In_685,In_844);
and U2014 (N_2014,In_1004,In_1485);
or U2015 (N_2015,In_926,In_98);
and U2016 (N_2016,In_1271,In_536);
nor U2017 (N_2017,In_1167,In_1452);
nor U2018 (N_2018,In_1301,In_565);
and U2019 (N_2019,In_559,In_391);
nor U2020 (N_2020,In_1172,In_1067);
nor U2021 (N_2021,In_122,In_385);
nor U2022 (N_2022,In_238,In_1372);
nand U2023 (N_2023,In_559,In_1339);
and U2024 (N_2024,In_1243,In_494);
and U2025 (N_2025,In_647,In_1203);
nor U2026 (N_2026,In_419,In_417);
nor U2027 (N_2027,In_1339,In_452);
nor U2028 (N_2028,In_204,In_680);
nor U2029 (N_2029,In_907,In_595);
nor U2030 (N_2030,In_437,In_1049);
or U2031 (N_2031,In_706,In_131);
or U2032 (N_2032,In_1322,In_1372);
nand U2033 (N_2033,In_1466,In_809);
or U2034 (N_2034,In_1173,In_804);
nor U2035 (N_2035,In_776,In_980);
or U2036 (N_2036,In_849,In_594);
or U2037 (N_2037,In_404,In_206);
nor U2038 (N_2038,In_403,In_704);
nand U2039 (N_2039,In_3,In_738);
nor U2040 (N_2040,In_977,In_61);
nand U2041 (N_2041,In_1180,In_709);
or U2042 (N_2042,In_569,In_1209);
and U2043 (N_2043,In_424,In_217);
and U2044 (N_2044,In_573,In_359);
nand U2045 (N_2045,In_420,In_1097);
or U2046 (N_2046,In_259,In_717);
or U2047 (N_2047,In_869,In_1320);
or U2048 (N_2048,In_108,In_961);
nor U2049 (N_2049,In_965,In_200);
nand U2050 (N_2050,In_132,In_153);
or U2051 (N_2051,In_70,In_19);
nand U2052 (N_2052,In_293,In_886);
nor U2053 (N_2053,In_186,In_1016);
nor U2054 (N_2054,In_502,In_184);
and U2055 (N_2055,In_123,In_1222);
and U2056 (N_2056,In_614,In_478);
nand U2057 (N_2057,In_1240,In_1112);
nor U2058 (N_2058,In_1046,In_1467);
nor U2059 (N_2059,In_849,In_1424);
or U2060 (N_2060,In_118,In_374);
and U2061 (N_2061,In_508,In_1028);
nor U2062 (N_2062,In_364,In_88);
and U2063 (N_2063,In_43,In_701);
or U2064 (N_2064,In_35,In_726);
nor U2065 (N_2065,In_211,In_821);
or U2066 (N_2066,In_1166,In_493);
nand U2067 (N_2067,In_159,In_404);
and U2068 (N_2068,In_8,In_1037);
and U2069 (N_2069,In_1307,In_1231);
nor U2070 (N_2070,In_637,In_1189);
nor U2071 (N_2071,In_1175,In_1051);
nor U2072 (N_2072,In_1327,In_24);
nand U2073 (N_2073,In_834,In_606);
and U2074 (N_2074,In_715,In_1418);
or U2075 (N_2075,In_1494,In_222);
nand U2076 (N_2076,In_362,In_878);
xnor U2077 (N_2077,In_1001,In_897);
nand U2078 (N_2078,In_1316,In_546);
nand U2079 (N_2079,In_1013,In_1108);
or U2080 (N_2080,In_1050,In_609);
nor U2081 (N_2081,In_780,In_1059);
nand U2082 (N_2082,In_466,In_871);
nand U2083 (N_2083,In_868,In_130);
or U2084 (N_2084,In_1220,In_255);
nor U2085 (N_2085,In_964,In_432);
and U2086 (N_2086,In_281,In_489);
nor U2087 (N_2087,In_1175,In_388);
nand U2088 (N_2088,In_780,In_400);
nand U2089 (N_2089,In_1322,In_814);
nand U2090 (N_2090,In_675,In_1137);
or U2091 (N_2091,In_1084,In_1418);
nor U2092 (N_2092,In_12,In_7);
nand U2093 (N_2093,In_1486,In_436);
nand U2094 (N_2094,In_577,In_237);
nor U2095 (N_2095,In_42,In_579);
nor U2096 (N_2096,In_249,In_1448);
nand U2097 (N_2097,In_925,In_1207);
nand U2098 (N_2098,In_433,In_59);
nor U2099 (N_2099,In_1200,In_1415);
nor U2100 (N_2100,In_690,In_1427);
nand U2101 (N_2101,In_1239,In_183);
nand U2102 (N_2102,In_1162,In_1248);
and U2103 (N_2103,In_1493,In_592);
nor U2104 (N_2104,In_1393,In_1333);
nor U2105 (N_2105,In_1000,In_1460);
or U2106 (N_2106,In_1405,In_742);
nand U2107 (N_2107,In_772,In_1133);
and U2108 (N_2108,In_1141,In_848);
or U2109 (N_2109,In_105,In_472);
and U2110 (N_2110,In_700,In_240);
and U2111 (N_2111,In_1397,In_1030);
nor U2112 (N_2112,In_685,In_355);
or U2113 (N_2113,In_1397,In_439);
nor U2114 (N_2114,In_1321,In_714);
and U2115 (N_2115,In_278,In_341);
and U2116 (N_2116,In_766,In_1421);
and U2117 (N_2117,In_53,In_1425);
and U2118 (N_2118,In_977,In_277);
nor U2119 (N_2119,In_1390,In_1054);
nor U2120 (N_2120,In_219,In_939);
nor U2121 (N_2121,In_1309,In_747);
or U2122 (N_2122,In_811,In_375);
xor U2123 (N_2123,In_1400,In_207);
nor U2124 (N_2124,In_261,In_863);
and U2125 (N_2125,In_11,In_1071);
or U2126 (N_2126,In_894,In_1101);
nor U2127 (N_2127,In_1460,In_708);
and U2128 (N_2128,In_1410,In_532);
and U2129 (N_2129,In_1344,In_753);
or U2130 (N_2130,In_901,In_1108);
and U2131 (N_2131,In_945,In_401);
nor U2132 (N_2132,In_1352,In_52);
and U2133 (N_2133,In_966,In_127);
nand U2134 (N_2134,In_1445,In_203);
or U2135 (N_2135,In_818,In_33);
nor U2136 (N_2136,In_718,In_985);
nor U2137 (N_2137,In_22,In_970);
and U2138 (N_2138,In_479,In_545);
or U2139 (N_2139,In_1167,In_921);
or U2140 (N_2140,In_494,In_399);
and U2141 (N_2141,In_1457,In_699);
and U2142 (N_2142,In_59,In_129);
nand U2143 (N_2143,In_1174,In_845);
nand U2144 (N_2144,In_1333,In_369);
or U2145 (N_2145,In_1075,In_854);
or U2146 (N_2146,In_40,In_1073);
or U2147 (N_2147,In_895,In_614);
nand U2148 (N_2148,In_1050,In_1369);
nor U2149 (N_2149,In_224,In_688);
nor U2150 (N_2150,In_827,In_5);
nand U2151 (N_2151,In_208,In_1397);
and U2152 (N_2152,In_701,In_1241);
and U2153 (N_2153,In_1286,In_1131);
nand U2154 (N_2154,In_1251,In_172);
nand U2155 (N_2155,In_500,In_282);
or U2156 (N_2156,In_394,In_248);
or U2157 (N_2157,In_34,In_1432);
nand U2158 (N_2158,In_689,In_353);
nand U2159 (N_2159,In_799,In_778);
nor U2160 (N_2160,In_355,In_1303);
and U2161 (N_2161,In_619,In_803);
nand U2162 (N_2162,In_771,In_66);
and U2163 (N_2163,In_1279,In_690);
or U2164 (N_2164,In_491,In_1220);
and U2165 (N_2165,In_869,In_1091);
nor U2166 (N_2166,In_1376,In_1232);
or U2167 (N_2167,In_140,In_1464);
and U2168 (N_2168,In_803,In_1391);
or U2169 (N_2169,In_272,In_633);
or U2170 (N_2170,In_1394,In_1123);
nand U2171 (N_2171,In_558,In_411);
nand U2172 (N_2172,In_244,In_916);
nor U2173 (N_2173,In_520,In_738);
nor U2174 (N_2174,In_98,In_1401);
nand U2175 (N_2175,In_119,In_1413);
or U2176 (N_2176,In_256,In_640);
nor U2177 (N_2177,In_52,In_528);
xnor U2178 (N_2178,In_1005,In_391);
nor U2179 (N_2179,In_959,In_645);
nor U2180 (N_2180,In_355,In_1051);
and U2181 (N_2181,In_650,In_342);
or U2182 (N_2182,In_656,In_613);
nand U2183 (N_2183,In_568,In_574);
and U2184 (N_2184,In_339,In_80);
and U2185 (N_2185,In_1168,In_727);
nor U2186 (N_2186,In_1118,In_789);
nor U2187 (N_2187,In_517,In_750);
or U2188 (N_2188,In_865,In_4);
or U2189 (N_2189,In_312,In_298);
or U2190 (N_2190,In_614,In_308);
or U2191 (N_2191,In_233,In_358);
or U2192 (N_2192,In_323,In_819);
nand U2193 (N_2193,In_696,In_319);
and U2194 (N_2194,In_1280,In_1393);
or U2195 (N_2195,In_345,In_413);
and U2196 (N_2196,In_806,In_1287);
or U2197 (N_2197,In_1257,In_885);
nor U2198 (N_2198,In_817,In_972);
and U2199 (N_2199,In_533,In_310);
nor U2200 (N_2200,In_322,In_461);
or U2201 (N_2201,In_916,In_768);
or U2202 (N_2202,In_522,In_978);
and U2203 (N_2203,In_1100,In_1414);
and U2204 (N_2204,In_473,In_1024);
nand U2205 (N_2205,In_644,In_577);
or U2206 (N_2206,In_960,In_781);
and U2207 (N_2207,In_1403,In_1224);
and U2208 (N_2208,In_110,In_1018);
or U2209 (N_2209,In_376,In_1034);
nor U2210 (N_2210,In_156,In_966);
nand U2211 (N_2211,In_529,In_1348);
and U2212 (N_2212,In_54,In_1499);
nand U2213 (N_2213,In_405,In_631);
nand U2214 (N_2214,In_759,In_772);
nand U2215 (N_2215,In_7,In_1181);
or U2216 (N_2216,In_103,In_1021);
or U2217 (N_2217,In_466,In_703);
nor U2218 (N_2218,In_508,In_1446);
nor U2219 (N_2219,In_968,In_239);
and U2220 (N_2220,In_15,In_608);
nand U2221 (N_2221,In_1350,In_776);
nor U2222 (N_2222,In_269,In_1140);
and U2223 (N_2223,In_1121,In_811);
and U2224 (N_2224,In_361,In_1315);
nor U2225 (N_2225,In_621,In_1258);
and U2226 (N_2226,In_1254,In_755);
and U2227 (N_2227,In_1467,In_807);
nor U2228 (N_2228,In_796,In_754);
nor U2229 (N_2229,In_657,In_1314);
xnor U2230 (N_2230,In_468,In_639);
nand U2231 (N_2231,In_1010,In_197);
nand U2232 (N_2232,In_1498,In_854);
and U2233 (N_2233,In_1121,In_483);
nand U2234 (N_2234,In_506,In_831);
and U2235 (N_2235,In_1360,In_709);
and U2236 (N_2236,In_711,In_1061);
nand U2237 (N_2237,In_146,In_466);
or U2238 (N_2238,In_515,In_738);
nor U2239 (N_2239,In_371,In_790);
or U2240 (N_2240,In_486,In_193);
and U2241 (N_2241,In_1425,In_455);
nand U2242 (N_2242,In_1357,In_61);
and U2243 (N_2243,In_181,In_1471);
and U2244 (N_2244,In_839,In_1245);
nand U2245 (N_2245,In_1276,In_123);
nor U2246 (N_2246,In_438,In_1163);
and U2247 (N_2247,In_1378,In_1385);
nor U2248 (N_2248,In_656,In_996);
nor U2249 (N_2249,In_55,In_178);
nor U2250 (N_2250,In_959,In_1090);
nand U2251 (N_2251,In_415,In_442);
or U2252 (N_2252,In_1334,In_1092);
nor U2253 (N_2253,In_849,In_1420);
or U2254 (N_2254,In_467,In_1434);
or U2255 (N_2255,In_1011,In_3);
or U2256 (N_2256,In_1411,In_628);
nand U2257 (N_2257,In_480,In_268);
nand U2258 (N_2258,In_1170,In_1049);
and U2259 (N_2259,In_458,In_585);
or U2260 (N_2260,In_566,In_1204);
nor U2261 (N_2261,In_1184,In_1155);
nand U2262 (N_2262,In_561,In_211);
or U2263 (N_2263,In_1141,In_302);
nor U2264 (N_2264,In_759,In_756);
or U2265 (N_2265,In_571,In_314);
and U2266 (N_2266,In_773,In_1227);
or U2267 (N_2267,In_824,In_412);
and U2268 (N_2268,In_837,In_420);
or U2269 (N_2269,In_428,In_1206);
or U2270 (N_2270,In_788,In_432);
nor U2271 (N_2271,In_73,In_538);
nand U2272 (N_2272,In_1386,In_1104);
nand U2273 (N_2273,In_443,In_451);
nor U2274 (N_2274,In_362,In_960);
nand U2275 (N_2275,In_831,In_1114);
nand U2276 (N_2276,In_1387,In_827);
or U2277 (N_2277,In_1158,In_458);
or U2278 (N_2278,In_548,In_1453);
nand U2279 (N_2279,In_216,In_760);
nor U2280 (N_2280,In_772,In_515);
and U2281 (N_2281,In_249,In_480);
xor U2282 (N_2282,In_311,In_1120);
nor U2283 (N_2283,In_1325,In_1044);
and U2284 (N_2284,In_647,In_1079);
nand U2285 (N_2285,In_209,In_1317);
and U2286 (N_2286,In_548,In_70);
and U2287 (N_2287,In_780,In_919);
nand U2288 (N_2288,In_970,In_346);
nor U2289 (N_2289,In_1357,In_1079);
and U2290 (N_2290,In_1304,In_1477);
nor U2291 (N_2291,In_1104,In_755);
or U2292 (N_2292,In_1181,In_1052);
nor U2293 (N_2293,In_976,In_969);
nand U2294 (N_2294,In_564,In_990);
xor U2295 (N_2295,In_880,In_915);
nand U2296 (N_2296,In_991,In_1070);
nand U2297 (N_2297,In_180,In_957);
nand U2298 (N_2298,In_756,In_987);
nor U2299 (N_2299,In_553,In_23);
nand U2300 (N_2300,In_1341,In_312);
or U2301 (N_2301,In_309,In_902);
nand U2302 (N_2302,In_423,In_701);
nand U2303 (N_2303,In_1052,In_141);
nor U2304 (N_2304,In_1424,In_1062);
nor U2305 (N_2305,In_1441,In_456);
and U2306 (N_2306,In_958,In_1462);
nand U2307 (N_2307,In_1417,In_1358);
nor U2308 (N_2308,In_814,In_82);
or U2309 (N_2309,In_278,In_227);
and U2310 (N_2310,In_352,In_423);
nand U2311 (N_2311,In_968,In_1448);
and U2312 (N_2312,In_302,In_1346);
or U2313 (N_2313,In_89,In_701);
or U2314 (N_2314,In_232,In_667);
or U2315 (N_2315,In_1246,In_1269);
or U2316 (N_2316,In_1082,In_747);
nor U2317 (N_2317,In_937,In_520);
nor U2318 (N_2318,In_999,In_719);
and U2319 (N_2319,In_300,In_945);
and U2320 (N_2320,In_52,In_1476);
nand U2321 (N_2321,In_639,In_1159);
and U2322 (N_2322,In_522,In_15);
nor U2323 (N_2323,In_909,In_1370);
and U2324 (N_2324,In_997,In_991);
or U2325 (N_2325,In_1010,In_230);
nor U2326 (N_2326,In_1445,In_1498);
or U2327 (N_2327,In_359,In_467);
nor U2328 (N_2328,In_185,In_383);
and U2329 (N_2329,In_928,In_1187);
and U2330 (N_2330,In_879,In_1202);
xor U2331 (N_2331,In_488,In_706);
nand U2332 (N_2332,In_556,In_877);
or U2333 (N_2333,In_404,In_826);
or U2334 (N_2334,In_975,In_1447);
nand U2335 (N_2335,In_165,In_704);
or U2336 (N_2336,In_68,In_382);
nand U2337 (N_2337,In_1243,In_1314);
nand U2338 (N_2338,In_1327,In_1454);
or U2339 (N_2339,In_1374,In_703);
nand U2340 (N_2340,In_491,In_1079);
nor U2341 (N_2341,In_1400,In_380);
and U2342 (N_2342,In_571,In_253);
and U2343 (N_2343,In_675,In_805);
and U2344 (N_2344,In_508,In_109);
or U2345 (N_2345,In_199,In_1123);
nor U2346 (N_2346,In_475,In_1011);
or U2347 (N_2347,In_1457,In_312);
nand U2348 (N_2348,In_379,In_408);
nand U2349 (N_2349,In_1266,In_1186);
or U2350 (N_2350,In_1176,In_1097);
nor U2351 (N_2351,In_685,In_447);
or U2352 (N_2352,In_35,In_584);
nor U2353 (N_2353,In_661,In_1076);
or U2354 (N_2354,In_356,In_520);
nor U2355 (N_2355,In_110,In_865);
nand U2356 (N_2356,In_1113,In_1045);
nor U2357 (N_2357,In_656,In_540);
and U2358 (N_2358,In_1298,In_132);
and U2359 (N_2359,In_29,In_1051);
nand U2360 (N_2360,In_1043,In_1496);
or U2361 (N_2361,In_611,In_316);
or U2362 (N_2362,In_195,In_109);
or U2363 (N_2363,In_1355,In_1322);
and U2364 (N_2364,In_553,In_1215);
or U2365 (N_2365,In_247,In_224);
or U2366 (N_2366,In_218,In_198);
and U2367 (N_2367,In_919,In_422);
nor U2368 (N_2368,In_190,In_1266);
and U2369 (N_2369,In_953,In_54);
nor U2370 (N_2370,In_175,In_563);
nor U2371 (N_2371,In_389,In_1390);
nand U2372 (N_2372,In_338,In_689);
or U2373 (N_2373,In_1020,In_485);
nand U2374 (N_2374,In_311,In_1306);
nand U2375 (N_2375,In_1021,In_366);
or U2376 (N_2376,In_419,In_1119);
or U2377 (N_2377,In_724,In_210);
or U2378 (N_2378,In_955,In_829);
nor U2379 (N_2379,In_925,In_642);
nor U2380 (N_2380,In_721,In_1236);
nor U2381 (N_2381,In_177,In_117);
nor U2382 (N_2382,In_774,In_65);
and U2383 (N_2383,In_186,In_1455);
xor U2384 (N_2384,In_695,In_146);
nand U2385 (N_2385,In_609,In_1128);
and U2386 (N_2386,In_42,In_207);
nor U2387 (N_2387,In_286,In_73);
or U2388 (N_2388,In_1378,In_953);
nor U2389 (N_2389,In_81,In_1433);
nand U2390 (N_2390,In_117,In_700);
and U2391 (N_2391,In_687,In_518);
and U2392 (N_2392,In_1291,In_179);
and U2393 (N_2393,In_339,In_449);
nand U2394 (N_2394,In_964,In_247);
nand U2395 (N_2395,In_250,In_363);
or U2396 (N_2396,In_1352,In_639);
or U2397 (N_2397,In_1364,In_147);
nor U2398 (N_2398,In_699,In_1086);
nand U2399 (N_2399,In_164,In_772);
and U2400 (N_2400,In_1059,In_995);
or U2401 (N_2401,In_481,In_1431);
nor U2402 (N_2402,In_1059,In_758);
nor U2403 (N_2403,In_1338,In_1218);
and U2404 (N_2404,In_1420,In_191);
nand U2405 (N_2405,In_248,In_1492);
nor U2406 (N_2406,In_1040,In_1078);
nor U2407 (N_2407,In_1186,In_387);
and U2408 (N_2408,In_668,In_1431);
and U2409 (N_2409,In_1279,In_864);
and U2410 (N_2410,In_213,In_1434);
nand U2411 (N_2411,In_661,In_996);
nand U2412 (N_2412,In_61,In_1204);
nor U2413 (N_2413,In_582,In_11);
or U2414 (N_2414,In_1230,In_886);
or U2415 (N_2415,In_1085,In_1180);
nor U2416 (N_2416,In_1261,In_867);
nand U2417 (N_2417,In_921,In_1484);
and U2418 (N_2418,In_1154,In_989);
or U2419 (N_2419,In_761,In_791);
and U2420 (N_2420,In_1155,In_907);
or U2421 (N_2421,In_1133,In_1487);
and U2422 (N_2422,In_271,In_943);
nand U2423 (N_2423,In_479,In_91);
nor U2424 (N_2424,In_731,In_884);
nand U2425 (N_2425,In_1280,In_591);
and U2426 (N_2426,In_1338,In_771);
nand U2427 (N_2427,In_1038,In_802);
nand U2428 (N_2428,In_941,In_1134);
nand U2429 (N_2429,In_250,In_1272);
nand U2430 (N_2430,In_1239,In_378);
and U2431 (N_2431,In_121,In_832);
nand U2432 (N_2432,In_299,In_955);
nor U2433 (N_2433,In_1314,In_1460);
or U2434 (N_2434,In_1097,In_1356);
and U2435 (N_2435,In_381,In_1192);
and U2436 (N_2436,In_1044,In_1236);
or U2437 (N_2437,In_1470,In_543);
or U2438 (N_2438,In_560,In_687);
and U2439 (N_2439,In_1127,In_763);
or U2440 (N_2440,In_764,In_644);
or U2441 (N_2441,In_1182,In_779);
and U2442 (N_2442,In_292,In_1450);
nor U2443 (N_2443,In_781,In_220);
or U2444 (N_2444,In_295,In_804);
or U2445 (N_2445,In_66,In_449);
xor U2446 (N_2446,In_697,In_33);
and U2447 (N_2447,In_434,In_1207);
nor U2448 (N_2448,In_68,In_289);
nand U2449 (N_2449,In_349,In_120);
nor U2450 (N_2450,In_413,In_801);
and U2451 (N_2451,In_607,In_1218);
xor U2452 (N_2452,In_864,In_833);
or U2453 (N_2453,In_551,In_661);
nand U2454 (N_2454,In_261,In_198);
nor U2455 (N_2455,In_605,In_139);
and U2456 (N_2456,In_222,In_992);
nor U2457 (N_2457,In_917,In_753);
nand U2458 (N_2458,In_439,In_1160);
or U2459 (N_2459,In_376,In_573);
nand U2460 (N_2460,In_236,In_952);
nor U2461 (N_2461,In_292,In_406);
and U2462 (N_2462,In_1204,In_279);
nand U2463 (N_2463,In_592,In_1255);
nor U2464 (N_2464,In_223,In_45);
nor U2465 (N_2465,In_1031,In_73);
nor U2466 (N_2466,In_1488,In_127);
nor U2467 (N_2467,In_1445,In_703);
nor U2468 (N_2468,In_1316,In_690);
nor U2469 (N_2469,In_30,In_859);
and U2470 (N_2470,In_877,In_398);
nand U2471 (N_2471,In_817,In_14);
or U2472 (N_2472,In_1321,In_162);
and U2473 (N_2473,In_424,In_1372);
or U2474 (N_2474,In_888,In_726);
nand U2475 (N_2475,In_46,In_1132);
nor U2476 (N_2476,In_131,In_1311);
and U2477 (N_2477,In_547,In_1038);
and U2478 (N_2478,In_525,In_327);
nor U2479 (N_2479,In_684,In_805);
nor U2480 (N_2480,In_1004,In_1169);
nand U2481 (N_2481,In_559,In_1367);
nand U2482 (N_2482,In_139,In_955);
and U2483 (N_2483,In_331,In_633);
and U2484 (N_2484,In_389,In_882);
or U2485 (N_2485,In_379,In_44);
nand U2486 (N_2486,In_1147,In_176);
xor U2487 (N_2487,In_1081,In_1159);
or U2488 (N_2488,In_554,In_549);
nor U2489 (N_2489,In_605,In_130);
nand U2490 (N_2490,In_1320,In_1012);
or U2491 (N_2491,In_762,In_130);
nand U2492 (N_2492,In_504,In_119);
or U2493 (N_2493,In_37,In_881);
or U2494 (N_2494,In_1383,In_1135);
and U2495 (N_2495,In_821,In_844);
nor U2496 (N_2496,In_907,In_485);
and U2497 (N_2497,In_949,In_518);
and U2498 (N_2498,In_176,In_454);
and U2499 (N_2499,In_545,In_1269);
nand U2500 (N_2500,In_168,In_1047);
and U2501 (N_2501,In_311,In_1465);
and U2502 (N_2502,In_845,In_1284);
or U2503 (N_2503,In_1493,In_994);
or U2504 (N_2504,In_337,In_124);
or U2505 (N_2505,In_604,In_669);
xor U2506 (N_2506,In_374,In_334);
nand U2507 (N_2507,In_267,In_1186);
nand U2508 (N_2508,In_74,In_1339);
nand U2509 (N_2509,In_245,In_1392);
or U2510 (N_2510,In_939,In_1494);
or U2511 (N_2511,In_347,In_1007);
and U2512 (N_2512,In_995,In_1234);
nor U2513 (N_2513,In_717,In_674);
nor U2514 (N_2514,In_132,In_368);
nand U2515 (N_2515,In_1275,In_12);
nand U2516 (N_2516,In_213,In_1456);
nand U2517 (N_2517,In_1048,In_127);
nand U2518 (N_2518,In_1067,In_701);
nor U2519 (N_2519,In_41,In_421);
and U2520 (N_2520,In_1340,In_1071);
or U2521 (N_2521,In_948,In_131);
nor U2522 (N_2522,In_848,In_130);
nor U2523 (N_2523,In_1420,In_435);
or U2524 (N_2524,In_1338,In_932);
nor U2525 (N_2525,In_1090,In_1274);
nand U2526 (N_2526,In_1314,In_190);
xor U2527 (N_2527,In_482,In_852);
or U2528 (N_2528,In_1286,In_77);
and U2529 (N_2529,In_929,In_1113);
nand U2530 (N_2530,In_423,In_138);
and U2531 (N_2531,In_317,In_217);
nor U2532 (N_2532,In_1004,In_1332);
nor U2533 (N_2533,In_530,In_145);
or U2534 (N_2534,In_1367,In_1361);
and U2535 (N_2535,In_223,In_1084);
or U2536 (N_2536,In_62,In_994);
and U2537 (N_2537,In_728,In_132);
nand U2538 (N_2538,In_554,In_1293);
nand U2539 (N_2539,In_888,In_1348);
xnor U2540 (N_2540,In_1124,In_551);
and U2541 (N_2541,In_1377,In_781);
and U2542 (N_2542,In_744,In_1201);
nand U2543 (N_2543,In_1211,In_462);
or U2544 (N_2544,In_305,In_283);
nor U2545 (N_2545,In_323,In_900);
nand U2546 (N_2546,In_838,In_911);
nand U2547 (N_2547,In_1301,In_801);
nor U2548 (N_2548,In_605,In_455);
nand U2549 (N_2549,In_247,In_287);
nand U2550 (N_2550,In_380,In_821);
and U2551 (N_2551,In_1295,In_1103);
nor U2552 (N_2552,In_499,In_1019);
nand U2553 (N_2553,In_1163,In_1286);
nor U2554 (N_2554,In_678,In_558);
or U2555 (N_2555,In_490,In_379);
nand U2556 (N_2556,In_902,In_1235);
nand U2557 (N_2557,In_719,In_526);
or U2558 (N_2558,In_159,In_333);
and U2559 (N_2559,In_152,In_685);
nand U2560 (N_2560,In_42,In_1167);
nor U2561 (N_2561,In_706,In_1190);
and U2562 (N_2562,In_1130,In_690);
and U2563 (N_2563,In_555,In_1356);
nor U2564 (N_2564,In_302,In_498);
nor U2565 (N_2565,In_629,In_601);
nand U2566 (N_2566,In_1261,In_1077);
nand U2567 (N_2567,In_163,In_431);
nor U2568 (N_2568,In_790,In_1406);
and U2569 (N_2569,In_337,In_364);
and U2570 (N_2570,In_860,In_45);
nand U2571 (N_2571,In_638,In_245);
nand U2572 (N_2572,In_1015,In_17);
and U2573 (N_2573,In_1298,In_648);
nand U2574 (N_2574,In_590,In_885);
and U2575 (N_2575,In_730,In_208);
nor U2576 (N_2576,In_977,In_1440);
or U2577 (N_2577,In_627,In_351);
and U2578 (N_2578,In_399,In_977);
nor U2579 (N_2579,In_272,In_834);
nor U2580 (N_2580,In_641,In_316);
or U2581 (N_2581,In_315,In_1037);
and U2582 (N_2582,In_726,In_540);
or U2583 (N_2583,In_684,In_1024);
or U2584 (N_2584,In_1355,In_97);
nand U2585 (N_2585,In_70,In_813);
xor U2586 (N_2586,In_1119,In_1117);
and U2587 (N_2587,In_1476,In_149);
nand U2588 (N_2588,In_1491,In_726);
and U2589 (N_2589,In_203,In_376);
nand U2590 (N_2590,In_158,In_222);
and U2591 (N_2591,In_1185,In_1191);
nand U2592 (N_2592,In_292,In_116);
or U2593 (N_2593,In_56,In_1204);
and U2594 (N_2594,In_1041,In_303);
xor U2595 (N_2595,In_229,In_594);
or U2596 (N_2596,In_643,In_1025);
nand U2597 (N_2597,In_1366,In_750);
and U2598 (N_2598,In_365,In_1104);
nand U2599 (N_2599,In_314,In_494);
or U2600 (N_2600,In_1364,In_945);
nor U2601 (N_2601,In_500,In_163);
or U2602 (N_2602,In_746,In_410);
and U2603 (N_2603,In_1341,In_765);
nand U2604 (N_2604,In_1012,In_1123);
or U2605 (N_2605,In_1005,In_103);
xnor U2606 (N_2606,In_445,In_1025);
and U2607 (N_2607,In_908,In_1402);
xnor U2608 (N_2608,In_735,In_1097);
and U2609 (N_2609,In_270,In_1449);
nand U2610 (N_2610,In_1085,In_1007);
and U2611 (N_2611,In_68,In_1119);
nand U2612 (N_2612,In_314,In_738);
and U2613 (N_2613,In_559,In_762);
nand U2614 (N_2614,In_503,In_484);
or U2615 (N_2615,In_566,In_892);
and U2616 (N_2616,In_58,In_1229);
nand U2617 (N_2617,In_1377,In_1358);
nor U2618 (N_2618,In_1497,In_249);
nand U2619 (N_2619,In_1172,In_220);
nor U2620 (N_2620,In_515,In_668);
or U2621 (N_2621,In_1132,In_933);
nor U2622 (N_2622,In_1367,In_579);
and U2623 (N_2623,In_31,In_1182);
or U2624 (N_2624,In_1349,In_769);
and U2625 (N_2625,In_175,In_1323);
or U2626 (N_2626,In_1296,In_1220);
or U2627 (N_2627,In_191,In_765);
and U2628 (N_2628,In_402,In_1141);
nand U2629 (N_2629,In_1351,In_958);
and U2630 (N_2630,In_497,In_992);
and U2631 (N_2631,In_832,In_823);
nand U2632 (N_2632,In_229,In_1096);
or U2633 (N_2633,In_415,In_533);
and U2634 (N_2634,In_1066,In_1098);
nand U2635 (N_2635,In_906,In_341);
and U2636 (N_2636,In_1338,In_512);
nor U2637 (N_2637,In_561,In_67);
nor U2638 (N_2638,In_730,In_88);
and U2639 (N_2639,In_1480,In_423);
or U2640 (N_2640,In_1146,In_824);
nand U2641 (N_2641,In_1225,In_615);
nand U2642 (N_2642,In_601,In_760);
nor U2643 (N_2643,In_844,In_60);
nor U2644 (N_2644,In_417,In_853);
and U2645 (N_2645,In_727,In_537);
nor U2646 (N_2646,In_366,In_261);
or U2647 (N_2647,In_448,In_1123);
nand U2648 (N_2648,In_1492,In_4);
and U2649 (N_2649,In_417,In_168);
nand U2650 (N_2650,In_1440,In_284);
or U2651 (N_2651,In_1332,In_599);
nand U2652 (N_2652,In_259,In_1279);
nor U2653 (N_2653,In_650,In_11);
or U2654 (N_2654,In_506,In_784);
and U2655 (N_2655,In_542,In_89);
nand U2656 (N_2656,In_883,In_552);
or U2657 (N_2657,In_235,In_1209);
nor U2658 (N_2658,In_590,In_350);
and U2659 (N_2659,In_363,In_428);
and U2660 (N_2660,In_799,In_547);
and U2661 (N_2661,In_153,In_100);
nand U2662 (N_2662,In_843,In_946);
or U2663 (N_2663,In_814,In_1212);
or U2664 (N_2664,In_1059,In_939);
nor U2665 (N_2665,In_35,In_822);
and U2666 (N_2666,In_795,In_770);
nor U2667 (N_2667,In_289,In_1040);
or U2668 (N_2668,In_295,In_1496);
nand U2669 (N_2669,In_1287,In_173);
nor U2670 (N_2670,In_1174,In_1000);
nor U2671 (N_2671,In_714,In_176);
and U2672 (N_2672,In_93,In_1251);
or U2673 (N_2673,In_458,In_626);
and U2674 (N_2674,In_137,In_1019);
nor U2675 (N_2675,In_177,In_1134);
nand U2676 (N_2676,In_766,In_1031);
nor U2677 (N_2677,In_88,In_1061);
nand U2678 (N_2678,In_654,In_130);
nor U2679 (N_2679,In_531,In_203);
or U2680 (N_2680,In_1491,In_1483);
or U2681 (N_2681,In_629,In_712);
and U2682 (N_2682,In_896,In_375);
nand U2683 (N_2683,In_683,In_206);
and U2684 (N_2684,In_226,In_662);
nand U2685 (N_2685,In_1230,In_88);
and U2686 (N_2686,In_849,In_211);
and U2687 (N_2687,In_1262,In_352);
nand U2688 (N_2688,In_988,In_1224);
nand U2689 (N_2689,In_1408,In_719);
nor U2690 (N_2690,In_412,In_945);
and U2691 (N_2691,In_312,In_96);
and U2692 (N_2692,In_831,In_412);
nand U2693 (N_2693,In_951,In_170);
nor U2694 (N_2694,In_1004,In_947);
nand U2695 (N_2695,In_330,In_284);
nor U2696 (N_2696,In_770,In_523);
nor U2697 (N_2697,In_1455,In_516);
and U2698 (N_2698,In_508,In_603);
or U2699 (N_2699,In_211,In_441);
nor U2700 (N_2700,In_1,In_12);
nor U2701 (N_2701,In_1313,In_1401);
nand U2702 (N_2702,In_414,In_1120);
nor U2703 (N_2703,In_1431,In_1035);
nor U2704 (N_2704,In_1485,In_434);
nor U2705 (N_2705,In_987,In_1027);
nor U2706 (N_2706,In_749,In_174);
xor U2707 (N_2707,In_603,In_1443);
or U2708 (N_2708,In_419,In_1387);
and U2709 (N_2709,In_399,In_668);
or U2710 (N_2710,In_436,In_144);
nor U2711 (N_2711,In_602,In_237);
and U2712 (N_2712,In_1131,In_1436);
or U2713 (N_2713,In_869,In_1239);
nand U2714 (N_2714,In_131,In_862);
and U2715 (N_2715,In_733,In_427);
nand U2716 (N_2716,In_1167,In_329);
nand U2717 (N_2717,In_279,In_1297);
nor U2718 (N_2718,In_80,In_1391);
nor U2719 (N_2719,In_1002,In_30);
and U2720 (N_2720,In_1021,In_1034);
and U2721 (N_2721,In_993,In_1089);
nand U2722 (N_2722,In_1261,In_1303);
nor U2723 (N_2723,In_256,In_410);
xnor U2724 (N_2724,In_1116,In_939);
or U2725 (N_2725,In_570,In_1398);
and U2726 (N_2726,In_276,In_127);
nand U2727 (N_2727,In_514,In_517);
or U2728 (N_2728,In_358,In_1437);
or U2729 (N_2729,In_1209,In_773);
or U2730 (N_2730,In_502,In_282);
and U2731 (N_2731,In_1378,In_930);
or U2732 (N_2732,In_677,In_738);
nand U2733 (N_2733,In_1167,In_511);
and U2734 (N_2734,In_767,In_361);
nor U2735 (N_2735,In_869,In_18);
nor U2736 (N_2736,In_734,In_1312);
nor U2737 (N_2737,In_1360,In_624);
or U2738 (N_2738,In_617,In_1336);
nand U2739 (N_2739,In_110,In_1381);
nand U2740 (N_2740,In_1313,In_1397);
nand U2741 (N_2741,In_851,In_362);
nand U2742 (N_2742,In_889,In_959);
and U2743 (N_2743,In_144,In_1312);
or U2744 (N_2744,In_558,In_446);
nor U2745 (N_2745,In_322,In_360);
or U2746 (N_2746,In_873,In_27);
or U2747 (N_2747,In_763,In_936);
nand U2748 (N_2748,In_958,In_646);
nand U2749 (N_2749,In_248,In_342);
or U2750 (N_2750,In_65,In_490);
nand U2751 (N_2751,In_185,In_522);
nand U2752 (N_2752,In_681,In_1482);
nand U2753 (N_2753,In_460,In_1427);
nand U2754 (N_2754,In_840,In_318);
nand U2755 (N_2755,In_559,In_645);
or U2756 (N_2756,In_212,In_1384);
or U2757 (N_2757,In_883,In_902);
nor U2758 (N_2758,In_1493,In_712);
nor U2759 (N_2759,In_1029,In_864);
nor U2760 (N_2760,In_953,In_1028);
nand U2761 (N_2761,In_316,In_247);
xor U2762 (N_2762,In_219,In_159);
xnor U2763 (N_2763,In_272,In_1494);
or U2764 (N_2764,In_1419,In_940);
and U2765 (N_2765,In_1129,In_1009);
nor U2766 (N_2766,In_628,In_1021);
or U2767 (N_2767,In_518,In_182);
or U2768 (N_2768,In_1056,In_120);
or U2769 (N_2769,In_678,In_326);
nand U2770 (N_2770,In_187,In_938);
nand U2771 (N_2771,In_153,In_70);
and U2772 (N_2772,In_429,In_1448);
nand U2773 (N_2773,In_945,In_1148);
or U2774 (N_2774,In_275,In_1331);
or U2775 (N_2775,In_872,In_9);
or U2776 (N_2776,In_829,In_473);
nor U2777 (N_2777,In_1349,In_1364);
nand U2778 (N_2778,In_813,In_628);
or U2779 (N_2779,In_1198,In_40);
xnor U2780 (N_2780,In_1010,In_252);
and U2781 (N_2781,In_923,In_801);
nand U2782 (N_2782,In_1154,In_669);
and U2783 (N_2783,In_864,In_1069);
and U2784 (N_2784,In_575,In_1218);
nand U2785 (N_2785,In_1464,In_55);
and U2786 (N_2786,In_706,In_445);
and U2787 (N_2787,In_1273,In_912);
or U2788 (N_2788,In_319,In_1209);
or U2789 (N_2789,In_831,In_390);
nand U2790 (N_2790,In_227,In_1116);
xor U2791 (N_2791,In_27,In_1250);
nand U2792 (N_2792,In_741,In_1403);
nor U2793 (N_2793,In_989,In_563);
nand U2794 (N_2794,In_234,In_1005);
and U2795 (N_2795,In_854,In_277);
nand U2796 (N_2796,In_899,In_265);
or U2797 (N_2797,In_493,In_689);
nor U2798 (N_2798,In_83,In_1432);
or U2799 (N_2799,In_916,In_1273);
nor U2800 (N_2800,In_494,In_934);
or U2801 (N_2801,In_613,In_671);
and U2802 (N_2802,In_1397,In_358);
nor U2803 (N_2803,In_908,In_983);
xor U2804 (N_2804,In_1390,In_838);
and U2805 (N_2805,In_443,In_405);
nor U2806 (N_2806,In_1247,In_291);
or U2807 (N_2807,In_305,In_1287);
or U2808 (N_2808,In_1297,In_408);
and U2809 (N_2809,In_428,In_822);
or U2810 (N_2810,In_499,In_1152);
and U2811 (N_2811,In_1397,In_1366);
nor U2812 (N_2812,In_429,In_610);
or U2813 (N_2813,In_883,In_867);
and U2814 (N_2814,In_363,In_422);
nor U2815 (N_2815,In_626,In_465);
nor U2816 (N_2816,In_1032,In_0);
nor U2817 (N_2817,In_1070,In_996);
nand U2818 (N_2818,In_865,In_560);
or U2819 (N_2819,In_251,In_1342);
nand U2820 (N_2820,In_165,In_768);
or U2821 (N_2821,In_1398,In_276);
nand U2822 (N_2822,In_199,In_659);
and U2823 (N_2823,In_794,In_538);
and U2824 (N_2824,In_1000,In_80);
nand U2825 (N_2825,In_647,In_110);
or U2826 (N_2826,In_1181,In_1378);
and U2827 (N_2827,In_1350,In_438);
and U2828 (N_2828,In_655,In_927);
nor U2829 (N_2829,In_1392,In_260);
or U2830 (N_2830,In_1365,In_302);
or U2831 (N_2831,In_201,In_344);
nor U2832 (N_2832,In_1395,In_91);
or U2833 (N_2833,In_597,In_542);
or U2834 (N_2834,In_399,In_810);
and U2835 (N_2835,In_824,In_790);
and U2836 (N_2836,In_1273,In_131);
nand U2837 (N_2837,In_771,In_804);
or U2838 (N_2838,In_470,In_296);
nand U2839 (N_2839,In_718,In_458);
nor U2840 (N_2840,In_238,In_976);
nand U2841 (N_2841,In_147,In_1256);
nor U2842 (N_2842,In_1077,In_9);
nand U2843 (N_2843,In_639,In_1247);
nand U2844 (N_2844,In_1164,In_943);
and U2845 (N_2845,In_330,In_732);
or U2846 (N_2846,In_1390,In_1227);
nand U2847 (N_2847,In_492,In_919);
or U2848 (N_2848,In_1369,In_1327);
nor U2849 (N_2849,In_1478,In_1006);
or U2850 (N_2850,In_12,In_280);
or U2851 (N_2851,In_1392,In_1450);
and U2852 (N_2852,In_1196,In_1294);
and U2853 (N_2853,In_869,In_1277);
and U2854 (N_2854,In_720,In_151);
and U2855 (N_2855,In_670,In_226);
or U2856 (N_2856,In_249,In_545);
nor U2857 (N_2857,In_20,In_1412);
nor U2858 (N_2858,In_1239,In_141);
and U2859 (N_2859,In_917,In_787);
and U2860 (N_2860,In_1247,In_513);
nand U2861 (N_2861,In_318,In_580);
nor U2862 (N_2862,In_435,In_318);
nor U2863 (N_2863,In_290,In_1141);
or U2864 (N_2864,In_20,In_680);
and U2865 (N_2865,In_1440,In_772);
and U2866 (N_2866,In_907,In_1338);
nor U2867 (N_2867,In_1014,In_356);
nor U2868 (N_2868,In_1373,In_629);
and U2869 (N_2869,In_1489,In_1313);
or U2870 (N_2870,In_1308,In_63);
and U2871 (N_2871,In_368,In_170);
nand U2872 (N_2872,In_571,In_582);
nand U2873 (N_2873,In_493,In_742);
nor U2874 (N_2874,In_1345,In_569);
nor U2875 (N_2875,In_1182,In_818);
or U2876 (N_2876,In_42,In_77);
nor U2877 (N_2877,In_700,In_102);
and U2878 (N_2878,In_1216,In_633);
or U2879 (N_2879,In_1237,In_747);
or U2880 (N_2880,In_1320,In_1051);
nor U2881 (N_2881,In_448,In_1055);
and U2882 (N_2882,In_1340,In_88);
nor U2883 (N_2883,In_923,In_34);
nand U2884 (N_2884,In_1298,In_653);
nor U2885 (N_2885,In_1202,In_919);
nor U2886 (N_2886,In_1398,In_220);
nor U2887 (N_2887,In_298,In_1282);
or U2888 (N_2888,In_339,In_792);
nand U2889 (N_2889,In_1439,In_168);
nor U2890 (N_2890,In_291,In_828);
and U2891 (N_2891,In_1242,In_578);
nor U2892 (N_2892,In_1295,In_730);
and U2893 (N_2893,In_759,In_692);
nand U2894 (N_2894,In_1301,In_179);
or U2895 (N_2895,In_52,In_1477);
nor U2896 (N_2896,In_1281,In_372);
nand U2897 (N_2897,In_441,In_862);
and U2898 (N_2898,In_1036,In_1473);
or U2899 (N_2899,In_186,In_524);
xnor U2900 (N_2900,In_880,In_825);
nor U2901 (N_2901,In_1454,In_1261);
and U2902 (N_2902,In_256,In_1078);
nand U2903 (N_2903,In_1434,In_1122);
nand U2904 (N_2904,In_777,In_989);
nand U2905 (N_2905,In_479,In_1267);
or U2906 (N_2906,In_473,In_1332);
and U2907 (N_2907,In_825,In_504);
nor U2908 (N_2908,In_375,In_817);
nand U2909 (N_2909,In_530,In_1187);
or U2910 (N_2910,In_485,In_1033);
and U2911 (N_2911,In_970,In_1199);
nand U2912 (N_2912,In_1398,In_432);
nand U2913 (N_2913,In_1376,In_777);
and U2914 (N_2914,In_944,In_62);
or U2915 (N_2915,In_1104,In_925);
or U2916 (N_2916,In_1386,In_819);
nand U2917 (N_2917,In_575,In_775);
or U2918 (N_2918,In_724,In_135);
nor U2919 (N_2919,In_1001,In_1317);
nand U2920 (N_2920,In_762,In_10);
and U2921 (N_2921,In_379,In_852);
nand U2922 (N_2922,In_430,In_748);
and U2923 (N_2923,In_1036,In_984);
or U2924 (N_2924,In_1329,In_649);
or U2925 (N_2925,In_888,In_1309);
and U2926 (N_2926,In_969,In_618);
or U2927 (N_2927,In_225,In_388);
and U2928 (N_2928,In_1333,In_1303);
or U2929 (N_2929,In_363,In_1146);
nor U2930 (N_2930,In_226,In_257);
nand U2931 (N_2931,In_287,In_375);
xor U2932 (N_2932,In_231,In_570);
nor U2933 (N_2933,In_435,In_134);
xor U2934 (N_2934,In_295,In_1410);
and U2935 (N_2935,In_1388,In_267);
nand U2936 (N_2936,In_826,In_179);
and U2937 (N_2937,In_615,In_1471);
nor U2938 (N_2938,In_109,In_916);
and U2939 (N_2939,In_8,In_539);
or U2940 (N_2940,In_1259,In_1039);
and U2941 (N_2941,In_1130,In_383);
and U2942 (N_2942,In_167,In_363);
nand U2943 (N_2943,In_781,In_11);
nor U2944 (N_2944,In_1202,In_1126);
and U2945 (N_2945,In_414,In_555);
or U2946 (N_2946,In_976,In_404);
and U2947 (N_2947,In_1341,In_1162);
or U2948 (N_2948,In_807,In_1050);
nand U2949 (N_2949,In_1317,In_1065);
and U2950 (N_2950,In_257,In_48);
nand U2951 (N_2951,In_138,In_317);
and U2952 (N_2952,In_1343,In_942);
or U2953 (N_2953,In_6,In_542);
nand U2954 (N_2954,In_888,In_564);
and U2955 (N_2955,In_34,In_924);
or U2956 (N_2956,In_1307,In_586);
nand U2957 (N_2957,In_233,In_1153);
or U2958 (N_2958,In_189,In_297);
and U2959 (N_2959,In_931,In_375);
or U2960 (N_2960,In_167,In_382);
nor U2961 (N_2961,In_1380,In_60);
nand U2962 (N_2962,In_570,In_530);
and U2963 (N_2963,In_1346,In_341);
and U2964 (N_2964,In_266,In_700);
and U2965 (N_2965,In_825,In_1482);
and U2966 (N_2966,In_562,In_1430);
nor U2967 (N_2967,In_1312,In_391);
and U2968 (N_2968,In_128,In_35);
nand U2969 (N_2969,In_21,In_343);
and U2970 (N_2970,In_1283,In_87);
nand U2971 (N_2971,In_841,In_410);
nor U2972 (N_2972,In_590,In_1117);
or U2973 (N_2973,In_253,In_561);
nor U2974 (N_2974,In_605,In_1115);
nor U2975 (N_2975,In_475,In_1199);
nor U2976 (N_2976,In_1041,In_1335);
nand U2977 (N_2977,In_729,In_1020);
nor U2978 (N_2978,In_102,In_237);
nor U2979 (N_2979,In_471,In_263);
nand U2980 (N_2980,In_101,In_5);
or U2981 (N_2981,In_809,In_155);
nor U2982 (N_2982,In_705,In_200);
nor U2983 (N_2983,In_1474,In_317);
nor U2984 (N_2984,In_644,In_6);
nand U2985 (N_2985,In_1441,In_826);
nor U2986 (N_2986,In_253,In_1011);
nor U2987 (N_2987,In_1493,In_236);
nor U2988 (N_2988,In_1040,In_65);
nand U2989 (N_2989,In_1375,In_243);
and U2990 (N_2990,In_1138,In_1495);
or U2991 (N_2991,In_973,In_1098);
nor U2992 (N_2992,In_666,In_1146);
and U2993 (N_2993,In_476,In_1214);
nor U2994 (N_2994,In_69,In_1364);
or U2995 (N_2995,In_1113,In_716);
nor U2996 (N_2996,In_163,In_868);
nor U2997 (N_2997,In_1324,In_853);
and U2998 (N_2998,In_1010,In_906);
and U2999 (N_2999,In_228,In_690);
and U3000 (N_3000,N_1894,N_2207);
nand U3001 (N_3001,N_652,N_2914);
and U3002 (N_3002,N_596,N_879);
and U3003 (N_3003,N_1217,N_1862);
nor U3004 (N_3004,N_1458,N_2783);
nand U3005 (N_3005,N_2334,N_2966);
nand U3006 (N_3006,N_1568,N_2851);
xnor U3007 (N_3007,N_2648,N_2912);
or U3008 (N_3008,N_1758,N_865);
nand U3009 (N_3009,N_972,N_261);
or U3010 (N_3010,N_912,N_66);
nand U3011 (N_3011,N_1275,N_96);
nand U3012 (N_3012,N_644,N_2714);
and U3013 (N_3013,N_2555,N_2995);
nand U3014 (N_3014,N_207,N_1768);
and U3015 (N_3015,N_907,N_759);
or U3016 (N_3016,N_806,N_1678);
nand U3017 (N_3017,N_12,N_2335);
nor U3018 (N_3018,N_924,N_1200);
or U3019 (N_3019,N_1770,N_638);
nand U3020 (N_3020,N_2168,N_567);
nor U3021 (N_3021,N_28,N_2541);
or U3022 (N_3022,N_634,N_2847);
nand U3023 (N_3023,N_250,N_2190);
and U3024 (N_3024,N_2142,N_2318);
nor U3025 (N_3025,N_1381,N_528);
xor U3026 (N_3026,N_1694,N_742);
or U3027 (N_3027,N_1571,N_492);
nor U3028 (N_3028,N_543,N_239);
nor U3029 (N_3029,N_80,N_2181);
and U3030 (N_3030,N_18,N_3);
nand U3031 (N_3031,N_2089,N_2617);
nand U3032 (N_3032,N_2809,N_1643);
or U3033 (N_3033,N_1882,N_1798);
and U3034 (N_3034,N_2401,N_350);
nor U3035 (N_3035,N_2515,N_2143);
and U3036 (N_3036,N_219,N_1548);
or U3037 (N_3037,N_578,N_2696);
nand U3038 (N_3038,N_1633,N_136);
and U3039 (N_3039,N_681,N_958);
or U3040 (N_3040,N_2650,N_1258);
nor U3041 (N_3041,N_1970,N_1473);
and U3042 (N_3042,N_304,N_372);
nand U3043 (N_3043,N_1712,N_1785);
or U3044 (N_3044,N_2016,N_977);
or U3045 (N_3045,N_792,N_14);
nand U3046 (N_3046,N_2742,N_485);
and U3047 (N_3047,N_1925,N_2432);
or U3048 (N_3048,N_1299,N_2057);
nand U3049 (N_3049,N_491,N_108);
xor U3050 (N_3050,N_2377,N_2965);
nand U3051 (N_3051,N_1595,N_2849);
and U3052 (N_3052,N_684,N_2928);
and U3053 (N_3053,N_637,N_2832);
and U3054 (N_3054,N_2102,N_2527);
and U3055 (N_3055,N_2684,N_710);
and U3056 (N_3056,N_1453,N_2224);
or U3057 (N_3057,N_1427,N_1727);
nor U3058 (N_3058,N_2305,N_833);
or U3059 (N_3059,N_2979,N_131);
nor U3060 (N_3060,N_1771,N_887);
or U3061 (N_3061,N_2306,N_377);
nand U3062 (N_3062,N_1435,N_1876);
or U3063 (N_3063,N_2268,N_293);
or U3064 (N_3064,N_2063,N_321);
and U3065 (N_3065,N_730,N_1869);
or U3066 (N_3066,N_1614,N_1684);
or U3067 (N_3067,N_1532,N_2571);
or U3068 (N_3068,N_2596,N_2895);
and U3069 (N_3069,N_768,N_902);
and U3070 (N_3070,N_1114,N_2256);
nand U3071 (N_3071,N_2546,N_698);
and U3072 (N_3072,N_2618,N_199);
nor U3073 (N_3073,N_1272,N_1877);
nand U3074 (N_3074,N_1604,N_712);
or U3075 (N_3075,N_606,N_2449);
xor U3076 (N_3076,N_1756,N_275);
and U3077 (N_3077,N_1985,N_1836);
nand U3078 (N_3078,N_691,N_2606);
or U3079 (N_3079,N_2872,N_271);
nand U3080 (N_3080,N_2670,N_2154);
nand U3081 (N_3081,N_206,N_1020);
or U3082 (N_3082,N_2139,N_1464);
nor U3083 (N_3083,N_2095,N_1372);
nor U3084 (N_3084,N_2624,N_1183);
and U3085 (N_3085,N_772,N_1500);
and U3086 (N_3086,N_1191,N_1971);
nor U3087 (N_3087,N_137,N_1597);
nand U3088 (N_3088,N_2623,N_421);
or U3089 (N_3089,N_138,N_1138);
nand U3090 (N_3090,N_514,N_944);
or U3091 (N_3091,N_1378,N_1454);
nand U3092 (N_3092,N_332,N_2262);
nand U3093 (N_3093,N_550,N_1361);
and U3094 (N_3094,N_1311,N_1920);
nand U3095 (N_3095,N_425,N_807);
or U3096 (N_3096,N_2397,N_1469);
nor U3097 (N_3097,N_397,N_2986);
nor U3098 (N_3098,N_1897,N_2289);
and U3099 (N_3099,N_564,N_2583);
or U3100 (N_3100,N_2850,N_1348);
nand U3101 (N_3101,N_2243,N_1497);
nand U3102 (N_3102,N_1959,N_1806);
nor U3103 (N_3103,N_830,N_1998);
nor U3104 (N_3104,N_437,N_2882);
and U3105 (N_3105,N_2183,N_2421);
or U3106 (N_3106,N_509,N_1105);
and U3107 (N_3107,N_1503,N_969);
nor U3108 (N_3108,N_1159,N_1800);
and U3109 (N_3109,N_2735,N_1573);
and U3110 (N_3110,N_2404,N_1239);
nor U3111 (N_3111,N_587,N_1111);
or U3112 (N_3112,N_410,N_1282);
and U3113 (N_3113,N_282,N_2414);
and U3114 (N_3114,N_1659,N_2941);
and U3115 (N_3115,N_20,N_2091);
nor U3116 (N_3116,N_1775,N_407);
nor U3117 (N_3117,N_2105,N_2343);
or U3118 (N_3118,N_2503,N_2630);
or U3119 (N_3119,N_2645,N_1474);
and U3120 (N_3120,N_486,N_2718);
nor U3121 (N_3121,N_391,N_1247);
nor U3122 (N_3122,N_2675,N_1574);
and U3123 (N_3123,N_458,N_2394);
or U3124 (N_3124,N_1506,N_1161);
and U3125 (N_3125,N_161,N_1695);
nor U3126 (N_3126,N_708,N_2138);
and U3127 (N_3127,N_1491,N_50);
or U3128 (N_3128,N_1011,N_815);
or U3129 (N_3129,N_990,N_975);
and U3130 (N_3130,N_1957,N_2493);
nand U3131 (N_3131,N_2798,N_633);
nand U3132 (N_3132,N_1018,N_2272);
and U3133 (N_3133,N_2940,N_2455);
and U3134 (N_3134,N_1778,N_1271);
or U3135 (N_3135,N_1585,N_1096);
or U3136 (N_3136,N_1001,N_2843);
and U3137 (N_3137,N_2613,N_1893);
and U3138 (N_3138,N_1683,N_2968);
nand U3139 (N_3139,N_754,N_1788);
nand U3140 (N_3140,N_449,N_2413);
and U3141 (N_3141,N_187,N_1617);
nand U3142 (N_3142,N_723,N_71);
or U3143 (N_3143,N_40,N_1637);
nand U3144 (N_3144,N_731,N_1730);
nor U3145 (N_3145,N_1377,N_1208);
and U3146 (N_3146,N_2426,N_429);
or U3147 (N_3147,N_1690,N_383);
or U3148 (N_3148,N_163,N_2944);
nand U3149 (N_3149,N_2549,N_1656);
or U3150 (N_3150,N_1108,N_1563);
or U3151 (N_3151,N_529,N_220);
and U3152 (N_3152,N_94,N_1080);
or U3153 (N_3153,N_2434,N_353);
and U3154 (N_3154,N_2737,N_1179);
nor U3155 (N_3155,N_1687,N_1210);
or U3156 (N_3156,N_2316,N_2239);
nand U3157 (N_3157,N_2865,N_1388);
and U3158 (N_3158,N_2700,N_1946);
and U3159 (N_3159,N_1227,N_547);
and U3160 (N_3160,N_2508,N_1718);
nor U3161 (N_3161,N_1629,N_2204);
or U3162 (N_3162,N_2734,N_2254);
or U3163 (N_3163,N_1205,N_1103);
and U3164 (N_3164,N_2788,N_287);
nor U3165 (N_3165,N_1787,N_1254);
nand U3166 (N_3166,N_2385,N_2892);
nand U3167 (N_3167,N_1776,N_1703);
nand U3168 (N_3168,N_2677,N_982);
nand U3169 (N_3169,N_60,N_1762);
nor U3170 (N_3170,N_2782,N_870);
and U3171 (N_3171,N_1366,N_1000);
nor U3172 (N_3172,N_1467,N_2984);
and U3173 (N_3173,N_249,N_473);
nand U3174 (N_3174,N_1870,N_2486);
nand U3175 (N_3175,N_668,N_517);
nor U3176 (N_3176,N_1655,N_1680);
nand U3177 (N_3177,N_313,N_1763);
and U3178 (N_3178,N_2641,N_1786);
nor U3179 (N_3179,N_1234,N_2667);
or U3180 (N_3180,N_1391,N_1207);
or U3181 (N_3181,N_2717,N_2135);
nand U3182 (N_3182,N_1740,N_1596);
or U3183 (N_3183,N_1173,N_33);
nand U3184 (N_3184,N_1068,N_341);
nand U3185 (N_3185,N_254,N_2857);
and U3186 (N_3186,N_460,N_2299);
nor U3187 (N_3187,N_2946,N_151);
or U3188 (N_3188,N_1074,N_921);
nand U3189 (N_3189,N_1566,N_1398);
or U3190 (N_3190,N_713,N_1496);
nand U3191 (N_3191,N_656,N_2856);
nor U3192 (N_3192,N_2821,N_607);
nand U3193 (N_3193,N_2038,N_677);
and U3194 (N_3194,N_1156,N_2322);
nand U3195 (N_3195,N_941,N_1580);
nor U3196 (N_3196,N_2516,N_843);
or U3197 (N_3197,N_2633,N_1866);
nand U3198 (N_3198,N_2283,N_2548);
and U3199 (N_3199,N_1196,N_305);
or U3200 (N_3200,N_2669,N_1057);
or U3201 (N_3201,N_1390,N_2161);
nand U3202 (N_3202,N_2627,N_1826);
nor U3203 (N_3203,N_1429,N_459);
or U3204 (N_3204,N_2149,N_2032);
nand U3205 (N_3205,N_2494,N_1902);
nor U3206 (N_3206,N_23,N_2147);
nor U3207 (N_3207,N_461,N_811);
xor U3208 (N_3208,N_1923,N_1514);
and U3209 (N_3209,N_300,N_1120);
or U3210 (N_3210,N_2829,N_917);
and U3211 (N_3211,N_2547,N_1991);
nor U3212 (N_3212,N_1859,N_1291);
and U3213 (N_3213,N_916,N_143);
and U3214 (N_3214,N_1641,N_1397);
nand U3215 (N_3215,N_1075,N_1393);
nand U3216 (N_3216,N_1416,N_512);
and U3217 (N_3217,N_808,N_651);
nor U3218 (N_3218,N_1949,N_2570);
and U3219 (N_3219,N_240,N_971);
and U3220 (N_3220,N_1169,N_2910);
nor U3221 (N_3221,N_2363,N_1024);
or U3222 (N_3222,N_1026,N_211);
and U3223 (N_3223,N_1600,N_2619);
and U3224 (N_3224,N_2565,N_292);
or U3225 (N_3225,N_1895,N_2015);
nand U3226 (N_3226,N_586,N_967);
or U3227 (N_3227,N_93,N_1293);
and U3228 (N_3228,N_2134,N_328);
and U3229 (N_3229,N_1852,N_336);
or U3230 (N_3230,N_988,N_2748);
or U3231 (N_3231,N_86,N_2279);
nand U3232 (N_3232,N_648,N_1996);
or U3233 (N_3233,N_537,N_2758);
nor U3234 (N_3234,N_2008,N_1578);
or U3235 (N_3235,N_1560,N_2048);
or U3236 (N_3236,N_2266,N_124);
and U3237 (N_3237,N_1302,N_1511);
and U3238 (N_3238,N_354,N_1967);
nor U3239 (N_3239,N_1968,N_822);
or U3240 (N_3240,N_168,N_72);
nand U3241 (N_3241,N_309,N_1019);
nand U3242 (N_3242,N_2826,N_2791);
nand U3243 (N_3243,N_2751,N_1848);
nand U3244 (N_3244,N_846,N_401);
and U3245 (N_3245,N_1155,N_15);
nand U3246 (N_3246,N_319,N_1766);
nand U3247 (N_3247,N_2698,N_1689);
and U3248 (N_3248,N_1016,N_2534);
or U3249 (N_3249,N_1347,N_2702);
nand U3250 (N_3250,N_1590,N_2248);
nor U3251 (N_3251,N_2635,N_2094);
and U3252 (N_3252,N_1493,N_1032);
nand U3253 (N_3253,N_834,N_1881);
xnor U3254 (N_3254,N_2461,N_976);
and U3255 (N_3255,N_281,N_568);
or U3256 (N_3256,N_1892,N_192);
and U3257 (N_3257,N_615,N_556);
and U3258 (N_3258,N_2766,N_1263);
nor U3259 (N_3259,N_2530,N_2108);
and U3260 (N_3260,N_148,N_2295);
and U3261 (N_3261,N_757,N_635);
and U3262 (N_3262,N_2173,N_1356);
nor U3263 (N_3263,N_1508,N_2164);
or U3264 (N_3264,N_2969,N_2390);
nor U3265 (N_3265,N_1536,N_2505);
nand U3266 (N_3266,N_330,N_1685);
xor U3267 (N_3267,N_2800,N_1874);
nor U3268 (N_3268,N_2054,N_1476);
xor U3269 (N_3269,N_2637,N_1448);
nand U3270 (N_3270,N_331,N_1420);
and U3271 (N_3271,N_1141,N_2992);
and U3272 (N_3272,N_500,N_2520);
and U3273 (N_3273,N_1402,N_1888);
or U3274 (N_3274,N_2802,N_621);
nand U3275 (N_3275,N_2216,N_953);
and U3276 (N_3276,N_358,N_2068);
nand U3277 (N_3277,N_2492,N_1827);
and U3278 (N_3278,N_378,N_2288);
or U3279 (N_3279,N_1171,N_1819);
and U3280 (N_3280,N_894,N_90);
nor U3281 (N_3281,N_1668,N_1821);
nand U3282 (N_3282,N_91,N_1663);
nand U3283 (N_3283,N_334,N_1250);
or U3284 (N_3284,N_73,N_1);
or U3285 (N_3285,N_2487,N_2481);
and U3286 (N_3286,N_1700,N_2287);
nand U3287 (N_3287,N_1228,N_630);
nor U3288 (N_3288,N_105,N_553);
nand U3289 (N_3289,N_1903,N_430);
nand U3290 (N_3290,N_873,N_262);
nor U3291 (N_3291,N_1449,N_1439);
or U3292 (N_3292,N_1808,N_1648);
nand U3293 (N_3293,N_2716,N_2719);
xor U3294 (N_3294,N_1910,N_2355);
nor U3295 (N_3295,N_2745,N_2059);
or U3296 (N_3296,N_75,N_1746);
and U3297 (N_3297,N_777,N_2017);
or U3298 (N_3298,N_2881,N_1833);
nand U3299 (N_3299,N_888,N_2431);
and U3300 (N_3300,N_2671,N_2093);
nand U3301 (N_3301,N_1657,N_2589);
nor U3302 (N_3302,N_346,N_2542);
and U3303 (N_3303,N_1613,N_1225);
or U3304 (N_3304,N_1886,N_1781);
or U3305 (N_3305,N_2250,N_1174);
or U3306 (N_3306,N_238,N_2364);
or U3307 (N_3307,N_783,N_215);
nand U3308 (N_3308,N_193,N_92);
or U3309 (N_3309,N_1615,N_899);
nor U3310 (N_3310,N_2418,N_1647);
and U3311 (N_3311,N_1212,N_302);
or U3312 (N_3312,N_2848,N_1445);
nand U3313 (N_3313,N_646,N_2314);
and U3314 (N_3314,N_244,N_2591);
and U3315 (N_3315,N_1256,N_157);
or U3316 (N_3316,N_2300,N_1463);
and U3317 (N_3317,N_946,N_2763);
nor U3318 (N_3318,N_2557,N_2592);
nor U3319 (N_3319,N_1583,N_403);
nand U3320 (N_3320,N_1344,N_2409);
nand U3321 (N_3321,N_2773,N_2771);
and U3322 (N_3322,N_195,N_411);
or U3323 (N_3323,N_1319,N_1995);
or U3324 (N_3324,N_258,N_2162);
and U3325 (N_3325,N_826,N_1209);
or U3326 (N_3326,N_2932,N_2935);
or U3327 (N_3327,N_2165,N_2581);
and U3328 (N_3328,N_2459,N_569);
or U3329 (N_3329,N_177,N_1734);
or U3330 (N_3330,N_595,N_1906);
or U3331 (N_3331,N_2704,N_2001);
and U3332 (N_3332,N_2496,N_1526);
nor U3333 (N_3333,N_2473,N_2009);
nand U3334 (N_3334,N_2896,N_1705);
nand U3335 (N_3335,N_167,N_2628);
nand U3336 (N_3336,N_2572,N_2395);
or U3337 (N_3337,N_1498,N_2269);
and U3338 (N_3338,N_591,N_1468);
nor U3339 (N_3339,N_314,N_2180);
nor U3340 (N_3340,N_735,N_1232);
nand U3341 (N_3341,N_1365,N_2133);
nor U3342 (N_3342,N_2000,N_2361);
nand U3343 (N_3343,N_2296,N_915);
nor U3344 (N_3344,N_1240,N_2382);
and U3345 (N_3345,N_482,N_2238);
or U3346 (N_3346,N_1460,N_802);
nor U3347 (N_3347,N_836,N_1070);
and U3348 (N_3348,N_526,N_2615);
or U3349 (N_3349,N_1799,N_2768);
nand U3350 (N_3350,N_2867,N_255);
nand U3351 (N_3351,N_88,N_2544);
and U3352 (N_3352,N_726,N_2044);
or U3353 (N_3353,N_1305,N_791);
or U3354 (N_3354,N_763,N_2835);
or U3355 (N_3355,N_2953,N_2833);
nand U3356 (N_3356,N_2086,N_1475);
nor U3357 (N_3357,N_1891,N_2778);
and U3358 (N_3358,N_495,N_229);
and U3359 (N_3359,N_922,N_2638);
nor U3360 (N_3360,N_2539,N_2304);
nand U3361 (N_3361,N_2075,N_2817);
and U3362 (N_3362,N_987,N_1287);
nand U3363 (N_3363,N_1741,N_1411);
nor U3364 (N_3364,N_371,N_74);
nand U3365 (N_3365,N_134,N_2998);
nor U3366 (N_3366,N_2131,N_2453);
nor U3367 (N_3367,N_2827,N_2976);
and U3368 (N_3368,N_474,N_1360);
nor U3369 (N_3369,N_2936,N_2200);
nand U3370 (N_3370,N_1274,N_2345);
or U3371 (N_3371,N_436,N_2987);
or U3372 (N_3372,N_1558,N_1117);
or U3373 (N_3373,N_1829,N_1593);
nor U3374 (N_3374,N_2729,N_1301);
or U3375 (N_3375,N_1851,N_2344);
or U3376 (N_3376,N_1831,N_2247);
nor U3377 (N_3377,N_1043,N_120);
and U3378 (N_3378,N_2490,N_1658);
nor U3379 (N_3379,N_1812,N_1328);
nor U3380 (N_3380,N_2241,N_1686);
or U3381 (N_3381,N_149,N_616);
nor U3382 (N_3382,N_573,N_1704);
and U3383 (N_3383,N_1129,N_2795);
nor U3384 (N_3384,N_1634,N_2902);
nand U3385 (N_3385,N_2649,N_2140);
nor U3386 (N_3386,N_1329,N_623);
and U3387 (N_3387,N_2518,N_1392);
and U3388 (N_3388,N_1181,N_542);
nor U3389 (N_3389,N_1144,N_2886);
nand U3390 (N_3390,N_1484,N_1928);
and U3391 (N_3391,N_1413,N_142);
or U3392 (N_3392,N_858,N_1048);
and U3393 (N_3393,N_365,N_1507);
or U3394 (N_3394,N_1150,N_2961);
or U3395 (N_3395,N_2107,N_950);
and U3396 (N_3396,N_2720,N_394);
nor U3397 (N_3397,N_2464,N_2297);
nand U3398 (N_3398,N_2340,N_2452);
nand U3399 (N_3399,N_1135,N_117);
and U3400 (N_3400,N_1950,N_715);
and U3401 (N_3401,N_1059,N_2739);
nor U3402 (N_3402,N_612,N_1364);
and U3403 (N_3403,N_876,N_1036);
nor U3404 (N_3404,N_2955,N_1285);
nor U3405 (N_3405,N_1056,N_642);
or U3406 (N_3406,N_1249,N_326);
or U3407 (N_3407,N_178,N_368);
nor U3408 (N_3408,N_582,N_584);
or U3409 (N_3409,N_1414,N_1029);
nand U3410 (N_3410,N_1544,N_1999);
nor U3411 (N_3411,N_1793,N_2184);
nand U3412 (N_3412,N_1853,N_427);
or U3413 (N_3413,N_2626,N_1002);
nand U3414 (N_3414,N_2721,N_2469);
or U3415 (N_3415,N_2166,N_2257);
nor U3416 (N_3416,N_536,N_805);
nand U3417 (N_3417,N_1660,N_1386);
or U3418 (N_3418,N_1719,N_2053);
nor U3419 (N_3419,N_1383,N_2952);
and U3420 (N_3420,N_1203,N_2488);
nand U3421 (N_3421,N_356,N_699);
or U3422 (N_3422,N_538,N_1031);
nor U3423 (N_3423,N_188,N_521);
or U3424 (N_3424,N_1373,N_1552);
or U3425 (N_3425,N_270,N_1084);
and U3426 (N_3426,N_2159,N_2625);
and U3427 (N_3427,N_579,N_643);
or U3428 (N_3428,N_1316,N_2981);
or U3429 (N_3429,N_2945,N_298);
and U3430 (N_3430,N_804,N_2810);
nand U3431 (N_3431,N_2972,N_2839);
and U3432 (N_3432,N_2824,N_1087);
or U3433 (N_3433,N_2400,N_2076);
nand U3434 (N_3434,N_1483,N_1102);
nor U3435 (N_3435,N_273,N_2997);
nand U3436 (N_3436,N_1623,N_357);
nor U3437 (N_3437,N_1528,N_2347);
or U3438 (N_3438,N_2387,N_1195);
nand U3439 (N_3439,N_2537,N_2310);
nor U3440 (N_3440,N_2609,N_566);
nor U3441 (N_3441,N_1735,N_2226);
and U3442 (N_3442,N_37,N_288);
nand U3443 (N_3443,N_1951,N_1535);
nor U3444 (N_3444,N_1098,N_711);
nand U3445 (N_3445,N_2622,N_1051);
or U3446 (N_3446,N_2668,N_1367);
nand U3447 (N_3447,N_2312,N_629);
xor U3448 (N_3448,N_997,N_2519);
and U3449 (N_3449,N_2512,N_1873);
nor U3450 (N_3450,N_1737,N_2175);
or U3451 (N_3451,N_284,N_795);
nand U3452 (N_3452,N_1178,N_1089);
and U3453 (N_3453,N_2203,N_498);
and U3454 (N_3454,N_996,N_1654);
and U3455 (N_3455,N_2273,N_1101);
xnor U3456 (N_3456,N_386,N_1533);
and U3457 (N_3457,N_1567,N_1666);
and U3458 (N_3458,N_2585,N_1118);
and U3459 (N_3459,N_1190,N_1947);
or U3460 (N_3460,N_1188,N_197);
or U3461 (N_3461,N_392,N_2365);
or U3462 (N_3462,N_2443,N_1309);
nor U3463 (N_3463,N_1269,N_471);
or U3464 (N_3464,N_1134,N_852);
nand U3465 (N_3465,N_611,N_1965);
or U3466 (N_3466,N_535,N_29);
nor U3467 (N_3467,N_692,N_1611);
and U3468 (N_3468,N_2258,N_1044);
nor U3469 (N_3469,N_17,N_2792);
and U3470 (N_3470,N_2457,N_1987);
and U3471 (N_3471,N_409,N_1027);
or U3472 (N_3472,N_1088,N_2422);
nor U3473 (N_3473,N_234,N_519);
nand U3474 (N_3474,N_2189,N_2521);
nor U3475 (N_3475,N_2383,N_2483);
nor U3476 (N_3476,N_2640,N_562);
nor U3477 (N_3477,N_935,N_1795);
or U3478 (N_3478,N_2568,N_2346);
nor U3479 (N_3479,N_1451,N_484);
nand U3480 (N_3480,N_2368,N_2003);
or U3481 (N_3481,N_1257,N_2261);
or U3482 (N_3482,N_658,N_2242);
and U3483 (N_3483,N_76,N_2909);
nor U3484 (N_3484,N_909,N_1674);
and U3485 (N_3485,N_515,N_2498);
nand U3486 (N_3486,N_1858,N_2412);
or U3487 (N_3487,N_1805,N_676);
xor U3488 (N_3488,N_116,N_1810);
nand U3489 (N_3489,N_2890,N_2104);
or U3490 (N_3490,N_2215,N_2513);
and U3491 (N_3491,N_109,N_2858);
nor U3492 (N_3492,N_57,N_2866);
nor U3493 (N_3493,N_1884,N_2212);
or U3494 (N_3494,N_2408,N_2417);
or U3495 (N_3495,N_2767,N_2073);
or U3496 (N_3496,N_2573,N_2553);
nor U3497 (N_3497,N_2903,N_2550);
nand U3498 (N_3498,N_373,N_2661);
nand U3499 (N_3499,N_2793,N_904);
nand U3500 (N_3500,N_1436,N_1885);
nand U3501 (N_3501,N_744,N_1350);
and U3502 (N_3502,N_248,N_2348);
nor U3503 (N_3503,N_1914,N_781);
and U3504 (N_3504,N_1880,N_548);
and U3505 (N_3505,N_1314,N_119);
or U3506 (N_3506,N_2564,N_627);
and U3507 (N_3507,N_1854,N_2072);
and U3508 (N_3508,N_2686,N_2179);
and U3509 (N_3509,N_693,N_21);
nor U3510 (N_3510,N_2924,N_1516);
and U3511 (N_3511,N_170,N_479);
nand U3512 (N_3512,N_1213,N_1266);
and U3513 (N_3513,N_1988,N_1455);
nor U3514 (N_3514,N_1222,N_849);
nand U3515 (N_3515,N_68,N_995);
and U3516 (N_3516,N_949,N_2081);
nor U3517 (N_3517,N_682,N_2301);
or U3518 (N_3518,N_191,N_2560);
or U3519 (N_3519,N_2580,N_481);
nand U3520 (N_3520,N_525,N_964);
and U3521 (N_3521,N_417,N_159);
and U3522 (N_3522,N_720,N_1342);
xor U3523 (N_3523,N_2085,N_2723);
and U3524 (N_3524,N_64,N_13);
and U3525 (N_3525,N_1149,N_2930);
nand U3526 (N_3526,N_2327,N_1481);
and U3527 (N_3527,N_79,N_83);
nand U3528 (N_3528,N_1845,N_1194);
or U3529 (N_3529,N_1417,N_2691);
and U3530 (N_3530,N_2750,N_649);
or U3531 (N_3531,N_121,N_2974);
nand U3532 (N_3532,N_1062,N_1284);
and U3533 (N_3533,N_2080,N_2141);
or U3534 (N_3534,N_182,N_1158);
and U3535 (N_3535,N_2219,N_1252);
nand U3536 (N_3536,N_1100,N_2970);
nand U3537 (N_3537,N_1519,N_1182);
and U3538 (N_3538,N_2373,N_2210);
or U3539 (N_3539,N_1248,N_1994);
nor U3540 (N_3540,N_2514,N_1045);
nand U3541 (N_3541,N_2045,N_1908);
nand U3542 (N_3542,N_58,N_2632);
or U3543 (N_3543,N_2764,N_2460);
nand U3544 (N_3544,N_2290,N_213);
nor U3545 (N_3545,N_2732,N_1006);
and U3546 (N_3546,N_2298,N_884);
or U3547 (N_3547,N_1530,N_1669);
nor U3548 (N_3548,N_565,N_1094);
and U3549 (N_3549,N_375,N_2706);
or U3550 (N_3550,N_1221,N_825);
nor U3551 (N_3551,N_599,N_1039);
and U3552 (N_3552,N_11,N_1446);
nor U3553 (N_3553,N_2244,N_1146);
and U3554 (N_3554,N_2883,N_717);
and U3555 (N_3555,N_1187,N_2034);
and U3556 (N_3556,N_268,N_2396);
nand U3557 (N_3557,N_98,N_2233);
and U3558 (N_3558,N_1198,N_130);
and U3559 (N_3559,N_674,N_2033);
nand U3560 (N_3560,N_2654,N_2427);
and U3561 (N_3561,N_2153,N_185);
and U3562 (N_3562,N_1022,N_874);
or U3563 (N_3563,N_2002,N_2436);
or U3564 (N_3564,N_2786,N_1049);
nor U3565 (N_3565,N_322,N_2779);
nor U3566 (N_3566,N_1792,N_1450);
or U3567 (N_3567,N_214,N_2420);
and U3568 (N_3568,N_1868,N_1014);
nor U3569 (N_3569,N_2898,N_2155);
or U3570 (N_3570,N_2249,N_2209);
nand U3571 (N_3571,N_264,N_2286);
nand U3572 (N_3572,N_228,N_2199);
and U3573 (N_3573,N_704,N_1706);
or U3574 (N_3574,N_2602,N_1325);
and U3575 (N_3575,N_1466,N_919);
nand U3576 (N_3576,N_885,N_1630);
nor U3577 (N_3577,N_572,N_1236);
nor U3578 (N_3578,N_1083,N_1412);
nand U3579 (N_3579,N_2814,N_2853);
nor U3580 (N_3580,N_1041,N_2389);
and U3581 (N_3581,N_2360,N_1864);
nand U3582 (N_3582,N_784,N_1355);
and U3583 (N_3583,N_2448,N_1421);
or U3584 (N_3584,N_2435,N_210);
or U3585 (N_3585,N_1082,N_1050);
and U3586 (N_3586,N_2776,N_2441);
and U3587 (N_3587,N_2523,N_2013);
or U3588 (N_3588,N_1277,N_1341);
nor U3589 (N_3589,N_2803,N_1241);
or U3590 (N_3590,N_1168,N_979);
nor U3591 (N_3591,N_1260,N_1961);
nand U3592 (N_3592,N_2062,N_785);
and U3593 (N_3593,N_813,N_466);
and U3594 (N_3594,N_180,N_2047);
or U3595 (N_3595,N_2820,N_2805);
and U3596 (N_3596,N_842,N_351);
or U3597 (N_3597,N_1953,N_5);
or U3598 (N_3598,N_2066,N_2709);
or U3599 (N_3599,N_560,N_1238);
and U3600 (N_3600,N_960,N_184);
nor U3601 (N_3601,N_2838,N_65);
nand U3602 (N_3602,N_423,N_103);
or U3603 (N_3603,N_1123,N_838);
or U3604 (N_3604,N_1964,N_452);
nand U3605 (N_3605,N_1261,N_2458);
and U3606 (N_3606,N_518,N_2846);
nor U3607 (N_3607,N_2681,N_10);
and U3608 (N_3608,N_1773,N_1140);
or U3609 (N_3609,N_819,N_1034);
nor U3610 (N_3610,N_1879,N_128);
and U3611 (N_3611,N_106,N_1612);
and U3612 (N_3612,N_345,N_235);
nor U3613 (N_3613,N_725,N_1116);
or U3614 (N_3614,N_2041,N_1564);
or U3615 (N_3615,N_110,N_2474);
nand U3616 (N_3616,N_2079,N_1984);
nand U3617 (N_3617,N_507,N_1797);
or U3618 (N_3618,N_47,N_818);
and U3619 (N_3619,N_2051,N_1760);
nand U3620 (N_3620,N_1843,N_1259);
or U3621 (N_3621,N_252,N_2574);
nor U3622 (N_3622,N_1755,N_2311);
nand U3623 (N_3623,N_2284,N_985);
nand U3624 (N_3624,N_2231,N_1707);
and U3625 (N_3625,N_154,N_99);
nor U3626 (N_3626,N_231,N_2816);
nor U3627 (N_3627,N_1547,N_1346);
nand U3628 (N_3628,N_533,N_2789);
or U3629 (N_3629,N_1432,N_402);
nand U3630 (N_3630,N_2566,N_112);
or U3631 (N_3631,N_2375,N_544);
and U3632 (N_3632,N_1731,N_728);
nand U3633 (N_3633,N_2963,N_1086);
and U3634 (N_3634,N_1697,N_1761);
nand U3635 (N_3635,N_2031,N_236);
and U3636 (N_3636,N_1610,N_1308);
nand U3637 (N_3637,N_1517,N_914);
nand U3638 (N_3638,N_695,N_212);
and U3639 (N_3639,N_1465,N_1307);
nor U3640 (N_3640,N_608,N_2738);
and U3641 (N_3641,N_2123,N_222);
nand U3642 (N_3642,N_256,N_1130);
nor U3643 (N_3643,N_1811,N_1370);
nor U3644 (N_3644,N_2634,N_1137);
nor U3645 (N_3645,N_2587,N_2479);
nand U3646 (N_3646,N_2959,N_415);
and U3647 (N_3647,N_2372,N_1176);
nand U3648 (N_3648,N_561,N_882);
nor U3649 (N_3649,N_2042,N_1005);
or U3650 (N_3650,N_1834,N_1113);
and U3651 (N_3651,N_1279,N_2);
nor U3652 (N_3652,N_1974,N_77);
and U3653 (N_3653,N_400,N_903);
nor U3654 (N_3654,N_1058,N_1579);
nor U3655 (N_3655,N_2774,N_202);
nor U3656 (N_3656,N_113,N_1440);
or U3657 (N_3657,N_739,N_200);
or U3658 (N_3658,N_1502,N_2307);
and U3659 (N_3659,N_1632,N_2501);
nand U3660 (N_3660,N_344,N_2507);
or U3661 (N_3661,N_2607,N_702);
and U3662 (N_3662,N_1716,N_1901);
nor U3663 (N_3663,N_738,N_324);
and U3664 (N_3664,N_1921,N_132);
or U3665 (N_3665,N_1061,N_1696);
nor U3666 (N_3666,N_2196,N_1067);
or U3667 (N_3667,N_297,N_39);
nand U3668 (N_3668,N_1926,N_1701);
and U3669 (N_3669,N_1015,N_1382);
or U3670 (N_3670,N_2021,N_869);
nor U3671 (N_3671,N_2235,N_102);
nor U3672 (N_3672,N_918,N_1433);
or U3673 (N_3673,N_1069,N_2251);
nor U3674 (N_3674,N_2888,N_1525);
and U3675 (N_3675,N_1817,N_934);
and U3676 (N_3676,N_217,N_1332);
nand U3677 (N_3677,N_1642,N_716);
or U3678 (N_3678,N_1504,N_1747);
nor U3679 (N_3679,N_2556,N_1423);
nor U3680 (N_3680,N_1969,N_1037);
or U3681 (N_3681,N_1667,N_1710);
nand U3682 (N_3682,N_2784,N_1231);
nand U3683 (N_3683,N_2978,N_1791);
xnor U3684 (N_3684,N_2274,N_2967);
nand U3685 (N_3685,N_1565,N_789);
nor U3686 (N_3686,N_2905,N_283);
or U3687 (N_3687,N_1932,N_1358);
and U3688 (N_3688,N_1471,N_675);
and U3689 (N_3689,N_1185,N_965);
nor U3690 (N_3690,N_1099,N_1907);
nor U3691 (N_3691,N_2983,N_454);
and U3692 (N_3692,N_1545,N_2915);
and U3693 (N_3693,N_510,N_442);
or U3694 (N_3694,N_1717,N_225);
or U3695 (N_3695,N_2957,N_1177);
and U3696 (N_3696,N_1431,N_2694);
nand U3697 (N_3697,N_444,N_844);
or U3698 (N_3698,N_2621,N_2119);
nor U3699 (N_3699,N_1830,N_2863);
nor U3700 (N_3700,N_1871,N_247);
nand U3701 (N_3701,N_1380,N_774);
and U3702 (N_3702,N_1981,N_898);
and U3703 (N_3703,N_347,N_1556);
or U3704 (N_3704,N_2354,N_1553);
or U3705 (N_3705,N_156,N_2907);
nand U3706 (N_3706,N_1167,N_1482);
nor U3707 (N_3707,N_1944,N_1013);
nor U3708 (N_3708,N_1399,N_1992);
nor U3709 (N_3709,N_2313,N_2191);
or U3710 (N_3710,N_456,N_705);
and U3711 (N_3711,N_1948,N_1142);
nand U3712 (N_3712,N_2949,N_1956);
or U3713 (N_3713,N_1505,N_2999);
and U3714 (N_3714,N_2176,N_396);
or U3715 (N_3715,N_1351,N_749);
or U3716 (N_3716,N_2315,N_2444);
and U3717 (N_3717,N_61,N_1649);
and U3718 (N_3718,N_1644,N_412);
nor U3719 (N_3719,N_278,N_2158);
and U3720 (N_3720,N_1550,N_1262);
nor U3721 (N_3721,N_2685,N_2900);
or U3722 (N_3722,N_2471,N_1244);
or U3723 (N_3723,N_532,N_2097);
xnor U3724 (N_3724,N_2908,N_1110);
nor U3725 (N_3725,N_1395,N_2018);
nor U3726 (N_3726,N_1352,N_2724);
or U3727 (N_3727,N_1721,N_718);
or U3728 (N_3728,N_2356,N_2639);
nor U3729 (N_3729,N_1197,N_753);
nor U3730 (N_3730,N_2939,N_756);
and U3731 (N_3731,N_952,N_285);
nand U3732 (N_3732,N_2120,N_729);
nand U3733 (N_3733,N_1330,N_370);
or U3734 (N_3734,N_2989,N_1333);
nor U3735 (N_3735,N_2925,N_743);
nor U3736 (N_3736,N_1023,N_158);
and U3737 (N_3737,N_1294,N_2911);
nor U3738 (N_3738,N_690,N_546);
or U3739 (N_3739,N_1624,N_1900);
nand U3740 (N_3740,N_2294,N_913);
and U3741 (N_3741,N_323,N_52);
and U3742 (N_3742,N_2058,N_111);
nor U3743 (N_3743,N_2177,N_613);
and U3744 (N_3744,N_1283,N_653);
nor U3745 (N_3745,N_340,N_2246);
or U3746 (N_3746,N_2938,N_1245);
or U3747 (N_3747,N_2703,N_1635);
or U3748 (N_3748,N_1861,N_385);
nor U3749 (N_3749,N_2472,N_1692);
or U3750 (N_3750,N_1489,N_2208);
nor U3751 (N_3751,N_905,N_600);
nor U3752 (N_3752,N_1281,N_2875);
nor U3753 (N_3753,N_272,N_2205);
or U3754 (N_3754,N_2065,N_1211);
and U3755 (N_3755,N_1204,N_2852);
or U3756 (N_3756,N_2064,N_1575);
nand U3757 (N_3757,N_1822,N_2323);
and U3758 (N_3758,N_104,N_307);
nor U3759 (N_3759,N_828,N_1172);
and U3760 (N_3760,N_1192,N_2926);
and U3761 (N_3761,N_2087,N_1499);
or U3762 (N_3762,N_2705,N_1754);
or U3763 (N_3763,N_2636,N_2575);
nand U3764 (N_3764,N_650,N_751);
or U3765 (N_3765,N_1983,N_927);
xnor U3766 (N_3766,N_2369,N_2082);
or U3767 (N_3767,N_520,N_2595);
and U3768 (N_3768,N_1816,N_2084);
and U3769 (N_3769,N_251,N_277);
nand U3770 (N_3770,N_2652,N_2005);
nand U3771 (N_3771,N_2710,N_1418);
nand U3772 (N_3772,N_2352,N_1828);
nand U3773 (N_3773,N_880,N_135);
and U3774 (N_3774,N_1555,N_1769);
or U3775 (N_3775,N_647,N_455);
nor U3776 (N_3776,N_100,N_639);
or U3777 (N_3777,N_380,N_661);
and U3778 (N_3778,N_2672,N_27);
or U3779 (N_3779,N_1699,N_957);
nor U3780 (N_3780,N_2780,N_2403);
and U3781 (N_3781,N_63,N_2916);
xor U3782 (N_3782,N_2263,N_2509);
nor U3783 (N_3783,N_2056,N_2679);
or U3784 (N_3784,N_798,N_1521);
nand U3785 (N_3785,N_1753,N_1682);
and U3786 (N_3786,N_1676,N_1963);
or U3787 (N_3787,N_2610,N_1419);
nand U3788 (N_3788,N_617,N_945);
nor U3789 (N_3789,N_2567,N_1035);
xor U3790 (N_3790,N_2195,N_2339);
or U3791 (N_3791,N_422,N_2206);
or U3792 (N_3792,N_2682,N_1860);
nand U3793 (N_3793,N_662,N_848);
nand U3794 (N_3794,N_803,N_451);
and U3795 (N_3795,N_511,N_2917);
nand U3796 (N_3796,N_221,N_1276);
nand U3797 (N_3797,N_1444,N_1943);
nor U3798 (N_3798,N_434,N_2787);
or U3799 (N_3799,N_1586,N_2442);
or U3800 (N_3800,N_446,N_631);
or U3801 (N_3801,N_2656,N_900);
or U3802 (N_3802,N_1608,N_2451);
nand U3803 (N_3803,N_776,N_1362);
and U3804 (N_3804,N_1779,N_1290);
and U3805 (N_3805,N_2759,N_2362);
nand U3806 (N_3806,N_605,N_685);
or U3807 (N_3807,N_859,N_745);
xor U3808 (N_3808,N_4,N_1518);
or U3809 (N_3809,N_2746,N_2285);
nor U3810 (N_3810,N_770,N_245);
or U3811 (N_3811,N_2217,N_2731);
or U3812 (N_3812,N_1904,N_1376);
or U3813 (N_3813,N_2576,N_796);
and U3814 (N_3814,N_2293,N_769);
nor U3815 (N_3815,N_2124,N_892);
and U3816 (N_3816,N_2897,N_1408);
nand U3817 (N_3817,N_475,N_194);
and U3818 (N_3818,N_82,N_2467);
or U3819 (N_3819,N_2524,N_1591);
and U3820 (N_3820,N_2880,N_989);
nor U3821 (N_3821,N_2605,N_1587);
or U3822 (N_3822,N_530,N_1640);
or U3823 (N_3823,N_673,N_2132);
and U3824 (N_3824,N_1814,N_172);
nand U3825 (N_3825,N_2741,N_655);
or U3826 (N_3826,N_1939,N_2713);
nand U3827 (N_3827,N_2725,N_1066);
and U3828 (N_3828,N_714,N_127);
nand U3829 (N_3829,N_1602,N_549);
or U3830 (N_3830,N_152,N_1359);
or U3831 (N_3831,N_2655,N_2597);
or U3832 (N_3832,N_147,N_1691);
nand U3833 (N_3833,N_133,N_126);
nand U3834 (N_3834,N_1226,N_2743);
nor U3835 (N_3835,N_59,N_999);
or U3836 (N_3836,N_223,N_1802);
nand U3837 (N_3837,N_1003,N_364);
and U3838 (N_3838,N_1157,N_2960);
nand U3839 (N_3839,N_1148,N_443);
nand U3840 (N_3840,N_2092,N_724);
and U3841 (N_3841,N_1976,N_1292);
and U3842 (N_3842,N_1220,N_2899);
or U3843 (N_3843,N_2933,N_2225);
nor U3844 (N_3844,N_118,N_2402);
nand U3845 (N_3845,N_2160,N_2423);
nor U3846 (N_3846,N_2326,N_2744);
nor U3847 (N_3847,N_2770,N_1820);
and U3848 (N_3848,N_2811,N_747);
and U3849 (N_3849,N_1732,N_1289);
and U3850 (N_3850,N_420,N_563);
or U3851 (N_3851,N_1855,N_1371);
and U3852 (N_3852,N_19,N_2845);
and U3853 (N_3853,N_2109,N_910);
nand U3854 (N_3854,N_1147,N_1905);
nor U3855 (N_3855,N_1599,N_1804);
and U3856 (N_3856,N_2887,N_1064);
nor U3857 (N_3857,N_2991,N_1338);
xnor U3858 (N_3858,N_2484,N_1052);
and U3859 (N_3859,N_1813,N_1645);
or U3860 (N_3860,N_2187,N_1520);
nor U3861 (N_3861,N_2370,N_1639);
nand U3862 (N_3862,N_1091,N_2071);
or U3863 (N_3863,N_1133,N_2415);
nand U3864 (N_3864,N_399,N_906);
nor U3865 (N_3865,N_289,N_1739);
and U3866 (N_3866,N_2980,N_1919);
nor U3867 (N_3867,N_1354,N_790);
nor U3868 (N_3868,N_1780,N_2985);
nor U3869 (N_3869,N_721,N_2475);
nor U3870 (N_3870,N_208,N_32);
and U3871 (N_3871,N_2708,N_267);
nor U3872 (N_3872,N_2993,N_1934);
and U3873 (N_3873,N_933,N_766);
nand U3874 (N_3874,N_2801,N_369);
and U3875 (N_3875,N_384,N_793);
and U3876 (N_3876,N_470,N_2411);
and U3877 (N_3877,N_457,N_1538);
or U3878 (N_3878,N_2854,N_467);
nor U3879 (N_3879,N_817,N_861);
or U3880 (N_3880,N_2439,N_663);
nor U3881 (N_3881,N_2061,N_2374);
nor U3882 (N_3882,N_1966,N_1401);
nand U3883 (N_3883,N_122,N_1835);
nor U3884 (N_3884,N_2799,N_592);
nand U3885 (N_3885,N_2871,N_2172);
or U3886 (N_3886,N_2877,N_2399);
or U3887 (N_3887,N_24,N_2036);
nor U3888 (N_3888,N_782,N_856);
and U3889 (N_3889,N_881,N_2577);
nand U3890 (N_3890,N_678,N_2099);
or U3891 (N_3891,N_2862,N_947);
or U3892 (N_3892,N_1430,N_688);
nor U3893 (N_3893,N_1164,N_2922);
nor U3894 (N_3894,N_2982,N_2535);
nand U3895 (N_3895,N_1154,N_970);
and U3896 (N_3896,N_2477,N_166);
nand U3897 (N_3897,N_2942,N_1515);
or U3898 (N_3898,N_2727,N_1929);
and U3899 (N_3899,N_2275,N_1783);
and U3900 (N_3900,N_1679,N_1404);
and U3901 (N_3901,N_1403,N_2973);
nor U3902 (N_3902,N_2163,N_2653);
or U3903 (N_3903,N_22,N_97);
or U3904 (N_3904,N_348,N_1751);
or U3905 (N_3905,N_926,N_1242);
and U3906 (N_3906,N_2230,N_2893);
nand U3907 (N_3907,N_333,N_2822);
nand U3908 (N_3908,N_890,N_107);
nand U3909 (N_3909,N_2951,N_476);
and U3910 (N_3910,N_2070,N_1750);
or U3911 (N_3911,N_594,N_2601);
or U3912 (N_3912,N_1652,N_1218);
and U3913 (N_3913,N_1915,N_2359);
or U3914 (N_3914,N_2971,N_320);
and U3915 (N_3915,N_1924,N_1145);
or U3916 (N_3916,N_857,N_2808);
nor U3917 (N_3917,N_1106,N_837);
and U3918 (N_3918,N_666,N_709);
and U3919 (N_3919,N_382,N_1752);
nand U3920 (N_3920,N_1219,N_1296);
nand U3921 (N_3921,N_2223,N_923);
or U3922 (N_3922,N_2582,N_672);
or U3923 (N_3923,N_1883,N_1856);
or U3924 (N_3924,N_2271,N_2281);
nor U3925 (N_3925,N_1650,N_951);
nor U3926 (N_3926,N_2529,N_2543);
or U3927 (N_3927,N_337,N_1562);
nand U3928 (N_3928,N_1542,N_2185);
nor U3929 (N_3929,N_2647,N_2665);
nor U3930 (N_3930,N_218,N_620);
nand U3931 (N_3931,N_1990,N_1288);
nor U3932 (N_3932,N_2631,N_1479);
nand U3933 (N_3933,N_2046,N_860);
and U3934 (N_3934,N_1912,N_1581);
and U3935 (N_3935,N_1008,N_349);
or U3936 (N_3936,N_1865,N_1962);
or U3937 (N_3937,N_2697,N_2678);
nor U3938 (N_3938,N_1713,N_1040);
and U3939 (N_3939,N_1646,N_516);
nand U3940 (N_3940,N_1742,N_1540);
or U3941 (N_3941,N_243,N_1424);
nor U3942 (N_3942,N_2014,N_1073);
nand U3943 (N_3943,N_1480,N_659);
and U3944 (N_3944,N_2765,N_868);
or U3945 (N_3945,N_2381,N_2074);
and U3946 (N_3946,N_1745,N_2220);
or U3947 (N_3947,N_2869,N_1215);
nand U3948 (N_3948,N_1935,N_2740);
nand U3949 (N_3949,N_405,N_2504);
nor U3950 (N_3950,N_404,N_366);
nor U3951 (N_3951,N_38,N_2425);
nand U3952 (N_3952,N_1318,N_812);
nor U3953 (N_3953,N_1572,N_1175);
and U3954 (N_3954,N_1636,N_1975);
and U3955 (N_3955,N_1317,N_2588);
or U3956 (N_3956,N_1495,N_1911);
nor U3957 (N_3957,N_114,N_583);
and U3958 (N_3958,N_664,N_1622);
and U3959 (N_3959,N_2478,N_1443);
nor U3960 (N_3960,N_1097,N_1004);
nand U3961 (N_3961,N_2463,N_559);
or U3962 (N_3962,N_2445,N_139);
or U3963 (N_3963,N_1396,N_308);
nand U3964 (N_3964,N_2357,N_1729);
and U3965 (N_3965,N_2237,N_280);
and U3966 (N_3966,N_506,N_95);
or U3967 (N_3967,N_2859,N_570);
or U3968 (N_3968,N_424,N_1104);
and U3969 (N_3969,N_854,N_469);
nand U3970 (N_3970,N_2830,N_722);
or U3971 (N_3971,N_1025,N_602);
or U3972 (N_3972,N_554,N_601);
or U3973 (N_3973,N_1163,N_1815);
nand U3974 (N_3974,N_746,N_1577);
nand U3975 (N_3975,N_707,N_2608);
and U3976 (N_3976,N_619,N_2349);
nor U3977 (N_3977,N_814,N_1486);
and U3978 (N_3978,N_431,N_984);
nor U3979 (N_3979,N_983,N_2186);
nand U3980 (N_3980,N_973,N_986);
and U3981 (N_3981,N_2885,N_2101);
and U3982 (N_3982,N_1878,N_2112);
nor U3983 (N_3983,N_2116,N_1092);
nor U3984 (N_3984,N_1310,N_1166);
nor U3985 (N_3985,N_1796,N_669);
and U3986 (N_3986,N_440,N_2167);
nand U3987 (N_3987,N_1509,N_1459);
nor U3988 (N_3988,N_2447,N_2687);
nor U3989 (N_3989,N_2760,N_1979);
and U3990 (N_3990,N_2188,N_1125);
or U3991 (N_3991,N_1807,N_51);
and U3992 (N_3992,N_2562,N_253);
or U3993 (N_3993,N_209,N_1917);
nand U3994 (N_3994,N_1989,N_1913);
nand U3995 (N_3995,N_1875,N_162);
nand U3996 (N_3996,N_1733,N_750);
nand U3997 (N_3997,N_306,N_1053);
nand U3998 (N_3998,N_1428,N_1076);
and U3999 (N_3999,N_787,N_832);
or U4000 (N_4000,N_6,N_2688);
and U4001 (N_4001,N_1407,N_1389);
nand U4002 (N_4002,N_1267,N_877);
and U4003 (N_4003,N_800,N_360);
nor U4004 (N_4004,N_867,N_527);
nor U4005 (N_4005,N_1126,N_2078);
or U4006 (N_4006,N_418,N_809);
nand U4007 (N_4007,N_286,N_46);
and U4008 (N_4008,N_1072,N_2069);
nand U4009 (N_4009,N_1112,N_179);
or U4010 (N_4010,N_48,N_2693);
nand U4011 (N_4011,N_1060,N_2879);
or U4012 (N_4012,N_2035,N_2775);
or U4013 (N_4013,N_2462,N_2096);
nand U4014 (N_4014,N_1278,N_2252);
nand U4015 (N_4015,N_1559,N_719);
nor U4016 (N_4016,N_165,N_908);
nand U4017 (N_4017,N_2690,N_2528);
nor U4018 (N_4018,N_1033,N_2392);
or U4019 (N_4019,N_2351,N_2692);
nor U4020 (N_4020,N_2990,N_2906);
and U4021 (N_4021,N_2405,N_2114);
nor U4022 (N_4022,N_1180,N_1300);
and U4023 (N_4023,N_2338,N_2122);
nand U4024 (N_4024,N_2532,N_1933);
and U4025 (N_4025,N_883,N_778);
and U4026 (N_4026,N_2117,N_2371);
and U4027 (N_4027,N_2282,N_1673);
nor U4028 (N_4028,N_2103,N_2569);
and U4029 (N_4029,N_1653,N_2837);
or U4030 (N_4030,N_453,N_327);
nor U4031 (N_4031,N_1777,N_2004);
nor U4032 (N_4032,N_767,N_361);
nand U4033 (N_4033,N_1038,N_2754);
or U4034 (N_4034,N_1487,N_1726);
or U4035 (N_4035,N_1457,N_1017);
and U4036 (N_4036,N_2506,N_2646);
nor U4037 (N_4037,N_701,N_1940);
nor U4038 (N_4038,N_1065,N_432);
and U4039 (N_4039,N_932,N_2753);
nor U4040 (N_4040,N_1010,N_1603);
and U4041 (N_4041,N_499,N_821);
or U4042 (N_4042,N_1594,N_1825);
nand U4043 (N_4043,N_936,N_2920);
or U4044 (N_4044,N_1237,N_1945);
or U4045 (N_4045,N_2255,N_925);
or U4046 (N_4046,N_2198,N_994);
and U4047 (N_4047,N_1368,N_845);
and U4048 (N_4048,N_2525,N_1824);
nor U4049 (N_4049,N_862,N_2026);
nor U4050 (N_4050,N_2868,N_311);
nand U4051 (N_4051,N_2536,N_123);
nand U4052 (N_4052,N_1744,N_1079);
nor U4053 (N_4053,N_610,N_551);
nor U4054 (N_4054,N_2121,N_85);
or U4055 (N_4055,N_2144,N_1627);
nand U4056 (N_4056,N_524,N_16);
nand U4057 (N_4057,N_169,N_1784);
or U4058 (N_4058,N_390,N_1569);
nor U4059 (N_4059,N_2860,N_761);
nand U4060 (N_4060,N_2715,N_1889);
nor U4061 (N_4061,N_1374,N_1028);
nand U4062 (N_4062,N_1757,N_472);
and U4063 (N_4063,N_609,N_2937);
and U4064 (N_4064,N_1152,N_2332);
and U4065 (N_4065,N_1109,N_618);
and U4066 (N_4066,N_55,N_1958);
nor U4067 (N_4067,N_175,N_1375);
nor U4068 (N_4068,N_2923,N_2476);
nor U4069 (N_4069,N_2019,N_1189);
nand U4070 (N_4070,N_2612,N_448);
nor U4071 (N_4071,N_463,N_539);
and U4072 (N_4072,N_260,N_2454);
and U4073 (N_4073,N_505,N_992);
nand U4074 (N_4074,N_144,N_181);
nor U4075 (N_4075,N_2253,N_1345);
and U4076 (N_4076,N_1510,N_1531);
and U4077 (N_4077,N_2222,N_2308);
and U4078 (N_4078,N_1162,N_2962);
nor U4079 (N_4079,N_216,N_2324);
and U4080 (N_4080,N_489,N_2380);
nor U4081 (N_4081,N_2278,N_2662);
nor U4082 (N_4082,N_1246,N_2674);
and U4083 (N_4083,N_2022,N_413);
nor U4084 (N_4084,N_2398,N_641);
nand U4085 (N_4085,N_1790,N_1223);
nand U4086 (N_4086,N_1379,N_89);
nand U4087 (N_4087,N_752,N_931);
and U4088 (N_4088,N_1782,N_2150);
nor U4089 (N_4089,N_2428,N_276);
and U4090 (N_4090,N_2028,N_414);
nand U4091 (N_4091,N_2037,N_1229);
and U4092 (N_4092,N_2864,N_978);
or U4093 (N_4093,N_1651,N_2620);
and U4094 (N_4094,N_2302,N_1916);
nor U4095 (N_4095,N_1725,N_508);
nor U4096 (N_4096,N_2806,N_1570);
or U4097 (N_4097,N_1708,N_30);
and U4098 (N_4098,N_2510,N_1541);
nor U4099 (N_4099,N_577,N_1336);
and U4100 (N_4100,N_764,N_1838);
nor U4101 (N_4101,N_998,N_1268);
nor U4102 (N_4102,N_2495,N_1115);
or U4103 (N_4103,N_2664,N_1199);
or U4104 (N_4104,N_2975,N_1136);
nand U4105 (N_4105,N_2842,N_1063);
and U4106 (N_4106,N_2115,N_2517);
nand U4107 (N_4107,N_2491,N_2211);
and U4108 (N_4108,N_190,N_1606);
and U4109 (N_4109,N_1738,N_2614);
nand U4110 (N_4110,N_2796,N_2919);
nand U4111 (N_4111,N_962,N_824);
nor U4112 (N_4112,N_389,N_41);
nor U4113 (N_4113,N_1702,N_755);
nor U4114 (N_4114,N_574,N_2870);
or U4115 (N_4115,N_342,N_956);
xor U4116 (N_4116,N_2192,N_1153);
nor U4117 (N_4117,N_2040,N_2736);
or U4118 (N_4118,N_1537,N_2593);
and U4119 (N_4119,N_942,N_2841);
or U4120 (N_4120,N_2170,N_35);
and U4121 (N_4121,N_1490,N_799);
or U4122 (N_4122,N_993,N_625);
nor U4123 (N_4123,N_56,N_1206);
or U4124 (N_4124,N_1139,N_2270);
and U4125 (N_4125,N_2777,N_2276);
nand U4126 (N_4126,N_593,N_1638);
nand U4127 (N_4127,N_2797,N_645);
and U4128 (N_4128,N_1312,N_2407);
and U4129 (N_4129,N_2011,N_2559);
or U4130 (N_4130,N_2812,N_727);
nor U4131 (N_4131,N_310,N_1315);
nor U4132 (N_4132,N_2934,N_1253);
or U4133 (N_4133,N_2511,N_352);
or U4134 (N_4134,N_176,N_2540);
or U4135 (N_4135,N_2280,N_683);
or U4136 (N_4136,N_445,N_2227);
or U4137 (N_4137,N_552,N_1513);
nand U4138 (N_4138,N_2157,N_2337);
or U4139 (N_4139,N_541,N_2499);
and U4140 (N_4140,N_233,N_1589);
or U4141 (N_4141,N_54,N_974);
or U4142 (N_4142,N_295,N_2193);
nor U4143 (N_4143,N_1214,N_2683);
and U4144 (N_4144,N_408,N_700);
nor U4145 (N_4145,N_2358,N_2563);
and U4146 (N_4146,N_2651,N_1598);
nand U4147 (N_4147,N_1477,N_2221);
nand U4148 (N_4148,N_2077,N_2336);
and U4149 (N_4149,N_1009,N_2410);
nor U4150 (N_4150,N_2277,N_628);
and U4151 (N_4151,N_387,N_1619);
xor U4152 (N_4152,N_2722,N_2419);
and U4153 (N_4153,N_2110,N_2531);
or U4154 (N_4154,N_146,N_680);
nand U4155 (N_4155,N_823,N_2050);
nor U4156 (N_4156,N_501,N_140);
and U4157 (N_4157,N_980,N_797);
nor U4158 (N_4158,N_291,N_1837);
or U4159 (N_4159,N_2234,N_2772);
nand U4160 (N_4160,N_125,N_2689);
and U4161 (N_4161,N_737,N_2813);
nor U4162 (N_4162,N_2666,N_2259);
nor U4163 (N_4163,N_2931,N_1306);
nand U4164 (N_4164,N_1986,N_1605);
or U4165 (N_4165,N_2755,N_1331);
nor U4166 (N_4166,N_820,N_2265);
nor U4167 (N_4167,N_45,N_227);
and U4168 (N_4168,N_1343,N_1922);
nor U4169 (N_4169,N_2446,N_1422);
or U4170 (N_4170,N_1954,N_2948);
xnor U4171 (N_4171,N_201,N_2707);
or U4172 (N_4172,N_2128,N_1534);
nor U4173 (N_4173,N_897,N_1931);
nor U4174 (N_4174,N_2680,N_2341);
or U4175 (N_4175,N_2927,N_929);
or U4176 (N_4176,N_2309,N_398);
nor U4177 (N_4177,N_1743,N_374);
or U4178 (N_4178,N_2701,N_2695);
and U4179 (N_4179,N_1224,N_2579);
or U4180 (N_4180,N_878,N_2039);
or U4181 (N_4181,N_1832,N_265);
nand U4182 (N_4182,N_706,N_1093);
or U4183 (N_4183,N_1523,N_2197);
nor U4184 (N_4184,N_2663,N_316);
nor U4185 (N_4185,N_1626,N_2913);
nand U4186 (N_4186,N_1672,N_2929);
and U4187 (N_4187,N_2456,N_388);
nand U4188 (N_4188,N_1774,N_1425);
nor U4189 (N_4189,N_1818,N_863);
or U4190 (N_4190,N_1151,N_355);
nor U4191 (N_4191,N_2804,N_955);
and U4192 (N_4192,N_2552,N_1601);
nor U4193 (N_4193,N_362,N_760);
and U4194 (N_4194,N_1918,N_670);
and U4195 (N_4195,N_2918,N_2367);
nor U4196 (N_4196,N_1047,N_2156);
nand U4197 (N_4197,N_480,N_1616);
nand U4198 (N_4198,N_1494,N_2485);
nor U4199 (N_4199,N_359,N_555);
nor U4200 (N_4200,N_2194,N_1789);
nor U4201 (N_4201,N_1794,N_891);
or U4202 (N_4202,N_433,N_1522);
nor U4203 (N_4203,N_1327,N_1529);
nand U4204 (N_4204,N_338,N_43);
and U4205 (N_4205,N_1369,N_242);
or U4206 (N_4206,N_2977,N_1930);
or U4207 (N_4207,N_428,N_2644);
or U4208 (N_4208,N_2586,N_2538);
and U4209 (N_4209,N_1326,N_1722);
nor U4210 (N_4210,N_343,N_2320);
and U4211 (N_4211,N_2876,N_1304);
and U4212 (N_4212,N_2465,N_847);
nor U4213 (N_4213,N_1582,N_2825);
or U4214 (N_4214,N_1625,N_1055);
or U4215 (N_4215,N_2201,N_2964);
and U4216 (N_4216,N_312,N_1415);
nand U4217 (N_4217,N_2267,N_1803);
and U4218 (N_4218,N_2781,N_2393);
and U4219 (N_4219,N_257,N_939);
nor U4220 (N_4220,N_2834,N_1973);
nand U4221 (N_4221,N_1512,N_968);
and U4222 (N_4222,N_145,N_2090);
and U4223 (N_4223,N_2145,N_363);
and U4224 (N_4224,N_1193,N_624);
nor U4225 (N_4225,N_603,N_1230);
or U4226 (N_4226,N_2214,N_2330);
nand U4227 (N_4227,N_241,N_654);
or U4228 (N_4228,N_1202,N_2292);
and U4229 (N_4229,N_2379,N_598);
and U4230 (N_4230,N_1549,N_335);
nor U4231 (N_4231,N_1840,N_1661);
or U4232 (N_4232,N_872,N_2100);
and U4233 (N_4233,N_1478,N_937);
and U4234 (N_4234,N_483,N_1938);
nand U4235 (N_4235,N_2561,N_2020);
or U4236 (N_4236,N_687,N_2350);
or U4237 (N_4237,N_2558,N_1942);
nand U4238 (N_4238,N_590,N_1670);
nand U4239 (N_4239,N_1233,N_290);
nand U4240 (N_4240,N_2321,N_597);
nand U4241 (N_4241,N_237,N_2291);
and U4242 (N_4242,N_2202,N_779);
nand U4243 (N_4243,N_943,N_1899);
nor U4244 (N_4244,N_954,N_1095);
and U4245 (N_4245,N_748,N_2761);
nor U4246 (N_4246,N_315,N_2947);
nand U4247 (N_4247,N_189,N_794);
nand U4248 (N_4248,N_1340,N_2629);
nand U4249 (N_4249,N_294,N_1119);
and U4250 (N_4250,N_462,N_1628);
nor U4251 (N_4251,N_67,N_2889);
xor U4252 (N_4252,N_640,N_1543);
nor U4253 (N_4253,N_2611,N_1823);
or U4254 (N_4254,N_1607,N_393);
or U4255 (N_4255,N_183,N_2616);
nand U4256 (N_4256,N_626,N_2264);
nand U4257 (N_4257,N_317,N_2470);
nor U4258 (N_4258,N_2526,N_1434);
xor U4259 (N_4259,N_1972,N_2333);
or U4260 (N_4260,N_49,N_1554);
nor U4261 (N_4261,N_2030,N_2232);
or U4262 (N_4262,N_2673,N_2151);
nor U4263 (N_4263,N_604,N_2130);
or U4264 (N_4264,N_1724,N_84);
and U4265 (N_4265,N_911,N_269);
nor U4266 (N_4266,N_274,N_1046);
and U4267 (N_4267,N_230,N_2733);
nor U4268 (N_4268,N_2260,N_2676);
nand U4269 (N_4269,N_1143,N_1090);
or U4270 (N_4270,N_1723,N_493);
or U4271 (N_4271,N_1909,N_540);
nor U4272 (N_4272,N_1385,N_2391);
and U4273 (N_4273,N_303,N_2894);
nor U4274 (N_4274,N_2424,N_1872);
and U4275 (N_4275,N_1078,N_1323);
xnor U4276 (N_4276,N_2388,N_2098);
nor U4277 (N_4277,N_1664,N_1337);
and U4278 (N_4278,N_2450,N_920);
nor U4279 (N_4279,N_9,N_2904);
nor U4280 (N_4280,N_1759,N_2590);
nor U4281 (N_4281,N_2384,N_2657);
nor U4282 (N_4282,N_1264,N_1551);
xor U4283 (N_4283,N_1748,N_2169);
nor U4284 (N_4284,N_1165,N_2440);
or U4285 (N_4285,N_2136,N_2545);
nor U4286 (N_4286,N_875,N_657);
nor U4287 (N_4287,N_733,N_1410);
and U4288 (N_4288,N_961,N_762);
and U4289 (N_4289,N_2728,N_889);
nor U4290 (N_4290,N_853,N_855);
nand U4291 (N_4291,N_1286,N_1927);
nor U4292 (N_4292,N_447,N_660);
or U4293 (N_4293,N_34,N_2416);
nor U4294 (N_4294,N_1890,N_622);
nand U4295 (N_4295,N_2137,N_2836);
nor U4296 (N_4296,N_589,N_198);
or U4297 (N_4297,N_2878,N_1665);
and U4298 (N_4298,N_2873,N_226);
and U4299 (N_4299,N_224,N_2489);
and U4300 (N_4300,N_2522,N_959);
and U4301 (N_4301,N_1107,N_2376);
or U4302 (N_4302,N_1127,N_502);
nor U4303 (N_4303,N_42,N_2769);
nand U4304 (N_4304,N_1339,N_2874);
or U4305 (N_4305,N_2594,N_2438);
nand U4306 (N_4306,N_325,N_671);
and U4307 (N_4307,N_1501,N_2466);
or U4308 (N_4308,N_1298,N_765);
or U4309 (N_4309,N_1030,N_31);
or U4310 (N_4310,N_775,N_1303);
nor U4311 (N_4311,N_1452,N_1736);
nand U4312 (N_4312,N_2366,N_2126);
or U4313 (N_4313,N_478,N_1576);
nand U4314 (N_4314,N_2643,N_204);
nand U4315 (N_4315,N_419,N_1863);
nand U4316 (N_4316,N_1887,N_696);
nand U4317 (N_4317,N_2502,N_1857);
nand U4318 (N_4318,N_786,N_205);
or U4319 (N_4319,N_810,N_395);
nand U4320 (N_4320,N_1335,N_1265);
or U4321 (N_4321,N_901,N_1085);
and U4322 (N_4322,N_2785,N_2006);
nand U4323 (N_4323,N_494,N_697);
and U4324 (N_4324,N_1488,N_2482);
and U4325 (N_4325,N_1131,N_2129);
and U4326 (N_4326,N_523,N_367);
nand U4327 (N_4327,N_2406,N_531);
nand U4328 (N_4328,N_36,N_1334);
nor U4329 (N_4329,N_703,N_129);
or U4330 (N_4330,N_2228,N_2325);
nand U4331 (N_4331,N_585,N_2303);
nor U4332 (N_4332,N_1714,N_439);
nand U4333 (N_4333,N_2319,N_490);
or U4334 (N_4334,N_2794,N_263);
nor U4335 (N_4335,N_1357,N_1472);
nor U4336 (N_4336,N_938,N_1313);
and U4337 (N_4337,N_1980,N_164);
or U4338 (N_4338,N_1977,N_841);
nand U4339 (N_4339,N_2757,N_81);
and U4340 (N_4340,N_2029,N_667);
or U4341 (N_4341,N_2551,N_2055);
nand U4342 (N_4342,N_1235,N_816);
or U4343 (N_4343,N_329,N_2600);
nand U4344 (N_4344,N_1321,N_734);
or U4345 (N_4345,N_948,N_1387);
or U4346 (N_4346,N_1273,N_1844);
and U4347 (N_4347,N_69,N_2353);
nand U4348 (N_4348,N_2762,N_1709);
and U4349 (N_4349,N_588,N_381);
nand U4350 (N_4350,N_2378,N_1662);
nor U4351 (N_4351,N_636,N_1251);
nor U4352 (N_4352,N_665,N_1846);
or U4353 (N_4353,N_2240,N_2752);
nand U4354 (N_4354,N_1170,N_1524);
nor U4355 (N_4355,N_174,N_1456);
or U4356 (N_4356,N_1592,N_1698);
and U4357 (N_4357,N_2010,N_1677);
and U4358 (N_4358,N_1438,N_1042);
nand U4359 (N_4359,N_299,N_1997);
nand U4360 (N_4360,N_1557,N_2726);
nand U4361 (N_4361,N_871,N_1546);
nand U4362 (N_4362,N_2146,N_1400);
nand U4363 (N_4363,N_2533,N_1693);
and U4364 (N_4364,N_1324,N_2497);
and U4365 (N_4365,N_557,N_1584);
nor U4366 (N_4366,N_771,N_2921);
and U4367 (N_4367,N_504,N_2171);
or U4368 (N_4368,N_1842,N_1485);
and U4369 (N_4369,N_1295,N_1186);
nor U4370 (N_4370,N_2113,N_893);
nor U4371 (N_4371,N_2807,N_1470);
or U4372 (N_4372,N_1809,N_1801);
or U4373 (N_4373,N_497,N_101);
nor U4374 (N_4374,N_1122,N_2658);
and U4375 (N_4375,N_1527,N_2599);
nor U4376 (N_4376,N_1406,N_2468);
and U4377 (N_4377,N_196,N_2052);
or U4378 (N_4378,N_1461,N_2437);
and U4379 (N_4379,N_7,N_441);
nand U4380 (N_4380,N_379,N_2844);
and U4381 (N_4381,N_930,N_301);
or U4382 (N_4382,N_773,N_2023);
and U4383 (N_4383,N_1320,N_2500);
nand U4384 (N_4384,N_895,N_2043);
and U4385 (N_4385,N_450,N_614);
nand U4386 (N_4386,N_2182,N_1270);
nor U4387 (N_4387,N_464,N_1681);
nand U4388 (N_4388,N_2328,N_740);
nand U4389 (N_4389,N_1621,N_62);
and U4390 (N_4390,N_1728,N_840);
nand U4391 (N_4391,N_2433,N_487);
nand U4392 (N_4392,N_2603,N_1978);
and U4393 (N_4393,N_171,N_2125);
nor U4394 (N_4394,N_558,N_2317);
xor U4395 (N_4395,N_488,N_1128);
or U4396 (N_4396,N_1715,N_1216);
xnor U4397 (N_4397,N_940,N_580);
and U4398 (N_4398,N_155,N_2988);
nand U4399 (N_4399,N_503,N_26);
nand U4400 (N_4400,N_835,N_780);
nand U4401 (N_4401,N_2954,N_2331);
and U4402 (N_4402,N_1394,N_1941);
nor U4403 (N_4403,N_576,N_963);
or U4404 (N_4404,N_1898,N_1850);
or U4405 (N_4405,N_2329,N_1936);
nor U4406 (N_4406,N_2236,N_2386);
xor U4407 (N_4407,N_435,N_1132);
or U4408 (N_4408,N_1867,N_2823);
or U4409 (N_4409,N_1749,N_2958);
nand U4410 (N_4410,N_70,N_2480);
nor U4411 (N_4411,N_1322,N_1405);
and U4412 (N_4412,N_1007,N_732);
nor U4413 (N_4413,N_2950,N_2088);
or U4414 (N_4414,N_991,N_981);
nor U4415 (N_4415,N_1021,N_1492);
or U4416 (N_4416,N_2996,N_1847);
and U4417 (N_4417,N_2024,N_1441);
nand U4418 (N_4418,N_1201,N_1243);
and U4419 (N_4419,N_1764,N_581);
nor U4420 (N_4420,N_1982,N_438);
and U4421 (N_4421,N_2749,N_2604);
or U4422 (N_4422,N_632,N_2747);
or U4423 (N_4423,N_1767,N_1937);
nor U4424 (N_4424,N_1184,N_2012);
xor U4425 (N_4425,N_1077,N_2584);
nor U4426 (N_4426,N_25,N_829);
nor U4427 (N_4427,N_2994,N_1561);
or U4428 (N_4428,N_850,N_1955);
nor U4429 (N_4429,N_2901,N_246);
or U4430 (N_4430,N_801,N_78);
or U4431 (N_4431,N_928,N_839);
nor U4432 (N_4432,N_2127,N_896);
and U4433 (N_4433,N_1849,N_465);
nor U4434 (N_4434,N_1711,N_571);
and U4435 (N_4435,N_2818,N_406);
or U4436 (N_4436,N_788,N_1081);
and U4437 (N_4437,N_2430,N_679);
or U4438 (N_4438,N_694,N_2660);
or U4439 (N_4439,N_2060,N_1349);
nor U4440 (N_4440,N_2578,N_522);
xnor U4441 (N_4441,N_689,N_376);
or U4442 (N_4442,N_1409,N_831);
and U4443 (N_4443,N_2342,N_1609);
or U4444 (N_4444,N_1620,N_150);
nor U4445 (N_4445,N_1012,N_2027);
nor U4446 (N_4446,N_1772,N_1124);
and U4447 (N_4447,N_2429,N_1539);
and U4448 (N_4448,N_2642,N_2598);
and U4449 (N_4449,N_160,N_1960);
or U4450 (N_4450,N_1618,N_2111);
or U4451 (N_4451,N_2699,N_141);
nand U4452 (N_4452,N_1280,N_2007);
and U4453 (N_4453,N_1353,N_2819);
nand U4454 (N_4454,N_2943,N_886);
and U4455 (N_4455,N_2840,N_741);
and U4456 (N_4456,N_279,N_1255);
nor U4457 (N_4457,N_686,N_53);
nand U4458 (N_4458,N_153,N_1426);
nor U4459 (N_4459,N_186,N_1671);
or U4460 (N_4460,N_2712,N_2790);
nand U4461 (N_4461,N_966,N_2049);
or U4462 (N_4462,N_2083,N_266);
and U4463 (N_4463,N_259,N_2855);
and U4464 (N_4464,N_2152,N_2815);
nand U4465 (N_4465,N_2891,N_426);
and U4466 (N_4466,N_2025,N_1839);
and U4467 (N_4467,N_1160,N_2730);
or U4468 (N_4468,N_468,N_2956);
nand U4469 (N_4469,N_1384,N_1720);
or U4470 (N_4470,N_575,N_851);
nor U4471 (N_4471,N_2148,N_0);
nand U4472 (N_4472,N_477,N_2711);
or U4473 (N_4473,N_1993,N_2229);
and U4474 (N_4474,N_2831,N_339);
and U4475 (N_4475,N_534,N_1462);
or U4476 (N_4476,N_1896,N_2118);
nor U4477 (N_4477,N_203,N_87);
nand U4478 (N_4478,N_115,N_1952);
or U4479 (N_4479,N_736,N_2756);
nor U4480 (N_4480,N_318,N_2213);
xor U4481 (N_4481,N_1442,N_2884);
and U4482 (N_4482,N_296,N_758);
nor U4483 (N_4483,N_1071,N_866);
and U4484 (N_4484,N_1841,N_416);
nor U4485 (N_4485,N_44,N_2245);
and U4486 (N_4486,N_2554,N_2174);
nand U4487 (N_4487,N_496,N_1121);
or U4488 (N_4488,N_2828,N_1631);
nand U4489 (N_4489,N_173,N_1437);
or U4490 (N_4490,N_1688,N_1675);
nand U4491 (N_4491,N_232,N_8);
nand U4492 (N_4492,N_1297,N_1363);
nor U4493 (N_4493,N_2659,N_2178);
and U4494 (N_4494,N_1447,N_1765);
and U4495 (N_4495,N_864,N_1054);
and U4496 (N_4496,N_545,N_827);
or U4497 (N_4497,N_1588,N_2106);
or U4498 (N_4498,N_2067,N_2861);
nand U4499 (N_4499,N_513,N_2218);
and U4500 (N_4500,N_2627,N_894);
or U4501 (N_4501,N_2484,N_1297);
nand U4502 (N_4502,N_1768,N_1783);
nand U4503 (N_4503,N_1716,N_777);
nand U4504 (N_4504,N_2227,N_339);
or U4505 (N_4505,N_1149,N_1942);
or U4506 (N_4506,N_1705,N_1386);
and U4507 (N_4507,N_847,N_1320);
or U4508 (N_4508,N_2006,N_441);
and U4509 (N_4509,N_2089,N_1385);
or U4510 (N_4510,N_2473,N_368);
or U4511 (N_4511,N_883,N_2645);
or U4512 (N_4512,N_2583,N_2557);
and U4513 (N_4513,N_2723,N_1919);
nand U4514 (N_4514,N_825,N_803);
or U4515 (N_4515,N_1468,N_802);
and U4516 (N_4516,N_933,N_534);
or U4517 (N_4517,N_2227,N_2566);
and U4518 (N_4518,N_2702,N_609);
nor U4519 (N_4519,N_2915,N_2218);
or U4520 (N_4520,N_2464,N_2225);
and U4521 (N_4521,N_2025,N_2393);
nand U4522 (N_4522,N_812,N_990);
nor U4523 (N_4523,N_107,N_1089);
nand U4524 (N_4524,N_2065,N_664);
and U4525 (N_4525,N_589,N_1980);
or U4526 (N_4526,N_2036,N_2427);
and U4527 (N_4527,N_1480,N_2195);
nor U4528 (N_4528,N_2513,N_2923);
nand U4529 (N_4529,N_81,N_393);
and U4530 (N_4530,N_1333,N_631);
or U4531 (N_4531,N_1416,N_1651);
and U4532 (N_4532,N_2739,N_2581);
or U4533 (N_4533,N_130,N_206);
nand U4534 (N_4534,N_2669,N_2567);
nand U4535 (N_4535,N_2184,N_1684);
nand U4536 (N_4536,N_1783,N_2937);
nor U4537 (N_4537,N_480,N_950);
nand U4538 (N_4538,N_36,N_379);
and U4539 (N_4539,N_309,N_1119);
or U4540 (N_4540,N_2844,N_1888);
or U4541 (N_4541,N_2402,N_779);
nand U4542 (N_4542,N_2117,N_218);
or U4543 (N_4543,N_2574,N_1701);
nor U4544 (N_4544,N_140,N_2280);
and U4545 (N_4545,N_1444,N_2597);
and U4546 (N_4546,N_1549,N_1262);
or U4547 (N_4547,N_820,N_2615);
or U4548 (N_4548,N_1312,N_2984);
nand U4549 (N_4549,N_2142,N_380);
nor U4550 (N_4550,N_985,N_226);
nor U4551 (N_4551,N_972,N_1539);
or U4552 (N_4552,N_1005,N_1070);
and U4553 (N_4553,N_139,N_418);
and U4554 (N_4554,N_1693,N_1103);
nor U4555 (N_4555,N_1114,N_2069);
or U4556 (N_4556,N_2430,N_2503);
nor U4557 (N_4557,N_977,N_1770);
nand U4558 (N_4558,N_2773,N_897);
nand U4559 (N_4559,N_1576,N_1507);
and U4560 (N_4560,N_2354,N_561);
nor U4561 (N_4561,N_103,N_1051);
or U4562 (N_4562,N_2126,N_1380);
nand U4563 (N_4563,N_2753,N_2272);
nor U4564 (N_4564,N_1520,N_1787);
nand U4565 (N_4565,N_1967,N_642);
and U4566 (N_4566,N_2580,N_1579);
nor U4567 (N_4567,N_515,N_686);
nand U4568 (N_4568,N_93,N_2687);
nor U4569 (N_4569,N_2116,N_1059);
and U4570 (N_4570,N_2930,N_1224);
and U4571 (N_4571,N_2866,N_1499);
or U4572 (N_4572,N_378,N_2148);
or U4573 (N_4573,N_1383,N_1854);
and U4574 (N_4574,N_894,N_2734);
and U4575 (N_4575,N_40,N_1572);
nand U4576 (N_4576,N_671,N_687);
nand U4577 (N_4577,N_1235,N_279);
and U4578 (N_4578,N_1290,N_1119);
nand U4579 (N_4579,N_2562,N_619);
or U4580 (N_4580,N_358,N_605);
or U4581 (N_4581,N_2874,N_2337);
nor U4582 (N_4582,N_2684,N_394);
nor U4583 (N_4583,N_1496,N_1159);
nor U4584 (N_4584,N_2728,N_958);
nor U4585 (N_4585,N_2238,N_703);
and U4586 (N_4586,N_2887,N_368);
and U4587 (N_4587,N_1105,N_1035);
nand U4588 (N_4588,N_2419,N_2822);
nand U4589 (N_4589,N_2172,N_46);
nand U4590 (N_4590,N_1880,N_188);
and U4591 (N_4591,N_1563,N_2520);
nand U4592 (N_4592,N_2142,N_1508);
or U4593 (N_4593,N_2115,N_2099);
and U4594 (N_4594,N_2731,N_1535);
and U4595 (N_4595,N_2397,N_28);
nand U4596 (N_4596,N_2415,N_2743);
or U4597 (N_4597,N_1633,N_587);
nor U4598 (N_4598,N_1838,N_2469);
and U4599 (N_4599,N_1508,N_1285);
nor U4600 (N_4600,N_2884,N_552);
nor U4601 (N_4601,N_1759,N_2922);
or U4602 (N_4602,N_448,N_489);
or U4603 (N_4603,N_1971,N_903);
nand U4604 (N_4604,N_629,N_266);
nand U4605 (N_4605,N_1164,N_2930);
or U4606 (N_4606,N_2909,N_352);
and U4607 (N_4607,N_2913,N_2091);
and U4608 (N_4608,N_2891,N_722);
nor U4609 (N_4609,N_749,N_1486);
and U4610 (N_4610,N_1733,N_755);
nor U4611 (N_4611,N_571,N_559);
or U4612 (N_4612,N_379,N_831);
and U4613 (N_4613,N_267,N_280);
nand U4614 (N_4614,N_2780,N_915);
and U4615 (N_4615,N_1014,N_1365);
or U4616 (N_4616,N_700,N_767);
and U4617 (N_4617,N_591,N_386);
nand U4618 (N_4618,N_1314,N_1040);
nor U4619 (N_4619,N_1357,N_2824);
or U4620 (N_4620,N_700,N_1077);
or U4621 (N_4621,N_938,N_1526);
nand U4622 (N_4622,N_2716,N_854);
nor U4623 (N_4623,N_496,N_783);
or U4624 (N_4624,N_2245,N_1393);
and U4625 (N_4625,N_2133,N_229);
nor U4626 (N_4626,N_2216,N_768);
and U4627 (N_4627,N_2668,N_2692);
or U4628 (N_4628,N_89,N_2695);
or U4629 (N_4629,N_217,N_1977);
and U4630 (N_4630,N_596,N_1702);
and U4631 (N_4631,N_776,N_770);
or U4632 (N_4632,N_1592,N_2277);
or U4633 (N_4633,N_1800,N_1509);
or U4634 (N_4634,N_598,N_2628);
nor U4635 (N_4635,N_2092,N_2808);
and U4636 (N_4636,N_419,N_1866);
nand U4637 (N_4637,N_1810,N_1442);
and U4638 (N_4638,N_1087,N_2759);
nor U4639 (N_4639,N_1450,N_1334);
nor U4640 (N_4640,N_380,N_1776);
and U4641 (N_4641,N_785,N_1995);
and U4642 (N_4642,N_99,N_1664);
or U4643 (N_4643,N_722,N_2828);
nand U4644 (N_4644,N_622,N_1812);
or U4645 (N_4645,N_1202,N_141);
nand U4646 (N_4646,N_324,N_1451);
or U4647 (N_4647,N_843,N_2925);
nand U4648 (N_4648,N_1326,N_710);
nand U4649 (N_4649,N_1177,N_1955);
or U4650 (N_4650,N_205,N_2992);
and U4651 (N_4651,N_2195,N_2832);
or U4652 (N_4652,N_1789,N_2106);
nor U4653 (N_4653,N_2297,N_995);
nand U4654 (N_4654,N_2856,N_2537);
and U4655 (N_4655,N_1054,N_1291);
or U4656 (N_4656,N_2375,N_1723);
and U4657 (N_4657,N_1059,N_2950);
nand U4658 (N_4658,N_1822,N_2992);
and U4659 (N_4659,N_2385,N_701);
or U4660 (N_4660,N_1612,N_1873);
nand U4661 (N_4661,N_2351,N_2685);
nand U4662 (N_4662,N_2652,N_1936);
or U4663 (N_4663,N_803,N_497);
and U4664 (N_4664,N_1995,N_1491);
or U4665 (N_4665,N_599,N_2982);
nand U4666 (N_4666,N_73,N_2744);
or U4667 (N_4667,N_1681,N_117);
or U4668 (N_4668,N_990,N_545);
or U4669 (N_4669,N_2470,N_2781);
nand U4670 (N_4670,N_1324,N_1823);
nand U4671 (N_4671,N_2061,N_2512);
and U4672 (N_4672,N_1289,N_935);
nor U4673 (N_4673,N_2772,N_1147);
nand U4674 (N_4674,N_282,N_734);
xor U4675 (N_4675,N_951,N_2213);
nor U4676 (N_4676,N_410,N_1626);
nor U4677 (N_4677,N_2458,N_208);
or U4678 (N_4678,N_1436,N_1797);
or U4679 (N_4679,N_306,N_914);
nand U4680 (N_4680,N_1073,N_349);
or U4681 (N_4681,N_2318,N_2499);
and U4682 (N_4682,N_2643,N_2432);
nor U4683 (N_4683,N_6,N_268);
nand U4684 (N_4684,N_2284,N_2738);
and U4685 (N_4685,N_701,N_268);
or U4686 (N_4686,N_2425,N_1987);
nand U4687 (N_4687,N_91,N_1052);
nor U4688 (N_4688,N_1965,N_970);
or U4689 (N_4689,N_1120,N_1852);
nand U4690 (N_4690,N_2141,N_1352);
and U4691 (N_4691,N_1706,N_2820);
nor U4692 (N_4692,N_616,N_2187);
nand U4693 (N_4693,N_527,N_445);
nor U4694 (N_4694,N_2447,N_2534);
nand U4695 (N_4695,N_2544,N_904);
or U4696 (N_4696,N_1670,N_874);
or U4697 (N_4697,N_1724,N_987);
nand U4698 (N_4698,N_1008,N_680);
nand U4699 (N_4699,N_425,N_2591);
and U4700 (N_4700,N_891,N_2971);
nand U4701 (N_4701,N_197,N_249);
nor U4702 (N_4702,N_2317,N_1416);
or U4703 (N_4703,N_2131,N_325);
nor U4704 (N_4704,N_2287,N_1476);
and U4705 (N_4705,N_1442,N_7);
nand U4706 (N_4706,N_2589,N_2106);
nor U4707 (N_4707,N_2065,N_2384);
and U4708 (N_4708,N_1359,N_2192);
or U4709 (N_4709,N_11,N_16);
or U4710 (N_4710,N_402,N_1745);
nand U4711 (N_4711,N_1144,N_629);
nand U4712 (N_4712,N_1726,N_539);
nand U4713 (N_4713,N_2779,N_2265);
or U4714 (N_4714,N_1891,N_692);
or U4715 (N_4715,N_2735,N_34);
nand U4716 (N_4716,N_2201,N_2348);
nor U4717 (N_4717,N_1137,N_461);
or U4718 (N_4718,N_2140,N_1976);
nor U4719 (N_4719,N_1870,N_459);
and U4720 (N_4720,N_1716,N_2919);
nor U4721 (N_4721,N_1329,N_2830);
nor U4722 (N_4722,N_1651,N_392);
nand U4723 (N_4723,N_674,N_609);
and U4724 (N_4724,N_2173,N_150);
nor U4725 (N_4725,N_822,N_2548);
or U4726 (N_4726,N_1475,N_1483);
nor U4727 (N_4727,N_1008,N_1430);
or U4728 (N_4728,N_2618,N_949);
and U4729 (N_4729,N_658,N_1838);
or U4730 (N_4730,N_716,N_2294);
and U4731 (N_4731,N_2359,N_2766);
and U4732 (N_4732,N_1544,N_1099);
and U4733 (N_4733,N_2230,N_1492);
and U4734 (N_4734,N_2086,N_512);
nor U4735 (N_4735,N_1151,N_2678);
or U4736 (N_4736,N_2119,N_445);
nand U4737 (N_4737,N_1579,N_1878);
nor U4738 (N_4738,N_2808,N_2543);
nor U4739 (N_4739,N_2189,N_427);
or U4740 (N_4740,N_1716,N_197);
nor U4741 (N_4741,N_2072,N_2471);
nand U4742 (N_4742,N_564,N_1409);
and U4743 (N_4743,N_235,N_712);
nand U4744 (N_4744,N_2003,N_91);
or U4745 (N_4745,N_188,N_960);
nand U4746 (N_4746,N_1435,N_279);
nand U4747 (N_4747,N_548,N_150);
nor U4748 (N_4748,N_1699,N_1630);
nand U4749 (N_4749,N_2230,N_1759);
nand U4750 (N_4750,N_1783,N_1521);
nor U4751 (N_4751,N_2550,N_2595);
nor U4752 (N_4752,N_1727,N_2129);
or U4753 (N_4753,N_1236,N_1063);
nand U4754 (N_4754,N_1487,N_2620);
or U4755 (N_4755,N_2015,N_2102);
nor U4756 (N_4756,N_610,N_1301);
and U4757 (N_4757,N_6,N_2126);
nor U4758 (N_4758,N_904,N_2151);
or U4759 (N_4759,N_1747,N_472);
and U4760 (N_4760,N_1242,N_2545);
and U4761 (N_4761,N_1799,N_2453);
and U4762 (N_4762,N_2009,N_41);
or U4763 (N_4763,N_1353,N_1254);
xor U4764 (N_4764,N_1656,N_2554);
nor U4765 (N_4765,N_2782,N_2322);
or U4766 (N_4766,N_1153,N_200);
and U4767 (N_4767,N_912,N_175);
and U4768 (N_4768,N_1651,N_461);
and U4769 (N_4769,N_624,N_2279);
or U4770 (N_4770,N_1542,N_1393);
nand U4771 (N_4771,N_658,N_2441);
and U4772 (N_4772,N_103,N_2954);
nor U4773 (N_4773,N_1105,N_665);
nor U4774 (N_4774,N_750,N_1501);
or U4775 (N_4775,N_2333,N_309);
or U4776 (N_4776,N_1847,N_2990);
nor U4777 (N_4777,N_1722,N_436);
nand U4778 (N_4778,N_1914,N_2035);
nor U4779 (N_4779,N_2468,N_2153);
nand U4780 (N_4780,N_753,N_411);
nor U4781 (N_4781,N_1075,N_1407);
nand U4782 (N_4782,N_1980,N_2055);
or U4783 (N_4783,N_1588,N_1141);
nor U4784 (N_4784,N_209,N_22);
nand U4785 (N_4785,N_2383,N_2951);
nor U4786 (N_4786,N_2116,N_416);
nor U4787 (N_4787,N_650,N_2702);
nor U4788 (N_4788,N_411,N_313);
and U4789 (N_4789,N_1603,N_799);
nor U4790 (N_4790,N_2080,N_2883);
nor U4791 (N_4791,N_1307,N_969);
and U4792 (N_4792,N_2726,N_163);
nand U4793 (N_4793,N_645,N_304);
nor U4794 (N_4794,N_319,N_375);
and U4795 (N_4795,N_1027,N_865);
and U4796 (N_4796,N_795,N_1004);
nand U4797 (N_4797,N_711,N_2368);
or U4798 (N_4798,N_353,N_935);
nor U4799 (N_4799,N_2094,N_803);
nand U4800 (N_4800,N_374,N_2115);
nor U4801 (N_4801,N_552,N_1293);
nand U4802 (N_4802,N_2482,N_747);
and U4803 (N_4803,N_210,N_324);
nand U4804 (N_4804,N_634,N_1625);
or U4805 (N_4805,N_999,N_2064);
or U4806 (N_4806,N_607,N_1025);
or U4807 (N_4807,N_2620,N_2723);
nor U4808 (N_4808,N_2511,N_1659);
nand U4809 (N_4809,N_2474,N_2560);
and U4810 (N_4810,N_2718,N_44);
nand U4811 (N_4811,N_716,N_2387);
nand U4812 (N_4812,N_693,N_2678);
nand U4813 (N_4813,N_2020,N_1594);
nand U4814 (N_4814,N_2350,N_1032);
and U4815 (N_4815,N_487,N_1860);
nand U4816 (N_4816,N_2356,N_1921);
nand U4817 (N_4817,N_1791,N_258);
nand U4818 (N_4818,N_1030,N_1900);
nor U4819 (N_4819,N_2707,N_1665);
nand U4820 (N_4820,N_2025,N_2665);
and U4821 (N_4821,N_2688,N_1000);
or U4822 (N_4822,N_2026,N_2350);
and U4823 (N_4823,N_2375,N_2644);
and U4824 (N_4824,N_2703,N_2456);
nand U4825 (N_4825,N_2789,N_1667);
xor U4826 (N_4826,N_769,N_2832);
nor U4827 (N_4827,N_2452,N_181);
or U4828 (N_4828,N_689,N_1850);
nand U4829 (N_4829,N_1054,N_2272);
and U4830 (N_4830,N_733,N_337);
nand U4831 (N_4831,N_265,N_2560);
and U4832 (N_4832,N_1801,N_1120);
nand U4833 (N_4833,N_360,N_98);
nand U4834 (N_4834,N_2119,N_2845);
nor U4835 (N_4835,N_2797,N_895);
nor U4836 (N_4836,N_1334,N_2640);
nand U4837 (N_4837,N_1978,N_1519);
and U4838 (N_4838,N_1861,N_2777);
nor U4839 (N_4839,N_2701,N_106);
nor U4840 (N_4840,N_194,N_2800);
nand U4841 (N_4841,N_1569,N_2687);
or U4842 (N_4842,N_708,N_441);
and U4843 (N_4843,N_124,N_2691);
and U4844 (N_4844,N_2868,N_2134);
nor U4845 (N_4845,N_37,N_1299);
and U4846 (N_4846,N_881,N_1909);
nor U4847 (N_4847,N_1219,N_1381);
nor U4848 (N_4848,N_2903,N_2176);
and U4849 (N_4849,N_1668,N_233);
and U4850 (N_4850,N_2448,N_2240);
nand U4851 (N_4851,N_1811,N_2217);
nor U4852 (N_4852,N_2584,N_874);
and U4853 (N_4853,N_87,N_2270);
nand U4854 (N_4854,N_384,N_726);
or U4855 (N_4855,N_1144,N_586);
or U4856 (N_4856,N_1989,N_1435);
nand U4857 (N_4857,N_1465,N_1962);
and U4858 (N_4858,N_532,N_2449);
or U4859 (N_4859,N_1190,N_1460);
nand U4860 (N_4860,N_34,N_938);
nor U4861 (N_4861,N_1282,N_1798);
or U4862 (N_4862,N_2252,N_1005);
and U4863 (N_4863,N_928,N_1378);
nor U4864 (N_4864,N_331,N_1417);
nor U4865 (N_4865,N_2179,N_1811);
or U4866 (N_4866,N_2738,N_1535);
nand U4867 (N_4867,N_2851,N_555);
or U4868 (N_4868,N_1446,N_2684);
and U4869 (N_4869,N_1098,N_2937);
or U4870 (N_4870,N_1024,N_947);
nand U4871 (N_4871,N_2368,N_945);
or U4872 (N_4872,N_2047,N_2629);
and U4873 (N_4873,N_579,N_1163);
and U4874 (N_4874,N_2418,N_108);
nand U4875 (N_4875,N_597,N_15);
nor U4876 (N_4876,N_1324,N_998);
nor U4877 (N_4877,N_2403,N_1614);
or U4878 (N_4878,N_2147,N_1366);
nor U4879 (N_4879,N_1522,N_362);
nand U4880 (N_4880,N_1965,N_541);
nor U4881 (N_4881,N_2197,N_2908);
nor U4882 (N_4882,N_2303,N_1232);
and U4883 (N_4883,N_2693,N_2273);
or U4884 (N_4884,N_2924,N_1951);
or U4885 (N_4885,N_2860,N_1385);
and U4886 (N_4886,N_1658,N_2171);
nand U4887 (N_4887,N_1827,N_2783);
and U4888 (N_4888,N_1437,N_2470);
and U4889 (N_4889,N_1691,N_2561);
and U4890 (N_4890,N_2345,N_2856);
or U4891 (N_4891,N_1763,N_323);
nor U4892 (N_4892,N_1029,N_2531);
or U4893 (N_4893,N_2059,N_2365);
nor U4894 (N_4894,N_2110,N_2579);
or U4895 (N_4895,N_2692,N_48);
and U4896 (N_4896,N_218,N_2408);
or U4897 (N_4897,N_895,N_1085);
or U4898 (N_4898,N_2972,N_1893);
nand U4899 (N_4899,N_733,N_2651);
and U4900 (N_4900,N_2059,N_2556);
nor U4901 (N_4901,N_616,N_400);
xor U4902 (N_4902,N_1949,N_207);
and U4903 (N_4903,N_820,N_1097);
and U4904 (N_4904,N_722,N_2627);
or U4905 (N_4905,N_2166,N_2141);
or U4906 (N_4906,N_1025,N_1382);
xnor U4907 (N_4907,N_1735,N_1725);
and U4908 (N_4908,N_1844,N_2687);
and U4909 (N_4909,N_1288,N_1017);
and U4910 (N_4910,N_534,N_1803);
or U4911 (N_4911,N_931,N_2201);
and U4912 (N_4912,N_1039,N_2204);
or U4913 (N_4913,N_1890,N_631);
or U4914 (N_4914,N_2423,N_529);
or U4915 (N_4915,N_2362,N_1666);
nand U4916 (N_4916,N_2075,N_1847);
and U4917 (N_4917,N_510,N_2978);
nor U4918 (N_4918,N_2050,N_284);
and U4919 (N_4919,N_1395,N_22);
nor U4920 (N_4920,N_2912,N_1776);
nor U4921 (N_4921,N_1377,N_1819);
nand U4922 (N_4922,N_1328,N_1742);
nand U4923 (N_4923,N_1676,N_68);
nand U4924 (N_4924,N_2461,N_206);
and U4925 (N_4925,N_230,N_956);
and U4926 (N_4926,N_1778,N_634);
nor U4927 (N_4927,N_2719,N_2963);
nor U4928 (N_4928,N_521,N_2648);
nand U4929 (N_4929,N_687,N_2745);
and U4930 (N_4930,N_1695,N_2111);
nand U4931 (N_4931,N_2089,N_694);
and U4932 (N_4932,N_128,N_1586);
nor U4933 (N_4933,N_2259,N_1555);
nand U4934 (N_4934,N_609,N_131);
nor U4935 (N_4935,N_1101,N_951);
nand U4936 (N_4936,N_2976,N_1756);
and U4937 (N_4937,N_2590,N_565);
or U4938 (N_4938,N_2114,N_2793);
and U4939 (N_4939,N_2322,N_2379);
nor U4940 (N_4940,N_126,N_1492);
nand U4941 (N_4941,N_547,N_2023);
and U4942 (N_4942,N_601,N_770);
nand U4943 (N_4943,N_923,N_1721);
and U4944 (N_4944,N_202,N_2895);
nand U4945 (N_4945,N_1775,N_1063);
nand U4946 (N_4946,N_509,N_1446);
and U4947 (N_4947,N_2735,N_1285);
and U4948 (N_4948,N_2430,N_1910);
nor U4949 (N_4949,N_1262,N_2021);
nor U4950 (N_4950,N_1772,N_1478);
nand U4951 (N_4951,N_2600,N_1548);
nor U4952 (N_4952,N_308,N_2325);
nor U4953 (N_4953,N_841,N_787);
or U4954 (N_4954,N_25,N_1241);
or U4955 (N_4955,N_1496,N_2486);
nand U4956 (N_4956,N_2316,N_498);
nor U4957 (N_4957,N_791,N_2769);
nand U4958 (N_4958,N_295,N_1965);
nor U4959 (N_4959,N_1231,N_1716);
nand U4960 (N_4960,N_858,N_1055);
nor U4961 (N_4961,N_1022,N_2232);
nand U4962 (N_4962,N_1146,N_2595);
and U4963 (N_4963,N_2569,N_908);
and U4964 (N_4964,N_827,N_1529);
or U4965 (N_4965,N_2732,N_1846);
nand U4966 (N_4966,N_53,N_496);
or U4967 (N_4967,N_1848,N_2656);
or U4968 (N_4968,N_295,N_434);
nand U4969 (N_4969,N_414,N_2594);
nor U4970 (N_4970,N_2342,N_1801);
nand U4971 (N_4971,N_1687,N_2878);
nor U4972 (N_4972,N_332,N_1188);
or U4973 (N_4973,N_1056,N_355);
nor U4974 (N_4974,N_2451,N_2101);
and U4975 (N_4975,N_2246,N_1331);
nand U4976 (N_4976,N_765,N_1765);
and U4977 (N_4977,N_1431,N_1323);
or U4978 (N_4978,N_1106,N_768);
nor U4979 (N_4979,N_1520,N_2356);
nor U4980 (N_4980,N_2225,N_1085);
or U4981 (N_4981,N_1758,N_1731);
and U4982 (N_4982,N_309,N_2884);
xor U4983 (N_4983,N_758,N_190);
or U4984 (N_4984,N_362,N_1961);
nor U4985 (N_4985,N_137,N_2924);
xnor U4986 (N_4986,N_134,N_644);
and U4987 (N_4987,N_986,N_454);
or U4988 (N_4988,N_427,N_1823);
or U4989 (N_4989,N_370,N_2376);
or U4990 (N_4990,N_406,N_2059);
nand U4991 (N_4991,N_972,N_1050);
or U4992 (N_4992,N_938,N_2469);
nor U4993 (N_4993,N_2304,N_850);
or U4994 (N_4994,N_760,N_2996);
nor U4995 (N_4995,N_1156,N_892);
and U4996 (N_4996,N_988,N_768);
or U4997 (N_4997,N_1490,N_1720);
nand U4998 (N_4998,N_1685,N_2908);
or U4999 (N_4999,N_2858,N_2743);
nor U5000 (N_5000,N_1059,N_163);
xnor U5001 (N_5001,N_1798,N_2767);
nor U5002 (N_5002,N_2657,N_2630);
nor U5003 (N_5003,N_2155,N_432);
nor U5004 (N_5004,N_2842,N_2454);
and U5005 (N_5005,N_2806,N_2073);
nand U5006 (N_5006,N_2667,N_322);
and U5007 (N_5007,N_591,N_433);
nand U5008 (N_5008,N_225,N_1343);
or U5009 (N_5009,N_1598,N_1466);
nor U5010 (N_5010,N_121,N_2595);
nor U5011 (N_5011,N_1619,N_1322);
or U5012 (N_5012,N_2624,N_1022);
and U5013 (N_5013,N_2707,N_1446);
nor U5014 (N_5014,N_2136,N_2382);
or U5015 (N_5015,N_822,N_2208);
or U5016 (N_5016,N_2413,N_2751);
xor U5017 (N_5017,N_2613,N_2031);
or U5018 (N_5018,N_357,N_1423);
or U5019 (N_5019,N_2748,N_1030);
and U5020 (N_5020,N_592,N_584);
and U5021 (N_5021,N_2582,N_2875);
nor U5022 (N_5022,N_2984,N_2832);
or U5023 (N_5023,N_828,N_126);
nand U5024 (N_5024,N_1189,N_770);
nand U5025 (N_5025,N_2327,N_2541);
nand U5026 (N_5026,N_2815,N_1617);
nand U5027 (N_5027,N_564,N_180);
and U5028 (N_5028,N_203,N_2380);
nand U5029 (N_5029,N_947,N_1304);
and U5030 (N_5030,N_13,N_1224);
and U5031 (N_5031,N_1246,N_1771);
nor U5032 (N_5032,N_2253,N_1805);
or U5033 (N_5033,N_1813,N_1408);
or U5034 (N_5034,N_1175,N_1765);
or U5035 (N_5035,N_758,N_300);
or U5036 (N_5036,N_428,N_1948);
and U5037 (N_5037,N_211,N_2992);
and U5038 (N_5038,N_1888,N_556);
nand U5039 (N_5039,N_1443,N_1287);
and U5040 (N_5040,N_1845,N_2803);
and U5041 (N_5041,N_2670,N_320);
nand U5042 (N_5042,N_2476,N_2169);
nand U5043 (N_5043,N_1931,N_2390);
nor U5044 (N_5044,N_2497,N_1608);
nand U5045 (N_5045,N_1547,N_1044);
nand U5046 (N_5046,N_2616,N_904);
or U5047 (N_5047,N_862,N_10);
and U5048 (N_5048,N_121,N_1675);
nand U5049 (N_5049,N_1968,N_2280);
nor U5050 (N_5050,N_2907,N_2699);
nand U5051 (N_5051,N_631,N_1507);
nand U5052 (N_5052,N_2959,N_1898);
nand U5053 (N_5053,N_1243,N_2137);
or U5054 (N_5054,N_311,N_731);
or U5055 (N_5055,N_2877,N_1047);
and U5056 (N_5056,N_1110,N_2754);
and U5057 (N_5057,N_1689,N_2966);
nand U5058 (N_5058,N_1526,N_2612);
nor U5059 (N_5059,N_546,N_994);
nor U5060 (N_5060,N_2496,N_1493);
and U5061 (N_5061,N_135,N_2044);
and U5062 (N_5062,N_1625,N_2855);
nand U5063 (N_5063,N_2434,N_1814);
nand U5064 (N_5064,N_1771,N_1457);
and U5065 (N_5065,N_907,N_57);
nand U5066 (N_5066,N_175,N_116);
nand U5067 (N_5067,N_1411,N_2769);
nand U5068 (N_5068,N_1452,N_1044);
nand U5069 (N_5069,N_275,N_767);
nor U5070 (N_5070,N_597,N_2426);
nor U5071 (N_5071,N_329,N_2738);
or U5072 (N_5072,N_902,N_375);
nor U5073 (N_5073,N_1932,N_52);
or U5074 (N_5074,N_2771,N_2656);
and U5075 (N_5075,N_1153,N_2876);
nand U5076 (N_5076,N_1825,N_612);
or U5077 (N_5077,N_1869,N_904);
and U5078 (N_5078,N_1889,N_1429);
nand U5079 (N_5079,N_2771,N_594);
nor U5080 (N_5080,N_575,N_389);
nand U5081 (N_5081,N_376,N_1730);
and U5082 (N_5082,N_2988,N_2118);
nand U5083 (N_5083,N_808,N_1327);
nor U5084 (N_5084,N_2087,N_2824);
and U5085 (N_5085,N_2964,N_1308);
or U5086 (N_5086,N_2204,N_844);
or U5087 (N_5087,N_634,N_1426);
or U5088 (N_5088,N_1448,N_2876);
nor U5089 (N_5089,N_844,N_1456);
nor U5090 (N_5090,N_1781,N_1789);
nand U5091 (N_5091,N_1726,N_677);
or U5092 (N_5092,N_1995,N_254);
nor U5093 (N_5093,N_487,N_2609);
nor U5094 (N_5094,N_853,N_2158);
or U5095 (N_5095,N_1252,N_1214);
and U5096 (N_5096,N_606,N_1767);
or U5097 (N_5097,N_337,N_2454);
and U5098 (N_5098,N_2793,N_1911);
nor U5099 (N_5099,N_1056,N_2747);
or U5100 (N_5100,N_115,N_1144);
nand U5101 (N_5101,N_874,N_2728);
nor U5102 (N_5102,N_2059,N_2366);
or U5103 (N_5103,N_2894,N_2819);
nand U5104 (N_5104,N_1253,N_246);
and U5105 (N_5105,N_1617,N_2);
and U5106 (N_5106,N_451,N_2440);
or U5107 (N_5107,N_2191,N_2908);
nor U5108 (N_5108,N_2925,N_1815);
nand U5109 (N_5109,N_1072,N_1476);
and U5110 (N_5110,N_2805,N_1882);
nand U5111 (N_5111,N_1248,N_1241);
and U5112 (N_5112,N_1106,N_2012);
nor U5113 (N_5113,N_1256,N_551);
nor U5114 (N_5114,N_2611,N_419);
nand U5115 (N_5115,N_2162,N_1770);
nand U5116 (N_5116,N_1142,N_770);
nor U5117 (N_5117,N_1902,N_2820);
or U5118 (N_5118,N_2042,N_2213);
nand U5119 (N_5119,N_453,N_227);
and U5120 (N_5120,N_774,N_1949);
and U5121 (N_5121,N_1317,N_991);
nand U5122 (N_5122,N_2322,N_227);
or U5123 (N_5123,N_1232,N_2128);
and U5124 (N_5124,N_1016,N_1836);
and U5125 (N_5125,N_62,N_2559);
nor U5126 (N_5126,N_2225,N_2616);
or U5127 (N_5127,N_585,N_1670);
nor U5128 (N_5128,N_1040,N_712);
or U5129 (N_5129,N_214,N_1450);
nand U5130 (N_5130,N_518,N_99);
nor U5131 (N_5131,N_1142,N_1194);
and U5132 (N_5132,N_1402,N_2872);
nor U5133 (N_5133,N_1424,N_1421);
nor U5134 (N_5134,N_2535,N_2102);
and U5135 (N_5135,N_2478,N_1214);
nand U5136 (N_5136,N_1195,N_1385);
and U5137 (N_5137,N_2171,N_2608);
nand U5138 (N_5138,N_1616,N_2618);
and U5139 (N_5139,N_276,N_71);
and U5140 (N_5140,N_349,N_1431);
and U5141 (N_5141,N_556,N_2735);
nor U5142 (N_5142,N_1910,N_157);
nand U5143 (N_5143,N_1007,N_1346);
or U5144 (N_5144,N_1589,N_480);
and U5145 (N_5145,N_452,N_691);
nor U5146 (N_5146,N_903,N_2404);
or U5147 (N_5147,N_1819,N_1345);
and U5148 (N_5148,N_1104,N_1752);
or U5149 (N_5149,N_1060,N_2443);
or U5150 (N_5150,N_1025,N_2051);
nand U5151 (N_5151,N_411,N_1671);
nand U5152 (N_5152,N_2637,N_2766);
and U5153 (N_5153,N_1066,N_2912);
nand U5154 (N_5154,N_2868,N_223);
nor U5155 (N_5155,N_322,N_2791);
nor U5156 (N_5156,N_2212,N_1986);
nor U5157 (N_5157,N_642,N_2877);
nand U5158 (N_5158,N_120,N_101);
nor U5159 (N_5159,N_2197,N_1827);
or U5160 (N_5160,N_2798,N_2151);
nand U5161 (N_5161,N_684,N_1587);
nor U5162 (N_5162,N_2228,N_2652);
nand U5163 (N_5163,N_372,N_118);
nor U5164 (N_5164,N_415,N_2321);
nor U5165 (N_5165,N_1012,N_368);
nor U5166 (N_5166,N_1564,N_2665);
and U5167 (N_5167,N_761,N_1035);
or U5168 (N_5168,N_2752,N_2652);
nor U5169 (N_5169,N_2736,N_2647);
nor U5170 (N_5170,N_1411,N_816);
or U5171 (N_5171,N_1671,N_1607);
and U5172 (N_5172,N_2887,N_708);
or U5173 (N_5173,N_1760,N_705);
nand U5174 (N_5174,N_2845,N_1696);
or U5175 (N_5175,N_1198,N_1529);
and U5176 (N_5176,N_2027,N_953);
nor U5177 (N_5177,N_553,N_2137);
nor U5178 (N_5178,N_697,N_1505);
or U5179 (N_5179,N_2269,N_804);
or U5180 (N_5180,N_2261,N_2034);
nand U5181 (N_5181,N_617,N_1545);
or U5182 (N_5182,N_1076,N_2451);
and U5183 (N_5183,N_943,N_1867);
and U5184 (N_5184,N_2875,N_612);
nand U5185 (N_5185,N_2850,N_726);
nor U5186 (N_5186,N_382,N_2147);
or U5187 (N_5187,N_2178,N_1488);
and U5188 (N_5188,N_898,N_912);
or U5189 (N_5189,N_1777,N_1268);
or U5190 (N_5190,N_568,N_2611);
and U5191 (N_5191,N_2603,N_1222);
or U5192 (N_5192,N_586,N_138);
nand U5193 (N_5193,N_2484,N_1122);
or U5194 (N_5194,N_1105,N_122);
and U5195 (N_5195,N_549,N_2976);
nor U5196 (N_5196,N_2824,N_2272);
nor U5197 (N_5197,N_393,N_2063);
nor U5198 (N_5198,N_1274,N_1996);
and U5199 (N_5199,N_958,N_1850);
nor U5200 (N_5200,N_1240,N_1025);
and U5201 (N_5201,N_1576,N_625);
nand U5202 (N_5202,N_1613,N_2829);
and U5203 (N_5203,N_1649,N_2165);
nor U5204 (N_5204,N_542,N_1307);
nor U5205 (N_5205,N_2907,N_1655);
or U5206 (N_5206,N_1133,N_902);
nand U5207 (N_5207,N_1786,N_252);
and U5208 (N_5208,N_2934,N_67);
and U5209 (N_5209,N_2353,N_809);
nor U5210 (N_5210,N_1544,N_2783);
or U5211 (N_5211,N_2980,N_1921);
nand U5212 (N_5212,N_502,N_2479);
nor U5213 (N_5213,N_732,N_1130);
nor U5214 (N_5214,N_1251,N_2136);
and U5215 (N_5215,N_866,N_1028);
and U5216 (N_5216,N_2968,N_396);
or U5217 (N_5217,N_2540,N_74);
and U5218 (N_5218,N_2446,N_1379);
nand U5219 (N_5219,N_93,N_944);
and U5220 (N_5220,N_2664,N_1539);
or U5221 (N_5221,N_797,N_1875);
nor U5222 (N_5222,N_2178,N_1818);
nand U5223 (N_5223,N_1564,N_1066);
and U5224 (N_5224,N_387,N_841);
and U5225 (N_5225,N_1501,N_1396);
nand U5226 (N_5226,N_59,N_1362);
or U5227 (N_5227,N_2950,N_2714);
and U5228 (N_5228,N_1700,N_144);
xnor U5229 (N_5229,N_2165,N_2702);
nor U5230 (N_5230,N_566,N_2398);
and U5231 (N_5231,N_2989,N_2108);
nand U5232 (N_5232,N_350,N_743);
and U5233 (N_5233,N_1763,N_2263);
nor U5234 (N_5234,N_2882,N_1719);
or U5235 (N_5235,N_1339,N_1072);
nor U5236 (N_5236,N_1436,N_128);
or U5237 (N_5237,N_497,N_1150);
nand U5238 (N_5238,N_736,N_468);
or U5239 (N_5239,N_2434,N_2448);
and U5240 (N_5240,N_522,N_1923);
and U5241 (N_5241,N_1428,N_113);
and U5242 (N_5242,N_845,N_2356);
or U5243 (N_5243,N_1991,N_841);
nor U5244 (N_5244,N_2525,N_346);
and U5245 (N_5245,N_2353,N_1309);
nand U5246 (N_5246,N_390,N_110);
nand U5247 (N_5247,N_164,N_1781);
nand U5248 (N_5248,N_1339,N_1349);
or U5249 (N_5249,N_1760,N_1571);
nor U5250 (N_5250,N_184,N_2848);
or U5251 (N_5251,N_1008,N_1575);
nand U5252 (N_5252,N_670,N_653);
and U5253 (N_5253,N_1644,N_945);
nand U5254 (N_5254,N_1883,N_1369);
or U5255 (N_5255,N_1112,N_2747);
nor U5256 (N_5256,N_34,N_742);
and U5257 (N_5257,N_1377,N_2113);
or U5258 (N_5258,N_1352,N_2954);
and U5259 (N_5259,N_1397,N_754);
or U5260 (N_5260,N_1808,N_2876);
or U5261 (N_5261,N_2305,N_1302);
nand U5262 (N_5262,N_2454,N_1256);
nor U5263 (N_5263,N_489,N_2872);
or U5264 (N_5264,N_18,N_792);
and U5265 (N_5265,N_1486,N_2025);
and U5266 (N_5266,N_1744,N_2293);
or U5267 (N_5267,N_21,N_2557);
and U5268 (N_5268,N_331,N_320);
or U5269 (N_5269,N_2464,N_333);
nor U5270 (N_5270,N_2059,N_2152);
or U5271 (N_5271,N_2330,N_1274);
nor U5272 (N_5272,N_1108,N_2524);
and U5273 (N_5273,N_433,N_2236);
nand U5274 (N_5274,N_1667,N_2014);
and U5275 (N_5275,N_784,N_2290);
nand U5276 (N_5276,N_2835,N_2611);
and U5277 (N_5277,N_383,N_1923);
nand U5278 (N_5278,N_520,N_1086);
or U5279 (N_5279,N_1545,N_2670);
nor U5280 (N_5280,N_211,N_1870);
nand U5281 (N_5281,N_404,N_2700);
or U5282 (N_5282,N_61,N_192);
and U5283 (N_5283,N_1952,N_344);
or U5284 (N_5284,N_1979,N_750);
and U5285 (N_5285,N_698,N_2277);
or U5286 (N_5286,N_1399,N_1842);
nand U5287 (N_5287,N_1139,N_563);
or U5288 (N_5288,N_238,N_1908);
nor U5289 (N_5289,N_371,N_2295);
and U5290 (N_5290,N_1754,N_558);
nand U5291 (N_5291,N_873,N_376);
nand U5292 (N_5292,N_700,N_1676);
and U5293 (N_5293,N_1684,N_1178);
and U5294 (N_5294,N_2577,N_1753);
nor U5295 (N_5295,N_1612,N_1027);
and U5296 (N_5296,N_1943,N_2708);
nor U5297 (N_5297,N_367,N_2566);
nand U5298 (N_5298,N_736,N_2796);
nor U5299 (N_5299,N_2824,N_30);
nor U5300 (N_5300,N_379,N_1126);
nor U5301 (N_5301,N_591,N_2008);
nand U5302 (N_5302,N_1774,N_1679);
or U5303 (N_5303,N_1603,N_1755);
nor U5304 (N_5304,N_465,N_2456);
and U5305 (N_5305,N_2337,N_1640);
nor U5306 (N_5306,N_1338,N_1390);
nor U5307 (N_5307,N_1644,N_2862);
nand U5308 (N_5308,N_1953,N_1860);
nand U5309 (N_5309,N_2826,N_1480);
or U5310 (N_5310,N_2218,N_421);
nand U5311 (N_5311,N_67,N_2145);
nand U5312 (N_5312,N_301,N_2098);
nor U5313 (N_5313,N_1023,N_1094);
and U5314 (N_5314,N_2798,N_1318);
and U5315 (N_5315,N_131,N_854);
nand U5316 (N_5316,N_844,N_1128);
or U5317 (N_5317,N_19,N_220);
and U5318 (N_5318,N_2391,N_1898);
or U5319 (N_5319,N_126,N_603);
and U5320 (N_5320,N_2720,N_140);
and U5321 (N_5321,N_2793,N_1914);
nor U5322 (N_5322,N_641,N_358);
and U5323 (N_5323,N_549,N_1317);
or U5324 (N_5324,N_2736,N_442);
nor U5325 (N_5325,N_1128,N_2244);
nand U5326 (N_5326,N_806,N_1636);
nor U5327 (N_5327,N_2236,N_2459);
nor U5328 (N_5328,N_821,N_1835);
nand U5329 (N_5329,N_296,N_2860);
and U5330 (N_5330,N_451,N_422);
nand U5331 (N_5331,N_1213,N_320);
nand U5332 (N_5332,N_67,N_2910);
nor U5333 (N_5333,N_2006,N_1418);
nand U5334 (N_5334,N_2133,N_2632);
and U5335 (N_5335,N_1559,N_983);
or U5336 (N_5336,N_2788,N_571);
nand U5337 (N_5337,N_1720,N_1310);
nor U5338 (N_5338,N_2745,N_2732);
nand U5339 (N_5339,N_2851,N_1822);
nor U5340 (N_5340,N_1882,N_2732);
nand U5341 (N_5341,N_548,N_1617);
nor U5342 (N_5342,N_1740,N_2860);
nor U5343 (N_5343,N_2081,N_843);
nand U5344 (N_5344,N_540,N_2149);
nor U5345 (N_5345,N_1993,N_1119);
and U5346 (N_5346,N_1136,N_1830);
nand U5347 (N_5347,N_9,N_2436);
and U5348 (N_5348,N_2972,N_2150);
and U5349 (N_5349,N_2112,N_2804);
nor U5350 (N_5350,N_387,N_103);
or U5351 (N_5351,N_1720,N_1035);
and U5352 (N_5352,N_480,N_2427);
and U5353 (N_5353,N_2770,N_1293);
nand U5354 (N_5354,N_2567,N_1487);
nand U5355 (N_5355,N_2092,N_2917);
or U5356 (N_5356,N_2490,N_336);
nand U5357 (N_5357,N_2915,N_1247);
nand U5358 (N_5358,N_21,N_1642);
or U5359 (N_5359,N_1789,N_2509);
and U5360 (N_5360,N_140,N_2031);
or U5361 (N_5361,N_448,N_1974);
nor U5362 (N_5362,N_1255,N_2576);
nand U5363 (N_5363,N_1339,N_41);
nor U5364 (N_5364,N_2847,N_326);
nor U5365 (N_5365,N_1428,N_2988);
nor U5366 (N_5366,N_2522,N_1829);
nor U5367 (N_5367,N_1170,N_2552);
nand U5368 (N_5368,N_2097,N_2475);
or U5369 (N_5369,N_2170,N_726);
nor U5370 (N_5370,N_828,N_1964);
nand U5371 (N_5371,N_1797,N_2935);
and U5372 (N_5372,N_1158,N_1858);
nand U5373 (N_5373,N_2181,N_1052);
nand U5374 (N_5374,N_2944,N_1844);
or U5375 (N_5375,N_546,N_2842);
nor U5376 (N_5376,N_915,N_318);
nor U5377 (N_5377,N_1612,N_731);
nand U5378 (N_5378,N_1888,N_762);
nor U5379 (N_5379,N_2323,N_2871);
nand U5380 (N_5380,N_968,N_126);
or U5381 (N_5381,N_2228,N_957);
or U5382 (N_5382,N_2193,N_918);
or U5383 (N_5383,N_2139,N_489);
or U5384 (N_5384,N_1401,N_1472);
nand U5385 (N_5385,N_2192,N_2551);
or U5386 (N_5386,N_424,N_1042);
nor U5387 (N_5387,N_2560,N_1936);
and U5388 (N_5388,N_2329,N_2273);
nor U5389 (N_5389,N_2280,N_1938);
nand U5390 (N_5390,N_2989,N_2205);
or U5391 (N_5391,N_1084,N_655);
and U5392 (N_5392,N_1756,N_1503);
and U5393 (N_5393,N_8,N_324);
or U5394 (N_5394,N_1657,N_2852);
nand U5395 (N_5395,N_317,N_243);
nand U5396 (N_5396,N_933,N_1048);
nor U5397 (N_5397,N_118,N_2128);
and U5398 (N_5398,N_292,N_1537);
and U5399 (N_5399,N_1570,N_1649);
nand U5400 (N_5400,N_498,N_429);
and U5401 (N_5401,N_1284,N_2005);
or U5402 (N_5402,N_2883,N_2063);
nand U5403 (N_5403,N_2060,N_1678);
nand U5404 (N_5404,N_1250,N_368);
nand U5405 (N_5405,N_2674,N_1359);
and U5406 (N_5406,N_550,N_1015);
or U5407 (N_5407,N_1295,N_1394);
and U5408 (N_5408,N_874,N_2311);
nand U5409 (N_5409,N_960,N_2219);
and U5410 (N_5410,N_2713,N_917);
or U5411 (N_5411,N_2918,N_172);
nor U5412 (N_5412,N_413,N_1135);
nand U5413 (N_5413,N_1355,N_2662);
nand U5414 (N_5414,N_2654,N_304);
or U5415 (N_5415,N_1304,N_132);
nor U5416 (N_5416,N_1999,N_2562);
nand U5417 (N_5417,N_831,N_2214);
and U5418 (N_5418,N_19,N_1313);
nand U5419 (N_5419,N_2240,N_1171);
and U5420 (N_5420,N_220,N_2683);
or U5421 (N_5421,N_196,N_717);
and U5422 (N_5422,N_639,N_2299);
or U5423 (N_5423,N_1175,N_2378);
nor U5424 (N_5424,N_2721,N_2229);
or U5425 (N_5425,N_628,N_1073);
nand U5426 (N_5426,N_2109,N_231);
nor U5427 (N_5427,N_1706,N_1128);
nand U5428 (N_5428,N_844,N_1529);
or U5429 (N_5429,N_1897,N_2858);
nand U5430 (N_5430,N_2592,N_2099);
nand U5431 (N_5431,N_1428,N_2656);
and U5432 (N_5432,N_633,N_2931);
and U5433 (N_5433,N_343,N_1619);
nand U5434 (N_5434,N_2397,N_102);
nor U5435 (N_5435,N_1461,N_684);
nand U5436 (N_5436,N_2786,N_2555);
nand U5437 (N_5437,N_789,N_246);
nor U5438 (N_5438,N_2499,N_1029);
or U5439 (N_5439,N_2219,N_1081);
or U5440 (N_5440,N_1668,N_1680);
and U5441 (N_5441,N_734,N_1749);
and U5442 (N_5442,N_47,N_1983);
nor U5443 (N_5443,N_2939,N_483);
nor U5444 (N_5444,N_607,N_1234);
or U5445 (N_5445,N_109,N_2563);
nand U5446 (N_5446,N_347,N_2968);
nor U5447 (N_5447,N_2638,N_359);
nor U5448 (N_5448,N_2380,N_948);
and U5449 (N_5449,N_1987,N_1569);
or U5450 (N_5450,N_1296,N_2206);
nand U5451 (N_5451,N_2322,N_49);
nor U5452 (N_5452,N_1972,N_1429);
nor U5453 (N_5453,N_1761,N_2251);
and U5454 (N_5454,N_408,N_1454);
or U5455 (N_5455,N_1292,N_1722);
or U5456 (N_5456,N_1292,N_1597);
nor U5457 (N_5457,N_2216,N_132);
nor U5458 (N_5458,N_1881,N_2530);
nor U5459 (N_5459,N_1616,N_1929);
nand U5460 (N_5460,N_13,N_2798);
or U5461 (N_5461,N_2254,N_1079);
nand U5462 (N_5462,N_77,N_1065);
nand U5463 (N_5463,N_2218,N_2324);
and U5464 (N_5464,N_705,N_160);
and U5465 (N_5465,N_2598,N_639);
nand U5466 (N_5466,N_2569,N_90);
nand U5467 (N_5467,N_184,N_1474);
and U5468 (N_5468,N_1756,N_1370);
or U5469 (N_5469,N_361,N_594);
or U5470 (N_5470,N_2999,N_2892);
and U5471 (N_5471,N_445,N_209);
nand U5472 (N_5472,N_829,N_864);
and U5473 (N_5473,N_1027,N_742);
or U5474 (N_5474,N_2917,N_684);
nor U5475 (N_5475,N_1999,N_636);
and U5476 (N_5476,N_2415,N_1645);
nand U5477 (N_5477,N_1320,N_1426);
and U5478 (N_5478,N_1728,N_1620);
and U5479 (N_5479,N_2046,N_2061);
nor U5480 (N_5480,N_333,N_939);
nand U5481 (N_5481,N_2709,N_1633);
or U5482 (N_5482,N_2493,N_1912);
or U5483 (N_5483,N_1763,N_862);
and U5484 (N_5484,N_1598,N_1871);
or U5485 (N_5485,N_2705,N_1759);
or U5486 (N_5486,N_2539,N_672);
nor U5487 (N_5487,N_730,N_1988);
and U5488 (N_5488,N_2262,N_532);
or U5489 (N_5489,N_1302,N_2132);
nor U5490 (N_5490,N_1385,N_1429);
nor U5491 (N_5491,N_409,N_1495);
nor U5492 (N_5492,N_1814,N_500);
or U5493 (N_5493,N_1654,N_804);
and U5494 (N_5494,N_2912,N_560);
nand U5495 (N_5495,N_2497,N_2475);
and U5496 (N_5496,N_2725,N_1115);
or U5497 (N_5497,N_1520,N_2063);
nor U5498 (N_5498,N_1094,N_23);
xor U5499 (N_5499,N_835,N_490);
or U5500 (N_5500,N_530,N_794);
or U5501 (N_5501,N_2449,N_167);
nand U5502 (N_5502,N_726,N_2974);
nor U5503 (N_5503,N_1512,N_2445);
nor U5504 (N_5504,N_101,N_653);
nor U5505 (N_5505,N_946,N_151);
and U5506 (N_5506,N_1510,N_795);
or U5507 (N_5507,N_202,N_2624);
or U5508 (N_5508,N_2373,N_1561);
or U5509 (N_5509,N_837,N_786);
nand U5510 (N_5510,N_576,N_792);
nand U5511 (N_5511,N_1893,N_2967);
nor U5512 (N_5512,N_1008,N_965);
or U5513 (N_5513,N_2840,N_1103);
nor U5514 (N_5514,N_1289,N_1530);
nor U5515 (N_5515,N_1628,N_845);
nor U5516 (N_5516,N_1481,N_1027);
nand U5517 (N_5517,N_2616,N_1959);
nand U5518 (N_5518,N_552,N_1580);
and U5519 (N_5519,N_1025,N_1326);
and U5520 (N_5520,N_161,N_1109);
and U5521 (N_5521,N_1521,N_2027);
nor U5522 (N_5522,N_825,N_2807);
or U5523 (N_5523,N_63,N_174);
and U5524 (N_5524,N_1698,N_2012);
and U5525 (N_5525,N_693,N_2084);
and U5526 (N_5526,N_1940,N_2301);
nor U5527 (N_5527,N_365,N_694);
nor U5528 (N_5528,N_1330,N_2988);
nand U5529 (N_5529,N_1779,N_1770);
nand U5530 (N_5530,N_1085,N_104);
or U5531 (N_5531,N_988,N_1142);
nand U5532 (N_5532,N_2916,N_1867);
or U5533 (N_5533,N_2364,N_1270);
or U5534 (N_5534,N_2328,N_1479);
and U5535 (N_5535,N_856,N_148);
nand U5536 (N_5536,N_1381,N_951);
and U5537 (N_5537,N_2598,N_2317);
or U5538 (N_5538,N_514,N_1795);
and U5539 (N_5539,N_353,N_251);
or U5540 (N_5540,N_2656,N_1541);
nand U5541 (N_5541,N_1258,N_2920);
and U5542 (N_5542,N_1043,N_110);
or U5543 (N_5543,N_2932,N_1816);
or U5544 (N_5544,N_68,N_1534);
nand U5545 (N_5545,N_82,N_2948);
nand U5546 (N_5546,N_2844,N_876);
nand U5547 (N_5547,N_2069,N_1123);
or U5548 (N_5548,N_2520,N_2756);
nand U5549 (N_5549,N_438,N_210);
nor U5550 (N_5550,N_52,N_502);
nor U5551 (N_5551,N_1783,N_496);
nand U5552 (N_5552,N_1924,N_1590);
and U5553 (N_5553,N_1083,N_836);
or U5554 (N_5554,N_2194,N_2243);
nor U5555 (N_5555,N_293,N_2189);
and U5556 (N_5556,N_1352,N_1305);
nor U5557 (N_5557,N_923,N_2185);
nand U5558 (N_5558,N_338,N_2147);
nor U5559 (N_5559,N_380,N_1436);
nor U5560 (N_5560,N_1563,N_393);
or U5561 (N_5561,N_715,N_685);
nand U5562 (N_5562,N_1227,N_170);
nand U5563 (N_5563,N_1421,N_2685);
nor U5564 (N_5564,N_1602,N_2224);
and U5565 (N_5565,N_1571,N_182);
and U5566 (N_5566,N_2277,N_741);
or U5567 (N_5567,N_999,N_1840);
nor U5568 (N_5568,N_209,N_2977);
and U5569 (N_5569,N_2788,N_1246);
nor U5570 (N_5570,N_1040,N_1829);
and U5571 (N_5571,N_1329,N_2790);
or U5572 (N_5572,N_933,N_2976);
and U5573 (N_5573,N_828,N_2498);
nand U5574 (N_5574,N_39,N_2519);
nand U5575 (N_5575,N_2563,N_2248);
nor U5576 (N_5576,N_2516,N_1115);
and U5577 (N_5577,N_1612,N_695);
or U5578 (N_5578,N_1364,N_267);
and U5579 (N_5579,N_213,N_2103);
nand U5580 (N_5580,N_1816,N_2859);
nor U5581 (N_5581,N_480,N_2036);
and U5582 (N_5582,N_2243,N_504);
and U5583 (N_5583,N_1926,N_2862);
and U5584 (N_5584,N_1415,N_60);
or U5585 (N_5585,N_2895,N_111);
nor U5586 (N_5586,N_1799,N_2713);
nand U5587 (N_5587,N_315,N_1659);
nand U5588 (N_5588,N_2123,N_1564);
or U5589 (N_5589,N_1068,N_1170);
or U5590 (N_5590,N_594,N_2630);
nor U5591 (N_5591,N_328,N_301);
nand U5592 (N_5592,N_1087,N_2690);
nand U5593 (N_5593,N_2510,N_1183);
nand U5594 (N_5594,N_322,N_1298);
and U5595 (N_5595,N_2817,N_2952);
and U5596 (N_5596,N_2860,N_1941);
nor U5597 (N_5597,N_799,N_601);
or U5598 (N_5598,N_912,N_2804);
or U5599 (N_5599,N_1167,N_2217);
nand U5600 (N_5600,N_1999,N_1548);
and U5601 (N_5601,N_348,N_2608);
or U5602 (N_5602,N_564,N_738);
and U5603 (N_5603,N_1798,N_1814);
or U5604 (N_5604,N_987,N_2508);
or U5605 (N_5605,N_2474,N_404);
nor U5606 (N_5606,N_2589,N_2065);
nand U5607 (N_5607,N_2644,N_358);
and U5608 (N_5608,N_36,N_403);
nand U5609 (N_5609,N_2846,N_2680);
nor U5610 (N_5610,N_1151,N_3);
nor U5611 (N_5611,N_576,N_896);
and U5612 (N_5612,N_1193,N_1548);
or U5613 (N_5613,N_1235,N_123);
or U5614 (N_5614,N_1574,N_900);
and U5615 (N_5615,N_305,N_1985);
nand U5616 (N_5616,N_1412,N_723);
and U5617 (N_5617,N_1105,N_2035);
or U5618 (N_5618,N_329,N_1941);
nand U5619 (N_5619,N_2744,N_2941);
and U5620 (N_5620,N_1631,N_1044);
and U5621 (N_5621,N_1625,N_2967);
or U5622 (N_5622,N_1499,N_1862);
and U5623 (N_5623,N_2692,N_1370);
nand U5624 (N_5624,N_2318,N_657);
nor U5625 (N_5625,N_1411,N_1878);
and U5626 (N_5626,N_238,N_1146);
nand U5627 (N_5627,N_1985,N_413);
and U5628 (N_5628,N_1246,N_2701);
and U5629 (N_5629,N_1210,N_138);
or U5630 (N_5630,N_718,N_45);
nand U5631 (N_5631,N_1851,N_1414);
nand U5632 (N_5632,N_1278,N_864);
and U5633 (N_5633,N_1469,N_1597);
nand U5634 (N_5634,N_874,N_2221);
nor U5635 (N_5635,N_2242,N_1188);
or U5636 (N_5636,N_1941,N_255);
nand U5637 (N_5637,N_2601,N_1514);
and U5638 (N_5638,N_1993,N_1255);
or U5639 (N_5639,N_411,N_1283);
nand U5640 (N_5640,N_703,N_1901);
or U5641 (N_5641,N_2377,N_1072);
and U5642 (N_5642,N_993,N_1021);
nor U5643 (N_5643,N_1789,N_1559);
nor U5644 (N_5644,N_653,N_1011);
nand U5645 (N_5645,N_154,N_2092);
or U5646 (N_5646,N_2384,N_2627);
nor U5647 (N_5647,N_2873,N_1679);
or U5648 (N_5648,N_479,N_1503);
nor U5649 (N_5649,N_1987,N_53);
and U5650 (N_5650,N_1391,N_901);
or U5651 (N_5651,N_1210,N_736);
or U5652 (N_5652,N_334,N_2404);
or U5653 (N_5653,N_2175,N_2728);
nor U5654 (N_5654,N_460,N_2210);
nand U5655 (N_5655,N_1723,N_1641);
or U5656 (N_5656,N_2749,N_1949);
and U5657 (N_5657,N_1370,N_2211);
and U5658 (N_5658,N_1665,N_130);
nor U5659 (N_5659,N_1629,N_1736);
nand U5660 (N_5660,N_1802,N_1435);
or U5661 (N_5661,N_348,N_2733);
and U5662 (N_5662,N_635,N_2435);
nor U5663 (N_5663,N_1745,N_1695);
or U5664 (N_5664,N_1373,N_909);
nand U5665 (N_5665,N_490,N_723);
nand U5666 (N_5666,N_2744,N_2800);
or U5667 (N_5667,N_2163,N_805);
nand U5668 (N_5668,N_1735,N_1697);
and U5669 (N_5669,N_1159,N_2348);
nor U5670 (N_5670,N_913,N_799);
nor U5671 (N_5671,N_200,N_2785);
nand U5672 (N_5672,N_2122,N_898);
nor U5673 (N_5673,N_2036,N_501);
nand U5674 (N_5674,N_2143,N_2456);
and U5675 (N_5675,N_1119,N_990);
or U5676 (N_5676,N_88,N_78);
nand U5677 (N_5677,N_1114,N_2597);
or U5678 (N_5678,N_527,N_1857);
nand U5679 (N_5679,N_2446,N_945);
nor U5680 (N_5680,N_1716,N_2686);
nand U5681 (N_5681,N_577,N_803);
and U5682 (N_5682,N_2909,N_782);
nand U5683 (N_5683,N_501,N_1485);
or U5684 (N_5684,N_2179,N_667);
nand U5685 (N_5685,N_2917,N_2340);
or U5686 (N_5686,N_1189,N_2031);
or U5687 (N_5687,N_1632,N_1408);
nor U5688 (N_5688,N_2742,N_662);
and U5689 (N_5689,N_432,N_1643);
nand U5690 (N_5690,N_783,N_813);
nand U5691 (N_5691,N_272,N_2177);
nand U5692 (N_5692,N_2265,N_1823);
nand U5693 (N_5693,N_2265,N_1485);
nand U5694 (N_5694,N_1727,N_2679);
nand U5695 (N_5695,N_644,N_2014);
or U5696 (N_5696,N_1484,N_477);
or U5697 (N_5697,N_371,N_2590);
and U5698 (N_5698,N_594,N_1370);
nor U5699 (N_5699,N_1343,N_2468);
nor U5700 (N_5700,N_1848,N_1286);
nand U5701 (N_5701,N_2151,N_54);
or U5702 (N_5702,N_1416,N_819);
nand U5703 (N_5703,N_710,N_1006);
or U5704 (N_5704,N_1184,N_1763);
or U5705 (N_5705,N_1296,N_146);
nor U5706 (N_5706,N_1234,N_1243);
and U5707 (N_5707,N_2540,N_2930);
and U5708 (N_5708,N_1042,N_1958);
and U5709 (N_5709,N_1884,N_1556);
nand U5710 (N_5710,N_259,N_2892);
and U5711 (N_5711,N_2925,N_145);
and U5712 (N_5712,N_1759,N_2410);
nand U5713 (N_5713,N_1552,N_1529);
nand U5714 (N_5714,N_1041,N_1431);
or U5715 (N_5715,N_1207,N_1538);
and U5716 (N_5716,N_1033,N_570);
and U5717 (N_5717,N_2402,N_1290);
or U5718 (N_5718,N_1636,N_1933);
nor U5719 (N_5719,N_2111,N_1540);
xnor U5720 (N_5720,N_1096,N_168);
nand U5721 (N_5721,N_2469,N_1116);
nand U5722 (N_5722,N_2747,N_1773);
nor U5723 (N_5723,N_96,N_656);
or U5724 (N_5724,N_2979,N_2932);
and U5725 (N_5725,N_2629,N_1535);
and U5726 (N_5726,N_81,N_458);
nand U5727 (N_5727,N_589,N_403);
or U5728 (N_5728,N_376,N_2464);
nor U5729 (N_5729,N_694,N_83);
nor U5730 (N_5730,N_2449,N_602);
or U5731 (N_5731,N_1302,N_2388);
nand U5732 (N_5732,N_2680,N_852);
nand U5733 (N_5733,N_406,N_354);
and U5734 (N_5734,N_2162,N_1284);
or U5735 (N_5735,N_1207,N_192);
nand U5736 (N_5736,N_1503,N_1930);
and U5737 (N_5737,N_596,N_254);
or U5738 (N_5738,N_2746,N_1220);
or U5739 (N_5739,N_470,N_1701);
nor U5740 (N_5740,N_1493,N_234);
nor U5741 (N_5741,N_1864,N_210);
and U5742 (N_5742,N_1200,N_1574);
and U5743 (N_5743,N_1397,N_1959);
and U5744 (N_5744,N_213,N_223);
nor U5745 (N_5745,N_2595,N_497);
nor U5746 (N_5746,N_2118,N_1132);
or U5747 (N_5747,N_2896,N_99);
nand U5748 (N_5748,N_1233,N_2859);
nand U5749 (N_5749,N_2437,N_115);
or U5750 (N_5750,N_776,N_1382);
or U5751 (N_5751,N_2561,N_1201);
nor U5752 (N_5752,N_2768,N_1452);
or U5753 (N_5753,N_320,N_1602);
and U5754 (N_5754,N_2202,N_2610);
nand U5755 (N_5755,N_2169,N_1601);
or U5756 (N_5756,N_2268,N_2139);
and U5757 (N_5757,N_1680,N_1324);
and U5758 (N_5758,N_398,N_1365);
nor U5759 (N_5759,N_177,N_182);
nor U5760 (N_5760,N_1370,N_2220);
nor U5761 (N_5761,N_1678,N_820);
and U5762 (N_5762,N_197,N_866);
or U5763 (N_5763,N_374,N_2454);
and U5764 (N_5764,N_1230,N_1088);
or U5765 (N_5765,N_1287,N_2246);
nand U5766 (N_5766,N_1453,N_417);
and U5767 (N_5767,N_318,N_1835);
or U5768 (N_5768,N_473,N_2249);
nand U5769 (N_5769,N_1089,N_2546);
and U5770 (N_5770,N_2867,N_2041);
and U5771 (N_5771,N_851,N_2587);
nand U5772 (N_5772,N_2853,N_1862);
or U5773 (N_5773,N_2878,N_553);
nor U5774 (N_5774,N_811,N_2517);
or U5775 (N_5775,N_1245,N_2143);
and U5776 (N_5776,N_1840,N_1646);
nand U5777 (N_5777,N_2216,N_702);
and U5778 (N_5778,N_2362,N_2215);
or U5779 (N_5779,N_2134,N_1175);
nand U5780 (N_5780,N_1211,N_1263);
nand U5781 (N_5781,N_1727,N_1856);
nand U5782 (N_5782,N_2602,N_354);
xnor U5783 (N_5783,N_114,N_1577);
or U5784 (N_5784,N_1121,N_2371);
nor U5785 (N_5785,N_874,N_1047);
and U5786 (N_5786,N_526,N_2856);
nor U5787 (N_5787,N_2376,N_2117);
nand U5788 (N_5788,N_1235,N_2811);
or U5789 (N_5789,N_2082,N_59);
nor U5790 (N_5790,N_804,N_2736);
nor U5791 (N_5791,N_2600,N_2438);
nor U5792 (N_5792,N_397,N_2050);
nor U5793 (N_5793,N_2605,N_1580);
nand U5794 (N_5794,N_1177,N_868);
nor U5795 (N_5795,N_268,N_2096);
or U5796 (N_5796,N_2515,N_541);
or U5797 (N_5797,N_2964,N_2609);
nor U5798 (N_5798,N_2500,N_1435);
nor U5799 (N_5799,N_1477,N_1199);
and U5800 (N_5800,N_2702,N_1899);
nand U5801 (N_5801,N_2569,N_1352);
nor U5802 (N_5802,N_690,N_446);
and U5803 (N_5803,N_2065,N_2533);
nor U5804 (N_5804,N_1584,N_1869);
and U5805 (N_5805,N_2292,N_626);
nand U5806 (N_5806,N_2245,N_2041);
or U5807 (N_5807,N_2877,N_377);
or U5808 (N_5808,N_1705,N_328);
or U5809 (N_5809,N_658,N_1456);
nor U5810 (N_5810,N_1828,N_34);
or U5811 (N_5811,N_2577,N_547);
or U5812 (N_5812,N_635,N_1677);
nor U5813 (N_5813,N_2001,N_1261);
nor U5814 (N_5814,N_2727,N_1148);
nand U5815 (N_5815,N_1224,N_2471);
and U5816 (N_5816,N_2036,N_2020);
nor U5817 (N_5817,N_2866,N_1956);
or U5818 (N_5818,N_23,N_2214);
or U5819 (N_5819,N_2184,N_2053);
nor U5820 (N_5820,N_680,N_546);
and U5821 (N_5821,N_2709,N_1139);
or U5822 (N_5822,N_1328,N_1539);
nor U5823 (N_5823,N_216,N_2929);
nand U5824 (N_5824,N_2559,N_1460);
or U5825 (N_5825,N_1710,N_239);
or U5826 (N_5826,N_537,N_372);
or U5827 (N_5827,N_2060,N_2214);
nor U5828 (N_5828,N_1648,N_1008);
nand U5829 (N_5829,N_2443,N_1657);
or U5830 (N_5830,N_727,N_892);
nor U5831 (N_5831,N_1770,N_1250);
and U5832 (N_5832,N_1763,N_1533);
nand U5833 (N_5833,N_96,N_454);
or U5834 (N_5834,N_64,N_2766);
or U5835 (N_5835,N_2608,N_1330);
and U5836 (N_5836,N_1066,N_1108);
nand U5837 (N_5837,N_1565,N_2864);
or U5838 (N_5838,N_157,N_2847);
or U5839 (N_5839,N_1158,N_438);
nor U5840 (N_5840,N_1588,N_622);
or U5841 (N_5841,N_863,N_849);
nand U5842 (N_5842,N_1158,N_1173);
nor U5843 (N_5843,N_2466,N_765);
nor U5844 (N_5844,N_1149,N_1204);
nor U5845 (N_5845,N_1143,N_585);
nand U5846 (N_5846,N_2274,N_558);
and U5847 (N_5847,N_2028,N_2433);
and U5848 (N_5848,N_1549,N_132);
or U5849 (N_5849,N_1635,N_1908);
and U5850 (N_5850,N_2421,N_1583);
and U5851 (N_5851,N_703,N_2155);
and U5852 (N_5852,N_1647,N_1891);
xnor U5853 (N_5853,N_1213,N_1737);
nor U5854 (N_5854,N_863,N_325);
and U5855 (N_5855,N_2084,N_232);
and U5856 (N_5856,N_2628,N_1697);
nand U5857 (N_5857,N_2862,N_1861);
and U5858 (N_5858,N_2299,N_1069);
and U5859 (N_5859,N_2857,N_301);
nand U5860 (N_5860,N_296,N_2784);
nand U5861 (N_5861,N_2547,N_741);
or U5862 (N_5862,N_1162,N_2672);
or U5863 (N_5863,N_689,N_1907);
and U5864 (N_5864,N_2599,N_2326);
nor U5865 (N_5865,N_1366,N_766);
nand U5866 (N_5866,N_657,N_2532);
nand U5867 (N_5867,N_2214,N_2172);
nor U5868 (N_5868,N_2948,N_2608);
nor U5869 (N_5869,N_2676,N_1562);
and U5870 (N_5870,N_496,N_1405);
or U5871 (N_5871,N_2020,N_770);
and U5872 (N_5872,N_160,N_2948);
nand U5873 (N_5873,N_2590,N_1613);
and U5874 (N_5874,N_63,N_2631);
and U5875 (N_5875,N_925,N_1748);
and U5876 (N_5876,N_620,N_2264);
or U5877 (N_5877,N_1366,N_1547);
xnor U5878 (N_5878,N_2154,N_19);
nand U5879 (N_5879,N_1529,N_1112);
nand U5880 (N_5880,N_2896,N_446);
and U5881 (N_5881,N_2265,N_1471);
or U5882 (N_5882,N_194,N_968);
and U5883 (N_5883,N_1523,N_2713);
and U5884 (N_5884,N_2293,N_771);
nor U5885 (N_5885,N_1223,N_161);
and U5886 (N_5886,N_1560,N_112);
nor U5887 (N_5887,N_911,N_1666);
nand U5888 (N_5888,N_492,N_773);
or U5889 (N_5889,N_2156,N_1136);
and U5890 (N_5890,N_1115,N_2870);
nand U5891 (N_5891,N_2511,N_494);
nor U5892 (N_5892,N_1485,N_739);
or U5893 (N_5893,N_414,N_978);
xor U5894 (N_5894,N_2436,N_301);
nand U5895 (N_5895,N_659,N_1168);
and U5896 (N_5896,N_1679,N_1966);
nand U5897 (N_5897,N_2765,N_793);
and U5898 (N_5898,N_1929,N_347);
nand U5899 (N_5899,N_1590,N_1468);
nand U5900 (N_5900,N_547,N_231);
nand U5901 (N_5901,N_2414,N_297);
and U5902 (N_5902,N_2875,N_704);
and U5903 (N_5903,N_2161,N_1675);
nor U5904 (N_5904,N_2836,N_1212);
nand U5905 (N_5905,N_1567,N_1337);
nand U5906 (N_5906,N_1643,N_1651);
or U5907 (N_5907,N_1557,N_2173);
nand U5908 (N_5908,N_1696,N_2732);
nand U5909 (N_5909,N_526,N_550);
or U5910 (N_5910,N_783,N_675);
and U5911 (N_5911,N_2355,N_2174);
or U5912 (N_5912,N_1078,N_1933);
nand U5913 (N_5913,N_2702,N_1588);
and U5914 (N_5914,N_1372,N_116);
nor U5915 (N_5915,N_643,N_873);
or U5916 (N_5916,N_1671,N_440);
nor U5917 (N_5917,N_407,N_2355);
nor U5918 (N_5918,N_2799,N_23);
nor U5919 (N_5919,N_1098,N_84);
or U5920 (N_5920,N_1213,N_673);
or U5921 (N_5921,N_1663,N_103);
nand U5922 (N_5922,N_188,N_1303);
nand U5923 (N_5923,N_2251,N_7);
nor U5924 (N_5924,N_1239,N_1746);
and U5925 (N_5925,N_132,N_313);
or U5926 (N_5926,N_2773,N_1589);
or U5927 (N_5927,N_2423,N_266);
and U5928 (N_5928,N_124,N_2970);
and U5929 (N_5929,N_2540,N_2247);
or U5930 (N_5930,N_1830,N_2996);
or U5931 (N_5931,N_2537,N_1354);
nor U5932 (N_5932,N_1870,N_2360);
nand U5933 (N_5933,N_2243,N_2745);
nand U5934 (N_5934,N_1953,N_1568);
or U5935 (N_5935,N_1746,N_2831);
nor U5936 (N_5936,N_1112,N_824);
and U5937 (N_5937,N_1208,N_574);
or U5938 (N_5938,N_978,N_2122);
nand U5939 (N_5939,N_2678,N_702);
nor U5940 (N_5940,N_2133,N_96);
nor U5941 (N_5941,N_564,N_1267);
and U5942 (N_5942,N_910,N_36);
and U5943 (N_5943,N_2165,N_653);
nand U5944 (N_5944,N_1714,N_1313);
nor U5945 (N_5945,N_528,N_1285);
and U5946 (N_5946,N_2884,N_2999);
nor U5947 (N_5947,N_1150,N_658);
or U5948 (N_5948,N_2762,N_416);
nor U5949 (N_5949,N_1733,N_2046);
or U5950 (N_5950,N_1297,N_1254);
nand U5951 (N_5951,N_1055,N_795);
nand U5952 (N_5952,N_1086,N_2889);
nand U5953 (N_5953,N_1449,N_1498);
or U5954 (N_5954,N_2034,N_2912);
nand U5955 (N_5955,N_2979,N_1461);
or U5956 (N_5956,N_2965,N_2014);
nand U5957 (N_5957,N_33,N_1870);
nand U5958 (N_5958,N_2651,N_789);
nor U5959 (N_5959,N_2687,N_795);
and U5960 (N_5960,N_277,N_1545);
and U5961 (N_5961,N_2811,N_1587);
nand U5962 (N_5962,N_2753,N_2107);
nor U5963 (N_5963,N_1166,N_1338);
nand U5964 (N_5964,N_1072,N_1643);
nand U5965 (N_5965,N_746,N_747);
or U5966 (N_5966,N_764,N_2932);
and U5967 (N_5967,N_2417,N_2626);
nand U5968 (N_5968,N_2810,N_2926);
or U5969 (N_5969,N_1842,N_339);
nor U5970 (N_5970,N_2700,N_517);
nor U5971 (N_5971,N_26,N_2327);
nand U5972 (N_5972,N_1046,N_481);
nor U5973 (N_5973,N_1135,N_2881);
and U5974 (N_5974,N_2698,N_1895);
or U5975 (N_5975,N_1624,N_966);
and U5976 (N_5976,N_1808,N_1574);
and U5977 (N_5977,N_2586,N_365);
nand U5978 (N_5978,N_1772,N_1158);
nand U5979 (N_5979,N_638,N_314);
and U5980 (N_5980,N_1610,N_1906);
or U5981 (N_5981,N_2030,N_2568);
nand U5982 (N_5982,N_703,N_205);
xor U5983 (N_5983,N_753,N_2745);
nor U5984 (N_5984,N_51,N_2497);
nor U5985 (N_5985,N_1226,N_1879);
or U5986 (N_5986,N_1173,N_1394);
and U5987 (N_5987,N_2921,N_10);
nand U5988 (N_5988,N_200,N_1343);
nor U5989 (N_5989,N_1299,N_1947);
nand U5990 (N_5990,N_2044,N_151);
and U5991 (N_5991,N_2812,N_2488);
nor U5992 (N_5992,N_2917,N_1856);
nand U5993 (N_5993,N_220,N_775);
xnor U5994 (N_5994,N_1131,N_2277);
or U5995 (N_5995,N_1913,N_28);
nand U5996 (N_5996,N_426,N_2082);
nand U5997 (N_5997,N_1095,N_2733);
and U5998 (N_5998,N_2695,N_981);
and U5999 (N_5999,N_860,N_522);
and U6000 (N_6000,N_3883,N_3654);
nor U6001 (N_6001,N_4237,N_3142);
or U6002 (N_6002,N_3065,N_5284);
nor U6003 (N_6003,N_3084,N_4418);
and U6004 (N_6004,N_3411,N_3891);
or U6005 (N_6005,N_5117,N_5872);
nand U6006 (N_6006,N_5314,N_3154);
and U6007 (N_6007,N_4700,N_4582);
nand U6008 (N_6008,N_3005,N_4484);
and U6009 (N_6009,N_5964,N_3683);
or U6010 (N_6010,N_4530,N_5026);
nand U6011 (N_6011,N_5688,N_5048);
nor U6012 (N_6012,N_3342,N_5833);
or U6013 (N_6013,N_4870,N_5669);
nor U6014 (N_6014,N_4283,N_3579);
nand U6015 (N_6015,N_5311,N_5654);
and U6016 (N_6016,N_3543,N_3536);
nand U6017 (N_6017,N_3261,N_3068);
nand U6018 (N_6018,N_4580,N_3196);
and U6019 (N_6019,N_3432,N_3774);
nand U6020 (N_6020,N_5751,N_3600);
or U6021 (N_6021,N_4810,N_3834);
xnor U6022 (N_6022,N_4533,N_5179);
and U6023 (N_6023,N_5736,N_4126);
and U6024 (N_6024,N_4316,N_5958);
and U6025 (N_6025,N_3726,N_3361);
or U6026 (N_6026,N_4058,N_3793);
or U6027 (N_6027,N_4224,N_5880);
nor U6028 (N_6028,N_5070,N_3472);
nor U6029 (N_6029,N_5816,N_5538);
nand U6030 (N_6030,N_5148,N_3340);
and U6031 (N_6031,N_5711,N_3431);
nand U6032 (N_6032,N_5400,N_5924);
and U6033 (N_6033,N_3466,N_3540);
nor U6034 (N_6034,N_5259,N_4414);
xnor U6035 (N_6035,N_4786,N_3019);
or U6036 (N_6036,N_3441,N_4758);
nor U6037 (N_6037,N_5365,N_3017);
and U6038 (N_6038,N_3000,N_5805);
nand U6039 (N_6039,N_5670,N_3969);
and U6040 (N_6040,N_4123,N_4965);
and U6041 (N_6041,N_5520,N_4937);
and U6042 (N_6042,N_3296,N_3684);
nand U6043 (N_6043,N_3563,N_5663);
nand U6044 (N_6044,N_4741,N_3162);
or U6045 (N_6045,N_5577,N_3483);
or U6046 (N_6046,N_5991,N_3460);
nand U6047 (N_6047,N_4183,N_4384);
nor U6048 (N_6048,N_3146,N_3632);
or U6049 (N_6049,N_5970,N_3604);
and U6050 (N_6050,N_3062,N_3486);
and U6051 (N_6051,N_5168,N_5348);
nor U6052 (N_6052,N_4903,N_5275);
nand U6053 (N_6053,N_5639,N_4361);
or U6054 (N_6054,N_3149,N_5856);
nand U6055 (N_6055,N_4492,N_5910);
nand U6056 (N_6056,N_4607,N_3766);
or U6057 (N_6057,N_4488,N_3822);
nor U6058 (N_6058,N_3456,N_3729);
and U6059 (N_6059,N_4685,N_3759);
or U6060 (N_6060,N_5007,N_4464);
and U6061 (N_6061,N_4841,N_3039);
nand U6062 (N_6062,N_4665,N_5749);
nand U6063 (N_6063,N_4048,N_5290);
or U6064 (N_6064,N_5362,N_5052);
nand U6065 (N_6065,N_4650,N_5427);
nand U6066 (N_6066,N_3918,N_3509);
or U6067 (N_6067,N_3275,N_4771);
or U6068 (N_6068,N_3699,N_4711);
or U6069 (N_6069,N_5730,N_4033);
nand U6070 (N_6070,N_3445,N_4856);
nand U6071 (N_6071,N_3026,N_4004);
nor U6072 (N_6072,N_4625,N_3475);
or U6073 (N_6073,N_4694,N_5793);
nor U6074 (N_6074,N_4606,N_5810);
nor U6075 (N_6075,N_4621,N_5900);
nand U6076 (N_6076,N_3878,N_4821);
nor U6077 (N_6077,N_4996,N_4335);
nand U6078 (N_6078,N_5491,N_4516);
nor U6079 (N_6079,N_4527,N_4457);
or U6080 (N_6080,N_5912,N_5943);
nand U6081 (N_6081,N_4267,N_3191);
nand U6082 (N_6082,N_3359,N_3896);
nor U6083 (N_6083,N_4654,N_5077);
nand U6084 (N_6084,N_5460,N_3870);
nand U6085 (N_6085,N_5761,N_5861);
or U6086 (N_6086,N_4997,N_4770);
or U6087 (N_6087,N_5118,N_4391);
and U6088 (N_6088,N_3095,N_5263);
or U6089 (N_6089,N_4556,N_3866);
and U6090 (N_6090,N_3665,N_5222);
nor U6091 (N_6091,N_5030,N_4578);
nand U6092 (N_6092,N_3393,N_3193);
or U6093 (N_6093,N_4523,N_5581);
xor U6094 (N_6094,N_4757,N_4295);
and U6095 (N_6095,N_4695,N_3354);
nand U6096 (N_6096,N_4348,N_4249);
or U6097 (N_6097,N_3897,N_4163);
and U6098 (N_6098,N_5554,N_3481);
nand U6099 (N_6099,N_5873,N_5074);
nand U6100 (N_6100,N_4636,N_5518);
and U6101 (N_6101,N_5496,N_4815);
and U6102 (N_6102,N_4838,N_4806);
nand U6103 (N_6103,N_4259,N_5997);
and U6104 (N_6104,N_3016,N_3150);
nor U6105 (N_6105,N_3349,N_5420);
nand U6106 (N_6106,N_4828,N_3298);
and U6107 (N_6107,N_5376,N_4489);
nor U6108 (N_6108,N_3782,N_4644);
or U6109 (N_6109,N_3381,N_5180);
nand U6110 (N_6110,N_3880,N_5944);
and U6111 (N_6111,N_5762,N_5599);
nor U6112 (N_6112,N_3879,N_4215);
and U6113 (N_6113,N_4710,N_4065);
and U6114 (N_6114,N_3144,N_4307);
and U6115 (N_6115,N_5422,N_3024);
and U6116 (N_6116,N_3974,N_3538);
and U6117 (N_6117,N_3605,N_4754);
nor U6118 (N_6118,N_3619,N_3471);
nor U6119 (N_6119,N_3407,N_4571);
or U6120 (N_6120,N_5398,N_4431);
or U6121 (N_6121,N_5937,N_4778);
nor U6122 (N_6122,N_4893,N_4794);
nor U6123 (N_6123,N_3187,N_5595);
nor U6124 (N_6124,N_5836,N_3272);
nand U6125 (N_6125,N_5646,N_3496);
or U6126 (N_6126,N_4887,N_5745);
or U6127 (N_6127,N_3979,N_4861);
or U6128 (N_6128,N_3165,N_5299);
or U6129 (N_6129,N_5563,N_4538);
nor U6130 (N_6130,N_3069,N_3728);
or U6131 (N_6131,N_3940,N_3614);
and U6132 (N_6132,N_4834,N_3723);
and U6133 (N_6133,N_5265,N_5760);
and U6134 (N_6134,N_5384,N_3670);
or U6135 (N_6135,N_3461,N_5813);
and U6136 (N_6136,N_5653,N_4882);
and U6137 (N_6137,N_5390,N_5616);
or U6138 (N_6138,N_5930,N_4385);
nor U6139 (N_6139,N_3963,N_3470);
nor U6140 (N_6140,N_5707,N_3109);
nor U6141 (N_6141,N_5378,N_5102);
or U6142 (N_6142,N_5177,N_3194);
xor U6143 (N_6143,N_5618,N_3955);
and U6144 (N_6144,N_4969,N_5915);
or U6145 (N_6145,N_5773,N_4467);
nor U6146 (N_6146,N_5236,N_4984);
and U6147 (N_6147,N_4880,N_4321);
nor U6148 (N_6148,N_4800,N_4749);
nor U6149 (N_6149,N_3508,N_4010);
and U6150 (N_6150,N_5975,N_5715);
nand U6151 (N_6151,N_3377,N_4509);
and U6152 (N_6152,N_3841,N_4963);
and U6153 (N_6153,N_5134,N_5374);
and U6154 (N_6154,N_4172,N_4862);
or U6155 (N_6155,N_3568,N_3111);
nand U6156 (N_6156,N_3678,N_4114);
or U6157 (N_6157,N_3716,N_3228);
nand U6158 (N_6158,N_4050,N_4765);
nand U6159 (N_6159,N_3888,N_3099);
and U6160 (N_6160,N_5338,N_5559);
and U6161 (N_6161,N_5774,N_4645);
nand U6162 (N_6162,N_3417,N_3707);
xnor U6163 (N_6163,N_4083,N_4909);
or U6164 (N_6164,N_4474,N_3698);
and U6165 (N_6165,N_5936,N_4293);
nor U6166 (N_6166,N_4734,N_3308);
nand U6167 (N_6167,N_4956,N_5887);
xnor U6168 (N_6168,N_3830,N_3003);
nand U6169 (N_6169,N_4426,N_5812);
or U6170 (N_6170,N_5747,N_3779);
nand U6171 (N_6171,N_4317,N_4136);
or U6172 (N_6172,N_5181,N_3552);
and U6173 (N_6173,N_5549,N_4929);
nor U6174 (N_6174,N_4857,N_4790);
nor U6175 (N_6175,N_3603,N_5297);
nand U6176 (N_6176,N_3862,N_4454);
or U6177 (N_6177,N_3905,N_4148);
nand U6178 (N_6178,N_3128,N_3567);
or U6179 (N_6179,N_5381,N_3971);
or U6180 (N_6180,N_5307,N_4078);
nand U6181 (N_6181,N_3249,N_3976);
or U6182 (N_6182,N_4389,N_5735);
nor U6183 (N_6183,N_4367,N_5136);
nand U6184 (N_6184,N_4167,N_4242);
or U6185 (N_6185,N_4742,N_5217);
nand U6186 (N_6186,N_4994,N_3337);
or U6187 (N_6187,N_5171,N_5324);
nor U6188 (N_6188,N_4539,N_3041);
and U6189 (N_6189,N_5462,N_4207);
nor U6190 (N_6190,N_5596,N_5661);
nor U6191 (N_6191,N_4737,N_3574);
nand U6192 (N_6192,N_3922,N_5459);
nand U6193 (N_6193,N_4152,N_4975);
and U6194 (N_6194,N_4440,N_3435);
nor U6195 (N_6195,N_5725,N_4192);
or U6196 (N_6196,N_4410,N_3789);
nor U6197 (N_6197,N_4420,N_3480);
and U6198 (N_6198,N_3843,N_5005);
nor U6199 (N_6199,N_5902,N_5218);
nand U6200 (N_6200,N_3220,N_5876);
and U6201 (N_6201,N_3242,N_4001);
or U6202 (N_6202,N_5124,N_4382);
nor U6203 (N_6203,N_4716,N_5457);
or U6204 (N_6204,N_4416,N_3184);
or U6205 (N_6205,N_3693,N_3070);
nor U6206 (N_6206,N_5527,N_5788);
or U6207 (N_6207,N_4564,N_5742);
or U6208 (N_6208,N_5929,N_5351);
or U6209 (N_6209,N_4455,N_4421);
nor U6210 (N_6210,N_4976,N_4917);
nand U6211 (N_6211,N_3833,N_5656);
nor U6212 (N_6212,N_4992,N_4659);
and U6213 (N_6213,N_5045,N_3842);
nor U6214 (N_6214,N_4236,N_3776);
nand U6215 (N_6215,N_3105,N_3190);
nand U6216 (N_6216,N_3088,N_3073);
nor U6217 (N_6217,N_5585,N_4681);
or U6218 (N_6218,N_5449,N_3036);
nand U6219 (N_6219,N_5027,N_4206);
nor U6220 (N_6220,N_3791,N_5032);
and U6221 (N_6221,N_5504,N_4752);
nor U6222 (N_6222,N_4042,N_4583);
or U6223 (N_6223,N_5184,N_5023);
and U6224 (N_6224,N_4931,N_4101);
and U6225 (N_6225,N_4477,N_5474);
nand U6226 (N_6226,N_4279,N_3704);
or U6227 (N_6227,N_4499,N_3264);
and U6228 (N_6228,N_5607,N_3973);
and U6229 (N_6229,N_5232,N_4386);
nor U6230 (N_6230,N_4679,N_5359);
and U6231 (N_6231,N_5128,N_3028);
xor U6232 (N_6232,N_3763,N_5723);
and U6233 (N_6233,N_5660,N_3288);
nor U6234 (N_6234,N_5874,N_5617);
nor U6235 (N_6235,N_5847,N_4543);
or U6236 (N_6236,N_5285,N_3322);
and U6237 (N_6237,N_5965,N_5739);
or U6238 (N_6238,N_4405,N_4823);
or U6239 (N_6239,N_4519,N_3437);
nand U6240 (N_6240,N_5315,N_4592);
nand U6241 (N_6241,N_3853,N_4220);
and U6242 (N_6242,N_4291,N_4993);
and U6243 (N_6243,N_5316,N_3629);
nand U6244 (N_6244,N_4461,N_3916);
and U6245 (N_6245,N_5811,N_4194);
and U6246 (N_6246,N_5093,N_5666);
and U6247 (N_6247,N_3688,N_5692);
or U6248 (N_6248,N_4038,N_4831);
nand U6249 (N_6249,N_4748,N_5984);
and U6250 (N_6250,N_4978,N_3239);
or U6251 (N_6251,N_3899,N_4891);
or U6252 (N_6252,N_5853,N_5208);
nand U6253 (N_6253,N_5310,N_4755);
and U6254 (N_6254,N_3383,N_3825);
and U6255 (N_6255,N_5994,N_5642);
and U6256 (N_6256,N_5101,N_4653);
or U6257 (N_6257,N_3283,N_4877);
nor U6258 (N_6258,N_3176,N_4198);
nand U6259 (N_6259,N_5100,N_4812);
and U6260 (N_6260,N_5200,N_3804);
or U6261 (N_6261,N_4103,N_4676);
nand U6262 (N_6262,N_5972,N_3932);
nor U6263 (N_6263,N_4719,N_3977);
and U6264 (N_6264,N_3387,N_4195);
or U6265 (N_6265,N_3355,N_3424);
or U6266 (N_6266,N_3625,N_5779);
and U6267 (N_6267,N_5354,N_4472);
or U6268 (N_6268,N_3281,N_5683);
and U6269 (N_6269,N_3198,N_4682);
nor U6270 (N_6270,N_5106,N_3867);
and U6271 (N_6271,N_5202,N_5963);
and U6272 (N_6272,N_4018,N_3443);
nor U6273 (N_6273,N_4008,N_3755);
or U6274 (N_6274,N_5056,N_5605);
nand U6275 (N_6275,N_4087,N_3076);
and U6276 (N_6276,N_3679,N_4166);
or U6277 (N_6277,N_4353,N_4478);
nand U6278 (N_6278,N_3170,N_4753);
or U6279 (N_6279,N_4113,N_4529);
nand U6280 (N_6280,N_5176,N_5840);
nand U6281 (N_6281,N_4261,N_5521);
and U6282 (N_6282,N_5417,N_3506);
nor U6283 (N_6283,N_4013,N_4190);
or U6284 (N_6284,N_3330,N_4160);
nor U6285 (N_6285,N_4034,N_5602);
nor U6286 (N_6286,N_3257,N_5305);
or U6287 (N_6287,N_5884,N_4112);
nand U6288 (N_6288,N_3391,N_3369);
and U6289 (N_6289,N_4573,N_5434);
nand U6290 (N_6290,N_5904,N_5705);
nand U6291 (N_6291,N_4450,N_3725);
or U6292 (N_6292,N_4155,N_4130);
and U6293 (N_6293,N_3663,N_3948);
nor U6294 (N_6294,N_5183,N_3912);
nand U6295 (N_6295,N_4832,N_5241);
or U6296 (N_6296,N_5868,N_5926);
or U6297 (N_6297,N_3999,N_5744);
nor U6298 (N_6298,N_3018,N_5204);
or U6299 (N_6299,N_4026,N_4272);
or U6300 (N_6300,N_5437,N_3380);
and U6301 (N_6301,N_3612,N_4497);
and U6302 (N_6302,N_4874,N_3490);
nand U6303 (N_6303,N_4505,N_4173);
and U6304 (N_6304,N_3245,N_3061);
nand U6305 (N_6305,N_4407,N_4429);
or U6306 (N_6306,N_5151,N_3054);
and U6307 (N_6307,N_5877,N_4177);
and U6308 (N_6308,N_5016,N_4156);
nor U6309 (N_6309,N_4235,N_4002);
and U6310 (N_6310,N_5546,N_3771);
nand U6311 (N_6311,N_5039,N_4954);
nor U6312 (N_6312,N_4175,N_4513);
nor U6313 (N_6313,N_5110,N_4133);
or U6314 (N_6314,N_3010,N_5846);
nor U6315 (N_6315,N_4853,N_4808);
and U6316 (N_6316,N_5619,N_3837);
and U6317 (N_6317,N_5716,N_4157);
nand U6318 (N_6318,N_5835,N_4390);
nor U6319 (N_6319,N_4756,N_4759);
or U6320 (N_6320,N_4071,N_3601);
or U6321 (N_6321,N_5541,N_4364);
nor U6322 (N_6322,N_5543,N_3967);
or U6323 (N_6323,N_3401,N_4964);
or U6324 (N_6324,N_3285,N_5610);
and U6325 (N_6325,N_5388,N_4159);
nand U6326 (N_6326,N_4022,N_4935);
nor U6327 (N_6327,N_5426,N_5651);
nand U6328 (N_6328,N_4671,N_4436);
or U6329 (N_6329,N_4922,N_4121);
and U6330 (N_6330,N_4397,N_5848);
nor U6331 (N_6331,N_3092,N_3739);
and U6332 (N_6332,N_3856,N_4433);
nor U6333 (N_6333,N_4995,N_5075);
and U6334 (N_6334,N_3012,N_3320);
nor U6335 (N_6335,N_5364,N_4186);
nand U6336 (N_6336,N_4016,N_5476);
and U6337 (N_6337,N_5678,N_4518);
and U6338 (N_6338,N_5797,N_4037);
nand U6339 (N_6339,N_4745,N_3127);
or U6340 (N_6340,N_4072,N_5503);
nand U6341 (N_6341,N_3964,N_3682);
nor U6342 (N_6342,N_5821,N_5588);
and U6343 (N_6343,N_4814,N_4938);
and U6344 (N_6344,N_3637,N_4313);
nor U6345 (N_6345,N_3748,N_3937);
nor U6346 (N_6346,N_4339,N_5274);
nand U6347 (N_6347,N_3179,N_5405);
and U6348 (N_6348,N_4168,N_5411);
or U6349 (N_6349,N_3892,N_4602);
nand U6350 (N_6350,N_4275,N_5624);
and U6351 (N_6351,N_4865,N_4662);
nor U6352 (N_6352,N_3367,N_3658);
nor U6353 (N_6353,N_5078,N_3675);
nor U6354 (N_6354,N_4377,N_5062);
nand U6355 (N_6355,N_4596,N_3474);
and U6356 (N_6356,N_3849,N_4804);
and U6357 (N_6357,N_5073,N_4998);
nand U6358 (N_6358,N_3415,N_5485);
and U6359 (N_6359,N_4598,N_4846);
or U6360 (N_6360,N_5794,N_4171);
or U6361 (N_6361,N_3767,N_5589);
or U6362 (N_6362,N_4302,N_5239);
nor U6363 (N_6363,N_3305,N_3643);
nand U6364 (N_6364,N_3284,N_4793);
nand U6365 (N_6365,N_3449,N_3809);
nor U6366 (N_6366,N_3364,N_3929);
or U6367 (N_6367,N_3520,N_3124);
nor U6368 (N_6368,N_3114,N_5412);
and U6369 (N_6369,N_3208,N_4552);
and U6370 (N_6370,N_5352,N_4306);
nand U6371 (N_6371,N_3232,N_3042);
nand U6372 (N_6372,N_5010,N_3983);
and U6373 (N_6373,N_5054,N_3130);
or U6374 (N_6374,N_3265,N_4061);
nor U6375 (N_6375,N_5780,N_4712);
nor U6376 (N_6376,N_4380,N_5233);
or U6377 (N_6377,N_3181,N_5011);
and U6378 (N_6378,N_5008,N_5450);
or U6379 (N_6379,N_5814,N_4240);
nand U6380 (N_6380,N_5867,N_5681);
nor U6381 (N_6381,N_5252,N_3622);
and U6382 (N_6382,N_3920,N_3332);
nor U6383 (N_6383,N_4945,N_5837);
nand U6384 (N_6384,N_3233,N_5419);
or U6385 (N_6385,N_5373,N_4280);
or U6386 (N_6386,N_5012,N_3510);
or U6387 (N_6387,N_4471,N_5031);
nor U6388 (N_6388,N_5555,N_3389);
nand U6389 (N_6389,N_3489,N_3172);
and U6390 (N_6390,N_3395,N_3950);
or U6391 (N_6391,N_3269,N_3203);
nor U6392 (N_6392,N_4179,N_4501);
nand U6393 (N_6393,N_3423,N_3901);
or U6394 (N_6394,N_4692,N_5757);
and U6395 (N_6395,N_4221,N_4941);
nand U6396 (N_6396,N_3593,N_3624);
nand U6397 (N_6397,N_3416,N_5264);
or U6398 (N_6398,N_5341,N_4350);
nand U6399 (N_6399,N_3497,N_4506);
nor U6400 (N_6400,N_5216,N_3338);
nand U6401 (N_6401,N_3734,N_3855);
or U6402 (N_6402,N_4647,N_4281);
and U6403 (N_6403,N_4773,N_3266);
or U6404 (N_6404,N_4904,N_4266);
or U6405 (N_6405,N_3202,N_4735);
nand U6406 (N_6406,N_3015,N_5603);
or U6407 (N_6407,N_3936,N_4025);
nor U6408 (N_6408,N_5754,N_4507);
nand U6409 (N_6409,N_5925,N_5143);
nor U6410 (N_6410,N_4864,N_3446);
or U6411 (N_6411,N_4491,N_3914);
nand U6412 (N_6412,N_3067,N_3171);
xnor U6413 (N_6413,N_5500,N_3764);
or U6414 (N_6414,N_4442,N_3794);
and U6415 (N_6415,N_3664,N_3487);
or U6416 (N_6416,N_5598,N_4041);
nor U6417 (N_6417,N_4381,N_3096);
nand U6418 (N_6418,N_4219,N_4906);
nand U6419 (N_6419,N_3174,N_3812);
nor U6420 (N_6420,N_3908,N_4709);
nand U6421 (N_6421,N_3805,N_5244);
nor U6422 (N_6422,N_3123,N_3797);
nor U6423 (N_6423,N_5892,N_4706);
nand U6424 (N_6424,N_5129,N_3676);
nand U6425 (N_6425,N_3363,N_5535);
or U6426 (N_6426,N_5006,N_3558);
or U6427 (N_6427,N_3956,N_5652);
and U6428 (N_6428,N_4035,N_5146);
nor U6429 (N_6429,N_4835,N_3255);
or U6430 (N_6430,N_3350,N_4928);
and U6431 (N_6431,N_5261,N_3134);
nand U6432 (N_6432,N_4690,N_5750);
or U6433 (N_6433,N_4926,N_3339);
nor U6434 (N_6434,N_4553,N_5104);
or U6435 (N_6435,N_5049,N_4624);
nand U6436 (N_6436,N_5854,N_3256);
and U6437 (N_6437,N_5098,N_3902);
or U6438 (N_6438,N_4446,N_5463);
xnor U6439 (N_6439,N_3136,N_5591);
xnor U6440 (N_6440,N_4840,N_4127);
and U6441 (N_6441,N_3692,N_4696);
nand U6442 (N_6442,N_5211,N_3104);
and U6443 (N_6443,N_5832,N_5905);
or U6444 (N_6444,N_5506,N_3572);
and U6445 (N_6445,N_3781,N_4108);
or U6446 (N_6446,N_5826,N_5022);
nand U6447 (N_6447,N_3260,N_5277);
or U6448 (N_6448,N_5825,N_3225);
nand U6449 (N_6449,N_5631,N_3680);
and U6450 (N_6450,N_4100,N_5532);
or U6451 (N_6451,N_5145,N_3083);
nand U6452 (N_6452,N_3863,N_5628);
and U6453 (N_6453,N_3773,N_5262);
and U6454 (N_6454,N_4122,N_3345);
or U6455 (N_6455,N_4554,N_3204);
and U6456 (N_6456,N_3981,N_5121);
nor U6457 (N_6457,N_3458,N_3169);
and U6458 (N_6458,N_3117,N_5433);
and U6459 (N_6459,N_5766,N_5186);
nand U6460 (N_6460,N_4579,N_4601);
nand U6461 (N_6461,N_4732,N_4591);
or U6462 (N_6462,N_5719,N_5404);
nor U6463 (N_6463,N_3941,N_5014);
and U6464 (N_6464,N_3711,N_4181);
or U6465 (N_6465,N_5295,N_4830);
and U6466 (N_6466,N_4054,N_3116);
nor U6467 (N_6467,N_4576,N_3851);
nor U6468 (N_6468,N_5511,N_5584);
nor U6469 (N_6469,N_3021,N_5334);
nor U6470 (N_6470,N_5668,N_5763);
nor U6471 (N_6471,N_5704,N_3493);
nor U6472 (N_6472,N_3697,N_4532);
or U6473 (N_6473,N_3120,N_4337);
nor U6474 (N_6474,N_5103,N_5732);
nand U6475 (N_6475,N_5718,N_4760);
nand U6476 (N_6476,N_3378,N_5621);
and U6477 (N_6477,N_4663,N_4845);
xor U6478 (N_6478,N_3178,N_4691);
nand U6479 (N_6479,N_3221,N_4044);
and U6480 (N_6480,N_4199,N_5492);
nor U6481 (N_6481,N_3397,N_5115);
nor U6482 (N_6482,N_5210,N_4608);
or U6483 (N_6483,N_4586,N_4310);
and U6484 (N_6484,N_3410,N_3262);
and U6485 (N_6485,N_5391,N_4727);
or U6486 (N_6486,N_5120,N_3998);
nor U6487 (N_6487,N_4762,N_3960);
nand U6488 (N_6488,N_3156,N_3945);
or U6489 (N_6489,N_3295,N_5230);
nor U6490 (N_6490,N_3219,N_3746);
nand U6491 (N_6491,N_4620,N_5069);
or U6492 (N_6492,N_3796,N_3695);
and U6493 (N_6493,N_3652,N_4971);
or U6494 (N_6494,N_4419,N_5679);
nand U6495 (N_6495,N_3714,N_5135);
and U6496 (N_6496,N_4378,N_4413);
or U6497 (N_6497,N_5772,N_4357);
or U6498 (N_6498,N_5323,N_3529);
or U6499 (N_6499,N_5094,N_4848);
nor U6500 (N_6500,N_3223,N_3669);
and U6501 (N_6501,N_5547,N_4558);
or U6502 (N_6502,N_3107,N_4656);
and U6503 (N_6503,N_5899,N_5424);
nor U6504 (N_6504,N_4398,N_3640);
nor U6505 (N_6505,N_5156,N_5820);
or U6506 (N_6506,N_3957,N_5565);
nand U6507 (N_6507,N_3653,N_3168);
or U6508 (N_6508,N_4705,N_5389);
and U6509 (N_6509,N_4686,N_4638);
nor U6510 (N_6510,N_5502,N_5795);
or U6511 (N_6511,N_4634,N_5697);
and U6512 (N_6512,N_4017,N_4792);
and U6513 (N_6513,N_4803,N_4504);
and U6514 (N_6514,N_5939,N_3408);
and U6515 (N_6515,N_4612,N_5672);
nor U6516 (N_6516,N_3659,N_3311);
nor U6517 (N_6517,N_5455,N_4162);
nand U6518 (N_6518,N_5920,N_3164);
nand U6519 (N_6519,N_3173,N_5785);
nor U6520 (N_6520,N_4807,N_5173);
nor U6521 (N_6521,N_4693,N_5286);
nand U6522 (N_6522,N_4508,N_3864);
and U6523 (N_6523,N_5472,N_5063);
nand U6524 (N_6524,N_3958,N_5144);
or U6525 (N_6525,N_3785,N_3591);
and U6526 (N_6526,N_4332,N_5933);
nor U6527 (N_6527,N_4435,N_3222);
nor U6528 (N_6528,N_4544,N_5465);
nor U6529 (N_6529,N_3677,N_5556);
nor U6530 (N_6530,N_4069,N_5843);
nor U6531 (N_6531,N_5320,N_5968);
nand U6532 (N_6532,N_3009,N_3523);
nor U6533 (N_6533,N_3869,N_5796);
or U6534 (N_6534,N_4067,N_5999);
and U6535 (N_6535,N_4725,N_5035);
and U6536 (N_6536,N_4842,N_4546);
nor U6537 (N_6537,N_4427,N_3872);
and U6538 (N_6538,N_3821,N_5830);
and U6539 (N_6539,N_3004,N_3690);
and U6540 (N_6540,N_3832,N_5524);
and U6541 (N_6541,N_5258,N_3278);
nand U6542 (N_6542,N_4209,N_5024);
or U6543 (N_6543,N_5907,N_4271);
or U6544 (N_6544,N_3947,N_3768);
nand U6545 (N_6545,N_3720,N_5765);
or U6546 (N_6546,N_5175,N_4081);
or U6547 (N_6547,N_5221,N_3206);
nand U6548 (N_6548,N_4697,N_5065);
nand U6549 (N_6549,N_3718,N_3343);
or U6550 (N_6550,N_3649,N_5980);
nor U6551 (N_6551,N_5629,N_5281);
or U6552 (N_6552,N_4940,N_5695);
nor U6553 (N_6553,N_4358,N_3696);
nor U6554 (N_6554,N_3077,N_3091);
nand U6555 (N_6555,N_4649,N_5300);
nand U6556 (N_6556,N_3362,N_4117);
nand U6557 (N_6557,N_5076,N_4816);
and U6558 (N_6558,N_3592,N_5844);
nand U6559 (N_6559,N_3059,N_5017);
nand U6560 (N_6560,N_3201,N_3399);
nand U6561 (N_6561,N_4324,N_3621);
nor U6562 (N_6562,N_3990,N_5278);
and U6563 (N_6563,N_4459,N_3344);
nor U6564 (N_6564,N_5392,N_5029);
or U6565 (N_6565,N_4363,N_4423);
nand U6566 (N_6566,N_5137,N_3501);
and U6567 (N_6567,N_3861,N_3951);
or U6568 (N_6568,N_5394,N_4943);
nand U6569 (N_6569,N_4104,N_5397);
or U6570 (N_6570,N_4777,N_3750);
or U6571 (N_6571,N_4424,N_3499);
and U6572 (N_6572,N_3770,N_4203);
or U6573 (N_6573,N_5347,N_3259);
and U6574 (N_6574,N_3882,N_4836);
or U6575 (N_6575,N_4919,N_5097);
nand U6576 (N_6576,N_5871,N_4228);
nand U6577 (N_6577,N_4524,N_3813);
nor U6578 (N_6578,N_3422,N_4541);
nor U6579 (N_6579,N_3072,N_4822);
or U6580 (N_6580,N_4388,N_3140);
and U6581 (N_6581,N_3597,N_3302);
or U6582 (N_6582,N_5706,N_4052);
or U6583 (N_6583,N_4406,N_5369);
and U6584 (N_6584,N_3559,N_5053);
xnor U6585 (N_6585,N_3743,N_5896);
nand U6586 (N_6586,N_5237,N_3735);
and U6587 (N_6587,N_4256,N_4570);
or U6588 (N_6588,N_5850,N_5140);
nor U6589 (N_6589,N_5978,N_4340);
nor U6590 (N_6590,N_5229,N_4918);
and U6591 (N_6591,N_4217,N_4566);
nand U6592 (N_6592,N_5256,N_3029);
nor U6593 (N_6593,N_4232,N_4779);
or U6594 (N_6594,N_3752,N_5522);
and U6595 (N_6595,N_5190,N_5615);
xor U6596 (N_6596,N_3442,N_3313);
nand U6597 (N_6597,N_5079,N_5823);
or U6598 (N_6598,N_5552,N_5335);
nor U6599 (N_6599,N_5199,N_3035);
or U6600 (N_6600,N_5990,N_3778);
nor U6601 (N_6601,N_5906,N_5649);
and U6602 (N_6602,N_3240,N_4051);
nor U6603 (N_6603,N_4642,N_5138);
nor U6604 (N_6604,N_5446,N_3189);
nand U6605 (N_6605,N_4927,N_4355);
or U6606 (N_6606,N_3814,N_4496);
nor U6607 (N_6607,N_4577,N_4912);
or U6608 (N_6608,N_3780,N_5717);
nand U6609 (N_6609,N_4952,N_4703);
nand U6610 (N_6610,N_4669,N_5699);
nor U6611 (N_6611,N_4730,N_5676);
nor U6612 (N_6612,N_3795,N_5312);
and U6613 (N_6613,N_5881,N_3907);
and U6614 (N_6614,N_4430,N_5674);
and U6615 (N_6615,N_3180,N_4677);
nand U6616 (N_6616,N_4520,N_3573);
nor U6617 (N_6617,N_4039,N_4374);
nand U6618 (N_6618,N_4110,N_3315);
and U6619 (N_6619,N_5081,N_4955);
nor U6620 (N_6620,N_3623,N_5611);
nand U6621 (N_6621,N_5575,N_5125);
nor U6622 (N_6622,N_5786,N_4327);
nor U6623 (N_6623,N_5822,N_3706);
nor U6624 (N_6624,N_4447,N_3001);
nor U6625 (N_6625,N_3721,N_5021);
and U6626 (N_6626,N_5042,N_5831);
nand U6627 (N_6627,N_4563,N_5336);
nor U6628 (N_6628,N_5122,N_5260);
and U6629 (N_6629,N_5291,N_4991);
nand U6630 (N_6630,N_4129,N_4057);
nor U6631 (N_6631,N_3808,N_3270);
or U6632 (N_6632,N_5321,N_5954);
and U6633 (N_6633,N_4107,N_4356);
or U6634 (N_6634,N_4908,N_4666);
or U6635 (N_6635,N_3943,N_3053);
and U6636 (N_6636,N_3935,N_4818);
or U6637 (N_6637,N_4920,N_3628);
and U6638 (N_6638,N_4032,N_5322);
nand U6639 (N_6639,N_4738,N_3984);
or U6640 (N_6640,N_5741,N_3463);
nor U6641 (N_6641,N_4802,N_5499);
nand U6642 (N_6642,N_4255,N_3419);
and U6643 (N_6643,N_5729,N_5440);
or U6644 (N_6644,N_4432,N_4837);
nand U6645 (N_6645,N_4796,N_3153);
nor U6646 (N_6646,N_5562,N_5174);
and U6647 (N_6647,N_4257,N_5004);
or U6648 (N_6648,N_3263,N_5254);
nand U6649 (N_6649,N_4049,N_4318);
nand U6650 (N_6650,N_3473,N_5977);
or U6651 (N_6651,N_4597,N_4149);
or U6652 (N_6652,N_5396,N_5934);
and U6653 (N_6653,N_4099,N_3336);
and U6654 (N_6654,N_5046,N_4750);
nand U6655 (N_6655,N_3583,N_3384);
nor U6656 (N_6656,N_5386,N_5519);
nor U6657 (N_6657,N_4096,N_4589);
nor U6658 (N_6658,N_3158,N_3754);
and U6659 (N_6659,N_3524,N_3844);
and U6660 (N_6660,N_4053,N_5266);
or U6661 (N_6661,N_4260,N_4066);
or U6662 (N_6662,N_5147,N_4486);
or U6663 (N_6663,N_3300,N_4417);
nor U6664 (N_6664,N_4784,N_4562);
nand U6665 (N_6665,N_5539,N_4886);
nand U6666 (N_6666,N_3148,N_3823);
nor U6667 (N_6667,N_5209,N_3216);
and U6668 (N_6668,N_4683,N_4141);
nand U6669 (N_6669,N_4131,N_3884);
nand U6670 (N_6670,N_3816,N_3900);
or U6671 (N_6671,N_3535,N_5303);
nand U6672 (N_6672,N_4522,N_5526);
nor U6673 (N_6673,N_4811,N_5090);
nor U6674 (N_6674,N_3209,N_5009);
and U6675 (N_6675,N_4603,N_4343);
nand U6676 (N_6676,N_5141,N_5667);
and U6677 (N_6677,N_4143,N_5448);
nand U6678 (N_6678,N_4086,N_5111);
nand U6679 (N_6679,N_4287,N_3968);
or U6680 (N_6680,N_4277,N_3102);
or U6681 (N_6681,N_5640,N_5720);
and U6682 (N_6682,N_3457,N_4820);
nor U6683 (N_6683,N_3824,N_5824);
nor U6684 (N_6684,N_5447,N_3465);
nand U6685 (N_6685,N_3512,N_3243);
nor U6686 (N_6686,N_3581,N_4320);
nor U6687 (N_6687,N_5185,N_5153);
and U6688 (N_6688,N_5438,N_5205);
nor U6689 (N_6689,N_4315,N_4019);
or U6690 (N_6690,N_4074,N_3719);
nand U6691 (N_6691,N_3118,N_5213);
nand U6692 (N_6692,N_5452,N_3093);
or U6693 (N_6693,N_5803,N_3141);
or U6694 (N_6694,N_3939,N_4568);
nand U6695 (N_6695,N_5306,N_4905);
and U6696 (N_6696,N_5623,N_5060);
nor U6697 (N_6697,N_4346,N_4411);
or U6698 (N_6698,N_5377,N_5159);
or U6699 (N_6699,N_4204,N_3758);
and U6700 (N_6700,N_4819,N_3006);
nor U6701 (N_6701,N_3331,N_4763);
and U6702 (N_6702,N_4897,N_4161);
and U6703 (N_6703,N_4899,N_5091);
or U6704 (N_6704,N_5531,N_3712);
nand U6705 (N_6705,N_4479,N_4664);
nand U6706 (N_6706,N_3548,N_3569);
nor U6707 (N_6707,N_5512,N_5142);
nor U6708 (N_6708,N_5249,N_5268);
nand U6709 (N_6709,N_3681,N_5545);
and U6710 (N_6710,N_4788,N_3056);
nor U6711 (N_6711,N_5356,N_3691);
or U6712 (N_6712,N_4670,N_4631);
nand U6713 (N_6713,N_5572,N_4623);
nor U6714 (N_6714,N_4714,N_4284);
or U6715 (N_6715,N_5878,N_4960);
nor U6716 (N_6716,N_5370,N_3551);
or U6717 (N_6717,N_4201,N_4744);
nor U6718 (N_6718,N_5080,N_4785);
and U6719 (N_6719,N_5182,N_5686);
and U6720 (N_6720,N_4463,N_4323);
nor U6721 (N_6721,N_3993,N_3404);
and U6722 (N_6722,N_5866,N_4005);
nand U6723 (N_6723,N_3710,N_5368);
nor U6724 (N_6724,N_4060,N_3358);
nor U6725 (N_6725,N_3644,N_5108);
nor U6726 (N_6726,N_3709,N_3661);
nor U6727 (N_6727,N_4613,N_5234);
nor U6728 (N_6728,N_3820,N_3555);
nand U6729 (N_6729,N_5188,N_3868);
or U6730 (N_6730,N_5408,N_3268);
nand U6731 (N_6731,N_4795,N_5033);
and U6732 (N_6732,N_3020,N_3143);
nor U6733 (N_6733,N_4000,N_4797);
or U6734 (N_6734,N_4341,N_3316);
and U6735 (N_6735,N_5809,N_5643);
and U6736 (N_6736,N_5331,N_4253);
nand U6737 (N_6737,N_5313,N_5085);
and U6738 (N_6738,N_3412,N_4898);
nor U6739 (N_6739,N_4813,N_3327);
nor U6740 (N_6740,N_3052,N_5895);
nor U6741 (N_6741,N_4376,N_4875);
and U6742 (N_6742,N_4957,N_4627);
or U6743 (N_6743,N_5992,N_4707);
nor U6744 (N_6744,N_5693,N_3089);
nand U6745 (N_6745,N_5072,N_4717);
nand U6746 (N_6746,N_3087,N_3112);
nor U6747 (N_6747,N_5326,N_4699);
or U6748 (N_6748,N_4510,N_4652);
and U6749 (N_6749,N_3732,N_5919);
xor U6750 (N_6750,N_4400,N_3230);
nor U6751 (N_6751,N_3532,N_3090);
nand U6752 (N_6752,N_3066,N_3894);
nand U6753 (N_6753,N_3045,N_4138);
nor U6754 (N_6754,N_3970,N_4024);
nand U6755 (N_6755,N_3959,N_3546);
nor U6756 (N_6756,N_3826,N_3986);
nor U6757 (N_6757,N_4154,N_3286);
xor U6758 (N_6758,N_5609,N_3515);
or U6759 (N_6759,N_3613,N_5413);
nand U6760 (N_6760,N_4443,N_4689);
nor U6761 (N_6761,N_3609,N_5731);
or U6762 (N_6762,N_4537,N_5701);
nor U6763 (N_6763,N_5827,N_3598);
or U6764 (N_6764,N_5219,N_5604);
and U6765 (N_6765,N_4614,N_3213);
nor U6766 (N_6766,N_4055,N_5487);
and U6767 (N_6767,N_5036,N_3989);
nand U6768 (N_6768,N_3836,N_3464);
and U6769 (N_6769,N_3876,N_3085);
and U6770 (N_6770,N_4628,N_3440);
or U6771 (N_6771,N_4672,N_5292);
and U6772 (N_6772,N_3803,N_5901);
and U6773 (N_6773,N_3611,N_4292);
nand U6774 (N_6774,N_4924,N_3137);
and U6775 (N_6775,N_4415,N_4263);
nor U6776 (N_6776,N_3040,N_4170);
and U6777 (N_6777,N_5909,N_3385);
nand U6778 (N_6778,N_5423,N_5633);
and U6779 (N_6779,N_4512,N_5586);
nand U6780 (N_6780,N_5296,N_4977);
or U6781 (N_6781,N_3329,N_3386);
and U6782 (N_6782,N_5673,N_4359);
and U6783 (N_6783,N_4393,N_5486);
nor U6784 (N_6784,N_4245,N_3476);
and U6785 (N_6785,N_3166,N_3846);
and U6786 (N_6786,N_5941,N_5540);
and U6787 (N_6787,N_4345,N_4056);
and U6788 (N_6788,N_4946,N_4799);
and U6789 (N_6789,N_3875,N_4789);
nor U6790 (N_6790,N_3537,N_3097);
or U6791 (N_6791,N_3627,N_4914);
nor U6792 (N_6792,N_4999,N_5453);
nand U6793 (N_6793,N_5451,N_4319);
and U6794 (N_6794,N_4982,N_3352);
nand U6795 (N_6795,N_5571,N_5196);
and U6796 (N_6796,N_5911,N_4787);
or U6797 (N_6797,N_4241,N_4495);
or U6798 (N_6798,N_4827,N_3185);
nor U6799 (N_6799,N_5636,N_5635);
or U6800 (N_6800,N_5366,N_4809);
nor U6801 (N_6801,N_4526,N_4604);
and U6802 (N_6802,N_3533,N_3375);
nor U6803 (N_6803,N_5342,N_3525);
nand U6804 (N_6804,N_5066,N_4366);
nand U6805 (N_6805,N_3616,N_4545);
xnor U6806 (N_6806,N_3662,N_3672);
or U6807 (N_6807,N_3046,N_4197);
or U6808 (N_6808,N_5682,N_4718);
nor U6809 (N_6809,N_3992,N_4879);
nor U6810 (N_6810,N_5787,N_4772);
nand U6811 (N_6811,N_3495,N_4401);
xor U6812 (N_6812,N_3588,N_4584);
nor U6813 (N_6813,N_4211,N_3370);
nor U6814 (N_6814,N_4180,N_4125);
nand U6815 (N_6815,N_4106,N_5890);
and U6816 (N_6816,N_4174,N_5626);
and U6817 (N_6817,N_4325,N_3571);
nor U6818 (N_6818,N_5996,N_4333);
or U6819 (N_6819,N_4238,N_3002);
nor U6820 (N_6820,N_3646,N_4517);
and U6821 (N_6821,N_3923,N_5570);
and U6822 (N_6822,N_5439,N_5139);
or U6823 (N_6823,N_4404,N_5922);
and U6824 (N_6824,N_3366,N_5214);
nand U6825 (N_6825,N_5484,N_5510);
nand U6826 (N_6826,N_4063,N_3451);
and U6827 (N_6827,N_4003,N_4187);
nand U6828 (N_6828,N_3252,N_4585);
and U6829 (N_6829,N_4134,N_5436);
nand U6830 (N_6830,N_4047,N_4896);
nand U6831 (N_6831,N_5375,N_3197);
and U6832 (N_6832,N_5340,N_5627);
and U6833 (N_6833,N_3639,N_5696);
or U6834 (N_6834,N_3772,N_5862);
or U6835 (N_6835,N_4801,N_3724);
and U6836 (N_6836,N_4502,N_5332);
xor U6837 (N_6837,N_3547,N_3078);
and U6838 (N_6838,N_3815,N_3008);
or U6839 (N_6839,N_4200,N_4322);
nand U6840 (N_6840,N_5415,N_4470);
or U6841 (N_6841,N_5838,N_3564);
and U6842 (N_6842,N_5864,N_4213);
or U6843 (N_6843,N_5298,N_5276);
nand U6844 (N_6844,N_4970,N_5777);
and U6845 (N_6845,N_3351,N_4723);
or U6846 (N_6846,N_5228,N_5505);
and U6847 (N_6847,N_4839,N_4967);
or U6848 (N_6848,N_3044,N_4036);
nand U6849 (N_6849,N_4581,N_5650);
nor U6850 (N_6850,N_3694,N_4089);
nand U6851 (N_6851,N_5702,N_5157);
or U6852 (N_6852,N_5908,N_5250);
or U6853 (N_6853,N_4768,N_5431);
nor U6854 (N_6854,N_4330,N_3100);
and U6855 (N_6855,N_5223,N_4867);
nor U6856 (N_6856,N_4439,N_4950);
and U6857 (N_6857,N_4702,N_5771);
nor U6858 (N_6858,N_3827,N_3211);
and U6859 (N_6859,N_3517,N_3271);
nor U6860 (N_6860,N_3231,N_4142);
nand U6861 (N_6861,N_4278,N_3713);
or U6862 (N_6862,N_5680,N_4902);
nand U6863 (N_6863,N_3835,N_5995);
nand U6864 (N_6864,N_3214,N_5852);
nand U6865 (N_6865,N_3910,N_3975);
nand U6866 (N_6866,N_3626,N_4782);
nor U6867 (N_6867,N_5123,N_5630);
nor U6868 (N_6868,N_4030,N_5025);
nor U6869 (N_6869,N_4866,N_3615);
xnor U6870 (N_6870,N_3101,N_3025);
nor U6871 (N_6871,N_3182,N_3365);
nor U6872 (N_6872,N_5560,N_3356);
nand U6873 (N_6873,N_3291,N_4305);
nand U6874 (N_6874,N_3094,N_3453);
and U6875 (N_6875,N_3048,N_3110);
nor U6876 (N_6876,N_4402,N_5957);
nor U6877 (N_6877,N_5429,N_3309);
or U6878 (N_6878,N_3060,N_3139);
nor U6879 (N_6879,N_5728,N_5224);
nand U6880 (N_6880,N_3513,N_3133);
and U6881 (N_6881,N_5947,N_3819);
nand U6882 (N_6882,N_4490,N_4265);
or U6883 (N_6883,N_3689,N_3433);
nand U6884 (N_6884,N_4375,N_4487);
or U6885 (N_6885,N_5245,N_3562);
and U6886 (N_6886,N_3398,N_3590);
and U6887 (N_6887,N_5665,N_3234);
nor U6888 (N_6888,N_5951,N_5304);
nand U6889 (N_6889,N_5869,N_3787);
nand U6890 (N_6890,N_3786,N_3687);
nor U6891 (N_6891,N_5383,N_3850);
nand U6892 (N_6892,N_5569,N_3982);
and U6893 (N_6893,N_3810,N_3392);
nand U6894 (N_6894,N_4214,N_4483);
and U6895 (N_6895,N_5067,N_5675);
and U6896 (N_6896,N_4395,N_5191);
and U6897 (N_6897,N_5482,N_4216);
or U6898 (N_6898,N_5644,N_3602);
or U6899 (N_6899,N_3273,N_4873);
or U6900 (N_6900,N_3942,N_3854);
or U6901 (N_6901,N_5817,N_3700);
or U6902 (N_6902,N_4883,N_4328);
and U6903 (N_6903,N_3650,N_5113);
and U6904 (N_6904,N_5410,N_5105);
nor U6905 (N_6905,N_4936,N_5960);
and U6906 (N_6906,N_5480,N_4888);
or U6907 (N_6907,N_5088,N_3403);
nor U6908 (N_6908,N_4588,N_3987);
and U6909 (N_6909,N_5952,N_4088);
or U6910 (N_6910,N_5150,N_5689);
nor U6911 (N_6911,N_3444,N_4210);
nand U6912 (N_6912,N_3917,N_3584);
nand U6913 (N_6913,N_5525,N_5255);
nand U6914 (N_6914,N_4262,N_4043);
or U6915 (N_6915,N_4521,N_3426);
or U6916 (N_6916,N_5165,N_3373);
nor U6917 (N_6917,N_3893,N_5523);
nand U6918 (N_6918,N_4668,N_5126);
and U6919 (N_6919,N_3954,N_4169);
nand U6920 (N_6920,N_5099,N_4274);
nor U6921 (N_6921,N_3642,N_5989);
nand U6922 (N_6922,N_3790,N_3634);
or U6923 (N_6923,N_5553,N_4860);
and U6924 (N_6924,N_3183,N_4942);
nor U6925 (N_6925,N_5253,N_5748);
nand U6926 (N_6926,N_3829,N_3554);
and U6927 (N_6927,N_5859,N_4480);
or U6928 (N_6928,N_4128,N_4503);
nand U6929 (N_6929,N_5658,N_4482);
nor U6930 (N_6930,N_5976,N_4660);
and U6931 (N_6931,N_3930,N_4064);
nand U6932 (N_6932,N_4599,N_3237);
nand U6933 (N_6933,N_5738,N_3668);
nand U6934 (N_6934,N_3762,N_5516);
nand U6935 (N_6935,N_3733,N_3292);
nand U6936 (N_6936,N_5040,N_3160);
nand U6937 (N_6937,N_3933,N_4244);
and U6938 (N_6938,N_3507,N_4090);
nor U6939 (N_6939,N_5573,N_3953);
or U6940 (N_6940,N_5568,N_3439);
nor U6941 (N_6941,N_5170,N_4233);
or U6942 (N_6942,N_4739,N_5068);
or U6943 (N_6943,N_3745,N_4408);
nand U6944 (N_6944,N_4643,N_3115);
nor U6945 (N_6945,N_5898,N_3454);
and U6946 (N_6946,N_4843,N_5597);
or U6947 (N_6947,N_4276,N_5966);
or U6948 (N_6948,N_3301,N_5612);
xor U6949 (N_6949,N_3757,N_3267);
nand U6950 (N_6950,N_4514,N_3570);
nor U6951 (N_6951,N_3889,N_3049);
and U6952 (N_6952,N_4297,N_4347);
nor U6953 (N_6953,N_5592,N_3560);
nor U6954 (N_6954,N_3860,N_5302);
and U6955 (N_6955,N_3526,N_4973);
nor U6956 (N_6956,N_5353,N_3769);
and U6957 (N_6957,N_5087,N_3753);
and U6958 (N_6958,N_4890,N_4139);
or U6959 (N_6959,N_5293,N_4269);
nor U6960 (N_6960,N_5421,N_4246);
nand U6961 (N_6961,N_3648,N_4329);
nand U6962 (N_6962,N_3541,N_4680);
and U6963 (N_6963,N_5647,N_5641);
or U6964 (N_6964,N_5659,N_3371);
and U6965 (N_6965,N_4428,N_3421);
nand U6966 (N_6966,N_4135,N_4569);
and U6967 (N_6967,N_4040,N_4176);
nor U6968 (N_6968,N_3561,N_3656);
and U6969 (N_6969,N_5799,N_4085);
or U6970 (N_6970,N_5393,N_4979);
nor U6971 (N_6971,N_3051,N_3106);
or U6972 (N_6972,N_5567,N_3119);
nor U6973 (N_6973,N_3557,N_3828);
nand U6974 (N_6974,N_5841,N_5301);
or U6975 (N_6975,N_3961,N_5212);
and U6976 (N_6976,N_4646,N_3038);
nor U6977 (N_6977,N_3436,N_4798);
and U6978 (N_6978,N_5530,N_4774);
nor U6979 (N_6979,N_5483,N_4561);
nor U6980 (N_6980,N_5769,N_5557);
nor U6981 (N_6981,N_4567,N_5467);
nor U6982 (N_6982,N_5133,N_3500);
or U6983 (N_6983,N_3666,N_3161);
or U6984 (N_6984,N_5703,N_5435);
nor U6985 (N_6985,N_3516,N_5346);
nand U6986 (N_6986,N_4540,N_4250);
and U6987 (N_6987,N_5201,N_5916);
or U6988 (N_6988,N_3946,N_4445);
and U6989 (N_6989,N_3199,N_4565);
and U6990 (N_6990,N_5095,N_5969);
nor U6991 (N_6991,N_4535,N_3368);
nand U6992 (N_6992,N_3931,N_5000);
nor U6993 (N_6993,N_4120,N_4178);
or U6994 (N_6994,N_3800,N_5402);
nor U6995 (N_6995,N_5444,N_4360);
and U6996 (N_6996,N_4968,N_5829);
or U6997 (N_6997,N_3839,N_4314);
nor U6998 (N_6998,N_5734,N_5536);
nand U6999 (N_6999,N_3919,N_3522);
nor U7000 (N_7000,N_4536,N_4422);
nor U7001 (N_7001,N_4743,N_3505);
and U7002 (N_7002,N_5481,N_4675);
nand U7003 (N_7003,N_5248,N_4202);
nand U7004 (N_7004,N_3258,N_4985);
nand U7005 (N_7005,N_3207,N_5220);
nor U7006 (N_7006,N_3542,N_3921);
and U7007 (N_7007,N_4234,N_5737);
and U7008 (N_7008,N_4222,N_5270);
nor U7009 (N_7009,N_3576,N_5594);
and U7010 (N_7010,N_3904,N_5923);
or U7011 (N_7011,N_4460,N_4549);
nor U7012 (N_7012,N_3756,N_3323);
xor U7013 (N_7013,N_3784,N_5194);
nor U7014 (N_7014,N_4290,N_4948);
nor U7015 (N_7015,N_5756,N_3147);
nand U7016 (N_7016,N_3731,N_5458);
nand U7017 (N_7017,N_3528,N_4892);
or U7018 (N_7018,N_3425,N_4326);
and U7019 (N_7019,N_5395,N_5935);
nor U7020 (N_7020,N_4409,N_5399);
or U7021 (N_7021,N_5514,N_3459);
nand U7022 (N_7022,N_5828,N_3071);
nor U7023 (N_7023,N_5700,N_5579);
and U7024 (N_7024,N_4988,N_4342);
nor U7025 (N_7025,N_5086,N_3577);
nand U7026 (N_7026,N_3818,N_3064);
nand U7027 (N_7027,N_5513,N_5187);
or U7028 (N_7028,N_5363,N_3450);
or U7029 (N_7029,N_5792,N_5019);
and U7030 (N_7030,N_5279,N_4387);
nand U7031 (N_7031,N_3630,N_4437);
nor U7032 (N_7032,N_3037,N_4006);
nand U7033 (N_7033,N_3589,N_4587);
and U7034 (N_7034,N_4633,N_3488);
nand U7035 (N_7035,N_3200,N_4655);
or U7036 (N_7036,N_5608,N_3409);
or U7037 (N_7037,N_5329,N_3788);
and U7038 (N_7038,N_4989,N_4910);
nor U7039 (N_7039,N_3324,N_4102);
or U7040 (N_7040,N_4311,N_3317);
or U7041 (N_7041,N_3840,N_5238);
nand U7042 (N_7042,N_3502,N_4379);
nor U7043 (N_7043,N_5517,N_5807);
or U7044 (N_7044,N_5548,N_5784);
nand U7045 (N_7045,N_3881,N_5698);
nor U7046 (N_7046,N_5294,N_5712);
nor U7047 (N_7047,N_4858,N_3503);
nand U7048 (N_7048,N_3877,N_3925);
and U7049 (N_7049,N_5897,N_5507);
nand U7050 (N_7050,N_3685,N_4595);
nor U7051 (N_7051,N_3596,N_4288);
nand U7052 (N_7052,N_5657,N_5215);
or U7053 (N_7053,N_4452,N_3521);
and U7054 (N_7054,N_3224,N_5037);
nor U7055 (N_7055,N_3701,N_4158);
nor U7056 (N_7056,N_4850,N_5114);
nor U7057 (N_7057,N_4494,N_3218);
nand U7058 (N_7058,N_3175,N_4678);
nand U7059 (N_7059,N_4118,N_3674);
nor U7060 (N_7060,N_5889,N_5724);
nand U7061 (N_7061,N_4029,N_4438);
nand U7062 (N_7062,N_4365,N_4273);
nand U7063 (N_7063,N_3469,N_3924);
or U7064 (N_7064,N_3477,N_5043);
and U7065 (N_7065,N_5606,N_3293);
nor U7066 (N_7066,N_4331,N_4894);
and U7067 (N_7067,N_3565,N_4684);
nor U7068 (N_7068,N_5464,N_5587);
nand U7069 (N_7069,N_4212,N_5013);
and U7070 (N_7070,N_3586,N_5882);
nor U7071 (N_7071,N_3708,N_5020);
nor U7072 (N_7072,N_3227,N_4987);
nand U7073 (N_7073,N_5050,N_5973);
and U7074 (N_7074,N_4466,N_4481);
nor U7075 (N_7075,N_5339,N_5089);
or U7076 (N_7076,N_4731,N_5337);
nor U7077 (N_7077,N_3727,N_3934);
nand U7078 (N_7078,N_3031,N_3742);
xor U7079 (N_7079,N_4825,N_3913);
and U7080 (N_7080,N_3909,N_4352);
and U7081 (N_7081,N_5684,N_4434);
and U7082 (N_7082,N_3396,N_5819);
nand U7083 (N_7083,N_4859,N_3594);
and U7084 (N_7084,N_3125,N_4630);
and U7085 (N_7085,N_3811,N_4304);
nand U7086 (N_7086,N_4884,N_3394);
nand U7087 (N_7087,N_5308,N_3238);
nand U7088 (N_7088,N_3430,N_5961);
or U7089 (N_7089,N_5534,N_3347);
or U7090 (N_7090,N_5379,N_5380);
nand U7091 (N_7091,N_3138,N_3282);
nor U7092 (N_7092,N_4299,N_4781);
or U7093 (N_7093,N_3599,N_3098);
or U7094 (N_7094,N_5454,N_5015);
nor U7095 (N_7095,N_4593,N_4226);
xor U7096 (N_7096,N_3388,N_5677);
nor U7097 (N_7097,N_4961,N_5330);
nand U7098 (N_7098,N_3462,N_4775);
or U7099 (N_7099,N_5109,N_4111);
and U7100 (N_7100,N_4729,N_5319);
or U7101 (N_7101,N_3730,N_4618);
and U7102 (N_7102,N_3413,N_5403);
nand U7103 (N_7103,N_4225,N_3082);
and U7104 (N_7104,N_4252,N_5409);
xnor U7105 (N_7105,N_4708,N_5955);
and U7106 (N_7106,N_3607,N_5967);
nor U7107 (N_7107,N_4344,N_4916);
nand U7108 (N_7108,N_5112,N_4247);
and U7109 (N_7109,N_3608,N_4109);
nor U7110 (N_7110,N_5443,N_3806);
nand U7111 (N_7111,N_3075,N_5888);
nand U7112 (N_7112,N_4915,N_5345);
nand U7113 (N_7113,N_3595,N_5834);
nand U7114 (N_7114,N_4640,N_4070);
nand U7115 (N_7115,N_3050,N_5946);
nor U7116 (N_7116,N_4009,N_5815);
or U7117 (N_7117,N_3585,N_4951);
nor U7118 (N_7118,N_4336,N_5456);
and U7119 (N_7119,N_5893,N_3702);
nand U7120 (N_7120,N_3667,N_3996);
nand U7121 (N_7121,N_5613,N_4747);
nor U7122 (N_7122,N_5921,N_3353);
nor U7123 (N_7123,N_3927,N_5582);
or U7124 (N_7124,N_5529,N_4124);
or U7125 (N_7125,N_4098,N_5280);
nor U7126 (N_7126,N_3129,N_3289);
nand U7127 (N_7127,N_3580,N_5428);
and U7128 (N_7128,N_5055,N_5344);
nor U7129 (N_7129,N_5061,N_3011);
or U7130 (N_7130,N_3376,N_4534);
nand U7131 (N_7131,N_3290,N_3379);
and U7132 (N_7132,N_4286,N_3241);
or U7133 (N_7133,N_4468,N_3578);
and U7134 (N_7134,N_3427,N_4205);
or U7135 (N_7135,N_4981,N_4594);
nor U7136 (N_7136,N_3749,N_5576);
xnor U7137 (N_7137,N_4045,N_5855);
or U7138 (N_7138,N_5493,N_4383);
or U7139 (N_7139,N_3467,N_5361);
or U7140 (N_7140,N_4907,N_5367);
nor U7141 (N_7141,N_4885,N_4673);
or U7142 (N_7142,N_4635,N_3550);
or U7143 (N_7143,N_5551,N_4824);
nand U7144 (N_7144,N_3871,N_4736);
and U7145 (N_7145,N_5564,N_4721);
nor U7146 (N_7146,N_4097,N_4188);
nand U7147 (N_7147,N_4062,N_3145);
xnor U7148 (N_7148,N_5498,N_4462);
nand U7149 (N_7149,N_5993,N_4733);
nand U7150 (N_7150,N_3215,N_3556);
nor U7151 (N_7151,N_4469,N_4441);
or U7152 (N_7152,N_3250,N_4144);
nor U7153 (N_7153,N_5743,N_5883);
or U7154 (N_7154,N_3086,N_5119);
and U7155 (N_7155,N_3997,N_5903);
nand U7156 (N_7156,N_3492,N_4934);
and U7157 (N_7157,N_5164,N_5158);
and U7158 (N_7158,N_3294,N_4394);
nor U7159 (N_7159,N_4849,N_3205);
nand U7160 (N_7160,N_4371,N_3485);
nor U7161 (N_7161,N_4575,N_5034);
nor U7162 (N_7162,N_5385,N_3831);
or U7163 (N_7163,N_3737,N_3188);
and U7164 (N_7164,N_4722,N_5600);
and U7165 (N_7165,N_4791,N_3022);
or U7166 (N_7166,N_5798,N_5489);
or U7167 (N_7167,N_3438,N_5478);
nand U7168 (N_7168,N_4615,N_4498);
and U7169 (N_7169,N_4667,N_4485);
nand U7170 (N_7170,N_3033,N_5632);
nor U7171 (N_7171,N_3798,N_3400);
and U7172 (N_7172,N_3553,N_5722);
nand U7173 (N_7173,N_4657,N_3455);
and U7174 (N_7174,N_5246,N_4303);
nand U7175 (N_7175,N_5953,N_5645);
or U7176 (N_7176,N_5981,N_5289);
or U7177 (N_7177,N_4572,N_4610);
nor U7178 (N_7178,N_3360,N_3135);
nor U7179 (N_7179,N_4740,N_3802);
and U7180 (N_7180,N_4559,N_3848);
or U7181 (N_7181,N_3448,N_4300);
and U7182 (N_7182,N_4476,N_4119);
or U7183 (N_7183,N_5207,N_5988);
nor U7184 (N_7184,N_5614,N_4243);
and U7185 (N_7185,N_5638,N_4590);
and U7186 (N_7186,N_5789,N_4079);
or U7187 (N_7187,N_5566,N_4425);
xor U7188 (N_7188,N_5288,N_3740);
or U7189 (N_7189,N_5387,N_3306);
or U7190 (N_7190,N_5740,N_4132);
nand U7191 (N_7191,N_3043,N_4465);
nand U7192 (N_7192,N_3303,N_3277);
and U7193 (N_7193,N_4115,N_5894);
nor U7194 (N_7194,N_5783,N_3527);
and U7195 (N_7195,N_5733,N_4027);
nor U7196 (N_7196,N_3926,N_5414);
nand U7197 (N_7197,N_3775,N_4091);
and U7198 (N_7198,N_3801,N_4334);
and U7199 (N_7199,N_3890,N_5860);
nand U7200 (N_7200,N_4116,N_4164);
or U7201 (N_7201,N_5318,N_4068);
or U7202 (N_7202,N_5710,N_3346);
nor U7203 (N_7203,N_3995,N_4766);
nor U7204 (N_7204,N_5620,N_3511);
or U7205 (N_7205,N_3985,N_4296);
nor U7206 (N_7206,N_3874,N_5622);
nor U7207 (N_7207,N_3341,N_4073);
or U7208 (N_7208,N_4231,N_4913);
nand U7209 (N_7209,N_5350,N_4312);
nor U7210 (N_7210,N_5441,N_3402);
and U7211 (N_7211,N_3906,N_5469);
nand U7212 (N_7212,N_4751,N_4855);
nand U7213 (N_7213,N_4184,N_5044);
or U7214 (N_7214,N_5770,N_4370);
or U7215 (N_7215,N_5727,N_4641);
and U7216 (N_7216,N_3751,N_3949);
or U7217 (N_7217,N_5802,N_5694);
or U7218 (N_7218,N_5857,N_5461);
nand U7219 (N_7219,N_4869,N_3530);
and U7220 (N_7220,N_3055,N_3229);
nand U7221 (N_7221,N_4551,N_5959);
nand U7222 (N_7222,N_4547,N_5949);
nand U7223 (N_7223,N_5561,N_5851);
nand U7224 (N_7224,N_3783,N_3638);
nand U7225 (N_7225,N_3657,N_3152);
nand U7226 (N_7226,N_3434,N_4605);
nor U7227 (N_7227,N_3063,N_4146);
nand U7228 (N_7228,N_3980,N_5328);
and U7229 (N_7229,N_5092,N_4616);
or U7230 (N_7230,N_4020,N_3747);
and U7231 (N_7231,N_4574,N_3186);
nor U7232 (N_7232,N_4720,N_4309);
nand U7233 (N_7233,N_5986,N_3514);
or U7234 (N_7234,N_5003,N_3299);
nand U7235 (N_7235,N_5528,N_5166);
nand U7236 (N_7236,N_4185,N_4528);
nor U7237 (N_7237,N_3328,N_4193);
nand U7238 (N_7238,N_5508,N_4550);
and U7239 (N_7239,N_5468,N_5637);
nand U7240 (N_7240,N_5082,N_5755);
or U7241 (N_7241,N_3857,N_3057);
or U7242 (N_7242,N_3321,N_5791);
nor U7243 (N_7243,N_5163,N_3254);
or U7244 (N_7244,N_5987,N_4872);
nor U7245 (N_7245,N_3314,N_5515);
and U7246 (N_7246,N_3817,N_4826);
and U7247 (N_7247,N_3647,N_3304);
or U7248 (N_7248,N_4218,N_4674);
or U7249 (N_7249,N_5913,N_4966);
and U7250 (N_7250,N_3617,N_3032);
and U7251 (N_7251,N_3792,N_3155);
or U7252 (N_7252,N_5051,N_5601);
or U7253 (N_7253,N_3518,N_5355);
and U7254 (N_7254,N_4511,N_3122);
xor U7255 (N_7255,N_4458,N_4629);
or U7256 (N_7256,N_4023,N_4456);
or U7257 (N_7257,N_5782,N_5418);
or U7258 (N_7258,N_5768,N_3248);
or U7259 (N_7259,N_4847,N_5808);
nand U7260 (N_7260,N_5084,N_3307);
nand U7261 (N_7261,N_5243,N_4369);
nand U7262 (N_7262,N_4046,N_3807);
nand U7263 (N_7263,N_4769,N_3962);
and U7264 (N_7264,N_3027,N_4844);
nand U7265 (N_7265,N_3545,N_4449);
and U7266 (N_7266,N_3660,N_4147);
nor U7267 (N_7267,N_3131,N_3132);
or U7268 (N_7268,N_4094,N_4294);
nor U7269 (N_7269,N_3549,N_3845);
and U7270 (N_7270,N_3744,N_3023);
or U7271 (N_7271,N_3765,N_3217);
nor U7272 (N_7272,N_4007,N_5583);
and U7273 (N_7273,N_5804,N_5430);
nand U7274 (N_7274,N_4444,N_5401);
and U7275 (N_7275,N_4362,N_4093);
and U7276 (N_7276,N_5154,N_5495);
nor U7277 (N_7277,N_3504,N_4953);
xnor U7278 (N_7278,N_4451,N_3244);
or U7279 (N_7279,N_5886,N_3318);
nor U7280 (N_7280,N_3297,N_3587);
nor U7281 (N_7281,N_5509,N_5477);
and U7282 (N_7282,N_5940,N_3741);
and U7283 (N_7283,N_5685,N_3312);
nand U7284 (N_7284,N_3761,N_3978);
and U7285 (N_7285,N_5713,N_4900);
or U7286 (N_7286,N_5247,N_4939);
nor U7287 (N_7287,N_3414,N_5127);
or U7288 (N_7288,N_5558,N_4105);
and U7289 (N_7289,N_4829,N_3885);
xor U7290 (N_7290,N_4031,N_4059);
or U7291 (N_7291,N_4701,N_3965);
and U7292 (N_7292,N_3671,N_3482);
or U7293 (N_7293,N_3406,N_5251);
nor U7294 (N_7294,N_4944,N_3279);
and U7295 (N_7295,N_3108,N_5634);
nand U7296 (N_7296,N_4493,N_3722);
or U7297 (N_7297,N_4600,N_5240);
nor U7298 (N_7298,N_4851,N_4637);
nand U7299 (N_7299,N_5160,N_4619);
and U7300 (N_7300,N_3760,N_5494);
nand U7301 (N_7301,N_5945,N_4626);
and U7302 (N_7302,N_5662,N_3944);
nand U7303 (N_7303,N_3246,N_3838);
and U7304 (N_7304,N_3859,N_4270);
nor U7305 (N_7305,N_3952,N_5193);
nand U7306 (N_7306,N_4661,N_5432);
nand U7307 (N_7307,N_4930,N_4972);
nor U7308 (N_7308,N_5059,N_5691);
and U7309 (N_7309,N_5479,N_4878);
or U7310 (N_7310,N_5071,N_5775);
nor U7311 (N_7311,N_3886,N_5842);
and U7312 (N_7312,N_5891,N_3192);
nor U7313 (N_7313,N_3428,N_3468);
and U7314 (N_7314,N_4911,N_4932);
nor U7315 (N_7315,N_4196,N_5131);
or U7316 (N_7316,N_5333,N_3103);
and U7317 (N_7317,N_5371,N_3079);
nand U7318 (N_7318,N_5758,N_3636);
and U7319 (N_7319,N_3717,N_3287);
nand U7320 (N_7320,N_3452,N_4223);
and U7321 (N_7321,N_3582,N_3738);
nor U7322 (N_7322,N_4392,N_4264);
nor U7323 (N_7323,N_5818,N_5282);
or U7324 (N_7324,N_4617,N_3703);
or U7325 (N_7325,N_5544,N_5875);
nand U7326 (N_7326,N_3334,N_3478);
nor U7327 (N_7327,N_5343,N_5574);
nand U7328 (N_7328,N_3852,N_5155);
nand U7329 (N_7329,N_3374,N_3058);
nor U7330 (N_7330,N_4704,N_3195);
nand U7331 (N_7331,N_4805,N_3007);
nor U7332 (N_7332,N_4990,N_4776);
nand U7333 (N_7333,N_3544,N_3606);
nor U7334 (N_7334,N_5537,N_3865);
or U7335 (N_7335,N_4075,N_3081);
or U7336 (N_7336,N_5226,N_5983);
and U7337 (N_7337,N_5470,N_4092);
and U7338 (N_7338,N_3418,N_4557);
and U7339 (N_7339,N_5152,N_4863);
or U7340 (N_7340,N_5149,N_4974);
or U7341 (N_7341,N_5488,N_3212);
nand U7342 (N_7342,N_4230,N_5938);
nor U7343 (N_7343,N_5998,N_4658);
nand U7344 (N_7344,N_5753,N_3167);
xnor U7345 (N_7345,N_4515,N_3705);
nand U7346 (N_7346,N_4298,N_3484);
nor U7347 (N_7347,N_5271,N_4817);
nor U7348 (N_7348,N_5948,N_4687);
nor U7349 (N_7349,N_4301,N_3357);
or U7350 (N_7350,N_3253,N_5726);
xnor U7351 (N_7351,N_3645,N_4980);
nand U7352 (N_7352,N_4150,N_4895);
nand U7353 (N_7353,N_4268,N_5001);
nor U7354 (N_7354,N_4833,N_5655);
nand U7355 (N_7355,N_3177,N_3210);
or U7356 (N_7356,N_4208,N_5038);
or U7357 (N_7357,N_3519,N_3531);
and U7358 (N_7358,N_4852,N_3333);
and U7359 (N_7359,N_4632,N_4373);
and U7360 (N_7360,N_4153,N_5690);
nor U7361 (N_7361,N_5407,N_5806);
nor U7362 (N_7362,N_3847,N_5776);
or U7363 (N_7363,N_4525,N_3858);
nand U7364 (N_7364,N_4349,N_4448);
or U7365 (N_7365,N_3651,N_3966);
xor U7366 (N_7366,N_5648,N_5116);
nand U7367 (N_7367,N_3325,N_5327);
and U7368 (N_7368,N_4475,N_3326);
or U7369 (N_7369,N_3251,N_3121);
and U7370 (N_7370,N_5928,N_5625);
or U7371 (N_7371,N_5203,N_5839);
nor U7372 (N_7372,N_5914,N_4028);
and U7373 (N_7373,N_5759,N_4854);
and U7374 (N_7374,N_3686,N_3610);
or U7375 (N_7375,N_5360,N_5132);
or U7376 (N_7376,N_5283,N_5041);
and U7377 (N_7377,N_5471,N_5257);
or U7378 (N_7378,N_4868,N_5971);
or U7379 (N_7379,N_5242,N_5781);
nand U7380 (N_7380,N_4308,N_5206);
and U7381 (N_7381,N_5501,N_4251);
nor U7382 (N_7382,N_4453,N_5083);
nand U7383 (N_7383,N_4724,N_4412);
or U7384 (N_7384,N_5942,N_5372);
nor U7385 (N_7385,N_5714,N_4077);
nand U7386 (N_7386,N_4258,N_3226);
nor U7387 (N_7387,N_3903,N_4182);
and U7388 (N_7388,N_4351,N_3151);
nand U7389 (N_7389,N_3938,N_4648);
and U7390 (N_7390,N_3335,N_4871);
or U7391 (N_7391,N_5687,N_5473);
nand U7392 (N_7392,N_5192,N_4746);
nand U7393 (N_7393,N_3047,N_3898);
or U7394 (N_7394,N_5002,N_5161);
nand U7395 (N_7395,N_3911,N_3673);
nand U7396 (N_7396,N_4881,N_5442);
nand U7397 (N_7397,N_5956,N_5982);
nor U7398 (N_7398,N_4651,N_3873);
or U7399 (N_7399,N_5227,N_3715);
or U7400 (N_7400,N_3247,N_3895);
nor U7401 (N_7401,N_5047,N_5267);
nand U7402 (N_7402,N_3641,N_4082);
and U7403 (N_7403,N_5550,N_5172);
nand U7404 (N_7404,N_5195,N_4622);
and U7405 (N_7405,N_3534,N_5130);
or U7406 (N_7406,N_4399,N_3799);
nand U7407 (N_7407,N_4876,N_5746);
nand U7408 (N_7408,N_4254,N_4715);
or U7409 (N_7409,N_5269,N_3777);
or U7410 (N_7410,N_4925,N_3113);
or U7411 (N_7411,N_5064,N_5863);
nand U7412 (N_7412,N_5096,N_5580);
nor U7413 (N_7413,N_4011,N_5382);
nand U7414 (N_7414,N_3539,N_4726);
and U7415 (N_7415,N_4639,N_4780);
nor U7416 (N_7416,N_4285,N_4239);
nor U7417 (N_7417,N_3887,N_5325);
nor U7418 (N_7418,N_4548,N_3390);
nand U7419 (N_7419,N_3280,N_4761);
nor U7420 (N_7420,N_3310,N_5708);
nand U7421 (N_7421,N_4014,N_3736);
or U7422 (N_7422,N_5169,N_4080);
or U7423 (N_7423,N_4921,N_3074);
nand U7424 (N_7424,N_4012,N_3928);
nand U7425 (N_7425,N_4282,N_5198);
nor U7426 (N_7426,N_4500,N_3159);
nor U7427 (N_7427,N_4713,N_3633);
or U7428 (N_7428,N_5974,N_4728);
and U7429 (N_7429,N_3013,N_4947);
or U7430 (N_7430,N_4555,N_4396);
nor U7431 (N_7431,N_4531,N_4084);
or U7432 (N_7432,N_5357,N_4901);
nor U7433 (N_7433,N_4145,N_5979);
and U7434 (N_7434,N_3479,N_3994);
nand U7435 (N_7435,N_3163,N_3276);
nand U7436 (N_7436,N_4609,N_5542);
nor U7437 (N_7437,N_3235,N_3988);
nor U7438 (N_7438,N_4137,N_3566);
nor U7439 (N_7439,N_3429,N_3635);
or U7440 (N_7440,N_5358,N_4151);
nor U7441 (N_7441,N_5752,N_4140);
nand U7442 (N_7442,N_3030,N_4021);
nand U7443 (N_7443,N_5445,N_3991);
nand U7444 (N_7444,N_5466,N_4933);
and U7445 (N_7445,N_5962,N_5885);
or U7446 (N_7446,N_5167,N_4698);
nand U7447 (N_7447,N_4165,N_5801);
nor U7448 (N_7448,N_4372,N_4354);
nor U7449 (N_7449,N_3420,N_5849);
nor U7450 (N_7450,N_4076,N_5918);
nand U7451 (N_7451,N_5475,N_5800);
and U7452 (N_7452,N_5879,N_3498);
or U7453 (N_7453,N_4783,N_4189);
or U7454 (N_7454,N_5931,N_5932);
and U7455 (N_7455,N_3972,N_3382);
nand U7456 (N_7456,N_5107,N_4403);
or U7457 (N_7457,N_4923,N_4542);
or U7458 (N_7458,N_5709,N_5197);
nor U7459 (N_7459,N_5593,N_3034);
or U7460 (N_7460,N_5985,N_5028);
or U7461 (N_7461,N_4958,N_3915);
nand U7462 (N_7462,N_3447,N_5778);
and U7463 (N_7463,N_5406,N_5865);
nand U7464 (N_7464,N_4560,N_4338);
and U7465 (N_7465,N_4368,N_5272);
and U7466 (N_7466,N_4986,N_5425);
and U7467 (N_7467,N_5235,N_5950);
nand U7468 (N_7468,N_5349,N_5664);
nand U7469 (N_7469,N_3274,N_5309);
xor U7470 (N_7470,N_4962,N_4289);
nor U7471 (N_7471,N_3491,N_4473);
or U7472 (N_7472,N_3618,N_3348);
nand U7473 (N_7473,N_5497,N_5057);
or U7474 (N_7474,N_5162,N_4959);
or U7475 (N_7475,N_5721,N_5790);
and U7476 (N_7476,N_5917,N_3655);
nor U7477 (N_7477,N_4764,N_4015);
nand U7478 (N_7478,N_5764,N_5273);
nand U7479 (N_7479,N_5671,N_3319);
nand U7480 (N_7480,N_4095,N_3126);
nand U7481 (N_7481,N_4227,N_3157);
and U7482 (N_7482,N_5767,N_5178);
nand U7483 (N_7483,N_5416,N_5578);
nor U7484 (N_7484,N_4983,N_5018);
or U7485 (N_7485,N_3236,N_3372);
nor U7486 (N_7486,N_5845,N_4688);
nand U7487 (N_7487,N_3405,N_5225);
nand U7488 (N_7488,N_5590,N_3080);
or U7489 (N_7489,N_4229,N_5231);
nand U7490 (N_7490,N_4191,N_4611);
nor U7491 (N_7491,N_5189,N_5927);
nor U7492 (N_7492,N_3494,N_5533);
nor U7493 (N_7493,N_3631,N_3575);
and U7494 (N_7494,N_4767,N_3014);
or U7495 (N_7495,N_4248,N_5058);
and U7496 (N_7496,N_4949,N_5858);
or U7497 (N_7497,N_5490,N_5317);
nor U7498 (N_7498,N_5287,N_5870);
and U7499 (N_7499,N_4889,N_3620);
or U7500 (N_7500,N_4662,N_4902);
and U7501 (N_7501,N_3842,N_5605);
or U7502 (N_7502,N_4700,N_5307);
nand U7503 (N_7503,N_4816,N_4845);
nor U7504 (N_7504,N_4993,N_4492);
or U7505 (N_7505,N_4645,N_3300);
and U7506 (N_7506,N_5522,N_5157);
nor U7507 (N_7507,N_4797,N_5221);
nand U7508 (N_7508,N_4642,N_3709);
or U7509 (N_7509,N_5711,N_3038);
nor U7510 (N_7510,N_5157,N_4680);
nand U7511 (N_7511,N_3856,N_5748);
or U7512 (N_7512,N_3765,N_4215);
or U7513 (N_7513,N_4926,N_3428);
nor U7514 (N_7514,N_3925,N_3322);
or U7515 (N_7515,N_4090,N_4611);
and U7516 (N_7516,N_4870,N_5696);
nand U7517 (N_7517,N_4447,N_3988);
or U7518 (N_7518,N_4752,N_3698);
and U7519 (N_7519,N_5900,N_4932);
nand U7520 (N_7520,N_3732,N_3335);
and U7521 (N_7521,N_3546,N_3177);
nand U7522 (N_7522,N_4999,N_3625);
and U7523 (N_7523,N_3658,N_4963);
nor U7524 (N_7524,N_3976,N_5665);
and U7525 (N_7525,N_5236,N_3219);
and U7526 (N_7526,N_3199,N_4878);
nor U7527 (N_7527,N_4418,N_4541);
and U7528 (N_7528,N_3443,N_4646);
nand U7529 (N_7529,N_3008,N_5403);
nor U7530 (N_7530,N_5284,N_5159);
and U7531 (N_7531,N_4283,N_5777);
nor U7532 (N_7532,N_3036,N_4893);
nor U7533 (N_7533,N_4365,N_4466);
and U7534 (N_7534,N_3193,N_3195);
nand U7535 (N_7535,N_3084,N_5863);
nor U7536 (N_7536,N_3846,N_4678);
nor U7537 (N_7537,N_3709,N_3202);
and U7538 (N_7538,N_3845,N_5214);
nor U7539 (N_7539,N_5351,N_3228);
or U7540 (N_7540,N_4927,N_3191);
and U7541 (N_7541,N_5280,N_3248);
nor U7542 (N_7542,N_3444,N_5551);
or U7543 (N_7543,N_3784,N_3856);
nor U7544 (N_7544,N_3679,N_3304);
and U7545 (N_7545,N_3837,N_3768);
nand U7546 (N_7546,N_4407,N_5671);
or U7547 (N_7547,N_3516,N_3664);
nand U7548 (N_7548,N_4784,N_5161);
and U7549 (N_7549,N_4798,N_5911);
or U7550 (N_7550,N_4862,N_4766);
or U7551 (N_7551,N_5940,N_4870);
nand U7552 (N_7552,N_3773,N_3655);
or U7553 (N_7553,N_3810,N_5645);
nor U7554 (N_7554,N_4005,N_3325);
nor U7555 (N_7555,N_5529,N_4343);
nand U7556 (N_7556,N_5545,N_5135);
nand U7557 (N_7557,N_3038,N_3097);
or U7558 (N_7558,N_4654,N_3803);
nor U7559 (N_7559,N_4624,N_3942);
or U7560 (N_7560,N_5028,N_5475);
or U7561 (N_7561,N_3277,N_5772);
or U7562 (N_7562,N_4511,N_3961);
nor U7563 (N_7563,N_5174,N_4318);
and U7564 (N_7564,N_4651,N_3324);
nand U7565 (N_7565,N_4042,N_5356);
nor U7566 (N_7566,N_3540,N_4017);
or U7567 (N_7567,N_4237,N_3002);
and U7568 (N_7568,N_3983,N_5763);
nand U7569 (N_7569,N_5445,N_3402);
and U7570 (N_7570,N_4167,N_4851);
and U7571 (N_7571,N_4012,N_4364);
nor U7572 (N_7572,N_4165,N_3406);
nor U7573 (N_7573,N_5898,N_4807);
nand U7574 (N_7574,N_5264,N_4526);
and U7575 (N_7575,N_4776,N_5828);
or U7576 (N_7576,N_3435,N_4050);
or U7577 (N_7577,N_3225,N_3527);
and U7578 (N_7578,N_5032,N_3547);
nor U7579 (N_7579,N_5648,N_4979);
and U7580 (N_7580,N_3360,N_5422);
nor U7581 (N_7581,N_4605,N_4401);
nand U7582 (N_7582,N_4013,N_3736);
nor U7583 (N_7583,N_3877,N_3682);
nor U7584 (N_7584,N_5784,N_4444);
nor U7585 (N_7585,N_4254,N_5235);
nand U7586 (N_7586,N_5324,N_5287);
or U7587 (N_7587,N_4830,N_5163);
nand U7588 (N_7588,N_3524,N_3788);
or U7589 (N_7589,N_3196,N_3515);
nand U7590 (N_7590,N_3955,N_4532);
nand U7591 (N_7591,N_3146,N_4716);
or U7592 (N_7592,N_3018,N_5016);
and U7593 (N_7593,N_3210,N_5514);
nor U7594 (N_7594,N_4828,N_4722);
and U7595 (N_7595,N_5252,N_4856);
nor U7596 (N_7596,N_5451,N_3302);
nand U7597 (N_7597,N_4286,N_3055);
nor U7598 (N_7598,N_3839,N_4248);
nand U7599 (N_7599,N_3956,N_5140);
nand U7600 (N_7600,N_4629,N_3097);
or U7601 (N_7601,N_4320,N_5004);
nor U7602 (N_7602,N_5532,N_4610);
and U7603 (N_7603,N_5187,N_5951);
or U7604 (N_7604,N_4025,N_5008);
nand U7605 (N_7605,N_5738,N_3374);
nor U7606 (N_7606,N_3796,N_5194);
nand U7607 (N_7607,N_3586,N_3244);
nand U7608 (N_7608,N_5002,N_5530);
and U7609 (N_7609,N_3141,N_4665);
or U7610 (N_7610,N_4504,N_3404);
nand U7611 (N_7611,N_3443,N_5678);
nor U7612 (N_7612,N_3737,N_3918);
nand U7613 (N_7613,N_3523,N_5273);
or U7614 (N_7614,N_4728,N_5328);
or U7615 (N_7615,N_4368,N_4025);
or U7616 (N_7616,N_5755,N_4020);
nor U7617 (N_7617,N_5733,N_4407);
nor U7618 (N_7618,N_5612,N_4630);
and U7619 (N_7619,N_5943,N_4482);
and U7620 (N_7620,N_5244,N_4092);
or U7621 (N_7621,N_3336,N_5729);
or U7622 (N_7622,N_3796,N_3557);
or U7623 (N_7623,N_3115,N_4709);
nand U7624 (N_7624,N_5616,N_4712);
or U7625 (N_7625,N_3947,N_4698);
nor U7626 (N_7626,N_3740,N_4687);
nor U7627 (N_7627,N_3057,N_4339);
or U7628 (N_7628,N_3995,N_5958);
and U7629 (N_7629,N_5699,N_5429);
and U7630 (N_7630,N_5657,N_4090);
nand U7631 (N_7631,N_4153,N_5530);
nor U7632 (N_7632,N_3774,N_5230);
and U7633 (N_7633,N_3080,N_5705);
or U7634 (N_7634,N_5631,N_4870);
nand U7635 (N_7635,N_4169,N_3334);
nand U7636 (N_7636,N_5044,N_5053);
or U7637 (N_7637,N_3878,N_5533);
nand U7638 (N_7638,N_4754,N_4579);
nor U7639 (N_7639,N_5486,N_4911);
and U7640 (N_7640,N_3799,N_3002);
and U7641 (N_7641,N_5652,N_3500);
or U7642 (N_7642,N_5224,N_3310);
or U7643 (N_7643,N_4557,N_4831);
nor U7644 (N_7644,N_5958,N_5183);
nand U7645 (N_7645,N_5718,N_3413);
nand U7646 (N_7646,N_4092,N_3152);
and U7647 (N_7647,N_3692,N_3849);
or U7648 (N_7648,N_4347,N_5361);
nand U7649 (N_7649,N_3705,N_3685);
or U7650 (N_7650,N_4602,N_4018);
nor U7651 (N_7651,N_4807,N_4939);
nand U7652 (N_7652,N_4645,N_4539);
nor U7653 (N_7653,N_4668,N_3746);
or U7654 (N_7654,N_5646,N_3843);
nor U7655 (N_7655,N_5455,N_4638);
nand U7656 (N_7656,N_4180,N_5138);
nor U7657 (N_7657,N_5548,N_5035);
nor U7658 (N_7658,N_3192,N_3185);
nand U7659 (N_7659,N_3857,N_4389);
nand U7660 (N_7660,N_4017,N_4513);
or U7661 (N_7661,N_4407,N_5481);
or U7662 (N_7662,N_3222,N_5393);
and U7663 (N_7663,N_4716,N_4181);
or U7664 (N_7664,N_4946,N_4229);
nor U7665 (N_7665,N_3901,N_4823);
and U7666 (N_7666,N_4967,N_4925);
nor U7667 (N_7667,N_5574,N_4498);
nand U7668 (N_7668,N_5140,N_3001);
or U7669 (N_7669,N_4899,N_4948);
nor U7670 (N_7670,N_5476,N_5700);
nand U7671 (N_7671,N_5172,N_3966);
nor U7672 (N_7672,N_3486,N_5338);
or U7673 (N_7673,N_5118,N_5267);
or U7674 (N_7674,N_5798,N_5996);
nor U7675 (N_7675,N_3147,N_4880);
nor U7676 (N_7676,N_5466,N_4051);
or U7677 (N_7677,N_4927,N_4095);
nor U7678 (N_7678,N_4274,N_4684);
nor U7679 (N_7679,N_3981,N_3715);
and U7680 (N_7680,N_5576,N_4672);
nand U7681 (N_7681,N_4573,N_5374);
nor U7682 (N_7682,N_5346,N_4022);
nand U7683 (N_7683,N_5492,N_3431);
or U7684 (N_7684,N_5643,N_3157);
nand U7685 (N_7685,N_3792,N_4426);
nand U7686 (N_7686,N_3283,N_5316);
and U7687 (N_7687,N_4529,N_5513);
nor U7688 (N_7688,N_5917,N_3239);
or U7689 (N_7689,N_3996,N_5036);
or U7690 (N_7690,N_4874,N_5503);
or U7691 (N_7691,N_3633,N_4047);
nor U7692 (N_7692,N_3466,N_4941);
nand U7693 (N_7693,N_5334,N_5661);
nand U7694 (N_7694,N_4676,N_3447);
nand U7695 (N_7695,N_4640,N_5418);
and U7696 (N_7696,N_5098,N_3691);
or U7697 (N_7697,N_5527,N_5829);
nor U7698 (N_7698,N_3911,N_4555);
nand U7699 (N_7699,N_3687,N_3324);
nand U7700 (N_7700,N_5682,N_3357);
nand U7701 (N_7701,N_3867,N_3309);
or U7702 (N_7702,N_5442,N_5691);
nor U7703 (N_7703,N_5580,N_5650);
or U7704 (N_7704,N_4103,N_3151);
nor U7705 (N_7705,N_5953,N_5526);
nand U7706 (N_7706,N_4158,N_3919);
nor U7707 (N_7707,N_5556,N_3321);
nand U7708 (N_7708,N_5628,N_3360);
and U7709 (N_7709,N_3008,N_4793);
and U7710 (N_7710,N_5733,N_3742);
and U7711 (N_7711,N_3328,N_4504);
or U7712 (N_7712,N_3384,N_4013);
nor U7713 (N_7713,N_5406,N_3188);
nor U7714 (N_7714,N_3927,N_5859);
nand U7715 (N_7715,N_4136,N_4500);
nor U7716 (N_7716,N_3574,N_3087);
or U7717 (N_7717,N_3981,N_4088);
nor U7718 (N_7718,N_3280,N_4110);
nand U7719 (N_7719,N_3600,N_5897);
nor U7720 (N_7720,N_4112,N_4656);
or U7721 (N_7721,N_4964,N_3144);
and U7722 (N_7722,N_4028,N_3103);
nand U7723 (N_7723,N_5578,N_5179);
nor U7724 (N_7724,N_3107,N_3182);
or U7725 (N_7725,N_4295,N_5185);
nand U7726 (N_7726,N_5629,N_4843);
and U7727 (N_7727,N_3657,N_4364);
nand U7728 (N_7728,N_4364,N_4150);
nand U7729 (N_7729,N_4930,N_3836);
nor U7730 (N_7730,N_4960,N_4323);
or U7731 (N_7731,N_3934,N_3464);
and U7732 (N_7732,N_5021,N_5906);
and U7733 (N_7733,N_5680,N_4970);
nor U7734 (N_7734,N_3236,N_5543);
or U7735 (N_7735,N_3597,N_4677);
nor U7736 (N_7736,N_4272,N_3762);
or U7737 (N_7737,N_3104,N_4864);
or U7738 (N_7738,N_5602,N_5849);
xor U7739 (N_7739,N_5342,N_5814);
nand U7740 (N_7740,N_5378,N_5410);
or U7741 (N_7741,N_4612,N_4501);
nand U7742 (N_7742,N_3486,N_4942);
and U7743 (N_7743,N_3941,N_4591);
and U7744 (N_7744,N_4692,N_5204);
nand U7745 (N_7745,N_3528,N_3199);
nand U7746 (N_7746,N_3942,N_5899);
nand U7747 (N_7747,N_4923,N_4964);
or U7748 (N_7748,N_5218,N_4209);
nand U7749 (N_7749,N_3586,N_5676);
and U7750 (N_7750,N_3118,N_4108);
nand U7751 (N_7751,N_4886,N_3931);
or U7752 (N_7752,N_5738,N_4503);
nand U7753 (N_7753,N_5115,N_3267);
nor U7754 (N_7754,N_3293,N_5396);
and U7755 (N_7755,N_4634,N_3588);
nand U7756 (N_7756,N_3214,N_5126);
and U7757 (N_7757,N_3513,N_3693);
or U7758 (N_7758,N_5706,N_4890);
nand U7759 (N_7759,N_3486,N_5394);
and U7760 (N_7760,N_3603,N_3470);
and U7761 (N_7761,N_3940,N_5008);
and U7762 (N_7762,N_5320,N_4563);
and U7763 (N_7763,N_5794,N_4038);
nor U7764 (N_7764,N_3907,N_5482);
or U7765 (N_7765,N_4768,N_3376);
or U7766 (N_7766,N_5756,N_4535);
nor U7767 (N_7767,N_3784,N_5012);
or U7768 (N_7768,N_5584,N_5957);
nand U7769 (N_7769,N_5490,N_5565);
and U7770 (N_7770,N_5439,N_3469);
and U7771 (N_7771,N_5032,N_5376);
or U7772 (N_7772,N_5259,N_3751);
nor U7773 (N_7773,N_5406,N_5852);
nor U7774 (N_7774,N_4391,N_4503);
nand U7775 (N_7775,N_3417,N_3479);
nand U7776 (N_7776,N_5687,N_4117);
and U7777 (N_7777,N_4055,N_4115);
nor U7778 (N_7778,N_3602,N_5834);
and U7779 (N_7779,N_4880,N_5725);
nor U7780 (N_7780,N_3162,N_3453);
nand U7781 (N_7781,N_5174,N_3567);
or U7782 (N_7782,N_5484,N_4787);
and U7783 (N_7783,N_5485,N_5803);
nand U7784 (N_7784,N_5944,N_3590);
nand U7785 (N_7785,N_3722,N_5803);
or U7786 (N_7786,N_3804,N_5367);
nor U7787 (N_7787,N_5131,N_5428);
or U7788 (N_7788,N_4044,N_3838);
and U7789 (N_7789,N_4031,N_3240);
or U7790 (N_7790,N_4456,N_5560);
and U7791 (N_7791,N_3771,N_3212);
nand U7792 (N_7792,N_4717,N_3700);
nand U7793 (N_7793,N_3328,N_4802);
nand U7794 (N_7794,N_5290,N_4996);
nor U7795 (N_7795,N_3428,N_4279);
or U7796 (N_7796,N_5279,N_3501);
and U7797 (N_7797,N_3640,N_3229);
nand U7798 (N_7798,N_5947,N_3581);
nor U7799 (N_7799,N_3383,N_5900);
nor U7800 (N_7800,N_4392,N_4949);
nor U7801 (N_7801,N_5627,N_5075);
or U7802 (N_7802,N_4365,N_4408);
nor U7803 (N_7803,N_5046,N_5359);
nor U7804 (N_7804,N_4896,N_5093);
and U7805 (N_7805,N_3673,N_5173);
nand U7806 (N_7806,N_3503,N_5456);
nand U7807 (N_7807,N_3371,N_4562);
nor U7808 (N_7808,N_4173,N_4704);
and U7809 (N_7809,N_3658,N_5671);
and U7810 (N_7810,N_5894,N_3295);
or U7811 (N_7811,N_4723,N_5284);
xor U7812 (N_7812,N_5246,N_4536);
nor U7813 (N_7813,N_3295,N_5387);
and U7814 (N_7814,N_5953,N_3016);
nor U7815 (N_7815,N_4875,N_4252);
and U7816 (N_7816,N_3133,N_3567);
nor U7817 (N_7817,N_3395,N_3979);
and U7818 (N_7818,N_3644,N_3839);
nor U7819 (N_7819,N_3219,N_4316);
and U7820 (N_7820,N_3157,N_4427);
nor U7821 (N_7821,N_4327,N_5847);
or U7822 (N_7822,N_3553,N_5531);
nor U7823 (N_7823,N_4660,N_4996);
or U7824 (N_7824,N_5162,N_4008);
nor U7825 (N_7825,N_4875,N_4233);
or U7826 (N_7826,N_5438,N_5836);
nand U7827 (N_7827,N_3261,N_5155);
nor U7828 (N_7828,N_3060,N_5749);
or U7829 (N_7829,N_5316,N_4872);
and U7830 (N_7830,N_4677,N_5732);
nand U7831 (N_7831,N_3694,N_3201);
and U7832 (N_7832,N_5591,N_3445);
and U7833 (N_7833,N_5995,N_4950);
or U7834 (N_7834,N_3087,N_4916);
or U7835 (N_7835,N_3360,N_4453);
nor U7836 (N_7836,N_4156,N_4757);
or U7837 (N_7837,N_5464,N_5972);
and U7838 (N_7838,N_5023,N_3057);
nor U7839 (N_7839,N_3232,N_4898);
nor U7840 (N_7840,N_4363,N_4589);
nand U7841 (N_7841,N_5357,N_3652);
nand U7842 (N_7842,N_5863,N_4237);
or U7843 (N_7843,N_4451,N_3022);
or U7844 (N_7844,N_3486,N_3099);
or U7845 (N_7845,N_3101,N_5124);
nand U7846 (N_7846,N_4191,N_4072);
and U7847 (N_7847,N_5456,N_5250);
nor U7848 (N_7848,N_5217,N_3590);
nand U7849 (N_7849,N_3625,N_3830);
nand U7850 (N_7850,N_4233,N_5220);
and U7851 (N_7851,N_3879,N_3545);
and U7852 (N_7852,N_4675,N_5821);
and U7853 (N_7853,N_3864,N_5170);
nand U7854 (N_7854,N_4715,N_4020);
nand U7855 (N_7855,N_5239,N_4335);
nor U7856 (N_7856,N_5418,N_4050);
nand U7857 (N_7857,N_3436,N_3741);
nand U7858 (N_7858,N_3571,N_4659);
or U7859 (N_7859,N_4629,N_3171);
or U7860 (N_7860,N_3088,N_4258);
nand U7861 (N_7861,N_5924,N_3537);
nor U7862 (N_7862,N_5632,N_3499);
and U7863 (N_7863,N_5892,N_3370);
or U7864 (N_7864,N_4130,N_5110);
nand U7865 (N_7865,N_3822,N_4668);
nor U7866 (N_7866,N_5589,N_4020);
nand U7867 (N_7867,N_3138,N_5623);
or U7868 (N_7868,N_3182,N_3926);
and U7869 (N_7869,N_4115,N_5502);
and U7870 (N_7870,N_3444,N_3627);
and U7871 (N_7871,N_5814,N_4962);
or U7872 (N_7872,N_5987,N_4819);
nand U7873 (N_7873,N_4369,N_4606);
or U7874 (N_7874,N_4912,N_3169);
nor U7875 (N_7875,N_5259,N_4740);
nand U7876 (N_7876,N_4594,N_5247);
nand U7877 (N_7877,N_3849,N_3758);
and U7878 (N_7878,N_3106,N_4060);
nand U7879 (N_7879,N_4093,N_3153);
nor U7880 (N_7880,N_5801,N_4758);
or U7881 (N_7881,N_5675,N_5010);
and U7882 (N_7882,N_3644,N_4437);
nand U7883 (N_7883,N_5769,N_4815);
nor U7884 (N_7884,N_5852,N_5784);
nand U7885 (N_7885,N_5889,N_3160);
or U7886 (N_7886,N_5106,N_3228);
nand U7887 (N_7887,N_4351,N_3611);
nand U7888 (N_7888,N_5157,N_5614);
nor U7889 (N_7889,N_3518,N_4801);
and U7890 (N_7890,N_5835,N_4211);
and U7891 (N_7891,N_4533,N_4716);
or U7892 (N_7892,N_3093,N_4088);
nand U7893 (N_7893,N_3353,N_5803);
nor U7894 (N_7894,N_3979,N_4863);
nand U7895 (N_7895,N_3896,N_5747);
nor U7896 (N_7896,N_3396,N_3552);
and U7897 (N_7897,N_3451,N_3141);
or U7898 (N_7898,N_3009,N_4439);
nor U7899 (N_7899,N_3041,N_4276);
nor U7900 (N_7900,N_4217,N_4101);
nand U7901 (N_7901,N_5897,N_5923);
nor U7902 (N_7902,N_3013,N_3578);
and U7903 (N_7903,N_3096,N_5545);
nor U7904 (N_7904,N_4010,N_5658);
nand U7905 (N_7905,N_4644,N_4059);
nand U7906 (N_7906,N_5241,N_3414);
and U7907 (N_7907,N_4729,N_3433);
nor U7908 (N_7908,N_3919,N_5268);
and U7909 (N_7909,N_3661,N_3804);
or U7910 (N_7910,N_5037,N_3457);
nor U7911 (N_7911,N_3846,N_5199);
nor U7912 (N_7912,N_3770,N_3439);
nor U7913 (N_7913,N_4278,N_3671);
or U7914 (N_7914,N_4032,N_3953);
and U7915 (N_7915,N_5750,N_4151);
and U7916 (N_7916,N_5517,N_4619);
and U7917 (N_7917,N_5883,N_3745);
nand U7918 (N_7918,N_5468,N_5472);
or U7919 (N_7919,N_3747,N_4354);
nand U7920 (N_7920,N_4934,N_4627);
nor U7921 (N_7921,N_4648,N_5755);
and U7922 (N_7922,N_3211,N_4803);
nor U7923 (N_7923,N_3091,N_4964);
and U7924 (N_7924,N_4996,N_3368);
nor U7925 (N_7925,N_5959,N_3872);
or U7926 (N_7926,N_4123,N_3601);
and U7927 (N_7927,N_3156,N_4393);
or U7928 (N_7928,N_3900,N_3798);
nand U7929 (N_7929,N_3718,N_3201);
and U7930 (N_7930,N_4167,N_5326);
nand U7931 (N_7931,N_5595,N_5278);
nor U7932 (N_7932,N_5015,N_5946);
xnor U7933 (N_7933,N_3523,N_3560);
nand U7934 (N_7934,N_5428,N_3763);
and U7935 (N_7935,N_5948,N_3000);
and U7936 (N_7936,N_5668,N_3902);
and U7937 (N_7937,N_3713,N_5535);
and U7938 (N_7938,N_3807,N_4472);
and U7939 (N_7939,N_3741,N_3159);
nand U7940 (N_7940,N_4853,N_4979);
nor U7941 (N_7941,N_4566,N_5469);
nand U7942 (N_7942,N_3061,N_5457);
or U7943 (N_7943,N_3622,N_3567);
and U7944 (N_7944,N_3876,N_3181);
nand U7945 (N_7945,N_5556,N_3259);
or U7946 (N_7946,N_4296,N_5062);
nor U7947 (N_7947,N_3132,N_5997);
or U7948 (N_7948,N_4293,N_3269);
and U7949 (N_7949,N_4875,N_3652);
and U7950 (N_7950,N_3417,N_5244);
nand U7951 (N_7951,N_3117,N_5581);
and U7952 (N_7952,N_3273,N_4669);
or U7953 (N_7953,N_3902,N_3374);
or U7954 (N_7954,N_3489,N_3375);
and U7955 (N_7955,N_5503,N_3414);
or U7956 (N_7956,N_5553,N_5123);
and U7957 (N_7957,N_4302,N_3253);
nor U7958 (N_7958,N_5523,N_5982);
nor U7959 (N_7959,N_3069,N_4668);
nand U7960 (N_7960,N_5639,N_3957);
and U7961 (N_7961,N_5307,N_5948);
nand U7962 (N_7962,N_4380,N_5444);
nor U7963 (N_7963,N_4556,N_4350);
nor U7964 (N_7964,N_4250,N_4213);
nand U7965 (N_7965,N_4793,N_4731);
or U7966 (N_7966,N_5780,N_4205);
or U7967 (N_7967,N_3815,N_4531);
nor U7968 (N_7968,N_3620,N_4701);
or U7969 (N_7969,N_3401,N_4241);
and U7970 (N_7970,N_3790,N_3631);
and U7971 (N_7971,N_3617,N_3849);
nor U7972 (N_7972,N_3078,N_5255);
nand U7973 (N_7973,N_4232,N_4274);
nor U7974 (N_7974,N_5923,N_3682);
and U7975 (N_7975,N_3962,N_5078);
or U7976 (N_7976,N_5771,N_5510);
and U7977 (N_7977,N_5293,N_3953);
nand U7978 (N_7978,N_4808,N_5356);
or U7979 (N_7979,N_5651,N_3618);
nor U7980 (N_7980,N_5073,N_5204);
and U7981 (N_7981,N_5415,N_5934);
nand U7982 (N_7982,N_4913,N_5609);
nor U7983 (N_7983,N_5490,N_3143);
or U7984 (N_7984,N_3185,N_4969);
xnor U7985 (N_7985,N_3113,N_5086);
and U7986 (N_7986,N_5363,N_5691);
nor U7987 (N_7987,N_3671,N_4440);
and U7988 (N_7988,N_3932,N_3554);
nor U7989 (N_7989,N_3646,N_5745);
or U7990 (N_7990,N_4106,N_3423);
and U7991 (N_7991,N_5632,N_4570);
nor U7992 (N_7992,N_5229,N_5845);
nor U7993 (N_7993,N_5221,N_4497);
nor U7994 (N_7994,N_4630,N_4303);
nor U7995 (N_7995,N_3637,N_5425);
nand U7996 (N_7996,N_5276,N_5647);
nand U7997 (N_7997,N_4651,N_4608);
nand U7998 (N_7998,N_4715,N_3069);
or U7999 (N_7999,N_5503,N_4738);
nand U8000 (N_8000,N_5548,N_3452);
or U8001 (N_8001,N_3316,N_4407);
nand U8002 (N_8002,N_5759,N_3490);
nand U8003 (N_8003,N_3867,N_5198);
nand U8004 (N_8004,N_4918,N_5848);
and U8005 (N_8005,N_3064,N_5494);
and U8006 (N_8006,N_4000,N_4510);
and U8007 (N_8007,N_3562,N_3879);
or U8008 (N_8008,N_3205,N_4392);
nor U8009 (N_8009,N_4440,N_5310);
or U8010 (N_8010,N_4881,N_5761);
nor U8011 (N_8011,N_3127,N_5332);
or U8012 (N_8012,N_5022,N_5704);
nor U8013 (N_8013,N_4842,N_4870);
nand U8014 (N_8014,N_5651,N_5283);
nor U8015 (N_8015,N_3904,N_4112);
or U8016 (N_8016,N_3722,N_4713);
nand U8017 (N_8017,N_5584,N_3913);
and U8018 (N_8018,N_3191,N_4500);
or U8019 (N_8019,N_3013,N_3315);
nor U8020 (N_8020,N_3720,N_5166);
or U8021 (N_8021,N_4020,N_5168);
nor U8022 (N_8022,N_5126,N_3018);
nor U8023 (N_8023,N_5240,N_4637);
nor U8024 (N_8024,N_5292,N_4281);
nor U8025 (N_8025,N_5373,N_4837);
or U8026 (N_8026,N_3887,N_5543);
nand U8027 (N_8027,N_3960,N_3332);
nand U8028 (N_8028,N_4047,N_5404);
and U8029 (N_8029,N_5875,N_4668);
nand U8030 (N_8030,N_5245,N_3492);
and U8031 (N_8031,N_3987,N_4268);
nor U8032 (N_8032,N_5203,N_3521);
and U8033 (N_8033,N_3634,N_5992);
nand U8034 (N_8034,N_5934,N_4358);
nor U8035 (N_8035,N_4320,N_5782);
nand U8036 (N_8036,N_3225,N_4824);
nor U8037 (N_8037,N_5366,N_5204);
nor U8038 (N_8038,N_5573,N_3837);
or U8039 (N_8039,N_4382,N_4474);
nor U8040 (N_8040,N_5533,N_3790);
nand U8041 (N_8041,N_5398,N_4470);
nand U8042 (N_8042,N_4259,N_5131);
or U8043 (N_8043,N_4263,N_3072);
nand U8044 (N_8044,N_5064,N_4165);
and U8045 (N_8045,N_4956,N_3752);
and U8046 (N_8046,N_5852,N_4586);
nand U8047 (N_8047,N_4820,N_3094);
or U8048 (N_8048,N_5454,N_5075);
nor U8049 (N_8049,N_3618,N_4503);
nand U8050 (N_8050,N_3324,N_4962);
nand U8051 (N_8051,N_4578,N_5245);
nor U8052 (N_8052,N_4114,N_5466);
or U8053 (N_8053,N_4365,N_4822);
xor U8054 (N_8054,N_3707,N_4868);
and U8055 (N_8055,N_3648,N_4828);
nor U8056 (N_8056,N_4046,N_5065);
nand U8057 (N_8057,N_3233,N_3164);
nand U8058 (N_8058,N_4126,N_3259);
or U8059 (N_8059,N_4866,N_3886);
nand U8060 (N_8060,N_3716,N_4302);
nor U8061 (N_8061,N_4043,N_5223);
nand U8062 (N_8062,N_4367,N_4038);
and U8063 (N_8063,N_3953,N_3667);
nand U8064 (N_8064,N_4142,N_5186);
and U8065 (N_8065,N_3591,N_3729);
or U8066 (N_8066,N_5059,N_3940);
xnor U8067 (N_8067,N_4133,N_4443);
or U8068 (N_8068,N_5258,N_3042);
nand U8069 (N_8069,N_4165,N_4263);
nor U8070 (N_8070,N_5182,N_3896);
or U8071 (N_8071,N_4632,N_4159);
nor U8072 (N_8072,N_5573,N_4747);
and U8073 (N_8073,N_3409,N_4840);
nand U8074 (N_8074,N_3322,N_3437);
nand U8075 (N_8075,N_3712,N_4645);
and U8076 (N_8076,N_4976,N_5093);
nand U8077 (N_8077,N_5199,N_5292);
nor U8078 (N_8078,N_5017,N_3501);
nor U8079 (N_8079,N_5960,N_4555);
and U8080 (N_8080,N_4456,N_3099);
nand U8081 (N_8081,N_4719,N_4512);
nand U8082 (N_8082,N_5099,N_4012);
nand U8083 (N_8083,N_5465,N_3666);
nand U8084 (N_8084,N_5378,N_4216);
or U8085 (N_8085,N_5912,N_4639);
nor U8086 (N_8086,N_4760,N_5282);
and U8087 (N_8087,N_3538,N_5997);
nor U8088 (N_8088,N_4567,N_4872);
nand U8089 (N_8089,N_5333,N_3774);
and U8090 (N_8090,N_4727,N_5474);
and U8091 (N_8091,N_4254,N_5373);
nand U8092 (N_8092,N_5297,N_5730);
nand U8093 (N_8093,N_3437,N_3890);
nor U8094 (N_8094,N_4440,N_4547);
and U8095 (N_8095,N_4551,N_4058);
nand U8096 (N_8096,N_5352,N_4156);
nand U8097 (N_8097,N_3944,N_5639);
nor U8098 (N_8098,N_4354,N_4051);
and U8099 (N_8099,N_5033,N_5613);
nor U8100 (N_8100,N_3080,N_3388);
nand U8101 (N_8101,N_4948,N_3049);
or U8102 (N_8102,N_3652,N_4015);
and U8103 (N_8103,N_5660,N_4085);
and U8104 (N_8104,N_4459,N_4008);
nand U8105 (N_8105,N_3714,N_5017);
or U8106 (N_8106,N_4035,N_5932);
and U8107 (N_8107,N_4194,N_3364);
and U8108 (N_8108,N_4425,N_3787);
nand U8109 (N_8109,N_3157,N_5948);
or U8110 (N_8110,N_4633,N_5201);
nand U8111 (N_8111,N_4232,N_5316);
nor U8112 (N_8112,N_4813,N_4945);
and U8113 (N_8113,N_5468,N_4324);
nor U8114 (N_8114,N_3634,N_5100);
nor U8115 (N_8115,N_3887,N_4771);
nand U8116 (N_8116,N_3829,N_4415);
or U8117 (N_8117,N_4166,N_4481);
or U8118 (N_8118,N_3784,N_4179);
and U8119 (N_8119,N_5039,N_5329);
or U8120 (N_8120,N_4039,N_5946);
or U8121 (N_8121,N_3736,N_3569);
or U8122 (N_8122,N_5844,N_5512);
nor U8123 (N_8123,N_4931,N_5299);
nand U8124 (N_8124,N_3231,N_4116);
xnor U8125 (N_8125,N_4320,N_4075);
nor U8126 (N_8126,N_5321,N_3563);
nand U8127 (N_8127,N_3531,N_5682);
and U8128 (N_8128,N_4259,N_3390);
nand U8129 (N_8129,N_3057,N_4851);
or U8130 (N_8130,N_5591,N_5907);
nand U8131 (N_8131,N_4503,N_3240);
or U8132 (N_8132,N_5322,N_3137);
and U8133 (N_8133,N_4774,N_5742);
nor U8134 (N_8134,N_3847,N_4193);
and U8135 (N_8135,N_5108,N_4807);
and U8136 (N_8136,N_3051,N_4819);
and U8137 (N_8137,N_5714,N_3354);
or U8138 (N_8138,N_3576,N_3328);
nand U8139 (N_8139,N_3622,N_3501);
and U8140 (N_8140,N_5589,N_3661);
or U8141 (N_8141,N_3855,N_4398);
and U8142 (N_8142,N_5287,N_3854);
nand U8143 (N_8143,N_4106,N_3030);
and U8144 (N_8144,N_3744,N_3303);
nor U8145 (N_8145,N_4009,N_4628);
xnor U8146 (N_8146,N_4795,N_3291);
nor U8147 (N_8147,N_5117,N_4754);
and U8148 (N_8148,N_5199,N_4120);
or U8149 (N_8149,N_3474,N_4659);
or U8150 (N_8150,N_5838,N_3086);
nor U8151 (N_8151,N_4485,N_5018);
and U8152 (N_8152,N_3302,N_4336);
and U8153 (N_8153,N_5549,N_3631);
nor U8154 (N_8154,N_4535,N_4502);
or U8155 (N_8155,N_4638,N_3987);
or U8156 (N_8156,N_5458,N_5253);
nand U8157 (N_8157,N_5135,N_5468);
nand U8158 (N_8158,N_4419,N_5991);
nor U8159 (N_8159,N_4642,N_3401);
nand U8160 (N_8160,N_4844,N_5515);
nand U8161 (N_8161,N_5700,N_4992);
nand U8162 (N_8162,N_4421,N_3499);
nand U8163 (N_8163,N_4966,N_4476);
nor U8164 (N_8164,N_4909,N_3466);
and U8165 (N_8165,N_5154,N_4624);
nand U8166 (N_8166,N_3385,N_3679);
nor U8167 (N_8167,N_3215,N_4749);
and U8168 (N_8168,N_5602,N_5697);
or U8169 (N_8169,N_4955,N_4081);
and U8170 (N_8170,N_3960,N_5726);
or U8171 (N_8171,N_4659,N_3160);
or U8172 (N_8172,N_3966,N_3256);
nor U8173 (N_8173,N_3568,N_4249);
and U8174 (N_8174,N_4541,N_5594);
and U8175 (N_8175,N_3276,N_3242);
nand U8176 (N_8176,N_3825,N_5664);
nor U8177 (N_8177,N_5209,N_5574);
nor U8178 (N_8178,N_5880,N_3596);
or U8179 (N_8179,N_5572,N_4867);
and U8180 (N_8180,N_3907,N_4437);
or U8181 (N_8181,N_5305,N_4114);
nand U8182 (N_8182,N_4119,N_5118);
nand U8183 (N_8183,N_5911,N_3666);
or U8184 (N_8184,N_5897,N_3106);
and U8185 (N_8185,N_4559,N_4577);
or U8186 (N_8186,N_3714,N_3978);
or U8187 (N_8187,N_4640,N_5040);
or U8188 (N_8188,N_3294,N_4312);
nor U8189 (N_8189,N_5524,N_5667);
and U8190 (N_8190,N_3669,N_5238);
and U8191 (N_8191,N_5428,N_4924);
or U8192 (N_8192,N_4892,N_4787);
and U8193 (N_8193,N_4323,N_3600);
nor U8194 (N_8194,N_4782,N_5453);
or U8195 (N_8195,N_4213,N_4085);
nor U8196 (N_8196,N_5149,N_3000);
and U8197 (N_8197,N_4683,N_3220);
or U8198 (N_8198,N_4996,N_3631);
and U8199 (N_8199,N_3955,N_3738);
and U8200 (N_8200,N_3987,N_4448);
nor U8201 (N_8201,N_4595,N_4545);
nor U8202 (N_8202,N_4056,N_3638);
nand U8203 (N_8203,N_4520,N_3161);
or U8204 (N_8204,N_5044,N_3844);
or U8205 (N_8205,N_3751,N_4612);
and U8206 (N_8206,N_3239,N_5329);
nor U8207 (N_8207,N_3472,N_5813);
and U8208 (N_8208,N_4009,N_5042);
nor U8209 (N_8209,N_5050,N_5462);
xor U8210 (N_8210,N_3475,N_4480);
and U8211 (N_8211,N_3318,N_5664);
or U8212 (N_8212,N_3181,N_4484);
or U8213 (N_8213,N_3092,N_5022);
or U8214 (N_8214,N_3899,N_4736);
and U8215 (N_8215,N_5817,N_5708);
or U8216 (N_8216,N_3933,N_3105);
nand U8217 (N_8217,N_4580,N_4304);
and U8218 (N_8218,N_5130,N_4842);
or U8219 (N_8219,N_5060,N_4304);
and U8220 (N_8220,N_5901,N_4539);
or U8221 (N_8221,N_4468,N_5994);
nand U8222 (N_8222,N_5863,N_5566);
nand U8223 (N_8223,N_3865,N_3384);
and U8224 (N_8224,N_5436,N_5228);
or U8225 (N_8225,N_4110,N_5162);
or U8226 (N_8226,N_4548,N_5969);
and U8227 (N_8227,N_5567,N_3933);
nor U8228 (N_8228,N_4224,N_3473);
nor U8229 (N_8229,N_5812,N_3701);
nor U8230 (N_8230,N_3669,N_5841);
or U8231 (N_8231,N_4196,N_3904);
nor U8232 (N_8232,N_4494,N_5442);
and U8233 (N_8233,N_5014,N_3730);
nor U8234 (N_8234,N_4485,N_5184);
and U8235 (N_8235,N_4238,N_3148);
and U8236 (N_8236,N_5279,N_3081);
nand U8237 (N_8237,N_4943,N_4558);
and U8238 (N_8238,N_4418,N_4660);
and U8239 (N_8239,N_4913,N_4461);
and U8240 (N_8240,N_5962,N_4603);
nor U8241 (N_8241,N_4420,N_3711);
nand U8242 (N_8242,N_4687,N_3412);
nor U8243 (N_8243,N_3243,N_5784);
nor U8244 (N_8244,N_5565,N_5104);
or U8245 (N_8245,N_4874,N_3230);
or U8246 (N_8246,N_3022,N_3617);
or U8247 (N_8247,N_5231,N_5995);
and U8248 (N_8248,N_5429,N_5696);
nor U8249 (N_8249,N_5005,N_3057);
and U8250 (N_8250,N_3288,N_5188);
nor U8251 (N_8251,N_5942,N_3933);
nand U8252 (N_8252,N_3289,N_3003);
nor U8253 (N_8253,N_3739,N_5981);
nor U8254 (N_8254,N_4747,N_5344);
and U8255 (N_8255,N_5064,N_3071);
or U8256 (N_8256,N_4728,N_3861);
or U8257 (N_8257,N_4677,N_4972);
nand U8258 (N_8258,N_3522,N_5839);
or U8259 (N_8259,N_3280,N_3583);
nor U8260 (N_8260,N_5420,N_4656);
and U8261 (N_8261,N_4293,N_5273);
or U8262 (N_8262,N_3047,N_4371);
nor U8263 (N_8263,N_4692,N_5508);
nor U8264 (N_8264,N_3279,N_3961);
nand U8265 (N_8265,N_5617,N_5916);
or U8266 (N_8266,N_3292,N_5144);
nor U8267 (N_8267,N_4025,N_5279);
and U8268 (N_8268,N_4519,N_4189);
or U8269 (N_8269,N_4278,N_3140);
nor U8270 (N_8270,N_3453,N_4050);
or U8271 (N_8271,N_5001,N_5200);
or U8272 (N_8272,N_3818,N_4870);
and U8273 (N_8273,N_5365,N_5320);
nand U8274 (N_8274,N_5027,N_3616);
nor U8275 (N_8275,N_5071,N_4886);
nand U8276 (N_8276,N_4624,N_3660);
nand U8277 (N_8277,N_5418,N_5107);
or U8278 (N_8278,N_4192,N_3745);
or U8279 (N_8279,N_5736,N_4032);
nand U8280 (N_8280,N_3440,N_5450);
and U8281 (N_8281,N_5882,N_3575);
or U8282 (N_8282,N_3986,N_4889);
nor U8283 (N_8283,N_5388,N_5718);
nor U8284 (N_8284,N_5713,N_3608);
nand U8285 (N_8285,N_4113,N_4063);
or U8286 (N_8286,N_5880,N_4129);
nor U8287 (N_8287,N_4542,N_5594);
nand U8288 (N_8288,N_3402,N_4681);
nor U8289 (N_8289,N_3822,N_3486);
and U8290 (N_8290,N_3021,N_3429);
or U8291 (N_8291,N_4708,N_4780);
nor U8292 (N_8292,N_4124,N_3610);
nand U8293 (N_8293,N_3108,N_4011);
or U8294 (N_8294,N_3597,N_4292);
and U8295 (N_8295,N_4943,N_3054);
nand U8296 (N_8296,N_5219,N_5081);
nand U8297 (N_8297,N_3506,N_3890);
nand U8298 (N_8298,N_3622,N_3749);
or U8299 (N_8299,N_4935,N_5895);
nand U8300 (N_8300,N_5992,N_4698);
nor U8301 (N_8301,N_4479,N_5730);
nand U8302 (N_8302,N_5779,N_5523);
or U8303 (N_8303,N_4011,N_3081);
and U8304 (N_8304,N_4710,N_5901);
nand U8305 (N_8305,N_5016,N_3120);
and U8306 (N_8306,N_4406,N_5969);
and U8307 (N_8307,N_4826,N_3592);
and U8308 (N_8308,N_5617,N_4374);
or U8309 (N_8309,N_3431,N_4706);
and U8310 (N_8310,N_5310,N_5159);
and U8311 (N_8311,N_5477,N_3712);
and U8312 (N_8312,N_5803,N_3794);
nor U8313 (N_8313,N_3325,N_5551);
nand U8314 (N_8314,N_5522,N_5832);
nand U8315 (N_8315,N_3400,N_5059);
nor U8316 (N_8316,N_4073,N_4618);
and U8317 (N_8317,N_3911,N_4141);
nand U8318 (N_8318,N_4922,N_3730);
and U8319 (N_8319,N_4082,N_5589);
or U8320 (N_8320,N_3794,N_4653);
nor U8321 (N_8321,N_4678,N_4256);
nor U8322 (N_8322,N_3310,N_4706);
or U8323 (N_8323,N_3809,N_5921);
nand U8324 (N_8324,N_4771,N_4783);
or U8325 (N_8325,N_4773,N_3172);
nor U8326 (N_8326,N_5701,N_4248);
nor U8327 (N_8327,N_5040,N_3569);
or U8328 (N_8328,N_5542,N_3661);
nor U8329 (N_8329,N_3909,N_5215);
nor U8330 (N_8330,N_3645,N_3746);
nor U8331 (N_8331,N_4330,N_3125);
nand U8332 (N_8332,N_5134,N_5462);
or U8333 (N_8333,N_3786,N_5968);
xnor U8334 (N_8334,N_3306,N_5518);
and U8335 (N_8335,N_3192,N_5729);
nand U8336 (N_8336,N_5202,N_4355);
nand U8337 (N_8337,N_4552,N_4614);
or U8338 (N_8338,N_3070,N_4405);
or U8339 (N_8339,N_4514,N_3060);
nor U8340 (N_8340,N_5008,N_3728);
and U8341 (N_8341,N_3393,N_3341);
or U8342 (N_8342,N_4456,N_5875);
nand U8343 (N_8343,N_3511,N_3386);
or U8344 (N_8344,N_3693,N_3592);
or U8345 (N_8345,N_4064,N_4908);
nor U8346 (N_8346,N_3547,N_4377);
nor U8347 (N_8347,N_4680,N_5851);
and U8348 (N_8348,N_5704,N_3224);
or U8349 (N_8349,N_3072,N_5516);
nand U8350 (N_8350,N_3851,N_4095);
and U8351 (N_8351,N_4228,N_4693);
nand U8352 (N_8352,N_3005,N_5249);
nor U8353 (N_8353,N_4468,N_5021);
nand U8354 (N_8354,N_3244,N_3521);
nand U8355 (N_8355,N_3029,N_4277);
or U8356 (N_8356,N_4443,N_3470);
and U8357 (N_8357,N_3519,N_3192);
or U8358 (N_8358,N_5960,N_4945);
and U8359 (N_8359,N_3779,N_4823);
or U8360 (N_8360,N_5422,N_4539);
or U8361 (N_8361,N_3347,N_4986);
and U8362 (N_8362,N_4837,N_5393);
or U8363 (N_8363,N_3582,N_4634);
and U8364 (N_8364,N_5343,N_5093);
and U8365 (N_8365,N_4389,N_4816);
xnor U8366 (N_8366,N_3423,N_4264);
or U8367 (N_8367,N_5712,N_3717);
and U8368 (N_8368,N_4585,N_5068);
nand U8369 (N_8369,N_3064,N_4259);
and U8370 (N_8370,N_4168,N_4567);
nand U8371 (N_8371,N_3141,N_5841);
or U8372 (N_8372,N_3491,N_4423);
and U8373 (N_8373,N_4990,N_3653);
nand U8374 (N_8374,N_4204,N_3931);
nor U8375 (N_8375,N_3525,N_3097);
nor U8376 (N_8376,N_3831,N_3577);
or U8377 (N_8377,N_5953,N_4564);
nand U8378 (N_8378,N_3934,N_3644);
nor U8379 (N_8379,N_3080,N_5853);
nor U8380 (N_8380,N_5225,N_5443);
or U8381 (N_8381,N_3269,N_4527);
xor U8382 (N_8382,N_4966,N_3195);
nor U8383 (N_8383,N_4465,N_4594);
and U8384 (N_8384,N_4825,N_3947);
nor U8385 (N_8385,N_4453,N_5986);
and U8386 (N_8386,N_3475,N_4752);
and U8387 (N_8387,N_4467,N_5728);
or U8388 (N_8388,N_3016,N_5916);
or U8389 (N_8389,N_5965,N_3064);
and U8390 (N_8390,N_3760,N_4546);
nand U8391 (N_8391,N_5409,N_4079);
or U8392 (N_8392,N_5319,N_3217);
and U8393 (N_8393,N_5778,N_3224);
nand U8394 (N_8394,N_3585,N_3270);
or U8395 (N_8395,N_5859,N_3510);
and U8396 (N_8396,N_3552,N_3672);
nand U8397 (N_8397,N_5789,N_3919);
and U8398 (N_8398,N_4617,N_5029);
and U8399 (N_8399,N_4212,N_5774);
nand U8400 (N_8400,N_5352,N_4226);
nand U8401 (N_8401,N_5060,N_3384);
or U8402 (N_8402,N_3850,N_5070);
or U8403 (N_8403,N_3321,N_3223);
and U8404 (N_8404,N_3843,N_4990);
nand U8405 (N_8405,N_4008,N_5216);
and U8406 (N_8406,N_3184,N_3818);
and U8407 (N_8407,N_3419,N_4748);
or U8408 (N_8408,N_3407,N_3682);
nand U8409 (N_8409,N_3656,N_3286);
nand U8410 (N_8410,N_5121,N_5158);
nor U8411 (N_8411,N_3482,N_3590);
nor U8412 (N_8412,N_4078,N_5960);
and U8413 (N_8413,N_3245,N_5381);
nor U8414 (N_8414,N_4494,N_5780);
or U8415 (N_8415,N_3593,N_5861);
and U8416 (N_8416,N_5479,N_4982);
nor U8417 (N_8417,N_5257,N_5476);
nor U8418 (N_8418,N_5801,N_4929);
nand U8419 (N_8419,N_3926,N_3404);
or U8420 (N_8420,N_5597,N_3678);
or U8421 (N_8421,N_3583,N_4663);
nor U8422 (N_8422,N_4239,N_3386);
nor U8423 (N_8423,N_3945,N_5562);
and U8424 (N_8424,N_3213,N_5395);
nand U8425 (N_8425,N_4271,N_4429);
and U8426 (N_8426,N_5375,N_3818);
nand U8427 (N_8427,N_3520,N_5850);
and U8428 (N_8428,N_4376,N_4451);
and U8429 (N_8429,N_5946,N_3265);
nand U8430 (N_8430,N_4711,N_4497);
or U8431 (N_8431,N_3559,N_4560);
nor U8432 (N_8432,N_4757,N_3910);
nor U8433 (N_8433,N_4433,N_4357);
and U8434 (N_8434,N_3825,N_3784);
and U8435 (N_8435,N_3284,N_4346);
and U8436 (N_8436,N_3283,N_5768);
nor U8437 (N_8437,N_5868,N_5969);
nor U8438 (N_8438,N_5019,N_5069);
and U8439 (N_8439,N_3101,N_3279);
and U8440 (N_8440,N_5540,N_4520);
or U8441 (N_8441,N_4831,N_5981);
or U8442 (N_8442,N_5852,N_3491);
nand U8443 (N_8443,N_4986,N_5913);
nand U8444 (N_8444,N_4751,N_5526);
or U8445 (N_8445,N_4224,N_3967);
and U8446 (N_8446,N_5363,N_5892);
nor U8447 (N_8447,N_4033,N_3368);
nand U8448 (N_8448,N_5490,N_4713);
nor U8449 (N_8449,N_5335,N_3561);
nor U8450 (N_8450,N_4948,N_4604);
nor U8451 (N_8451,N_4154,N_5452);
or U8452 (N_8452,N_4551,N_4366);
nor U8453 (N_8453,N_5871,N_4320);
nor U8454 (N_8454,N_5287,N_5676);
and U8455 (N_8455,N_5994,N_4928);
nand U8456 (N_8456,N_5666,N_5805);
nor U8457 (N_8457,N_3479,N_3205);
nor U8458 (N_8458,N_3968,N_3459);
nand U8459 (N_8459,N_5796,N_4751);
nand U8460 (N_8460,N_4222,N_5827);
nand U8461 (N_8461,N_5696,N_3149);
nor U8462 (N_8462,N_3176,N_4964);
nand U8463 (N_8463,N_4355,N_4795);
nand U8464 (N_8464,N_4260,N_4235);
and U8465 (N_8465,N_3225,N_3027);
and U8466 (N_8466,N_5220,N_3886);
nor U8467 (N_8467,N_5877,N_5804);
or U8468 (N_8468,N_5396,N_3768);
nor U8469 (N_8469,N_5655,N_4178);
nand U8470 (N_8470,N_3045,N_3736);
and U8471 (N_8471,N_5604,N_4248);
or U8472 (N_8472,N_5041,N_3057);
or U8473 (N_8473,N_3900,N_3475);
nor U8474 (N_8474,N_3218,N_4394);
nand U8475 (N_8475,N_4046,N_3641);
nand U8476 (N_8476,N_5232,N_4185);
nand U8477 (N_8477,N_4859,N_4812);
xnor U8478 (N_8478,N_4214,N_4618);
and U8479 (N_8479,N_4847,N_3254);
nand U8480 (N_8480,N_4966,N_5531);
nand U8481 (N_8481,N_5837,N_5669);
or U8482 (N_8482,N_4087,N_3449);
or U8483 (N_8483,N_5823,N_3858);
nand U8484 (N_8484,N_3586,N_3242);
or U8485 (N_8485,N_3894,N_3873);
nand U8486 (N_8486,N_3568,N_5840);
nand U8487 (N_8487,N_3620,N_4297);
and U8488 (N_8488,N_5472,N_4135);
or U8489 (N_8489,N_3861,N_3743);
or U8490 (N_8490,N_4413,N_3555);
and U8491 (N_8491,N_5021,N_4991);
nand U8492 (N_8492,N_5989,N_3261);
and U8493 (N_8493,N_5588,N_4672);
or U8494 (N_8494,N_3493,N_5345);
nand U8495 (N_8495,N_4507,N_4478);
nor U8496 (N_8496,N_3375,N_4133);
nor U8497 (N_8497,N_5216,N_3514);
nor U8498 (N_8498,N_5214,N_5047);
nor U8499 (N_8499,N_5561,N_4240);
and U8500 (N_8500,N_3090,N_5617);
nand U8501 (N_8501,N_5332,N_3515);
nand U8502 (N_8502,N_4761,N_3805);
nor U8503 (N_8503,N_3214,N_4438);
and U8504 (N_8504,N_5946,N_5028);
and U8505 (N_8505,N_4839,N_4528);
and U8506 (N_8506,N_3981,N_5017);
nand U8507 (N_8507,N_4207,N_4334);
nand U8508 (N_8508,N_3605,N_4722);
and U8509 (N_8509,N_4445,N_5168);
nor U8510 (N_8510,N_3295,N_3871);
nand U8511 (N_8511,N_3882,N_3372);
and U8512 (N_8512,N_5303,N_4853);
nand U8513 (N_8513,N_5175,N_5394);
or U8514 (N_8514,N_4618,N_4174);
and U8515 (N_8515,N_3329,N_4534);
or U8516 (N_8516,N_3465,N_5541);
or U8517 (N_8517,N_4634,N_5262);
nor U8518 (N_8518,N_4445,N_5486);
or U8519 (N_8519,N_4868,N_5296);
and U8520 (N_8520,N_3073,N_4634);
nand U8521 (N_8521,N_3833,N_4550);
nand U8522 (N_8522,N_5099,N_4681);
and U8523 (N_8523,N_3592,N_5661);
nor U8524 (N_8524,N_3909,N_5555);
nand U8525 (N_8525,N_3320,N_5985);
or U8526 (N_8526,N_5457,N_4220);
or U8527 (N_8527,N_5652,N_3396);
nand U8528 (N_8528,N_3885,N_3673);
or U8529 (N_8529,N_3149,N_5778);
and U8530 (N_8530,N_4425,N_4863);
and U8531 (N_8531,N_3467,N_4158);
nand U8532 (N_8532,N_3742,N_3728);
and U8533 (N_8533,N_4744,N_4027);
or U8534 (N_8534,N_5671,N_4092);
nor U8535 (N_8535,N_5553,N_3623);
nand U8536 (N_8536,N_5170,N_5405);
or U8537 (N_8537,N_3090,N_5855);
or U8538 (N_8538,N_4710,N_5404);
nor U8539 (N_8539,N_4403,N_4345);
nand U8540 (N_8540,N_4576,N_5928);
or U8541 (N_8541,N_3007,N_5257);
nand U8542 (N_8542,N_3462,N_4741);
and U8543 (N_8543,N_3667,N_5620);
nand U8544 (N_8544,N_3735,N_4078);
nor U8545 (N_8545,N_3197,N_4731);
and U8546 (N_8546,N_4147,N_5663);
nor U8547 (N_8547,N_4273,N_5450);
nand U8548 (N_8548,N_3338,N_4888);
nand U8549 (N_8549,N_5320,N_3493);
and U8550 (N_8550,N_4430,N_4069);
nand U8551 (N_8551,N_5421,N_5434);
and U8552 (N_8552,N_5087,N_4042);
nand U8553 (N_8553,N_5678,N_5661);
nand U8554 (N_8554,N_4397,N_3553);
or U8555 (N_8555,N_3508,N_3782);
or U8556 (N_8556,N_3444,N_5174);
or U8557 (N_8557,N_3355,N_4377);
nand U8558 (N_8558,N_4556,N_3677);
nor U8559 (N_8559,N_5856,N_5656);
nand U8560 (N_8560,N_4970,N_4265);
nor U8561 (N_8561,N_3657,N_3246);
nor U8562 (N_8562,N_3794,N_4706);
or U8563 (N_8563,N_3822,N_4959);
nor U8564 (N_8564,N_4659,N_4260);
and U8565 (N_8565,N_5039,N_3491);
nor U8566 (N_8566,N_5115,N_4198);
nand U8567 (N_8567,N_3103,N_5768);
or U8568 (N_8568,N_4801,N_3107);
and U8569 (N_8569,N_3153,N_5051);
nand U8570 (N_8570,N_3419,N_3077);
and U8571 (N_8571,N_3111,N_3199);
nor U8572 (N_8572,N_3666,N_4537);
and U8573 (N_8573,N_3424,N_5550);
or U8574 (N_8574,N_4370,N_4264);
nor U8575 (N_8575,N_5721,N_4756);
nand U8576 (N_8576,N_4067,N_5918);
and U8577 (N_8577,N_3630,N_4407);
nand U8578 (N_8578,N_5805,N_5698);
nor U8579 (N_8579,N_3130,N_5083);
nor U8580 (N_8580,N_3577,N_5186);
nand U8581 (N_8581,N_5061,N_3961);
and U8582 (N_8582,N_3108,N_5090);
xor U8583 (N_8583,N_3882,N_5790);
and U8584 (N_8584,N_5145,N_4080);
or U8585 (N_8585,N_5960,N_3555);
or U8586 (N_8586,N_5811,N_4520);
nand U8587 (N_8587,N_4728,N_4811);
xnor U8588 (N_8588,N_3690,N_3940);
and U8589 (N_8589,N_3425,N_3059);
nor U8590 (N_8590,N_4398,N_4921);
nand U8591 (N_8591,N_5787,N_3203);
nor U8592 (N_8592,N_3762,N_4169);
nor U8593 (N_8593,N_3896,N_5223);
nand U8594 (N_8594,N_5845,N_4215);
nor U8595 (N_8595,N_4817,N_3894);
and U8596 (N_8596,N_4415,N_5486);
or U8597 (N_8597,N_3116,N_4690);
and U8598 (N_8598,N_5995,N_3411);
nand U8599 (N_8599,N_3635,N_4898);
nor U8600 (N_8600,N_3502,N_4804);
nor U8601 (N_8601,N_5600,N_3979);
nand U8602 (N_8602,N_3731,N_5084);
nand U8603 (N_8603,N_3076,N_4003);
nor U8604 (N_8604,N_3062,N_4507);
nand U8605 (N_8605,N_4253,N_5364);
nand U8606 (N_8606,N_3095,N_4959);
or U8607 (N_8607,N_3501,N_4595);
or U8608 (N_8608,N_5447,N_4367);
or U8609 (N_8609,N_4900,N_4680);
nor U8610 (N_8610,N_4788,N_4640);
or U8611 (N_8611,N_5269,N_4552);
or U8612 (N_8612,N_5076,N_4552);
nand U8613 (N_8613,N_3096,N_5336);
and U8614 (N_8614,N_3868,N_5693);
nor U8615 (N_8615,N_4145,N_4108);
nor U8616 (N_8616,N_3516,N_5633);
nor U8617 (N_8617,N_4111,N_4422);
and U8618 (N_8618,N_4198,N_4813);
or U8619 (N_8619,N_4187,N_4770);
nand U8620 (N_8620,N_5290,N_3863);
or U8621 (N_8621,N_3759,N_3062);
nand U8622 (N_8622,N_5561,N_4990);
and U8623 (N_8623,N_5924,N_3710);
xor U8624 (N_8624,N_5134,N_3822);
nor U8625 (N_8625,N_4659,N_4086);
nand U8626 (N_8626,N_5859,N_3479);
nor U8627 (N_8627,N_4379,N_4545);
nor U8628 (N_8628,N_3631,N_4345);
nor U8629 (N_8629,N_4790,N_5449);
or U8630 (N_8630,N_4851,N_4718);
nand U8631 (N_8631,N_3507,N_3308);
nor U8632 (N_8632,N_5394,N_4621);
or U8633 (N_8633,N_3230,N_5474);
nand U8634 (N_8634,N_4641,N_5045);
nor U8635 (N_8635,N_3022,N_3435);
or U8636 (N_8636,N_3642,N_4762);
nand U8637 (N_8637,N_3580,N_5336);
and U8638 (N_8638,N_4029,N_4456);
nand U8639 (N_8639,N_4182,N_5436);
nand U8640 (N_8640,N_5987,N_4607);
nor U8641 (N_8641,N_3150,N_5083);
or U8642 (N_8642,N_3370,N_4012);
and U8643 (N_8643,N_3496,N_5869);
or U8644 (N_8644,N_5638,N_5076);
or U8645 (N_8645,N_5298,N_4323);
nor U8646 (N_8646,N_5672,N_4703);
and U8647 (N_8647,N_5958,N_3546);
nor U8648 (N_8648,N_3574,N_5371);
or U8649 (N_8649,N_5730,N_3224);
nand U8650 (N_8650,N_4171,N_3316);
nor U8651 (N_8651,N_3619,N_3893);
and U8652 (N_8652,N_5791,N_4841);
and U8653 (N_8653,N_3174,N_3688);
nand U8654 (N_8654,N_3396,N_4077);
nor U8655 (N_8655,N_3300,N_3731);
or U8656 (N_8656,N_3811,N_4244);
nand U8657 (N_8657,N_4844,N_4360);
and U8658 (N_8658,N_5539,N_5191);
and U8659 (N_8659,N_5721,N_3157);
nor U8660 (N_8660,N_5744,N_5754);
nand U8661 (N_8661,N_3841,N_3307);
or U8662 (N_8662,N_4323,N_4047);
or U8663 (N_8663,N_5286,N_3249);
and U8664 (N_8664,N_5928,N_3513);
or U8665 (N_8665,N_5219,N_3820);
or U8666 (N_8666,N_4587,N_3467);
nand U8667 (N_8667,N_4500,N_5566);
or U8668 (N_8668,N_5158,N_4814);
and U8669 (N_8669,N_5441,N_5920);
and U8670 (N_8670,N_3634,N_5944);
or U8671 (N_8671,N_5625,N_4175);
and U8672 (N_8672,N_5637,N_3756);
nor U8673 (N_8673,N_3039,N_5904);
nand U8674 (N_8674,N_3938,N_4365);
and U8675 (N_8675,N_4405,N_4134);
and U8676 (N_8676,N_5972,N_3504);
and U8677 (N_8677,N_5522,N_5282);
or U8678 (N_8678,N_4932,N_3294);
nand U8679 (N_8679,N_5658,N_3991);
or U8680 (N_8680,N_3716,N_4847);
nor U8681 (N_8681,N_4465,N_4928);
nor U8682 (N_8682,N_5520,N_5881);
and U8683 (N_8683,N_3094,N_4668);
and U8684 (N_8684,N_5283,N_5512);
nor U8685 (N_8685,N_4004,N_4488);
nor U8686 (N_8686,N_3551,N_4595);
or U8687 (N_8687,N_4752,N_4413);
or U8688 (N_8688,N_4336,N_3447);
nand U8689 (N_8689,N_5383,N_3333);
nor U8690 (N_8690,N_5611,N_4017);
and U8691 (N_8691,N_4824,N_4767);
and U8692 (N_8692,N_5444,N_4719);
and U8693 (N_8693,N_3857,N_3092);
and U8694 (N_8694,N_3462,N_5792);
nand U8695 (N_8695,N_4120,N_4782);
nor U8696 (N_8696,N_5985,N_3829);
nand U8697 (N_8697,N_5828,N_4803);
and U8698 (N_8698,N_3656,N_4965);
nand U8699 (N_8699,N_3698,N_4029);
nand U8700 (N_8700,N_5937,N_3558);
or U8701 (N_8701,N_3754,N_5741);
or U8702 (N_8702,N_3685,N_3267);
nor U8703 (N_8703,N_5917,N_5398);
nand U8704 (N_8704,N_5634,N_4026);
or U8705 (N_8705,N_4930,N_4011);
nand U8706 (N_8706,N_4387,N_3201);
and U8707 (N_8707,N_5531,N_4438);
nand U8708 (N_8708,N_5425,N_5559);
or U8709 (N_8709,N_3510,N_4641);
and U8710 (N_8710,N_4077,N_3213);
nand U8711 (N_8711,N_5429,N_4340);
or U8712 (N_8712,N_5324,N_5729);
or U8713 (N_8713,N_5377,N_3646);
and U8714 (N_8714,N_4990,N_4006);
nor U8715 (N_8715,N_4742,N_4821);
and U8716 (N_8716,N_4130,N_3107);
nand U8717 (N_8717,N_4295,N_3926);
or U8718 (N_8718,N_3677,N_4082);
and U8719 (N_8719,N_5510,N_4840);
nand U8720 (N_8720,N_4708,N_4520);
nor U8721 (N_8721,N_5058,N_4997);
nor U8722 (N_8722,N_5195,N_5002);
and U8723 (N_8723,N_3441,N_5937);
and U8724 (N_8724,N_3469,N_5036);
nand U8725 (N_8725,N_5598,N_3368);
nor U8726 (N_8726,N_4760,N_4069);
nor U8727 (N_8727,N_5080,N_3145);
nand U8728 (N_8728,N_4737,N_4542);
or U8729 (N_8729,N_5941,N_5796);
nor U8730 (N_8730,N_3264,N_3742);
nand U8731 (N_8731,N_5778,N_3060);
or U8732 (N_8732,N_3257,N_4782);
nor U8733 (N_8733,N_5467,N_3924);
and U8734 (N_8734,N_5012,N_3588);
nand U8735 (N_8735,N_4815,N_3000);
nand U8736 (N_8736,N_4416,N_5971);
or U8737 (N_8737,N_3078,N_4989);
and U8738 (N_8738,N_5034,N_4264);
or U8739 (N_8739,N_3077,N_4494);
or U8740 (N_8740,N_3594,N_3144);
or U8741 (N_8741,N_4707,N_4936);
or U8742 (N_8742,N_4918,N_4690);
nor U8743 (N_8743,N_5413,N_5016);
and U8744 (N_8744,N_4504,N_5652);
or U8745 (N_8745,N_5659,N_4632);
nand U8746 (N_8746,N_5478,N_3426);
or U8747 (N_8747,N_5426,N_3632);
nand U8748 (N_8748,N_4609,N_4970);
nor U8749 (N_8749,N_3023,N_3557);
nor U8750 (N_8750,N_4074,N_4305);
or U8751 (N_8751,N_4859,N_5441);
or U8752 (N_8752,N_5995,N_3913);
nor U8753 (N_8753,N_5943,N_5180);
nand U8754 (N_8754,N_5982,N_5763);
or U8755 (N_8755,N_4196,N_4795);
nand U8756 (N_8756,N_3203,N_3722);
nand U8757 (N_8757,N_3674,N_4601);
nor U8758 (N_8758,N_5732,N_4334);
or U8759 (N_8759,N_5869,N_3930);
nor U8760 (N_8760,N_5404,N_3376);
nor U8761 (N_8761,N_3266,N_3140);
or U8762 (N_8762,N_3559,N_5283);
and U8763 (N_8763,N_5039,N_3946);
nand U8764 (N_8764,N_3224,N_3954);
nor U8765 (N_8765,N_3268,N_4574);
nor U8766 (N_8766,N_3571,N_3384);
nand U8767 (N_8767,N_5799,N_5581);
or U8768 (N_8768,N_3395,N_3091);
or U8769 (N_8769,N_5839,N_3055);
nor U8770 (N_8770,N_4943,N_4116);
nor U8771 (N_8771,N_5510,N_4967);
nand U8772 (N_8772,N_5139,N_4952);
nor U8773 (N_8773,N_3496,N_5037);
and U8774 (N_8774,N_4790,N_5383);
nand U8775 (N_8775,N_5772,N_3393);
nor U8776 (N_8776,N_5356,N_3397);
nor U8777 (N_8777,N_3769,N_5955);
nor U8778 (N_8778,N_3787,N_5809);
xnor U8779 (N_8779,N_5432,N_3421);
and U8780 (N_8780,N_3625,N_4471);
nor U8781 (N_8781,N_5630,N_5599);
nand U8782 (N_8782,N_4497,N_3016);
or U8783 (N_8783,N_5928,N_3636);
nand U8784 (N_8784,N_4365,N_4473);
or U8785 (N_8785,N_4446,N_3580);
nor U8786 (N_8786,N_4148,N_3031);
or U8787 (N_8787,N_4917,N_5136);
nand U8788 (N_8788,N_4244,N_4970);
nor U8789 (N_8789,N_3779,N_3234);
and U8790 (N_8790,N_3344,N_5508);
nand U8791 (N_8791,N_3893,N_4878);
nand U8792 (N_8792,N_3286,N_5830);
nand U8793 (N_8793,N_3132,N_4277);
or U8794 (N_8794,N_3172,N_3300);
nand U8795 (N_8795,N_4058,N_3144);
or U8796 (N_8796,N_3537,N_3295);
or U8797 (N_8797,N_3150,N_4091);
or U8798 (N_8798,N_4876,N_3757);
nor U8799 (N_8799,N_3890,N_5830);
nand U8800 (N_8800,N_5001,N_4783);
nand U8801 (N_8801,N_5588,N_4731);
nor U8802 (N_8802,N_4078,N_3610);
or U8803 (N_8803,N_5744,N_5822);
or U8804 (N_8804,N_5211,N_4101);
or U8805 (N_8805,N_5749,N_4664);
and U8806 (N_8806,N_3604,N_5441);
nor U8807 (N_8807,N_3283,N_4049);
or U8808 (N_8808,N_5701,N_5361);
nor U8809 (N_8809,N_5951,N_4370);
or U8810 (N_8810,N_4921,N_5467);
or U8811 (N_8811,N_4345,N_5100);
or U8812 (N_8812,N_5844,N_3385);
and U8813 (N_8813,N_3873,N_5348);
nor U8814 (N_8814,N_3898,N_3341);
nor U8815 (N_8815,N_3854,N_3700);
and U8816 (N_8816,N_5573,N_3373);
nor U8817 (N_8817,N_5829,N_5094);
xnor U8818 (N_8818,N_4517,N_3278);
nor U8819 (N_8819,N_5328,N_4640);
or U8820 (N_8820,N_5256,N_3968);
nor U8821 (N_8821,N_3698,N_4961);
or U8822 (N_8822,N_4201,N_3055);
or U8823 (N_8823,N_3640,N_3776);
or U8824 (N_8824,N_4274,N_5180);
nand U8825 (N_8825,N_4275,N_3004);
nor U8826 (N_8826,N_4935,N_3270);
nor U8827 (N_8827,N_3665,N_4842);
xnor U8828 (N_8828,N_3988,N_4933);
or U8829 (N_8829,N_5932,N_5266);
nand U8830 (N_8830,N_5742,N_4842);
nand U8831 (N_8831,N_3050,N_5238);
or U8832 (N_8832,N_5921,N_3570);
or U8833 (N_8833,N_5062,N_5110);
nand U8834 (N_8834,N_5819,N_3805);
or U8835 (N_8835,N_5382,N_3354);
nand U8836 (N_8836,N_4499,N_3272);
and U8837 (N_8837,N_4592,N_4156);
nor U8838 (N_8838,N_5434,N_4128);
or U8839 (N_8839,N_3982,N_3679);
nor U8840 (N_8840,N_5617,N_3681);
nand U8841 (N_8841,N_4812,N_3294);
and U8842 (N_8842,N_4006,N_3036);
or U8843 (N_8843,N_5645,N_4287);
nor U8844 (N_8844,N_4150,N_4590);
or U8845 (N_8845,N_3446,N_4460);
and U8846 (N_8846,N_3661,N_5434);
and U8847 (N_8847,N_4899,N_4006);
and U8848 (N_8848,N_3408,N_3881);
nor U8849 (N_8849,N_4046,N_4938);
or U8850 (N_8850,N_5175,N_3117);
or U8851 (N_8851,N_5603,N_5610);
nand U8852 (N_8852,N_3741,N_4235);
or U8853 (N_8853,N_5331,N_4213);
and U8854 (N_8854,N_4867,N_5429);
or U8855 (N_8855,N_4906,N_3405);
nand U8856 (N_8856,N_5842,N_4330);
nand U8857 (N_8857,N_3206,N_4087);
and U8858 (N_8858,N_4924,N_4318);
nor U8859 (N_8859,N_3075,N_5188);
and U8860 (N_8860,N_4380,N_4866);
or U8861 (N_8861,N_4557,N_4388);
or U8862 (N_8862,N_3198,N_4796);
and U8863 (N_8863,N_4431,N_3115);
xor U8864 (N_8864,N_4686,N_3775);
nor U8865 (N_8865,N_5205,N_3214);
nor U8866 (N_8866,N_3204,N_4667);
or U8867 (N_8867,N_4714,N_5443);
or U8868 (N_8868,N_3684,N_3093);
and U8869 (N_8869,N_5280,N_4562);
or U8870 (N_8870,N_5488,N_5437);
nor U8871 (N_8871,N_5586,N_4523);
and U8872 (N_8872,N_4117,N_5989);
nand U8873 (N_8873,N_3816,N_5657);
nand U8874 (N_8874,N_4180,N_3340);
and U8875 (N_8875,N_5600,N_3629);
or U8876 (N_8876,N_4929,N_3649);
and U8877 (N_8877,N_4779,N_3260);
or U8878 (N_8878,N_5726,N_4606);
nand U8879 (N_8879,N_4292,N_5511);
and U8880 (N_8880,N_3130,N_3881);
nand U8881 (N_8881,N_3244,N_3501);
and U8882 (N_8882,N_4866,N_5967);
or U8883 (N_8883,N_4819,N_4013);
and U8884 (N_8884,N_4213,N_5801);
xor U8885 (N_8885,N_3302,N_3931);
nand U8886 (N_8886,N_5257,N_3170);
nor U8887 (N_8887,N_3974,N_3674);
nand U8888 (N_8888,N_4476,N_5580);
nor U8889 (N_8889,N_5123,N_4105);
and U8890 (N_8890,N_4562,N_5475);
or U8891 (N_8891,N_5650,N_3746);
or U8892 (N_8892,N_3664,N_5494);
nand U8893 (N_8893,N_3715,N_3025);
nand U8894 (N_8894,N_5771,N_5609);
nand U8895 (N_8895,N_5931,N_3317);
nand U8896 (N_8896,N_5341,N_3964);
nor U8897 (N_8897,N_5715,N_5674);
and U8898 (N_8898,N_5608,N_4937);
nor U8899 (N_8899,N_5931,N_5958);
nand U8900 (N_8900,N_3754,N_5120);
nand U8901 (N_8901,N_3909,N_4257);
and U8902 (N_8902,N_5890,N_5747);
nor U8903 (N_8903,N_3104,N_4212);
nand U8904 (N_8904,N_3484,N_4383);
nor U8905 (N_8905,N_4696,N_4479);
and U8906 (N_8906,N_4085,N_3540);
nor U8907 (N_8907,N_4055,N_4313);
nor U8908 (N_8908,N_4387,N_5098);
nand U8909 (N_8909,N_4907,N_4882);
or U8910 (N_8910,N_3913,N_4743);
or U8911 (N_8911,N_3348,N_4458);
nor U8912 (N_8912,N_3889,N_4262);
or U8913 (N_8913,N_3057,N_3707);
nor U8914 (N_8914,N_3399,N_3925);
nor U8915 (N_8915,N_3477,N_5911);
nor U8916 (N_8916,N_4806,N_4654);
nand U8917 (N_8917,N_4549,N_3537);
or U8918 (N_8918,N_3540,N_5659);
and U8919 (N_8919,N_5794,N_5503);
or U8920 (N_8920,N_5113,N_3949);
nand U8921 (N_8921,N_4875,N_4487);
nor U8922 (N_8922,N_3095,N_3039);
nor U8923 (N_8923,N_4168,N_4105);
nor U8924 (N_8924,N_5149,N_5667);
and U8925 (N_8925,N_4425,N_4959);
nand U8926 (N_8926,N_4559,N_5229);
nor U8927 (N_8927,N_5124,N_3125);
and U8928 (N_8928,N_3261,N_5920);
nor U8929 (N_8929,N_3673,N_5400);
or U8930 (N_8930,N_4795,N_3500);
or U8931 (N_8931,N_4745,N_4845);
or U8932 (N_8932,N_3807,N_3546);
nor U8933 (N_8933,N_5391,N_5014);
nor U8934 (N_8934,N_4730,N_3573);
nor U8935 (N_8935,N_4931,N_3967);
and U8936 (N_8936,N_4492,N_5446);
nor U8937 (N_8937,N_4363,N_4847);
or U8938 (N_8938,N_3623,N_4141);
and U8939 (N_8939,N_4215,N_3560);
and U8940 (N_8940,N_3117,N_3869);
or U8941 (N_8941,N_5365,N_4417);
or U8942 (N_8942,N_4956,N_5896);
or U8943 (N_8943,N_5809,N_4225);
and U8944 (N_8944,N_5501,N_5178);
nand U8945 (N_8945,N_5997,N_5055);
and U8946 (N_8946,N_5686,N_5930);
nand U8947 (N_8947,N_3866,N_5417);
xnor U8948 (N_8948,N_3102,N_5675);
nand U8949 (N_8949,N_4278,N_4329);
and U8950 (N_8950,N_4599,N_5880);
and U8951 (N_8951,N_4165,N_5719);
nor U8952 (N_8952,N_4709,N_3249);
and U8953 (N_8953,N_3304,N_5065);
nor U8954 (N_8954,N_4699,N_4888);
and U8955 (N_8955,N_5685,N_3057);
and U8956 (N_8956,N_4468,N_5711);
nor U8957 (N_8957,N_4590,N_5362);
nand U8958 (N_8958,N_3735,N_3494);
or U8959 (N_8959,N_5211,N_4985);
nor U8960 (N_8960,N_3896,N_5761);
nor U8961 (N_8961,N_4770,N_5671);
nor U8962 (N_8962,N_3202,N_5638);
and U8963 (N_8963,N_3258,N_3410);
and U8964 (N_8964,N_5433,N_4392);
and U8965 (N_8965,N_5499,N_5461);
nand U8966 (N_8966,N_4792,N_5239);
nor U8967 (N_8967,N_3331,N_4523);
nand U8968 (N_8968,N_5823,N_3152);
nand U8969 (N_8969,N_5907,N_4087);
and U8970 (N_8970,N_3669,N_5318);
nand U8971 (N_8971,N_4850,N_5586);
nor U8972 (N_8972,N_5876,N_3977);
and U8973 (N_8973,N_4768,N_3627);
and U8974 (N_8974,N_4041,N_3248);
nor U8975 (N_8975,N_3717,N_4532);
and U8976 (N_8976,N_3979,N_5441);
nor U8977 (N_8977,N_4260,N_5743);
and U8978 (N_8978,N_3545,N_5854);
nor U8979 (N_8979,N_4755,N_4233);
nand U8980 (N_8980,N_3029,N_3738);
nor U8981 (N_8981,N_3643,N_3181);
and U8982 (N_8982,N_4712,N_5843);
and U8983 (N_8983,N_3315,N_5346);
nand U8984 (N_8984,N_5588,N_3367);
and U8985 (N_8985,N_3986,N_5061);
or U8986 (N_8986,N_5233,N_5792);
nand U8987 (N_8987,N_4403,N_4153);
nor U8988 (N_8988,N_5636,N_3750);
and U8989 (N_8989,N_3191,N_5724);
or U8990 (N_8990,N_3892,N_3143);
nand U8991 (N_8991,N_3532,N_3873);
nand U8992 (N_8992,N_3977,N_4716);
and U8993 (N_8993,N_5779,N_5087);
and U8994 (N_8994,N_4800,N_5694);
nor U8995 (N_8995,N_5059,N_5353);
and U8996 (N_8996,N_5157,N_4567);
and U8997 (N_8997,N_3956,N_5603);
nor U8998 (N_8998,N_3348,N_5807);
nand U8999 (N_8999,N_4925,N_5447);
nor U9000 (N_9000,N_7702,N_7205);
and U9001 (N_9001,N_8834,N_7429);
or U9002 (N_9002,N_7575,N_6524);
nor U9003 (N_9003,N_7379,N_8388);
nor U9004 (N_9004,N_8888,N_6233);
and U9005 (N_9005,N_6422,N_6353);
nor U9006 (N_9006,N_6779,N_7123);
or U9007 (N_9007,N_8634,N_8345);
nor U9008 (N_9008,N_8746,N_8279);
nor U9009 (N_9009,N_7440,N_8587);
nand U9010 (N_9010,N_8170,N_6606);
nand U9011 (N_9011,N_6411,N_7744);
nor U9012 (N_9012,N_8195,N_6658);
nor U9013 (N_9013,N_8353,N_7571);
or U9014 (N_9014,N_6224,N_7244);
xor U9015 (N_9015,N_8306,N_6197);
nand U9016 (N_9016,N_7452,N_7489);
and U9017 (N_9017,N_8946,N_6941);
or U9018 (N_9018,N_7284,N_8928);
nor U9019 (N_9019,N_6786,N_7255);
and U9020 (N_9020,N_6818,N_6426);
and U9021 (N_9021,N_6871,N_7032);
nor U9022 (N_9022,N_6169,N_7209);
and U9023 (N_9023,N_7014,N_8258);
or U9024 (N_9024,N_7406,N_7331);
and U9025 (N_9025,N_8537,N_8357);
nand U9026 (N_9026,N_6063,N_6024);
and U9027 (N_9027,N_6351,N_6093);
nand U9028 (N_9028,N_7795,N_6053);
nor U9029 (N_9029,N_7319,N_8288);
or U9030 (N_9030,N_6827,N_8425);
nor U9031 (N_9031,N_8990,N_8988);
nand U9032 (N_9032,N_7347,N_7404);
and U9033 (N_9033,N_6472,N_6129);
and U9034 (N_9034,N_6593,N_6320);
or U9035 (N_9035,N_7986,N_8086);
nand U9036 (N_9036,N_8497,N_6223);
nand U9037 (N_9037,N_8320,N_8368);
or U9038 (N_9038,N_8160,N_7106);
nand U9039 (N_9039,N_7105,N_8082);
or U9040 (N_9040,N_8821,N_6898);
and U9041 (N_9041,N_8630,N_6925);
or U9042 (N_9042,N_8885,N_6916);
nand U9043 (N_9043,N_7859,N_7761);
or U9044 (N_9044,N_6300,N_6058);
and U9045 (N_9045,N_8807,N_7860);
nand U9046 (N_9046,N_6112,N_8073);
or U9047 (N_9047,N_7625,N_8131);
nand U9048 (N_9048,N_7771,N_7349);
or U9049 (N_9049,N_8934,N_7982);
nor U9050 (N_9050,N_6635,N_7926);
nor U9051 (N_9051,N_6948,N_6376);
xor U9052 (N_9052,N_7763,N_6346);
and U9053 (N_9053,N_7350,N_8054);
nor U9054 (N_9054,N_6480,N_7346);
nor U9055 (N_9055,N_6153,N_7536);
or U9056 (N_9056,N_8406,N_8595);
nor U9057 (N_9057,N_8047,N_7131);
or U9058 (N_9058,N_7647,N_8509);
nand U9059 (N_9059,N_6111,N_7493);
and U9060 (N_9060,N_8840,N_7089);
and U9061 (N_9061,N_8230,N_6036);
nor U9062 (N_9062,N_7765,N_6288);
nor U9063 (N_9063,N_7740,N_6164);
nand U9064 (N_9064,N_7392,N_8499);
nand U9065 (N_9065,N_8691,N_7138);
nor U9066 (N_9066,N_8111,N_6578);
and U9067 (N_9067,N_7259,N_7360);
or U9068 (N_9068,N_6421,N_7001);
nor U9069 (N_9069,N_7964,N_7760);
nor U9070 (N_9070,N_6445,N_7621);
and U9071 (N_9071,N_6231,N_8447);
and U9072 (N_9072,N_7983,N_6767);
or U9073 (N_9073,N_8496,N_6051);
nand U9074 (N_9074,N_8226,N_6553);
nor U9075 (N_9075,N_7203,N_6564);
or U9076 (N_9076,N_8590,N_6208);
and U9077 (N_9077,N_8552,N_7516);
and U9078 (N_9078,N_6056,N_6436);
and U9079 (N_9079,N_6872,N_8680);
nor U9080 (N_9080,N_7335,N_7509);
and U9081 (N_9081,N_6294,N_7037);
nor U9082 (N_9082,N_8655,N_6530);
and U9083 (N_9083,N_6584,N_7042);
and U9084 (N_9084,N_6444,N_6694);
nand U9085 (N_9085,N_6017,N_8322);
or U9086 (N_9086,N_6810,N_7401);
and U9087 (N_9087,N_7325,N_6859);
or U9088 (N_9088,N_7507,N_8905);
and U9089 (N_9089,N_7112,N_7181);
nor U9090 (N_9090,N_6020,N_6567);
nand U9091 (N_9091,N_8823,N_6640);
and U9092 (N_9092,N_6760,N_7180);
nand U9093 (N_9093,N_8392,N_7544);
or U9094 (N_9094,N_7371,N_7249);
nor U9095 (N_9095,N_7035,N_6711);
or U9096 (N_9096,N_6725,N_7864);
nand U9097 (N_9097,N_8294,N_7616);
nand U9098 (N_9098,N_8531,N_8972);
and U9099 (N_9099,N_8025,N_7425);
nor U9100 (N_9100,N_8610,N_6212);
nor U9101 (N_9101,N_6579,N_7899);
nor U9102 (N_9102,N_7879,N_7052);
and U9103 (N_9103,N_8040,N_6296);
nand U9104 (N_9104,N_8663,N_8962);
or U9105 (N_9105,N_6149,N_8613);
or U9106 (N_9106,N_7091,N_8204);
nor U9107 (N_9107,N_8700,N_6004);
or U9108 (N_9108,N_8185,N_6176);
or U9109 (N_9109,N_6536,N_7756);
nor U9110 (N_9110,N_6778,N_7020);
and U9111 (N_9111,N_6964,N_8423);
and U9112 (N_9112,N_7132,N_8601);
xnor U9113 (N_9113,N_6309,N_7329);
nor U9114 (N_9114,N_8546,N_7301);
or U9115 (N_9115,N_7681,N_7364);
and U9116 (N_9116,N_6631,N_7258);
nand U9117 (N_9117,N_6045,N_6371);
nor U9118 (N_9118,N_6209,N_6693);
or U9119 (N_9119,N_6367,N_7537);
or U9120 (N_9120,N_6338,N_8362);
nor U9121 (N_9121,N_8057,N_6868);
or U9122 (N_9122,N_7519,N_6756);
nor U9123 (N_9123,N_8354,N_6406);
and U9124 (N_9124,N_8352,N_7597);
or U9125 (N_9125,N_6213,N_7328);
nor U9126 (N_9126,N_7520,N_8830);
nand U9127 (N_9127,N_6393,N_7423);
nor U9128 (N_9128,N_6886,N_7158);
or U9129 (N_9129,N_6404,N_7311);
or U9130 (N_9130,N_7247,N_6830);
or U9131 (N_9131,N_6229,N_8019);
or U9132 (N_9132,N_7114,N_6260);
or U9133 (N_9133,N_7805,N_8666);
and U9134 (N_9134,N_8557,N_7380);
and U9135 (N_9135,N_6379,N_8660);
and U9136 (N_9136,N_6959,N_8402);
nand U9137 (N_9137,N_8163,N_8287);
nand U9138 (N_9138,N_8745,N_6982);
nor U9139 (N_9139,N_6425,N_8408);
and U9140 (N_9140,N_7831,N_7093);
and U9141 (N_9141,N_8200,N_8790);
or U9142 (N_9142,N_6005,N_7248);
nand U9143 (N_9143,N_6442,N_8524);
and U9144 (N_9144,N_7028,N_7774);
and U9145 (N_9145,N_8451,N_6549);
nand U9146 (N_9146,N_8097,N_6597);
nand U9147 (N_9147,N_7736,N_8028);
nand U9148 (N_9148,N_7821,N_7517);
nor U9149 (N_9149,N_8310,N_8029);
nand U9150 (N_9150,N_7000,N_6280);
or U9151 (N_9151,N_6855,N_8330);
and U9152 (N_9152,N_8887,N_7826);
or U9153 (N_9153,N_6754,N_8624);
or U9154 (N_9154,N_7835,N_7602);
or U9155 (N_9155,N_8867,N_7278);
nand U9156 (N_9156,N_7746,N_6595);
or U9157 (N_9157,N_7709,N_8898);
or U9158 (N_9158,N_6980,N_8532);
or U9159 (N_9159,N_8386,N_6021);
or U9160 (N_9160,N_8658,N_6569);
or U9161 (N_9161,N_6732,N_6849);
nor U9162 (N_9162,N_7629,N_6313);
or U9163 (N_9163,N_8023,N_6576);
and U9164 (N_9164,N_7593,N_6254);
nor U9165 (N_9165,N_7355,N_8014);
and U9166 (N_9166,N_7776,N_7530);
nor U9167 (N_9167,N_7045,N_6744);
nand U9168 (N_9168,N_6327,N_6455);
and U9169 (N_9169,N_8038,N_7121);
or U9170 (N_9170,N_7660,N_7356);
and U9171 (N_9171,N_8882,N_7690);
nor U9172 (N_9172,N_8827,N_7897);
nor U9173 (N_9173,N_7006,N_6440);
or U9174 (N_9174,N_8498,N_7149);
or U9175 (N_9175,N_7584,N_6001);
nor U9176 (N_9176,N_7451,N_6811);
or U9177 (N_9177,N_6594,N_7395);
nand U9178 (N_9178,N_6883,N_6081);
nand U9179 (N_9179,N_8804,N_7747);
nor U9180 (N_9180,N_8802,N_6022);
nand U9181 (N_9181,N_7172,N_8342);
or U9182 (N_9182,N_7876,N_6906);
nor U9183 (N_9183,N_6347,N_6032);
and U9184 (N_9184,N_7476,N_7657);
nand U9185 (N_9185,N_8329,N_8224);
nor U9186 (N_9186,N_8366,N_8635);
nand U9187 (N_9187,N_8578,N_6620);
and U9188 (N_9188,N_6207,N_6145);
nand U9189 (N_9189,N_8449,N_7454);
nor U9190 (N_9190,N_8314,N_8800);
and U9191 (N_9191,N_6873,N_8120);
nor U9192 (N_9192,N_8332,N_6281);
and U9193 (N_9193,N_6533,N_7898);
or U9194 (N_9194,N_7612,N_8187);
nor U9195 (N_9195,N_7310,N_7990);
nor U9196 (N_9196,N_7388,N_6104);
nand U9197 (N_9197,N_6630,N_7659);
nand U9198 (N_9198,N_8511,N_7743);
nor U9199 (N_9199,N_8782,N_7783);
nand U9200 (N_9200,N_7521,N_7296);
nand U9201 (N_9201,N_7101,N_8237);
nand U9202 (N_9202,N_6844,N_6014);
nand U9203 (N_9203,N_8442,N_6375);
nand U9204 (N_9204,N_8290,N_6326);
nor U9205 (N_9205,N_8466,N_7762);
and U9206 (N_9206,N_6088,N_7884);
nand U9207 (N_9207,N_8156,N_7506);
nor U9208 (N_9208,N_8521,N_7769);
nor U9209 (N_9209,N_8334,N_7855);
and U9210 (N_9210,N_6646,N_7485);
nand U9211 (N_9211,N_8923,N_7154);
nor U9212 (N_9212,N_8883,N_8145);
and U9213 (N_9213,N_7268,N_6957);
nor U9214 (N_9214,N_7845,N_6716);
and U9215 (N_9215,N_6683,N_7633);
nor U9216 (N_9216,N_8444,N_6938);
nand U9217 (N_9217,N_7386,N_6203);
or U9218 (N_9218,N_7303,N_8062);
nand U9219 (N_9219,N_7717,N_7193);
or U9220 (N_9220,N_6166,N_6124);
or U9221 (N_9221,N_6082,N_8340);
nor U9222 (N_9222,N_6554,N_6879);
nor U9223 (N_9223,N_8953,N_6540);
and U9224 (N_9224,N_8103,N_7062);
or U9225 (N_9225,N_7246,N_8303);
and U9226 (N_9226,N_7279,N_7607);
and U9227 (N_9227,N_7133,N_8238);
nor U9228 (N_9228,N_8084,N_6848);
or U9229 (N_9229,N_8707,N_8126);
nand U9230 (N_9230,N_7320,N_8067);
or U9231 (N_9231,N_7232,N_8912);
nand U9232 (N_9232,N_6641,N_8030);
and U9233 (N_9233,N_7167,N_6775);
nand U9234 (N_9234,N_8036,N_6158);
nor U9235 (N_9235,N_7420,N_8275);
nor U9236 (N_9236,N_6971,N_6537);
and U9237 (N_9237,N_8041,N_8661);
or U9238 (N_9238,N_6465,N_6136);
nor U9239 (N_9239,N_6986,N_8347);
and U9240 (N_9240,N_6705,N_7599);
nand U9241 (N_9241,N_8034,N_6193);
nand U9242 (N_9242,N_8374,N_8809);
nand U9243 (N_9243,N_7984,N_6621);
nand U9244 (N_9244,N_7147,N_8850);
or U9245 (N_9245,N_8223,N_6023);
nand U9246 (N_9246,N_8172,N_6660);
nand U9247 (N_9247,N_6127,N_6282);
nand U9248 (N_9248,N_7642,N_8794);
or U9249 (N_9249,N_7885,N_6741);
or U9250 (N_9250,N_6628,N_6071);
and U9251 (N_9251,N_7354,N_6330);
nor U9252 (N_9252,N_7806,N_8201);
or U9253 (N_9253,N_6463,N_8066);
or U9254 (N_9254,N_7413,N_8569);
and U9255 (N_9255,N_7004,N_7711);
nor U9256 (N_9256,N_6601,N_6459);
and U9257 (N_9257,N_7935,N_8064);
or U9258 (N_9258,N_7729,N_7908);
or U9259 (N_9259,N_8920,N_8665);
and U9260 (N_9260,N_6479,N_8174);
and U9261 (N_9261,N_7491,N_6847);
nand U9262 (N_9262,N_7973,N_6667);
nand U9263 (N_9263,N_7095,N_8829);
nor U9264 (N_9264,N_7389,N_7471);
and U9265 (N_9265,N_7160,N_7965);
nor U9266 (N_9266,N_7804,N_8280);
or U9267 (N_9267,N_7499,N_6780);
or U9268 (N_9268,N_7883,N_7110);
nor U9269 (N_9269,N_7666,N_7226);
or U9270 (N_9270,N_8319,N_8991);
or U9271 (N_9271,N_6261,N_7713);
nand U9272 (N_9272,N_6672,N_6441);
or U9273 (N_9273,N_8616,N_8048);
and U9274 (N_9274,N_8902,N_6325);
nand U9275 (N_9275,N_8731,N_8476);
nor U9276 (N_9276,N_6889,N_6246);
nand U9277 (N_9277,N_6015,N_7923);
or U9278 (N_9278,N_8186,N_7472);
nand U9279 (N_9279,N_8735,N_8525);
nand U9280 (N_9280,N_8563,N_8878);
nor U9281 (N_9281,N_8118,N_6543);
nand U9282 (N_9282,N_6988,N_8012);
nand U9283 (N_9283,N_6615,N_8718);
nor U9284 (N_9284,N_7915,N_6717);
nand U9285 (N_9285,N_6752,N_6388);
or U9286 (N_9286,N_8672,N_7460);
nand U9287 (N_9287,N_8367,N_6216);
or U9288 (N_9288,N_7615,N_6098);
and U9289 (N_9289,N_7641,N_8930);
or U9290 (N_9290,N_8083,N_6336);
or U9291 (N_9291,N_7048,N_6570);
and U9292 (N_9292,N_7526,N_8936);
and U9293 (N_9293,N_8094,N_7239);
nand U9294 (N_9294,N_7757,N_8440);
or U9295 (N_9295,N_7085,N_8424);
nor U9296 (N_9296,N_8693,N_8191);
nor U9297 (N_9297,N_8924,N_6893);
nor U9298 (N_9298,N_6324,N_7564);
nand U9299 (N_9299,N_7409,N_6605);
or U9300 (N_9300,N_6293,N_7689);
or U9301 (N_9301,N_8608,N_8101);
nor U9302 (N_9302,N_8371,N_6839);
nand U9303 (N_9303,N_8968,N_7730);
and U9304 (N_9304,N_6414,N_6235);
or U9305 (N_9305,N_6782,N_7870);
or U9306 (N_9306,N_7387,N_8671);
or U9307 (N_9307,N_7925,N_7691);
and U9308 (N_9308,N_6908,N_8326);
or U9309 (N_9309,N_8382,N_8207);
or U9310 (N_9310,N_6538,N_8542);
and U9311 (N_9311,N_6924,N_7549);
nor U9312 (N_9312,N_6663,N_8974);
nor U9313 (N_9313,N_6712,N_8229);
nor U9314 (N_9314,N_6757,N_7777);
nand U9315 (N_9315,N_6973,N_7144);
nand U9316 (N_9316,N_8045,N_7924);
nor U9317 (N_9317,N_6688,N_6115);
nand U9318 (N_9318,N_8777,N_7545);
nand U9319 (N_9319,N_8032,N_6653);
nand U9320 (N_9320,N_7358,N_6386);
and U9321 (N_9321,N_8245,N_7291);
and U9322 (N_9322,N_8337,N_6496);
nor U9323 (N_9323,N_6151,N_6909);
and U9324 (N_9324,N_6837,N_7527);
and U9325 (N_9325,N_7953,N_6460);
or U9326 (N_9326,N_6170,N_7941);
nand U9327 (N_9327,N_8098,N_7723);
and U9328 (N_9328,N_8594,N_8265);
and U9329 (N_9329,N_6905,N_6755);
nand U9330 (N_9330,N_7937,N_8137);
or U9331 (N_9331,N_8584,N_7435);
nand U9332 (N_9332,N_7415,N_7759);
nor U9333 (N_9333,N_8318,N_6534);
xnor U9334 (N_9334,N_6027,N_7672);
nor U9335 (N_9335,N_7685,N_8432);
and U9336 (N_9336,N_8977,N_6194);
or U9337 (N_9337,N_8916,N_7515);
and U9338 (N_9338,N_7288,N_7008);
and U9339 (N_9339,N_6639,N_7210);
or U9340 (N_9340,N_7061,N_6532);
or U9341 (N_9341,N_7766,N_7862);
and U9342 (N_9342,N_6997,N_7518);
nor U9343 (N_9343,N_6991,N_8293);
or U9344 (N_9344,N_8538,N_6950);
or U9345 (N_9345,N_6845,N_6299);
and U9346 (N_9346,N_6344,N_6644);
and U9347 (N_9347,N_6877,N_7251);
nor U9348 (N_9348,N_7720,N_6928);
nand U9349 (N_9349,N_8622,N_8133);
nand U9350 (N_9350,N_6042,N_6146);
and U9351 (N_9351,N_6177,N_7921);
or U9352 (N_9352,N_6896,N_7846);
nand U9353 (N_9353,N_7630,N_7531);
and U9354 (N_9354,N_8379,N_8443);
nand U9355 (N_9355,N_7443,N_8022);
nand U9356 (N_9356,N_8218,N_8446);
nor U9357 (N_9357,N_8952,N_6400);
nor U9358 (N_9358,N_6996,N_8161);
and U9359 (N_9359,N_7731,N_6163);
and U9360 (N_9360,N_6439,N_8754);
nand U9361 (N_9361,N_6935,N_6978);
nor U9362 (N_9362,N_7861,N_7137);
or U9363 (N_9363,N_6831,N_6793);
nand U9364 (N_9364,N_8096,N_8717);
nor U9365 (N_9365,N_7150,N_6652);
nor U9366 (N_9366,N_6800,N_7171);
nand U9367 (N_9367,N_7715,N_8157);
and U9368 (N_9368,N_6587,N_7620);
or U9369 (N_9369,N_7794,N_8602);
and U9370 (N_9370,N_8792,N_7113);
and U9371 (N_9371,N_7719,N_8831);
nor U9372 (N_9372,N_8506,N_6188);
nand U9373 (N_9373,N_8647,N_6514);
or U9374 (N_9374,N_6154,N_6858);
or U9375 (N_9375,N_8772,N_6581);
nand U9376 (N_9376,N_8260,N_7002);
or U9377 (N_9377,N_6995,N_8771);
nand U9378 (N_9378,N_7751,N_8768);
nor U9379 (N_9379,N_6801,N_8242);
nand U9380 (N_9380,N_8020,N_7697);
nand U9381 (N_9381,N_7153,N_8356);
nor U9382 (N_9382,N_6897,N_6284);
and U9383 (N_9383,N_6817,N_6315);
nor U9384 (N_9384,N_7140,N_8397);
nand U9385 (N_9385,N_8895,N_7287);
nand U9386 (N_9386,N_8960,N_7212);
or U9387 (N_9387,N_7250,N_6061);
or U9388 (N_9388,N_7285,N_7975);
nand U9389 (N_9389,N_6006,N_7817);
nor U9390 (N_9390,N_8766,N_8938);
or U9391 (N_9391,N_7490,N_8927);
nor U9392 (N_9392,N_6623,N_8167);
or U9393 (N_9393,N_6237,N_8404);
nor U9394 (N_9394,N_8272,N_7605);
nand U9395 (N_9395,N_8349,N_7240);
nor U9396 (N_9396,N_8135,N_8562);
and U9397 (N_9397,N_8738,N_7922);
nand U9398 (N_9398,N_8958,N_6018);
or U9399 (N_9399,N_7053,N_6499);
or U9400 (N_9400,N_8657,N_6632);
nand U9401 (N_9401,N_6415,N_7822);
or U9402 (N_9402,N_6501,N_7145);
nand U9403 (N_9403,N_8209,N_7635);
and U9404 (N_9404,N_8596,N_6637);
and U9405 (N_9405,N_7555,N_7779);
nor U9406 (N_9406,N_7036,N_7116);
nand U9407 (N_9407,N_6762,N_8818);
nand U9408 (N_9408,N_6077,N_7894);
or U9409 (N_9409,N_8641,N_6678);
nor U9410 (N_9410,N_8421,N_6539);
and U9411 (N_9411,N_8278,N_8035);
nor U9412 (N_9412,N_7069,N_7465);
or U9413 (N_9413,N_6390,N_6328);
or U9414 (N_9414,N_6487,N_7758);
nand U9415 (N_9415,N_7634,N_8615);
and U9416 (N_9416,N_8803,N_8626);
and U9417 (N_9417,N_7445,N_7046);
or U9418 (N_9418,N_6967,N_6220);
nand U9419 (N_9419,N_7265,N_6795);
nor U9420 (N_9420,N_8913,N_8171);
or U9421 (N_9421,N_8791,N_6475);
or U9422 (N_9422,N_6825,N_6427);
and U9423 (N_9423,N_8510,N_8274);
nor U9424 (N_9424,N_6087,N_6590);
and U9425 (N_9425,N_6332,N_7800);
nor U9426 (N_9426,N_8142,N_6529);
nor U9427 (N_9427,N_8418,N_8919);
nand U9428 (N_9428,N_8428,N_8950);
or U9429 (N_9429,N_6128,N_6713);
and U9430 (N_9430,N_6408,N_8307);
or U9431 (N_9431,N_8598,N_8132);
and U9432 (N_9432,N_6160,N_6832);
nand U9433 (N_9433,N_7122,N_7955);
or U9434 (N_9434,N_6552,N_6733);
nand U9435 (N_9435,N_8776,N_6887);
and U9436 (N_9436,N_6798,N_8964);
and U9437 (N_9437,N_6304,N_7222);
and U9438 (N_9438,N_8080,N_8026);
nor U9439 (N_9439,N_7913,N_8909);
nand U9440 (N_9440,N_7688,N_6221);
nor U9441 (N_9441,N_6147,N_8529);
and U9442 (N_9442,N_8997,N_7565);
nand U9443 (N_9443,N_8037,N_7466);
and U9444 (N_9444,N_7896,N_8890);
nor U9445 (N_9445,N_6108,N_7289);
and U9446 (N_9446,N_6205,N_6714);
and U9447 (N_9447,N_8703,N_6274);
nand U9448 (N_9448,N_7993,N_6041);
and U9449 (N_9449,N_8677,N_6616);
nand U9450 (N_9450,N_7414,N_7591);
nor U9451 (N_9451,N_7871,N_6642);
or U9452 (N_9452,N_6784,N_6271);
nand U9453 (N_9453,N_7182,N_6114);
or U9454 (N_9454,N_7559,N_6586);
and U9455 (N_9455,N_6109,N_7437);
nand U9456 (N_9456,N_7535,N_7770);
nand U9457 (N_9457,N_7159,N_6503);
nor U9458 (N_9458,N_8998,N_8117);
or U9459 (N_9459,N_8536,N_8730);
nor U9460 (N_9460,N_7475,N_7943);
nor U9461 (N_9461,N_8859,N_8090);
nand U9462 (N_9462,N_6574,N_6904);
nand U9463 (N_9463,N_8273,N_8180);
nor U9464 (N_9464,N_7393,N_7534);
or U9465 (N_9465,N_6990,N_6738);
nor U9466 (N_9466,N_8785,N_6086);
nor U9467 (N_9467,N_7547,N_7829);
nand U9468 (N_9468,N_7063,N_7999);
and U9469 (N_9469,N_7818,N_6322);
nor U9470 (N_9470,N_8249,N_8300);
nand U9471 (N_9471,N_7722,N_6308);
or U9472 (N_9472,N_7865,N_8961);
and U9473 (N_9473,N_8549,N_6240);
and U9474 (N_9474,N_6185,N_8670);
and U9475 (N_9475,N_7906,N_6876);
nand U9476 (N_9476,N_6596,N_8148);
or U9477 (N_9477,N_6002,N_8130);
nor U9478 (N_9478,N_7514,N_6416);
nand U9479 (N_9479,N_8001,N_7236);
and U9480 (N_9480,N_7676,N_6159);
nand U9481 (N_9481,N_6121,N_7151);
or U9482 (N_9482,N_6335,N_6003);
xor U9483 (N_9483,N_8749,N_6947);
nand U9484 (N_9484,N_8775,N_7496);
and U9485 (N_9485,N_7995,N_7312);
xnor U9486 (N_9486,N_6310,N_7726);
or U9487 (N_9487,N_6525,N_6458);
and U9488 (N_9488,N_7143,N_8146);
and U9489 (N_9489,N_8741,N_8826);
nor U9490 (N_9490,N_7361,N_8454);
nor U9491 (N_9491,N_6946,N_8505);
and U9492 (N_9492,N_8574,N_7868);
and U9493 (N_9493,N_6851,N_8586);
or U9494 (N_9494,N_8740,N_6936);
nand U9495 (N_9495,N_6664,N_7293);
nand U9496 (N_9496,N_8884,N_6341);
nor U9497 (N_9497,N_6860,N_8774);
and U9498 (N_9498,N_8087,N_7257);
or U9499 (N_9499,N_7337,N_7919);
or U9500 (N_9500,N_6462,N_8076);
or U9501 (N_9501,N_8119,N_7980);
and U9502 (N_9502,N_7877,N_8734);
and U9503 (N_9503,N_7566,N_7773);
nor U9504 (N_9504,N_6676,N_8589);
or U9505 (N_9505,N_8695,N_6821);
or U9506 (N_9506,N_6403,N_6944);
or U9507 (N_9507,N_6482,N_6278);
or U9508 (N_9508,N_7343,N_8860);
and U9509 (N_9509,N_7416,N_7674);
xnor U9510 (N_9510,N_6250,N_7775);
or U9511 (N_9511,N_8981,N_8752);
or U9512 (N_9512,N_6276,N_6417);
nor U9513 (N_9513,N_6378,N_7658);
or U9514 (N_9514,N_7914,N_6437);
and U9515 (N_9515,N_6366,N_8407);
nor U9516 (N_9516,N_7314,N_8996);
and U9517 (N_9517,N_8267,N_7589);
or U9518 (N_9518,N_6766,N_7680);
nor U9519 (N_9519,N_7714,N_7376);
nor U9520 (N_9520,N_7199,N_8013);
nand U9521 (N_9521,N_8857,N_8491);
nand U9522 (N_9522,N_7148,N_8004);
nand U9523 (N_9523,N_7206,N_7185);
and U9524 (N_9524,N_7211,N_7315);
or U9525 (N_9525,N_6096,N_6057);
and U9526 (N_9526,N_6577,N_8870);
nor U9527 (N_9527,N_8748,N_8365);
nor U9528 (N_9528,N_7015,N_6443);
nor U9529 (N_9529,N_6999,N_6720);
nand U9530 (N_9530,N_8007,N_8378);
and U9531 (N_9531,N_6046,N_8351);
or U9532 (N_9532,N_7434,N_6392);
nand U9533 (N_9533,N_8954,N_6228);
or U9534 (N_9534,N_8464,N_8617);
nor U9535 (N_9535,N_7074,N_8292);
xor U9536 (N_9536,N_8079,N_8475);
or U9537 (N_9537,N_6091,N_6239);
and U9538 (N_9538,N_7608,N_8175);
or U9539 (N_9539,N_7622,N_6661);
or U9540 (N_9540,N_8116,N_8868);
nor U9541 (N_9541,N_7394,N_7058);
nor U9542 (N_9542,N_7825,N_8892);
nand U9543 (N_9543,N_8907,N_6449);
and U9544 (N_9544,N_6070,N_7699);
nand U9545 (N_9545,N_7594,N_7976);
and U9546 (N_9546,N_7784,N_6794);
or U9547 (N_9547,N_6191,N_6187);
nand U9548 (N_9548,N_8618,N_7368);
nor U9549 (N_9549,N_6974,N_6970);
and U9550 (N_9550,N_7592,N_8701);
and U9551 (N_9551,N_7348,N_7936);
and U9552 (N_9552,N_6867,N_6917);
nand U9553 (N_9553,N_7272,N_8176);
nand U9554 (N_9554,N_6608,N_8383);
or U9555 (N_9555,N_8605,N_6419);
and U9556 (N_9556,N_6342,N_8266);
and U9557 (N_9557,N_6105,N_7117);
nor U9558 (N_9558,N_6613,N_7778);
nand U9559 (N_9559,N_8526,N_7484);
and U9560 (N_9560,N_8642,N_7245);
or U9561 (N_9561,N_8871,N_7202);
or U9562 (N_9562,N_6617,N_8712);
or U9563 (N_9563,N_8983,N_7056);
or U9564 (N_9564,N_6588,N_8197);
nor U9565 (N_9565,N_7686,N_8561);
nand U9566 (N_9566,N_8869,N_7334);
and U9567 (N_9567,N_8283,N_8102);
nor U9568 (N_9568,N_8935,N_6609);
and U9569 (N_9569,N_7651,N_8335);
nor U9570 (N_9570,N_6138,N_6181);
nand U9571 (N_9571,N_7422,N_6542);
or U9572 (N_9572,N_8305,N_7606);
nand U9573 (N_9573,N_7803,N_8984);
nor U9574 (N_9574,N_8816,N_8989);
or U9575 (N_9575,N_8387,N_7649);
nor U9576 (N_9576,N_7170,N_7269);
nand U9577 (N_9577,N_7673,N_7080);
nand U9578 (N_9578,N_6709,N_8697);
nor U9579 (N_9579,N_6526,N_8801);
nand U9580 (N_9580,N_8941,N_6387);
and U9581 (N_9581,N_6984,N_7039);
or U9582 (N_9582,N_7242,N_8944);
nor U9583 (N_9583,N_8591,N_7836);
nor U9584 (N_9584,N_7667,N_6504);
nand U9585 (N_9585,N_8417,N_7120);
nand U9586 (N_9586,N_6295,N_6826);
or U9587 (N_9587,N_6927,N_7560);
nor U9588 (N_9588,N_7235,N_6556);
or U9589 (N_9589,N_6771,N_6636);
nor U9590 (N_9590,N_7909,N_6824);
or U9591 (N_9591,N_8762,N_8742);
nand U9592 (N_9592,N_8298,N_7059);
nand U9593 (N_9593,N_6610,N_8519);
and U9594 (N_9594,N_6788,N_8252);
and U9595 (N_9595,N_7377,N_6279);
or U9596 (N_9596,N_8192,N_6433);
nor U9597 (N_9597,N_6037,N_8481);
or U9598 (N_9598,N_8289,N_7742);
nor U9599 (N_9599,N_8385,N_7843);
or U9600 (N_9600,N_7292,N_8547);
or U9601 (N_9601,N_7109,N_6702);
or U9602 (N_9602,N_7588,N_8106);
nand U9603 (N_9603,N_8582,N_6424);
or U9604 (N_9604,N_6930,N_6648);
and U9605 (N_9605,N_6783,N_7963);
nor U9606 (N_9606,N_8018,N_6345);
nand U9607 (N_9607,N_8183,N_6696);
nand U9608 (N_9608,N_6157,N_6369);
or U9609 (N_9609,N_8553,N_8508);
nand U9610 (N_9610,N_8810,N_6662);
and U9611 (N_9611,N_7031,N_6007);
xnor U9612 (N_9612,N_7650,N_7665);
nor U9613 (N_9613,N_8603,N_8675);
nand U9614 (N_9614,N_8324,N_6384);
nor U9615 (N_9615,N_6464,N_8971);
nand U9616 (N_9616,N_6891,N_6079);
or U9617 (N_9617,N_8328,N_6728);
and U9618 (N_9618,N_8761,N_6226);
and U9619 (N_9619,N_6446,N_6700);
and U9620 (N_9620,N_7807,N_8939);
or U9621 (N_9621,N_8473,N_6684);
nor U9622 (N_9622,N_6888,N_8993);
or U9623 (N_9623,N_7971,N_8270);
or U9624 (N_9624,N_8254,N_7989);
and U9625 (N_9625,N_7886,N_6506);
or U9626 (N_9626,N_6477,N_7581);
nor U9627 (N_9627,N_7463,N_8728);
or U9628 (N_9628,N_7345,N_6302);
and U9629 (N_9629,N_7900,N_6451);
nand U9630 (N_9630,N_8405,N_8904);
nand U9631 (N_9631,N_7017,N_7256);
or U9632 (N_9632,N_8959,N_6225);
nor U9633 (N_9633,N_8211,N_7603);
or U9634 (N_9634,N_8951,N_8495);
or U9635 (N_9635,N_8704,N_7146);
nor U9636 (N_9636,N_7332,N_8049);
or U9637 (N_9637,N_7184,N_8429);
or U9638 (N_9638,N_8769,N_8908);
or U9639 (N_9639,N_7512,N_7529);
nand U9640 (N_9640,N_6488,N_8674);
nand U9641 (N_9641,N_7933,N_7190);
xor U9642 (N_9642,N_6306,N_8459);
and U9643 (N_9643,N_7483,N_6806);
nor U9644 (N_9644,N_7942,N_6232);
nor U9645 (N_9645,N_8350,N_8844);
nor U9646 (N_9646,N_8441,N_6998);
nand U9647 (N_9647,N_7799,N_7433);
and U9648 (N_9648,N_6179,N_8389);
nand U9649 (N_9649,N_7801,N_7668);
nand U9650 (N_9650,N_6708,N_8808);
nor U9651 (N_9651,N_8750,N_7179);
nor U9652 (N_9652,N_6816,N_6764);
nor U9653 (N_9653,N_6823,N_8522);
or U9654 (N_9654,N_6707,N_6268);
and U9655 (N_9655,N_8753,N_8842);
nand U9656 (N_9656,N_6189,N_8259);
and U9657 (N_9657,N_6283,N_8688);
nand U9658 (N_9658,N_8263,N_6494);
nor U9659 (N_9659,N_7598,N_7838);
or U9660 (N_9660,N_8956,N_7186);
nand U9661 (N_9661,N_8492,N_8685);
or U9662 (N_9662,N_7441,N_8162);
nor U9663 (N_9663,N_8614,N_6726);
or U9664 (N_9664,N_8394,N_6380);
nor U9665 (N_9665,N_7282,N_8121);
nand U9666 (N_9666,N_7175,N_7075);
and U9667 (N_9667,N_6643,N_6582);
or U9668 (N_9668,N_8757,N_7436);
or U9669 (N_9669,N_8839,N_6355);
nor U9670 (N_9670,N_6430,N_7840);
nand U9671 (N_9671,N_6028,N_8338);
and U9672 (N_9672,N_6039,N_8559);
nand U9673 (N_9673,N_7583,N_7724);
nor U9674 (N_9674,N_6192,N_6550);
or U9675 (N_9675,N_7716,N_6937);
nor U9676 (N_9676,N_6370,N_8795);
xor U9677 (N_9677,N_8922,N_8656);
nor U9678 (N_9678,N_8551,N_7277);
nand U9679 (N_9679,N_7189,N_7967);
or U9680 (N_9680,N_7732,N_8416);
nor U9681 (N_9681,N_8755,N_8937);
or U9682 (N_9682,N_6902,N_8632);
nand U9683 (N_9683,N_7271,N_8445);
nor U9684 (N_9684,N_6357,N_6011);
or U9685 (N_9685,N_7839,N_8756);
nor U9686 (N_9686,N_8751,N_8471);
and U9687 (N_9687,N_8431,N_7064);
nor U9688 (N_9688,N_6418,N_8250);
nand U9689 (N_9689,N_8081,N_7573);
and U9690 (N_9690,N_6675,N_8364);
and U9691 (N_9691,N_6214,N_7934);
or U9692 (N_9692,N_8227,N_6983);
and U9693 (N_9693,N_6535,N_8363);
and U9694 (N_9694,N_7164,N_7950);
nor U9695 (N_9695,N_6478,N_6407);
and U9696 (N_9696,N_6354,N_6152);
or U9697 (N_9697,N_6808,N_7224);
or U9698 (N_9698,N_7243,N_8344);
and U9699 (N_9699,N_7461,N_6059);
or U9700 (N_9700,N_8784,N_6373);
nor U9701 (N_9701,N_7338,N_6666);
nor U9702 (N_9702,N_7007,N_7026);
nor U9703 (N_9703,N_7972,N_8609);
nor U9704 (N_9704,N_6956,N_6915);
or U9705 (N_9705,N_6361,N_7352);
or U9706 (N_9706,N_6172,N_7546);
nand U9707 (N_9707,N_7797,N_7939);
nand U9708 (N_9708,N_7582,N_7892);
or U9709 (N_9709,N_8659,N_6343);
nand U9710 (N_9710,N_7944,N_7539);
and U9711 (N_9711,N_6923,N_7959);
or U9712 (N_9712,N_6715,N_8060);
nand U9713 (N_9713,N_7796,N_6691);
nor U9714 (N_9714,N_6804,N_6572);
and U9715 (N_9715,N_6833,N_7927);
nand U9716 (N_9716,N_6196,N_8653);
nand U9717 (N_9717,N_7308,N_8676);
or U9718 (N_9718,N_6523,N_6627);
nor U9719 (N_9719,N_8600,N_7077);
or U9720 (N_9720,N_8843,N_6050);
and U9721 (N_9721,N_8391,N_7671);
and U9722 (N_9722,N_6682,N_8686);
nand U9723 (N_9723,N_6669,N_8360);
or U9724 (N_9724,N_6123,N_6773);
nor U9725 (N_9725,N_6107,N_6655);
and U9726 (N_9726,N_7359,N_6687);
and U9727 (N_9727,N_7533,N_6611);
nand U9728 (N_9728,N_6072,N_7567);
and U9729 (N_9729,N_7562,N_8095);
xor U9730 (N_9730,N_6319,N_6852);
or U9731 (N_9731,N_6894,N_7764);
nand U9732 (N_9732,N_8743,N_7099);
nor U9733 (N_9733,N_6218,N_7019);
and U9734 (N_9734,N_8419,N_8005);
nand U9735 (N_9735,N_7962,N_6362);
or U9736 (N_9736,N_7813,N_8339);
nor U9737 (N_9737,N_8501,N_7609);
nand U9738 (N_9738,N_7554,N_8193);
nand U9739 (N_9739,N_8872,N_8918);
nor U9740 (N_9740,N_7841,N_7169);
or U9741 (N_9741,N_7494,N_8286);
nor U9742 (N_9742,N_7270,N_6918);
or U9743 (N_9743,N_6981,N_6679);
or U9744 (N_9744,N_6555,N_7018);
or U9745 (N_9745,N_6413,N_6505);
or U9746 (N_9746,N_6518,N_8056);
or U9747 (N_9747,N_7351,N_8516);
and U9748 (N_9748,N_6763,N_7503);
nor U9749 (N_9749,N_7012,N_7188);
or U9750 (N_9750,N_7220,N_7785);
nor U9751 (N_9751,N_7492,N_7442);
nor U9752 (N_9752,N_6869,N_7501);
and U9753 (N_9753,N_7572,N_8556);
and U9754 (N_9754,N_7094,N_6318);
and U9755 (N_9755,N_6466,N_8422);
nand U9756 (N_9756,N_8629,N_8327);
nand U9757 (N_9757,N_6979,N_8520);
and U9758 (N_9758,N_7595,N_7540);
nand U9759 (N_9759,N_8125,N_7444);
or U9760 (N_9760,N_6242,N_8945);
nor U9761 (N_9761,N_7382,N_8886);
and U9762 (N_9762,N_6992,N_7357);
nor U9763 (N_9763,N_6878,N_8448);
and U9764 (N_9764,N_7684,N_8219);
and U9765 (N_9765,N_8699,N_7558);
nor U9766 (N_9766,N_8855,N_6659);
nor U9767 (N_9767,N_7166,N_7737);
and U9768 (N_9768,N_7459,N_6993);
nor U9769 (N_9769,N_6273,N_7979);
nand U9770 (N_9770,N_6863,N_6485);
and U9771 (N_9771,N_7419,N_7872);
and U9772 (N_9772,N_6634,N_6389);
nand U9773 (N_9773,N_8706,N_8107);
nand U9774 (N_9774,N_6677,N_7905);
nor U9775 (N_9775,N_6960,N_8411);
or U9776 (N_9776,N_8213,N_8926);
and U9777 (N_9777,N_8184,N_7791);
nand U9778 (N_9778,N_8648,N_6656);
or U9779 (N_9779,N_7192,N_7991);
nor U9780 (N_9780,N_8243,N_6751);
or U9781 (N_9781,N_7648,N_6243);
nor U9782 (N_9782,N_6802,N_8812);
nor U9783 (N_9783,N_7115,N_6090);
nand U9784 (N_9784,N_6975,N_7692);
nand U9785 (N_9785,N_6874,N_7851);
nor U9786 (N_9786,N_6234,N_7468);
nor U9787 (N_9787,N_8806,N_7313);
and U9788 (N_9788,N_8302,N_7336);
or U9789 (N_9789,N_7707,N_6903);
nand U9790 (N_9790,N_8925,N_6772);
or U9791 (N_9791,N_8541,N_6789);
nor U9792 (N_9792,N_8251,N_7678);
nand U9793 (N_9793,N_7467,N_7430);
nor U9794 (N_9794,N_6933,N_8480);
or U9795 (N_9795,N_6339,N_7013);
and U9796 (N_9796,N_8637,N_7011);
and U9797 (N_9797,N_6076,N_7833);
and U9798 (N_9798,N_6178,N_8323);
and U9799 (N_9799,N_7852,N_6383);
and U9800 (N_9800,N_7752,N_7640);
and U9801 (N_9801,N_7623,N_8426);
and U9802 (N_9802,N_6167,N_6805);
xor U9803 (N_9803,N_6272,N_7217);
nor U9804 (N_9804,N_7134,N_7275);
and U9805 (N_9805,N_8845,N_8535);
nand U9806 (N_9806,N_8963,N_8694);
nor U9807 (N_9807,N_8088,N_7097);
and U9808 (N_9808,N_8151,N_6931);
nor U9809 (N_9809,N_6065,N_8114);
nor U9810 (N_9810,N_8815,N_8343);
or U9811 (N_9811,N_8141,N_6372);
or U9812 (N_9812,N_8246,N_8150);
nor U9813 (N_9813,N_7780,N_7478);
or U9814 (N_9814,N_7010,N_8716);
and U9815 (N_9815,N_6803,N_7215);
nor U9816 (N_9816,N_7618,N_8739);
and U9817 (N_9817,N_7073,N_7874);
or U9818 (N_9818,N_8858,N_8619);
or U9819 (N_9819,N_7016,N_8138);
nor U9820 (N_9820,N_8767,N_7636);
and U9821 (N_9821,N_8235,N_7958);
nor U9822 (N_9822,N_7111,N_7997);
nor U9823 (N_9823,N_6381,N_8539);
and U9824 (N_9824,N_8380,N_8268);
or U9825 (N_9825,N_7808,N_7005);
and U9826 (N_9826,N_8413,N_7297);
or U9827 (N_9827,N_7426,N_6965);
nand U9828 (N_9828,N_8100,N_8031);
nor U9829 (N_9829,N_6265,N_7086);
and U9830 (N_9830,N_6068,N_8865);
nand U9831 (N_9831,N_6131,N_6008);
nor U9832 (N_9832,N_6531,N_6340);
and U9833 (N_9833,N_7194,N_6350);
or U9834 (N_9834,N_8401,N_7479);
and U9835 (N_9835,N_7745,N_8282);
or U9836 (N_9836,N_7788,N_8099);
nor U9837 (N_9837,N_7195,N_8438);
nor U9838 (N_9838,N_6814,N_6113);
nand U9839 (N_9839,N_8819,N_6141);
and U9840 (N_9840,N_7066,N_8470);
nand U9841 (N_9841,N_7847,N_7304);
nand U9842 (N_9842,N_8377,N_8372);
nand U9843 (N_9843,N_8077,N_7378);
or U9844 (N_9844,N_8225,N_6566);
nor U9845 (N_9845,N_7911,N_8468);
nor U9846 (N_9846,N_7300,N_6428);
or U9847 (N_9847,N_8046,N_8838);
or U9848 (N_9848,N_6391,N_7372);
and U9849 (N_9849,N_6311,N_6737);
nor U9850 (N_9850,N_6084,N_8970);
nand U9851 (N_9851,N_8856,N_7610);
nand U9852 (N_9852,N_7043,N_7286);
nor U9853 (N_9853,N_6750,N_8091);
nand U9854 (N_9854,N_7421,N_7396);
or U9855 (N_9855,N_7306,N_6670);
nor U9856 (N_9856,N_8427,N_7333);
nor U9857 (N_9857,N_7706,N_8376);
nor U9858 (N_9858,N_7753,N_6547);
and U9859 (N_9859,N_6049,N_6612);
nand U9860 (N_9860,N_8932,N_7079);
or U9861 (N_9861,N_8579,N_6512);
or U9862 (N_9862,N_6807,N_8072);
and U9863 (N_9863,N_6297,N_7948);
nor U9864 (N_9864,N_7219,N_6215);
or U9865 (N_9865,N_7299,N_8240);
nand U9866 (N_9866,N_8649,N_7165);
and U9867 (N_9867,N_6710,N_7646);
or U9868 (N_9868,N_6175,N_7174);
or U9869 (N_9869,N_7366,N_7809);
and U9870 (N_9870,N_6173,N_6657);
nor U9871 (N_9871,N_7469,N_6060);
nand U9872 (N_9872,N_6052,N_6573);
and U9873 (N_9873,N_7034,N_8628);
and U9874 (N_9874,N_8866,N_8381);
nand U9875 (N_9875,N_6094,N_8957);
nand U9876 (N_9876,N_6323,N_7455);
nand U9877 (N_9877,N_6953,N_6680);
or U9878 (N_9878,N_7917,N_7410);
and U9879 (N_9879,N_8361,N_7510);
or U9880 (N_9880,N_7104,N_6092);
or U9881 (N_9881,N_7952,N_8625);
nand U9882 (N_9882,N_8159,N_6850);
and U9883 (N_9883,N_7241,N_6922);
nor U9884 (N_9884,N_6934,N_6029);
nor U9885 (N_9885,N_6650,N_7302);
nor U9886 (N_9886,N_6412,N_8727);
nand U9887 (N_9887,N_6792,N_8112);
and U9888 (N_9888,N_6592,N_7542);
nor U9889 (N_9889,N_6200,N_8269);
nor U9890 (N_9890,N_8059,N_8092);
nand U9891 (N_9891,N_6749,N_7626);
nor U9892 (N_9892,N_8021,N_7163);
nand U9893 (N_9893,N_6363,N_8849);
nand U9894 (N_9894,N_7341,N_6571);
or U9895 (N_9895,N_6892,N_7065);
nand U9896 (N_9896,N_8331,N_6962);
nor U9897 (N_9897,N_8841,N_7464);
or U9898 (N_9898,N_8917,N_6186);
nand U9899 (N_9899,N_7637,N_8975);
nand U9900 (N_9900,N_6075,N_7907);
and U9901 (N_9901,N_6777,N_8705);
and U9902 (N_9902,N_7569,N_6204);
nand U9903 (N_9903,N_7187,N_6467);
nand U9904 (N_9904,N_8316,N_8783);
nor U9905 (N_9905,N_7994,N_7050);
or U9906 (N_9906,N_7579,N_7446);
nand U9907 (N_9907,N_7294,N_8122);
or U9908 (N_9908,N_6399,N_6600);
nor U9909 (N_9909,N_7231,N_8644);
and U9910 (N_9910,N_8550,N_8832);
or U9911 (N_9911,N_6560,N_7624);
and U9912 (N_9912,N_7947,N_6150);
and U9913 (N_9913,N_7996,N_6010);
or U9914 (N_9914,N_7233,N_8173);
nand U9915 (N_9915,N_6491,N_7135);
and U9916 (N_9916,N_6614,N_7644);
and U9917 (N_9917,N_8304,N_7728);
and U9918 (N_9918,N_6912,N_8571);
nor U9919 (N_9919,N_7087,N_7548);
or U9920 (N_9920,N_7107,N_7488);
and U9921 (N_9921,N_7022,N_7932);
or U9922 (N_9922,N_6119,N_7473);
or U9923 (N_9923,N_8931,N_7694);
nor U9924 (N_9924,N_6420,N_6043);
or U9925 (N_9925,N_7810,N_6155);
or U9926 (N_9926,N_6781,N_8296);
and U9927 (N_9927,N_6073,N_7670);
nand U9928 (N_9928,N_8987,N_8620);
nand U9929 (N_9929,N_8504,N_6942);
nor U9930 (N_9930,N_8244,N_8284);
nand U9931 (N_9931,N_7453,N_6314);
or U9932 (N_9932,N_8709,N_7238);
and U9933 (N_9933,N_6476,N_7497);
nor U9934 (N_9934,N_8713,N_8667);
nor U9935 (N_9935,N_6622,N_8852);
or U9936 (N_9936,N_7596,N_7428);
nand U9937 (N_9937,N_7196,N_8724);
or U9938 (N_9938,N_6966,N_8285);
nor U9939 (N_9939,N_6862,N_8576);
and U9940 (N_9940,N_7438,N_7532);
and U9941 (N_9941,N_7088,N_6557);
and U9942 (N_9942,N_7261,N_6180);
xor U9943 (N_9943,N_6731,N_7701);
or U9944 (N_9944,N_6718,N_6125);
and U9945 (N_9945,N_7856,N_6292);
and U9946 (N_9946,N_7570,N_7888);
or U9947 (N_9947,N_8643,N_7142);
nand U9948 (N_9948,N_6759,N_8164);
and U9949 (N_9949,N_8113,N_6066);
or U9950 (N_9950,N_8486,N_8627);
and U9951 (N_9951,N_6397,N_8462);
nand U9952 (N_9952,N_8210,N_7655);
nand U9953 (N_9953,N_7051,N_6522);
nor U9954 (N_9954,N_8881,N_8540);
and U9955 (N_9955,N_6585,N_8992);
and U9956 (N_9956,N_8297,N_6447);
nor U9957 (N_9957,N_8607,N_7735);
nand U9958 (N_9958,N_7168,N_7362);
nor U9959 (N_9959,N_6401,N_6519);
or U9960 (N_9960,N_8568,N_6394);
and U9961 (N_9961,N_7384,N_8638);
nor U9962 (N_9962,N_8003,N_7639);
or U9963 (N_9963,N_6649,N_6665);
nand U9964 (N_9964,N_8315,N_8071);
nand U9965 (N_9965,N_7627,N_8291);
or U9966 (N_9966,N_6822,N_7067);
or U9967 (N_9967,N_6134,N_7912);
or U9968 (N_9968,N_7966,N_8140);
and U9969 (N_9969,N_7663,N_8942);
or U9970 (N_9970,N_8502,N_8669);
nand U9971 (N_9971,N_8277,N_7710);
and U9972 (N_9972,N_6248,N_7887);
or U9973 (N_9973,N_7344,N_8978);
and U9974 (N_9974,N_6333,N_8636);
and U9975 (N_9975,N_7266,N_7578);
and U9976 (N_9976,N_7857,N_6719);
and U9977 (N_9977,N_7949,N_7654);
nand U9978 (N_9978,N_8985,N_6236);
nor U9979 (N_9979,N_7230,N_8894);
nand U9980 (N_9980,N_6747,N_8078);
and U9981 (N_9981,N_7687,N_7309);
or U9982 (N_9982,N_8847,N_7889);
and U9983 (N_9983,N_8554,N_7956);
or U9984 (N_9984,N_8747,N_8055);
and U9985 (N_9985,N_8239,N_8764);
and U9986 (N_9986,N_7968,N_6697);
nor U9987 (N_9987,N_8436,N_6165);
nor U9988 (N_9988,N_7252,N_7873);
or U9989 (N_9989,N_7216,N_8015);
nor U9990 (N_9990,N_8948,N_7792);
and U9991 (N_9991,N_7025,N_7815);
nand U9992 (N_9992,N_8645,N_6103);
nor U9993 (N_9993,N_7693,N_6921);
nand U9994 (N_9994,N_6729,N_8543);
nor U9995 (N_9995,N_7072,N_8410);
and U9996 (N_9996,N_7487,N_7495);
or U9997 (N_9997,N_8264,N_7456);
nor U9998 (N_9998,N_7904,N_6358);
nand U9999 (N_9999,N_6195,N_7318);
nor U10000 (N_10000,N_6565,N_6758);
and U10001 (N_10001,N_6130,N_6210);
nor U10002 (N_10002,N_8217,N_7070);
nand U10003 (N_10003,N_8458,N_8597);
nor U10004 (N_10004,N_6253,N_8188);
nor U10005 (N_10005,N_7881,N_7207);
nor U10006 (N_10006,N_8915,N_6866);
nand U10007 (N_10007,N_8507,N_8500);
nand U10008 (N_10008,N_8369,N_7978);
or U10009 (N_10009,N_7399,N_7957);
nand U10010 (N_10010,N_8317,N_6033);
nand U10011 (N_10011,N_8247,N_8786);
xor U10012 (N_10012,N_8679,N_7373);
or U10013 (N_10013,N_8682,N_8166);
nand U10014 (N_10014,N_6468,N_6047);
and U10015 (N_10015,N_7367,N_7586);
and U10016 (N_10016,N_8232,N_8409);
and U10017 (N_10017,N_7157,N_6484);
nand U10018 (N_10018,N_8256,N_6647);
nand U10019 (N_10019,N_7477,N_6580);
or U10020 (N_10020,N_7895,N_6943);
or U10021 (N_10021,N_6301,N_6721);
or U10022 (N_10022,N_6626,N_6761);
or U10023 (N_10023,N_6558,N_6454);
nor U10024 (N_10024,N_8897,N_7431);
and U10025 (N_10025,N_7449,N_6030);
nor U10026 (N_10026,N_6875,N_8308);
and U10027 (N_10027,N_8104,N_8450);
nor U10028 (N_10028,N_6285,N_6645);
nand U10029 (N_10029,N_8472,N_6252);
nor U10030 (N_10030,N_7552,N_6453);
and U10031 (N_10031,N_8982,N_8683);
nor U10032 (N_10032,N_8070,N_8965);
and U10033 (N_10033,N_6730,N_7047);
and U10034 (N_10034,N_8797,N_6834);
nand U10035 (N_10035,N_6820,N_7910);
nor U10036 (N_10036,N_8127,N_7457);
nor U10037 (N_10037,N_6461,N_6206);
or U10038 (N_10038,N_8154,N_7832);
or U10039 (N_10039,N_6148,N_7055);
or U10040 (N_10040,N_8836,N_7100);
nor U10041 (N_10041,N_6727,N_8359);
nand U10042 (N_10042,N_6945,N_6334);
nor U10043 (N_10043,N_8262,N_6184);
nor U10044 (N_10044,N_6009,N_6607);
or U10045 (N_10045,N_7823,N_6940);
or U10046 (N_10046,N_7786,N_6040);
or U10047 (N_10047,N_7858,N_6735);
nor U10048 (N_10048,N_6349,N_6563);
and U10049 (N_10049,N_6815,N_8560);
nand U10050 (N_10050,N_6785,N_7076);
or U10051 (N_10051,N_6901,N_6143);
xor U10052 (N_10052,N_6132,N_7850);
nand U10053 (N_10053,N_7863,N_7090);
and U10054 (N_10054,N_6633,N_6987);
and U10055 (N_10055,N_8969,N_8311);
xor U10056 (N_10056,N_8011,N_8514);
and U10057 (N_10057,N_6083,N_8355);
and U10058 (N_10058,N_7511,N_8177);
nand U10059 (N_10059,N_8650,N_8732);
nor U10060 (N_10060,N_8570,N_8876);
and U10061 (N_10061,N_7009,N_7214);
and U10062 (N_10062,N_8781,N_6673);
or U10063 (N_10063,N_8862,N_6117);
and U10064 (N_10064,N_7375,N_8955);
or U10065 (N_10065,N_8710,N_8006);
and U10066 (N_10066,N_8517,N_7054);
or U10067 (N_10067,N_6190,N_6835);
nand U10068 (N_10068,N_7044,N_8215);
or U10069 (N_10069,N_8189,N_6085);
nor U10070 (N_10070,N_7397,N_8069);
or U10071 (N_10071,N_6742,N_7204);
or U10072 (N_10072,N_8583,N_6256);
or U10073 (N_10073,N_8430,N_7408);
or U10074 (N_10074,N_6267,N_6069);
and U10075 (N_10075,N_7225,N_7893);
nor U10076 (N_10076,N_7508,N_6048);
nand U10077 (N_10077,N_7749,N_8152);
or U10078 (N_10078,N_7407,N_6511);
nor U10079 (N_10079,N_6396,N_7556);
or U10080 (N_10080,N_8465,N_7551);
nor U10081 (N_10081,N_7398,N_6575);
and U10082 (N_10082,N_8910,N_8879);
nand U10083 (N_10083,N_7869,N_8592);
and U10084 (N_10084,N_7124,N_8453);
nor U10085 (N_10085,N_7916,N_6140);
and U10086 (N_10086,N_6368,N_8490);
nand U10087 (N_10087,N_6277,N_7802);
nor U10088 (N_10088,N_6122,N_8976);
nand U10089 (N_10089,N_6836,N_8725);
and U10090 (N_10090,N_7108,N_7317);
nand U10091 (N_10091,N_7550,N_7754);
nand U10092 (N_10092,N_7027,N_8488);
xor U10093 (N_10093,N_7611,N_7830);
and U10094 (N_10094,N_8640,N_8375);
nand U10095 (N_10095,N_8530,N_8370);
and U10096 (N_10096,N_6360,N_6095);
or U10097 (N_10097,N_8052,N_7585);
and U10098 (N_10098,N_6241,N_7208);
nor U10099 (N_10099,N_6797,N_6471);
nand U10100 (N_10100,N_8469,N_7082);
and U10101 (N_10101,N_6541,N_8271);
and U10102 (N_10102,N_6929,N_8853);
or U10103 (N_10103,N_8002,N_7954);
xnor U10104 (N_10104,N_7854,N_6972);
or U10105 (N_10105,N_8433,N_6685);
nor U10106 (N_10106,N_7946,N_8312);
nand U10107 (N_10107,N_6490,N_7176);
and U10108 (N_10108,N_8109,N_8390);
and U10109 (N_10109,N_6654,N_7793);
or U10110 (N_10110,N_7866,N_6230);
nand U10111 (N_10111,N_7538,N_6838);
and U10112 (N_10112,N_7652,N_8943);
nor U10113 (N_10113,N_6118,N_8896);
nor U10114 (N_10114,N_6211,N_6864);
xor U10115 (N_10115,N_8580,N_6842);
and U10116 (N_10116,N_8093,N_8558);
and U10117 (N_10117,N_6671,N_7712);
and U10118 (N_10118,N_8780,N_7696);
nand U10119 (N_10119,N_8384,N_8900);
and U10120 (N_10120,N_6275,N_6080);
and U10121 (N_10121,N_6900,N_7931);
and U10122 (N_10122,N_8577,N_6013);
nand U10123 (N_10123,N_8129,N_6409);
nand U10124 (N_10124,N_7374,N_7698);
and U10125 (N_10125,N_6920,N_8817);
nor U10126 (N_10126,N_6110,N_7734);
nand U10127 (N_10127,N_6385,N_6890);
nor U10128 (N_10128,N_7580,N_8973);
and U10129 (N_10129,N_8198,N_8182);
and U10130 (N_10130,N_8461,N_6619);
and U10131 (N_10131,N_7703,N_6559);
and U10132 (N_10132,N_8050,N_6312);
nand U10133 (N_10133,N_7161,N_7383);
nand U10134 (N_10134,N_8581,N_8058);
nor U10135 (N_10135,N_7365,N_8714);
or U10136 (N_10136,N_6474,N_7750);
nand U10137 (N_10137,N_7324,N_6120);
and U10138 (N_10138,N_6739,N_6161);
or U10139 (N_10139,N_6142,N_8398);
and U10140 (N_10140,N_6101,N_7156);
or U10141 (N_10141,N_8692,N_7675);
nor U10142 (N_10142,N_8478,N_8696);
and U10143 (N_10143,N_8395,N_6919);
nand U10144 (N_10144,N_7385,N_6846);
xor U10145 (N_10145,N_6337,N_8527);
and U10146 (N_10146,N_8206,N_8236);
nor U10147 (N_10147,N_8039,N_6162);
nor U10148 (N_10148,N_8299,N_6331);
nand U10149 (N_10149,N_6217,N_8875);
or U10150 (N_10150,N_7273,N_6365);
or U10151 (N_10151,N_8241,N_8528);
nor U10152 (N_10152,N_7960,N_8000);
nor U10153 (N_10153,N_8123,N_8873);
and U10154 (N_10154,N_6377,N_8044);
or U10155 (N_10155,N_7481,N_8565);
and U10156 (N_10156,N_8222,N_7427);
xor U10157 (N_10157,N_6026,N_8947);
nand U10158 (N_10158,N_6245,N_6508);
nand U10159 (N_10159,N_7504,N_8798);
nand U10160 (N_10160,N_6809,N_7191);
and U10161 (N_10161,N_6382,N_6000);
nand U10162 (N_10162,N_7340,N_7557);
or U10163 (N_10163,N_7523,N_6133);
and U10164 (N_10164,N_8822,N_7462);
or U10165 (N_10165,N_8833,N_6753);
and U10166 (N_10166,N_6489,N_6955);
and U10167 (N_10167,N_7162,N_7218);
nor U10168 (N_10168,N_6509,N_6486);
or U10169 (N_10169,N_6269,N_8008);
and U10170 (N_10170,N_7024,N_6963);
and U10171 (N_10171,N_8053,N_7418);
nor U10172 (N_10172,N_7819,N_8533);
nand U10173 (N_10173,N_6668,N_8124);
nor U10174 (N_10174,N_7201,N_6168);
or U10175 (N_10175,N_6969,N_6448);
or U10176 (N_10176,N_7038,N_7083);
or U10177 (N_10177,N_6251,N_8763);
nand U10178 (N_10178,N_8033,N_6745);
nand U10179 (N_10179,N_7631,N_6227);
and U10180 (N_10180,N_7322,N_6977);
or U10181 (N_10181,N_6583,N_8396);
nor U10182 (N_10182,N_8848,N_7229);
nand U10183 (N_10183,N_8295,N_7812);
or U10184 (N_10184,N_8837,N_6952);
nor U10185 (N_10185,N_7767,N_8515);
nor U10186 (N_10186,N_8009,N_8455);
or U10187 (N_10187,N_7628,N_7103);
and U10188 (N_10188,N_8134,N_8348);
or U10189 (N_10189,N_7390,N_6958);
nand U10190 (N_10190,N_6787,N_8437);
nor U10191 (N_10191,N_7522,N_6321);
nand U10192 (N_10192,N_6932,N_7276);
or U10193 (N_10193,N_7283,N_8253);
and U10194 (N_10194,N_6291,N_8545);
nor U10195 (N_10195,N_7128,N_6199);
or U10196 (N_10196,N_7985,N_7951);
and U10197 (N_10197,N_7574,N_6171);
and U10198 (N_10198,N_7600,N_7391);
nor U10199 (N_10199,N_6495,N_6856);
nand U10200 (N_10200,N_6507,N_7470);
nor U10201 (N_10201,N_8105,N_6262);
and U10202 (N_10202,N_7679,N_6521);
or U10203 (N_10203,N_6144,N_6044);
nand U10204 (N_10204,N_7040,N_7342);
nor U10205 (N_10205,N_6182,N_7563);
or U10206 (N_10206,N_6513,N_7370);
or U10207 (N_10207,N_8085,N_8759);
and U10208 (N_10208,N_7021,N_8089);
or U10209 (N_10209,N_8301,N_6910);
nand U10210 (N_10210,N_8633,N_6723);
and U10211 (N_10211,N_6264,N_8155);
nor U10212 (N_10212,N_6895,N_6674);
nor U10213 (N_10213,N_7781,N_7738);
and U10214 (N_10214,N_8729,N_6062);
or U10215 (N_10215,N_6951,N_8621);
and U10216 (N_10216,N_8726,N_8593);
or U10217 (N_10217,N_8813,N_6100);
or U10218 (N_10218,N_6078,N_8414);
nor U10219 (N_10219,N_6840,N_8980);
and U10220 (N_10220,N_8708,N_7081);
or U10221 (N_10221,N_8063,N_8194);
nand U10222 (N_10222,N_6202,N_7848);
and U10223 (N_10223,N_7789,N_6624);
or U10224 (N_10224,N_7448,N_7695);
nand U10225 (N_10225,N_8487,N_7305);
and U10226 (N_10226,N_7141,N_7814);
and U10227 (N_10227,N_6517,N_7590);
nand U10228 (N_10228,N_6748,N_6681);
nand U10229 (N_10229,N_6316,N_7928);
and U10230 (N_10230,N_6603,N_6602);
or U10231 (N_10231,N_8646,N_7824);
nand U10232 (N_10232,N_8673,N_6258);
nand U10233 (N_10233,N_7198,N_6812);
and U10234 (N_10234,N_8864,N_7613);
nand U10235 (N_10235,N_6690,N_8744);
nand U10236 (N_10236,N_8027,N_7638);
or U10237 (N_10237,N_6116,N_8489);
or U10238 (N_10238,N_6884,N_6829);
xor U10239 (N_10239,N_6352,N_6139);
nor U10240 (N_10240,N_6074,N_6604);
nor U10241 (N_10241,N_6861,N_8325);
and U10242 (N_10242,N_6290,N_8689);
and U10243 (N_10243,N_6527,N_8181);
nand U10244 (N_10244,N_8043,N_6520);
nand U10245 (N_10245,N_6135,N_7274);
and U10246 (N_10246,N_7920,N_8901);
nor U10247 (N_10247,N_8452,N_8199);
nand U10248 (N_10248,N_8214,N_7576);
nor U10249 (N_10249,N_8457,N_6497);
nand U10250 (N_10250,N_8863,N_8820);
nor U10251 (N_10251,N_7323,N_6790);
and U10252 (N_10252,N_6736,N_7057);
nor U10253 (N_10253,N_8016,N_7450);
or U10254 (N_10254,N_6689,N_7125);
and U10255 (N_10255,N_8835,N_8203);
nor U10256 (N_10256,N_8010,N_6546);
nand U10257 (N_10257,N_7553,N_8439);
nand U10258 (N_10258,N_6799,N_6695);
nand U10259 (N_10259,N_7118,N_7772);
and U10260 (N_10260,N_7741,N_7363);
nand U10261 (N_10261,N_7432,N_8787);
nor U10262 (N_10262,N_8828,N_6939);
or U10263 (N_10263,N_7601,N_8358);
or U10264 (N_10264,N_7653,N_8276);
nand U10265 (N_10265,N_7152,N_8420);
and U10266 (N_10266,N_7992,N_8403);
nor U10267 (N_10267,N_6359,N_7974);
nand U10268 (N_10268,N_8068,N_7400);
and U10269 (N_10269,N_6949,N_8075);
nand U10270 (N_10270,N_8846,N_8479);
and U10271 (N_10271,N_6651,N_8588);
nand U10272 (N_10272,N_7918,N_7782);
or U10273 (N_10273,N_7768,N_7525);
and U10274 (N_10274,N_6102,N_7619);
or U10275 (N_10275,N_6183,N_8147);
or U10276 (N_10276,N_8733,N_6686);
nor U10277 (N_10277,N_6768,N_6740);
nor U10278 (N_10278,N_7970,N_7987);
nor U10279 (N_10279,N_7029,N_8678);
and U10280 (N_10280,N_8721,N_6410);
nand U10281 (N_10281,N_8723,N_8760);
and U10282 (N_10282,N_8814,N_8599);
xor U10283 (N_10283,N_7844,N_7945);
or U10284 (N_10284,N_6307,N_6638);
nand U10285 (N_10285,N_6429,N_8460);
and U10286 (N_10286,N_8861,N_8796);
nor U10287 (N_10287,N_6174,N_6423);
or U10288 (N_10288,N_7500,N_7502);
or U10289 (N_10289,N_7223,N_6796);
nand U10290 (N_10290,N_8877,N_8967);
or U10291 (N_10291,N_6926,N_8024);
and U10292 (N_10292,N_8548,N_8400);
and U10293 (N_10293,N_7891,N_7880);
xor U10294 (N_10294,N_8255,N_6064);
and U10295 (N_10295,N_8778,N_7447);
or U10296 (N_10296,N_7092,N_8346);
nand U10297 (N_10297,N_6911,N_7411);
nand U10298 (N_10298,N_6976,N_6865);
or U10299 (N_10299,N_8523,N_6599);
nor U10300 (N_10300,N_6544,N_8687);
nand U10301 (N_10301,N_7402,N_8758);
and U10302 (N_10302,N_6263,N_7718);
or U10303 (N_10303,N_6317,N_8779);
and U10304 (N_10304,N_6067,N_7482);
or U10305 (N_10305,N_6881,N_8143);
and U10306 (N_10306,N_6452,N_7339);
nand U10307 (N_10307,N_7119,N_8179);
nor U10308 (N_10308,N_8208,N_6989);
nand U10309 (N_10309,N_7084,N_7988);
nor U10310 (N_10310,N_8573,N_7281);
nand U10311 (N_10311,N_8668,N_8720);
or U10312 (N_10312,N_7617,N_6054);
and U10313 (N_10313,N_7568,N_6701);
and U10314 (N_10314,N_6961,N_8631);
or U10315 (N_10315,N_6432,N_7505);
or U10316 (N_10316,N_7280,N_6097);
or U10317 (N_10317,N_6238,N_6398);
and U10318 (N_10318,N_6348,N_7253);
nand U10319 (N_10319,N_6510,N_7403);
and U10320 (N_10320,N_8995,N_6198);
nor U10321 (N_10321,N_8373,N_6629);
and U10322 (N_10322,N_7632,N_7664);
and U10323 (N_10323,N_8513,N_8722);
or U10324 (N_10324,N_8212,N_7901);
or U10325 (N_10325,N_7853,N_7260);
nand U10326 (N_10326,N_7327,N_7677);
nand U10327 (N_10327,N_6598,N_6706);
nor U10328 (N_10328,N_8503,N_7577);
and U10329 (N_10329,N_6914,N_6734);
nand U10330 (N_10330,N_7307,N_6774);
or U10331 (N_10331,N_7878,N_7071);
nor U10332 (N_10332,N_7173,N_7902);
nor U10333 (N_10333,N_7842,N_7790);
nand U10334 (N_10334,N_7129,N_8248);
and U10335 (N_10335,N_7228,N_7748);
or U10336 (N_10336,N_7643,N_7023);
nand U10337 (N_10337,N_6035,N_6857);
nor U10338 (N_10338,N_8168,N_8736);
nand U10339 (N_10339,N_6724,N_8933);
or U10340 (N_10340,N_8770,N_6395);
and U10341 (N_10341,N_7940,N_7458);
nor U10342 (N_10342,N_6843,N_7041);
nor U10343 (N_10343,N_6329,N_7669);
nor U10344 (N_10344,N_6870,N_8891);
or U10345 (N_10345,N_7604,N_7130);
or U10346 (N_10346,N_7721,N_7683);
nor U10347 (N_10347,N_6528,N_6483);
nor U10348 (N_10348,N_8914,N_8623);
nor U10349 (N_10349,N_6791,N_7330);
or U10350 (N_10350,N_6298,N_6722);
nor U10351 (N_10351,N_8110,N_8534);
or U10352 (N_10352,N_6703,N_6249);
nor U10353 (N_10353,N_6219,N_6776);
nand U10354 (N_10354,N_6156,N_6492);
or U10355 (N_10355,N_7127,N_8567);
nand U10356 (N_10356,N_8205,N_7969);
nand U10357 (N_10357,N_8261,N_6882);
nor U10358 (N_10358,N_8483,N_8880);
nor U10359 (N_10359,N_7003,N_8196);
or U10360 (N_10360,N_8662,N_7656);
nor U10361 (N_10361,N_8702,N_6498);
or U10362 (N_10362,N_6913,N_8435);
xnor U10363 (N_10363,N_6450,N_8606);
nor U10364 (N_10364,N_6828,N_7682);
and U10365 (N_10365,N_7882,N_7700);
or U10366 (N_10366,N_7405,N_8824);
nand U10367 (N_10367,N_8136,N_6222);
nor U10368 (N_10368,N_8257,N_6954);
or U10369 (N_10369,N_8415,N_8144);
nand U10370 (N_10370,N_7096,N_6099);
nand U10371 (N_10371,N_6819,N_8216);
nand U10372 (N_10372,N_8966,N_7126);
and U10373 (N_10373,N_7254,N_6692);
or U10374 (N_10374,N_7727,N_6968);
nor U10375 (N_10375,N_8788,N_8169);
nor U10376 (N_10376,N_6770,N_8979);
or U10377 (N_10377,N_7060,N_6589);
or U10378 (N_10378,N_8811,N_8139);
nand U10379 (N_10379,N_7733,N_7213);
or U10380 (N_10380,N_7705,N_8893);
nand U10381 (N_10381,N_7353,N_8474);
or U10382 (N_10382,N_7890,N_7262);
nand U10383 (N_10383,N_8929,N_7561);
nor U10384 (N_10384,N_7827,N_8165);
or U10385 (N_10385,N_8341,N_8854);
nand U10386 (N_10386,N_8393,N_7078);
and U10387 (N_10387,N_6055,N_8889);
nand U10388 (N_10388,N_7178,N_7068);
nor U10389 (N_10389,N_8313,N_6270);
nor U10390 (N_10390,N_7513,N_6089);
nor U10391 (N_10391,N_7298,N_8681);
and U10392 (N_10392,N_6568,N_8604);
nand U10393 (N_10393,N_7480,N_6434);
and U10394 (N_10394,N_6841,N_6907);
nand U10395 (N_10395,N_6431,N_8221);
or U10396 (N_10396,N_6853,N_7708);
or U10397 (N_10397,N_7030,N_8544);
nor U10398 (N_10398,N_7811,N_7725);
nor U10399 (N_10399,N_6019,N_8233);
and U10400 (N_10400,N_8566,N_6247);
or U10401 (N_10401,N_7929,N_7424);
xnor U10402 (N_10402,N_7234,N_7587);
nand U10403 (N_10403,N_8399,N_6481);
and U10404 (N_10404,N_6356,N_6038);
and U10405 (N_10405,N_8518,N_7474);
nand U10406 (N_10406,N_8799,N_6287);
nand U10407 (N_10407,N_6500,N_7828);
and U10408 (N_10408,N_8467,N_8711);
and U10409 (N_10409,N_6899,N_8434);
and U10410 (N_10410,N_8202,N_7486);
and U10411 (N_10411,N_8108,N_6244);
or U10412 (N_10412,N_7237,N_7849);
nand U10413 (N_10413,N_7867,N_7098);
nand U10414 (N_10414,N_6704,N_8921);
nand U10415 (N_10415,N_7834,N_7326);
nand U10416 (N_10416,N_7998,N_6137);
nand U10417 (N_10417,N_8220,N_7528);
or U10418 (N_10418,N_6502,N_8575);
nand U10419 (N_10419,N_7439,N_7417);
and U10420 (N_10420,N_8949,N_6435);
or U10421 (N_10421,N_6126,N_8484);
nor U10422 (N_10422,N_8190,N_8639);
or U10423 (N_10423,N_7816,N_7264);
or U10424 (N_10424,N_6106,N_7381);
or U10425 (N_10425,N_6402,N_8765);
nand U10426 (N_10426,N_6374,N_8654);
nor U10427 (N_10427,N_7263,N_8017);
and U10428 (N_10428,N_6562,N_7977);
nand U10429 (N_10429,N_8789,N_8564);
nor U10430 (N_10430,N_8994,N_6438);
nor U10431 (N_10431,N_6025,N_7295);
nand U10432 (N_10432,N_8719,N_6765);
and U10433 (N_10433,N_7930,N_7961);
or U10434 (N_10434,N_8493,N_7903);
nor U10435 (N_10435,N_6201,N_8999);
or U10436 (N_10436,N_6880,N_7369);
nand U10437 (N_10437,N_6813,N_7755);
and U10438 (N_10438,N_8482,N_8463);
and U10439 (N_10439,N_7614,N_8153);
and U10440 (N_10440,N_6699,N_8698);
or U10441 (N_10441,N_7197,N_8333);
nand U10442 (N_10442,N_8555,N_6473);
nand U10443 (N_10443,N_8512,N_8281);
or U10444 (N_10444,N_6545,N_6305);
or U10445 (N_10445,N_6854,N_7049);
nand U10446 (N_10446,N_8851,N_8690);
nor U10447 (N_10447,N_8128,N_6405);
nand U10448 (N_10448,N_8906,N_7798);
nand U10449 (N_10449,N_8178,N_6994);
or U10450 (N_10450,N_8477,N_6286);
nand U10451 (N_10451,N_7981,N_6031);
or U10452 (N_10452,N_6698,N_8825);
nand U10453 (N_10453,N_6016,N_7136);
nand U10454 (N_10454,N_8652,N_7662);
nand U10455 (N_10455,N_8903,N_7033);
and U10456 (N_10456,N_8494,N_7787);
nor U10457 (N_10457,N_7267,N_8773);
or U10458 (N_10458,N_8611,N_8234);
or U10459 (N_10459,N_8684,N_8149);
nand U10460 (N_10460,N_8115,N_8412);
and U10461 (N_10461,N_7498,N_6743);
nand U10462 (N_10462,N_8321,N_6885);
and U10463 (N_10463,N_7227,N_8940);
nor U10464 (N_10464,N_6257,N_6457);
and U10465 (N_10465,N_8074,N_8485);
nand U10466 (N_10466,N_8651,N_8805);
nor U10467 (N_10467,N_8336,N_8793);
and U10468 (N_10468,N_8065,N_8715);
and U10469 (N_10469,N_7290,N_6985);
xnor U10470 (N_10470,N_7661,N_6034);
and U10471 (N_10471,N_8986,N_6625);
or U10472 (N_10472,N_8456,N_6746);
nor U10473 (N_10473,N_7155,N_7200);
nor U10474 (N_10474,N_8231,N_6618);
and U10475 (N_10475,N_7102,N_6364);
or U10476 (N_10476,N_7875,N_7412);
or U10477 (N_10477,N_8612,N_8737);
and U10478 (N_10478,N_8158,N_7321);
nor U10479 (N_10479,N_7739,N_7820);
nand U10480 (N_10480,N_7316,N_8899);
or U10481 (N_10481,N_7837,N_7177);
nor U10482 (N_10482,N_6255,N_6591);
and U10483 (N_10483,N_6259,N_8585);
nand U10484 (N_10484,N_7541,N_8228);
nand U10485 (N_10485,N_6266,N_6469);
and U10486 (N_10486,N_6289,N_8061);
nand U10487 (N_10487,N_8874,N_6470);
and U10488 (N_10488,N_7938,N_6515);
nor U10489 (N_10489,N_7524,N_6493);
and U10490 (N_10490,N_7704,N_7221);
nand U10491 (N_10491,N_8911,N_6012);
and U10492 (N_10492,N_6769,N_6548);
nor U10493 (N_10493,N_7183,N_7543);
nor U10494 (N_10494,N_6456,N_6561);
or U10495 (N_10495,N_8572,N_7645);
nor U10496 (N_10496,N_7139,N_8042);
nor U10497 (N_10497,N_6303,N_8309);
or U10498 (N_10498,N_6551,N_6516);
or U10499 (N_10499,N_8664,N_8051);
and U10500 (N_10500,N_6805,N_7293);
nor U10501 (N_10501,N_6891,N_8952);
nor U10502 (N_10502,N_7930,N_7854);
nand U10503 (N_10503,N_6127,N_8354);
or U10504 (N_10504,N_7572,N_6756);
nor U10505 (N_10505,N_8890,N_8648);
xor U10506 (N_10506,N_7162,N_8200);
xnor U10507 (N_10507,N_6625,N_6810);
nor U10508 (N_10508,N_8774,N_6125);
and U10509 (N_10509,N_6293,N_8928);
nor U10510 (N_10510,N_8452,N_6197);
or U10511 (N_10511,N_8839,N_8416);
or U10512 (N_10512,N_8601,N_8798);
or U10513 (N_10513,N_8601,N_8910);
or U10514 (N_10514,N_8147,N_6032);
nor U10515 (N_10515,N_6975,N_6158);
and U10516 (N_10516,N_7783,N_6341);
nand U10517 (N_10517,N_7184,N_6055);
nor U10518 (N_10518,N_8233,N_8966);
nand U10519 (N_10519,N_6236,N_7617);
nand U10520 (N_10520,N_6857,N_6647);
nor U10521 (N_10521,N_8248,N_7694);
and U10522 (N_10522,N_7613,N_7388);
nor U10523 (N_10523,N_7967,N_6826);
and U10524 (N_10524,N_7419,N_7906);
nor U10525 (N_10525,N_8456,N_6253);
nor U10526 (N_10526,N_7577,N_7222);
nor U10527 (N_10527,N_8161,N_8119);
and U10528 (N_10528,N_6678,N_8940);
nand U10529 (N_10529,N_8488,N_6022);
and U10530 (N_10530,N_8727,N_8460);
or U10531 (N_10531,N_8310,N_7889);
nor U10532 (N_10532,N_6427,N_8312);
and U10533 (N_10533,N_7041,N_6352);
nor U10534 (N_10534,N_8144,N_6291);
nor U10535 (N_10535,N_8406,N_6473);
nand U10536 (N_10536,N_8630,N_7273);
or U10537 (N_10537,N_6090,N_6725);
nor U10538 (N_10538,N_8890,N_7822);
and U10539 (N_10539,N_8284,N_6959);
or U10540 (N_10540,N_7357,N_6100);
or U10541 (N_10541,N_7225,N_8717);
and U10542 (N_10542,N_7156,N_7596);
nor U10543 (N_10543,N_7012,N_6245);
or U10544 (N_10544,N_6710,N_6499);
and U10545 (N_10545,N_7875,N_8815);
nand U10546 (N_10546,N_7505,N_6759);
nand U10547 (N_10547,N_7982,N_6201);
or U10548 (N_10548,N_7475,N_7016);
or U10549 (N_10549,N_8660,N_8214);
nand U10550 (N_10550,N_7513,N_6589);
and U10551 (N_10551,N_8845,N_6073);
and U10552 (N_10552,N_6378,N_8498);
nor U10553 (N_10553,N_6821,N_6364);
and U10554 (N_10554,N_7149,N_7629);
nor U10555 (N_10555,N_6822,N_8442);
and U10556 (N_10556,N_7732,N_6347);
or U10557 (N_10557,N_6035,N_6992);
and U10558 (N_10558,N_8438,N_8595);
and U10559 (N_10559,N_8659,N_8607);
nand U10560 (N_10560,N_8199,N_7523);
or U10561 (N_10561,N_7274,N_8755);
and U10562 (N_10562,N_8803,N_7401);
nor U10563 (N_10563,N_7582,N_6943);
or U10564 (N_10564,N_8095,N_7314);
nand U10565 (N_10565,N_8596,N_7210);
nor U10566 (N_10566,N_7716,N_6633);
nor U10567 (N_10567,N_8200,N_8982);
or U10568 (N_10568,N_6467,N_8404);
or U10569 (N_10569,N_7448,N_6485);
nor U10570 (N_10570,N_8818,N_7626);
or U10571 (N_10571,N_7694,N_6691);
nand U10572 (N_10572,N_6462,N_8905);
or U10573 (N_10573,N_6669,N_6965);
and U10574 (N_10574,N_7862,N_8113);
and U10575 (N_10575,N_8620,N_6369);
nand U10576 (N_10576,N_7647,N_8256);
and U10577 (N_10577,N_6728,N_7567);
and U10578 (N_10578,N_7986,N_7999);
xnor U10579 (N_10579,N_7024,N_6818);
or U10580 (N_10580,N_7509,N_7636);
and U10581 (N_10581,N_7438,N_6258);
and U10582 (N_10582,N_6762,N_6144);
nor U10583 (N_10583,N_6988,N_6276);
or U10584 (N_10584,N_8462,N_8565);
nand U10585 (N_10585,N_6159,N_7223);
and U10586 (N_10586,N_7789,N_6558);
or U10587 (N_10587,N_6156,N_8749);
nand U10588 (N_10588,N_7586,N_8775);
and U10589 (N_10589,N_6171,N_6794);
nor U10590 (N_10590,N_7916,N_8052);
or U10591 (N_10591,N_8312,N_8150);
or U10592 (N_10592,N_7726,N_6524);
or U10593 (N_10593,N_8988,N_6269);
nand U10594 (N_10594,N_7585,N_6563);
or U10595 (N_10595,N_7673,N_6518);
nor U10596 (N_10596,N_8364,N_6074);
and U10597 (N_10597,N_8695,N_8496);
nand U10598 (N_10598,N_7869,N_7636);
or U10599 (N_10599,N_8677,N_6017);
or U10600 (N_10600,N_8923,N_7957);
nand U10601 (N_10601,N_8367,N_8709);
nand U10602 (N_10602,N_8057,N_7615);
and U10603 (N_10603,N_7358,N_6471);
or U10604 (N_10604,N_6169,N_7647);
nand U10605 (N_10605,N_7482,N_6778);
nand U10606 (N_10606,N_6092,N_6390);
or U10607 (N_10607,N_6101,N_7707);
nand U10608 (N_10608,N_8321,N_8158);
or U10609 (N_10609,N_6089,N_6844);
nand U10610 (N_10610,N_7431,N_7823);
and U10611 (N_10611,N_6911,N_6658);
nand U10612 (N_10612,N_6267,N_8966);
nand U10613 (N_10613,N_6036,N_7486);
and U10614 (N_10614,N_6371,N_8934);
or U10615 (N_10615,N_8459,N_6930);
nor U10616 (N_10616,N_6760,N_6092);
and U10617 (N_10617,N_6444,N_6859);
or U10618 (N_10618,N_8614,N_7148);
nand U10619 (N_10619,N_6746,N_6126);
and U10620 (N_10620,N_8403,N_8385);
nor U10621 (N_10621,N_8616,N_8862);
nand U10622 (N_10622,N_8320,N_8796);
nor U10623 (N_10623,N_8290,N_8280);
or U10624 (N_10624,N_6260,N_7412);
nor U10625 (N_10625,N_7742,N_6102);
and U10626 (N_10626,N_6491,N_7911);
or U10627 (N_10627,N_6394,N_6397);
or U10628 (N_10628,N_8173,N_7411);
xor U10629 (N_10629,N_8641,N_8800);
nor U10630 (N_10630,N_8518,N_7868);
nor U10631 (N_10631,N_6874,N_8092);
nor U10632 (N_10632,N_8588,N_6229);
or U10633 (N_10633,N_7561,N_8096);
nand U10634 (N_10634,N_8923,N_7749);
or U10635 (N_10635,N_6243,N_8503);
or U10636 (N_10636,N_6179,N_7303);
or U10637 (N_10637,N_8479,N_7834);
nand U10638 (N_10638,N_8183,N_7749);
nand U10639 (N_10639,N_7996,N_7955);
and U10640 (N_10640,N_6867,N_6025);
or U10641 (N_10641,N_6842,N_6577);
nand U10642 (N_10642,N_8649,N_6032);
nand U10643 (N_10643,N_8236,N_8759);
and U10644 (N_10644,N_6751,N_8153);
xor U10645 (N_10645,N_7542,N_8636);
nand U10646 (N_10646,N_8162,N_6508);
and U10647 (N_10647,N_7358,N_6248);
nor U10648 (N_10648,N_8994,N_7591);
nor U10649 (N_10649,N_8154,N_7844);
or U10650 (N_10650,N_7292,N_6359);
or U10651 (N_10651,N_6352,N_8007);
nand U10652 (N_10652,N_8173,N_7724);
or U10653 (N_10653,N_8008,N_8393);
or U10654 (N_10654,N_8153,N_7090);
nor U10655 (N_10655,N_7905,N_7837);
or U10656 (N_10656,N_6229,N_8527);
nand U10657 (N_10657,N_6918,N_7194);
nand U10658 (N_10658,N_6470,N_7503);
nor U10659 (N_10659,N_7333,N_8409);
nand U10660 (N_10660,N_6530,N_7963);
nand U10661 (N_10661,N_7690,N_8730);
and U10662 (N_10662,N_7518,N_6216);
and U10663 (N_10663,N_6677,N_6419);
nand U10664 (N_10664,N_8534,N_6695);
or U10665 (N_10665,N_6168,N_8298);
nand U10666 (N_10666,N_8352,N_7375);
nor U10667 (N_10667,N_7294,N_6874);
nand U10668 (N_10668,N_6904,N_7202);
or U10669 (N_10669,N_7894,N_8359);
nand U10670 (N_10670,N_8323,N_8373);
nand U10671 (N_10671,N_6525,N_6301);
and U10672 (N_10672,N_8312,N_7207);
nand U10673 (N_10673,N_6891,N_6554);
nand U10674 (N_10674,N_7715,N_8224);
or U10675 (N_10675,N_6395,N_8861);
or U10676 (N_10676,N_8643,N_6189);
nor U10677 (N_10677,N_6687,N_7908);
nor U10678 (N_10678,N_6861,N_8086);
or U10679 (N_10679,N_6927,N_6068);
nand U10680 (N_10680,N_6120,N_7327);
and U10681 (N_10681,N_7440,N_8890);
nor U10682 (N_10682,N_7854,N_8814);
nor U10683 (N_10683,N_8997,N_7361);
and U10684 (N_10684,N_8035,N_6683);
or U10685 (N_10685,N_7635,N_6547);
nor U10686 (N_10686,N_8382,N_6725);
nor U10687 (N_10687,N_7001,N_8501);
nand U10688 (N_10688,N_8831,N_7289);
or U10689 (N_10689,N_7416,N_7277);
and U10690 (N_10690,N_7158,N_6077);
xor U10691 (N_10691,N_8644,N_8156);
nand U10692 (N_10692,N_7458,N_8506);
or U10693 (N_10693,N_6785,N_7620);
and U10694 (N_10694,N_7566,N_6947);
or U10695 (N_10695,N_7723,N_6565);
and U10696 (N_10696,N_8615,N_7067);
or U10697 (N_10697,N_6854,N_7261);
and U10698 (N_10698,N_6330,N_6832);
and U10699 (N_10699,N_7269,N_7900);
or U10700 (N_10700,N_7248,N_7440);
and U10701 (N_10701,N_6891,N_6917);
or U10702 (N_10702,N_7145,N_6122);
nand U10703 (N_10703,N_6032,N_8027);
and U10704 (N_10704,N_6019,N_7560);
nand U10705 (N_10705,N_7595,N_8623);
and U10706 (N_10706,N_8192,N_6483);
nor U10707 (N_10707,N_7948,N_6826);
nor U10708 (N_10708,N_8694,N_6436);
nand U10709 (N_10709,N_6916,N_8787);
nor U10710 (N_10710,N_7184,N_6530);
nor U10711 (N_10711,N_6709,N_7195);
nor U10712 (N_10712,N_6613,N_7343);
or U10713 (N_10713,N_8807,N_6135);
nor U10714 (N_10714,N_6077,N_8100);
and U10715 (N_10715,N_7894,N_8007);
nor U10716 (N_10716,N_7153,N_8127);
and U10717 (N_10717,N_8118,N_7859);
nand U10718 (N_10718,N_6637,N_8990);
or U10719 (N_10719,N_7146,N_8966);
nor U10720 (N_10720,N_7844,N_7561);
nor U10721 (N_10721,N_7034,N_6973);
nand U10722 (N_10722,N_6586,N_6819);
or U10723 (N_10723,N_6472,N_6687);
nor U10724 (N_10724,N_8722,N_6249);
nor U10725 (N_10725,N_6027,N_6307);
nand U10726 (N_10726,N_6117,N_6536);
nor U10727 (N_10727,N_7311,N_6920);
nand U10728 (N_10728,N_8927,N_7509);
nand U10729 (N_10729,N_6862,N_6371);
nor U10730 (N_10730,N_7281,N_7267);
nand U10731 (N_10731,N_7202,N_7353);
or U10732 (N_10732,N_8150,N_6007);
and U10733 (N_10733,N_8321,N_6916);
nand U10734 (N_10734,N_8902,N_7690);
and U10735 (N_10735,N_8806,N_8605);
or U10736 (N_10736,N_7917,N_6296);
and U10737 (N_10737,N_6221,N_6066);
or U10738 (N_10738,N_7719,N_6457);
or U10739 (N_10739,N_8207,N_8853);
nand U10740 (N_10740,N_7051,N_7993);
or U10741 (N_10741,N_8905,N_7569);
and U10742 (N_10742,N_7323,N_8126);
or U10743 (N_10743,N_7034,N_7053);
nand U10744 (N_10744,N_6182,N_6781);
or U10745 (N_10745,N_7131,N_8032);
nand U10746 (N_10746,N_7508,N_6958);
and U10747 (N_10747,N_8967,N_7731);
and U10748 (N_10748,N_6185,N_8012);
and U10749 (N_10749,N_6133,N_7491);
nand U10750 (N_10750,N_8756,N_7880);
nand U10751 (N_10751,N_8695,N_6027);
and U10752 (N_10752,N_8781,N_6524);
nand U10753 (N_10753,N_7237,N_7993);
and U10754 (N_10754,N_7685,N_7712);
and U10755 (N_10755,N_6311,N_7133);
xnor U10756 (N_10756,N_6840,N_8016);
nand U10757 (N_10757,N_6247,N_7167);
or U10758 (N_10758,N_8191,N_6525);
nor U10759 (N_10759,N_7964,N_8587);
nand U10760 (N_10760,N_8677,N_8198);
nor U10761 (N_10761,N_6179,N_6847);
and U10762 (N_10762,N_6334,N_8979);
or U10763 (N_10763,N_8751,N_8463);
and U10764 (N_10764,N_8384,N_6215);
nor U10765 (N_10765,N_8832,N_8999);
or U10766 (N_10766,N_6090,N_7706);
and U10767 (N_10767,N_7050,N_8791);
nor U10768 (N_10768,N_7922,N_7444);
nand U10769 (N_10769,N_8561,N_8484);
nor U10770 (N_10770,N_7093,N_7287);
or U10771 (N_10771,N_8877,N_7739);
nand U10772 (N_10772,N_8744,N_6341);
nand U10773 (N_10773,N_8864,N_8534);
nor U10774 (N_10774,N_7895,N_6696);
and U10775 (N_10775,N_8881,N_7253);
nand U10776 (N_10776,N_7922,N_7091);
or U10777 (N_10777,N_7408,N_6301);
and U10778 (N_10778,N_7458,N_6742);
nand U10779 (N_10779,N_6025,N_8282);
nand U10780 (N_10780,N_7040,N_7898);
nor U10781 (N_10781,N_7844,N_6383);
and U10782 (N_10782,N_6410,N_8168);
nor U10783 (N_10783,N_8692,N_6636);
or U10784 (N_10784,N_7451,N_6309);
and U10785 (N_10785,N_7094,N_8582);
or U10786 (N_10786,N_8833,N_8357);
and U10787 (N_10787,N_6354,N_7970);
and U10788 (N_10788,N_7847,N_7595);
and U10789 (N_10789,N_8783,N_6346);
nand U10790 (N_10790,N_7301,N_6096);
or U10791 (N_10791,N_8114,N_7670);
and U10792 (N_10792,N_6042,N_8169);
and U10793 (N_10793,N_6558,N_8163);
nor U10794 (N_10794,N_7398,N_6267);
and U10795 (N_10795,N_8851,N_7799);
nor U10796 (N_10796,N_8349,N_6345);
nor U10797 (N_10797,N_6538,N_6310);
or U10798 (N_10798,N_6834,N_7450);
and U10799 (N_10799,N_8099,N_7132);
nor U10800 (N_10800,N_7580,N_7436);
nor U10801 (N_10801,N_8862,N_7265);
nor U10802 (N_10802,N_8311,N_6536);
nand U10803 (N_10803,N_7665,N_6438);
or U10804 (N_10804,N_7511,N_8816);
or U10805 (N_10805,N_8239,N_7753);
nand U10806 (N_10806,N_7833,N_6241);
and U10807 (N_10807,N_8931,N_7800);
nor U10808 (N_10808,N_8120,N_8008);
or U10809 (N_10809,N_7260,N_7298);
and U10810 (N_10810,N_8100,N_6642);
nand U10811 (N_10811,N_8023,N_6645);
and U10812 (N_10812,N_8280,N_6939);
and U10813 (N_10813,N_8298,N_8819);
nor U10814 (N_10814,N_8955,N_7591);
nor U10815 (N_10815,N_8396,N_7321);
nor U10816 (N_10816,N_7681,N_8372);
nand U10817 (N_10817,N_8673,N_7293);
nor U10818 (N_10818,N_8968,N_8402);
nor U10819 (N_10819,N_8064,N_7696);
or U10820 (N_10820,N_6148,N_6535);
and U10821 (N_10821,N_6211,N_6175);
or U10822 (N_10822,N_6919,N_6682);
nand U10823 (N_10823,N_7685,N_7817);
xor U10824 (N_10824,N_8403,N_8846);
or U10825 (N_10825,N_7337,N_7963);
nand U10826 (N_10826,N_6663,N_7388);
or U10827 (N_10827,N_8204,N_8893);
or U10828 (N_10828,N_8241,N_7200);
nand U10829 (N_10829,N_7628,N_7250);
nand U10830 (N_10830,N_7146,N_6610);
or U10831 (N_10831,N_8518,N_8433);
nand U10832 (N_10832,N_6861,N_6784);
nor U10833 (N_10833,N_7453,N_7055);
and U10834 (N_10834,N_7907,N_6711);
nor U10835 (N_10835,N_8299,N_7245);
nor U10836 (N_10836,N_6131,N_8266);
nor U10837 (N_10837,N_7429,N_8789);
or U10838 (N_10838,N_8191,N_7277);
and U10839 (N_10839,N_7352,N_6262);
nor U10840 (N_10840,N_6179,N_6505);
nor U10841 (N_10841,N_7517,N_7184);
and U10842 (N_10842,N_8205,N_8897);
nand U10843 (N_10843,N_6067,N_7770);
or U10844 (N_10844,N_8707,N_7570);
nand U10845 (N_10845,N_6054,N_8265);
nand U10846 (N_10846,N_6436,N_6793);
and U10847 (N_10847,N_7822,N_7589);
nand U10848 (N_10848,N_8704,N_6084);
nor U10849 (N_10849,N_8528,N_8771);
nor U10850 (N_10850,N_7905,N_7237);
nand U10851 (N_10851,N_8346,N_7635);
and U10852 (N_10852,N_6797,N_6887);
and U10853 (N_10853,N_7129,N_7139);
or U10854 (N_10854,N_7279,N_6570);
nor U10855 (N_10855,N_6238,N_8541);
xor U10856 (N_10856,N_6479,N_7680);
nand U10857 (N_10857,N_8512,N_6906);
and U10858 (N_10858,N_6823,N_7384);
nor U10859 (N_10859,N_6140,N_6509);
or U10860 (N_10860,N_7554,N_8924);
and U10861 (N_10861,N_7100,N_8141);
or U10862 (N_10862,N_7115,N_8661);
nor U10863 (N_10863,N_6977,N_7480);
nand U10864 (N_10864,N_6329,N_6459);
or U10865 (N_10865,N_6917,N_7345);
or U10866 (N_10866,N_8398,N_8353);
and U10867 (N_10867,N_6308,N_6499);
and U10868 (N_10868,N_6821,N_6890);
nor U10869 (N_10869,N_6520,N_7789);
nand U10870 (N_10870,N_7846,N_7720);
and U10871 (N_10871,N_6847,N_7158);
nand U10872 (N_10872,N_6456,N_8627);
or U10873 (N_10873,N_6513,N_7390);
nor U10874 (N_10874,N_6436,N_8290);
nor U10875 (N_10875,N_8969,N_8839);
or U10876 (N_10876,N_8941,N_8799);
or U10877 (N_10877,N_8049,N_7717);
and U10878 (N_10878,N_6839,N_7429);
nor U10879 (N_10879,N_6646,N_6894);
nand U10880 (N_10880,N_6965,N_8724);
nand U10881 (N_10881,N_6846,N_6105);
or U10882 (N_10882,N_8411,N_6437);
or U10883 (N_10883,N_7857,N_6357);
or U10884 (N_10884,N_6539,N_6585);
and U10885 (N_10885,N_7730,N_8251);
nand U10886 (N_10886,N_6643,N_7006);
nor U10887 (N_10887,N_8474,N_7514);
and U10888 (N_10888,N_7971,N_7585);
or U10889 (N_10889,N_8896,N_6414);
and U10890 (N_10890,N_8531,N_6367);
and U10891 (N_10891,N_7166,N_8217);
nor U10892 (N_10892,N_7292,N_7984);
nor U10893 (N_10893,N_8391,N_8780);
nand U10894 (N_10894,N_8665,N_7000);
and U10895 (N_10895,N_8521,N_7322);
and U10896 (N_10896,N_7243,N_6881);
or U10897 (N_10897,N_7506,N_7242);
nor U10898 (N_10898,N_7689,N_7798);
nand U10899 (N_10899,N_6949,N_7809);
nor U10900 (N_10900,N_7512,N_7351);
nand U10901 (N_10901,N_7840,N_6498);
and U10902 (N_10902,N_8840,N_6665);
nand U10903 (N_10903,N_7679,N_6058);
or U10904 (N_10904,N_6455,N_8387);
nand U10905 (N_10905,N_7459,N_8133);
and U10906 (N_10906,N_8712,N_7914);
nand U10907 (N_10907,N_8398,N_8575);
nor U10908 (N_10908,N_7076,N_6202);
nand U10909 (N_10909,N_6506,N_6158);
or U10910 (N_10910,N_6913,N_6874);
nor U10911 (N_10911,N_8524,N_8359);
and U10912 (N_10912,N_7992,N_8893);
and U10913 (N_10913,N_6521,N_7358);
nor U10914 (N_10914,N_8789,N_6703);
or U10915 (N_10915,N_6935,N_6500);
nand U10916 (N_10916,N_8937,N_8464);
and U10917 (N_10917,N_8544,N_8822);
nor U10918 (N_10918,N_8495,N_8185);
nor U10919 (N_10919,N_6439,N_7004);
nor U10920 (N_10920,N_7236,N_8808);
nand U10921 (N_10921,N_6446,N_7445);
and U10922 (N_10922,N_7858,N_8715);
and U10923 (N_10923,N_8837,N_6991);
or U10924 (N_10924,N_8978,N_7161);
and U10925 (N_10925,N_7584,N_7276);
nand U10926 (N_10926,N_8111,N_8604);
or U10927 (N_10927,N_6113,N_8507);
and U10928 (N_10928,N_6120,N_7762);
or U10929 (N_10929,N_7711,N_6906);
or U10930 (N_10930,N_7467,N_6831);
or U10931 (N_10931,N_6232,N_6893);
nand U10932 (N_10932,N_7534,N_6068);
or U10933 (N_10933,N_6990,N_7423);
and U10934 (N_10934,N_6319,N_8861);
nand U10935 (N_10935,N_7567,N_8369);
nor U10936 (N_10936,N_6950,N_7978);
nand U10937 (N_10937,N_7003,N_7485);
and U10938 (N_10938,N_6509,N_7583);
nor U10939 (N_10939,N_7805,N_7215);
nand U10940 (N_10940,N_7650,N_6412);
or U10941 (N_10941,N_7363,N_8159);
nand U10942 (N_10942,N_8488,N_6920);
and U10943 (N_10943,N_7226,N_6069);
nand U10944 (N_10944,N_8483,N_6998);
and U10945 (N_10945,N_7908,N_6915);
nor U10946 (N_10946,N_7866,N_8143);
nand U10947 (N_10947,N_7380,N_6642);
and U10948 (N_10948,N_8063,N_7280);
and U10949 (N_10949,N_7269,N_8041);
nand U10950 (N_10950,N_7005,N_7592);
and U10951 (N_10951,N_7435,N_7892);
or U10952 (N_10952,N_8029,N_6195);
and U10953 (N_10953,N_8993,N_8699);
or U10954 (N_10954,N_8824,N_7374);
nand U10955 (N_10955,N_7269,N_8399);
and U10956 (N_10956,N_7163,N_6998);
and U10957 (N_10957,N_6375,N_8972);
or U10958 (N_10958,N_7129,N_8768);
nand U10959 (N_10959,N_6796,N_6699);
nor U10960 (N_10960,N_7332,N_7474);
or U10961 (N_10961,N_8193,N_8839);
nand U10962 (N_10962,N_7623,N_7916);
or U10963 (N_10963,N_8696,N_6485);
or U10964 (N_10964,N_8263,N_7380);
nor U10965 (N_10965,N_6881,N_8504);
and U10966 (N_10966,N_6059,N_6271);
or U10967 (N_10967,N_7387,N_8949);
or U10968 (N_10968,N_8403,N_6534);
and U10969 (N_10969,N_8689,N_6080);
nand U10970 (N_10970,N_6657,N_8805);
nor U10971 (N_10971,N_8963,N_6501);
nand U10972 (N_10972,N_8811,N_7901);
and U10973 (N_10973,N_7810,N_8528);
nand U10974 (N_10974,N_6006,N_7814);
nand U10975 (N_10975,N_6698,N_6056);
and U10976 (N_10976,N_7131,N_6646);
nand U10977 (N_10977,N_7470,N_7399);
and U10978 (N_10978,N_6660,N_8612);
or U10979 (N_10979,N_7773,N_8139);
and U10980 (N_10980,N_6957,N_6769);
nand U10981 (N_10981,N_8057,N_6574);
and U10982 (N_10982,N_8533,N_6618);
and U10983 (N_10983,N_6987,N_8118);
and U10984 (N_10984,N_7291,N_7692);
and U10985 (N_10985,N_6420,N_8748);
and U10986 (N_10986,N_6417,N_8958);
or U10987 (N_10987,N_7175,N_8747);
nor U10988 (N_10988,N_8928,N_7599);
nor U10989 (N_10989,N_7228,N_7682);
and U10990 (N_10990,N_6072,N_7684);
or U10991 (N_10991,N_7591,N_8956);
xnor U10992 (N_10992,N_6175,N_7073);
or U10993 (N_10993,N_8177,N_8509);
or U10994 (N_10994,N_6938,N_6293);
xnor U10995 (N_10995,N_7200,N_7318);
and U10996 (N_10996,N_7832,N_8447);
xor U10997 (N_10997,N_7377,N_8959);
nor U10998 (N_10998,N_6323,N_6371);
nand U10999 (N_10999,N_8155,N_8946);
and U11000 (N_11000,N_6228,N_7211);
nor U11001 (N_11001,N_7723,N_8275);
or U11002 (N_11002,N_7334,N_6832);
nand U11003 (N_11003,N_6080,N_8242);
and U11004 (N_11004,N_6309,N_6048);
or U11005 (N_11005,N_7599,N_8178);
nand U11006 (N_11006,N_8147,N_8223);
nor U11007 (N_11007,N_7576,N_7289);
and U11008 (N_11008,N_7177,N_7108);
and U11009 (N_11009,N_6314,N_7833);
nor U11010 (N_11010,N_8151,N_8247);
xnor U11011 (N_11011,N_7198,N_8588);
and U11012 (N_11012,N_6653,N_7600);
or U11013 (N_11013,N_8438,N_7437);
or U11014 (N_11014,N_7137,N_6645);
nand U11015 (N_11015,N_8829,N_8034);
nand U11016 (N_11016,N_7667,N_8660);
nor U11017 (N_11017,N_8775,N_7512);
and U11018 (N_11018,N_8284,N_7233);
or U11019 (N_11019,N_7074,N_7526);
or U11020 (N_11020,N_7099,N_8034);
or U11021 (N_11021,N_7358,N_8690);
and U11022 (N_11022,N_8618,N_6136);
nor U11023 (N_11023,N_7164,N_6745);
or U11024 (N_11024,N_8399,N_8084);
nor U11025 (N_11025,N_7391,N_8593);
nand U11026 (N_11026,N_6398,N_8299);
and U11027 (N_11027,N_6899,N_7233);
nand U11028 (N_11028,N_7580,N_6224);
and U11029 (N_11029,N_7594,N_6226);
nand U11030 (N_11030,N_6606,N_8351);
or U11031 (N_11031,N_6769,N_7167);
and U11032 (N_11032,N_8171,N_6675);
nand U11033 (N_11033,N_8081,N_8920);
or U11034 (N_11034,N_8212,N_7079);
xor U11035 (N_11035,N_8640,N_8008);
nand U11036 (N_11036,N_6654,N_8365);
nor U11037 (N_11037,N_8080,N_8024);
nand U11038 (N_11038,N_7751,N_8078);
or U11039 (N_11039,N_8184,N_6818);
or U11040 (N_11040,N_8183,N_7898);
nor U11041 (N_11041,N_8928,N_7942);
or U11042 (N_11042,N_6806,N_6389);
or U11043 (N_11043,N_7129,N_6258);
and U11044 (N_11044,N_6815,N_8864);
nand U11045 (N_11045,N_7395,N_6489);
nor U11046 (N_11046,N_8224,N_6638);
nand U11047 (N_11047,N_6981,N_8515);
and U11048 (N_11048,N_6372,N_8806);
nor U11049 (N_11049,N_6221,N_8840);
nand U11050 (N_11050,N_7177,N_8472);
nor U11051 (N_11051,N_6180,N_7999);
nor U11052 (N_11052,N_8911,N_8372);
and U11053 (N_11053,N_7172,N_7901);
nor U11054 (N_11054,N_7433,N_7146);
nand U11055 (N_11055,N_8202,N_8166);
nor U11056 (N_11056,N_7152,N_8745);
nor U11057 (N_11057,N_8422,N_8661);
or U11058 (N_11058,N_8291,N_7006);
and U11059 (N_11059,N_7099,N_7809);
or U11060 (N_11060,N_7257,N_6051);
and U11061 (N_11061,N_7007,N_6946);
and U11062 (N_11062,N_8002,N_6887);
or U11063 (N_11063,N_8439,N_8978);
or U11064 (N_11064,N_7758,N_6558);
xor U11065 (N_11065,N_7025,N_7247);
and U11066 (N_11066,N_8124,N_6622);
and U11067 (N_11067,N_8822,N_7841);
nand U11068 (N_11068,N_8752,N_8891);
or U11069 (N_11069,N_8206,N_8284);
nand U11070 (N_11070,N_6413,N_8218);
or U11071 (N_11071,N_8566,N_7530);
nor U11072 (N_11072,N_8439,N_6467);
or U11073 (N_11073,N_7768,N_7617);
or U11074 (N_11074,N_7761,N_6349);
and U11075 (N_11075,N_8509,N_7278);
and U11076 (N_11076,N_8034,N_7280);
nand U11077 (N_11077,N_6731,N_8153);
nor U11078 (N_11078,N_8787,N_6151);
nor U11079 (N_11079,N_8745,N_7159);
nand U11080 (N_11080,N_6788,N_7406);
nand U11081 (N_11081,N_8099,N_8103);
and U11082 (N_11082,N_7262,N_6418);
or U11083 (N_11083,N_6986,N_8078);
or U11084 (N_11084,N_8220,N_6596);
nand U11085 (N_11085,N_6623,N_8281);
and U11086 (N_11086,N_8341,N_6789);
nand U11087 (N_11087,N_8154,N_7473);
nand U11088 (N_11088,N_6132,N_8538);
xnor U11089 (N_11089,N_8494,N_8919);
or U11090 (N_11090,N_6735,N_8690);
and U11091 (N_11091,N_8841,N_8953);
nor U11092 (N_11092,N_7435,N_8131);
or U11093 (N_11093,N_6199,N_7458);
and U11094 (N_11094,N_7155,N_7531);
nor U11095 (N_11095,N_6442,N_7431);
or U11096 (N_11096,N_7408,N_8112);
nand U11097 (N_11097,N_6748,N_7366);
or U11098 (N_11098,N_8784,N_6893);
and U11099 (N_11099,N_6169,N_7967);
nor U11100 (N_11100,N_6462,N_7172);
nor U11101 (N_11101,N_7301,N_7854);
or U11102 (N_11102,N_7092,N_6689);
nand U11103 (N_11103,N_6995,N_6476);
nor U11104 (N_11104,N_8582,N_7863);
or U11105 (N_11105,N_6399,N_8225);
or U11106 (N_11106,N_8169,N_8551);
nand U11107 (N_11107,N_8923,N_7178);
or U11108 (N_11108,N_7729,N_6565);
or U11109 (N_11109,N_8253,N_8783);
xnor U11110 (N_11110,N_8829,N_7034);
or U11111 (N_11111,N_6047,N_7624);
and U11112 (N_11112,N_7150,N_6226);
and U11113 (N_11113,N_7807,N_7224);
nor U11114 (N_11114,N_7397,N_7787);
and U11115 (N_11115,N_6663,N_8844);
nand U11116 (N_11116,N_6657,N_7431);
nand U11117 (N_11117,N_7420,N_7682);
or U11118 (N_11118,N_6384,N_7893);
nand U11119 (N_11119,N_6948,N_7343);
nand U11120 (N_11120,N_7212,N_7286);
nand U11121 (N_11121,N_6224,N_6292);
nand U11122 (N_11122,N_7846,N_8376);
and U11123 (N_11123,N_7963,N_8684);
and U11124 (N_11124,N_8700,N_6685);
nand U11125 (N_11125,N_8170,N_8507);
nor U11126 (N_11126,N_6383,N_8852);
or U11127 (N_11127,N_8823,N_7273);
and U11128 (N_11128,N_8423,N_8858);
nor U11129 (N_11129,N_8621,N_7780);
nand U11130 (N_11130,N_8285,N_7571);
xor U11131 (N_11131,N_6627,N_6883);
nor U11132 (N_11132,N_6884,N_6826);
nor U11133 (N_11133,N_8080,N_7207);
and U11134 (N_11134,N_7279,N_6332);
or U11135 (N_11135,N_6462,N_6972);
or U11136 (N_11136,N_7502,N_6861);
nor U11137 (N_11137,N_6953,N_8410);
xor U11138 (N_11138,N_8488,N_6378);
or U11139 (N_11139,N_6589,N_7476);
or U11140 (N_11140,N_8529,N_6601);
nand U11141 (N_11141,N_7606,N_7409);
nand U11142 (N_11142,N_8051,N_8670);
or U11143 (N_11143,N_7231,N_6297);
and U11144 (N_11144,N_7317,N_6084);
or U11145 (N_11145,N_8627,N_7105);
and U11146 (N_11146,N_6416,N_8665);
and U11147 (N_11147,N_7068,N_6392);
or U11148 (N_11148,N_6453,N_8276);
xor U11149 (N_11149,N_6940,N_8715);
and U11150 (N_11150,N_6165,N_7477);
nand U11151 (N_11151,N_6941,N_6327);
or U11152 (N_11152,N_6296,N_8953);
or U11153 (N_11153,N_8495,N_7562);
or U11154 (N_11154,N_6698,N_7661);
or U11155 (N_11155,N_6058,N_6478);
nor U11156 (N_11156,N_7600,N_8093);
and U11157 (N_11157,N_7433,N_8465);
or U11158 (N_11158,N_8207,N_8935);
or U11159 (N_11159,N_6325,N_7302);
nand U11160 (N_11160,N_8839,N_8204);
and U11161 (N_11161,N_7218,N_7846);
nand U11162 (N_11162,N_6883,N_6039);
or U11163 (N_11163,N_6319,N_6342);
nand U11164 (N_11164,N_8784,N_6231);
or U11165 (N_11165,N_6848,N_6721);
nand U11166 (N_11166,N_7055,N_6372);
nand U11167 (N_11167,N_6661,N_6309);
or U11168 (N_11168,N_7989,N_6990);
nor U11169 (N_11169,N_8474,N_6949);
nor U11170 (N_11170,N_8195,N_7788);
and U11171 (N_11171,N_6078,N_7288);
and U11172 (N_11172,N_8519,N_7236);
nand U11173 (N_11173,N_6456,N_7543);
nand U11174 (N_11174,N_6543,N_7104);
or U11175 (N_11175,N_7551,N_7897);
nand U11176 (N_11176,N_6861,N_6590);
and U11177 (N_11177,N_6770,N_7930);
or U11178 (N_11178,N_8133,N_6407);
or U11179 (N_11179,N_7038,N_7380);
nand U11180 (N_11180,N_6380,N_7142);
nand U11181 (N_11181,N_7755,N_6148);
nand U11182 (N_11182,N_8786,N_7663);
nor U11183 (N_11183,N_8972,N_7863);
nor U11184 (N_11184,N_6730,N_7783);
or U11185 (N_11185,N_8929,N_7578);
and U11186 (N_11186,N_7527,N_7471);
and U11187 (N_11187,N_7795,N_8962);
nand U11188 (N_11188,N_6717,N_8999);
or U11189 (N_11189,N_6814,N_6004);
nand U11190 (N_11190,N_8220,N_6653);
or U11191 (N_11191,N_6111,N_6284);
nand U11192 (N_11192,N_6434,N_7863);
or U11193 (N_11193,N_7483,N_8171);
or U11194 (N_11194,N_7238,N_8969);
or U11195 (N_11195,N_6485,N_8163);
and U11196 (N_11196,N_7883,N_6971);
nand U11197 (N_11197,N_8046,N_7547);
nand U11198 (N_11198,N_8369,N_6590);
and U11199 (N_11199,N_8824,N_8384);
nand U11200 (N_11200,N_8515,N_6212);
and U11201 (N_11201,N_8392,N_6000);
nand U11202 (N_11202,N_6244,N_8516);
nor U11203 (N_11203,N_6120,N_6203);
and U11204 (N_11204,N_6527,N_7292);
nor U11205 (N_11205,N_6532,N_7395);
nor U11206 (N_11206,N_8850,N_8784);
or U11207 (N_11207,N_6154,N_7369);
and U11208 (N_11208,N_8936,N_7418);
or U11209 (N_11209,N_6687,N_7954);
or U11210 (N_11210,N_8409,N_6259);
and U11211 (N_11211,N_8659,N_7966);
nand U11212 (N_11212,N_8975,N_8114);
or U11213 (N_11213,N_8633,N_6978);
or U11214 (N_11214,N_6947,N_6376);
nor U11215 (N_11215,N_8070,N_7081);
nor U11216 (N_11216,N_7439,N_8806);
nand U11217 (N_11217,N_8051,N_7974);
or U11218 (N_11218,N_7322,N_7209);
nor U11219 (N_11219,N_6731,N_8042);
or U11220 (N_11220,N_8028,N_7094);
and U11221 (N_11221,N_7952,N_6441);
nand U11222 (N_11222,N_7845,N_6072);
or U11223 (N_11223,N_7885,N_7493);
nor U11224 (N_11224,N_7245,N_7710);
or U11225 (N_11225,N_6818,N_7638);
or U11226 (N_11226,N_8191,N_6506);
or U11227 (N_11227,N_8336,N_6282);
nand U11228 (N_11228,N_7510,N_7834);
or U11229 (N_11229,N_7326,N_8296);
and U11230 (N_11230,N_7628,N_6580);
nand U11231 (N_11231,N_6445,N_7100);
xor U11232 (N_11232,N_6352,N_8395);
or U11233 (N_11233,N_7388,N_6652);
nor U11234 (N_11234,N_7650,N_8569);
nand U11235 (N_11235,N_6942,N_6421);
or U11236 (N_11236,N_8040,N_6588);
or U11237 (N_11237,N_7966,N_6939);
or U11238 (N_11238,N_6277,N_8939);
or U11239 (N_11239,N_6522,N_7931);
or U11240 (N_11240,N_7740,N_6445);
and U11241 (N_11241,N_6040,N_7271);
or U11242 (N_11242,N_6692,N_7723);
nand U11243 (N_11243,N_7108,N_6253);
nand U11244 (N_11244,N_7716,N_6151);
nor U11245 (N_11245,N_8776,N_7876);
nand U11246 (N_11246,N_7371,N_7914);
nor U11247 (N_11247,N_7002,N_7344);
and U11248 (N_11248,N_7420,N_8120);
nor U11249 (N_11249,N_8167,N_6304);
nand U11250 (N_11250,N_6496,N_8652);
and U11251 (N_11251,N_8338,N_7140);
or U11252 (N_11252,N_8154,N_8526);
nor U11253 (N_11253,N_6789,N_7660);
nand U11254 (N_11254,N_6319,N_8341);
or U11255 (N_11255,N_8295,N_6213);
nand U11256 (N_11256,N_8890,N_6959);
and U11257 (N_11257,N_7242,N_7138);
and U11258 (N_11258,N_6131,N_8420);
nand U11259 (N_11259,N_8008,N_6260);
and U11260 (N_11260,N_6240,N_7779);
nor U11261 (N_11261,N_8081,N_8892);
or U11262 (N_11262,N_8346,N_8575);
or U11263 (N_11263,N_7052,N_8827);
and U11264 (N_11264,N_6577,N_6819);
nand U11265 (N_11265,N_7300,N_7194);
or U11266 (N_11266,N_8442,N_8751);
nor U11267 (N_11267,N_6623,N_6124);
and U11268 (N_11268,N_8913,N_8438);
nand U11269 (N_11269,N_8262,N_8716);
nand U11270 (N_11270,N_6208,N_8969);
and U11271 (N_11271,N_7037,N_6102);
nand U11272 (N_11272,N_6800,N_6497);
and U11273 (N_11273,N_6822,N_8941);
nor U11274 (N_11274,N_7569,N_7585);
and U11275 (N_11275,N_7117,N_6915);
nor U11276 (N_11276,N_8827,N_7765);
or U11277 (N_11277,N_6120,N_7558);
or U11278 (N_11278,N_8676,N_6802);
or U11279 (N_11279,N_8148,N_8200);
or U11280 (N_11280,N_8291,N_6148);
nand U11281 (N_11281,N_6271,N_8205);
nand U11282 (N_11282,N_6280,N_7035);
and U11283 (N_11283,N_6790,N_8594);
or U11284 (N_11284,N_7419,N_6208);
nor U11285 (N_11285,N_7719,N_6330);
and U11286 (N_11286,N_6665,N_8997);
or U11287 (N_11287,N_6441,N_8491);
or U11288 (N_11288,N_7592,N_8146);
nand U11289 (N_11289,N_6465,N_7413);
nor U11290 (N_11290,N_6385,N_6127);
nor U11291 (N_11291,N_8143,N_8111);
or U11292 (N_11292,N_7052,N_8215);
nor U11293 (N_11293,N_7045,N_7901);
or U11294 (N_11294,N_8078,N_6324);
nor U11295 (N_11295,N_6225,N_7239);
nor U11296 (N_11296,N_6271,N_7540);
nor U11297 (N_11297,N_8875,N_8785);
and U11298 (N_11298,N_7400,N_6670);
or U11299 (N_11299,N_7228,N_6348);
and U11300 (N_11300,N_6830,N_7156);
nor U11301 (N_11301,N_8982,N_8573);
and U11302 (N_11302,N_7495,N_7703);
or U11303 (N_11303,N_6201,N_8929);
nor U11304 (N_11304,N_7614,N_7052);
nor U11305 (N_11305,N_8321,N_6595);
or U11306 (N_11306,N_6911,N_8333);
or U11307 (N_11307,N_6741,N_6721);
nor U11308 (N_11308,N_8521,N_6051);
nor U11309 (N_11309,N_7496,N_8589);
or U11310 (N_11310,N_6791,N_8087);
or U11311 (N_11311,N_6984,N_7028);
nand U11312 (N_11312,N_7283,N_7501);
and U11313 (N_11313,N_8064,N_8978);
and U11314 (N_11314,N_6510,N_8180);
or U11315 (N_11315,N_7189,N_7691);
and U11316 (N_11316,N_8788,N_8075);
nor U11317 (N_11317,N_8532,N_7622);
nor U11318 (N_11318,N_8668,N_6656);
nor U11319 (N_11319,N_6868,N_7923);
or U11320 (N_11320,N_7692,N_6555);
or U11321 (N_11321,N_6161,N_8234);
nor U11322 (N_11322,N_8167,N_7946);
nor U11323 (N_11323,N_7109,N_7773);
nand U11324 (N_11324,N_7190,N_6449);
and U11325 (N_11325,N_6204,N_7850);
or U11326 (N_11326,N_6142,N_7485);
nand U11327 (N_11327,N_8858,N_8751);
nand U11328 (N_11328,N_8760,N_7914);
or U11329 (N_11329,N_7829,N_7822);
and U11330 (N_11330,N_8186,N_8822);
and U11331 (N_11331,N_6643,N_7200);
or U11332 (N_11332,N_7504,N_6838);
or U11333 (N_11333,N_8927,N_8279);
and U11334 (N_11334,N_7415,N_7085);
nor U11335 (N_11335,N_7739,N_6797);
and U11336 (N_11336,N_8784,N_8682);
nand U11337 (N_11337,N_8846,N_8014);
or U11338 (N_11338,N_8025,N_8058);
nand U11339 (N_11339,N_8041,N_7685);
and U11340 (N_11340,N_8956,N_6947);
or U11341 (N_11341,N_6414,N_7738);
nor U11342 (N_11342,N_7845,N_6743);
or U11343 (N_11343,N_6103,N_7371);
nand U11344 (N_11344,N_6894,N_8119);
or U11345 (N_11345,N_8068,N_8627);
and U11346 (N_11346,N_8207,N_6912);
and U11347 (N_11347,N_8417,N_7308);
nand U11348 (N_11348,N_7119,N_6765);
xnor U11349 (N_11349,N_8985,N_6416);
and U11350 (N_11350,N_8250,N_8676);
or U11351 (N_11351,N_6702,N_6219);
and U11352 (N_11352,N_6041,N_8592);
nor U11353 (N_11353,N_7316,N_6587);
and U11354 (N_11354,N_8825,N_7635);
nand U11355 (N_11355,N_6153,N_7636);
or U11356 (N_11356,N_8963,N_7909);
or U11357 (N_11357,N_6629,N_6928);
and U11358 (N_11358,N_7787,N_7758);
nor U11359 (N_11359,N_8769,N_7779);
nor U11360 (N_11360,N_6325,N_6246);
or U11361 (N_11361,N_8993,N_8425);
and U11362 (N_11362,N_6204,N_7828);
and U11363 (N_11363,N_7002,N_8899);
nor U11364 (N_11364,N_7201,N_7586);
or U11365 (N_11365,N_6057,N_7881);
nor U11366 (N_11366,N_7336,N_7413);
and U11367 (N_11367,N_7444,N_8900);
and U11368 (N_11368,N_7866,N_6527);
nor U11369 (N_11369,N_7199,N_8660);
or U11370 (N_11370,N_6231,N_7294);
xnor U11371 (N_11371,N_7118,N_6056);
and U11372 (N_11372,N_6666,N_6208);
and U11373 (N_11373,N_7793,N_8931);
and U11374 (N_11374,N_8542,N_6670);
or U11375 (N_11375,N_8359,N_8614);
nand U11376 (N_11376,N_7180,N_6804);
nand U11377 (N_11377,N_8692,N_8777);
nand U11378 (N_11378,N_7381,N_8916);
nand U11379 (N_11379,N_7863,N_6049);
nand U11380 (N_11380,N_7374,N_8297);
and U11381 (N_11381,N_7193,N_6032);
nand U11382 (N_11382,N_8896,N_7822);
and U11383 (N_11383,N_6812,N_8321);
nand U11384 (N_11384,N_8555,N_7917);
or U11385 (N_11385,N_7465,N_8060);
nand U11386 (N_11386,N_6166,N_7768);
nor U11387 (N_11387,N_6404,N_7735);
or U11388 (N_11388,N_8921,N_6823);
and U11389 (N_11389,N_8727,N_8408);
nand U11390 (N_11390,N_7761,N_6063);
or U11391 (N_11391,N_8979,N_6564);
or U11392 (N_11392,N_7487,N_7579);
or U11393 (N_11393,N_6430,N_6669);
nor U11394 (N_11394,N_7771,N_7794);
or U11395 (N_11395,N_7966,N_7723);
nor U11396 (N_11396,N_6129,N_8798);
nand U11397 (N_11397,N_8366,N_6521);
nand U11398 (N_11398,N_7198,N_6429);
nor U11399 (N_11399,N_7485,N_7053);
and U11400 (N_11400,N_8043,N_7374);
and U11401 (N_11401,N_8828,N_6999);
nand U11402 (N_11402,N_8597,N_6990);
and U11403 (N_11403,N_8100,N_7639);
and U11404 (N_11404,N_6229,N_6374);
and U11405 (N_11405,N_7800,N_7292);
nor U11406 (N_11406,N_8552,N_7486);
or U11407 (N_11407,N_6999,N_7316);
and U11408 (N_11408,N_8282,N_7358);
nand U11409 (N_11409,N_8815,N_6154);
and U11410 (N_11410,N_7185,N_6504);
or U11411 (N_11411,N_7281,N_7328);
and U11412 (N_11412,N_7049,N_7538);
or U11413 (N_11413,N_8609,N_7086);
and U11414 (N_11414,N_8095,N_6570);
nor U11415 (N_11415,N_6303,N_6932);
and U11416 (N_11416,N_6213,N_8833);
or U11417 (N_11417,N_6346,N_7649);
nand U11418 (N_11418,N_7412,N_6640);
nor U11419 (N_11419,N_8964,N_7524);
nand U11420 (N_11420,N_7366,N_8912);
nor U11421 (N_11421,N_7706,N_6176);
nor U11422 (N_11422,N_7981,N_8731);
and U11423 (N_11423,N_8215,N_6390);
or U11424 (N_11424,N_8024,N_7667);
and U11425 (N_11425,N_8092,N_8869);
and U11426 (N_11426,N_6346,N_7807);
or U11427 (N_11427,N_8448,N_6957);
nor U11428 (N_11428,N_7596,N_7120);
and U11429 (N_11429,N_7320,N_8008);
nand U11430 (N_11430,N_6567,N_8909);
and U11431 (N_11431,N_7504,N_6229);
and U11432 (N_11432,N_8642,N_6219);
or U11433 (N_11433,N_6863,N_6536);
or U11434 (N_11434,N_8272,N_6991);
and U11435 (N_11435,N_7909,N_7366);
nor U11436 (N_11436,N_8661,N_6921);
nand U11437 (N_11437,N_6997,N_6534);
nand U11438 (N_11438,N_7916,N_8573);
and U11439 (N_11439,N_8353,N_7144);
nand U11440 (N_11440,N_6122,N_6762);
nor U11441 (N_11441,N_6561,N_6483);
xor U11442 (N_11442,N_7530,N_6605);
or U11443 (N_11443,N_7931,N_8708);
and U11444 (N_11444,N_7090,N_8312);
nand U11445 (N_11445,N_8332,N_6777);
and U11446 (N_11446,N_8387,N_6199);
or U11447 (N_11447,N_7944,N_8033);
and U11448 (N_11448,N_8583,N_8358);
nand U11449 (N_11449,N_7397,N_7405);
and U11450 (N_11450,N_8365,N_8225);
and U11451 (N_11451,N_6102,N_8757);
and U11452 (N_11452,N_6207,N_7195);
and U11453 (N_11453,N_7359,N_6303);
nand U11454 (N_11454,N_6102,N_6192);
xnor U11455 (N_11455,N_8335,N_7903);
and U11456 (N_11456,N_8134,N_7303);
nor U11457 (N_11457,N_6288,N_8364);
or U11458 (N_11458,N_8589,N_6159);
nand U11459 (N_11459,N_8128,N_7864);
and U11460 (N_11460,N_6959,N_7710);
and U11461 (N_11461,N_7933,N_7141);
nor U11462 (N_11462,N_6679,N_6130);
or U11463 (N_11463,N_8471,N_7964);
nor U11464 (N_11464,N_8152,N_8595);
nand U11465 (N_11465,N_7720,N_8399);
nand U11466 (N_11466,N_8620,N_6164);
nor U11467 (N_11467,N_7238,N_7989);
or U11468 (N_11468,N_7502,N_6253);
nor U11469 (N_11469,N_6162,N_6923);
nand U11470 (N_11470,N_6880,N_7822);
nor U11471 (N_11471,N_6916,N_6658);
nor U11472 (N_11472,N_8098,N_7531);
xnor U11473 (N_11473,N_7000,N_7771);
or U11474 (N_11474,N_7116,N_8342);
and U11475 (N_11475,N_6406,N_7695);
nor U11476 (N_11476,N_8487,N_7534);
nor U11477 (N_11477,N_7035,N_7497);
nor U11478 (N_11478,N_7598,N_7988);
or U11479 (N_11479,N_7602,N_7176);
and U11480 (N_11480,N_8098,N_6486);
nor U11481 (N_11481,N_6086,N_7968);
and U11482 (N_11482,N_8818,N_8655);
nand U11483 (N_11483,N_8510,N_8900);
nor U11484 (N_11484,N_7716,N_7517);
and U11485 (N_11485,N_7881,N_6476);
or U11486 (N_11486,N_7627,N_8004);
nor U11487 (N_11487,N_7306,N_7914);
and U11488 (N_11488,N_7813,N_8493);
or U11489 (N_11489,N_6653,N_7069);
nor U11490 (N_11490,N_7878,N_8034);
nand U11491 (N_11491,N_8199,N_8296);
nor U11492 (N_11492,N_6868,N_6461);
and U11493 (N_11493,N_7187,N_6898);
nand U11494 (N_11494,N_6250,N_7984);
nand U11495 (N_11495,N_7313,N_8337);
xnor U11496 (N_11496,N_7593,N_6587);
nor U11497 (N_11497,N_8277,N_6928);
nor U11498 (N_11498,N_8741,N_8940);
and U11499 (N_11499,N_6253,N_6799);
nor U11500 (N_11500,N_6689,N_7319);
nand U11501 (N_11501,N_6624,N_6598);
nand U11502 (N_11502,N_8075,N_6079);
nand U11503 (N_11503,N_6741,N_6596);
nor U11504 (N_11504,N_6679,N_6170);
and U11505 (N_11505,N_7508,N_7109);
nor U11506 (N_11506,N_6248,N_6011);
nand U11507 (N_11507,N_6103,N_6277);
or U11508 (N_11508,N_7283,N_7114);
or U11509 (N_11509,N_7927,N_8947);
and U11510 (N_11510,N_8815,N_6550);
or U11511 (N_11511,N_6393,N_8441);
and U11512 (N_11512,N_8089,N_8833);
and U11513 (N_11513,N_6015,N_8952);
and U11514 (N_11514,N_7531,N_8779);
nor U11515 (N_11515,N_6450,N_7382);
nand U11516 (N_11516,N_7138,N_6256);
or U11517 (N_11517,N_7274,N_8904);
nand U11518 (N_11518,N_7401,N_6647);
or U11519 (N_11519,N_6202,N_7338);
or U11520 (N_11520,N_6304,N_7752);
nand U11521 (N_11521,N_6394,N_6287);
and U11522 (N_11522,N_6482,N_8592);
and U11523 (N_11523,N_7928,N_8820);
nand U11524 (N_11524,N_8559,N_6693);
nand U11525 (N_11525,N_6179,N_7796);
and U11526 (N_11526,N_8071,N_7848);
or U11527 (N_11527,N_7276,N_6436);
nand U11528 (N_11528,N_8584,N_6990);
and U11529 (N_11529,N_7940,N_6802);
or U11530 (N_11530,N_7907,N_8551);
nor U11531 (N_11531,N_6514,N_8169);
nor U11532 (N_11532,N_8394,N_7255);
nor U11533 (N_11533,N_6103,N_6254);
or U11534 (N_11534,N_7190,N_6019);
nor U11535 (N_11535,N_6081,N_7368);
nor U11536 (N_11536,N_6414,N_6098);
and U11537 (N_11537,N_7928,N_8302);
nor U11538 (N_11538,N_8317,N_8107);
nor U11539 (N_11539,N_8461,N_6459);
or U11540 (N_11540,N_6174,N_8511);
nor U11541 (N_11541,N_8278,N_7901);
nor U11542 (N_11542,N_6080,N_8658);
or U11543 (N_11543,N_6343,N_8695);
nor U11544 (N_11544,N_7179,N_6325);
nand U11545 (N_11545,N_6958,N_6769);
nand U11546 (N_11546,N_6566,N_8061);
or U11547 (N_11547,N_7119,N_8201);
nor U11548 (N_11548,N_7936,N_8506);
nand U11549 (N_11549,N_8072,N_6691);
nor U11550 (N_11550,N_8440,N_6248);
nor U11551 (N_11551,N_6799,N_7088);
nand U11552 (N_11552,N_8018,N_6074);
or U11553 (N_11553,N_7007,N_7225);
nand U11554 (N_11554,N_7465,N_6431);
and U11555 (N_11555,N_6883,N_8165);
nand U11556 (N_11556,N_8489,N_8460);
nor U11557 (N_11557,N_6865,N_7735);
or U11558 (N_11558,N_7853,N_8209);
nor U11559 (N_11559,N_7773,N_8246);
nor U11560 (N_11560,N_8434,N_8581);
and U11561 (N_11561,N_6838,N_6399);
and U11562 (N_11562,N_8729,N_6351);
nand U11563 (N_11563,N_6885,N_7414);
and U11564 (N_11564,N_6789,N_7474);
nor U11565 (N_11565,N_6916,N_6882);
or U11566 (N_11566,N_7624,N_8684);
or U11567 (N_11567,N_6110,N_8652);
or U11568 (N_11568,N_8575,N_7817);
nor U11569 (N_11569,N_7461,N_8664);
and U11570 (N_11570,N_8665,N_7263);
or U11571 (N_11571,N_8944,N_8985);
nand U11572 (N_11572,N_6530,N_7263);
and U11573 (N_11573,N_8003,N_7185);
or U11574 (N_11574,N_7380,N_7195);
and U11575 (N_11575,N_7389,N_7729);
nand U11576 (N_11576,N_6072,N_7521);
or U11577 (N_11577,N_8313,N_6161);
and U11578 (N_11578,N_6280,N_8263);
nor U11579 (N_11579,N_7592,N_6981);
and U11580 (N_11580,N_7001,N_6913);
or U11581 (N_11581,N_8754,N_7270);
nor U11582 (N_11582,N_8362,N_6672);
and U11583 (N_11583,N_7258,N_8032);
and U11584 (N_11584,N_7222,N_7762);
or U11585 (N_11585,N_6728,N_6139);
and U11586 (N_11586,N_8058,N_7017);
nor U11587 (N_11587,N_6756,N_7729);
and U11588 (N_11588,N_7854,N_6705);
and U11589 (N_11589,N_8040,N_6939);
nor U11590 (N_11590,N_8717,N_6043);
and U11591 (N_11591,N_7241,N_8975);
or U11592 (N_11592,N_8151,N_6825);
nor U11593 (N_11593,N_7582,N_7751);
nand U11594 (N_11594,N_7397,N_6500);
or U11595 (N_11595,N_8896,N_7402);
or U11596 (N_11596,N_7211,N_8324);
and U11597 (N_11597,N_8832,N_8836);
and U11598 (N_11598,N_6100,N_7432);
nor U11599 (N_11599,N_7165,N_8485);
or U11600 (N_11600,N_7925,N_7621);
nand U11601 (N_11601,N_6594,N_6001);
nand U11602 (N_11602,N_6990,N_8225);
and U11603 (N_11603,N_7898,N_6546);
and U11604 (N_11604,N_8080,N_7904);
and U11605 (N_11605,N_7149,N_6825);
nand U11606 (N_11606,N_8423,N_8056);
nand U11607 (N_11607,N_7617,N_7728);
nand U11608 (N_11608,N_6793,N_8008);
nand U11609 (N_11609,N_7564,N_6968);
nor U11610 (N_11610,N_7244,N_8202);
nor U11611 (N_11611,N_7663,N_8970);
or U11612 (N_11612,N_7795,N_8348);
nand U11613 (N_11613,N_7642,N_7822);
nor U11614 (N_11614,N_8614,N_8958);
or U11615 (N_11615,N_7504,N_8812);
nor U11616 (N_11616,N_7786,N_8096);
or U11617 (N_11617,N_8462,N_6339);
and U11618 (N_11618,N_6473,N_7561);
nor U11619 (N_11619,N_6129,N_8805);
and U11620 (N_11620,N_6892,N_6003);
or U11621 (N_11621,N_7523,N_7749);
nand U11622 (N_11622,N_8488,N_7216);
or U11623 (N_11623,N_7791,N_7931);
and U11624 (N_11624,N_6896,N_6222);
nor U11625 (N_11625,N_6523,N_8729);
nand U11626 (N_11626,N_8840,N_7712);
or U11627 (N_11627,N_8965,N_8508);
and U11628 (N_11628,N_7483,N_8391);
and U11629 (N_11629,N_7121,N_6375);
and U11630 (N_11630,N_6529,N_8053);
nand U11631 (N_11631,N_6099,N_7938);
nor U11632 (N_11632,N_8693,N_7566);
nor U11633 (N_11633,N_6112,N_8674);
or U11634 (N_11634,N_6518,N_7371);
or U11635 (N_11635,N_8278,N_8992);
nand U11636 (N_11636,N_8676,N_6827);
and U11637 (N_11637,N_7491,N_6443);
nand U11638 (N_11638,N_6072,N_7497);
or U11639 (N_11639,N_7911,N_6505);
or U11640 (N_11640,N_6673,N_7928);
or U11641 (N_11641,N_6356,N_8355);
and U11642 (N_11642,N_8409,N_7297);
and U11643 (N_11643,N_6695,N_6597);
or U11644 (N_11644,N_6833,N_7962);
and U11645 (N_11645,N_7495,N_7465);
or U11646 (N_11646,N_6738,N_7483);
nor U11647 (N_11647,N_6404,N_6367);
nor U11648 (N_11648,N_8355,N_6520);
and U11649 (N_11649,N_6027,N_6687);
or U11650 (N_11650,N_8249,N_6273);
nor U11651 (N_11651,N_8213,N_8895);
or U11652 (N_11652,N_8268,N_6523);
nor U11653 (N_11653,N_8493,N_7238);
nor U11654 (N_11654,N_7963,N_6734);
nand U11655 (N_11655,N_7103,N_7481);
nand U11656 (N_11656,N_6814,N_6395);
and U11657 (N_11657,N_8931,N_6744);
nand U11658 (N_11658,N_6408,N_6649);
or U11659 (N_11659,N_6587,N_8411);
or U11660 (N_11660,N_8929,N_6890);
nand U11661 (N_11661,N_6889,N_7793);
and U11662 (N_11662,N_7717,N_8214);
or U11663 (N_11663,N_7632,N_8424);
nand U11664 (N_11664,N_7048,N_6390);
nor U11665 (N_11665,N_7765,N_8838);
nand U11666 (N_11666,N_6135,N_6745);
nand U11667 (N_11667,N_7169,N_8288);
or U11668 (N_11668,N_6946,N_7201);
or U11669 (N_11669,N_7773,N_6431);
or U11670 (N_11670,N_8871,N_7068);
nor U11671 (N_11671,N_7340,N_6046);
and U11672 (N_11672,N_7312,N_6645);
and U11673 (N_11673,N_8036,N_6750);
nand U11674 (N_11674,N_8627,N_6552);
nand U11675 (N_11675,N_8961,N_7668);
nand U11676 (N_11676,N_6766,N_8141);
nor U11677 (N_11677,N_6934,N_7393);
nor U11678 (N_11678,N_6498,N_7489);
nand U11679 (N_11679,N_8771,N_6452);
and U11680 (N_11680,N_7314,N_6422);
nand U11681 (N_11681,N_7994,N_7814);
or U11682 (N_11682,N_8283,N_8748);
and U11683 (N_11683,N_6141,N_7438);
and U11684 (N_11684,N_7800,N_6468);
and U11685 (N_11685,N_6980,N_7671);
or U11686 (N_11686,N_7747,N_7601);
nand U11687 (N_11687,N_6780,N_7232);
nand U11688 (N_11688,N_7688,N_8816);
or U11689 (N_11689,N_7780,N_6176);
or U11690 (N_11690,N_8807,N_8323);
nor U11691 (N_11691,N_7453,N_6240);
and U11692 (N_11692,N_8257,N_6199);
nor U11693 (N_11693,N_6177,N_6064);
and U11694 (N_11694,N_7318,N_6296);
or U11695 (N_11695,N_8564,N_7061);
xor U11696 (N_11696,N_8511,N_6370);
nor U11697 (N_11697,N_8776,N_7541);
and U11698 (N_11698,N_6582,N_7282);
nor U11699 (N_11699,N_8916,N_6480);
and U11700 (N_11700,N_6534,N_6866);
or U11701 (N_11701,N_6356,N_7765);
or U11702 (N_11702,N_6615,N_6944);
or U11703 (N_11703,N_6995,N_8370);
nor U11704 (N_11704,N_6459,N_7602);
or U11705 (N_11705,N_7072,N_7999);
and U11706 (N_11706,N_8078,N_6494);
or U11707 (N_11707,N_8486,N_6820);
and U11708 (N_11708,N_8688,N_8008);
nor U11709 (N_11709,N_6296,N_8262);
nand U11710 (N_11710,N_8545,N_8008);
nand U11711 (N_11711,N_7318,N_7419);
and U11712 (N_11712,N_8430,N_8962);
and U11713 (N_11713,N_6747,N_8820);
and U11714 (N_11714,N_8249,N_6432);
or U11715 (N_11715,N_8060,N_7188);
nand U11716 (N_11716,N_7915,N_8846);
or U11717 (N_11717,N_6037,N_8623);
nand U11718 (N_11718,N_6680,N_8581);
and U11719 (N_11719,N_7580,N_8437);
and U11720 (N_11720,N_8975,N_7809);
and U11721 (N_11721,N_8369,N_6186);
or U11722 (N_11722,N_6119,N_8631);
nand U11723 (N_11723,N_7599,N_8182);
and U11724 (N_11724,N_7250,N_7306);
xnor U11725 (N_11725,N_6321,N_6368);
and U11726 (N_11726,N_6253,N_8601);
nand U11727 (N_11727,N_7071,N_7068);
or U11728 (N_11728,N_6656,N_8636);
nor U11729 (N_11729,N_6532,N_6436);
or U11730 (N_11730,N_7248,N_6052);
nand U11731 (N_11731,N_8717,N_7373);
nand U11732 (N_11732,N_8438,N_7775);
or U11733 (N_11733,N_7366,N_6920);
or U11734 (N_11734,N_6315,N_7843);
nor U11735 (N_11735,N_8473,N_6779);
nor U11736 (N_11736,N_6442,N_6206);
or U11737 (N_11737,N_8531,N_8578);
or U11738 (N_11738,N_8740,N_8922);
or U11739 (N_11739,N_8087,N_6003);
and U11740 (N_11740,N_7105,N_7216);
nor U11741 (N_11741,N_6051,N_8805);
and U11742 (N_11742,N_7310,N_7386);
nor U11743 (N_11743,N_7942,N_6513);
nand U11744 (N_11744,N_6282,N_7466);
nand U11745 (N_11745,N_7088,N_6781);
and U11746 (N_11746,N_8408,N_8868);
or U11747 (N_11747,N_8392,N_7161);
or U11748 (N_11748,N_8548,N_8921);
and U11749 (N_11749,N_7873,N_6772);
or U11750 (N_11750,N_8003,N_7831);
nand U11751 (N_11751,N_8426,N_8394);
or U11752 (N_11752,N_6462,N_6267);
nor U11753 (N_11753,N_6667,N_7207);
nor U11754 (N_11754,N_8386,N_7006);
nand U11755 (N_11755,N_7876,N_8928);
nand U11756 (N_11756,N_6990,N_6556);
nor U11757 (N_11757,N_6821,N_8420);
or U11758 (N_11758,N_6236,N_6092);
nor U11759 (N_11759,N_8567,N_7655);
nor U11760 (N_11760,N_6162,N_7280);
or U11761 (N_11761,N_7217,N_8767);
nand U11762 (N_11762,N_8442,N_8129);
nor U11763 (N_11763,N_7730,N_7783);
nor U11764 (N_11764,N_8045,N_8296);
nand U11765 (N_11765,N_7014,N_7351);
nand U11766 (N_11766,N_8332,N_8854);
xnor U11767 (N_11767,N_6696,N_7898);
and U11768 (N_11768,N_8172,N_6578);
and U11769 (N_11769,N_8617,N_8886);
nor U11770 (N_11770,N_7526,N_8533);
or U11771 (N_11771,N_7889,N_8861);
nor U11772 (N_11772,N_7166,N_6332);
or U11773 (N_11773,N_6221,N_7677);
nand U11774 (N_11774,N_6811,N_7389);
or U11775 (N_11775,N_6104,N_8016);
or U11776 (N_11776,N_6764,N_6223);
and U11777 (N_11777,N_8407,N_8563);
or U11778 (N_11778,N_6959,N_6275);
nand U11779 (N_11779,N_8944,N_6939);
nand U11780 (N_11780,N_8318,N_6109);
and U11781 (N_11781,N_7012,N_7981);
and U11782 (N_11782,N_7696,N_8860);
nor U11783 (N_11783,N_8469,N_7350);
and U11784 (N_11784,N_7061,N_8355);
and U11785 (N_11785,N_8146,N_6712);
or U11786 (N_11786,N_7546,N_8871);
nand U11787 (N_11787,N_7996,N_7474);
or U11788 (N_11788,N_8268,N_6554);
and U11789 (N_11789,N_8561,N_8650);
nand U11790 (N_11790,N_7976,N_6986);
nand U11791 (N_11791,N_8715,N_6983);
nor U11792 (N_11792,N_6976,N_7919);
nand U11793 (N_11793,N_8015,N_7332);
nand U11794 (N_11794,N_8268,N_7749);
nor U11795 (N_11795,N_6912,N_6844);
and U11796 (N_11796,N_8393,N_7918);
and U11797 (N_11797,N_7500,N_7203);
and U11798 (N_11798,N_7995,N_8050);
and U11799 (N_11799,N_6152,N_6436);
or U11800 (N_11800,N_7386,N_7907);
and U11801 (N_11801,N_8303,N_6625);
and U11802 (N_11802,N_6608,N_8749);
and U11803 (N_11803,N_8319,N_6789);
nor U11804 (N_11804,N_6824,N_6882);
nor U11805 (N_11805,N_6434,N_8269);
and U11806 (N_11806,N_7885,N_8470);
nor U11807 (N_11807,N_8693,N_8120);
xor U11808 (N_11808,N_7447,N_7271);
and U11809 (N_11809,N_7766,N_8791);
or U11810 (N_11810,N_6469,N_8139);
or U11811 (N_11811,N_7868,N_8672);
and U11812 (N_11812,N_6693,N_8639);
nand U11813 (N_11813,N_7931,N_7003);
nor U11814 (N_11814,N_7570,N_6898);
xor U11815 (N_11815,N_8994,N_6877);
nor U11816 (N_11816,N_6845,N_8610);
nor U11817 (N_11817,N_6440,N_6645);
nand U11818 (N_11818,N_8537,N_8358);
and U11819 (N_11819,N_7296,N_8096);
nand U11820 (N_11820,N_8530,N_8188);
or U11821 (N_11821,N_6209,N_7622);
and U11822 (N_11822,N_6406,N_8597);
nor U11823 (N_11823,N_8993,N_6426);
or U11824 (N_11824,N_7527,N_6972);
and U11825 (N_11825,N_8288,N_8337);
and U11826 (N_11826,N_6455,N_7019);
nor U11827 (N_11827,N_6990,N_8182);
nor U11828 (N_11828,N_7990,N_8499);
or U11829 (N_11829,N_7179,N_8793);
and U11830 (N_11830,N_7697,N_6180);
and U11831 (N_11831,N_6119,N_8250);
and U11832 (N_11832,N_6770,N_6768);
or U11833 (N_11833,N_8020,N_8328);
and U11834 (N_11834,N_8482,N_7438);
and U11835 (N_11835,N_6278,N_7513);
nor U11836 (N_11836,N_8696,N_6879);
xnor U11837 (N_11837,N_8385,N_6465);
or U11838 (N_11838,N_7923,N_6168);
or U11839 (N_11839,N_7206,N_8582);
or U11840 (N_11840,N_8140,N_7946);
and U11841 (N_11841,N_8943,N_6386);
nand U11842 (N_11842,N_7719,N_7543);
and U11843 (N_11843,N_6661,N_6462);
or U11844 (N_11844,N_7669,N_8944);
and U11845 (N_11845,N_8536,N_7359);
nor U11846 (N_11846,N_8322,N_8415);
or U11847 (N_11847,N_7003,N_7766);
nand U11848 (N_11848,N_6582,N_8641);
and U11849 (N_11849,N_7551,N_7495);
nand U11850 (N_11850,N_7344,N_8739);
nand U11851 (N_11851,N_8378,N_6204);
nor U11852 (N_11852,N_6385,N_7869);
nor U11853 (N_11853,N_6782,N_6115);
nand U11854 (N_11854,N_6329,N_8022);
nand U11855 (N_11855,N_8635,N_8959);
or U11856 (N_11856,N_7554,N_8418);
or U11857 (N_11857,N_6986,N_7407);
or U11858 (N_11858,N_6330,N_8291);
or U11859 (N_11859,N_7408,N_7968);
nor U11860 (N_11860,N_7936,N_6320);
and U11861 (N_11861,N_7679,N_7452);
and U11862 (N_11862,N_8684,N_8732);
or U11863 (N_11863,N_8012,N_7301);
or U11864 (N_11864,N_6043,N_8760);
nand U11865 (N_11865,N_8699,N_7100);
xor U11866 (N_11866,N_6874,N_6646);
and U11867 (N_11867,N_8661,N_7875);
or U11868 (N_11868,N_7517,N_8414);
or U11869 (N_11869,N_7866,N_8347);
or U11870 (N_11870,N_7075,N_8362);
and U11871 (N_11871,N_7230,N_8399);
nor U11872 (N_11872,N_8058,N_7191);
nor U11873 (N_11873,N_7929,N_7856);
and U11874 (N_11874,N_8692,N_8829);
nand U11875 (N_11875,N_7172,N_7152);
nor U11876 (N_11876,N_6478,N_8691);
or U11877 (N_11877,N_6199,N_8166);
nand U11878 (N_11878,N_8070,N_6979);
and U11879 (N_11879,N_7394,N_6010);
and U11880 (N_11880,N_6772,N_8715);
and U11881 (N_11881,N_6429,N_7331);
nor U11882 (N_11882,N_6314,N_7510);
nand U11883 (N_11883,N_8000,N_6095);
and U11884 (N_11884,N_8170,N_6599);
and U11885 (N_11885,N_7089,N_7911);
nor U11886 (N_11886,N_6245,N_8234);
nor U11887 (N_11887,N_7446,N_6483);
or U11888 (N_11888,N_6504,N_6730);
and U11889 (N_11889,N_6529,N_7266);
nand U11890 (N_11890,N_6872,N_8850);
nor U11891 (N_11891,N_6900,N_8985);
or U11892 (N_11892,N_6000,N_7201);
nand U11893 (N_11893,N_8275,N_7353);
nand U11894 (N_11894,N_6892,N_6798);
and U11895 (N_11895,N_6354,N_6006);
nand U11896 (N_11896,N_7046,N_8451);
nand U11897 (N_11897,N_8820,N_6746);
or U11898 (N_11898,N_7871,N_8275);
nor U11899 (N_11899,N_7506,N_6548);
and U11900 (N_11900,N_7616,N_6815);
nand U11901 (N_11901,N_8377,N_6689);
or U11902 (N_11902,N_8464,N_7466);
nor U11903 (N_11903,N_6786,N_7498);
nand U11904 (N_11904,N_8955,N_6650);
or U11905 (N_11905,N_6871,N_6513);
nand U11906 (N_11906,N_8846,N_7710);
and U11907 (N_11907,N_8517,N_8601);
nand U11908 (N_11908,N_7303,N_6495);
or U11909 (N_11909,N_7697,N_8561);
and U11910 (N_11910,N_6511,N_8513);
nor U11911 (N_11911,N_6820,N_7408);
nor U11912 (N_11912,N_6092,N_7155);
and U11913 (N_11913,N_7657,N_7819);
nor U11914 (N_11914,N_6521,N_6646);
nor U11915 (N_11915,N_8717,N_6142);
nor U11916 (N_11916,N_6655,N_6114);
and U11917 (N_11917,N_8338,N_6434);
nor U11918 (N_11918,N_7670,N_8016);
nor U11919 (N_11919,N_6072,N_6364);
nor U11920 (N_11920,N_7297,N_8436);
nor U11921 (N_11921,N_8532,N_6820);
or U11922 (N_11922,N_7996,N_8708);
nand U11923 (N_11923,N_8832,N_6027);
nand U11924 (N_11924,N_7877,N_8211);
nand U11925 (N_11925,N_8887,N_7092);
nor U11926 (N_11926,N_7761,N_7998);
nand U11927 (N_11927,N_7892,N_8329);
or U11928 (N_11928,N_8059,N_7112);
or U11929 (N_11929,N_8407,N_6122);
nand U11930 (N_11930,N_8345,N_6811);
or U11931 (N_11931,N_6509,N_7564);
nand U11932 (N_11932,N_6526,N_6279);
nor U11933 (N_11933,N_7261,N_8302);
and U11934 (N_11934,N_6824,N_6311);
and U11935 (N_11935,N_8940,N_6706);
or U11936 (N_11936,N_8526,N_6844);
xor U11937 (N_11937,N_7751,N_7571);
and U11938 (N_11938,N_8827,N_7959);
nand U11939 (N_11939,N_8145,N_8050);
nor U11940 (N_11940,N_6193,N_8674);
or U11941 (N_11941,N_7538,N_7406);
nor U11942 (N_11942,N_7015,N_6421);
nor U11943 (N_11943,N_7200,N_7500);
nor U11944 (N_11944,N_8049,N_7386);
nor U11945 (N_11945,N_7126,N_8836);
nand U11946 (N_11946,N_6779,N_8574);
and U11947 (N_11947,N_6823,N_7241);
or U11948 (N_11948,N_7713,N_8282);
and U11949 (N_11949,N_7767,N_6085);
nor U11950 (N_11950,N_8878,N_8643);
and U11951 (N_11951,N_6335,N_8189);
or U11952 (N_11952,N_7331,N_8600);
nor U11953 (N_11953,N_8773,N_7882);
nand U11954 (N_11954,N_7536,N_8617);
and U11955 (N_11955,N_7421,N_8553);
xnor U11956 (N_11956,N_6646,N_7424);
or U11957 (N_11957,N_7715,N_6957);
or U11958 (N_11958,N_8069,N_6147);
or U11959 (N_11959,N_6328,N_6533);
and U11960 (N_11960,N_8672,N_6862);
nor U11961 (N_11961,N_8477,N_7290);
nor U11962 (N_11962,N_6379,N_7220);
or U11963 (N_11963,N_7235,N_6435);
nand U11964 (N_11964,N_6756,N_6903);
and U11965 (N_11965,N_7148,N_7572);
and U11966 (N_11966,N_7499,N_8923);
nand U11967 (N_11967,N_8901,N_7859);
nand U11968 (N_11968,N_8821,N_6963);
and U11969 (N_11969,N_8625,N_7417);
xnor U11970 (N_11970,N_7651,N_7618);
or U11971 (N_11971,N_7115,N_7027);
or U11972 (N_11972,N_8559,N_6858);
and U11973 (N_11973,N_8614,N_7719);
or U11974 (N_11974,N_7245,N_6307);
nor U11975 (N_11975,N_7342,N_6482);
or U11976 (N_11976,N_7220,N_6293);
and U11977 (N_11977,N_7620,N_7785);
or U11978 (N_11978,N_6681,N_6631);
nor U11979 (N_11979,N_7860,N_6686);
or U11980 (N_11980,N_7270,N_8953);
or U11981 (N_11981,N_7379,N_7946);
nor U11982 (N_11982,N_7694,N_8880);
nor U11983 (N_11983,N_6913,N_6084);
nand U11984 (N_11984,N_8497,N_7778);
and U11985 (N_11985,N_7907,N_7523);
and U11986 (N_11986,N_8807,N_6787);
or U11987 (N_11987,N_7673,N_7260);
nand U11988 (N_11988,N_7245,N_6506);
nand U11989 (N_11989,N_7217,N_7767);
nor U11990 (N_11990,N_6816,N_8757);
nand U11991 (N_11991,N_6054,N_7281);
nor U11992 (N_11992,N_8580,N_7250);
nor U11993 (N_11993,N_7022,N_6797);
or U11994 (N_11994,N_7577,N_6065);
and U11995 (N_11995,N_6995,N_8859);
or U11996 (N_11996,N_6642,N_8762);
or U11997 (N_11997,N_8500,N_7883);
and U11998 (N_11998,N_7232,N_6519);
nand U11999 (N_11999,N_6598,N_7086);
or U12000 (N_12000,N_9762,N_10851);
nor U12001 (N_12001,N_11064,N_9318);
nand U12002 (N_12002,N_11596,N_9114);
nand U12003 (N_12003,N_11438,N_11855);
nor U12004 (N_12004,N_9194,N_10526);
nand U12005 (N_12005,N_11789,N_10675);
and U12006 (N_12006,N_11829,N_9814);
nand U12007 (N_12007,N_11737,N_11535);
nor U12008 (N_12008,N_9604,N_10177);
nand U12009 (N_12009,N_11575,N_10844);
nor U12010 (N_12010,N_9475,N_9163);
or U12011 (N_12011,N_10965,N_10218);
and U12012 (N_12012,N_10959,N_9880);
nand U12013 (N_12013,N_11477,N_10673);
or U12014 (N_12014,N_11331,N_10827);
nor U12015 (N_12015,N_9268,N_9101);
nor U12016 (N_12016,N_10100,N_9132);
and U12017 (N_12017,N_10627,N_10683);
or U12018 (N_12018,N_9892,N_11788);
and U12019 (N_12019,N_9579,N_10752);
nor U12020 (N_12020,N_11715,N_10832);
xor U12021 (N_12021,N_10754,N_9255);
nor U12022 (N_12022,N_9742,N_11927);
or U12023 (N_12023,N_11791,N_11419);
or U12024 (N_12024,N_11548,N_10693);
nand U12025 (N_12025,N_9747,N_10369);
nand U12026 (N_12026,N_11595,N_11199);
nand U12027 (N_12027,N_11197,N_11570);
or U12028 (N_12028,N_9083,N_11490);
nand U12029 (N_12029,N_11882,N_11917);
nor U12030 (N_12030,N_10976,N_10839);
nor U12031 (N_12031,N_10488,N_11301);
nand U12032 (N_12032,N_9497,N_10637);
nor U12033 (N_12033,N_10953,N_11128);
and U12034 (N_12034,N_9055,N_10642);
and U12035 (N_12035,N_11978,N_11183);
and U12036 (N_12036,N_9175,N_11192);
and U12037 (N_12037,N_11292,N_10812);
nor U12038 (N_12038,N_10424,N_11452);
nor U12039 (N_12039,N_9238,N_10698);
or U12040 (N_12040,N_10457,N_9458);
or U12041 (N_12041,N_9613,N_9451);
nor U12042 (N_12042,N_11985,N_9694);
or U12043 (N_12043,N_9011,N_11445);
nor U12044 (N_12044,N_10681,N_9303);
or U12045 (N_12045,N_10934,N_9938);
and U12046 (N_12046,N_11956,N_10875);
and U12047 (N_12047,N_11071,N_10454);
and U12048 (N_12048,N_10774,N_10896);
or U12049 (N_12049,N_9206,N_9187);
nand U12050 (N_12050,N_11954,N_9663);
or U12051 (N_12051,N_10075,N_10977);
nor U12052 (N_12052,N_10757,N_9772);
and U12053 (N_12053,N_9510,N_11053);
nor U12054 (N_12054,N_9505,N_10746);
nor U12055 (N_12055,N_11514,N_9671);
and U12056 (N_12056,N_10301,N_9700);
and U12057 (N_12057,N_10196,N_9727);
nor U12058 (N_12058,N_11965,N_11754);
nand U12059 (N_12059,N_9855,N_10336);
or U12060 (N_12060,N_10314,N_10141);
nor U12061 (N_12061,N_9617,N_9491);
nor U12062 (N_12062,N_11902,N_9020);
and U12063 (N_12063,N_9724,N_10522);
nand U12064 (N_12064,N_9217,N_9974);
and U12065 (N_12065,N_11177,N_10281);
or U12066 (N_12066,N_9788,N_9627);
or U12067 (N_12067,N_10884,N_9254);
or U12068 (N_12068,N_11214,N_10227);
nand U12069 (N_12069,N_11929,N_10157);
and U12070 (N_12070,N_9882,N_11337);
and U12071 (N_12071,N_9684,N_10855);
nor U12072 (N_12072,N_9036,N_10840);
and U12073 (N_12073,N_10663,N_9328);
or U12074 (N_12074,N_11534,N_11850);
nand U12075 (N_12075,N_11624,N_10067);
and U12076 (N_12076,N_10188,N_10463);
nor U12077 (N_12077,N_9369,N_10047);
nand U12078 (N_12078,N_10327,N_9988);
and U12079 (N_12079,N_10872,N_10871);
nor U12080 (N_12080,N_11690,N_10018);
nor U12081 (N_12081,N_11792,N_10242);
nand U12082 (N_12082,N_11826,N_11479);
or U12083 (N_12083,N_10544,N_9917);
and U12084 (N_12084,N_10362,N_10672);
or U12085 (N_12085,N_10927,N_9162);
nor U12086 (N_12086,N_10116,N_11330);
nor U12087 (N_12087,N_10012,N_10248);
and U12088 (N_12088,N_10946,N_11253);
or U12089 (N_12089,N_11079,N_11375);
xor U12090 (N_12090,N_11924,N_10226);
or U12091 (N_12091,N_11151,N_9498);
nand U12092 (N_12092,N_10980,N_9360);
or U12093 (N_12093,N_9168,N_10858);
nor U12094 (N_12094,N_9751,N_9079);
or U12095 (N_12095,N_11734,N_11097);
nor U12096 (N_12096,N_9801,N_9234);
and U12097 (N_12097,N_10269,N_9810);
or U12098 (N_12098,N_10000,N_10169);
or U12099 (N_12099,N_11576,N_11951);
nand U12100 (N_12100,N_9553,N_11092);
nand U12101 (N_12101,N_11244,N_9013);
nor U12102 (N_12102,N_11362,N_11102);
nand U12103 (N_12103,N_11091,N_9651);
and U12104 (N_12104,N_9999,N_11594);
or U12105 (N_12105,N_9316,N_10077);
nand U12106 (N_12106,N_9593,N_11047);
xnor U12107 (N_12107,N_9874,N_11138);
or U12108 (N_12108,N_9386,N_11294);
and U12109 (N_12109,N_9569,N_11308);
nand U12110 (N_12110,N_10236,N_10056);
or U12111 (N_12111,N_10793,N_11495);
or U12112 (N_12112,N_9464,N_9240);
nor U12113 (N_12113,N_10559,N_11153);
nand U12114 (N_12114,N_11778,N_10496);
nand U12115 (N_12115,N_11557,N_10966);
nor U12116 (N_12116,N_10250,N_10365);
and U12117 (N_12117,N_9448,N_10553);
nor U12118 (N_12118,N_10868,N_10937);
nand U12119 (N_12119,N_10049,N_11824);
nand U12120 (N_12120,N_10631,N_9518);
nand U12121 (N_12121,N_10228,N_10005);
nand U12122 (N_12122,N_10703,N_10968);
and U12123 (N_12123,N_10473,N_10278);
nor U12124 (N_12124,N_9203,N_10607);
or U12125 (N_12125,N_9930,N_11974);
nand U12126 (N_12126,N_10195,N_9023);
or U12127 (N_12127,N_11195,N_11061);
and U12128 (N_12128,N_10468,N_10450);
nor U12129 (N_12129,N_11806,N_9567);
nor U12130 (N_12130,N_9753,N_9073);
nand U12131 (N_12131,N_10520,N_9461);
and U12132 (N_12132,N_11204,N_10514);
and U12133 (N_12133,N_9302,N_11469);
and U12134 (N_12134,N_11234,N_9147);
nand U12135 (N_12135,N_10412,N_10733);
nand U12136 (N_12136,N_10864,N_9872);
nand U12137 (N_12137,N_11921,N_9247);
nor U12138 (N_12138,N_10493,N_10790);
or U12139 (N_12139,N_11519,N_9253);
nand U12140 (N_12140,N_11649,N_10474);
and U12141 (N_12141,N_11720,N_11843);
nor U12142 (N_12142,N_10178,N_10736);
nor U12143 (N_12143,N_9285,N_10458);
nand U12144 (N_12144,N_11232,N_11820);
and U12145 (N_12145,N_11878,N_11193);
or U12146 (N_12146,N_11381,N_9289);
nand U12147 (N_12147,N_10778,N_11009);
or U12148 (N_12148,N_9967,N_10765);
nor U12149 (N_12149,N_9306,N_10616);
nand U12150 (N_12150,N_9152,N_10716);
and U12151 (N_12151,N_9260,N_10209);
nor U12152 (N_12152,N_10099,N_11545);
or U12153 (N_12153,N_11074,N_9249);
nand U12154 (N_12154,N_11834,N_10411);
and U12155 (N_12155,N_10926,N_10013);
nor U12156 (N_12156,N_11486,N_10601);
or U12157 (N_12157,N_11285,N_9725);
and U12158 (N_12158,N_9525,N_9923);
nor U12159 (N_12159,N_11683,N_9915);
or U12160 (N_12160,N_9324,N_9982);
nand U12161 (N_12161,N_11196,N_11320);
xor U12162 (N_12162,N_10329,N_10655);
and U12163 (N_12163,N_11746,N_9941);
nand U12164 (N_12164,N_10330,N_10262);
nand U12165 (N_12165,N_9435,N_11623);
and U12166 (N_12166,N_9117,N_9668);
nor U12167 (N_12167,N_11708,N_11868);
and U12168 (N_12168,N_10780,N_11993);
or U12169 (N_12169,N_10221,N_11571);
nand U12170 (N_12170,N_11742,N_11260);
and U12171 (N_12171,N_10154,N_11706);
nor U12172 (N_12172,N_9598,N_11520);
nor U12173 (N_12173,N_10313,N_9232);
nor U12174 (N_12174,N_10619,N_9825);
nand U12175 (N_12175,N_10785,N_10867);
and U12176 (N_12176,N_11202,N_11466);
nor U12177 (N_12177,N_10094,N_11815);
nand U12178 (N_12178,N_9108,N_9947);
or U12179 (N_12179,N_9250,N_9992);
nand U12180 (N_12180,N_11861,N_11240);
and U12181 (N_12181,N_9068,N_11989);
nand U12182 (N_12182,N_10279,N_10521);
and U12183 (N_12183,N_9913,N_9638);
and U12184 (N_12184,N_11547,N_9533);
or U12185 (N_12185,N_9682,N_11089);
or U12186 (N_12186,N_10376,N_11421);
and U12187 (N_12187,N_10605,N_10433);
and U12188 (N_12188,N_11030,N_11586);
nor U12189 (N_12189,N_11425,N_9688);
or U12190 (N_12190,N_9105,N_10095);
or U12191 (N_12191,N_9916,N_10555);
nand U12192 (N_12192,N_9080,N_11664);
nand U12193 (N_12193,N_10027,N_9634);
or U12194 (N_12194,N_9978,N_10986);
nand U12195 (N_12195,N_11562,N_9970);
nand U12196 (N_12196,N_11341,N_10658);
nor U12197 (N_12197,N_9259,N_10728);
and U12198 (N_12198,N_10015,N_9502);
nor U12199 (N_12199,N_10888,N_10023);
nand U12200 (N_12200,N_11536,N_10264);
and U12201 (N_12201,N_11748,N_11357);
nor U12202 (N_12202,N_11002,N_11284);
or U12203 (N_12203,N_11710,N_10661);
and U12204 (N_12204,N_11396,N_9170);
or U12205 (N_12205,N_11465,N_10233);
nor U12206 (N_12206,N_10384,N_10291);
nor U12207 (N_12207,N_10261,N_9675);
nand U12208 (N_12208,N_11581,N_9805);
or U12209 (N_12209,N_9102,N_9844);
nand U12210 (N_12210,N_9368,N_11532);
or U12211 (N_12211,N_10639,N_9831);
nand U12212 (N_12212,N_9580,N_11609);
or U12213 (N_12213,N_10951,N_11981);
nand U12214 (N_12214,N_11654,N_10659);
or U12215 (N_12215,N_10779,N_10448);
nand U12216 (N_12216,N_10371,N_10210);
and U12217 (N_12217,N_9099,N_9439);
nor U12218 (N_12218,N_10597,N_11145);
or U12219 (N_12219,N_10708,N_9798);
nand U12220 (N_12220,N_9802,N_11027);
nor U12221 (N_12221,N_11884,N_10536);
nand U12222 (N_12222,N_9721,N_11923);
nand U12223 (N_12223,N_9057,N_10540);
and U12224 (N_12224,N_10964,N_11697);
nor U12225 (N_12225,N_10957,N_11444);
nand U12226 (N_12226,N_10660,N_9574);
nor U12227 (N_12227,N_9066,N_10272);
nor U12228 (N_12228,N_11173,N_11448);
or U12229 (N_12229,N_9791,N_9568);
nand U12230 (N_12230,N_9779,N_10442);
nand U12231 (N_12231,N_9050,N_10328);
and U12232 (N_12232,N_10092,N_11961);
and U12233 (N_12233,N_11267,N_11579);
or U12234 (N_12234,N_10344,N_9002);
or U12235 (N_12235,N_10907,N_9446);
and U12236 (N_12236,N_10600,N_10182);
and U12237 (N_12237,N_10789,N_10428);
nand U12238 (N_12238,N_10014,N_10909);
nor U12239 (N_12239,N_9756,N_10970);
nor U12240 (N_12240,N_9927,N_10837);
nor U12241 (N_12241,N_11109,N_11691);
nor U12242 (N_12242,N_10685,N_9883);
nand U12243 (N_12243,N_9933,N_11982);
nand U12244 (N_12244,N_11123,N_10691);
or U12245 (N_12245,N_9975,N_11502);
and U12246 (N_12246,N_11704,N_11328);
or U12247 (N_12247,N_10383,N_9431);
or U12248 (N_12248,N_11758,N_9596);
or U12249 (N_12249,N_9618,N_9354);
xor U12250 (N_12250,N_10657,N_10158);
nor U12251 (N_12251,N_11271,N_10721);
nor U12252 (N_12252,N_11573,N_10594);
xor U12253 (N_12253,N_9048,N_11959);
or U12254 (N_12254,N_9224,N_9884);
nand U12255 (N_12255,N_10198,N_11297);
nand U12256 (N_12256,N_11043,N_10944);
nor U12257 (N_12257,N_10375,N_9331);
nand U12258 (N_12258,N_11431,N_11887);
and U12259 (N_12259,N_9655,N_9806);
nand U12260 (N_12260,N_9961,N_11401);
xor U12261 (N_12261,N_10398,N_9936);
and U12262 (N_12262,N_10849,N_11756);
or U12263 (N_12263,N_10595,N_10997);
nand U12264 (N_12264,N_9847,N_10469);
nand U12265 (N_12265,N_9739,N_11101);
or U12266 (N_12266,N_10205,N_10820);
and U12267 (N_12267,N_11616,N_9078);
nor U12268 (N_12268,N_11120,N_11058);
or U12269 (N_12269,N_11456,N_9873);
nand U12270 (N_12270,N_9144,N_9284);
or U12271 (N_12271,N_10300,N_9662);
or U12272 (N_12272,N_11392,N_9846);
nand U12273 (N_12273,N_10282,N_9134);
or U12274 (N_12274,N_11430,N_11026);
and U12275 (N_12275,N_9001,N_10679);
or U12276 (N_12276,N_9614,N_10400);
or U12277 (N_12277,N_9922,N_10317);
nor U12278 (N_12278,N_9047,N_10443);
and U12279 (N_12279,N_10294,N_11871);
or U12280 (N_12280,N_11941,N_10768);
nor U12281 (N_12281,N_10308,N_10471);
and U12282 (N_12282,N_9524,N_10394);
and U12283 (N_12283,N_10397,N_11363);
nor U12284 (N_12284,N_9706,N_10666);
and U12285 (N_12285,N_11937,N_11345);
nand U12286 (N_12286,N_9130,N_11672);
and U12287 (N_12287,N_11158,N_9543);
or U12288 (N_12288,N_11447,N_10366);
or U12289 (N_12289,N_9030,N_9071);
or U12290 (N_12290,N_9243,N_10819);
or U12291 (N_12291,N_11491,N_10713);
or U12292 (N_12292,N_9755,N_10273);
or U12293 (N_12293,N_9490,N_10569);
and U12294 (N_12294,N_9636,N_9990);
and U12295 (N_12295,N_11650,N_9319);
nor U12296 (N_12296,N_10485,N_9904);
and U12297 (N_12297,N_10583,N_10147);
and U12298 (N_12298,N_11633,N_11618);
and U12299 (N_12299,N_9501,N_10602);
nand U12300 (N_12300,N_9834,N_10709);
nor U12301 (N_12301,N_10423,N_9186);
and U12302 (N_12302,N_11528,N_9022);
and U12303 (N_12303,N_9179,N_10061);
and U12304 (N_12304,N_11783,N_9353);
nand U12305 (N_12305,N_9167,N_9345);
nor U12306 (N_12306,N_10073,N_11740);
and U12307 (N_12307,N_11095,N_11004);
or U12308 (N_12308,N_11118,N_10197);
nand U12309 (N_12309,N_11877,N_9852);
nor U12310 (N_12310,N_11793,N_11743);
nand U12311 (N_12311,N_9287,N_11728);
or U12312 (N_12312,N_11449,N_9746);
nor U12313 (N_12313,N_9777,N_11684);
and U12314 (N_12314,N_10303,N_11296);
and U12315 (N_12315,N_9212,N_11760);
or U12316 (N_12316,N_10504,N_11327);
nor U12317 (N_12317,N_10413,N_11156);
or U12318 (N_12318,N_10382,N_9723);
or U12319 (N_12319,N_9423,N_11358);
or U12320 (N_12320,N_11821,N_9198);
and U12321 (N_12321,N_10935,N_10761);
nor U12322 (N_12322,N_10647,N_10582);
nor U12323 (N_12323,N_10035,N_10542);
or U12324 (N_12324,N_11913,N_9375);
nand U12325 (N_12325,N_9304,N_9886);
nor U12326 (N_12326,N_10089,N_10948);
and U12327 (N_12327,N_10750,N_10356);
nor U12328 (N_12328,N_11673,N_11588);
or U12329 (N_12329,N_10432,N_9157);
nand U12330 (N_12330,N_11818,N_9716);
or U12331 (N_12331,N_11011,N_10741);
nand U12332 (N_12332,N_9561,N_9955);
or U12333 (N_12333,N_11352,N_10247);
and U12334 (N_12334,N_10760,N_10950);
nand U12335 (N_12335,N_10472,N_9398);
and U12336 (N_12336,N_11224,N_11852);
and U12337 (N_12337,N_11897,N_10155);
and U12338 (N_12338,N_9330,N_11918);
or U12339 (N_12339,N_10203,N_11418);
nand U12340 (N_12340,N_10490,N_11797);
or U12341 (N_12341,N_11745,N_9093);
nand U12342 (N_12342,N_11104,N_10123);
or U12343 (N_12343,N_10387,N_9493);
and U12344 (N_12344,N_11607,N_11784);
and U12345 (N_12345,N_9028,N_10500);
nand U12346 (N_12346,N_9665,N_10083);
nor U12347 (N_12347,N_9400,N_10910);
or U12348 (N_12348,N_10088,N_11134);
and U12349 (N_12349,N_11459,N_9529);
nand U12350 (N_12350,N_11409,N_9744);
and U12351 (N_12351,N_10380,N_10845);
or U12352 (N_12352,N_11919,N_9571);
or U12353 (N_12353,N_11346,N_10924);
nand U12354 (N_12354,N_11835,N_9476);
nor U12355 (N_12355,N_11597,N_11473);
nand U12356 (N_12356,N_10190,N_11147);
nand U12357 (N_12357,N_11638,N_10091);
nand U12358 (N_12358,N_9632,N_9804);
nand U12359 (N_12359,N_11901,N_11050);
and U12360 (N_12360,N_11786,N_11731);
nand U12361 (N_12361,N_9348,N_9090);
or U12362 (N_12362,N_10406,N_9843);
and U12363 (N_12363,N_11537,N_10148);
nor U12364 (N_12364,N_11798,N_10710);
and U12365 (N_12365,N_10925,N_9086);
nor U12366 (N_12366,N_11667,N_9519);
or U12367 (N_12367,N_11216,N_10489);
and U12368 (N_12368,N_11239,N_9729);
and U12369 (N_12369,N_10696,N_9278);
and U12370 (N_12370,N_11540,N_10363);
nor U12371 (N_12371,N_11119,N_10447);
nor U12372 (N_12372,N_9358,N_11274);
nand U12373 (N_12373,N_11481,N_9550);
nand U12374 (N_12374,N_10286,N_9311);
nand U12375 (N_12375,N_9044,N_9708);
and U12376 (N_12376,N_9542,N_11254);
and U12377 (N_12377,N_10256,N_9236);
and U12378 (N_12378,N_10813,N_9293);
and U12379 (N_12379,N_9600,N_10360);
or U12380 (N_12380,N_9312,N_10802);
nor U12381 (N_12381,N_11242,N_10921);
nor U12382 (N_12382,N_10905,N_10004);
and U12383 (N_12383,N_9956,N_11642);
or U12384 (N_12384,N_9678,N_9893);
nand U12385 (N_12385,N_9004,N_11437);
or U12386 (N_12386,N_10404,N_11413);
nor U12387 (N_12387,N_11154,N_11659);
and U12388 (N_12388,N_9887,N_9760);
and U12389 (N_12389,N_9648,N_9784);
nor U12390 (N_12390,N_9637,N_9546);
and U12391 (N_12391,N_9709,N_10331);
or U12392 (N_12392,N_11155,N_11827);
nor U12393 (N_12393,N_9996,N_10632);
and U12394 (N_12394,N_9213,N_10873);
and U12395 (N_12395,N_9943,N_9871);
nand U12396 (N_12396,N_11550,N_11805);
nor U12397 (N_12397,N_10348,N_9558);
and U12398 (N_12398,N_10146,N_9181);
nand U12399 (N_12399,N_9365,N_11839);
nand U12400 (N_12400,N_11893,N_11368);
and U12401 (N_12401,N_11142,N_11257);
and U12402 (N_12402,N_9095,N_9372);
and U12403 (N_12403,N_9926,N_9677);
nand U12404 (N_12404,N_10150,N_11360);
and U12405 (N_12405,N_9667,N_9738);
or U12406 (N_12406,N_11217,N_11457);
or U12407 (N_12407,N_11367,N_9585);
nand U12408 (N_12408,N_9195,N_9067);
nand U12409 (N_12409,N_9087,N_9531);
nor U12410 (N_12410,N_10343,N_10243);
nor U12411 (N_12411,N_10829,N_11181);
and U12412 (N_12412,N_10641,N_10949);
nor U12413 (N_12413,N_11630,N_11212);
nand U12414 (N_12414,N_10296,N_10168);
nor U12415 (N_12415,N_10044,N_10347);
and U12416 (N_12416,N_10487,N_9998);
and U12417 (N_12417,N_10821,N_10912);
nand U12418 (N_12418,N_11404,N_9381);
and U12419 (N_12419,N_10687,N_11166);
and U12420 (N_12420,N_10625,N_10340);
or U12421 (N_12421,N_10747,N_10219);
or U12422 (N_12422,N_10885,N_9816);
or U12423 (N_12423,N_11905,N_10119);
nor U12424 (N_12424,N_9628,N_9957);
or U12425 (N_12425,N_9699,N_9024);
or U12426 (N_12426,N_9428,N_11023);
or U12427 (N_12427,N_10870,N_10224);
or U12428 (N_12428,N_9853,N_10734);
and U12429 (N_12429,N_9754,N_11524);
or U12430 (N_12430,N_11231,N_11387);
or U12431 (N_12431,N_11022,N_10016);
and U12432 (N_12432,N_11316,N_11435);
nor U12433 (N_12433,N_9256,N_9601);
or U12434 (N_12434,N_11938,N_10087);
and U12435 (N_12435,N_11577,N_9572);
nor U12436 (N_12436,N_9630,N_9749);
nor U12437 (N_12437,N_11000,N_10263);
nor U12438 (N_12438,N_10050,N_10517);
nor U12439 (N_12439,N_9797,N_9719);
nor U12440 (N_12440,N_11964,N_9356);
or U12441 (N_12441,N_9530,N_10824);
or U12442 (N_12442,N_11580,N_11032);
or U12443 (N_12443,N_9623,N_9468);
nand U12444 (N_12444,N_10998,N_10152);
or U12445 (N_12445,N_9277,N_10108);
or U12446 (N_12446,N_9714,N_11464);
or U12447 (N_12447,N_10952,N_10556);
and U12448 (N_12448,N_11458,N_9064);
or U12449 (N_12449,N_9308,N_11015);
or U12450 (N_12450,N_9391,N_10097);
nor U12451 (N_12451,N_9041,N_10904);
or U12452 (N_12452,N_10677,N_11380);
and U12453 (N_12453,N_10836,N_10310);
and U12454 (N_12454,N_10550,N_11933);
nor U12455 (N_12455,N_11189,N_10357);
and U12456 (N_12456,N_10598,N_11812);
nand U12457 (N_12457,N_10571,N_11478);
or U12458 (N_12458,N_10001,N_10938);
nand U12459 (N_12459,N_10766,N_9965);
and U12460 (N_12460,N_10311,N_9454);
and U12461 (N_12461,N_9690,N_11828);
nand U12462 (N_12462,N_11476,N_10808);
and U12463 (N_12463,N_9033,N_9921);
xor U12464 (N_12464,N_10903,N_11687);
nand U12465 (N_12465,N_9472,N_10564);
nand U12466 (N_12466,N_9968,N_10249);
nor U12467 (N_12467,N_10498,N_9467);
or U12468 (N_12468,N_11972,N_10161);
nor U12469 (N_12469,N_9803,N_9265);
and U12470 (N_12470,N_9774,N_10702);
or U12471 (N_12471,N_11757,N_10561);
or U12472 (N_12472,N_9412,N_11077);
nand U12473 (N_12473,N_10610,N_10011);
nor U12474 (N_12474,N_11218,N_9397);
and U12475 (N_12475,N_10305,N_11637);
nor U12476 (N_12476,N_11621,N_9214);
nor U12477 (N_12477,N_11522,N_11084);
and U12478 (N_12478,N_11349,N_9740);
nor U12479 (N_12479,N_11045,N_9326);
nand U12480 (N_12480,N_9889,N_10620);
nor U12481 (N_12481,N_9859,N_10777);
nand U12482 (N_12482,N_11903,N_11526);
and U12483 (N_12483,N_11914,N_11865);
nor U12484 (N_12484,N_10794,N_10973);
and U12485 (N_12485,N_10889,N_9511);
nor U12486 (N_12486,N_10159,N_9333);
nand U12487 (N_12487,N_9931,N_11561);
nand U12488 (N_12488,N_10505,N_11583);
nor U12489 (N_12489,N_11178,N_10739);
nand U12490 (N_12490,N_9879,N_9424);
and U12491 (N_12491,N_9065,N_9314);
or U12492 (N_12492,N_9017,N_10299);
or U12493 (N_12493,N_11261,N_9752);
nor U12494 (N_12494,N_9649,N_11144);
and U12495 (N_12495,N_9626,N_9046);
or U12496 (N_12496,N_9937,N_11034);
nand U12497 (N_12497,N_10367,N_11338);
or U12498 (N_12498,N_9566,N_10235);
nor U12499 (N_12499,N_9387,N_11497);
or U12500 (N_12500,N_9656,N_10399);
and U12501 (N_12501,N_10078,N_9625);
and U12502 (N_12502,N_9782,N_11415);
or U12503 (N_12503,N_10984,N_9257);
nor U12504 (N_12504,N_9141,N_10309);
and U12505 (N_12505,N_11627,N_9014);
and U12506 (N_12506,N_9989,N_11773);
nand U12507 (N_12507,N_11107,N_11593);
nor U12508 (N_12508,N_11810,N_11932);
nor U12509 (N_12509,N_10315,N_10288);
nor U12510 (N_12510,N_10525,N_11001);
and U12511 (N_12511,N_11480,N_9091);
nor U12512 (N_12512,N_10609,N_9414);
or U12513 (N_12513,N_9404,N_11010);
nor U12514 (N_12514,N_11373,N_9683);
and U12515 (N_12515,N_10758,N_11724);
nand U12516 (N_12516,N_9680,N_9420);
and U12517 (N_12517,N_11056,N_9647);
and U12518 (N_12518,N_9315,N_10461);
or U12519 (N_12519,N_11270,N_9878);
or U12520 (N_12520,N_10546,N_11321);
nor U12521 (N_12521,N_10694,N_10831);
nor U12522 (N_12522,N_10990,N_10391);
and U12523 (N_12523,N_11970,N_10081);
and U12524 (N_12524,N_11774,N_9201);
nor U12525 (N_12525,N_9135,N_10538);
or U12526 (N_12526,N_11958,N_11279);
and U12527 (N_12527,N_9757,N_10316);
or U12528 (N_12528,N_9606,N_10876);
or U12529 (N_12529,N_11999,N_9881);
nand U12530 (N_12530,N_11287,N_10143);
or U12531 (N_12531,N_11682,N_9018);
nand U12532 (N_12532,N_11198,N_9443);
nor U12533 (N_12533,N_10194,N_10617);
or U12534 (N_12534,N_11949,N_11552);
or U12535 (N_12535,N_11006,N_10459);
nor U12536 (N_12536,N_9864,N_9622);
nand U12537 (N_12537,N_9687,N_9590);
and U12538 (N_12538,N_10478,N_11335);
and U12539 (N_12539,N_11751,N_11483);
nand U12540 (N_12540,N_9440,N_11008);
nor U12541 (N_12541,N_10920,N_10287);
or U12542 (N_12542,N_9115,N_10402);
and U12543 (N_12543,N_9164,N_10674);
or U12544 (N_12544,N_9426,N_11059);
nand U12545 (N_12545,N_11159,N_11446);
and U12546 (N_12546,N_10913,N_10621);
and U12547 (N_12547,N_10689,N_9058);
and U12548 (N_12548,N_11334,N_9935);
nor U12549 (N_12549,N_10006,N_10635);
nor U12550 (N_12550,N_9189,N_10320);
and U12551 (N_12551,N_10307,N_11587);
nand U12552 (N_12552,N_9849,N_10640);
nand U12553 (N_12553,N_11152,N_11076);
and U12554 (N_12554,N_11622,N_9096);
or U12555 (N_12555,N_10690,N_10656);
xnor U12556 (N_12556,N_10437,N_9573);
or U12557 (N_12557,N_11794,N_10535);
nor U12558 (N_12558,N_10271,N_9045);
and U12559 (N_12559,N_10711,N_9126);
nand U12560 (N_12560,N_10401,N_9340);
nor U12561 (N_12561,N_10989,N_9075);
and U12562 (N_12562,N_11694,N_11809);
nand U12563 (N_12563,N_11796,N_9327);
nand U12564 (N_12564,N_11831,N_11420);
and U12565 (N_12565,N_9726,N_10999);
nand U12566 (N_12566,N_11213,N_10592);
nand U12567 (N_12567,N_11188,N_9089);
and U12568 (N_12568,N_9823,N_9799);
nand U12569 (N_12569,N_10629,N_10901);
nor U12570 (N_12570,N_10932,N_10445);
nand U12571 (N_12571,N_9748,N_9390);
nand U12572 (N_12572,N_9292,N_10455);
nor U12573 (N_12573,N_10895,N_9143);
nor U12574 (N_12574,N_11613,N_10654);
and U12575 (N_12575,N_11851,N_10026);
or U12576 (N_12576,N_10568,N_10270);
nand U12577 (N_12577,N_9070,N_11663);
nand U12578 (N_12578,N_11612,N_11347);
or U12579 (N_12579,N_10850,N_11976);
and U12580 (N_12580,N_10054,N_9246);
nor U12581 (N_12581,N_10804,N_9685);
nor U12582 (N_12582,N_9639,N_10134);
nand U12583 (N_12583,N_9953,N_9172);
and U12584 (N_12584,N_10866,N_9200);
and U12585 (N_12585,N_10881,N_10572);
nor U12586 (N_12586,N_9657,N_11533);
or U12587 (N_12587,N_10892,N_10763);
nor U12588 (N_12588,N_11604,N_11962);
nor U12589 (N_12589,N_9359,N_9669);
nand U12590 (N_12590,N_9417,N_11636);
or U12591 (N_12591,N_10470,N_11717);
and U12592 (N_12592,N_9890,N_9952);
and U12593 (N_12593,N_11598,N_10603);
or U12594 (N_12594,N_11310,N_11379);
nand U12595 (N_12595,N_11823,N_10545);
or U12596 (N_12596,N_11036,N_9650);
nand U12597 (N_12597,N_9960,N_11556);
nor U12598 (N_12598,N_10695,N_11228);
or U12599 (N_12599,N_9589,N_10416);
and U12600 (N_12600,N_11220,N_10306);
nand U12601 (N_12601,N_9948,N_11922);
nor U12602 (N_12602,N_9098,N_10865);
or U12603 (N_12603,N_9581,N_11499);
nand U12604 (N_12604,N_10584,N_11995);
or U12605 (N_12605,N_9824,N_11062);
nor U12606 (N_12606,N_9793,N_11911);
nand U12607 (N_12607,N_11222,N_10070);
nand U12608 (N_12608,N_9891,N_11149);
nand U12609 (N_12609,N_9262,N_11558);
and U12610 (N_12610,N_10125,N_9088);
and U12611 (N_12611,N_11700,N_11237);
or U12612 (N_12612,N_11660,N_9672);
nor U12613 (N_12613,N_9140,N_9540);
or U12614 (N_12614,N_9396,N_9251);
nand U12615 (N_12615,N_9266,N_9934);
or U12616 (N_12616,N_10987,N_11614);
and U12617 (N_12617,N_10847,N_9032);
or U12618 (N_12618,N_11675,N_10604);
or U12619 (N_12619,N_9517,N_11864);
or U12620 (N_12620,N_11866,N_10033);
nand U12621 (N_12621,N_11723,N_9072);
nand U12622 (N_12622,N_9334,N_9969);
nand U12623 (N_12623,N_9300,N_11920);
or U12624 (N_12624,N_9123,N_10843);
and U12625 (N_12625,N_9447,N_10644);
and U12626 (N_12626,N_10992,N_9868);
nor U12627 (N_12627,N_10646,N_11677);
and U12628 (N_12628,N_11035,N_9858);
or U12629 (N_12629,N_11772,N_9405);
and U12630 (N_12630,N_11889,N_11945);
and U12631 (N_12631,N_10722,N_11280);
and U12632 (N_12632,N_9282,N_9124);
nor U12633 (N_12633,N_10121,N_9015);
nor U12634 (N_12634,N_11139,N_10991);
or U12635 (N_12635,N_10122,N_9139);
or U12636 (N_12636,N_11521,N_9983);
or U12637 (N_12637,N_11785,N_11709);
nor U12638 (N_12638,N_10180,N_9842);
nand U12639 (N_12639,N_11750,N_10576);
nand U12640 (N_12640,N_9310,N_9811);
and U12641 (N_12641,N_10202,N_10373);
and U12642 (N_12642,N_10890,N_9856);
nor U12643 (N_12643,N_11775,N_10030);
nor U12644 (N_12644,N_10491,N_9279);
or U12645 (N_12645,N_9950,N_11203);
xor U12646 (N_12646,N_9895,N_9759);
nand U12647 (N_12647,N_11135,N_9794);
or U12648 (N_12648,N_11681,N_10007);
or U12649 (N_12649,N_10480,N_9731);
nor U12650 (N_12650,N_9100,N_10040);
nor U12651 (N_12651,N_10395,N_9703);
and U12652 (N_12652,N_10649,N_10295);
and U12653 (N_12653,N_10943,N_9346);
and U12654 (N_12654,N_10481,N_10213);
or U12655 (N_12655,N_11225,N_9538);
nand U12656 (N_12656,N_11566,N_11289);
and U12657 (N_12657,N_9790,N_11620);
nand U12658 (N_12658,N_9837,N_10995);
nor U12659 (N_12659,N_11844,N_11863);
or U12660 (N_12660,N_11325,N_11883);
or U12661 (N_12661,N_11565,N_10811);
or U12662 (N_12662,N_9808,N_11702);
or U12663 (N_12663,N_9673,N_11055);
nor U12664 (N_12664,N_9363,N_11243);
nand U12665 (N_12665,N_10427,N_11635);
nor U12666 (N_12666,N_11223,N_9735);
nand U12667 (N_12667,N_11619,N_11944);
and U12668 (N_12668,N_10879,N_11894);
nor U12669 (N_12669,N_11482,N_11209);
nor U12670 (N_12670,N_11606,N_9336);
nor U12671 (N_12671,N_10128,N_10834);
nor U12672 (N_12672,N_9129,N_10274);
nor U12673 (N_12673,N_11443,N_11979);
and U12674 (N_12674,N_9038,N_11766);
and U12675 (N_12675,N_11996,N_11355);
and U12676 (N_12676,N_11572,N_10374);
or U12677 (N_12677,N_10096,N_9775);
or U12678 (N_12678,N_10453,N_10547);
and U12679 (N_12679,N_10893,N_9705);
and U12680 (N_12680,N_9870,N_11721);
and U12681 (N_12681,N_11066,N_11813);
or U12682 (N_12682,N_11265,N_11029);
nor U12683 (N_12683,N_11653,N_10636);
nor U12684 (N_12684,N_10072,N_9460);
nor U12685 (N_12685,N_11408,N_9288);
or U12686 (N_12686,N_11508,N_11185);
nand U12687 (N_12687,N_11811,N_10010);
or U12688 (N_12688,N_10071,N_11259);
nor U12689 (N_12689,N_9393,N_10434);
or U12690 (N_12690,N_9679,N_10586);
nor U12691 (N_12691,N_9401,N_10479);
xnor U12692 (N_12692,N_9654,N_10429);
and U12693 (N_12693,N_11701,N_9900);
nand U12694 (N_12694,N_9441,N_10537);
or U12695 (N_12695,N_10297,N_9357);
nand U12696 (N_12696,N_9325,N_11611);
nor U12697 (N_12697,N_9621,N_9081);
nor U12698 (N_12698,N_9539,N_9388);
nor U12699 (N_12699,N_11657,N_10246);
or U12700 (N_12700,N_11303,N_10339);
and U12701 (N_12701,N_9026,N_10529);
and U12702 (N_12702,N_10509,N_11065);
nand U12703 (N_12703,N_11171,N_11311);
and U12704 (N_12704,N_11639,N_11674);
nand U12705 (N_12705,N_10981,N_11752);
or U12706 (N_12706,N_10039,N_11527);
and U12707 (N_12707,N_10494,N_11680);
nand U12708 (N_12708,N_11862,N_9773);
nand U12709 (N_12709,N_9160,N_10032);
nor U12710 (N_12710,N_9136,N_9261);
nand U12711 (N_12711,N_10438,N_11140);
nand U12712 (N_12712,N_11439,N_9697);
nor U12713 (N_12713,N_11801,N_9605);
and U12714 (N_12714,N_9016,N_11021);
nand U12715 (N_12715,N_11406,N_10059);
nor U12716 (N_12716,N_9885,N_10038);
or U12717 (N_12717,N_10165,N_11819);
nor U12718 (N_12718,N_9764,N_9541);
and U12719 (N_12719,N_11041,N_10080);
nor U12720 (N_12720,N_10217,N_11890);
or U12721 (N_12721,N_11656,N_11983);
or U12722 (N_12722,N_9552,N_10066);
nor U12723 (N_12723,N_11269,N_10350);
nor U12724 (N_12724,N_11148,N_11290);
or U12725 (N_12725,N_11936,N_11190);
and U12726 (N_12726,N_10185,N_10497);
or U12727 (N_12727,N_11384,N_9291);
nand U12728 (N_12728,N_9392,N_9204);
and U12729 (N_12729,N_10818,N_9222);
and U12730 (N_12730,N_11046,N_10823);
or U12731 (N_12731,N_10129,N_10828);
and U12732 (N_12732,N_10947,N_9534);
or U12733 (N_12733,N_11351,N_10201);
or U12734 (N_12734,N_9695,N_9118);
or U12735 (N_12735,N_11388,N_10861);
or U12736 (N_12736,N_10321,N_9199);
and U12737 (N_12737,N_10179,N_10941);
or U12738 (N_12738,N_9394,N_10682);
or U12739 (N_12739,N_9111,N_11169);
nand U12740 (N_12740,N_11105,N_10173);
nand U12741 (N_12741,N_9551,N_9640);
and U12742 (N_12742,N_9180,N_10916);
xnor U12743 (N_12743,N_9732,N_9449);
and U12744 (N_12744,N_10599,N_11605);
nor U12745 (N_12745,N_9670,N_9205);
and U12746 (N_12746,N_10822,N_10506);
or U12747 (N_12747,N_11393,N_9629);
nand U12748 (N_12748,N_10955,N_11984);
and U12749 (N_12749,N_10749,N_9252);
nand U12750 (N_12750,N_10846,N_11732);
or U12751 (N_12751,N_10359,N_11711);
nor U12752 (N_12752,N_9062,N_10755);
nor U12753 (N_12753,N_11389,N_11969);
xor U12754 (N_12754,N_10737,N_9298);
nand U12755 (N_12755,N_11150,N_9182);
or U12756 (N_12756,N_9317,N_10676);
or U12757 (N_12757,N_11676,N_10869);
nor U12758 (N_12758,N_10567,N_10945);
nor U12759 (N_12759,N_11525,N_10806);
or U12760 (N_12760,N_10688,N_9231);
or U12761 (N_12761,N_11846,N_10863);
nand U12762 (N_12762,N_10764,N_10136);
nor U12763 (N_12763,N_11170,N_10956);
nand U12764 (N_12764,N_9765,N_9631);
nand U12765 (N_12765,N_11451,N_11727);
and U12766 (N_12766,N_11286,N_11250);
and U12767 (N_12767,N_10612,N_11329);
nor U12768 (N_12768,N_9054,N_11096);
or U12769 (N_12769,N_10112,N_11264);
nand U12770 (N_12770,N_9459,N_11293);
nor U12771 (N_12771,N_10345,N_9554);
or U12772 (N_12772,N_11374,N_11990);
nor U12773 (N_12773,N_11168,N_11837);
nand U12774 (N_12774,N_11753,N_10697);
or U12775 (N_12775,N_9122,N_11833);
or U12776 (N_12776,N_9836,N_10551);
and U12777 (N_12777,N_10163,N_11295);
nor U12778 (N_12778,N_10954,N_9177);
nor U12779 (N_12779,N_11494,N_11641);
nor U12780 (N_12780,N_11313,N_10385);
and U12781 (N_12781,N_9743,N_9432);
nor U12782 (N_12782,N_10204,N_10853);
nand U12783 (N_12783,N_10680,N_11033);
and U12784 (N_12784,N_10502,N_9897);
nor U12785 (N_12785,N_10238,N_10292);
or U12786 (N_12786,N_11688,N_9496);
nand U12787 (N_12787,N_9169,N_9211);
nand U12788 (N_12788,N_9052,N_10717);
nor U12789 (N_12789,N_10118,N_9728);
nor U12790 (N_12790,N_9042,N_10460);
or U12791 (N_12791,N_10613,N_11383);
nand U12792 (N_12792,N_9283,N_11405);
and U12793 (N_12793,N_10451,N_10748);
or U12794 (N_12794,N_11402,N_11907);
nor U12795 (N_12795,N_11574,N_11288);
nand U12796 (N_12796,N_9207,N_11957);
nand U12797 (N_12797,N_11226,N_10055);
or U12798 (N_12798,N_10389,N_10043);
xnor U12799 (N_12799,N_11086,N_10918);
or U12800 (N_12800,N_9466,N_9866);
and U12801 (N_12801,N_10113,N_9275);
and U12802 (N_12802,N_11679,N_10063);
and U12803 (N_12803,N_10390,N_11143);
nor U12804 (N_12804,N_10266,N_9763);
nand U12805 (N_12805,N_10192,N_9299);
nor U12806 (N_12806,N_11886,N_10743);
nor U12807 (N_12807,N_11044,N_9444);
and U12808 (N_12808,N_9437,N_11007);
and U12809 (N_12809,N_11211,N_11137);
nand U12810 (N_12810,N_9106,N_10114);
or U12811 (N_12811,N_11429,N_10131);
nand U12812 (N_12812,N_9615,N_11698);
nand U12813 (N_12813,N_9039,N_9389);
and U12814 (N_12814,N_10475,N_11973);
and U12815 (N_12815,N_10421,N_11912);
nor U12816 (N_12816,N_10254,N_10628);
xor U12817 (N_12817,N_10939,N_10467);
nand U12818 (N_12818,N_10523,N_11559);
or U12819 (N_12819,N_11879,N_9792);
nor U12820 (N_12820,N_9660,N_10267);
and U12821 (N_12821,N_11336,N_10231);
nand U12822 (N_12822,N_10335,N_11515);
nand U12823 (N_12823,N_9151,N_10996);
nor U12824 (N_12824,N_9051,N_10531);
and U12825 (N_12825,N_9809,N_9620);
nand U12826 (N_12826,N_9138,N_10988);
or U12827 (N_12827,N_10825,N_9219);
and U12828 (N_12828,N_11236,N_11503);
nor U12829 (N_12829,N_9902,N_9196);
and U12830 (N_12830,N_9379,N_11093);
nor U12831 (N_12831,N_9481,N_10648);
nand U12832 (N_12832,N_9981,N_9845);
and U12833 (N_12833,N_11426,N_10978);
nor U12834 (N_12834,N_11146,N_9215);
nand U12835 (N_12835,N_11665,N_11343);
and U12836 (N_12836,N_11591,N_9929);
nor U12837 (N_12837,N_11963,N_10234);
nor U12838 (N_12838,N_11634,N_9966);
and U12839 (N_12839,N_9239,N_11493);
and U12840 (N_12840,N_11590,N_9305);
and U12841 (N_12841,N_10024,N_10908);
and U12842 (N_12842,N_10312,N_11233);
nor U12843 (N_12843,N_10880,N_9061);
or U12844 (N_12844,N_10548,N_11398);
or U12845 (N_12845,N_10403,N_9851);
nand U12846 (N_12846,N_10857,N_11194);
or U12847 (N_12847,N_11926,N_11629);
or U12848 (N_12848,N_9607,N_11207);
nand U12849 (N_12849,N_11496,N_11391);
nand U12850 (N_12850,N_10776,N_9833);
nand U12851 (N_12851,N_9486,N_11488);
or U12852 (N_12852,N_11057,N_11909);
or U12853 (N_12853,N_11372,N_9689);
or U12854 (N_12854,N_9165,N_9007);
or U12855 (N_12855,N_9819,N_11505);
nor U12856 (N_12856,N_11551,N_10796);
or U12857 (N_12857,N_11780,N_9761);
nor U12858 (N_12858,N_9241,N_10492);
nor U12859 (N_12859,N_11427,N_10140);
and U12860 (N_12860,N_10482,N_9119);
and U12861 (N_12861,N_11689,N_11795);
nor U12862 (N_12862,N_11885,N_9329);
nor U12863 (N_12863,N_10144,N_11263);
nor U12864 (N_12864,N_11005,N_9991);
xor U12865 (N_12865,N_9920,N_9994);
or U12866 (N_12866,N_10557,N_11948);
nand U12867 (N_12867,N_11930,N_10735);
and U12868 (N_12868,N_9413,N_10265);
or U12869 (N_12869,N_9576,N_11584);
or U12870 (N_12870,N_9320,N_9821);
or U12871 (N_12871,N_11900,N_11068);
nor U12872 (N_12872,N_11098,N_9380);
nor U12873 (N_12873,N_10623,N_9076);
nor U12874 (N_12874,N_9616,N_9549);
nor U12875 (N_12875,N_9603,N_11880);
nor U12876 (N_12876,N_9899,N_9820);
or U12877 (N_12877,N_11980,N_10753);
nand U12878 (N_12878,N_11906,N_9269);
or U12879 (N_12879,N_10971,N_9995);
or U12880 (N_12880,N_10770,N_9583);
and U12881 (N_12881,N_10277,N_11668);
and U12882 (N_12882,N_10215,N_10914);
nand U12883 (N_12883,N_11162,N_9815);
nand U12884 (N_12884,N_11655,N_11807);
or U12885 (N_12885,N_9059,N_9125);
nand U12886 (N_12886,N_11423,N_9113);
or U12887 (N_12887,N_11312,N_10606);
nor U12888 (N_12888,N_10532,N_10499);
and U12889 (N_12889,N_10358,N_9280);
or U12890 (N_12890,N_11771,N_10392);
nand U12891 (N_12891,N_10515,N_11201);
or U12892 (N_12892,N_10326,N_11424);
or U12893 (N_12893,N_9408,N_10126);
nor U12894 (N_12894,N_11157,N_11782);
or U12895 (N_12895,N_10142,N_11977);
and U12896 (N_12896,N_11048,N_10706);
or U12897 (N_12897,N_9226,N_10630);
and U12898 (N_12898,N_9562,N_10052);
nand U12899 (N_12899,N_10512,N_11730);
and U12900 (N_12900,N_9565,N_10503);
or U12901 (N_12901,N_9350,N_11516);
or U12902 (N_12902,N_9958,N_9227);
or U12903 (N_12903,N_9645,N_10486);
nand U12904 (N_12904,N_9976,N_9597);
nand U12905 (N_12905,N_9807,N_10719);
or U12906 (N_12906,N_9906,N_9120);
or U12907 (N_12907,N_10767,N_11713);
nor U12908 (N_12908,N_10283,N_9575);
and U12909 (N_12909,N_11315,N_10060);
nor U12910 (N_12910,N_11208,N_10810);
nor U12911 (N_12911,N_10138,N_9294);
and U12912 (N_12912,N_9854,N_10216);
nand U12913 (N_12913,N_10200,N_10911);
or U12914 (N_12914,N_11781,N_11054);
or U12915 (N_12915,N_11966,N_10137);
and U12916 (N_12916,N_11440,N_10124);
nor U12917 (N_12917,N_9710,N_10171);
xnor U12918 (N_12918,N_9693,N_9865);
nand U12919 (N_12919,N_10501,N_9563);
or U12920 (N_12920,N_9544,N_11410);
nand U12921 (N_12921,N_10788,N_9185);
or U12922 (N_12922,N_10664,N_10149);
and U12923 (N_12923,N_11394,N_11859);
or U12924 (N_12924,N_9862,N_9653);
or U12925 (N_12925,N_9962,N_10560);
nand U12926 (N_12926,N_11895,N_11960);
nand U12927 (N_12927,N_10508,N_11998);
and U12928 (N_12928,N_10456,N_10036);
or U12929 (N_12929,N_10172,N_9750);
nand U12930 (N_12930,N_9867,N_11686);
and U12931 (N_12931,N_11695,N_10684);
or U12932 (N_12932,N_10958,N_11247);
and U12933 (N_12933,N_10034,N_9237);
and U12934 (N_12934,N_9416,N_10167);
nand U12935 (N_12935,N_10645,N_10132);
and U12936 (N_12936,N_10106,N_11474);
nor U12937 (N_12937,N_10626,N_9480);
and U12938 (N_12938,N_11470,N_11416);
nand U12939 (N_12939,N_11817,N_10883);
nand U12940 (N_12940,N_9686,N_9578);
nand U12941 (N_12941,N_9349,N_10332);
nor U12942 (N_12942,N_10527,N_10573);
nand U12943 (N_12943,N_9216,N_10730);
and U12944 (N_12944,N_11869,N_10549);
nand U12945 (N_12945,N_10678,N_11377);
or U12946 (N_12946,N_11648,N_10530);
nor U12947 (N_12947,N_11354,N_9901);
nor U12948 (N_12948,N_11020,N_9343);
nor U12949 (N_12949,N_9110,N_10111);
nor U12950 (N_12950,N_9455,N_10430);
nand U12951 (N_12951,N_10960,N_11417);
and U12952 (N_12952,N_9276,N_11205);
and U12953 (N_12953,N_11888,N_11543);
or U12954 (N_12954,N_10009,N_11276);
nor U12955 (N_12955,N_10704,N_11433);
nor U12956 (N_12956,N_10723,N_9385);
and U12957 (N_12957,N_9352,N_9031);
and U12958 (N_12958,N_10791,N_11881);
nand U12959 (N_12959,N_11741,N_9430);
nor U12960 (N_12960,N_10585,N_11762);
nor U12961 (N_12961,N_9527,N_9235);
and U12962 (N_12962,N_9339,N_10175);
nand U12963 (N_12963,N_9951,N_9131);
and U12964 (N_12964,N_10252,N_9783);
nand U12965 (N_12965,N_9582,N_9442);
or U12966 (N_12966,N_9652,N_11765);
nor U12967 (N_12967,N_9395,N_11024);
or U12968 (N_12968,N_11848,N_9370);
and U12969 (N_12969,N_9445,N_11072);
nand U12970 (N_12970,N_11436,N_11210);
and U12971 (N_12971,N_10284,N_11569);
or U12972 (N_12972,N_11567,N_9484);
or U12973 (N_12973,N_11761,N_10251);
and U12974 (N_12974,N_10346,N_11318);
nand U12975 (N_12975,N_9382,N_11645);
and U12976 (N_12976,N_11003,N_11492);
and U12977 (N_12977,N_9471,N_10232);
or U12978 (N_12978,N_10396,N_9209);
and U12979 (N_12979,N_10334,N_11317);
and U12980 (N_12980,N_11353,N_10002);
nor U12981 (N_12981,N_11787,N_10045);
nand U12982 (N_12982,N_11407,N_9371);
and U12983 (N_12983,N_9698,N_9875);
and U12984 (N_12984,N_9184,N_11814);
nor U12985 (N_12985,N_10420,N_10562);
nor U12986 (N_12986,N_11873,N_10727);
nand U12987 (N_12987,N_11165,N_9910);
or U12988 (N_12988,N_9818,N_10405);
or U12989 (N_12989,N_10516,N_9335);
and U12990 (N_12990,N_11541,N_9153);
and U12991 (N_12991,N_10341,N_11132);
nor U12992 (N_12992,N_9924,N_11115);
or U12993 (N_12993,N_9406,N_11187);
nand U12994 (N_12994,N_11161,N_9069);
or U12995 (N_12995,N_9785,N_9309);
and U12996 (N_12996,N_9161,N_10074);
or U12997 (N_12997,N_10841,N_11019);
nand U12998 (N_12998,N_11872,N_11658);
nor U12999 (N_12999,N_10579,N_9178);
nand U13000 (N_13000,N_11080,N_11385);
and U13001 (N_13001,N_11141,N_9940);
nand U13002 (N_13002,N_11272,N_10651);
and U13003 (N_13003,N_9155,N_11662);
nor U13004 (N_13004,N_9676,N_9366);
nor U13005 (N_13005,N_9556,N_9005);
or U13006 (N_13006,N_11163,N_9012);
nand U13007 (N_13007,N_10731,N_11114);
nand U13008 (N_13008,N_10372,N_10588);
nand U13009 (N_13009,N_11099,N_11414);
nor U13010 (N_13010,N_9399,N_9273);
nor U13011 (N_13011,N_10426,N_11640);
nor U13012 (N_13012,N_11738,N_11309);
and U13013 (N_13013,N_11854,N_10902);
or U13014 (N_13014,N_10738,N_11255);
nand U13015 (N_13015,N_11403,N_10983);
nand U13016 (N_13016,N_10994,N_11460);
and U13017 (N_13017,N_11770,N_10507);
nand U13018 (N_13018,N_9483,N_11726);
and U13019 (N_13019,N_9896,N_11485);
nand U13020 (N_13020,N_9504,N_11200);
nand U13021 (N_13021,N_10436,N_10848);
nor U13022 (N_13022,N_9827,N_10732);
and U13023 (N_13023,N_10351,N_9488);
nand U13024 (N_13024,N_10222,N_9861);
or U13025 (N_13025,N_11304,N_11400);
nor U13026 (N_13026,N_9116,N_11666);
and U13027 (N_13027,N_10025,N_11986);
xor U13028 (N_13028,N_10667,N_11432);
nor U13029 (N_13029,N_10422,N_9599);
or U13030 (N_13030,N_10589,N_9470);
nand U13031 (N_13031,N_10379,N_11246);
nor U13032 (N_13032,N_9642,N_10982);
and U13033 (N_13033,N_9508,N_9342);
nor U13034 (N_13034,N_9949,N_9560);
and U13035 (N_13035,N_10440,N_9084);
and U13036 (N_13036,N_9228,N_10275);
and U13037 (N_13037,N_10255,N_10415);
nand U13038 (N_13038,N_9290,N_10856);
nand U13039 (N_13039,N_11235,N_10917);
nor U13040 (N_13040,N_11472,N_9800);
nand U13041 (N_13041,N_10618,N_11858);
nand U13042 (N_13042,N_9520,N_9987);
and U13043 (N_13043,N_10759,N_10744);
nor U13044 (N_13044,N_10199,N_9586);
nand U13045 (N_13045,N_10386,N_10668);
or U13046 (N_13046,N_10707,N_11078);
and U13047 (N_13047,N_11646,N_11307);
and U13048 (N_13048,N_10862,N_11042);
and U13049 (N_13049,N_11245,N_11025);
and U13050 (N_13050,N_11227,N_10462);
and U13051 (N_13051,N_11553,N_11248);
nor U13052 (N_13052,N_11991,N_10558);
or U13053 (N_13053,N_11131,N_10260);
or U13054 (N_13054,N_11258,N_10285);
nor U13055 (N_13055,N_11361,N_9409);
or U13056 (N_13056,N_11230,N_11278);
nor U13057 (N_13057,N_9281,N_11510);
or U13058 (N_13058,N_10624,N_9925);
nor U13059 (N_13059,N_10414,N_9817);
and U13060 (N_13060,N_10253,N_9564);
nand U13061 (N_13061,N_9229,N_9733);
nand U13062 (N_13062,N_9786,N_10223);
nand U13063 (N_13063,N_11122,N_9351);
and U13064 (N_13064,N_10922,N_9008);
nand U13065 (N_13065,N_10280,N_10653);
nor U13066 (N_13066,N_9374,N_11707);
xor U13067 (N_13067,N_11366,N_9997);
and U13068 (N_13068,N_10574,N_10318);
nor U13069 (N_13069,N_11931,N_11892);
nor U13070 (N_13070,N_10830,N_9107);
nand U13071 (N_13071,N_10388,N_9344);
and U13072 (N_13072,N_11925,N_9332);
and U13073 (N_13073,N_9297,N_11950);
xor U13074 (N_13074,N_11955,N_11300);
nor U13075 (N_13075,N_11028,N_10102);
nand U13076 (N_13076,N_9121,N_9009);
nor U13077 (N_13077,N_10093,N_9720);
nor U13078 (N_13078,N_11842,N_10775);
nand U13079 (N_13079,N_10511,N_9835);
or U13080 (N_13080,N_10800,N_10444);
or U13081 (N_13081,N_11849,N_10109);
and U13082 (N_13082,N_11108,N_9734);
or U13083 (N_13083,N_11229,N_9474);
nor U13084 (N_13084,N_11518,N_10076);
or U13085 (N_13085,N_11442,N_10068);
nand U13086 (N_13086,N_9869,N_10352);
nor U13087 (N_13087,N_9027,N_11051);
or U13088 (N_13088,N_10225,N_10323);
nor U13089 (N_13089,N_10700,N_11103);
and U13090 (N_13090,N_9453,N_11378);
or U13091 (N_13091,N_10008,N_9919);
nor U13092 (N_13092,N_9402,N_9770);
or U13093 (N_13093,N_9848,N_10290);
or U13094 (N_13094,N_9034,N_9701);
nor U13095 (N_13095,N_11511,N_9361);
and U13096 (N_13096,N_9307,N_11455);
nand U13097 (N_13097,N_11910,N_11489);
nand U13098 (N_13098,N_9220,N_10377);
nand U13099 (N_13099,N_10425,N_10289);
nor U13100 (N_13100,N_9056,N_11599);
nor U13101 (N_13101,N_9477,N_10833);
nor U13102 (N_13102,N_11428,N_10590);
or U13103 (N_13103,N_10740,N_10795);
and U13104 (N_13104,N_9980,N_9128);
nand U13105 (N_13105,N_11625,N_11971);
and U13106 (N_13106,N_11365,N_11356);
nand U13107 (N_13107,N_10104,N_11749);
nand U13108 (N_13108,N_9715,N_10714);
nor U13109 (N_13109,N_9322,N_9337);
or U13110 (N_13110,N_9218,N_11090);
and U13111 (N_13111,N_11719,N_11507);
nand U13112 (N_13112,N_10891,N_9681);
nand U13113 (N_13113,N_10554,N_9202);
and U13114 (N_13114,N_10441,N_11946);
nor U13115 (N_13115,N_9646,N_10786);
or U13116 (N_13116,N_11517,N_9964);
or U13117 (N_13117,N_11136,N_10985);
and U13118 (N_13118,N_11916,N_11238);
and U13119 (N_13119,N_9094,N_10803);
nor U13120 (N_13120,N_11670,N_9977);
or U13121 (N_13121,N_9173,N_9898);
nand U13122 (N_13122,N_11314,N_11685);
nand U13123 (N_13123,N_11904,N_11206);
or U13124 (N_13124,N_11544,N_9577);
nand U13125 (N_13125,N_9795,N_9513);
and U13126 (N_13126,N_10524,N_9347);
nor U13127 (N_13127,N_11693,N_10439);
and U13128 (N_13128,N_10781,N_11127);
xor U13129 (N_13129,N_9495,N_9528);
xnor U13130 (N_13130,N_10591,N_9644);
nand U13131 (N_13131,N_11870,N_10634);
nand U13132 (N_13132,N_10041,N_10725);
or U13133 (N_13133,N_10064,N_10361);
and U13134 (N_13134,N_11075,N_10929);
or U13135 (N_13135,N_10886,N_11344);
nand U13136 (N_13136,N_10115,N_11182);
or U13137 (N_13137,N_11935,N_11617);
nand U13138 (N_13138,N_10543,N_11386);
nor U13139 (N_13139,N_11487,N_11186);
nor U13140 (N_13140,N_9154,N_9197);
or U13141 (N_13141,N_10174,N_10936);
and U13142 (N_13142,N_9674,N_9608);
and U13143 (N_13143,N_11500,N_11012);
and U13144 (N_13144,N_9526,N_9378);
nand U13145 (N_13145,N_9296,N_11453);
nand U13146 (N_13146,N_10449,N_11769);
nand U13147 (N_13147,N_11841,N_11179);
or U13148 (N_13148,N_11467,N_9166);
nor U13149 (N_13149,N_9971,N_9522);
or U13150 (N_13150,N_11615,N_10139);
nor U13151 (N_13151,N_10805,N_11085);
xnor U13152 (N_13152,N_11471,N_9376);
and U13153 (N_13153,N_9766,N_9010);
or U13154 (N_13154,N_9029,N_11282);
nor U13155 (N_13155,N_11117,N_9713);
or U13156 (N_13156,N_11221,N_10319);
nand U13157 (N_13157,N_10276,N_10349);
and U13158 (N_13158,N_9954,N_10972);
and U13159 (N_13159,N_9082,N_9712);
and U13160 (N_13160,N_9737,N_9959);
and U13161 (N_13161,N_11498,N_10797);
xor U13162 (N_13162,N_10211,N_11484);
nor U13163 (N_13163,N_10079,N_9863);
or U13164 (N_13164,N_10187,N_10686);
and U13165 (N_13165,N_9641,N_11087);
or U13166 (N_13166,N_10860,N_11529);
or U13167 (N_13167,N_9537,N_11899);
or U13168 (N_13168,N_9159,N_11759);
and U13169 (N_13169,N_9104,N_11722);
and U13170 (N_13170,N_9473,N_10368);
nor U13171 (N_13171,N_10915,N_9485);
nand U13172 (N_13172,N_10712,N_11631);
nand U13173 (N_13173,N_10446,N_10726);
and U13174 (N_13174,N_11968,N_10575);
and U13175 (N_13175,N_9503,N_9421);
or U13176 (N_13176,N_11790,N_11038);
nor U13177 (N_13177,N_9611,N_11016);
and U13178 (N_13178,N_9928,N_10720);
and U13179 (N_13179,N_11940,N_9244);
and U13180 (N_13180,N_10206,N_11411);
and U13181 (N_13181,N_9411,N_9338);
and U13182 (N_13182,N_10887,N_9410);
or U13183 (N_13183,N_11928,N_9436);
nor U13184 (N_13184,N_9223,N_11705);
and U13185 (N_13185,N_11768,N_9840);
or U13186 (N_13186,N_10364,N_11626);
nor U13187 (N_13187,N_10541,N_9191);
nor U13188 (N_13188,N_11040,N_11506);
nand U13189 (N_13189,N_11324,N_9512);
nor U13190 (N_13190,N_11652,N_10476);
xor U13191 (N_13191,N_9594,N_11875);
nor U13192 (N_13192,N_9973,N_10563);
nand U13193 (N_13193,N_9323,N_11718);
nor U13194 (N_13194,N_10153,N_11608);
or U13195 (N_13195,N_11857,N_10151);
or U13196 (N_13196,N_9450,N_9912);
and U13197 (N_13197,N_10967,N_11273);
nand U13198 (N_13198,N_11342,N_11441);
or U13199 (N_13199,N_10608,N_10814);
or U13200 (N_13200,N_9903,N_10581);
or U13201 (N_13201,N_9362,N_10090);
nor U13202 (N_13202,N_11319,N_11376);
nand U13203 (N_13203,N_11874,N_10207);
nand U13204 (N_13204,N_10183,N_11563);
and U13205 (N_13205,N_11610,N_9469);
or U13206 (N_13206,N_11628,N_9272);
or U13207 (N_13207,N_10098,N_10669);
or U13208 (N_13208,N_10874,N_10611);
and U13209 (N_13209,N_11249,N_11509);
and U13210 (N_13210,N_9137,N_11512);
nand U13211 (N_13211,N_10435,N_11167);
and U13212 (N_13212,N_9429,N_11692);
or U13213 (N_13213,N_11298,N_9545);
nor U13214 (N_13214,N_9591,N_11130);
nor U13215 (N_13215,N_10643,N_10338);
nor U13216 (N_13216,N_10580,N_11017);
nand U13217 (N_13217,N_9758,N_11339);
and U13218 (N_13218,N_9730,N_9245);
nor U13219 (N_13219,N_11124,N_9482);
nand U13220 (N_13220,N_9148,N_9478);
and U13221 (N_13221,N_9985,N_10120);
or U13222 (N_13222,N_10048,N_9225);
nand U13223 (N_13223,N_11129,N_11729);
nand U13224 (N_13224,N_9158,N_9841);
and U13225 (N_13225,N_11845,N_9183);
nand U13226 (N_13226,N_11853,N_10241);
and U13227 (N_13227,N_10477,N_9557);
nor U13228 (N_13228,N_9666,N_9711);
nand U13229 (N_13229,N_10852,N_9321);
or U13230 (N_13230,N_11184,N_11822);
or U13231 (N_13231,N_9221,N_10593);
nor U13232 (N_13232,N_9932,N_9828);
nor U13233 (N_13233,N_10784,N_9174);
or U13234 (N_13234,N_10191,N_11350);
and U13235 (N_13235,N_10940,N_9515);
nor U13236 (N_13236,N_10622,N_10692);
and U13237 (N_13237,N_11256,N_11549);
or U13238 (N_13238,N_9830,N_11450);
or U13239 (N_13239,N_10465,N_10882);
nand U13240 (N_13240,N_10894,N_11082);
nand U13241 (N_13241,N_9506,N_9619);
or U13242 (N_13242,N_10378,N_11840);
or U13243 (N_13243,N_10431,N_10518);
nor U13244 (N_13244,N_10962,N_9142);
and U13245 (N_13245,N_11546,N_10164);
nor U13246 (N_13246,N_10815,N_10212);
nand U13247 (N_13247,N_10189,N_9074);
nor U13248 (N_13248,N_10483,N_9661);
nand U13249 (N_13249,N_10534,N_10407);
nand U13250 (N_13250,N_9979,N_10370);
and U13251 (N_13251,N_11747,N_9425);
or U13252 (N_13252,N_11860,N_10993);
nor U13253 (N_13253,N_9355,N_11716);
nor U13254 (N_13254,N_10587,N_11997);
or U13255 (N_13255,N_11501,N_10570);
or U13256 (N_13256,N_11735,N_10230);
nor U13257 (N_13257,N_11725,N_10729);
nand U13258 (N_13258,N_10652,N_11219);
or U13259 (N_13259,N_11382,N_9993);
nand U13260 (N_13260,N_11081,N_9271);
nand U13261 (N_13261,N_9043,N_11952);
nor U13262 (N_13262,N_10170,N_10495);
nand U13263 (N_13263,N_9857,N_11763);
and U13264 (N_13264,N_10355,N_11100);
and U13265 (N_13265,N_9171,N_10464);
nand U13266 (N_13266,N_11764,N_9829);
nor U13267 (N_13267,N_9176,N_9745);
or U13268 (N_13268,N_11542,N_10816);
or U13269 (N_13269,N_11369,N_9021);
nand U13270 (N_13270,N_10809,N_10186);
nor U13271 (N_13271,N_11830,N_9274);
nor U13272 (N_13272,N_10237,N_9025);
nand U13273 (N_13273,N_9918,N_9415);
xor U13274 (N_13274,N_10942,N_10671);
nand U13275 (N_13275,N_9602,N_10565);
xor U13276 (N_13276,N_10854,N_11994);
or U13277 (N_13277,N_9905,N_9514);
and U13278 (N_13278,N_10110,N_11323);
and U13279 (N_13279,N_10298,N_9768);
or U13280 (N_13280,N_11523,N_9210);
or U13281 (N_13281,N_10566,N_10408);
or U13282 (N_13282,N_9633,N_10257);
nor U13283 (N_13283,N_11031,N_9492);
nor U13284 (N_13284,N_10633,N_11816);
and U13285 (N_13285,N_10897,N_11643);
and U13286 (N_13286,N_10181,N_9463);
and U13287 (N_13287,N_11669,N_11014);
nor U13288 (N_13288,N_11992,N_9063);
and U13289 (N_13289,N_11847,N_10101);
nand U13290 (N_13290,N_11589,N_11083);
and U13291 (N_13291,N_9780,N_9149);
and U13292 (N_13292,N_10065,N_11538);
nand U13293 (N_13293,N_9489,N_11602);
and U13294 (N_13294,N_11073,N_9767);
and U13295 (N_13295,N_11736,N_11776);
or U13296 (N_13296,N_9146,N_11975);
or U13297 (N_13297,N_10931,N_9914);
nor U13298 (N_13298,N_9778,N_11632);
nor U13299 (N_13299,N_11322,N_10961);
or U13300 (N_13300,N_11268,N_9109);
and U13301 (N_13301,N_10670,N_10176);
nor U13302 (N_13302,N_10381,N_10240);
or U13303 (N_13303,N_9407,N_10022);
nand U13304 (N_13304,N_11395,N_9876);
nor U13305 (N_13305,N_9877,N_9085);
nand U13306 (N_13306,N_9000,N_9911);
and U13307 (N_13307,N_10745,N_11121);
or U13308 (N_13308,N_10042,N_10293);
nor U13309 (N_13309,N_11302,N_11275);
and U13310 (N_13310,N_10801,N_11164);
xor U13311 (N_13311,N_9664,N_10792);
nand U13312 (N_13312,N_11013,N_9494);
nand U13313 (N_13313,N_10539,N_11592);
and U13314 (N_13314,N_9377,N_9584);
nor U13315 (N_13315,N_11110,N_9418);
or U13316 (N_13316,N_10665,N_11876);
and U13317 (N_13317,N_10930,N_9643);
and U13318 (N_13318,N_11802,N_9776);
nor U13319 (N_13319,N_10756,N_9612);
or U13320 (N_13320,N_10105,N_9462);
nor U13321 (N_13321,N_10650,N_9035);
and U13322 (N_13322,N_9208,N_11804);
and U13323 (N_13323,N_9736,N_9301);
nand U13324 (N_13324,N_10333,N_9103);
and U13325 (N_13325,N_9984,N_11251);
and U13326 (N_13326,N_9233,N_11934);
and U13327 (N_13327,N_9796,N_10085);
nor U13328 (N_13328,N_11052,N_11397);
or U13329 (N_13329,N_9270,N_10029);
and U13330 (N_13330,N_9092,N_10718);
or U13331 (N_13331,N_10578,N_11564);
or U13332 (N_13332,N_10062,N_9894);
nor U13333 (N_13333,N_9624,N_11399);
nand U13334 (N_13334,N_9781,N_11867);
and U13335 (N_13335,N_10928,N_9945);
nand U13336 (N_13336,N_9373,N_10053);
nand U13337 (N_13337,N_10058,N_9133);
and U13338 (N_13338,N_11800,N_9341);
nand U13339 (N_13339,N_11539,N_10742);
xnor U13340 (N_13340,N_10699,N_10145);
xnor U13341 (N_13341,N_11333,N_10799);
or U13342 (N_13342,N_11252,N_10899);
nand U13343 (N_13343,N_10130,N_9438);
and U13344 (N_13344,N_10974,N_11908);
nor U13345 (N_13345,N_10969,N_9487);
or U13346 (N_13346,N_11585,N_11126);
nor U13347 (N_13347,N_11060,N_9812);
nand U13348 (N_13348,N_11291,N_9367);
and U13349 (N_13349,N_9507,N_10239);
and U13350 (N_13350,N_11600,N_10838);
nor U13351 (N_13351,N_10409,N_9193);
or U13352 (N_13352,N_9150,N_11582);
and U13353 (N_13353,N_10046,N_9702);
and U13354 (N_13354,N_9258,N_9500);
nor U13355 (N_13355,N_9826,N_9787);
nand U13356 (N_13356,N_11856,N_11191);
or U13357 (N_13357,N_10724,N_10086);
or U13358 (N_13358,N_11049,N_10807);
nand U13359 (N_13359,N_9986,N_10528);
nor U13360 (N_13360,N_11988,N_9263);
or U13361 (N_13361,N_9434,N_11671);
or U13362 (N_13362,N_9049,N_10107);
nor U13363 (N_13363,N_11390,N_10552);
xor U13364 (N_13364,N_11703,N_11712);
nor U13365 (N_13365,N_11651,N_9838);
and U13366 (N_13366,N_10773,N_9313);
or U13367 (N_13367,N_11838,N_10084);
or U13368 (N_13368,N_11661,N_9789);
or U13369 (N_13369,N_10417,N_9555);
and U13370 (N_13370,N_9427,N_9403);
and U13371 (N_13371,N_11088,N_10715);
nand U13372 (N_13372,N_10782,N_10762);
and U13373 (N_13373,N_10156,N_11578);
nand U13374 (N_13374,N_11125,N_10028);
nand U13375 (N_13375,N_11306,N_9588);
and U13376 (N_13376,N_9003,N_9595);
nor U13377 (N_13377,N_10577,N_10258);
nand U13378 (N_13378,N_9532,N_9908);
nand U13379 (N_13379,N_10166,N_9704);
or U13380 (N_13380,N_9942,N_9707);
or U13381 (N_13381,N_9242,N_9946);
nor U13382 (N_13382,N_11241,N_9559);
and U13383 (N_13383,N_11568,N_10510);
and U13384 (N_13384,N_9813,N_9127);
nor U13385 (N_13385,N_9659,N_9944);
nand U13386 (N_13386,N_9384,N_11370);
and U13387 (N_13387,N_9077,N_11283);
or U13388 (N_13388,N_11739,N_11560);
nor U13389 (N_13389,N_11215,N_9939);
or U13390 (N_13390,N_9832,N_11832);
and U13391 (N_13391,N_11176,N_11422);
and U13392 (N_13392,N_11939,N_11112);
and U13393 (N_13393,N_9717,N_9457);
nor U13394 (N_13394,N_9295,N_10103);
nor U13395 (N_13395,N_11915,N_10127);
and U13396 (N_13396,N_11678,N_9692);
or U13397 (N_13397,N_11475,N_9156);
nand U13398 (N_13398,N_11180,N_9535);
or U13399 (N_13399,N_9286,N_11174);
nor U13400 (N_13400,N_10324,N_11777);
nor U13401 (N_13401,N_11037,N_9909);
nor U13402 (N_13402,N_10979,N_11733);
nor U13403 (N_13403,N_10245,N_11468);
or U13404 (N_13404,N_10452,N_10519);
nand U13405 (N_13405,N_11696,N_11299);
nor U13406 (N_13406,N_9383,N_10133);
nor U13407 (N_13407,N_11371,N_10963);
or U13408 (N_13408,N_9587,N_9006);
or U13409 (N_13409,N_11755,N_10354);
or U13410 (N_13410,N_10878,N_10353);
or U13411 (N_13411,N_10259,N_10325);
and U13412 (N_13412,N_11530,N_9188);
and U13413 (N_13413,N_9419,N_10842);
and U13414 (N_13414,N_9972,N_11281);
nand U13415 (N_13415,N_9963,N_10614);
nand U13416 (N_13416,N_10322,N_11348);
or U13417 (N_13417,N_9548,N_11172);
or U13418 (N_13418,N_10751,N_11699);
nor U13419 (N_13419,N_10135,N_11340);
or U13420 (N_13420,N_11070,N_10513);
nor U13421 (N_13421,N_9037,N_10705);
and U13422 (N_13422,N_11531,N_11987);
nand U13423 (N_13423,N_10769,N_11714);
nor U13424 (N_13424,N_11018,N_10019);
nand U13425 (N_13425,N_9040,N_11063);
nor U13426 (N_13426,N_10533,N_9888);
nor U13427 (N_13427,N_10337,N_9264);
nand U13428 (N_13428,N_10162,N_10021);
and U13429 (N_13429,N_11160,N_9509);
and U13430 (N_13430,N_9610,N_10701);
nor U13431 (N_13431,N_11967,N_11111);
nor U13432 (N_13432,N_11067,N_10057);
nand U13433 (N_13433,N_9658,N_10342);
and U13434 (N_13434,N_11332,N_10772);
nand U13435 (N_13435,N_9112,N_9053);
and U13436 (N_13436,N_9850,N_11803);
or U13437 (N_13437,N_11116,N_11601);
nand U13438 (N_13438,N_10244,N_11744);
nand U13439 (N_13439,N_10826,N_10037);
and U13440 (N_13440,N_11953,N_11364);
or U13441 (N_13441,N_10933,N_9499);
nand U13442 (N_13442,N_11094,N_10787);
and U13443 (N_13443,N_9741,N_10771);
and U13444 (N_13444,N_10082,N_11891);
nand U13445 (N_13445,N_11262,N_9536);
or U13446 (N_13446,N_9771,N_11504);
nand U13447 (N_13447,N_11836,N_9860);
nor U13448 (N_13448,N_11434,N_9547);
nand U13449 (N_13449,N_10466,N_9718);
nor U13450 (N_13450,N_9364,N_10304);
and U13451 (N_13451,N_10410,N_11133);
or U13452 (N_13452,N_11513,N_10003);
nor U13453 (N_13453,N_10919,N_9422);
and U13454 (N_13454,N_10596,N_10220);
nor U13455 (N_13455,N_9570,N_10835);
or U13456 (N_13456,N_11175,N_9907);
or U13457 (N_13457,N_10615,N_10817);
and U13458 (N_13458,N_10783,N_10069);
nor U13459 (N_13459,N_9433,N_10160);
nand U13460 (N_13460,N_11896,N_10419);
nand U13461 (N_13461,N_9696,N_10900);
nor U13462 (N_13462,N_9190,N_11644);
or U13463 (N_13463,N_11039,N_10877);
and U13464 (N_13464,N_11898,N_10051);
nand U13465 (N_13465,N_10923,N_10798);
or U13466 (N_13466,N_11603,N_9097);
nand U13467 (N_13467,N_9192,N_11454);
nor U13468 (N_13468,N_11942,N_10898);
or U13469 (N_13469,N_10229,N_9060);
nor U13470 (N_13470,N_11947,N_11305);
and U13471 (N_13471,N_10393,N_11799);
nand U13472 (N_13472,N_11113,N_11943);
and U13473 (N_13473,N_9592,N_9267);
or U13474 (N_13474,N_10268,N_11463);
or U13475 (N_13475,N_10208,N_10975);
nand U13476 (N_13476,N_10638,N_10184);
xnor U13477 (N_13477,N_9839,N_9523);
nand U13478 (N_13478,N_11069,N_9230);
nor U13479 (N_13479,N_10484,N_10117);
or U13480 (N_13480,N_10302,N_9456);
nand U13481 (N_13481,N_10193,N_11825);
or U13482 (N_13482,N_10662,N_9145);
and U13483 (N_13483,N_11359,N_9691);
or U13484 (N_13484,N_9479,N_10017);
or U13485 (N_13485,N_9769,N_11277);
and U13486 (N_13486,N_11808,N_9248);
nor U13487 (N_13487,N_11779,N_9465);
nor U13488 (N_13488,N_11555,N_11266);
nand U13489 (N_13489,N_9722,N_11554);
nor U13490 (N_13490,N_9609,N_9452);
nor U13491 (N_13491,N_9019,N_10214);
nand U13492 (N_13492,N_11461,N_11326);
or U13493 (N_13493,N_10906,N_9822);
and U13494 (N_13494,N_10020,N_11767);
nor U13495 (N_13495,N_10031,N_11462);
and U13496 (N_13496,N_9635,N_9521);
nand U13497 (N_13497,N_11647,N_10859);
or U13498 (N_13498,N_11106,N_10418);
or U13499 (N_13499,N_9516,N_11412);
and U13500 (N_13500,N_9441,N_11515);
and U13501 (N_13501,N_10929,N_11135);
or U13502 (N_13502,N_11113,N_10053);
nor U13503 (N_13503,N_10896,N_11917);
and U13504 (N_13504,N_9093,N_9770);
nor U13505 (N_13505,N_9773,N_9892);
or U13506 (N_13506,N_9444,N_11038);
nor U13507 (N_13507,N_10990,N_11155);
and U13508 (N_13508,N_9097,N_10274);
and U13509 (N_13509,N_11146,N_10498);
or U13510 (N_13510,N_11798,N_9807);
nor U13511 (N_13511,N_11683,N_11692);
nand U13512 (N_13512,N_9183,N_10429);
nor U13513 (N_13513,N_10040,N_11352);
nand U13514 (N_13514,N_11912,N_11697);
and U13515 (N_13515,N_10099,N_9010);
nor U13516 (N_13516,N_9688,N_11099);
and U13517 (N_13517,N_11503,N_9052);
or U13518 (N_13518,N_11880,N_9933);
and U13519 (N_13519,N_10107,N_11050);
or U13520 (N_13520,N_9599,N_11950);
or U13521 (N_13521,N_10283,N_10992);
nor U13522 (N_13522,N_11470,N_10735);
and U13523 (N_13523,N_10743,N_11008);
nor U13524 (N_13524,N_9704,N_11701);
nor U13525 (N_13525,N_11737,N_11463);
or U13526 (N_13526,N_11180,N_10726);
or U13527 (N_13527,N_9475,N_10868);
or U13528 (N_13528,N_11312,N_9692);
nand U13529 (N_13529,N_10219,N_9624);
nand U13530 (N_13530,N_9879,N_10638);
nor U13531 (N_13531,N_11684,N_10722);
or U13532 (N_13532,N_9338,N_11937);
and U13533 (N_13533,N_10276,N_10834);
nor U13534 (N_13534,N_11502,N_11513);
or U13535 (N_13535,N_9949,N_11502);
or U13536 (N_13536,N_9382,N_11937);
nor U13537 (N_13537,N_9782,N_10542);
or U13538 (N_13538,N_9889,N_10920);
nor U13539 (N_13539,N_11331,N_11127);
nor U13540 (N_13540,N_11683,N_9505);
or U13541 (N_13541,N_11885,N_9214);
nor U13542 (N_13542,N_9124,N_10893);
nand U13543 (N_13543,N_9661,N_10467);
or U13544 (N_13544,N_9661,N_9808);
or U13545 (N_13545,N_11469,N_10646);
nand U13546 (N_13546,N_9110,N_11519);
or U13547 (N_13547,N_11817,N_10790);
or U13548 (N_13548,N_9367,N_9286);
nand U13549 (N_13549,N_11755,N_11480);
nand U13550 (N_13550,N_10395,N_9847);
or U13551 (N_13551,N_11765,N_10342);
nand U13552 (N_13552,N_11718,N_9668);
and U13553 (N_13553,N_10259,N_11538);
nand U13554 (N_13554,N_11166,N_10108);
and U13555 (N_13555,N_11738,N_11045);
nor U13556 (N_13556,N_9316,N_11369);
and U13557 (N_13557,N_9438,N_11941);
or U13558 (N_13558,N_9735,N_11370);
nor U13559 (N_13559,N_9521,N_10508);
and U13560 (N_13560,N_11250,N_10448);
or U13561 (N_13561,N_10087,N_11558);
nand U13562 (N_13562,N_9766,N_10250);
or U13563 (N_13563,N_10508,N_9713);
and U13564 (N_13564,N_11203,N_11388);
nor U13565 (N_13565,N_11245,N_9705);
and U13566 (N_13566,N_10324,N_10918);
nand U13567 (N_13567,N_9291,N_10099);
and U13568 (N_13568,N_11274,N_11644);
nand U13569 (N_13569,N_11646,N_10477);
or U13570 (N_13570,N_11237,N_9642);
or U13571 (N_13571,N_9754,N_10206);
nor U13572 (N_13572,N_11476,N_10370);
nand U13573 (N_13573,N_9201,N_10556);
nor U13574 (N_13574,N_10847,N_9220);
nor U13575 (N_13575,N_11929,N_10646);
and U13576 (N_13576,N_10054,N_10120);
nor U13577 (N_13577,N_10316,N_9591);
and U13578 (N_13578,N_11963,N_11208);
nor U13579 (N_13579,N_11255,N_10862);
or U13580 (N_13580,N_10794,N_10769);
and U13581 (N_13581,N_10059,N_11084);
nor U13582 (N_13582,N_11116,N_9997);
nor U13583 (N_13583,N_10334,N_9837);
or U13584 (N_13584,N_10106,N_11205);
xor U13585 (N_13585,N_11887,N_10138);
or U13586 (N_13586,N_9736,N_11062);
and U13587 (N_13587,N_10067,N_11336);
nand U13588 (N_13588,N_11506,N_9949);
nand U13589 (N_13589,N_9839,N_9193);
nand U13590 (N_13590,N_9260,N_9417);
xor U13591 (N_13591,N_9995,N_11433);
nor U13592 (N_13592,N_10090,N_11377);
nand U13593 (N_13593,N_9198,N_9685);
nor U13594 (N_13594,N_9028,N_9635);
and U13595 (N_13595,N_10048,N_10428);
nor U13596 (N_13596,N_10804,N_10286);
and U13597 (N_13597,N_10633,N_11879);
nand U13598 (N_13598,N_9858,N_11967);
and U13599 (N_13599,N_10038,N_11636);
or U13600 (N_13600,N_11169,N_10485);
or U13601 (N_13601,N_9291,N_10266);
nor U13602 (N_13602,N_10324,N_11733);
nor U13603 (N_13603,N_11874,N_10495);
nor U13604 (N_13604,N_9243,N_11956);
or U13605 (N_13605,N_10843,N_10410);
nor U13606 (N_13606,N_10706,N_11301);
nand U13607 (N_13607,N_11834,N_10187);
and U13608 (N_13608,N_10543,N_11210);
nand U13609 (N_13609,N_9501,N_10854);
nor U13610 (N_13610,N_10983,N_11225);
nor U13611 (N_13611,N_11229,N_10051);
and U13612 (N_13612,N_11614,N_10604);
and U13613 (N_13613,N_10387,N_11496);
and U13614 (N_13614,N_10376,N_10408);
and U13615 (N_13615,N_9474,N_11988);
and U13616 (N_13616,N_11482,N_10281);
or U13617 (N_13617,N_9306,N_11505);
nor U13618 (N_13618,N_9475,N_10230);
or U13619 (N_13619,N_10208,N_9750);
nand U13620 (N_13620,N_10941,N_9952);
nor U13621 (N_13621,N_10421,N_9461);
nor U13622 (N_13622,N_10219,N_11846);
nor U13623 (N_13623,N_11733,N_11700);
nand U13624 (N_13624,N_10538,N_11261);
xnor U13625 (N_13625,N_9101,N_9449);
or U13626 (N_13626,N_9771,N_11048);
nand U13627 (N_13627,N_10304,N_10045);
and U13628 (N_13628,N_9044,N_10395);
and U13629 (N_13629,N_11190,N_11359);
nand U13630 (N_13630,N_10562,N_9868);
nand U13631 (N_13631,N_11316,N_9505);
and U13632 (N_13632,N_11294,N_9626);
or U13633 (N_13633,N_11915,N_11280);
nor U13634 (N_13634,N_9729,N_11961);
nor U13635 (N_13635,N_9699,N_11068);
nand U13636 (N_13636,N_10866,N_9336);
nand U13637 (N_13637,N_9060,N_9989);
or U13638 (N_13638,N_10162,N_10768);
nand U13639 (N_13639,N_11670,N_10560);
or U13640 (N_13640,N_10681,N_9842);
nand U13641 (N_13641,N_10821,N_9962);
nor U13642 (N_13642,N_9378,N_10092);
or U13643 (N_13643,N_9648,N_9982);
xnor U13644 (N_13644,N_10024,N_9819);
and U13645 (N_13645,N_9198,N_10123);
and U13646 (N_13646,N_9618,N_9111);
and U13647 (N_13647,N_11636,N_11019);
nand U13648 (N_13648,N_10766,N_9769);
and U13649 (N_13649,N_10055,N_10320);
or U13650 (N_13650,N_11733,N_11713);
or U13651 (N_13651,N_9576,N_11694);
nor U13652 (N_13652,N_9000,N_9283);
nand U13653 (N_13653,N_9081,N_10255);
nand U13654 (N_13654,N_9848,N_11010);
or U13655 (N_13655,N_10882,N_9130);
nand U13656 (N_13656,N_10600,N_11294);
and U13657 (N_13657,N_9602,N_9566);
nand U13658 (N_13658,N_9006,N_10822);
and U13659 (N_13659,N_9032,N_11282);
and U13660 (N_13660,N_11454,N_11260);
or U13661 (N_13661,N_10979,N_11957);
nor U13662 (N_13662,N_9825,N_11422);
nor U13663 (N_13663,N_9941,N_9900);
nor U13664 (N_13664,N_10507,N_10123);
and U13665 (N_13665,N_10985,N_10281);
nand U13666 (N_13666,N_10306,N_10279);
nor U13667 (N_13667,N_10754,N_11560);
nand U13668 (N_13668,N_9553,N_11987);
and U13669 (N_13669,N_10281,N_11099);
nand U13670 (N_13670,N_9824,N_11046);
nand U13671 (N_13671,N_9884,N_10641);
or U13672 (N_13672,N_10997,N_10553);
or U13673 (N_13673,N_11638,N_9913);
nor U13674 (N_13674,N_9452,N_9115);
nor U13675 (N_13675,N_11336,N_10540);
nor U13676 (N_13676,N_9902,N_9529);
or U13677 (N_13677,N_10449,N_9279);
or U13678 (N_13678,N_9368,N_9868);
nand U13679 (N_13679,N_11395,N_10520);
nor U13680 (N_13680,N_9515,N_10470);
nor U13681 (N_13681,N_9499,N_10531);
or U13682 (N_13682,N_11960,N_10749);
or U13683 (N_13683,N_11563,N_11355);
nand U13684 (N_13684,N_9348,N_9699);
and U13685 (N_13685,N_11106,N_11768);
or U13686 (N_13686,N_11196,N_9633);
nor U13687 (N_13687,N_9087,N_9693);
or U13688 (N_13688,N_9330,N_10956);
nand U13689 (N_13689,N_10063,N_9816);
and U13690 (N_13690,N_9458,N_10436);
nor U13691 (N_13691,N_10269,N_9744);
nand U13692 (N_13692,N_9370,N_10481);
or U13693 (N_13693,N_10373,N_10436);
nor U13694 (N_13694,N_11280,N_10235);
and U13695 (N_13695,N_9043,N_9894);
nand U13696 (N_13696,N_11236,N_9105);
or U13697 (N_13697,N_11496,N_11850);
nand U13698 (N_13698,N_11229,N_10503);
nand U13699 (N_13699,N_11086,N_9248);
nand U13700 (N_13700,N_10606,N_9851);
and U13701 (N_13701,N_9451,N_10726);
and U13702 (N_13702,N_11808,N_9587);
nor U13703 (N_13703,N_10147,N_11790);
nor U13704 (N_13704,N_11183,N_10246);
nand U13705 (N_13705,N_11183,N_11914);
nor U13706 (N_13706,N_11958,N_10285);
nand U13707 (N_13707,N_11552,N_10162);
or U13708 (N_13708,N_11879,N_11396);
or U13709 (N_13709,N_9629,N_11924);
or U13710 (N_13710,N_10767,N_9817);
nand U13711 (N_13711,N_11795,N_10859);
and U13712 (N_13712,N_10340,N_9696);
nor U13713 (N_13713,N_9939,N_9682);
and U13714 (N_13714,N_11675,N_11114);
or U13715 (N_13715,N_11366,N_9653);
or U13716 (N_13716,N_11411,N_11965);
nor U13717 (N_13717,N_11679,N_10368);
nor U13718 (N_13718,N_11953,N_9936);
and U13719 (N_13719,N_9360,N_9038);
nand U13720 (N_13720,N_10571,N_9794);
and U13721 (N_13721,N_9048,N_9774);
or U13722 (N_13722,N_9498,N_11897);
or U13723 (N_13723,N_9619,N_11421);
and U13724 (N_13724,N_9731,N_11866);
nand U13725 (N_13725,N_10512,N_9804);
or U13726 (N_13726,N_11433,N_10908);
nor U13727 (N_13727,N_10412,N_11534);
nand U13728 (N_13728,N_11824,N_9590);
or U13729 (N_13729,N_11765,N_11028);
and U13730 (N_13730,N_9574,N_10972);
nor U13731 (N_13731,N_11372,N_9379);
nor U13732 (N_13732,N_11173,N_10312);
nor U13733 (N_13733,N_11383,N_10080);
or U13734 (N_13734,N_9382,N_10156);
or U13735 (N_13735,N_11029,N_11166);
nor U13736 (N_13736,N_10542,N_11885);
or U13737 (N_13737,N_9912,N_10575);
and U13738 (N_13738,N_9121,N_11180);
and U13739 (N_13739,N_9522,N_9445);
nand U13740 (N_13740,N_9361,N_10954);
nand U13741 (N_13741,N_11159,N_10363);
nand U13742 (N_13742,N_9866,N_10136);
and U13743 (N_13743,N_9008,N_10867);
and U13744 (N_13744,N_9490,N_10271);
nor U13745 (N_13745,N_11631,N_10693);
nand U13746 (N_13746,N_10055,N_9087);
nor U13747 (N_13747,N_9488,N_10929);
nor U13748 (N_13748,N_11520,N_11926);
nor U13749 (N_13749,N_9837,N_10551);
nor U13750 (N_13750,N_9827,N_11730);
nand U13751 (N_13751,N_11830,N_10886);
or U13752 (N_13752,N_10054,N_11714);
nand U13753 (N_13753,N_10893,N_11486);
nand U13754 (N_13754,N_9271,N_11266);
and U13755 (N_13755,N_11592,N_10669);
or U13756 (N_13756,N_11112,N_10162);
nand U13757 (N_13757,N_11448,N_9005);
or U13758 (N_13758,N_11298,N_9764);
nand U13759 (N_13759,N_11722,N_10414);
and U13760 (N_13760,N_11468,N_10907);
nor U13761 (N_13761,N_9052,N_9057);
and U13762 (N_13762,N_9790,N_11202);
or U13763 (N_13763,N_10989,N_9059);
and U13764 (N_13764,N_10129,N_10520);
nor U13765 (N_13765,N_11328,N_11197);
and U13766 (N_13766,N_10018,N_10492);
nor U13767 (N_13767,N_9922,N_9658);
nand U13768 (N_13768,N_11960,N_9140);
nand U13769 (N_13769,N_11115,N_9553);
nor U13770 (N_13770,N_10221,N_10508);
and U13771 (N_13771,N_9842,N_10207);
and U13772 (N_13772,N_9570,N_10448);
nor U13773 (N_13773,N_10669,N_10020);
and U13774 (N_13774,N_11609,N_9268);
nand U13775 (N_13775,N_11185,N_9338);
nor U13776 (N_13776,N_9489,N_10764);
nor U13777 (N_13777,N_9393,N_11276);
nand U13778 (N_13778,N_11640,N_11200);
nand U13779 (N_13779,N_10406,N_10629);
or U13780 (N_13780,N_9921,N_9653);
nand U13781 (N_13781,N_10386,N_11106);
nor U13782 (N_13782,N_10218,N_11982);
or U13783 (N_13783,N_10607,N_9342);
nor U13784 (N_13784,N_11597,N_11572);
nor U13785 (N_13785,N_11592,N_10186);
and U13786 (N_13786,N_10155,N_9507);
and U13787 (N_13787,N_9189,N_11580);
or U13788 (N_13788,N_10929,N_10022);
nor U13789 (N_13789,N_11771,N_11700);
and U13790 (N_13790,N_10853,N_10563);
nor U13791 (N_13791,N_11682,N_11901);
or U13792 (N_13792,N_9503,N_9188);
nor U13793 (N_13793,N_11421,N_9422);
nor U13794 (N_13794,N_11604,N_9894);
or U13795 (N_13795,N_9785,N_9190);
and U13796 (N_13796,N_11469,N_9614);
and U13797 (N_13797,N_11633,N_9876);
or U13798 (N_13798,N_10205,N_11164);
nor U13799 (N_13799,N_10535,N_10423);
and U13800 (N_13800,N_11025,N_10840);
and U13801 (N_13801,N_9560,N_11068);
and U13802 (N_13802,N_9061,N_9755);
and U13803 (N_13803,N_10067,N_11578);
and U13804 (N_13804,N_11780,N_9004);
and U13805 (N_13805,N_11055,N_9428);
nor U13806 (N_13806,N_10962,N_10126);
or U13807 (N_13807,N_10740,N_10896);
nor U13808 (N_13808,N_11471,N_11355);
and U13809 (N_13809,N_11227,N_11908);
and U13810 (N_13810,N_11634,N_9233);
or U13811 (N_13811,N_9824,N_10891);
or U13812 (N_13812,N_11265,N_9848);
nand U13813 (N_13813,N_10858,N_11152);
and U13814 (N_13814,N_10385,N_11530);
nor U13815 (N_13815,N_9345,N_9476);
nor U13816 (N_13816,N_10614,N_10271);
and U13817 (N_13817,N_11999,N_9874);
nand U13818 (N_13818,N_10033,N_9150);
nor U13819 (N_13819,N_10565,N_10525);
nand U13820 (N_13820,N_9065,N_10381);
and U13821 (N_13821,N_11782,N_11848);
or U13822 (N_13822,N_9561,N_10465);
or U13823 (N_13823,N_9809,N_10437);
nor U13824 (N_13824,N_10394,N_10800);
or U13825 (N_13825,N_10719,N_10016);
xor U13826 (N_13826,N_10419,N_10908);
and U13827 (N_13827,N_10997,N_9844);
or U13828 (N_13828,N_9935,N_10104);
and U13829 (N_13829,N_11052,N_10080);
nand U13830 (N_13830,N_10545,N_10080);
nand U13831 (N_13831,N_11184,N_11382);
and U13832 (N_13832,N_10146,N_10177);
nor U13833 (N_13833,N_11750,N_9208);
nand U13834 (N_13834,N_9250,N_10554);
and U13835 (N_13835,N_10452,N_9583);
and U13836 (N_13836,N_9402,N_10797);
or U13837 (N_13837,N_9300,N_9611);
and U13838 (N_13838,N_11335,N_9488);
or U13839 (N_13839,N_9596,N_9149);
xor U13840 (N_13840,N_9662,N_11968);
nor U13841 (N_13841,N_9619,N_9565);
nand U13842 (N_13842,N_10321,N_9419);
and U13843 (N_13843,N_10277,N_10093);
nor U13844 (N_13844,N_10290,N_10208);
nand U13845 (N_13845,N_10592,N_9640);
and U13846 (N_13846,N_11435,N_9143);
or U13847 (N_13847,N_9806,N_10541);
xor U13848 (N_13848,N_11418,N_9427);
or U13849 (N_13849,N_10763,N_10932);
nor U13850 (N_13850,N_9971,N_11354);
and U13851 (N_13851,N_9451,N_10164);
nor U13852 (N_13852,N_10852,N_10298);
or U13853 (N_13853,N_11447,N_10082);
and U13854 (N_13854,N_11809,N_9974);
nand U13855 (N_13855,N_10859,N_11154);
or U13856 (N_13856,N_11684,N_11947);
or U13857 (N_13857,N_10321,N_9544);
nand U13858 (N_13858,N_10341,N_10918);
and U13859 (N_13859,N_11482,N_11072);
nor U13860 (N_13860,N_11647,N_9932);
or U13861 (N_13861,N_10885,N_9727);
nand U13862 (N_13862,N_9609,N_11927);
or U13863 (N_13863,N_11045,N_9685);
nor U13864 (N_13864,N_9179,N_11664);
nand U13865 (N_13865,N_9907,N_9369);
and U13866 (N_13866,N_10800,N_11395);
or U13867 (N_13867,N_10416,N_9596);
and U13868 (N_13868,N_11788,N_9552);
or U13869 (N_13869,N_10800,N_10086);
and U13870 (N_13870,N_10538,N_9695);
or U13871 (N_13871,N_10126,N_9839);
nand U13872 (N_13872,N_10118,N_11741);
nor U13873 (N_13873,N_11863,N_10606);
nand U13874 (N_13874,N_10998,N_9397);
or U13875 (N_13875,N_11084,N_10023);
or U13876 (N_13876,N_10821,N_10235);
or U13877 (N_13877,N_9932,N_10287);
nand U13878 (N_13878,N_9917,N_11164);
and U13879 (N_13879,N_9668,N_11564);
nor U13880 (N_13880,N_9616,N_10062);
and U13881 (N_13881,N_11182,N_10842);
and U13882 (N_13882,N_9358,N_10660);
or U13883 (N_13883,N_9306,N_9349);
nand U13884 (N_13884,N_11134,N_10857);
and U13885 (N_13885,N_11009,N_10106);
or U13886 (N_13886,N_11080,N_11376);
or U13887 (N_13887,N_9729,N_9376);
or U13888 (N_13888,N_9286,N_10211);
nand U13889 (N_13889,N_9530,N_9208);
nor U13890 (N_13890,N_9787,N_10451);
or U13891 (N_13891,N_11723,N_11879);
or U13892 (N_13892,N_11392,N_10953);
and U13893 (N_13893,N_9082,N_11100);
nor U13894 (N_13894,N_10612,N_11252);
or U13895 (N_13895,N_10254,N_9841);
and U13896 (N_13896,N_10227,N_11610);
nand U13897 (N_13897,N_9459,N_11930);
or U13898 (N_13898,N_9681,N_9731);
nor U13899 (N_13899,N_11752,N_11870);
and U13900 (N_13900,N_11527,N_11922);
nand U13901 (N_13901,N_10211,N_9110);
nand U13902 (N_13902,N_10214,N_9021);
or U13903 (N_13903,N_11236,N_11553);
and U13904 (N_13904,N_10944,N_9967);
or U13905 (N_13905,N_9761,N_9118);
or U13906 (N_13906,N_10290,N_11839);
or U13907 (N_13907,N_11893,N_9064);
nor U13908 (N_13908,N_11030,N_11796);
or U13909 (N_13909,N_11797,N_10241);
nand U13910 (N_13910,N_11823,N_10912);
nand U13911 (N_13911,N_10651,N_10300);
nand U13912 (N_13912,N_9284,N_11083);
nand U13913 (N_13913,N_11616,N_10206);
and U13914 (N_13914,N_11372,N_11341);
and U13915 (N_13915,N_11532,N_9763);
nor U13916 (N_13916,N_11250,N_11730);
and U13917 (N_13917,N_11262,N_11412);
and U13918 (N_13918,N_11316,N_11794);
or U13919 (N_13919,N_11195,N_9387);
nor U13920 (N_13920,N_9426,N_11339);
nor U13921 (N_13921,N_11863,N_10348);
xor U13922 (N_13922,N_11760,N_11200);
or U13923 (N_13923,N_10395,N_11640);
and U13924 (N_13924,N_11906,N_10870);
or U13925 (N_13925,N_11477,N_11159);
nand U13926 (N_13926,N_11207,N_11252);
and U13927 (N_13927,N_9565,N_9085);
nand U13928 (N_13928,N_11432,N_11940);
or U13929 (N_13929,N_10671,N_11755);
and U13930 (N_13930,N_11444,N_9933);
nor U13931 (N_13931,N_9420,N_10913);
or U13932 (N_13932,N_9186,N_10685);
and U13933 (N_13933,N_10321,N_9910);
and U13934 (N_13934,N_11673,N_11272);
nand U13935 (N_13935,N_9212,N_9217);
nor U13936 (N_13936,N_9234,N_11381);
nand U13937 (N_13937,N_11456,N_9866);
nor U13938 (N_13938,N_11846,N_9110);
nor U13939 (N_13939,N_10756,N_11230);
and U13940 (N_13940,N_9944,N_10025);
and U13941 (N_13941,N_10833,N_11349);
nand U13942 (N_13942,N_11679,N_10635);
or U13943 (N_13943,N_11184,N_9183);
nand U13944 (N_13944,N_9256,N_9250);
nor U13945 (N_13945,N_9727,N_11317);
nand U13946 (N_13946,N_11154,N_9980);
or U13947 (N_13947,N_10910,N_9199);
or U13948 (N_13948,N_11818,N_9730);
nand U13949 (N_13949,N_9891,N_10159);
and U13950 (N_13950,N_11271,N_11227);
or U13951 (N_13951,N_11956,N_10140);
and U13952 (N_13952,N_11847,N_11149);
or U13953 (N_13953,N_9317,N_9060);
nor U13954 (N_13954,N_10141,N_11383);
nor U13955 (N_13955,N_10348,N_9599);
or U13956 (N_13956,N_10521,N_11727);
nand U13957 (N_13957,N_9865,N_10337);
and U13958 (N_13958,N_9412,N_10160);
and U13959 (N_13959,N_9648,N_9595);
and U13960 (N_13960,N_9784,N_11491);
nor U13961 (N_13961,N_9818,N_11666);
and U13962 (N_13962,N_9136,N_11161);
and U13963 (N_13963,N_9618,N_10534);
nand U13964 (N_13964,N_10060,N_9738);
and U13965 (N_13965,N_9119,N_11014);
and U13966 (N_13966,N_10563,N_11591);
and U13967 (N_13967,N_9847,N_10043);
nor U13968 (N_13968,N_11127,N_11581);
nor U13969 (N_13969,N_10754,N_11354);
nor U13970 (N_13970,N_10760,N_11710);
nand U13971 (N_13971,N_10944,N_10785);
nor U13972 (N_13972,N_9536,N_11800);
nand U13973 (N_13973,N_10057,N_10092);
nor U13974 (N_13974,N_10128,N_11995);
or U13975 (N_13975,N_9605,N_11253);
nor U13976 (N_13976,N_9555,N_11294);
or U13977 (N_13977,N_10234,N_10435);
nor U13978 (N_13978,N_10788,N_9937);
and U13979 (N_13979,N_11773,N_11824);
nor U13980 (N_13980,N_9036,N_10083);
nor U13981 (N_13981,N_9775,N_9014);
nand U13982 (N_13982,N_11842,N_9254);
nand U13983 (N_13983,N_11837,N_10625);
nor U13984 (N_13984,N_11674,N_9782);
or U13985 (N_13985,N_9387,N_11951);
or U13986 (N_13986,N_11082,N_10122);
or U13987 (N_13987,N_9296,N_10712);
nor U13988 (N_13988,N_9216,N_11687);
nor U13989 (N_13989,N_11091,N_9307);
nand U13990 (N_13990,N_10006,N_9881);
nand U13991 (N_13991,N_10437,N_11365);
nor U13992 (N_13992,N_10395,N_10772);
nor U13993 (N_13993,N_10355,N_10542);
or U13994 (N_13994,N_9058,N_9315);
or U13995 (N_13995,N_9159,N_9481);
and U13996 (N_13996,N_10782,N_11189);
nand U13997 (N_13997,N_9230,N_11300);
nand U13998 (N_13998,N_10835,N_11512);
xnor U13999 (N_13999,N_10020,N_9620);
nor U14000 (N_14000,N_10195,N_9371);
and U14001 (N_14001,N_11020,N_11986);
or U14002 (N_14002,N_11538,N_10473);
and U14003 (N_14003,N_10213,N_11406);
nand U14004 (N_14004,N_9625,N_11803);
nand U14005 (N_14005,N_10047,N_11355);
nor U14006 (N_14006,N_11865,N_11636);
nor U14007 (N_14007,N_9076,N_11130);
nand U14008 (N_14008,N_11720,N_11170);
or U14009 (N_14009,N_10838,N_10571);
nor U14010 (N_14010,N_10914,N_11346);
or U14011 (N_14011,N_10575,N_11339);
xor U14012 (N_14012,N_10200,N_9042);
nor U14013 (N_14013,N_9396,N_11075);
or U14014 (N_14014,N_11679,N_11574);
nand U14015 (N_14015,N_11905,N_9629);
or U14016 (N_14016,N_11942,N_10764);
or U14017 (N_14017,N_10228,N_9397);
and U14018 (N_14018,N_11509,N_11906);
nand U14019 (N_14019,N_10721,N_10287);
or U14020 (N_14020,N_10184,N_11284);
and U14021 (N_14021,N_10314,N_10810);
nor U14022 (N_14022,N_9297,N_11495);
and U14023 (N_14023,N_11495,N_9159);
or U14024 (N_14024,N_9742,N_9354);
and U14025 (N_14025,N_9788,N_9298);
and U14026 (N_14026,N_11361,N_10838);
and U14027 (N_14027,N_10452,N_10083);
and U14028 (N_14028,N_9950,N_10920);
or U14029 (N_14029,N_11509,N_10768);
nand U14030 (N_14030,N_11286,N_10191);
nand U14031 (N_14031,N_9755,N_9255);
or U14032 (N_14032,N_9138,N_9363);
and U14033 (N_14033,N_11246,N_9791);
nand U14034 (N_14034,N_10376,N_11564);
and U14035 (N_14035,N_9034,N_9794);
nor U14036 (N_14036,N_10566,N_11417);
nor U14037 (N_14037,N_10353,N_11617);
and U14038 (N_14038,N_11802,N_9954);
and U14039 (N_14039,N_10286,N_10748);
or U14040 (N_14040,N_11135,N_11283);
or U14041 (N_14041,N_10839,N_10000);
and U14042 (N_14042,N_9418,N_9910);
nand U14043 (N_14043,N_11058,N_11257);
and U14044 (N_14044,N_10259,N_11386);
or U14045 (N_14045,N_9220,N_10928);
and U14046 (N_14046,N_9203,N_10704);
nand U14047 (N_14047,N_10131,N_9357);
or U14048 (N_14048,N_9596,N_11064);
or U14049 (N_14049,N_11854,N_9413);
nor U14050 (N_14050,N_10254,N_11642);
nor U14051 (N_14051,N_9981,N_11316);
nor U14052 (N_14052,N_10099,N_10487);
nor U14053 (N_14053,N_9070,N_10952);
and U14054 (N_14054,N_9572,N_11558);
nand U14055 (N_14055,N_9247,N_9777);
nor U14056 (N_14056,N_10171,N_11867);
and U14057 (N_14057,N_11608,N_9660);
nor U14058 (N_14058,N_11282,N_10401);
nand U14059 (N_14059,N_10749,N_10760);
or U14060 (N_14060,N_9341,N_10774);
and U14061 (N_14061,N_11464,N_10246);
nand U14062 (N_14062,N_11878,N_9515);
nor U14063 (N_14063,N_9618,N_10366);
or U14064 (N_14064,N_10630,N_9616);
nor U14065 (N_14065,N_11300,N_11071);
nor U14066 (N_14066,N_11034,N_9881);
nor U14067 (N_14067,N_11035,N_9753);
or U14068 (N_14068,N_10663,N_10078);
and U14069 (N_14069,N_11833,N_9630);
xor U14070 (N_14070,N_9113,N_9815);
nand U14071 (N_14071,N_10084,N_11197);
nor U14072 (N_14072,N_10374,N_11605);
and U14073 (N_14073,N_11673,N_9530);
nor U14074 (N_14074,N_11700,N_9134);
nor U14075 (N_14075,N_11658,N_11979);
nor U14076 (N_14076,N_9088,N_10323);
nor U14077 (N_14077,N_9284,N_11819);
nand U14078 (N_14078,N_11448,N_10141);
nand U14079 (N_14079,N_10322,N_10617);
nand U14080 (N_14080,N_9831,N_9296);
and U14081 (N_14081,N_11498,N_9127);
or U14082 (N_14082,N_9192,N_11964);
and U14083 (N_14083,N_9855,N_11202);
nor U14084 (N_14084,N_9635,N_9190);
nand U14085 (N_14085,N_10184,N_10853);
and U14086 (N_14086,N_9258,N_11906);
and U14087 (N_14087,N_10844,N_10777);
nor U14088 (N_14088,N_9243,N_11363);
or U14089 (N_14089,N_9660,N_9675);
and U14090 (N_14090,N_9381,N_9603);
nor U14091 (N_14091,N_10636,N_10573);
nand U14092 (N_14092,N_11393,N_11730);
nand U14093 (N_14093,N_10404,N_10465);
and U14094 (N_14094,N_11510,N_10871);
or U14095 (N_14095,N_10850,N_10820);
and U14096 (N_14096,N_9700,N_10215);
and U14097 (N_14097,N_11877,N_10037);
nor U14098 (N_14098,N_11105,N_10352);
nor U14099 (N_14099,N_11151,N_10993);
nor U14100 (N_14100,N_11549,N_10175);
or U14101 (N_14101,N_11684,N_9723);
and U14102 (N_14102,N_10734,N_11135);
xnor U14103 (N_14103,N_9072,N_10469);
nand U14104 (N_14104,N_11522,N_11337);
nor U14105 (N_14105,N_9161,N_10797);
and U14106 (N_14106,N_11449,N_10349);
nor U14107 (N_14107,N_11548,N_9360);
and U14108 (N_14108,N_9825,N_10595);
nand U14109 (N_14109,N_9858,N_10516);
and U14110 (N_14110,N_9372,N_11710);
nor U14111 (N_14111,N_10764,N_9570);
nand U14112 (N_14112,N_9010,N_11896);
and U14113 (N_14113,N_10279,N_10827);
nor U14114 (N_14114,N_11442,N_9390);
or U14115 (N_14115,N_9838,N_9834);
nand U14116 (N_14116,N_10208,N_11121);
nor U14117 (N_14117,N_10350,N_9264);
and U14118 (N_14118,N_9228,N_10801);
nand U14119 (N_14119,N_10268,N_10384);
nor U14120 (N_14120,N_10209,N_9472);
nand U14121 (N_14121,N_10012,N_11158);
nor U14122 (N_14122,N_9583,N_10765);
nor U14123 (N_14123,N_10835,N_9441);
nand U14124 (N_14124,N_9368,N_9785);
nor U14125 (N_14125,N_9808,N_11302);
nand U14126 (N_14126,N_10295,N_9425);
and U14127 (N_14127,N_10660,N_11537);
and U14128 (N_14128,N_11037,N_9510);
or U14129 (N_14129,N_10159,N_10717);
or U14130 (N_14130,N_9712,N_9987);
nand U14131 (N_14131,N_11262,N_9853);
nand U14132 (N_14132,N_10226,N_10162);
nand U14133 (N_14133,N_11309,N_9677);
nand U14134 (N_14134,N_10051,N_10424);
and U14135 (N_14135,N_9159,N_10089);
or U14136 (N_14136,N_10160,N_10545);
or U14137 (N_14137,N_10637,N_9854);
or U14138 (N_14138,N_10545,N_10371);
and U14139 (N_14139,N_11108,N_9676);
nor U14140 (N_14140,N_9097,N_9924);
nand U14141 (N_14141,N_10751,N_11626);
and U14142 (N_14142,N_10375,N_10340);
xnor U14143 (N_14143,N_10250,N_10155);
and U14144 (N_14144,N_10002,N_9090);
nor U14145 (N_14145,N_9205,N_9196);
or U14146 (N_14146,N_10393,N_10289);
or U14147 (N_14147,N_9885,N_10399);
or U14148 (N_14148,N_10723,N_10784);
nor U14149 (N_14149,N_10237,N_11560);
and U14150 (N_14150,N_9080,N_11366);
nand U14151 (N_14151,N_9789,N_11882);
or U14152 (N_14152,N_10715,N_10480);
nor U14153 (N_14153,N_10841,N_9954);
nor U14154 (N_14154,N_10240,N_10194);
nand U14155 (N_14155,N_11248,N_9131);
or U14156 (N_14156,N_11062,N_10763);
or U14157 (N_14157,N_9380,N_9211);
nor U14158 (N_14158,N_11278,N_11830);
nor U14159 (N_14159,N_9467,N_9495);
and U14160 (N_14160,N_10744,N_9812);
nand U14161 (N_14161,N_10579,N_11080);
nand U14162 (N_14162,N_10415,N_9800);
nand U14163 (N_14163,N_11991,N_11904);
nor U14164 (N_14164,N_9965,N_10501);
nor U14165 (N_14165,N_9045,N_9169);
nand U14166 (N_14166,N_11968,N_9679);
nand U14167 (N_14167,N_11138,N_9896);
nor U14168 (N_14168,N_9206,N_9915);
nand U14169 (N_14169,N_11900,N_9535);
nor U14170 (N_14170,N_11552,N_9137);
or U14171 (N_14171,N_10102,N_10507);
and U14172 (N_14172,N_9066,N_9607);
or U14173 (N_14173,N_9173,N_11292);
nor U14174 (N_14174,N_10604,N_11048);
xnor U14175 (N_14175,N_10376,N_11200);
or U14176 (N_14176,N_11666,N_9406);
and U14177 (N_14177,N_9147,N_9854);
and U14178 (N_14178,N_11144,N_11250);
nand U14179 (N_14179,N_10727,N_9941);
nor U14180 (N_14180,N_11339,N_10443);
nand U14181 (N_14181,N_10637,N_10134);
and U14182 (N_14182,N_11749,N_11986);
and U14183 (N_14183,N_10680,N_10528);
nor U14184 (N_14184,N_10348,N_11265);
or U14185 (N_14185,N_11454,N_11489);
and U14186 (N_14186,N_10887,N_10876);
nand U14187 (N_14187,N_10795,N_11448);
and U14188 (N_14188,N_10355,N_11536);
or U14189 (N_14189,N_11921,N_11586);
or U14190 (N_14190,N_10247,N_10291);
and U14191 (N_14191,N_9694,N_9521);
nand U14192 (N_14192,N_11807,N_11382);
nand U14193 (N_14193,N_11699,N_11725);
nand U14194 (N_14194,N_10642,N_11576);
nor U14195 (N_14195,N_9552,N_9465);
nand U14196 (N_14196,N_11838,N_10112);
nand U14197 (N_14197,N_11938,N_10942);
or U14198 (N_14198,N_9181,N_10021);
nand U14199 (N_14199,N_9751,N_10871);
or U14200 (N_14200,N_9088,N_10727);
or U14201 (N_14201,N_11072,N_10092);
and U14202 (N_14202,N_9989,N_10834);
or U14203 (N_14203,N_9926,N_10233);
or U14204 (N_14204,N_11273,N_9029);
xor U14205 (N_14205,N_10505,N_10521);
or U14206 (N_14206,N_9452,N_11228);
and U14207 (N_14207,N_9220,N_11422);
and U14208 (N_14208,N_10252,N_9922);
and U14209 (N_14209,N_10050,N_9135);
or U14210 (N_14210,N_11746,N_9061);
and U14211 (N_14211,N_10422,N_10713);
nand U14212 (N_14212,N_9171,N_11378);
nor U14213 (N_14213,N_9004,N_11403);
nor U14214 (N_14214,N_11636,N_11882);
nand U14215 (N_14215,N_11358,N_11654);
and U14216 (N_14216,N_9292,N_9289);
nor U14217 (N_14217,N_9477,N_9175);
and U14218 (N_14218,N_10426,N_9599);
and U14219 (N_14219,N_10242,N_11197);
and U14220 (N_14220,N_11159,N_10431);
or U14221 (N_14221,N_11134,N_10348);
nand U14222 (N_14222,N_9284,N_11701);
nand U14223 (N_14223,N_9060,N_9136);
or U14224 (N_14224,N_10034,N_10166);
nor U14225 (N_14225,N_10578,N_9246);
nor U14226 (N_14226,N_11759,N_11591);
or U14227 (N_14227,N_11282,N_11157);
and U14228 (N_14228,N_11285,N_10282);
nor U14229 (N_14229,N_10799,N_11907);
nand U14230 (N_14230,N_9067,N_9457);
nand U14231 (N_14231,N_10760,N_10981);
xor U14232 (N_14232,N_11972,N_11751);
and U14233 (N_14233,N_11112,N_11697);
nor U14234 (N_14234,N_11979,N_11594);
nand U14235 (N_14235,N_9588,N_9719);
nor U14236 (N_14236,N_10503,N_10037);
and U14237 (N_14237,N_10073,N_10759);
nor U14238 (N_14238,N_10971,N_9943);
and U14239 (N_14239,N_9006,N_11435);
nand U14240 (N_14240,N_9499,N_11163);
and U14241 (N_14241,N_10750,N_9716);
and U14242 (N_14242,N_11394,N_9961);
nand U14243 (N_14243,N_10189,N_11768);
or U14244 (N_14244,N_11431,N_9797);
and U14245 (N_14245,N_11215,N_11726);
nor U14246 (N_14246,N_9683,N_11458);
nand U14247 (N_14247,N_11910,N_9247);
nand U14248 (N_14248,N_10941,N_10404);
or U14249 (N_14249,N_9185,N_11490);
nor U14250 (N_14250,N_11872,N_10964);
nand U14251 (N_14251,N_11857,N_11878);
nor U14252 (N_14252,N_9122,N_9695);
and U14253 (N_14253,N_10229,N_10702);
and U14254 (N_14254,N_10992,N_9701);
nand U14255 (N_14255,N_10522,N_10361);
and U14256 (N_14256,N_9371,N_9960);
nand U14257 (N_14257,N_11332,N_9048);
nand U14258 (N_14258,N_9963,N_11417);
nand U14259 (N_14259,N_11521,N_10850);
nor U14260 (N_14260,N_11686,N_11015);
and U14261 (N_14261,N_10863,N_10191);
nor U14262 (N_14262,N_9706,N_11498);
nor U14263 (N_14263,N_11845,N_10452);
nor U14264 (N_14264,N_9823,N_10397);
nand U14265 (N_14265,N_10121,N_11600);
nor U14266 (N_14266,N_11339,N_10007);
nand U14267 (N_14267,N_11626,N_9826);
or U14268 (N_14268,N_10711,N_10548);
nand U14269 (N_14269,N_11982,N_10968);
nor U14270 (N_14270,N_10303,N_9703);
nor U14271 (N_14271,N_9858,N_11694);
and U14272 (N_14272,N_10402,N_9767);
or U14273 (N_14273,N_10303,N_9128);
nand U14274 (N_14274,N_9620,N_10108);
or U14275 (N_14275,N_9185,N_11736);
or U14276 (N_14276,N_10716,N_10694);
nand U14277 (N_14277,N_11869,N_10737);
nand U14278 (N_14278,N_9506,N_10183);
or U14279 (N_14279,N_11717,N_10211);
and U14280 (N_14280,N_11707,N_10435);
and U14281 (N_14281,N_9701,N_10861);
and U14282 (N_14282,N_10136,N_11551);
xnor U14283 (N_14283,N_9106,N_9416);
nand U14284 (N_14284,N_10657,N_11577);
nand U14285 (N_14285,N_11028,N_9893);
and U14286 (N_14286,N_10718,N_9727);
and U14287 (N_14287,N_9703,N_9637);
nor U14288 (N_14288,N_9177,N_11252);
nand U14289 (N_14289,N_11251,N_11133);
or U14290 (N_14290,N_11302,N_11187);
nor U14291 (N_14291,N_9221,N_9915);
nand U14292 (N_14292,N_9553,N_9297);
or U14293 (N_14293,N_9121,N_9075);
and U14294 (N_14294,N_9584,N_10255);
nand U14295 (N_14295,N_9839,N_10820);
nand U14296 (N_14296,N_9173,N_10844);
nor U14297 (N_14297,N_9028,N_10211);
and U14298 (N_14298,N_10467,N_9967);
nor U14299 (N_14299,N_9219,N_9726);
and U14300 (N_14300,N_9704,N_10202);
or U14301 (N_14301,N_11368,N_11664);
nand U14302 (N_14302,N_9432,N_11113);
and U14303 (N_14303,N_9581,N_9622);
and U14304 (N_14304,N_11638,N_10308);
nand U14305 (N_14305,N_9082,N_10036);
and U14306 (N_14306,N_10685,N_10465);
or U14307 (N_14307,N_11295,N_10161);
nor U14308 (N_14308,N_10531,N_11315);
nor U14309 (N_14309,N_9637,N_9520);
and U14310 (N_14310,N_9857,N_9560);
nand U14311 (N_14311,N_11101,N_11467);
and U14312 (N_14312,N_10080,N_10453);
and U14313 (N_14313,N_11984,N_10153);
or U14314 (N_14314,N_10025,N_10940);
or U14315 (N_14315,N_10025,N_10342);
nor U14316 (N_14316,N_9172,N_9079);
nor U14317 (N_14317,N_9373,N_9396);
or U14318 (N_14318,N_10736,N_9003);
or U14319 (N_14319,N_11306,N_11238);
nand U14320 (N_14320,N_11568,N_9147);
nor U14321 (N_14321,N_9426,N_10119);
nand U14322 (N_14322,N_11645,N_11749);
nor U14323 (N_14323,N_10168,N_11708);
nor U14324 (N_14324,N_9169,N_11540);
and U14325 (N_14325,N_10964,N_9755);
and U14326 (N_14326,N_11906,N_11815);
and U14327 (N_14327,N_10387,N_9154);
or U14328 (N_14328,N_10937,N_9724);
or U14329 (N_14329,N_10735,N_11747);
or U14330 (N_14330,N_9320,N_10001);
nand U14331 (N_14331,N_9804,N_9245);
and U14332 (N_14332,N_11067,N_9473);
nand U14333 (N_14333,N_11868,N_11756);
or U14334 (N_14334,N_11139,N_11527);
and U14335 (N_14335,N_11875,N_11369);
nor U14336 (N_14336,N_9827,N_11483);
nor U14337 (N_14337,N_11871,N_9358);
nor U14338 (N_14338,N_11523,N_9331);
or U14339 (N_14339,N_10681,N_10021);
nor U14340 (N_14340,N_11789,N_9305);
nand U14341 (N_14341,N_11259,N_11753);
nand U14342 (N_14342,N_11246,N_11107);
nand U14343 (N_14343,N_9127,N_10990);
or U14344 (N_14344,N_10101,N_11026);
nor U14345 (N_14345,N_10023,N_10421);
nand U14346 (N_14346,N_10419,N_9647);
nand U14347 (N_14347,N_11798,N_10002);
nor U14348 (N_14348,N_9071,N_9056);
and U14349 (N_14349,N_11484,N_10273);
nor U14350 (N_14350,N_11543,N_9386);
nor U14351 (N_14351,N_9067,N_10201);
nor U14352 (N_14352,N_10456,N_10337);
or U14353 (N_14353,N_11913,N_11277);
or U14354 (N_14354,N_10931,N_11844);
and U14355 (N_14355,N_9982,N_9078);
nand U14356 (N_14356,N_9261,N_11177);
nand U14357 (N_14357,N_11824,N_9370);
or U14358 (N_14358,N_10116,N_9228);
nor U14359 (N_14359,N_10251,N_11777);
and U14360 (N_14360,N_11220,N_10222);
xnor U14361 (N_14361,N_11429,N_9337);
nor U14362 (N_14362,N_10596,N_11567);
or U14363 (N_14363,N_10254,N_11094);
nor U14364 (N_14364,N_11963,N_11207);
nor U14365 (N_14365,N_11042,N_10526);
nor U14366 (N_14366,N_9968,N_9921);
and U14367 (N_14367,N_11615,N_11782);
nand U14368 (N_14368,N_9736,N_9553);
nand U14369 (N_14369,N_10004,N_11311);
nand U14370 (N_14370,N_9205,N_10637);
or U14371 (N_14371,N_10364,N_11269);
and U14372 (N_14372,N_9760,N_9481);
nand U14373 (N_14373,N_9820,N_10920);
nor U14374 (N_14374,N_9538,N_11052);
and U14375 (N_14375,N_11703,N_11463);
and U14376 (N_14376,N_10455,N_10772);
nor U14377 (N_14377,N_10912,N_10132);
or U14378 (N_14378,N_11888,N_10349);
or U14379 (N_14379,N_10152,N_11314);
nand U14380 (N_14380,N_11507,N_11239);
nand U14381 (N_14381,N_9447,N_11486);
nand U14382 (N_14382,N_9673,N_11870);
nor U14383 (N_14383,N_9023,N_11914);
nand U14384 (N_14384,N_9932,N_10138);
nor U14385 (N_14385,N_9349,N_9158);
and U14386 (N_14386,N_9301,N_9435);
and U14387 (N_14387,N_11033,N_11429);
nor U14388 (N_14388,N_9074,N_10845);
nor U14389 (N_14389,N_11439,N_9728);
or U14390 (N_14390,N_9846,N_9038);
and U14391 (N_14391,N_9685,N_11195);
or U14392 (N_14392,N_11208,N_11039);
nor U14393 (N_14393,N_11349,N_11114);
nand U14394 (N_14394,N_9398,N_10227);
nor U14395 (N_14395,N_10194,N_9530);
and U14396 (N_14396,N_11497,N_9062);
nor U14397 (N_14397,N_10649,N_11351);
and U14398 (N_14398,N_11632,N_9075);
nor U14399 (N_14399,N_10673,N_9386);
nor U14400 (N_14400,N_11718,N_9020);
nor U14401 (N_14401,N_9059,N_10201);
nor U14402 (N_14402,N_9398,N_11747);
nand U14403 (N_14403,N_11272,N_9115);
and U14404 (N_14404,N_11360,N_9913);
nor U14405 (N_14405,N_10226,N_9222);
nand U14406 (N_14406,N_11927,N_10574);
and U14407 (N_14407,N_11225,N_9092);
nand U14408 (N_14408,N_9304,N_10388);
nand U14409 (N_14409,N_11094,N_9680);
nor U14410 (N_14410,N_9000,N_9599);
and U14411 (N_14411,N_11617,N_10782);
or U14412 (N_14412,N_9411,N_10808);
or U14413 (N_14413,N_11767,N_11394);
nor U14414 (N_14414,N_9060,N_10917);
nor U14415 (N_14415,N_10259,N_11999);
or U14416 (N_14416,N_11196,N_10689);
nand U14417 (N_14417,N_10030,N_10534);
nor U14418 (N_14418,N_9012,N_9403);
and U14419 (N_14419,N_10429,N_11465);
nand U14420 (N_14420,N_9995,N_9434);
and U14421 (N_14421,N_10381,N_10030);
nand U14422 (N_14422,N_9430,N_11312);
nor U14423 (N_14423,N_10942,N_10727);
and U14424 (N_14424,N_11997,N_9996);
or U14425 (N_14425,N_10647,N_11837);
nor U14426 (N_14426,N_9096,N_11179);
nand U14427 (N_14427,N_10585,N_9402);
xnor U14428 (N_14428,N_9728,N_11452);
or U14429 (N_14429,N_9374,N_10954);
nor U14430 (N_14430,N_11988,N_10383);
or U14431 (N_14431,N_11429,N_9544);
and U14432 (N_14432,N_10595,N_10839);
or U14433 (N_14433,N_11896,N_10999);
nand U14434 (N_14434,N_9418,N_9009);
nand U14435 (N_14435,N_9674,N_10753);
or U14436 (N_14436,N_10110,N_9407);
nor U14437 (N_14437,N_11134,N_10327);
or U14438 (N_14438,N_10117,N_9649);
nor U14439 (N_14439,N_11983,N_10070);
nor U14440 (N_14440,N_9131,N_9108);
or U14441 (N_14441,N_9707,N_11785);
nand U14442 (N_14442,N_10960,N_9713);
or U14443 (N_14443,N_11385,N_10945);
or U14444 (N_14444,N_9493,N_10982);
nor U14445 (N_14445,N_9716,N_11220);
or U14446 (N_14446,N_11943,N_11836);
nand U14447 (N_14447,N_11700,N_11060);
nor U14448 (N_14448,N_9651,N_9833);
nor U14449 (N_14449,N_11528,N_9227);
or U14450 (N_14450,N_11108,N_10323);
nor U14451 (N_14451,N_10960,N_10967);
or U14452 (N_14452,N_11452,N_11457);
nor U14453 (N_14453,N_10450,N_10698);
or U14454 (N_14454,N_10920,N_10465);
or U14455 (N_14455,N_11144,N_10123);
nand U14456 (N_14456,N_9602,N_10919);
and U14457 (N_14457,N_9259,N_9364);
nand U14458 (N_14458,N_11890,N_10637);
nor U14459 (N_14459,N_11460,N_9132);
nor U14460 (N_14460,N_9166,N_9011);
and U14461 (N_14461,N_10306,N_10459);
or U14462 (N_14462,N_11193,N_10934);
and U14463 (N_14463,N_10991,N_11306);
or U14464 (N_14464,N_11831,N_11284);
and U14465 (N_14465,N_11507,N_10037);
and U14466 (N_14466,N_9360,N_9763);
or U14467 (N_14467,N_10279,N_11752);
or U14468 (N_14468,N_9671,N_9076);
nand U14469 (N_14469,N_10622,N_11999);
or U14470 (N_14470,N_11516,N_9001);
and U14471 (N_14471,N_11047,N_11906);
nand U14472 (N_14472,N_9268,N_10339);
and U14473 (N_14473,N_10817,N_11331);
nand U14474 (N_14474,N_10798,N_11588);
nor U14475 (N_14475,N_11210,N_9820);
nor U14476 (N_14476,N_10878,N_9585);
or U14477 (N_14477,N_10218,N_11056);
xor U14478 (N_14478,N_9140,N_10341);
nor U14479 (N_14479,N_11733,N_10789);
and U14480 (N_14480,N_10531,N_10306);
and U14481 (N_14481,N_11839,N_9717);
or U14482 (N_14482,N_11307,N_10937);
or U14483 (N_14483,N_11424,N_11378);
or U14484 (N_14484,N_9742,N_10652);
or U14485 (N_14485,N_11203,N_10032);
nor U14486 (N_14486,N_10566,N_9966);
or U14487 (N_14487,N_10967,N_9615);
nor U14488 (N_14488,N_11010,N_9712);
nand U14489 (N_14489,N_10883,N_10705);
nor U14490 (N_14490,N_9508,N_10167);
or U14491 (N_14491,N_11971,N_11306);
nand U14492 (N_14492,N_11473,N_11381);
xor U14493 (N_14493,N_11413,N_11334);
or U14494 (N_14494,N_9885,N_9188);
nor U14495 (N_14495,N_10664,N_9448);
and U14496 (N_14496,N_10773,N_9175);
and U14497 (N_14497,N_11663,N_9019);
nand U14498 (N_14498,N_11627,N_9186);
and U14499 (N_14499,N_9473,N_10875);
or U14500 (N_14500,N_11057,N_9126);
nand U14501 (N_14501,N_11088,N_11586);
nand U14502 (N_14502,N_10777,N_10062);
nand U14503 (N_14503,N_10510,N_10779);
or U14504 (N_14504,N_10715,N_11324);
or U14505 (N_14505,N_11992,N_11205);
and U14506 (N_14506,N_11497,N_10340);
and U14507 (N_14507,N_11007,N_9524);
nand U14508 (N_14508,N_9848,N_10564);
nor U14509 (N_14509,N_10832,N_10827);
and U14510 (N_14510,N_9304,N_10163);
and U14511 (N_14511,N_9677,N_10364);
nand U14512 (N_14512,N_10726,N_11312);
nand U14513 (N_14513,N_10331,N_9297);
and U14514 (N_14514,N_9607,N_10078);
and U14515 (N_14515,N_10493,N_9100);
and U14516 (N_14516,N_11863,N_11693);
or U14517 (N_14517,N_10843,N_11265);
and U14518 (N_14518,N_11236,N_11133);
nand U14519 (N_14519,N_10299,N_11266);
nor U14520 (N_14520,N_10970,N_11657);
nor U14521 (N_14521,N_9169,N_10039);
nand U14522 (N_14522,N_9200,N_9011);
and U14523 (N_14523,N_10614,N_11631);
nand U14524 (N_14524,N_10111,N_11755);
nor U14525 (N_14525,N_10917,N_9398);
nor U14526 (N_14526,N_9288,N_11994);
nand U14527 (N_14527,N_9914,N_10395);
nor U14528 (N_14528,N_10774,N_9836);
nand U14529 (N_14529,N_11389,N_10400);
nor U14530 (N_14530,N_9368,N_9485);
and U14531 (N_14531,N_9622,N_9927);
and U14532 (N_14532,N_11566,N_11517);
nand U14533 (N_14533,N_11873,N_10709);
nand U14534 (N_14534,N_10291,N_11074);
and U14535 (N_14535,N_10213,N_10060);
nor U14536 (N_14536,N_10180,N_9236);
and U14537 (N_14537,N_9349,N_10719);
nor U14538 (N_14538,N_9524,N_11365);
or U14539 (N_14539,N_9628,N_9753);
or U14540 (N_14540,N_11941,N_11974);
and U14541 (N_14541,N_11172,N_9148);
nor U14542 (N_14542,N_11762,N_10708);
or U14543 (N_14543,N_10410,N_10943);
nand U14544 (N_14544,N_11113,N_11315);
and U14545 (N_14545,N_11628,N_10526);
or U14546 (N_14546,N_11583,N_9851);
nor U14547 (N_14547,N_11634,N_9003);
nand U14548 (N_14548,N_9199,N_9860);
or U14549 (N_14549,N_9297,N_9848);
and U14550 (N_14550,N_11160,N_10518);
nor U14551 (N_14551,N_10793,N_9661);
nand U14552 (N_14552,N_11403,N_9770);
and U14553 (N_14553,N_9737,N_10479);
nor U14554 (N_14554,N_9622,N_10054);
nor U14555 (N_14555,N_11404,N_10974);
nor U14556 (N_14556,N_11401,N_11299);
or U14557 (N_14557,N_9085,N_11557);
nor U14558 (N_14558,N_10166,N_11608);
nand U14559 (N_14559,N_10262,N_11255);
nand U14560 (N_14560,N_11390,N_10295);
and U14561 (N_14561,N_11413,N_11050);
nand U14562 (N_14562,N_10725,N_10674);
nor U14563 (N_14563,N_10832,N_10409);
or U14564 (N_14564,N_11666,N_9102);
nor U14565 (N_14565,N_11885,N_11085);
or U14566 (N_14566,N_11974,N_10602);
nand U14567 (N_14567,N_11488,N_10880);
or U14568 (N_14568,N_11296,N_11805);
or U14569 (N_14569,N_10489,N_9664);
or U14570 (N_14570,N_11079,N_10794);
nor U14571 (N_14571,N_10565,N_9144);
nand U14572 (N_14572,N_9364,N_10784);
or U14573 (N_14573,N_10653,N_9159);
xor U14574 (N_14574,N_10425,N_11624);
and U14575 (N_14575,N_10814,N_11030);
nor U14576 (N_14576,N_9584,N_9070);
and U14577 (N_14577,N_10371,N_9929);
nor U14578 (N_14578,N_10424,N_10308);
and U14579 (N_14579,N_10969,N_9974);
nand U14580 (N_14580,N_11307,N_10993);
xor U14581 (N_14581,N_11146,N_9889);
nor U14582 (N_14582,N_11834,N_10559);
nor U14583 (N_14583,N_10464,N_10657);
nand U14584 (N_14584,N_11382,N_11303);
nor U14585 (N_14585,N_10662,N_11625);
or U14586 (N_14586,N_11095,N_10406);
nand U14587 (N_14587,N_11359,N_11867);
or U14588 (N_14588,N_10739,N_9611);
nand U14589 (N_14589,N_11354,N_10090);
or U14590 (N_14590,N_11296,N_9919);
or U14591 (N_14591,N_11310,N_10278);
nor U14592 (N_14592,N_9561,N_10884);
nor U14593 (N_14593,N_11440,N_9440);
nand U14594 (N_14594,N_11312,N_11161);
nor U14595 (N_14595,N_11057,N_11732);
and U14596 (N_14596,N_11934,N_10450);
nand U14597 (N_14597,N_11774,N_9063);
nand U14598 (N_14598,N_10660,N_11709);
nor U14599 (N_14599,N_9905,N_11960);
nand U14600 (N_14600,N_10030,N_11861);
or U14601 (N_14601,N_9241,N_11410);
nor U14602 (N_14602,N_9316,N_9813);
nor U14603 (N_14603,N_11493,N_11033);
nor U14604 (N_14604,N_9360,N_9690);
nand U14605 (N_14605,N_9288,N_9997);
or U14606 (N_14606,N_9013,N_9897);
or U14607 (N_14607,N_11233,N_10843);
nor U14608 (N_14608,N_9512,N_10109);
or U14609 (N_14609,N_11658,N_9243);
or U14610 (N_14610,N_11503,N_9808);
nand U14611 (N_14611,N_9018,N_11644);
nor U14612 (N_14612,N_9414,N_10590);
nor U14613 (N_14613,N_11287,N_10039);
nand U14614 (N_14614,N_10696,N_10456);
or U14615 (N_14615,N_10796,N_11770);
and U14616 (N_14616,N_11089,N_11116);
nor U14617 (N_14617,N_10947,N_10244);
nor U14618 (N_14618,N_9811,N_11820);
nand U14619 (N_14619,N_9660,N_11004);
xnor U14620 (N_14620,N_9979,N_10714);
nand U14621 (N_14621,N_9029,N_10121);
and U14622 (N_14622,N_10662,N_10933);
nor U14623 (N_14623,N_11673,N_10783);
and U14624 (N_14624,N_10623,N_9532);
nor U14625 (N_14625,N_10837,N_9988);
and U14626 (N_14626,N_10599,N_11718);
nor U14627 (N_14627,N_9189,N_9789);
nand U14628 (N_14628,N_10867,N_10256);
nor U14629 (N_14629,N_10273,N_11678);
and U14630 (N_14630,N_9222,N_9975);
nor U14631 (N_14631,N_9978,N_10099);
nor U14632 (N_14632,N_11349,N_10613);
nand U14633 (N_14633,N_9419,N_9159);
and U14634 (N_14634,N_10047,N_9371);
nand U14635 (N_14635,N_11013,N_10000);
or U14636 (N_14636,N_9360,N_9140);
nor U14637 (N_14637,N_10721,N_10427);
and U14638 (N_14638,N_11471,N_9769);
nor U14639 (N_14639,N_11527,N_11083);
and U14640 (N_14640,N_10723,N_11255);
nand U14641 (N_14641,N_10352,N_11667);
or U14642 (N_14642,N_9009,N_9707);
or U14643 (N_14643,N_10948,N_9611);
or U14644 (N_14644,N_11136,N_11425);
nand U14645 (N_14645,N_10393,N_11314);
and U14646 (N_14646,N_9874,N_10304);
nor U14647 (N_14647,N_10221,N_9250);
nand U14648 (N_14648,N_9829,N_9261);
and U14649 (N_14649,N_10853,N_9622);
nand U14650 (N_14650,N_11609,N_9076);
and U14651 (N_14651,N_11472,N_11648);
nor U14652 (N_14652,N_11742,N_11685);
nand U14653 (N_14653,N_9118,N_11437);
and U14654 (N_14654,N_9092,N_11548);
nand U14655 (N_14655,N_11905,N_9208);
nand U14656 (N_14656,N_10244,N_11541);
nor U14657 (N_14657,N_11929,N_10415);
nand U14658 (N_14658,N_9697,N_9324);
nand U14659 (N_14659,N_10028,N_10132);
and U14660 (N_14660,N_9603,N_11888);
xnor U14661 (N_14661,N_11814,N_10175);
nor U14662 (N_14662,N_9623,N_9141);
nand U14663 (N_14663,N_11286,N_10515);
nor U14664 (N_14664,N_11887,N_11804);
nor U14665 (N_14665,N_10358,N_11221);
and U14666 (N_14666,N_11041,N_11429);
and U14667 (N_14667,N_10984,N_10870);
and U14668 (N_14668,N_11594,N_9115);
nor U14669 (N_14669,N_9415,N_9093);
nand U14670 (N_14670,N_11273,N_9254);
and U14671 (N_14671,N_10846,N_9506);
and U14672 (N_14672,N_9530,N_11243);
and U14673 (N_14673,N_11736,N_11853);
nor U14674 (N_14674,N_10659,N_9087);
and U14675 (N_14675,N_9510,N_9375);
and U14676 (N_14676,N_11990,N_11533);
and U14677 (N_14677,N_11402,N_11924);
and U14678 (N_14678,N_9111,N_9059);
or U14679 (N_14679,N_10944,N_10303);
nand U14680 (N_14680,N_10049,N_11274);
and U14681 (N_14681,N_11046,N_10450);
or U14682 (N_14682,N_10272,N_11725);
or U14683 (N_14683,N_9059,N_11837);
nor U14684 (N_14684,N_10980,N_10184);
nor U14685 (N_14685,N_10081,N_11980);
or U14686 (N_14686,N_10585,N_11123);
or U14687 (N_14687,N_11932,N_11717);
or U14688 (N_14688,N_11032,N_11094);
or U14689 (N_14689,N_9330,N_9842);
nor U14690 (N_14690,N_10227,N_11970);
nor U14691 (N_14691,N_11930,N_9687);
xor U14692 (N_14692,N_9592,N_11801);
nand U14693 (N_14693,N_9643,N_9541);
nor U14694 (N_14694,N_9044,N_10728);
and U14695 (N_14695,N_9643,N_10500);
nor U14696 (N_14696,N_10269,N_9892);
xor U14697 (N_14697,N_10156,N_9615);
nand U14698 (N_14698,N_9866,N_9840);
and U14699 (N_14699,N_9138,N_9321);
and U14700 (N_14700,N_11517,N_9878);
or U14701 (N_14701,N_11615,N_10592);
and U14702 (N_14702,N_10934,N_11352);
nor U14703 (N_14703,N_9110,N_9309);
and U14704 (N_14704,N_10100,N_11125);
or U14705 (N_14705,N_11718,N_9286);
and U14706 (N_14706,N_10066,N_10844);
xor U14707 (N_14707,N_10551,N_11433);
and U14708 (N_14708,N_9886,N_10855);
or U14709 (N_14709,N_10676,N_10670);
and U14710 (N_14710,N_9009,N_9563);
and U14711 (N_14711,N_9973,N_9759);
and U14712 (N_14712,N_10135,N_10767);
or U14713 (N_14713,N_11642,N_9957);
and U14714 (N_14714,N_11833,N_10550);
nor U14715 (N_14715,N_9730,N_9795);
and U14716 (N_14716,N_10869,N_10865);
nand U14717 (N_14717,N_10800,N_9364);
nand U14718 (N_14718,N_9496,N_10126);
or U14719 (N_14719,N_11311,N_9388);
nand U14720 (N_14720,N_10147,N_10988);
and U14721 (N_14721,N_10761,N_9250);
nor U14722 (N_14722,N_10274,N_9514);
or U14723 (N_14723,N_10734,N_11877);
nor U14724 (N_14724,N_10900,N_11365);
nor U14725 (N_14725,N_11906,N_9877);
or U14726 (N_14726,N_9126,N_11467);
or U14727 (N_14727,N_9763,N_11921);
nor U14728 (N_14728,N_11621,N_10026);
nand U14729 (N_14729,N_11846,N_11553);
or U14730 (N_14730,N_9874,N_9327);
and U14731 (N_14731,N_9604,N_9934);
and U14732 (N_14732,N_9458,N_9962);
and U14733 (N_14733,N_9143,N_9148);
or U14734 (N_14734,N_11983,N_9724);
xnor U14735 (N_14735,N_10911,N_11777);
nand U14736 (N_14736,N_9747,N_11327);
nand U14737 (N_14737,N_11981,N_10095);
nand U14738 (N_14738,N_9302,N_10271);
and U14739 (N_14739,N_9750,N_9297);
nor U14740 (N_14740,N_9660,N_10516);
and U14741 (N_14741,N_9726,N_9162);
or U14742 (N_14742,N_11714,N_9062);
or U14743 (N_14743,N_11092,N_11724);
nor U14744 (N_14744,N_9480,N_9271);
nor U14745 (N_14745,N_9428,N_11037);
or U14746 (N_14746,N_11559,N_11102);
nand U14747 (N_14747,N_10033,N_11116);
nor U14748 (N_14748,N_9465,N_11493);
nand U14749 (N_14749,N_10883,N_9546);
nand U14750 (N_14750,N_9235,N_10768);
nand U14751 (N_14751,N_10336,N_10233);
or U14752 (N_14752,N_9933,N_10751);
or U14753 (N_14753,N_11609,N_11157);
nand U14754 (N_14754,N_9419,N_11381);
and U14755 (N_14755,N_10194,N_10308);
nand U14756 (N_14756,N_10088,N_9684);
nand U14757 (N_14757,N_11208,N_9654);
nor U14758 (N_14758,N_11183,N_11780);
and U14759 (N_14759,N_9252,N_11178);
nand U14760 (N_14760,N_10155,N_11020);
or U14761 (N_14761,N_10412,N_9714);
nand U14762 (N_14762,N_10565,N_11778);
nor U14763 (N_14763,N_11279,N_10448);
nand U14764 (N_14764,N_11942,N_10283);
and U14765 (N_14765,N_9855,N_10224);
nor U14766 (N_14766,N_10649,N_10085);
nand U14767 (N_14767,N_11740,N_9256);
nor U14768 (N_14768,N_11343,N_10374);
or U14769 (N_14769,N_11706,N_11562);
and U14770 (N_14770,N_9112,N_10319);
nor U14771 (N_14771,N_10912,N_9081);
and U14772 (N_14772,N_10299,N_9803);
or U14773 (N_14773,N_9928,N_10464);
and U14774 (N_14774,N_10113,N_11409);
or U14775 (N_14775,N_11649,N_10264);
nand U14776 (N_14776,N_11205,N_11174);
and U14777 (N_14777,N_10088,N_11732);
nor U14778 (N_14778,N_11481,N_10341);
or U14779 (N_14779,N_11443,N_10016);
or U14780 (N_14780,N_10797,N_11274);
or U14781 (N_14781,N_11964,N_9786);
nand U14782 (N_14782,N_11030,N_10094);
nand U14783 (N_14783,N_11410,N_10496);
or U14784 (N_14784,N_9287,N_11718);
and U14785 (N_14785,N_10990,N_10124);
and U14786 (N_14786,N_10528,N_10482);
nand U14787 (N_14787,N_10962,N_10561);
nor U14788 (N_14788,N_9426,N_10338);
nor U14789 (N_14789,N_9899,N_10348);
and U14790 (N_14790,N_10863,N_10982);
nor U14791 (N_14791,N_11510,N_10463);
or U14792 (N_14792,N_9605,N_9302);
or U14793 (N_14793,N_10261,N_10768);
or U14794 (N_14794,N_10508,N_10646);
nand U14795 (N_14795,N_11404,N_9365);
and U14796 (N_14796,N_11798,N_9065);
nor U14797 (N_14797,N_10018,N_10505);
or U14798 (N_14798,N_10862,N_11376);
or U14799 (N_14799,N_10054,N_10262);
nor U14800 (N_14800,N_11661,N_11780);
or U14801 (N_14801,N_9047,N_10882);
or U14802 (N_14802,N_10963,N_10703);
or U14803 (N_14803,N_10445,N_10711);
nand U14804 (N_14804,N_11199,N_9757);
nand U14805 (N_14805,N_10023,N_11175);
and U14806 (N_14806,N_11320,N_10483);
or U14807 (N_14807,N_10367,N_11799);
nand U14808 (N_14808,N_9213,N_10517);
nand U14809 (N_14809,N_10339,N_9263);
nor U14810 (N_14810,N_10732,N_10240);
or U14811 (N_14811,N_9024,N_11204);
or U14812 (N_14812,N_10781,N_9145);
nand U14813 (N_14813,N_11818,N_9335);
nand U14814 (N_14814,N_9338,N_11230);
and U14815 (N_14815,N_9540,N_11235);
nor U14816 (N_14816,N_10103,N_10368);
nand U14817 (N_14817,N_11966,N_10088);
and U14818 (N_14818,N_9497,N_9301);
nor U14819 (N_14819,N_11612,N_10132);
nor U14820 (N_14820,N_10450,N_9243);
and U14821 (N_14821,N_11965,N_11085);
nor U14822 (N_14822,N_9837,N_10813);
nor U14823 (N_14823,N_9877,N_11470);
nor U14824 (N_14824,N_10192,N_9745);
and U14825 (N_14825,N_9014,N_9508);
and U14826 (N_14826,N_9386,N_10326);
xor U14827 (N_14827,N_9073,N_10227);
nand U14828 (N_14828,N_11600,N_10658);
or U14829 (N_14829,N_9013,N_9545);
nand U14830 (N_14830,N_11107,N_9849);
nand U14831 (N_14831,N_11648,N_10828);
or U14832 (N_14832,N_9236,N_10328);
and U14833 (N_14833,N_9016,N_9766);
and U14834 (N_14834,N_11086,N_10736);
nor U14835 (N_14835,N_11063,N_11413);
nor U14836 (N_14836,N_9779,N_9124);
nor U14837 (N_14837,N_11469,N_9180);
nor U14838 (N_14838,N_11740,N_9480);
nand U14839 (N_14839,N_11441,N_10297);
and U14840 (N_14840,N_11381,N_10252);
nand U14841 (N_14841,N_10337,N_10758);
and U14842 (N_14842,N_11491,N_10533);
and U14843 (N_14843,N_11546,N_9176);
and U14844 (N_14844,N_10999,N_9764);
and U14845 (N_14845,N_10169,N_9346);
or U14846 (N_14846,N_9110,N_10093);
and U14847 (N_14847,N_9965,N_11248);
nand U14848 (N_14848,N_9592,N_9642);
and U14849 (N_14849,N_9746,N_9495);
nor U14850 (N_14850,N_10504,N_9945);
and U14851 (N_14851,N_9059,N_10975);
or U14852 (N_14852,N_10742,N_9490);
and U14853 (N_14853,N_10195,N_9018);
nor U14854 (N_14854,N_11625,N_9823);
nor U14855 (N_14855,N_9962,N_10784);
nor U14856 (N_14856,N_9713,N_11489);
nand U14857 (N_14857,N_9101,N_9556);
or U14858 (N_14858,N_10864,N_9103);
nand U14859 (N_14859,N_9493,N_9439);
nand U14860 (N_14860,N_9770,N_10716);
or U14861 (N_14861,N_11028,N_9458);
nand U14862 (N_14862,N_11434,N_10696);
or U14863 (N_14863,N_10488,N_9581);
nand U14864 (N_14864,N_9854,N_11347);
and U14865 (N_14865,N_9202,N_9267);
nor U14866 (N_14866,N_11120,N_10235);
nand U14867 (N_14867,N_9755,N_9778);
or U14868 (N_14868,N_11956,N_11584);
and U14869 (N_14869,N_11544,N_9045);
nor U14870 (N_14870,N_11258,N_9205);
or U14871 (N_14871,N_10992,N_9068);
xor U14872 (N_14872,N_11276,N_10980);
and U14873 (N_14873,N_9067,N_11391);
nand U14874 (N_14874,N_11455,N_9144);
or U14875 (N_14875,N_9583,N_9483);
and U14876 (N_14876,N_11260,N_10893);
nor U14877 (N_14877,N_11263,N_9974);
nor U14878 (N_14878,N_9614,N_9067);
xnor U14879 (N_14879,N_10294,N_9631);
nor U14880 (N_14880,N_9032,N_9361);
and U14881 (N_14881,N_11859,N_10494);
nand U14882 (N_14882,N_9954,N_10851);
or U14883 (N_14883,N_9014,N_10351);
and U14884 (N_14884,N_10126,N_10604);
nand U14885 (N_14885,N_10812,N_10158);
and U14886 (N_14886,N_11719,N_10516);
or U14887 (N_14887,N_11318,N_9787);
nor U14888 (N_14888,N_10247,N_9469);
nand U14889 (N_14889,N_10007,N_9329);
or U14890 (N_14890,N_11338,N_9523);
or U14891 (N_14891,N_10470,N_10837);
nand U14892 (N_14892,N_9629,N_9579);
and U14893 (N_14893,N_9325,N_10248);
or U14894 (N_14894,N_11356,N_9066);
and U14895 (N_14895,N_10525,N_10200);
and U14896 (N_14896,N_10281,N_10601);
and U14897 (N_14897,N_10818,N_9716);
nand U14898 (N_14898,N_9664,N_10910);
or U14899 (N_14899,N_9398,N_10451);
xor U14900 (N_14900,N_11939,N_11428);
and U14901 (N_14901,N_10612,N_9121);
and U14902 (N_14902,N_10194,N_11485);
and U14903 (N_14903,N_11060,N_9621);
nand U14904 (N_14904,N_11528,N_10168);
and U14905 (N_14905,N_9250,N_9881);
or U14906 (N_14906,N_11100,N_10709);
nand U14907 (N_14907,N_10016,N_10545);
or U14908 (N_14908,N_10847,N_10895);
nand U14909 (N_14909,N_10919,N_10499);
or U14910 (N_14910,N_9907,N_11282);
and U14911 (N_14911,N_9842,N_10509);
or U14912 (N_14912,N_10682,N_11401);
and U14913 (N_14913,N_9451,N_11855);
nand U14914 (N_14914,N_10426,N_9748);
nand U14915 (N_14915,N_11464,N_9319);
or U14916 (N_14916,N_11977,N_11236);
nand U14917 (N_14917,N_10216,N_10630);
or U14918 (N_14918,N_9562,N_9728);
and U14919 (N_14919,N_9574,N_9588);
and U14920 (N_14920,N_10638,N_11628);
nand U14921 (N_14921,N_10662,N_9935);
and U14922 (N_14922,N_10879,N_10358);
nand U14923 (N_14923,N_9783,N_11374);
nor U14924 (N_14924,N_9306,N_11530);
nand U14925 (N_14925,N_10700,N_11321);
or U14926 (N_14926,N_11993,N_10973);
nand U14927 (N_14927,N_10825,N_10375);
and U14928 (N_14928,N_11805,N_10897);
or U14929 (N_14929,N_9178,N_9702);
and U14930 (N_14930,N_11624,N_11415);
nand U14931 (N_14931,N_10228,N_11176);
or U14932 (N_14932,N_9579,N_11188);
nor U14933 (N_14933,N_11166,N_9861);
and U14934 (N_14934,N_9013,N_10916);
or U14935 (N_14935,N_9412,N_9718);
and U14936 (N_14936,N_11171,N_9617);
xor U14937 (N_14937,N_10661,N_10756);
or U14938 (N_14938,N_11439,N_9252);
nand U14939 (N_14939,N_9320,N_11897);
nor U14940 (N_14940,N_9170,N_11011);
or U14941 (N_14941,N_10050,N_11648);
nand U14942 (N_14942,N_9784,N_11550);
or U14943 (N_14943,N_9148,N_9625);
nand U14944 (N_14944,N_11168,N_11135);
or U14945 (N_14945,N_10537,N_11609);
nand U14946 (N_14946,N_11794,N_10627);
nand U14947 (N_14947,N_9010,N_9455);
and U14948 (N_14948,N_10442,N_10579);
nor U14949 (N_14949,N_11895,N_9636);
and U14950 (N_14950,N_9219,N_9211);
or U14951 (N_14951,N_10381,N_10060);
nor U14952 (N_14952,N_9270,N_10162);
and U14953 (N_14953,N_11876,N_10531);
nand U14954 (N_14954,N_9841,N_9515);
and U14955 (N_14955,N_11119,N_10264);
nand U14956 (N_14956,N_11007,N_10314);
and U14957 (N_14957,N_11317,N_11110);
nand U14958 (N_14958,N_9980,N_9453);
nand U14959 (N_14959,N_9288,N_11024);
nor U14960 (N_14960,N_9162,N_11569);
nand U14961 (N_14961,N_11053,N_10646);
or U14962 (N_14962,N_10617,N_11241);
nor U14963 (N_14963,N_9944,N_10781);
or U14964 (N_14964,N_11040,N_10734);
nand U14965 (N_14965,N_11958,N_10308);
and U14966 (N_14966,N_9443,N_11655);
or U14967 (N_14967,N_10026,N_10130);
nor U14968 (N_14968,N_9979,N_9246);
nor U14969 (N_14969,N_10084,N_9893);
or U14970 (N_14970,N_9915,N_11960);
nand U14971 (N_14971,N_9831,N_11753);
and U14972 (N_14972,N_11483,N_11384);
or U14973 (N_14973,N_9189,N_11643);
and U14974 (N_14974,N_11055,N_10719);
nor U14975 (N_14975,N_10434,N_11447);
nand U14976 (N_14976,N_9705,N_9289);
and U14977 (N_14977,N_10786,N_10625);
nand U14978 (N_14978,N_11791,N_10823);
and U14979 (N_14979,N_10457,N_10951);
or U14980 (N_14980,N_10287,N_10440);
and U14981 (N_14981,N_10573,N_11624);
nor U14982 (N_14982,N_10529,N_11186);
nand U14983 (N_14983,N_11790,N_9554);
or U14984 (N_14984,N_9296,N_9906);
nor U14985 (N_14985,N_11213,N_9035);
nand U14986 (N_14986,N_10490,N_9259);
nand U14987 (N_14987,N_10072,N_11748);
and U14988 (N_14988,N_9638,N_10774);
nand U14989 (N_14989,N_10913,N_10157);
nand U14990 (N_14990,N_11829,N_9134);
or U14991 (N_14991,N_10475,N_9544);
or U14992 (N_14992,N_11861,N_9456);
or U14993 (N_14993,N_9264,N_11095);
or U14994 (N_14994,N_10083,N_11620);
nor U14995 (N_14995,N_9931,N_9707);
nor U14996 (N_14996,N_10672,N_11126);
nor U14997 (N_14997,N_9997,N_11520);
nand U14998 (N_14998,N_11210,N_10831);
nand U14999 (N_14999,N_11622,N_11958);
nand UO_0 (O_0,N_14282,N_12948);
nand UO_1 (O_1,N_13831,N_12726);
xor UO_2 (O_2,N_12893,N_14267);
nor UO_3 (O_3,N_12698,N_12258);
or UO_4 (O_4,N_12507,N_14692);
nor UO_5 (O_5,N_13094,N_12461);
and UO_6 (O_6,N_12191,N_13272);
or UO_7 (O_7,N_13593,N_14166);
nor UO_8 (O_8,N_14578,N_12694);
and UO_9 (O_9,N_14288,N_14489);
nor UO_10 (O_10,N_12632,N_14758);
and UO_11 (O_11,N_12284,N_13257);
nor UO_12 (O_12,N_13001,N_14082);
or UO_13 (O_13,N_13059,N_14813);
and UO_14 (O_14,N_12285,N_13469);
or UO_15 (O_15,N_14073,N_13218);
nand UO_16 (O_16,N_14897,N_12722);
nor UO_17 (O_17,N_12878,N_14907);
nand UO_18 (O_18,N_13570,N_12394);
nor UO_19 (O_19,N_12445,N_14121);
or UO_20 (O_20,N_13173,N_14273);
and UO_21 (O_21,N_13460,N_14732);
and UO_22 (O_22,N_12424,N_12660);
and UO_23 (O_23,N_12491,N_12506);
nor UO_24 (O_24,N_13418,N_14217);
nand UO_25 (O_25,N_12370,N_13387);
nand UO_26 (O_26,N_14490,N_12346);
nor UO_27 (O_27,N_13860,N_13800);
nor UO_28 (O_28,N_14803,N_14629);
nor UO_29 (O_29,N_14967,N_14355);
nand UO_30 (O_30,N_14548,N_12876);
nand UO_31 (O_31,N_13102,N_14036);
nand UO_32 (O_32,N_14475,N_12431);
and UO_33 (O_33,N_12044,N_13176);
nor UO_34 (O_34,N_12655,N_14038);
or UO_35 (O_35,N_12913,N_12451);
or UO_36 (O_36,N_13214,N_14942);
nand UO_37 (O_37,N_14497,N_14766);
nand UO_38 (O_38,N_12832,N_14191);
and UO_39 (O_39,N_14078,N_12155);
and UO_40 (O_40,N_14672,N_12756);
and UO_41 (O_41,N_12412,N_12686);
and UO_42 (O_42,N_12669,N_14301);
and UO_43 (O_43,N_13975,N_12723);
nand UO_44 (O_44,N_13522,N_12077);
or UO_45 (O_45,N_13091,N_14498);
nand UO_46 (O_46,N_14914,N_14583);
nand UO_47 (O_47,N_13133,N_14248);
or UO_48 (O_48,N_13096,N_12217);
nor UO_49 (O_49,N_14747,N_13380);
nand UO_50 (O_50,N_13752,N_13519);
nand UO_51 (O_51,N_14581,N_14561);
nand UO_52 (O_52,N_13347,N_13857);
nand UO_53 (O_53,N_12634,N_12513);
and UO_54 (O_54,N_13787,N_14620);
xor UO_55 (O_55,N_13164,N_12956);
nand UO_56 (O_56,N_13285,N_12069);
or UO_57 (O_57,N_13103,N_14249);
nor UO_58 (O_58,N_12001,N_13117);
nand UO_59 (O_59,N_13234,N_12021);
or UO_60 (O_60,N_12706,N_12964);
and UO_61 (O_61,N_13331,N_13660);
and UO_62 (O_62,N_14253,N_12281);
nor UO_63 (O_63,N_12314,N_14387);
or UO_64 (O_64,N_14095,N_13672);
xnor UO_65 (O_65,N_12407,N_12817);
nor UO_66 (O_66,N_12218,N_12159);
or UO_67 (O_67,N_14965,N_14409);
and UO_68 (O_68,N_12958,N_13303);
and UO_69 (O_69,N_14065,N_14171);
and UO_70 (O_70,N_12846,N_14389);
and UO_71 (O_71,N_13187,N_13210);
or UO_72 (O_72,N_12869,N_12783);
nor UO_73 (O_73,N_12758,N_12481);
and UO_74 (O_74,N_13410,N_12633);
and UO_75 (O_75,N_13919,N_12983);
or UO_76 (O_76,N_13815,N_13475);
or UO_77 (O_77,N_13918,N_14087);
and UO_78 (O_78,N_12170,N_13360);
or UO_79 (O_79,N_13119,N_13172);
nand UO_80 (O_80,N_12172,N_14710);
nor UO_81 (O_81,N_13627,N_14990);
or UO_82 (O_82,N_12049,N_13629);
or UO_83 (O_83,N_14635,N_13625);
nor UO_84 (O_84,N_12564,N_14882);
and UO_85 (O_85,N_12204,N_12608);
nor UO_86 (O_86,N_14901,N_14983);
or UO_87 (O_87,N_14592,N_13146);
nor UO_88 (O_88,N_13706,N_14568);
and UO_89 (O_89,N_12676,N_14039);
and UO_90 (O_90,N_13022,N_12476);
and UO_91 (O_91,N_14450,N_12656);
nand UO_92 (O_92,N_14676,N_12363);
and UO_93 (O_93,N_13619,N_12561);
nor UO_94 (O_94,N_14064,N_12436);
and UO_95 (O_95,N_13808,N_13614);
nor UO_96 (O_96,N_13048,N_13714);
and UO_97 (O_97,N_12068,N_14091);
nor UO_98 (O_98,N_13878,N_12665);
nor UO_99 (O_99,N_14595,N_13306);
and UO_100 (O_100,N_14812,N_14216);
or UO_101 (O_101,N_14247,N_14778);
and UO_102 (O_102,N_13325,N_12724);
and UO_103 (O_103,N_14051,N_13192);
and UO_104 (O_104,N_13058,N_12425);
or UO_105 (O_105,N_14337,N_12764);
or UO_106 (O_106,N_14430,N_13830);
and UO_107 (O_107,N_13236,N_12496);
or UO_108 (O_108,N_13676,N_12442);
or UO_109 (O_109,N_13940,N_14846);
nor UO_110 (O_110,N_12975,N_14896);
nand UO_111 (O_111,N_12380,N_14440);
nor UO_112 (O_112,N_12057,N_13177);
and UO_113 (O_113,N_12969,N_13917);
and UO_114 (O_114,N_12587,N_13602);
nand UO_115 (O_115,N_12345,N_13631);
nand UO_116 (O_116,N_14514,N_12508);
nand UO_117 (O_117,N_14386,N_13992);
and UO_118 (O_118,N_14843,N_14239);
or UO_119 (O_119,N_14571,N_13204);
nand UO_120 (O_120,N_14610,N_14969);
or UO_121 (O_121,N_13350,N_14099);
nand UO_122 (O_122,N_12470,N_14259);
or UO_123 (O_123,N_14853,N_14458);
and UO_124 (O_124,N_14176,N_14344);
or UO_125 (O_125,N_14600,N_14545);
nor UO_126 (O_126,N_13559,N_12158);
or UO_127 (O_127,N_12238,N_12937);
or UO_128 (O_128,N_13926,N_14984);
and UO_129 (O_129,N_12965,N_13092);
nand UO_130 (O_130,N_13948,N_14372);
or UO_131 (O_131,N_14512,N_13757);
or UO_132 (O_132,N_13729,N_12884);
nor UO_133 (O_133,N_13216,N_13265);
nand UO_134 (O_134,N_13313,N_12213);
and UO_135 (O_135,N_12031,N_13343);
and UO_136 (O_136,N_13376,N_13184);
and UO_137 (O_137,N_14981,N_13338);
and UO_138 (O_138,N_13613,N_14768);
or UO_139 (O_139,N_12701,N_14238);
or UO_140 (O_140,N_13320,N_13888);
nand UO_141 (O_141,N_12984,N_14560);
nand UO_142 (O_142,N_12120,N_12798);
nand UO_143 (O_143,N_12458,N_12991);
and UO_144 (O_144,N_12544,N_13244);
and UO_145 (O_145,N_13209,N_14013);
nand UO_146 (O_146,N_14636,N_12672);
and UO_147 (O_147,N_14360,N_12328);
nor UO_148 (O_148,N_13561,N_13299);
and UO_149 (O_149,N_14689,N_13984);
nor UO_150 (O_150,N_14056,N_14009);
nand UO_151 (O_151,N_13304,N_13776);
or UO_152 (O_152,N_14417,N_12611);
nor UO_153 (O_153,N_12418,N_13771);
nand UO_154 (O_154,N_13828,N_14502);
nand UO_155 (O_155,N_14885,N_14791);
and UO_156 (O_156,N_13390,N_14572);
nand UO_157 (O_157,N_12624,N_14619);
and UO_158 (O_158,N_14993,N_13007);
or UO_159 (O_159,N_13267,N_12304);
or UO_160 (O_160,N_14785,N_14991);
and UO_161 (O_161,N_13950,N_14305);
nand UO_162 (O_162,N_12319,N_12560);
and UO_163 (O_163,N_14938,N_13520);
or UO_164 (O_164,N_14648,N_13314);
nor UO_165 (O_165,N_13993,N_13795);
nand UO_166 (O_166,N_14792,N_13716);
or UO_167 (O_167,N_12820,N_12171);
and UO_168 (O_168,N_12322,N_14264);
nor UO_169 (O_169,N_14613,N_13446);
nor UO_170 (O_170,N_12642,N_13741);
or UO_171 (O_171,N_12121,N_12497);
nand UO_172 (O_172,N_13862,N_14102);
and UO_173 (O_173,N_13889,N_14204);
nand UO_174 (O_174,N_13089,N_13689);
nor UO_175 (O_175,N_14042,N_12145);
nand UO_176 (O_176,N_14043,N_14839);
nor UO_177 (O_177,N_13432,N_14870);
and UO_178 (O_178,N_12678,N_13363);
nand UO_179 (O_179,N_13675,N_12742);
or UO_180 (O_180,N_12105,N_13989);
or UO_181 (O_181,N_13999,N_13219);
and UO_182 (O_182,N_12427,N_13324);
and UO_183 (O_183,N_13786,N_13105);
nand UO_184 (O_184,N_13620,N_12657);
or UO_185 (O_185,N_14281,N_12341);
nand UO_186 (O_186,N_13130,N_14531);
nand UO_187 (O_187,N_14989,N_12428);
nor UO_188 (O_188,N_12510,N_12840);
nand UO_189 (O_189,N_14861,N_14678);
nor UO_190 (O_190,N_14866,N_14992);
nor UO_191 (O_191,N_13849,N_14006);
nand UO_192 (O_192,N_14937,N_14765);
and UO_193 (O_193,N_14149,N_12269);
xor UO_194 (O_194,N_14911,N_14887);
and UO_195 (O_195,N_13052,N_13760);
nand UO_196 (O_196,N_12162,N_14685);
or UO_197 (O_197,N_13928,N_12195);
and UO_198 (O_198,N_13093,N_12233);
nor UO_199 (O_199,N_13990,N_13384);
nor UO_200 (O_200,N_13241,N_12810);
and UO_201 (O_201,N_14585,N_13822);
nor UO_202 (O_202,N_13348,N_12192);
nor UO_203 (O_203,N_12602,N_13077);
nor UO_204 (O_204,N_12762,N_12550);
or UO_205 (O_205,N_12229,N_12264);
nand UO_206 (O_206,N_12531,N_13796);
and UO_207 (O_207,N_14432,N_12457);
nand UO_208 (O_208,N_14977,N_14284);
nor UO_209 (O_209,N_14342,N_12179);
nor UO_210 (O_210,N_14564,N_13047);
nand UO_211 (O_211,N_14256,N_14873);
nand UO_212 (O_212,N_12467,N_14123);
and UO_213 (O_213,N_14225,N_13755);
nor UO_214 (O_214,N_14241,N_13974);
nand UO_215 (O_215,N_12640,N_14903);
nor UO_216 (O_216,N_13886,N_13961);
and UO_217 (O_217,N_14963,N_12901);
nand UO_218 (O_218,N_13339,N_13353);
nor UO_219 (O_219,N_14328,N_12551);
nor UO_220 (O_220,N_12148,N_14665);
nand UO_221 (O_221,N_12117,N_14508);
and UO_222 (O_222,N_13083,N_13226);
nand UO_223 (O_223,N_14606,N_12851);
nand UO_224 (O_224,N_14702,N_13767);
nor UO_225 (O_225,N_13044,N_14031);
and UO_226 (O_226,N_13062,N_13066);
or UO_227 (O_227,N_13557,N_12912);
nand UO_228 (O_228,N_14515,N_14669);
and UO_229 (O_229,N_12957,N_14666);
and UO_230 (O_230,N_13289,N_13663);
or UO_231 (O_231,N_14876,N_12881);
or UO_232 (O_232,N_12146,N_12946);
xnor UO_233 (O_233,N_13232,N_14567);
or UO_234 (O_234,N_13869,N_14913);
nand UO_235 (O_235,N_13131,N_12244);
nand UO_236 (O_236,N_12711,N_12525);
and UO_237 (O_237,N_12997,N_14457);
and UO_238 (O_238,N_13742,N_14308);
and UO_239 (O_239,N_13169,N_13791);
nand UO_240 (O_240,N_13259,N_14940);
and UO_241 (O_241,N_13581,N_14001);
nand UO_242 (O_242,N_13161,N_14173);
xor UO_243 (O_243,N_13401,N_14811);
nor UO_244 (O_244,N_12278,N_14598);
or UO_245 (O_245,N_12393,N_13181);
nor UO_246 (O_246,N_14334,N_14005);
nor UO_247 (O_247,N_14032,N_14010);
nor UO_248 (O_248,N_12230,N_12520);
nor UO_249 (O_249,N_12571,N_12708);
and UO_250 (O_250,N_13027,N_13690);
nand UO_251 (O_251,N_13158,N_13197);
nand UO_252 (O_252,N_13175,N_12422);
nor UO_253 (O_253,N_12921,N_12466);
nor UO_254 (O_254,N_12562,N_13877);
nor UO_255 (O_255,N_14319,N_12592);
or UO_256 (O_256,N_13659,N_14451);
or UO_257 (O_257,N_14017,N_12241);
nor UO_258 (O_258,N_13108,N_14162);
and UO_259 (O_259,N_12329,N_14482);
nand UO_260 (O_260,N_14202,N_14733);
nand UO_261 (O_261,N_12088,N_12201);
nand UO_262 (O_262,N_14760,N_14639);
nor UO_263 (O_263,N_14607,N_14327);
nand UO_264 (O_264,N_14879,N_14975);
and UO_265 (O_265,N_13318,N_13517);
nand UO_266 (O_266,N_14071,N_13621);
and UO_267 (O_267,N_13275,N_13142);
nand UO_268 (O_268,N_13769,N_12149);
and UO_269 (O_269,N_12749,N_14226);
nor UO_270 (O_270,N_14467,N_13424);
or UO_271 (O_271,N_14605,N_14452);
nand UO_272 (O_272,N_13407,N_13470);
or UO_273 (O_273,N_12164,N_14856);
and UO_274 (O_274,N_13650,N_13783);
or UO_275 (O_275,N_13703,N_14054);
and UO_276 (O_276,N_13431,N_14426);
nand UO_277 (O_277,N_14357,N_14481);
or UO_278 (O_278,N_13388,N_14019);
nor UO_279 (O_279,N_14033,N_12070);
nor UO_280 (O_280,N_14686,N_12400);
nand UO_281 (O_281,N_12033,N_12081);
nand UO_282 (O_282,N_13827,N_12863);
and UO_283 (O_283,N_13647,N_13977);
or UO_284 (O_284,N_13588,N_12440);
nand UO_285 (O_285,N_14961,N_13435);
nor UO_286 (O_286,N_12821,N_13101);
or UO_287 (O_287,N_12740,N_12260);
or UO_288 (O_288,N_14401,N_12504);
and UO_289 (O_289,N_12653,N_13558);
or UO_290 (O_290,N_14919,N_12927);
nor UO_291 (O_291,N_14850,N_12514);
nor UO_292 (O_292,N_13897,N_13991);
nor UO_293 (O_293,N_13834,N_14931);
nand UO_294 (O_294,N_12659,N_12778);
and UO_295 (O_295,N_12537,N_14004);
and UO_296 (O_296,N_13549,N_14077);
and UO_297 (O_297,N_13213,N_13768);
or UO_298 (O_298,N_12344,N_13321);
and UO_299 (O_299,N_12209,N_12112);
nor UO_300 (O_300,N_12011,N_12649);
or UO_301 (O_301,N_14047,N_14706);
nor UO_302 (O_302,N_12478,N_12986);
nor UO_303 (O_303,N_13514,N_14845);
nand UO_304 (O_304,N_12459,N_14982);
nand UO_305 (O_305,N_13453,N_13429);
and UO_306 (O_306,N_13262,N_14194);
nand UO_307 (O_307,N_14858,N_12035);
or UO_308 (O_308,N_13692,N_13616);
or UO_309 (O_309,N_14464,N_13296);
nor UO_310 (O_310,N_12046,N_12480);
and UO_311 (O_311,N_13641,N_12372);
or UO_312 (O_312,N_13451,N_13775);
or UO_313 (O_313,N_14245,N_13139);
and UO_314 (O_314,N_12861,N_14820);
and UO_315 (O_315,N_14278,N_12430);
and UO_316 (O_316,N_14641,N_13811);
nand UO_317 (O_317,N_14966,N_12833);
nor UO_318 (O_318,N_14011,N_12064);
nand UO_319 (O_319,N_14331,N_13594);
nor UO_320 (O_320,N_12239,N_14111);
or UO_321 (O_321,N_12194,N_14721);
and UO_322 (O_322,N_13894,N_12890);
nand UO_323 (O_323,N_14045,N_13615);
and UO_324 (O_324,N_12111,N_14024);
nand UO_325 (O_325,N_12596,N_14129);
and UO_326 (O_326,N_13686,N_14616);
and UO_327 (O_327,N_12809,N_13053);
nand UO_328 (O_328,N_13399,N_13893);
or UO_329 (O_329,N_12133,N_12962);
nor UO_330 (O_330,N_14591,N_14987);
or UO_331 (O_331,N_14941,N_12588);
or UO_332 (O_332,N_14016,N_12736);
nand UO_333 (O_333,N_13070,N_12570);
and UO_334 (O_334,N_12763,N_14872);
and UO_335 (O_335,N_13400,N_13402);
and UO_336 (O_336,N_14729,N_14418);
or UO_337 (O_337,N_12293,N_13416);
or UO_338 (O_338,N_12384,N_13736);
nand UO_339 (O_339,N_13719,N_13705);
nand UO_340 (O_340,N_12565,N_13605);
and UO_341 (O_341,N_13854,N_14549);
or UO_342 (O_342,N_13847,N_14754);
nand UO_343 (O_343,N_14974,N_12774);
and UO_344 (O_344,N_14378,N_14465);
nand UO_345 (O_345,N_13334,N_12186);
and UO_346 (O_346,N_14518,N_14220);
nor UO_347 (O_347,N_13088,N_13927);
and UO_348 (O_348,N_14207,N_12794);
or UO_349 (O_349,N_12853,N_12801);
nand UO_350 (O_350,N_14246,N_13525);
nor UO_351 (O_351,N_14783,N_12323);
or UO_352 (O_352,N_14761,N_14716);
or UO_353 (O_353,N_12073,N_13954);
nand UO_354 (O_354,N_14155,N_13297);
and UO_355 (O_355,N_13511,N_13646);
or UO_356 (O_356,N_13507,N_13700);
or UO_357 (O_357,N_13978,N_13987);
nor UO_358 (O_358,N_13589,N_13931);
or UO_359 (O_359,N_12808,N_14103);
nand UO_360 (O_360,N_12232,N_12482);
or UO_361 (O_361,N_12301,N_13277);
and UO_362 (O_362,N_12242,N_14838);
or UO_363 (O_363,N_14244,N_12787);
nor UO_364 (O_364,N_13601,N_14623);
nor UO_365 (O_365,N_13753,N_12750);
nand UO_366 (O_366,N_12932,N_13821);
or UO_367 (O_367,N_12718,N_13471);
xnor UO_368 (O_368,N_12292,N_12362);
and UO_369 (O_369,N_13668,N_13064);
or UO_370 (O_370,N_12594,N_13555);
nor UO_371 (O_371,N_13098,N_13493);
nand UO_372 (O_372,N_14526,N_14384);
nand UO_373 (O_373,N_14924,N_13282);
nor UO_374 (O_374,N_13150,N_13191);
and UO_375 (O_375,N_13051,N_14088);
nand UO_376 (O_376,N_14898,N_12777);
or UO_377 (O_377,N_14435,N_12388);
and UO_378 (O_378,N_13712,N_12533);
xor UO_379 (O_379,N_13127,N_12545);
and UO_380 (O_380,N_13566,N_13071);
nor UO_381 (O_381,N_14317,N_14883);
or UO_382 (O_382,N_13042,N_12006);
nand UO_383 (O_383,N_13569,N_12169);
nor UO_384 (O_384,N_13916,N_14958);
nor UO_385 (O_385,N_14664,N_13134);
and UO_386 (O_386,N_12308,N_12943);
nor UO_387 (O_387,N_14988,N_13554);
nand UO_388 (O_388,N_13655,N_12004);
nor UO_389 (O_389,N_13009,N_14090);
and UO_390 (O_390,N_13844,N_14014);
nand UO_391 (O_391,N_12167,N_13495);
nor UO_392 (O_392,N_13415,N_13510);
or UO_393 (O_393,N_13693,N_14611);
and UO_394 (O_394,N_12406,N_14737);
nor UO_395 (O_395,N_14133,N_13899);
nor UO_396 (O_396,N_14260,N_14744);
nand UO_397 (O_397,N_14651,N_14849);
nand UO_398 (O_398,N_13112,N_14841);
or UO_399 (O_399,N_14832,N_14139);
nor UO_400 (O_400,N_12036,N_12931);
nor UO_401 (O_401,N_14848,N_13190);
or UO_402 (O_402,N_13374,N_13669);
nand UO_403 (O_403,N_13372,N_13643);
and UO_404 (O_404,N_12432,N_14823);
nand UO_405 (O_405,N_13015,N_13163);
xor UO_406 (O_406,N_13368,N_14799);
nor UO_407 (O_407,N_12168,N_14169);
nor UO_408 (O_408,N_13801,N_13509);
nand UO_409 (O_409,N_13361,N_13281);
nor UO_410 (O_410,N_14151,N_13963);
and UO_411 (O_411,N_14622,N_14801);
and UO_412 (O_412,N_13033,N_13385);
nor UO_413 (O_413,N_12843,N_13486);
and UO_414 (O_414,N_13463,N_14892);
nor UO_415 (O_415,N_13002,N_14098);
and UO_416 (O_416,N_14910,N_14356);
nor UO_417 (O_417,N_13707,N_12536);
nand UO_418 (O_418,N_14684,N_14478);
and UO_419 (O_419,N_14617,N_14730);
nand UO_420 (O_420,N_12741,N_14309);
and UO_421 (O_421,N_12748,N_14057);
or UO_422 (O_422,N_13538,N_14347);
and UO_423 (O_423,N_13573,N_14240);
nor UO_424 (O_424,N_12099,N_14373);
nand UO_425 (O_425,N_13922,N_13503);
nand UO_426 (O_426,N_13872,N_13995);
or UO_427 (O_427,N_14985,N_13254);
or UO_428 (O_428,N_12612,N_14302);
nand UO_429 (O_429,N_14330,N_13125);
or UO_430 (O_430,N_12267,N_12548);
and UO_431 (O_431,N_14303,N_12096);
nor UO_432 (O_432,N_14696,N_12027);
nor UO_433 (O_433,N_13651,N_13779);
and UO_434 (O_434,N_14724,N_13260);
and UO_435 (O_435,N_12039,N_14780);
nand UO_436 (O_436,N_14703,N_12371);
and UO_437 (O_437,N_12617,N_12631);
nand UO_438 (O_438,N_14816,N_12176);
or UO_439 (O_439,N_13207,N_14637);
and UO_440 (O_440,N_12381,N_12349);
and UO_441 (O_441,N_14135,N_13017);
nor UO_442 (O_442,N_12993,N_12343);
and UO_443 (O_443,N_12091,N_13711);
nor UO_444 (O_444,N_12391,N_13206);
nand UO_445 (O_445,N_14973,N_12223);
nand UO_446 (O_446,N_12063,N_13667);
nor UO_447 (O_447,N_13049,N_14343);
and UO_448 (O_448,N_12834,N_12585);
or UO_449 (O_449,N_14749,N_14723);
or UO_450 (O_450,N_12187,N_14424);
and UO_451 (O_451,N_13344,N_13225);
and UO_452 (O_452,N_12463,N_14537);
nand UO_453 (O_453,N_14367,N_13898);
nand UO_454 (O_454,N_12203,N_12788);
nand UO_455 (O_455,N_14374,N_14609);
and UO_456 (O_456,N_14211,N_13936);
and UO_457 (O_457,N_12386,N_13300);
nor UO_458 (O_458,N_14423,N_13247);
or UO_459 (O_459,N_14370,N_13544);
nand UO_460 (O_460,N_12735,N_14037);
or UO_461 (O_461,N_14881,N_13542);
nand UO_462 (O_462,N_13883,N_12009);
and UO_463 (O_463,N_13080,N_13696);
nand UO_464 (O_464,N_14986,N_14945);
or UO_465 (O_465,N_14626,N_12909);
or UO_466 (O_466,N_12423,N_12212);
nor UO_467 (O_467,N_13996,N_14270);
or UO_468 (O_468,N_14053,N_12591);
and UO_469 (O_469,N_14510,N_14385);
and UO_470 (O_470,N_13205,N_13654);
nor UO_471 (O_471,N_13737,N_14884);
nor UO_472 (O_472,N_12572,N_12226);
nor UO_473 (O_473,N_12206,N_12517);
and UO_474 (O_474,N_12829,N_14833);
nand UO_475 (O_475,N_13761,N_13312);
or UO_476 (O_476,N_12673,N_14486);
nand UO_477 (O_477,N_14840,N_12252);
nor UO_478 (O_478,N_13371,N_13732);
xnor UO_479 (O_479,N_14955,N_13104);
or UO_480 (O_480,N_12717,N_12056);
and UO_481 (O_481,N_13426,N_12523);
and UO_482 (O_482,N_13807,N_14679);
and UO_483 (O_483,N_12920,N_13114);
nand UO_484 (O_484,N_12126,N_12732);
nand UO_485 (O_485,N_13307,N_14500);
nor UO_486 (O_486,N_13684,N_13452);
nor UO_487 (O_487,N_13118,N_13905);
or UO_488 (O_488,N_14871,N_13496);
nor UO_489 (O_489,N_13656,N_13797);
and UO_490 (O_490,N_14081,N_12435);
or UO_491 (O_491,N_13208,N_14142);
nor UO_492 (O_492,N_13870,N_12390);
or UO_493 (O_493,N_12397,N_12988);
or UO_494 (O_494,N_14704,N_12526);
nand UO_495 (O_495,N_13095,N_14741);
and UO_496 (O_496,N_14757,N_12101);
xnor UO_497 (O_497,N_13082,N_12154);
nor UO_498 (O_498,N_12488,N_12302);
and UO_499 (O_499,N_12376,N_14891);
or UO_500 (O_500,N_12468,N_12198);
or UO_501 (O_501,N_14709,N_12689);
and UO_502 (O_502,N_12879,N_14713);
or UO_503 (O_503,N_13280,N_13358);
and UO_504 (O_504,N_14563,N_13292);
nor UO_505 (O_505,N_13653,N_12803);
nand UO_506 (O_506,N_12464,N_13227);
or UO_507 (O_507,N_12753,N_12651);
nand UO_508 (O_508,N_14376,N_13512);
and UO_509 (O_509,N_12874,N_14122);
or UO_510 (O_510,N_14770,N_13043);
nand UO_511 (O_511,N_14493,N_12797);
nor UO_512 (O_512,N_13938,N_13739);
and UO_513 (O_513,N_14283,N_12306);
or UO_514 (O_514,N_14154,N_14864);
nor UO_515 (O_515,N_14677,N_14285);
nand UO_516 (O_516,N_13516,N_13523);
nor UO_517 (O_517,N_13110,N_13481);
or UO_518 (O_518,N_14925,N_12950);
and UO_519 (O_519,N_12528,N_13930);
nand UO_520 (O_520,N_13381,N_14738);
and UO_521 (O_521,N_13147,N_12297);
nor UO_522 (O_522,N_14772,N_13454);
nand UO_523 (O_523,N_14000,N_13547);
nand UO_524 (O_524,N_12043,N_13245);
and UO_525 (O_525,N_14559,N_13962);
or UO_526 (O_526,N_12502,N_13682);
nand UO_527 (O_527,N_12581,N_14597);
nor UO_528 (O_528,N_13445,N_14405);
and UO_529 (O_529,N_13162,N_14003);
nand UO_530 (O_530,N_12288,N_13240);
or UO_531 (O_531,N_14735,N_14353);
or UO_532 (O_532,N_14177,N_14008);
and UO_533 (O_533,N_12967,N_12348);
nor UO_534 (O_534,N_12826,N_12462);
or UO_535 (O_535,N_12791,N_12013);
nand UO_536 (O_536,N_12650,N_12981);
and UO_537 (O_537,N_14124,N_14449);
or UO_538 (O_538,N_14059,N_12871);
or UO_539 (O_539,N_14854,N_13909);
nor UO_540 (O_540,N_12253,N_13759);
nand UO_541 (O_541,N_14711,N_12320);
nor UO_542 (O_542,N_12107,N_14773);
nand UO_543 (O_543,N_13305,N_12854);
and UO_544 (O_544,N_12116,N_12702);
and UO_545 (O_545,N_14222,N_13490);
and UO_546 (O_546,N_12939,N_13274);
nor UO_547 (O_547,N_14543,N_14119);
or UO_548 (O_548,N_14048,N_12709);
and UO_549 (O_549,N_12438,N_12755);
or UO_550 (O_550,N_12163,N_14774);
and UO_551 (O_551,N_13998,N_12729);
nor UO_552 (O_552,N_13489,N_14532);
and UO_553 (O_553,N_14690,N_12141);
and UO_554 (O_554,N_13021,N_12799);
nand UO_555 (O_555,N_12477,N_13423);
nand UO_556 (O_556,N_12350,N_14752);
and UO_557 (O_557,N_14137,N_13784);
or UO_558 (O_558,N_12225,N_12305);
nand UO_559 (O_559,N_14215,N_13580);
nor UO_560 (O_560,N_12471,N_13140);
and UO_561 (O_561,N_12772,N_12638);
nand UO_562 (O_562,N_14821,N_13935);
and UO_563 (O_563,N_14668,N_13957);
or UO_564 (O_564,N_13369,N_13541);
or UO_565 (O_565,N_12614,N_14455);
and UO_566 (O_566,N_14022,N_12910);
and UO_567 (O_567,N_13546,N_13328);
nand UO_568 (O_568,N_12752,N_12365);
and UO_569 (O_569,N_13268,N_14759);
or UO_570 (O_570,N_13604,N_13107);
nor UO_571 (O_571,N_14717,N_13461);
nand UO_572 (O_572,N_14573,N_13330);
or UO_573 (O_573,N_12222,N_13953);
or UO_574 (O_574,N_13242,N_12016);
or UO_575 (O_575,N_14277,N_14740);
nand UO_576 (O_576,N_13124,N_12535);
or UO_577 (O_577,N_14999,N_14391);
and UO_578 (O_578,N_14371,N_12071);
nand UO_579 (O_579,N_12818,N_13421);
nor UO_580 (O_580,N_14203,N_12746);
or UO_581 (O_581,N_13840,N_13911);
nor UO_582 (O_582,N_12886,N_13430);
or UO_583 (O_583,N_14701,N_14818);
nor UO_584 (O_584,N_14186,N_13763);
nand UO_585 (O_585,N_12093,N_14496);
or UO_586 (O_586,N_14025,N_13032);
nand UO_587 (O_587,N_13626,N_14547);
nand UO_588 (O_588,N_13061,N_13717);
nand UO_589 (O_589,N_13859,N_12625);
nand UO_590 (O_590,N_13988,N_12613);
nor UO_591 (O_591,N_13266,N_12351);
nor UO_592 (O_592,N_13725,N_13195);
or UO_593 (O_593,N_14831,N_12739);
and UO_594 (O_594,N_12254,N_12483);
xnor UO_595 (O_595,N_13960,N_13074);
or UO_596 (O_596,N_14089,N_12237);
nand UO_597 (O_597,N_12999,N_12547);
nor UO_598 (O_598,N_12161,N_14243);
nor UO_599 (O_599,N_14590,N_12796);
nand UO_600 (O_600,N_13476,N_13762);
nand UO_601 (O_601,N_13342,N_14113);
nand UO_602 (O_602,N_14187,N_13835);
and UO_603 (O_603,N_14300,N_12361);
nor UO_604 (O_604,N_12900,N_12490);
or UO_605 (O_605,N_12472,N_12479);
nand UO_606 (O_606,N_14175,N_13636);
nand UO_607 (O_607,N_13290,N_14809);
or UO_608 (O_608,N_13772,N_12555);
nand UO_609 (O_609,N_13271,N_14847);
nor UO_610 (O_610,N_12845,N_12715);
nor UO_611 (O_611,N_14380,N_14228);
and UO_612 (O_612,N_13749,N_12012);
nor UO_613 (O_613,N_13167,N_14654);
nor UO_614 (O_614,N_12693,N_14462);
nor UO_615 (O_615,N_13720,N_12054);
nand UO_616 (O_616,N_12682,N_14978);
or UO_617 (O_617,N_14921,N_14638);
nor UO_618 (O_618,N_13582,N_13518);
and UO_619 (O_619,N_14511,N_14555);
nor UO_620 (O_620,N_14979,N_13097);
and UO_621 (O_621,N_13011,N_13188);
and UO_622 (O_622,N_12247,N_14063);
nand UO_623 (O_623,N_14787,N_12289);
and UO_624 (O_624,N_12994,N_14437);
and UO_625 (O_625,N_12335,N_14698);
or UO_626 (O_626,N_12662,N_14888);
nor UO_627 (O_627,N_13329,N_13805);
nand UO_628 (O_628,N_14232,N_14425);
nand UO_629 (O_629,N_13237,N_12731);
and UO_630 (O_630,N_12971,N_14310);
nor UO_631 (O_631,N_12727,N_13456);
nor UO_632 (O_632,N_14096,N_12804);
nand UO_633 (O_633,N_14525,N_13311);
and UO_634 (O_634,N_13144,N_14414);
and UO_635 (O_635,N_12737,N_14722);
nand UO_636 (O_636,N_14867,N_12103);
nand UO_637 (O_637,N_14516,N_14649);
or UO_638 (O_638,N_12474,N_13644);
nor UO_639 (O_639,N_13484,N_13864);
nor UO_640 (O_640,N_12277,N_12705);
and UO_641 (O_641,N_12949,N_14134);
or UO_642 (O_642,N_13848,N_13825);
nand UO_643 (O_643,N_13947,N_14851);
nor UO_644 (O_644,N_13906,N_14381);
nor UO_645 (O_645,N_13332,N_13501);
nand UO_646 (O_646,N_12664,N_13068);
and UO_647 (O_647,N_12100,N_13843);
nor UO_648 (O_648,N_12963,N_13944);
nor UO_649 (O_649,N_14562,N_12626);
nand UO_650 (O_650,N_12897,N_13069);
nor UO_651 (O_651,N_14052,N_14807);
and UO_652 (O_652,N_14411,N_13436);
nor UO_653 (O_653,N_14815,N_12529);
nand UO_654 (O_654,N_13160,N_13592);
nor UO_655 (O_655,N_14050,N_12398);
and UO_656 (O_656,N_12211,N_14108);
and UO_657 (O_657,N_12885,N_14029);
nand UO_658 (O_658,N_13224,N_12867);
xnor UO_659 (O_659,N_14970,N_13536);
or UO_660 (O_660,N_12800,N_14200);
nor UO_661 (O_661,N_14307,N_12118);
or UO_662 (O_662,N_13976,N_12639);
nand UO_663 (O_663,N_12152,N_14551);
nor UO_664 (O_664,N_13661,N_14822);
or UO_665 (O_665,N_12272,N_12839);
nor UO_666 (O_666,N_12954,N_12903);
or UO_667 (O_667,N_14530,N_14196);
or UO_668 (O_668,N_13740,N_13099);
nand UO_669 (O_669,N_12907,N_13276);
and UO_670 (O_670,N_12697,N_13852);
or UO_671 (O_671,N_13585,N_14201);
nand UO_672 (O_672,N_14322,N_12973);
or UO_673 (O_673,N_12844,N_13478);
nand UO_674 (O_674,N_14026,N_14960);
nand UO_675 (O_675,N_13386,N_12316);
nor UO_676 (O_676,N_12002,N_14643);
nor UO_677 (O_677,N_12864,N_14333);
nor UO_678 (O_678,N_14923,N_13803);
and UO_679 (O_679,N_14115,N_14209);
nor UO_680 (O_680,N_12008,N_12875);
and UO_681 (O_681,N_14157,N_13462);
and UO_682 (O_682,N_12299,N_13395);
nand UO_683 (O_683,N_14136,N_14265);
xnor UO_684 (O_684,N_13466,N_12607);
and UO_685 (O_685,N_14292,N_14902);
nand UO_686 (O_686,N_13364,N_13437);
xnor UO_687 (O_687,N_13038,N_14295);
or UO_688 (O_688,N_14601,N_14436);
nor UO_689 (O_689,N_12872,N_14379);
nand UO_690 (O_690,N_12034,N_14316);
nand UO_691 (O_691,N_13050,N_14614);
or UO_692 (O_692,N_12977,N_13359);
nand UO_693 (O_693,N_12786,N_12790);
nor UO_694 (O_694,N_14060,N_14030);
nor UO_695 (O_695,N_12029,N_13551);
and UO_696 (O_696,N_12865,N_13157);
or UO_697 (O_697,N_13850,N_12644);
and UO_698 (O_698,N_12618,N_12360);
or UO_699 (O_699,N_13724,N_13008);
and UO_700 (O_700,N_13004,N_13326);
and UO_701 (O_701,N_13562,N_12894);
and UO_702 (O_702,N_12603,N_13041);
or UO_703 (O_703,N_13081,N_12899);
and UO_704 (O_704,N_13243,N_13836);
or UO_705 (O_705,N_12645,N_13599);
or UO_706 (O_706,N_13201,N_13617);
and UO_707 (O_707,N_13315,N_13873);
or UO_708 (O_708,N_12147,N_14213);
or UO_709 (O_709,N_14165,N_14361);
nor UO_710 (O_710,N_14527,N_12714);
nor UO_711 (O_711,N_12024,N_13316);
nor UO_712 (O_712,N_14459,N_13648);
nand UO_713 (O_713,N_13751,N_14427);
or UO_714 (O_714,N_14350,N_14582);
nand UO_715 (O_715,N_14181,N_13174);
nor UO_716 (O_716,N_12761,N_14105);
or UO_717 (O_717,N_14140,N_14900);
and UO_718 (O_718,N_14229,N_13483);
nor UO_719 (O_719,N_14326,N_14494);
nand UO_720 (O_720,N_13657,N_12530);
nand UO_721 (O_721,N_12266,N_12415);
and UO_722 (O_722,N_14577,N_14068);
nand UO_723 (O_723,N_13447,N_12926);
nor UO_724 (O_724,N_12569,N_13392);
and UO_725 (O_725,N_13718,N_12989);
and UO_726 (O_726,N_14148,N_13346);
nand UO_727 (O_727,N_13055,N_13393);
or UO_728 (O_728,N_13945,N_14167);
or UO_729 (O_729,N_13085,N_13745);
and UO_730 (O_730,N_12768,N_12160);
and UO_731 (O_731,N_13362,N_14662);
nand UO_732 (O_732,N_13031,N_12789);
xor UO_733 (O_733,N_14487,N_12933);
nor UO_734 (O_734,N_13612,N_14304);
nor UO_735 (O_735,N_14894,N_14506);
and UO_736 (O_736,N_13880,N_14340);
and UO_737 (O_737,N_13571,N_12542);
and UO_738 (O_738,N_12830,N_13709);
and UO_739 (O_739,N_12166,N_12413);
and UO_740 (O_740,N_12795,N_12157);
and UO_741 (O_741,N_12733,N_13301);
or UO_742 (O_742,N_14074,N_13833);
and UO_743 (O_743,N_13005,N_14456);
nor UO_744 (O_744,N_12610,N_12219);
and UO_745 (O_745,N_12028,N_13550);
or UO_746 (O_746,N_12579,N_14114);
nand UO_747 (O_747,N_14554,N_12690);
nand UO_748 (O_748,N_12240,N_14550);
or UO_749 (O_749,N_13335,N_14509);
nor UO_750 (O_750,N_12859,N_14956);
nand UO_751 (O_751,N_14415,N_13560);
or UO_752 (O_752,N_14584,N_14877);
or UO_753 (O_753,N_13389,N_13106);
or UO_754 (O_754,N_13710,N_14477);
nand UO_755 (O_755,N_14388,N_12200);
nor UO_756 (O_756,N_12387,N_12904);
or UO_757 (O_757,N_12086,N_14860);
nor UO_758 (O_758,N_12945,N_14104);
or UO_759 (O_759,N_13171,N_13502);
and UO_760 (O_760,N_12583,N_14764);
nor UO_761 (O_761,N_13448,N_14393);
nand UO_762 (O_762,N_12465,N_14466);
nand UO_763 (O_763,N_13273,N_14964);
or UO_764 (O_764,N_13010,N_13375);
nor UO_765 (O_765,N_13904,N_12616);
nand UO_766 (O_766,N_12667,N_12340);
or UO_767 (O_767,N_13365,N_13220);
or UO_768 (O_768,N_13499,N_12566);
or UO_769 (O_769,N_12215,N_13168);
nand UO_770 (O_770,N_13820,N_12456);
nor UO_771 (O_771,N_13153,N_12104);
and UO_772 (O_772,N_14874,N_13468);
nor UO_773 (O_773,N_14976,N_14407);
or UO_774 (O_774,N_12058,N_13084);
or UO_775 (O_775,N_14618,N_14364);
nand UO_776 (O_776,N_14857,N_14018);
or UO_777 (O_777,N_13215,N_14290);
or UO_778 (O_778,N_12134,N_13508);
nand UO_779 (O_779,N_12042,N_14021);
nor UO_780 (O_780,N_13479,N_14748);
or UO_781 (O_781,N_12182,N_12243);
and UO_782 (O_782,N_14700,N_13874);
nor UO_783 (O_783,N_12072,N_13649);
and UO_784 (O_784,N_14130,N_13185);
nor UO_785 (O_785,N_13319,N_14184);
nand UO_786 (O_786,N_12728,N_14802);
and UO_787 (O_787,N_12460,N_13212);
or UO_788 (O_788,N_12641,N_12411);
nor UO_789 (O_789,N_12473,N_14223);
nand UO_790 (O_790,N_14044,N_13148);
nand UO_791 (O_791,N_12666,N_14321);
nand UO_792 (O_792,N_14869,N_14612);
nor UO_793 (O_793,N_13540,N_13046);
or UO_794 (O_794,N_14743,N_14895);
or UO_795 (O_795,N_13750,N_13634);
and UO_796 (O_796,N_12590,N_12037);
nand UO_797 (O_797,N_13428,N_14254);
nand UO_798 (O_798,N_12019,N_13871);
and UO_799 (O_799,N_14375,N_14640);
and UO_800 (O_800,N_13628,N_13885);
or UO_801 (O_801,N_12017,N_13826);
nor UO_802 (O_802,N_13521,N_13896);
and UO_803 (O_803,N_12409,N_12685);
nand UO_804 (O_804,N_13258,N_14058);
nor UO_805 (O_805,N_14280,N_12674);
or UO_806 (O_806,N_13366,N_14944);
nor UO_807 (O_807,N_12891,N_12775);
and UO_808 (O_808,N_12982,N_12475);
and UO_809 (O_809,N_13054,N_14189);
and UO_810 (O_810,N_12868,N_14170);
nand UO_811 (O_811,N_12515,N_13933);
and UO_812 (O_812,N_12576,N_13915);
and UO_813 (O_813,N_14274,N_13673);
nand UO_814 (O_814,N_14072,N_12546);
or UO_815 (O_815,N_12061,N_13638);
nor UO_816 (O_816,N_14447,N_13728);
or UO_817 (O_817,N_12040,N_14715);
or UO_818 (O_818,N_13973,N_12824);
and UO_819 (O_819,N_14311,N_12270);
nand UO_820 (O_820,N_14306,N_12883);
nand UO_821 (O_821,N_14836,N_13506);
or UO_822 (O_822,N_12574,N_14644);
nor UO_823 (O_823,N_14588,N_12448);
nor UO_824 (O_824,N_12995,N_13708);
or UO_825 (O_825,N_14168,N_14541);
or UO_826 (O_826,N_14667,N_13420);
and UO_827 (O_827,N_12827,N_13982);
nor UO_828 (O_828,N_13966,N_12695);
or UO_829 (O_829,N_12765,N_14994);
or UO_830 (O_830,N_13925,N_12359);
or UO_831 (O_831,N_13702,N_12097);
nand UO_832 (O_832,N_12298,N_13920);
or UO_833 (O_833,N_14727,N_14746);
nand UO_834 (O_834,N_14699,N_14416);
or UO_835 (O_835,N_14844,N_14492);
and UO_836 (O_836,N_13060,N_12048);
or UO_837 (O_837,N_12747,N_13310);
or UO_838 (O_838,N_12793,N_14726);
and UO_839 (O_839,N_14779,N_13802);
nor UO_840 (O_840,N_14110,N_13291);
or UO_841 (O_841,N_13000,N_12178);
and UO_842 (O_842,N_13178,N_14908);
or UO_843 (O_843,N_14255,N_14396);
or UO_844 (O_844,N_12582,N_12823);
nor UO_845 (O_845,N_14538,N_14227);
nor UO_846 (O_846,N_12654,N_14781);
nand UO_847 (O_847,N_14540,N_13256);
or UO_848 (O_848,N_12144,N_13743);
nor UO_849 (O_849,N_12586,N_13863);
and UO_850 (O_850,N_12129,N_12032);
and UO_851 (O_851,N_13527,N_13851);
or UO_852 (O_852,N_12300,N_13970);
nor UO_853 (O_853,N_13798,N_14824);
nor UO_854 (O_854,N_13255,N_14995);
nand UO_855 (O_855,N_14429,N_12888);
nand UO_856 (O_856,N_14185,N_14659);
and UO_857 (O_857,N_13284,N_14106);
nand UO_858 (O_858,N_13866,N_13793);
nor UO_859 (O_859,N_14474,N_13156);
or UO_860 (O_860,N_14015,N_14671);
nor UO_861 (O_861,N_12511,N_12730);
nor UO_862 (O_862,N_14753,N_12095);
nor UO_863 (O_863,N_13697,N_12819);
nand UO_864 (O_864,N_12866,N_12452);
nor UO_865 (O_865,N_12487,N_14507);
nand UO_866 (O_866,N_12892,N_13867);
and UO_867 (O_867,N_14835,N_13837);
and UO_868 (O_868,N_13391,N_14251);
nor UO_869 (O_869,N_13111,N_14928);
or UO_870 (O_870,N_14890,N_14624);
nor UO_871 (O_871,N_13597,N_12842);
nor UO_872 (O_872,N_13295,N_12952);
nor UO_873 (O_873,N_14804,N_12030);
nor UO_874 (O_874,N_14513,N_13270);
and UO_875 (O_875,N_12960,N_14889);
or UO_876 (O_876,N_12175,N_13203);
nand UO_877 (O_877,N_13327,N_12113);
nand UO_878 (O_878,N_13608,N_12369);
and UO_879 (O_879,N_12870,N_13913);
and UO_880 (O_880,N_13901,N_14172);
nor UO_881 (O_881,N_12917,N_13678);
and UO_882 (O_882,N_13003,N_14469);
nor UO_883 (O_883,N_12014,N_13794);
or UO_884 (O_884,N_13671,N_13194);
and UO_885 (O_885,N_13515,N_13079);
and UO_886 (O_886,N_14762,N_13138);
nor UO_887 (O_887,N_14160,N_14599);
or UO_888 (O_888,N_13744,N_13136);
nor UO_889 (O_889,N_13881,N_13383);
or UO_890 (O_890,N_14040,N_13685);
and UO_891 (O_891,N_14161,N_12807);
nor UO_892 (O_892,N_13528,N_13414);
nand UO_893 (O_893,N_12110,N_14615);
nor UO_894 (O_894,N_13238,N_12084);
or UO_895 (O_895,N_13396,N_13914);
nand UO_896 (O_896,N_14829,N_13378);
and UO_897 (O_897,N_14463,N_14188);
and UO_898 (O_898,N_13100,N_14377);
and UO_899 (O_899,N_13704,N_12090);
nor UO_900 (O_900,N_14461,N_12108);
and UO_901 (O_901,N_12696,N_14433);
or UO_902 (O_902,N_13971,N_12373);
nor UO_903 (O_903,N_13838,N_14646);
nand UO_904 (O_904,N_13856,N_12130);
or UO_905 (O_905,N_12623,N_12822);
and UO_906 (O_906,N_14179,N_14473);
and UO_907 (O_907,N_13983,N_13606);
or UO_908 (O_908,N_14745,N_12426);
and UO_909 (O_909,N_12534,N_12814);
or UO_910 (O_910,N_14390,N_12700);
or UO_911 (O_911,N_13861,N_12643);
nor UO_912 (O_912,N_12679,N_14904);
nor UO_913 (O_913,N_12855,N_13765);
xnor UO_914 (O_914,N_13679,N_12668);
nor UO_915 (O_915,N_14066,N_14927);
nand UO_916 (O_916,N_13855,N_12972);
and UO_917 (O_917,N_13036,N_13781);
nand UO_918 (O_918,N_13072,N_12326);
nand UO_919 (O_919,N_14454,N_13485);
and UO_920 (O_920,N_14602,N_13526);
or UO_921 (O_921,N_13574,N_14445);
and UO_922 (O_922,N_12710,N_12131);
and UO_923 (O_923,N_13858,N_12911);
or UO_924 (O_924,N_14164,N_12489);
nor UO_925 (O_925,N_12401,N_14705);
nand UO_926 (O_926,N_12251,N_12224);
nand UO_927 (O_927,N_12124,N_12287);
or UO_928 (O_928,N_14797,N_12966);
and UO_929 (O_929,N_14061,N_14147);
nor UO_930 (O_930,N_13799,N_14935);
or UO_931 (O_931,N_12268,N_14453);
or UO_932 (O_932,N_13487,N_14658);
nor UO_933 (O_933,N_13443,N_14120);
xor UO_934 (O_934,N_13450,N_13876);
or UO_935 (O_935,N_13427,N_12681);
or UO_936 (O_936,N_14932,N_12106);
nor UO_937 (O_937,N_12493,N_14868);
and UO_938 (O_938,N_12652,N_13969);
nand UO_939 (O_939,N_13747,N_13535);
nand UO_940 (O_940,N_12806,N_12671);
and UO_941 (O_941,N_13231,N_12196);
and UO_942 (O_942,N_12433,N_13584);
nor UO_943 (O_943,N_12595,N_12439);
and UO_944 (O_944,N_12067,N_12185);
and UO_945 (O_945,N_13438,N_13419);
nand UO_946 (O_946,N_13151,N_14100);
nor UO_947 (O_947,N_14291,N_13229);
and UO_948 (O_948,N_13723,N_12228);
or UO_949 (O_949,N_12339,N_12449);
and UO_950 (O_950,N_12637,N_14276);
nor UO_951 (O_951,N_12246,N_12687);
nand UO_952 (O_952,N_14298,N_14790);
or UO_953 (O_953,N_13687,N_12554);
nand UO_954 (O_954,N_12738,N_14346);
nor UO_955 (O_955,N_12540,N_13556);
and UO_956 (O_956,N_13349,N_13773);
and UO_957 (O_957,N_13500,N_14438);
or UO_958 (O_958,N_13233,N_12085);
or UO_959 (O_959,N_12557,N_13477);
or UO_960 (O_960,N_12757,N_13379);
and UO_961 (O_961,N_14275,N_14912);
or UO_962 (O_962,N_12342,N_13018);
or UO_963 (O_963,N_12895,N_14997);
and UO_964 (O_964,N_12220,N_13037);
nor UO_965 (O_965,N_13590,N_13370);
nor UO_966 (O_966,N_14817,N_14234);
and UO_967 (O_967,N_14693,N_13024);
nor UO_968 (O_968,N_12265,N_14863);
or UO_969 (O_969,N_12896,N_13730);
and UO_970 (O_970,N_13439,N_14587);
nor UO_971 (O_971,N_12076,N_14529);
or UO_972 (O_972,N_12469,N_14674);
or UO_973 (O_973,N_12584,N_12151);
and UO_974 (O_974,N_13063,N_13611);
and UO_975 (O_975,N_12902,N_12441);
nor UO_976 (O_976,N_13530,N_14776);
and UO_977 (O_977,N_14287,N_12405);
or UO_978 (O_978,N_13929,N_14020);
and UO_979 (O_979,N_13895,N_14918);
or UO_980 (O_980,N_12609,N_13691);
and UO_981 (O_981,N_14153,N_14394);
or UO_982 (O_982,N_12309,N_12416);
or UO_983 (O_983,N_12050,N_12498);
and UO_984 (O_984,N_14673,N_13572);
nand UO_985 (O_985,N_12060,N_14268);
and UO_986 (O_986,N_14421,N_13618);
or UO_987 (O_987,N_13308,N_12915);
nor UO_988 (O_988,N_12143,N_12628);
nor UO_989 (O_989,N_12382,N_12751);
nand UO_990 (O_990,N_13853,N_12916);
and UO_991 (O_991,N_14972,N_14893);
nor UO_992 (O_992,N_12813,N_14794);
and UO_993 (O_993,N_12378,N_12485);
and UO_994 (O_994,N_14939,N_13713);
nand UO_995 (O_995,N_13624,N_14795);
nand UO_996 (O_996,N_12837,N_12139);
or UO_997 (O_997,N_14756,N_12353);
and UO_998 (O_998,N_13778,N_14589);
or UO_999 (O_999,N_12527,N_13610);
or UO_1000 (O_1000,N_14782,N_13942);
and UO_1001 (O_1001,N_14533,N_14329);
or UO_1002 (O_1002,N_12317,N_12691);
and UO_1003 (O_1003,N_14771,N_13818);
and UO_1004 (O_1004,N_13846,N_14996);
and UO_1005 (O_1005,N_12303,N_13949);
or UO_1006 (O_1006,N_12446,N_13698);
nand UO_1007 (O_1007,N_13113,N_12720);
nand UO_1008 (O_1008,N_14112,N_14210);
nor UO_1009 (O_1009,N_14439,N_13135);
nor UO_1010 (O_1010,N_14523,N_12337);
and UO_1011 (O_1011,N_14320,N_12447);
nor UO_1012 (O_1012,N_13946,N_13155);
and UO_1013 (O_1013,N_13603,N_12444);
nand UO_1014 (O_1014,N_13035,N_12990);
and UO_1015 (O_1015,N_13141,N_12330);
or UO_1016 (O_1016,N_13126,N_14132);
nand UO_1017 (O_1017,N_14557,N_13680);
nor UO_1018 (O_1018,N_13924,N_14315);
nand UO_1019 (O_1019,N_13023,N_14798);
and UO_1020 (O_1020,N_14544,N_12683);
or UO_1021 (O_1021,N_13159,N_14528);
and UO_1022 (O_1022,N_12862,N_13642);
nand UO_1023 (O_1023,N_12038,N_14725);
and UO_1024 (O_1024,N_13025,N_14174);
nor UO_1025 (O_1025,N_13149,N_13986);
nor UO_1026 (O_1026,N_12354,N_12109);
nand UO_1027 (O_1027,N_13965,N_14579);
nor UO_1028 (O_1028,N_13200,N_14712);
and UO_1029 (O_1029,N_13694,N_13842);
and UO_1030 (O_1030,N_14448,N_13677);
nor UO_1031 (O_1031,N_12140,N_13221);
nand UO_1032 (O_1032,N_14468,N_13756);
nor UO_1033 (O_1033,N_12970,N_14631);
nand UO_1034 (O_1034,N_14093,N_13565);
nor UO_1035 (O_1035,N_14266,N_13397);
nor UO_1036 (O_1036,N_12978,N_14392);
and UO_1037 (O_1037,N_13411,N_14569);
nand UO_1038 (O_1038,N_14943,N_12083);
and UO_1039 (O_1039,N_14657,N_14929);
or UO_1040 (O_1040,N_13341,N_12856);
nand UO_1041 (O_1041,N_12286,N_13832);
nand UO_1042 (O_1042,N_13578,N_14446);
nor UO_1043 (O_1043,N_14195,N_12275);
nand UO_1044 (O_1044,N_13449,N_12395);
and UO_1045 (O_1045,N_13122,N_13355);
and UO_1046 (O_1046,N_12005,N_12919);
nand UO_1047 (O_1047,N_12454,N_14954);
or UO_1048 (O_1048,N_13652,N_12421);
nand UO_1049 (O_1049,N_14208,N_14230);
or UO_1050 (O_1050,N_14719,N_14906);
or UO_1051 (O_1051,N_14271,N_13727);
or UO_1052 (O_1052,N_12620,N_14936);
nand UO_1053 (O_1053,N_13943,N_12291);
xnor UO_1054 (O_1054,N_14633,N_14810);
and UO_1055 (O_1055,N_14109,N_14878);
or UO_1056 (O_1056,N_12338,N_13813);
or UO_1057 (O_1057,N_14959,N_13211);
or UO_1058 (O_1058,N_12098,N_13985);
or UO_1059 (O_1059,N_12630,N_12847);
or UO_1060 (O_1060,N_13492,N_12273);
and UO_1061 (O_1061,N_13980,N_13317);
or UO_1062 (O_1062,N_12276,N_13937);
or UO_1063 (O_1063,N_12563,N_13564);
or UO_1064 (O_1064,N_12816,N_12597);
nand UO_1065 (O_1065,N_14297,N_14852);
and UO_1066 (O_1066,N_14742,N_14413);
and UO_1067 (O_1067,N_12692,N_12331);
nand UO_1068 (O_1068,N_14419,N_14402);
nor UO_1069 (O_1069,N_14552,N_14198);
nor UO_1070 (O_1070,N_13640,N_13269);
or UO_1071 (O_1071,N_13223,N_13777);
or UO_1072 (O_1072,N_13524,N_14534);
nand UO_1073 (O_1073,N_14708,N_12519);
and UO_1074 (O_1074,N_14076,N_12184);
nor UO_1075 (O_1075,N_13065,N_12935);
nor UO_1076 (O_1076,N_12150,N_14775);
nor UO_1077 (O_1077,N_12857,N_12538);
nand UO_1078 (O_1078,N_14366,N_13340);
or UO_1079 (O_1079,N_14286,N_12245);
nand UO_1080 (O_1080,N_13189,N_12882);
nand UO_1081 (O_1081,N_13735,N_13302);
nor UO_1082 (O_1082,N_14953,N_14728);
nor UO_1083 (O_1083,N_14398,N_13180);
or UO_1084 (O_1084,N_14470,N_13406);
nand UO_1085 (O_1085,N_13595,N_14621);
or UO_1086 (O_1086,N_13804,N_14118);
nor UO_1087 (O_1087,N_12663,N_12358);
and UO_1088 (O_1088,N_14826,N_12713);
nor UO_1089 (O_1089,N_12082,N_13403);
nor UO_1090 (O_1090,N_14442,N_14206);
nand UO_1091 (O_1091,N_12249,N_13721);
and UO_1092 (O_1092,N_13972,N_14397);
nand UO_1093 (O_1093,N_13533,N_12998);
nor UO_1094 (O_1094,N_12128,N_13674);
or UO_1095 (O_1095,N_12003,N_14949);
and UO_1096 (O_1096,N_14575,N_12953);
and UO_1097 (O_1097,N_14777,N_14697);
and UO_1098 (O_1098,N_14428,N_14049);
and UO_1099 (O_1099,N_13457,N_14630);
or UO_1100 (O_1100,N_12333,N_12188);
nor UO_1101 (O_1101,N_13532,N_12938);
nor UO_1102 (O_1102,N_14143,N_12835);
and UO_1103 (O_1103,N_12357,N_14593);
or UO_1104 (O_1104,N_13294,N_12996);
nand UO_1105 (O_1105,N_14231,N_12961);
nand UO_1106 (O_1106,N_12347,N_12255);
or UO_1107 (O_1107,N_13288,N_12403);
or UO_1108 (O_1108,N_13337,N_14012);
nand UO_1109 (O_1109,N_12181,N_14193);
nor UO_1110 (O_1110,N_12295,N_12841);
and UO_1111 (O_1111,N_13045,N_14125);
nand UO_1112 (O_1112,N_13090,N_12636);
or UO_1113 (O_1113,N_13921,N_14349);
and UO_1114 (O_1114,N_12532,N_14695);
nand UO_1115 (O_1115,N_13683,N_14412);
nor UO_1116 (O_1116,N_12074,N_13586);
nor UO_1117 (O_1117,N_13137,N_14083);
and UO_1118 (O_1118,N_13543,N_13016);
and UO_1119 (O_1119,N_14859,N_13444);
or UO_1120 (O_1120,N_12051,N_13664);
nor UO_1121 (O_1121,N_12648,N_12712);
and UO_1122 (O_1122,N_13075,N_14410);
nand UO_1123 (O_1123,N_14218,N_12290);
nand UO_1124 (O_1124,N_14369,N_12605);
nand UO_1125 (O_1125,N_12716,N_14116);
nand UO_1126 (O_1126,N_12780,N_14926);
and UO_1127 (O_1127,N_13731,N_14947);
and UO_1128 (O_1128,N_14358,N_13196);
and UO_1129 (O_1129,N_14503,N_13907);
or UO_1130 (O_1130,N_13405,N_12703);
nand UO_1131 (O_1131,N_13912,N_14546);
and UO_1132 (O_1132,N_14505,N_12207);
or UO_1133 (O_1133,N_12183,N_13623);
and UO_1134 (O_1134,N_13109,N_12486);
or UO_1135 (O_1135,N_14235,N_13013);
nand UO_1136 (O_1136,N_14205,N_12367);
or UO_1137 (O_1137,N_12541,N_14504);
or UO_1138 (O_1138,N_14952,N_14980);
nor UO_1139 (O_1139,N_12568,N_12053);
and UO_1140 (O_1140,N_14880,N_13182);
nor UO_1141 (O_1141,N_12976,N_13504);
or UO_1142 (O_1142,N_13513,N_13491);
nor UO_1143 (O_1143,N_12873,N_13591);
nand UO_1144 (O_1144,N_13699,N_13746);
and UO_1145 (O_1145,N_12941,N_12521);
nor UO_1146 (O_1146,N_12383,N_14827);
nor UO_1147 (O_1147,N_13823,N_14080);
xnor UO_1148 (O_1148,N_13806,N_13073);
nor UO_1149 (O_1149,N_12221,N_12779);
or UO_1150 (O_1150,N_14484,N_14720);
or UO_1151 (O_1151,N_14731,N_12327);
or UO_1152 (O_1152,N_13123,N_13910);
and UO_1153 (O_1153,N_12396,N_13816);
or UO_1154 (O_1154,N_13198,N_14524);
nand UO_1155 (O_1155,N_13951,N_12924);
nor UO_1156 (O_1156,N_12860,N_13230);
and UO_1157 (O_1157,N_13956,N_14097);
and UO_1158 (O_1158,N_14313,N_12589);
nor UO_1159 (O_1159,N_14257,N_12908);
and UO_1160 (O_1160,N_12078,N_13545);
nand UO_1161 (O_1161,N_13132,N_13412);
nor UO_1162 (O_1162,N_12041,N_12216);
nand UO_1163 (O_1163,N_12558,N_14092);
nor UO_1164 (O_1164,N_12389,N_13228);
or UO_1165 (O_1165,N_14694,N_13812);
or UO_1166 (O_1166,N_13994,N_12015);
or UO_1167 (O_1167,N_14886,N_12974);
or UO_1168 (O_1168,N_12173,N_12484);
or UO_1169 (O_1169,N_12580,N_12368);
and UO_1170 (O_1170,N_12235,N_12905);
nor UO_1171 (O_1171,N_12135,N_14345);
and UO_1172 (O_1172,N_12047,N_12959);
and UO_1173 (O_1173,N_12936,N_12324);
and UO_1174 (O_1174,N_13087,N_14819);
nor UO_1175 (O_1175,N_12784,N_12271);
nand UO_1176 (O_1176,N_12923,N_13766);
or UO_1177 (O_1177,N_14224,N_13179);
or UO_1178 (O_1178,N_13548,N_14293);
nor UO_1179 (O_1179,N_13019,N_14406);
and UO_1180 (O_1180,N_14336,N_14002);
nand UO_1181 (O_1181,N_14661,N_13754);
nor UO_1182 (O_1182,N_13824,N_12619);
or UO_1183 (O_1183,N_14178,N_13086);
nand UO_1184 (O_1184,N_12450,N_12087);
nor UO_1185 (O_1185,N_14750,N_13567);
nor UO_1186 (O_1186,N_12066,N_14650);
and UO_1187 (O_1187,N_12744,N_13967);
nand UO_1188 (O_1188,N_14382,N_13129);
nand UO_1189 (O_1189,N_13293,N_14834);
or UO_1190 (O_1190,N_12190,N_14107);
nor UO_1191 (O_1191,N_14751,N_14736);
xnor UO_1192 (O_1192,N_13774,N_13121);
nor UO_1193 (O_1193,N_14046,N_13404);
nand UO_1194 (O_1194,N_13979,N_13425);
or UO_1195 (O_1195,N_13440,N_12836);
or UO_1196 (O_1196,N_13183,N_13600);
and UO_1197 (O_1197,N_14535,N_14755);
or UO_1198 (O_1198,N_13632,N_12259);
nor UO_1199 (O_1199,N_12825,N_14670);
or UO_1200 (O_1200,N_13286,N_14399);
nand UO_1201 (O_1201,N_12719,N_13537);
or UO_1202 (O_1202,N_13845,N_13964);
nor UO_1203 (O_1203,N_12199,N_12307);
or UO_1204 (O_1204,N_13076,N_14094);
or UO_1205 (O_1205,N_12567,N_12010);
or UO_1206 (O_1206,N_13434,N_14855);
nor UO_1207 (O_1207,N_12670,N_12539);
nand UO_1208 (O_1208,N_12492,N_12503);
nor UO_1209 (O_1209,N_12296,N_13662);
nor UO_1210 (O_1210,N_14786,N_12052);
or UO_1211 (O_1211,N_13433,N_13250);
or UO_1212 (O_1212,N_12189,N_12505);
nand UO_1213 (O_1213,N_13809,N_13829);
and UO_1214 (O_1214,N_14479,N_12677);
nand UO_1215 (O_1215,N_12559,N_12310);
or UO_1216 (O_1216,N_12236,N_13222);
nor UO_1217 (O_1217,N_13958,N_12615);
nor UO_1218 (O_1218,N_14212,N_13186);
or UO_1219 (O_1219,N_12501,N_14354);
or UO_1220 (O_1220,N_14250,N_14634);
nand UO_1221 (O_1221,N_12334,N_13498);
or UO_1222 (O_1222,N_13251,N_14476);
and UO_1223 (O_1223,N_13734,N_14294);
nor UO_1224 (O_1224,N_14152,N_13553);
nand UO_1225 (O_1225,N_13722,N_12156);
nand UO_1226 (O_1226,N_13635,N_13356);
nand UO_1227 (O_1227,N_12197,N_13377);
nand UO_1228 (O_1228,N_13067,N_13030);
nor UO_1229 (O_1229,N_13287,N_13665);
or UO_1230 (O_1230,N_14828,N_14789);
or UO_1231 (O_1231,N_13473,N_13166);
nor UO_1232 (O_1232,N_14594,N_12434);
nor UO_1233 (O_1233,N_12193,N_12930);
nor UO_1234 (O_1234,N_12499,N_14628);
or UO_1235 (O_1235,N_12621,N_12055);
nand UO_1236 (O_1236,N_14341,N_14395);
nand UO_1237 (O_1237,N_12231,N_12018);
nor UO_1238 (O_1238,N_13026,N_14718);
nand UO_1239 (O_1239,N_14128,N_12745);
or UO_1240 (O_1240,N_13531,N_13645);
nor UO_1241 (O_1241,N_12500,N_12721);
or UO_1242 (O_1242,N_14808,N_12940);
nand UO_1243 (O_1243,N_14948,N_13165);
nor UO_1244 (O_1244,N_12918,N_13968);
nor UO_1245 (O_1245,N_14566,N_14055);
nor UO_1246 (O_1246,N_12760,N_12979);
and UO_1247 (O_1247,N_14642,N_14814);
or UO_1248 (O_1248,N_13246,N_14069);
and UO_1249 (O_1249,N_13154,N_13394);
nand UO_1250 (O_1250,N_14663,N_13028);
nor UO_1251 (O_1251,N_14420,N_12992);
and UO_1252 (O_1252,N_12776,N_12379);
nor UO_1253 (O_1253,N_13890,N_14800);
and UO_1254 (O_1254,N_12356,N_13577);
and UO_1255 (O_1255,N_12781,N_14521);
or UO_1256 (O_1256,N_12404,N_14084);
and UO_1257 (O_1257,N_12274,N_13782);
and UO_1258 (O_1258,N_14574,N_13923);
or UO_1259 (O_1259,N_13465,N_13367);
and UO_1260 (O_1260,N_12955,N_14408);
nand UO_1261 (O_1261,N_13607,N_12399);
nand UO_1262 (O_1262,N_14365,N_14352);
nor UO_1263 (O_1263,N_12811,N_13006);
or UO_1264 (O_1264,N_12516,N_13202);
nand UO_1265 (O_1265,N_14909,N_12377);
and UO_1266 (O_1266,N_12675,N_12075);
and UO_1267 (O_1267,N_13738,N_13934);
and UO_1268 (O_1268,N_13817,N_12355);
and UO_1269 (O_1269,N_13639,N_14192);
nand UO_1270 (O_1270,N_14520,N_13464);
nand UO_1271 (O_1271,N_13309,N_14580);
nand UO_1272 (O_1272,N_14920,N_13057);
and UO_1273 (O_1273,N_13408,N_14660);
nor UO_1274 (O_1274,N_13637,N_13941);
and UO_1275 (O_1275,N_14683,N_13441);
nand UO_1276 (O_1276,N_13034,N_14962);
nand UO_1277 (O_1277,N_14269,N_13633);
and UO_1278 (O_1278,N_14324,N_12627);
nand UO_1279 (O_1279,N_14182,N_12601);
nor UO_1280 (O_1280,N_14570,N_14645);
or UO_1281 (O_1281,N_14146,N_12375);
nand UO_1282 (O_1282,N_12889,N_14158);
nand UO_1283 (O_1283,N_13128,N_14272);
and UO_1284 (O_1284,N_12262,N_13497);
and UO_1285 (O_1285,N_13482,N_13354);
nor UO_1286 (O_1286,N_13868,N_13939);
and UO_1287 (O_1287,N_14522,N_14252);
nand UO_1288 (O_1288,N_12089,N_12280);
nand UO_1289 (O_1289,N_12321,N_14444);
nor UO_1290 (O_1290,N_13598,N_14862);
or UO_1291 (O_1291,N_12318,N_14443);
and UO_1292 (O_1292,N_14998,N_13217);
nor UO_1293 (O_1293,N_13908,N_14915);
nor UO_1294 (O_1294,N_12102,N_13249);
nand UO_1295 (O_1295,N_14586,N_13039);
nor UO_1296 (O_1296,N_13688,N_13040);
and UO_1297 (O_1297,N_13357,N_13263);
nand UO_1298 (O_1298,N_14488,N_14767);
or UO_1299 (O_1299,N_14023,N_13952);
nand UO_1300 (O_1300,N_14258,N_14403);
nand UO_1301 (O_1301,N_14363,N_14934);
and UO_1302 (O_1302,N_13014,N_13056);
nand UO_1303 (O_1303,N_14647,N_13336);
or UO_1304 (O_1304,N_14197,N_14517);
and UO_1305 (O_1305,N_12887,N_13681);
or UO_1306 (O_1306,N_12142,N_14806);
nor UO_1307 (O_1307,N_12234,N_14183);
or UO_1308 (O_1308,N_13839,N_12352);
or UO_1309 (O_1309,N_12848,N_12707);
and UO_1310 (O_1310,N_13814,N_14067);
nor UO_1311 (O_1311,N_14608,N_12647);
or UO_1312 (O_1312,N_14875,N_12769);
nor UO_1313 (O_1313,N_12914,N_14793);
nand UO_1314 (O_1314,N_13199,N_14763);
and UO_1315 (O_1315,N_12374,N_13882);
nand UO_1316 (O_1316,N_14335,N_12122);
nor UO_1317 (O_1317,N_14075,N_14495);
nand UO_1318 (O_1318,N_14837,N_12443);
and UO_1319 (O_1319,N_14632,N_12248);
or UO_1320 (O_1320,N_12092,N_13568);
nor UO_1321 (O_1321,N_13442,N_12279);
nand UO_1322 (O_1322,N_12838,N_13459);
or UO_1323 (O_1323,N_14951,N_12684);
or UO_1324 (O_1324,N_13152,N_14957);
and UO_1325 (O_1325,N_12137,N_12214);
and UO_1326 (O_1326,N_14519,N_14400);
or UO_1327 (O_1327,N_12045,N_12000);
nand UO_1328 (O_1328,N_12417,N_13472);
nor UO_1329 (O_1329,N_14101,N_12782);
nand UO_1330 (O_1330,N_12680,N_13012);
xnor UO_1331 (O_1331,N_12257,N_14262);
nand UO_1332 (O_1332,N_14131,N_12704);
nand UO_1333 (O_1333,N_12815,N_13981);
nand UO_1334 (O_1334,N_13467,N_13120);
nand UO_1335 (O_1335,N_14739,N_13788);
or UO_1336 (O_1336,N_12606,N_14163);
or UO_1337 (O_1337,N_12132,N_13278);
nand UO_1338 (O_1338,N_14434,N_12622);
or UO_1339 (O_1339,N_12453,N_12364);
nor UO_1340 (O_1340,N_12877,N_13298);
or UO_1341 (O_1341,N_13575,N_12925);
and UO_1342 (O_1342,N_13666,N_12629);
nor UO_1343 (O_1343,N_12402,N_14734);
or UO_1344 (O_1344,N_12725,N_12773);
or UO_1345 (O_1345,N_12025,N_14769);
or UO_1346 (O_1346,N_12922,N_12332);
nand UO_1347 (O_1347,N_13563,N_14236);
and UO_1348 (O_1348,N_12408,N_12059);
or UO_1349 (O_1349,N_14968,N_14190);
and UO_1350 (O_1350,N_14656,N_13733);
nand UO_1351 (O_1351,N_14460,N_14830);
nor UO_1352 (O_1352,N_13409,N_14652);
and UO_1353 (O_1353,N_14035,N_13879);
nand UO_1354 (O_1354,N_12898,N_14339);
or UO_1355 (O_1355,N_13748,N_14289);
nor UO_1356 (O_1356,N_12256,N_13248);
and UO_1357 (O_1357,N_14922,N_14144);
nor UO_1358 (O_1358,N_14299,N_14682);
or UO_1359 (O_1359,N_13758,N_14933);
nand UO_1360 (O_1360,N_12598,N_12577);
and UO_1361 (O_1361,N_14553,N_13494);
and UO_1362 (O_1362,N_14499,N_14653);
and UO_1363 (O_1363,N_12437,N_13505);
or UO_1364 (O_1364,N_14971,N_12509);
or UO_1365 (O_1365,N_12646,N_13792);
and UO_1366 (O_1366,N_14688,N_13622);
or UO_1367 (O_1367,N_14916,N_14404);
nor UO_1368 (O_1368,N_14681,N_13701);
and UO_1369 (O_1369,N_12573,N_14332);
and UO_1370 (O_1370,N_13789,N_12658);
or UO_1371 (O_1371,N_12968,N_12315);
nor UO_1372 (O_1372,N_12208,N_13900);
and UO_1373 (O_1373,N_12261,N_12852);
or UO_1374 (O_1374,N_12250,N_12928);
nand UO_1375 (O_1375,N_12020,N_12942);
and UO_1376 (O_1376,N_12934,N_12127);
or UO_1377 (O_1377,N_14314,N_14028);
or UO_1378 (O_1378,N_13455,N_14279);
and UO_1379 (O_1379,N_13596,N_12759);
nor UO_1380 (O_1380,N_13417,N_12136);
nand UO_1381 (O_1381,N_12553,N_12980);
or UO_1382 (O_1382,N_14899,N_12414);
and UO_1383 (O_1383,N_14596,N_14930);
or UO_1384 (O_1384,N_14950,N_12429);
nand UO_1385 (O_1385,N_13323,N_12858);
or UO_1386 (O_1386,N_13658,N_13726);
and UO_1387 (O_1387,N_12699,N_14086);
nand UO_1388 (O_1388,N_13534,N_12165);
nand UO_1389 (O_1389,N_14296,N_13695);
nor UO_1390 (O_1390,N_14242,N_14471);
nor UO_1391 (O_1391,N_13413,N_14117);
or UO_1392 (O_1392,N_12947,N_14127);
and UO_1393 (O_1393,N_12079,N_12599);
nand UO_1394 (O_1394,N_14627,N_12138);
or UO_1395 (O_1395,N_12743,N_12065);
nand UO_1396 (O_1396,N_14325,N_12026);
nor UO_1397 (O_1397,N_13474,N_12227);
or UO_1398 (O_1398,N_12495,N_14714);
and UO_1399 (O_1399,N_14034,N_12119);
and UO_1400 (O_1400,N_14219,N_12177);
or UO_1401 (O_1401,N_12951,N_12849);
nor UO_1402 (O_1402,N_12294,N_13670);
and UO_1403 (O_1403,N_14576,N_13583);
nand UO_1404 (O_1404,N_12518,N_12420);
xnor UO_1405 (O_1405,N_13997,N_12180);
nand UO_1406 (O_1406,N_13264,N_13770);
nand UO_1407 (O_1407,N_13892,N_13279);
nand UO_1408 (O_1408,N_14655,N_12336);
and UO_1409 (O_1409,N_14214,N_13351);
and UO_1410 (O_1410,N_12385,N_12313);
or UO_1411 (O_1411,N_12210,N_14536);
nand UO_1412 (O_1412,N_14138,N_13333);
nor UO_1413 (O_1413,N_13283,N_13422);
nor UO_1414 (O_1414,N_13819,N_12419);
nor UO_1415 (O_1415,N_14221,N_12635);
or UO_1416 (O_1416,N_13764,N_13488);
nor UO_1417 (O_1417,N_12325,N_13902);
or UO_1418 (O_1418,N_14542,N_14233);
or UO_1419 (O_1419,N_12556,N_13029);
nand UO_1420 (O_1420,N_14788,N_13078);
nor UO_1421 (O_1421,N_13529,N_13115);
nand UO_1422 (O_1422,N_14825,N_12311);
nor UO_1423 (O_1423,N_14318,N_14348);
nor UO_1424 (O_1424,N_12766,N_12007);
and UO_1425 (O_1425,N_12263,N_14312);
and UO_1426 (O_1426,N_14359,N_14368);
nand UO_1427 (O_1427,N_12543,N_14501);
nor UO_1428 (O_1428,N_12174,N_12366);
and UO_1429 (O_1429,N_13785,N_13253);
or UO_1430 (O_1430,N_13587,N_14070);
and UO_1431 (O_1431,N_13576,N_13193);
or UO_1432 (O_1432,N_13239,N_12880);
or UO_1433 (O_1433,N_13116,N_14338);
and UO_1434 (O_1434,N_13398,N_14062);
nor UO_1435 (O_1435,N_14180,N_12410);
nand UO_1436 (O_1436,N_13715,N_12785);
and UO_1437 (O_1437,N_14085,N_12283);
and UO_1438 (O_1438,N_13539,N_13252);
nand UO_1439 (O_1439,N_13235,N_13810);
nand UO_1440 (O_1440,N_12123,N_13143);
and UO_1441 (O_1441,N_13170,N_12578);
nor UO_1442 (O_1442,N_13887,N_12944);
nor UO_1443 (O_1443,N_12987,N_14007);
and UO_1444 (O_1444,N_14805,N_12022);
nor UO_1445 (O_1445,N_14480,N_12593);
nor UO_1446 (O_1446,N_14441,N_14141);
nor UO_1447 (O_1447,N_12600,N_12805);
nor UO_1448 (O_1448,N_14263,N_12522);
and UO_1449 (O_1449,N_13955,N_13865);
and UO_1450 (O_1450,N_14865,N_14431);
and UO_1451 (O_1451,N_14603,N_13959);
and UO_1452 (O_1452,N_12202,N_12767);
or UO_1453 (O_1453,N_12455,N_14565);
nor UO_1454 (O_1454,N_14362,N_13373);
and UO_1455 (O_1455,N_12114,N_13480);
nand UO_1456 (O_1456,N_12734,N_12524);
and UO_1457 (O_1457,N_14604,N_14491);
or UO_1458 (O_1458,N_12153,N_14558);
and UO_1459 (O_1459,N_14691,N_12812);
or UO_1460 (O_1460,N_12770,N_13352);
nor UO_1461 (O_1461,N_14351,N_14485);
nand UO_1462 (O_1462,N_14237,N_14159);
or UO_1463 (O_1463,N_13145,N_13884);
nand UO_1464 (O_1464,N_13345,N_14041);
and UO_1465 (O_1465,N_12205,N_13458);
and UO_1466 (O_1466,N_13630,N_13020);
nand UO_1467 (O_1467,N_14199,N_12688);
nand UO_1468 (O_1468,N_14946,N_12771);
or UO_1469 (O_1469,N_12850,N_14483);
nor UO_1470 (O_1470,N_13932,N_14680);
nand UO_1471 (O_1471,N_12282,N_12312);
nor UO_1472 (O_1472,N_12575,N_14079);
nand UO_1473 (O_1473,N_12661,N_13552);
and UO_1474 (O_1474,N_14784,N_12080);
nand UO_1475 (O_1475,N_14383,N_12831);
nand UO_1476 (O_1476,N_12906,N_13841);
nand UO_1477 (O_1477,N_14472,N_12604);
nor UO_1478 (O_1478,N_12115,N_13579);
or UO_1479 (O_1479,N_13903,N_12802);
nor UO_1480 (O_1480,N_13891,N_14027);
and UO_1481 (O_1481,N_14539,N_12985);
nor UO_1482 (O_1482,N_14905,N_14625);
nand UO_1483 (O_1483,N_13322,N_14707);
xor UO_1484 (O_1484,N_14796,N_14150);
and UO_1485 (O_1485,N_12125,N_13382);
nand UO_1486 (O_1486,N_12552,N_14261);
and UO_1487 (O_1487,N_14917,N_12062);
nor UO_1488 (O_1488,N_14556,N_12494);
nand UO_1489 (O_1489,N_12094,N_12549);
nor UO_1490 (O_1490,N_12512,N_14323);
and UO_1491 (O_1491,N_13875,N_13609);
and UO_1492 (O_1492,N_14126,N_13780);
nor UO_1493 (O_1493,N_14687,N_13790);
nand UO_1494 (O_1494,N_12023,N_12828);
nand UO_1495 (O_1495,N_12929,N_12392);
nand UO_1496 (O_1496,N_12792,N_12754);
nor UO_1497 (O_1497,N_14675,N_14145);
nor UO_1498 (O_1498,N_14156,N_14842);
nor UO_1499 (O_1499,N_14422,N_13261);
and UO_1500 (O_1500,N_13149,N_12071);
and UO_1501 (O_1501,N_14546,N_13076);
nand UO_1502 (O_1502,N_13191,N_13491);
and UO_1503 (O_1503,N_13509,N_13928);
or UO_1504 (O_1504,N_14275,N_12846);
nand UO_1505 (O_1505,N_14879,N_12155);
nor UO_1506 (O_1506,N_14925,N_12465);
nor UO_1507 (O_1507,N_14976,N_14479);
and UO_1508 (O_1508,N_13232,N_14833);
and UO_1509 (O_1509,N_13216,N_12298);
or UO_1510 (O_1510,N_13530,N_14481);
or UO_1511 (O_1511,N_13889,N_13007);
nor UO_1512 (O_1512,N_14183,N_13217);
and UO_1513 (O_1513,N_14789,N_14817);
or UO_1514 (O_1514,N_13030,N_13805);
nand UO_1515 (O_1515,N_12679,N_14508);
and UO_1516 (O_1516,N_14021,N_12559);
and UO_1517 (O_1517,N_13650,N_14263);
nor UO_1518 (O_1518,N_12450,N_13736);
or UO_1519 (O_1519,N_13260,N_13034);
or UO_1520 (O_1520,N_14223,N_13595);
nand UO_1521 (O_1521,N_12836,N_12317);
and UO_1522 (O_1522,N_14695,N_12070);
or UO_1523 (O_1523,N_13235,N_13988);
and UO_1524 (O_1524,N_12285,N_13416);
and UO_1525 (O_1525,N_12168,N_14496);
or UO_1526 (O_1526,N_14092,N_13423);
and UO_1527 (O_1527,N_13109,N_13286);
and UO_1528 (O_1528,N_14556,N_13095);
nand UO_1529 (O_1529,N_13280,N_12904);
and UO_1530 (O_1530,N_13157,N_13929);
or UO_1531 (O_1531,N_12435,N_13139);
nor UO_1532 (O_1532,N_13947,N_13551);
xnor UO_1533 (O_1533,N_14823,N_12681);
nor UO_1534 (O_1534,N_13107,N_14067);
nor UO_1535 (O_1535,N_14718,N_14002);
and UO_1536 (O_1536,N_14189,N_12079);
nand UO_1537 (O_1537,N_12952,N_14732);
nor UO_1538 (O_1538,N_13792,N_14379);
nor UO_1539 (O_1539,N_12216,N_12153);
and UO_1540 (O_1540,N_14635,N_12018);
nor UO_1541 (O_1541,N_12066,N_13155);
nand UO_1542 (O_1542,N_12449,N_12065);
nand UO_1543 (O_1543,N_14507,N_13861);
or UO_1544 (O_1544,N_14312,N_14804);
or UO_1545 (O_1545,N_14248,N_14752);
or UO_1546 (O_1546,N_12756,N_12940);
or UO_1547 (O_1547,N_12348,N_14984);
nor UO_1548 (O_1548,N_14030,N_14588);
or UO_1549 (O_1549,N_13420,N_12728);
and UO_1550 (O_1550,N_12795,N_14505);
nor UO_1551 (O_1551,N_13687,N_14563);
and UO_1552 (O_1552,N_13326,N_14170);
or UO_1553 (O_1553,N_14871,N_14959);
nand UO_1554 (O_1554,N_14462,N_14750);
nand UO_1555 (O_1555,N_12143,N_14927);
and UO_1556 (O_1556,N_13465,N_12682);
or UO_1557 (O_1557,N_14067,N_13349);
nor UO_1558 (O_1558,N_14723,N_13042);
or UO_1559 (O_1559,N_14051,N_13788);
and UO_1560 (O_1560,N_12968,N_14979);
xor UO_1561 (O_1561,N_12126,N_12617);
and UO_1562 (O_1562,N_14961,N_14219);
xor UO_1563 (O_1563,N_14251,N_14359);
nor UO_1564 (O_1564,N_14638,N_13800);
nand UO_1565 (O_1565,N_14530,N_13187);
nand UO_1566 (O_1566,N_14259,N_12459);
nand UO_1567 (O_1567,N_12567,N_13358);
or UO_1568 (O_1568,N_13651,N_12259);
and UO_1569 (O_1569,N_13474,N_13880);
or UO_1570 (O_1570,N_12820,N_12361);
or UO_1571 (O_1571,N_13950,N_13601);
nand UO_1572 (O_1572,N_14650,N_13137);
and UO_1573 (O_1573,N_12407,N_12222);
nor UO_1574 (O_1574,N_13448,N_14008);
nand UO_1575 (O_1575,N_12138,N_12960);
or UO_1576 (O_1576,N_14361,N_12479);
nor UO_1577 (O_1577,N_14278,N_12730);
and UO_1578 (O_1578,N_14385,N_13599);
nor UO_1579 (O_1579,N_12323,N_14707);
nor UO_1580 (O_1580,N_12403,N_13457);
nor UO_1581 (O_1581,N_13582,N_12678);
nor UO_1582 (O_1582,N_14237,N_14431);
nand UO_1583 (O_1583,N_12272,N_13727);
or UO_1584 (O_1584,N_13309,N_12888);
and UO_1585 (O_1585,N_12312,N_14841);
nor UO_1586 (O_1586,N_13475,N_12850);
or UO_1587 (O_1587,N_12037,N_14072);
nand UO_1588 (O_1588,N_13239,N_12458);
nor UO_1589 (O_1589,N_13406,N_13255);
nand UO_1590 (O_1590,N_13528,N_14598);
or UO_1591 (O_1591,N_13779,N_14325);
or UO_1592 (O_1592,N_14735,N_12702);
nand UO_1593 (O_1593,N_14151,N_13609);
xor UO_1594 (O_1594,N_12175,N_13362);
or UO_1595 (O_1595,N_12240,N_13293);
nor UO_1596 (O_1596,N_14129,N_13483);
and UO_1597 (O_1597,N_13420,N_13022);
nand UO_1598 (O_1598,N_12230,N_14660);
and UO_1599 (O_1599,N_14316,N_14568);
and UO_1600 (O_1600,N_12808,N_12348);
nand UO_1601 (O_1601,N_14452,N_13160);
and UO_1602 (O_1602,N_14737,N_14662);
nand UO_1603 (O_1603,N_12765,N_13978);
nor UO_1604 (O_1604,N_14588,N_12166);
nand UO_1605 (O_1605,N_13164,N_13583);
and UO_1606 (O_1606,N_14622,N_14991);
nor UO_1607 (O_1607,N_13984,N_13987);
nand UO_1608 (O_1608,N_13933,N_14696);
or UO_1609 (O_1609,N_14409,N_14188);
nor UO_1610 (O_1610,N_12560,N_13412);
or UO_1611 (O_1611,N_12762,N_12735);
and UO_1612 (O_1612,N_12808,N_13085);
or UO_1613 (O_1613,N_13901,N_13346);
or UO_1614 (O_1614,N_13392,N_12903);
or UO_1615 (O_1615,N_14379,N_14471);
or UO_1616 (O_1616,N_14760,N_14385);
and UO_1617 (O_1617,N_14288,N_13457);
nand UO_1618 (O_1618,N_14667,N_14902);
nor UO_1619 (O_1619,N_14024,N_12585);
and UO_1620 (O_1620,N_14581,N_14320);
or UO_1621 (O_1621,N_14077,N_14918);
or UO_1622 (O_1622,N_13243,N_13161);
nor UO_1623 (O_1623,N_14044,N_12598);
nor UO_1624 (O_1624,N_12983,N_12011);
and UO_1625 (O_1625,N_14803,N_12499);
nor UO_1626 (O_1626,N_13517,N_13540);
nor UO_1627 (O_1627,N_14237,N_12110);
nor UO_1628 (O_1628,N_13406,N_13857);
and UO_1629 (O_1629,N_13193,N_13048);
and UO_1630 (O_1630,N_12451,N_14003);
and UO_1631 (O_1631,N_12764,N_13069);
nor UO_1632 (O_1632,N_13535,N_14119);
and UO_1633 (O_1633,N_12134,N_13774);
and UO_1634 (O_1634,N_13085,N_14220);
and UO_1635 (O_1635,N_14032,N_14936);
nand UO_1636 (O_1636,N_14936,N_13756);
nor UO_1637 (O_1637,N_14264,N_12483);
and UO_1638 (O_1638,N_13278,N_12116);
and UO_1639 (O_1639,N_12043,N_13343);
or UO_1640 (O_1640,N_13974,N_14290);
or UO_1641 (O_1641,N_12511,N_12223);
and UO_1642 (O_1642,N_13936,N_14679);
nand UO_1643 (O_1643,N_13667,N_12251);
or UO_1644 (O_1644,N_12241,N_14150);
and UO_1645 (O_1645,N_14279,N_13274);
and UO_1646 (O_1646,N_12351,N_13591);
nor UO_1647 (O_1647,N_14525,N_13957);
or UO_1648 (O_1648,N_14383,N_14792);
nand UO_1649 (O_1649,N_14111,N_12104);
nor UO_1650 (O_1650,N_13860,N_13987);
and UO_1651 (O_1651,N_12908,N_13027);
nand UO_1652 (O_1652,N_12126,N_13313);
and UO_1653 (O_1653,N_14487,N_14091);
or UO_1654 (O_1654,N_12000,N_14905);
nand UO_1655 (O_1655,N_12148,N_13626);
and UO_1656 (O_1656,N_12461,N_12949);
nor UO_1657 (O_1657,N_12466,N_14058);
and UO_1658 (O_1658,N_12718,N_14673);
nand UO_1659 (O_1659,N_12595,N_13859);
and UO_1660 (O_1660,N_12263,N_12606);
nand UO_1661 (O_1661,N_12937,N_12507);
and UO_1662 (O_1662,N_12777,N_14300);
nor UO_1663 (O_1663,N_13419,N_12568);
nor UO_1664 (O_1664,N_13931,N_14684);
or UO_1665 (O_1665,N_12955,N_12776);
and UO_1666 (O_1666,N_13348,N_14120);
nor UO_1667 (O_1667,N_12696,N_14099);
and UO_1668 (O_1668,N_14553,N_13292);
or UO_1669 (O_1669,N_13550,N_12778);
nand UO_1670 (O_1670,N_12846,N_13829);
nand UO_1671 (O_1671,N_13203,N_12477);
nand UO_1672 (O_1672,N_13651,N_14472);
or UO_1673 (O_1673,N_14166,N_14454);
nor UO_1674 (O_1674,N_12915,N_12613);
nor UO_1675 (O_1675,N_12758,N_14375);
or UO_1676 (O_1676,N_14122,N_12834);
and UO_1677 (O_1677,N_12040,N_12368);
or UO_1678 (O_1678,N_13674,N_14444);
nor UO_1679 (O_1679,N_12069,N_13940);
and UO_1680 (O_1680,N_14626,N_14560);
nand UO_1681 (O_1681,N_14413,N_14493);
or UO_1682 (O_1682,N_14462,N_12369);
and UO_1683 (O_1683,N_12354,N_14968);
nand UO_1684 (O_1684,N_14519,N_13559);
or UO_1685 (O_1685,N_14828,N_12577);
and UO_1686 (O_1686,N_12337,N_12513);
or UO_1687 (O_1687,N_12124,N_14642);
and UO_1688 (O_1688,N_12582,N_13989);
nand UO_1689 (O_1689,N_12415,N_13266);
nor UO_1690 (O_1690,N_13206,N_12169);
or UO_1691 (O_1691,N_14023,N_14628);
and UO_1692 (O_1692,N_13444,N_13368);
nor UO_1693 (O_1693,N_13023,N_14245);
or UO_1694 (O_1694,N_12291,N_12415);
or UO_1695 (O_1695,N_12691,N_13493);
nor UO_1696 (O_1696,N_13543,N_13239);
or UO_1697 (O_1697,N_12589,N_14374);
nand UO_1698 (O_1698,N_12964,N_12071);
nand UO_1699 (O_1699,N_13258,N_12617);
nand UO_1700 (O_1700,N_12951,N_12190);
nand UO_1701 (O_1701,N_14666,N_14990);
nand UO_1702 (O_1702,N_13139,N_13803);
nor UO_1703 (O_1703,N_14286,N_14027);
nand UO_1704 (O_1704,N_14748,N_14843);
nor UO_1705 (O_1705,N_12296,N_14848);
nand UO_1706 (O_1706,N_14541,N_12804);
or UO_1707 (O_1707,N_13861,N_12128);
nand UO_1708 (O_1708,N_13373,N_12337);
or UO_1709 (O_1709,N_12122,N_14879);
and UO_1710 (O_1710,N_14088,N_14006);
and UO_1711 (O_1711,N_12288,N_12599);
nor UO_1712 (O_1712,N_13048,N_14702);
nand UO_1713 (O_1713,N_14655,N_13227);
or UO_1714 (O_1714,N_12931,N_13611);
nand UO_1715 (O_1715,N_14589,N_14080);
and UO_1716 (O_1716,N_14534,N_13760);
and UO_1717 (O_1717,N_14938,N_13021);
or UO_1718 (O_1718,N_14177,N_14226);
nor UO_1719 (O_1719,N_13391,N_13032);
or UO_1720 (O_1720,N_12493,N_12930);
or UO_1721 (O_1721,N_14609,N_14296);
nor UO_1722 (O_1722,N_13821,N_14667);
nor UO_1723 (O_1723,N_13192,N_13079);
nand UO_1724 (O_1724,N_12356,N_13750);
or UO_1725 (O_1725,N_12850,N_14249);
nor UO_1726 (O_1726,N_14770,N_14624);
and UO_1727 (O_1727,N_12683,N_13421);
or UO_1728 (O_1728,N_13329,N_14648);
nand UO_1729 (O_1729,N_13366,N_14981);
nor UO_1730 (O_1730,N_12926,N_12340);
nor UO_1731 (O_1731,N_12876,N_12423);
or UO_1732 (O_1732,N_14066,N_13818);
nor UO_1733 (O_1733,N_12236,N_12500);
nor UO_1734 (O_1734,N_12878,N_12186);
and UO_1735 (O_1735,N_13484,N_12990);
nand UO_1736 (O_1736,N_14141,N_13308);
nor UO_1737 (O_1737,N_12333,N_12386);
or UO_1738 (O_1738,N_13316,N_13924);
or UO_1739 (O_1739,N_12340,N_12932);
or UO_1740 (O_1740,N_14194,N_13121);
or UO_1741 (O_1741,N_12590,N_14013);
xor UO_1742 (O_1742,N_14421,N_12150);
and UO_1743 (O_1743,N_14113,N_14430);
and UO_1744 (O_1744,N_13013,N_13860);
nand UO_1745 (O_1745,N_13168,N_12649);
nor UO_1746 (O_1746,N_14238,N_14393);
nand UO_1747 (O_1747,N_13271,N_14732);
or UO_1748 (O_1748,N_13851,N_12760);
or UO_1749 (O_1749,N_14646,N_12871);
and UO_1750 (O_1750,N_12731,N_13724);
nor UO_1751 (O_1751,N_14041,N_12737);
nand UO_1752 (O_1752,N_12518,N_12556);
nand UO_1753 (O_1753,N_12209,N_14394);
nor UO_1754 (O_1754,N_13179,N_12476);
or UO_1755 (O_1755,N_12835,N_13152);
nand UO_1756 (O_1756,N_13831,N_13092);
and UO_1757 (O_1757,N_14351,N_13493);
nand UO_1758 (O_1758,N_12878,N_13867);
nor UO_1759 (O_1759,N_13564,N_14036);
nor UO_1760 (O_1760,N_12254,N_14501);
nor UO_1761 (O_1761,N_12572,N_12197);
nor UO_1762 (O_1762,N_13609,N_14510);
nand UO_1763 (O_1763,N_12547,N_12428);
or UO_1764 (O_1764,N_13948,N_13920);
and UO_1765 (O_1765,N_14238,N_13280);
nor UO_1766 (O_1766,N_14423,N_13677);
nor UO_1767 (O_1767,N_14945,N_13745);
nor UO_1768 (O_1768,N_13607,N_13826);
nand UO_1769 (O_1769,N_14830,N_12760);
or UO_1770 (O_1770,N_13808,N_12411);
and UO_1771 (O_1771,N_14805,N_13375);
nor UO_1772 (O_1772,N_13376,N_14724);
nand UO_1773 (O_1773,N_12884,N_12230);
or UO_1774 (O_1774,N_12970,N_13044);
and UO_1775 (O_1775,N_12754,N_12577);
nand UO_1776 (O_1776,N_12653,N_14757);
nor UO_1777 (O_1777,N_14953,N_12624);
or UO_1778 (O_1778,N_12182,N_12095);
nor UO_1779 (O_1779,N_14726,N_14443);
and UO_1780 (O_1780,N_14040,N_14671);
nor UO_1781 (O_1781,N_14448,N_13740);
and UO_1782 (O_1782,N_12316,N_14663);
nor UO_1783 (O_1783,N_13929,N_12805);
nand UO_1784 (O_1784,N_13285,N_14479);
and UO_1785 (O_1785,N_13368,N_12660);
nor UO_1786 (O_1786,N_12898,N_14766);
or UO_1787 (O_1787,N_13174,N_14886);
and UO_1788 (O_1788,N_13286,N_14205);
nand UO_1789 (O_1789,N_14199,N_14651);
nor UO_1790 (O_1790,N_13913,N_12086);
nor UO_1791 (O_1791,N_14525,N_13539);
nand UO_1792 (O_1792,N_13611,N_12364);
and UO_1793 (O_1793,N_13160,N_12481);
nand UO_1794 (O_1794,N_12419,N_12562);
and UO_1795 (O_1795,N_13684,N_14512);
nand UO_1796 (O_1796,N_14662,N_13573);
nand UO_1797 (O_1797,N_12753,N_12363);
and UO_1798 (O_1798,N_12047,N_14741);
nand UO_1799 (O_1799,N_14397,N_13550);
nand UO_1800 (O_1800,N_14653,N_14438);
nor UO_1801 (O_1801,N_13957,N_12438);
nand UO_1802 (O_1802,N_13324,N_14911);
nor UO_1803 (O_1803,N_14337,N_13872);
or UO_1804 (O_1804,N_13937,N_14651);
or UO_1805 (O_1805,N_14887,N_13823);
nor UO_1806 (O_1806,N_12230,N_14890);
nand UO_1807 (O_1807,N_14897,N_12485);
or UO_1808 (O_1808,N_12157,N_13016);
and UO_1809 (O_1809,N_13559,N_13594);
nor UO_1810 (O_1810,N_13520,N_12214);
nand UO_1811 (O_1811,N_12409,N_13175);
nor UO_1812 (O_1812,N_13762,N_14072);
and UO_1813 (O_1813,N_12849,N_14780);
nor UO_1814 (O_1814,N_12862,N_13468);
nand UO_1815 (O_1815,N_14139,N_13900);
nor UO_1816 (O_1816,N_14116,N_14387);
nand UO_1817 (O_1817,N_14078,N_13922);
nand UO_1818 (O_1818,N_14289,N_12028);
nor UO_1819 (O_1819,N_14606,N_13063);
and UO_1820 (O_1820,N_14992,N_12220);
nor UO_1821 (O_1821,N_12932,N_14442);
nor UO_1822 (O_1822,N_12656,N_13803);
nand UO_1823 (O_1823,N_12117,N_12820);
nor UO_1824 (O_1824,N_14012,N_14457);
nand UO_1825 (O_1825,N_12910,N_13028);
or UO_1826 (O_1826,N_12530,N_13376);
nand UO_1827 (O_1827,N_12073,N_12318);
and UO_1828 (O_1828,N_12056,N_13244);
or UO_1829 (O_1829,N_14156,N_13215);
nor UO_1830 (O_1830,N_13434,N_14214);
and UO_1831 (O_1831,N_14894,N_12899);
and UO_1832 (O_1832,N_14728,N_14710);
and UO_1833 (O_1833,N_13520,N_13864);
and UO_1834 (O_1834,N_14531,N_13058);
and UO_1835 (O_1835,N_12422,N_12816);
or UO_1836 (O_1836,N_14471,N_13303);
nor UO_1837 (O_1837,N_14427,N_14768);
and UO_1838 (O_1838,N_12873,N_12936);
nor UO_1839 (O_1839,N_13006,N_13072);
nand UO_1840 (O_1840,N_12063,N_13968);
nand UO_1841 (O_1841,N_13205,N_14665);
nor UO_1842 (O_1842,N_14303,N_12042);
or UO_1843 (O_1843,N_14196,N_13605);
and UO_1844 (O_1844,N_13639,N_13975);
or UO_1845 (O_1845,N_13650,N_14062);
nor UO_1846 (O_1846,N_13573,N_12294);
or UO_1847 (O_1847,N_14562,N_12668);
or UO_1848 (O_1848,N_13324,N_13552);
nand UO_1849 (O_1849,N_12990,N_12854);
xor UO_1850 (O_1850,N_12609,N_12128);
nor UO_1851 (O_1851,N_13865,N_12771);
nand UO_1852 (O_1852,N_12724,N_12658);
and UO_1853 (O_1853,N_12668,N_14359);
and UO_1854 (O_1854,N_13342,N_12608);
nand UO_1855 (O_1855,N_13681,N_14457);
nor UO_1856 (O_1856,N_13944,N_14038);
nor UO_1857 (O_1857,N_12478,N_14120);
and UO_1858 (O_1858,N_12545,N_14214);
nor UO_1859 (O_1859,N_13356,N_13708);
nor UO_1860 (O_1860,N_14113,N_13516);
or UO_1861 (O_1861,N_13514,N_12525);
or UO_1862 (O_1862,N_14614,N_13505);
and UO_1863 (O_1863,N_12541,N_13839);
or UO_1864 (O_1864,N_13905,N_12903);
nor UO_1865 (O_1865,N_13079,N_14945);
nand UO_1866 (O_1866,N_13159,N_12072);
nor UO_1867 (O_1867,N_12570,N_12155);
nand UO_1868 (O_1868,N_14883,N_12381);
or UO_1869 (O_1869,N_12828,N_13345);
and UO_1870 (O_1870,N_13262,N_13679);
nor UO_1871 (O_1871,N_13324,N_14170);
or UO_1872 (O_1872,N_14928,N_12560);
nand UO_1873 (O_1873,N_14650,N_13642);
nor UO_1874 (O_1874,N_14150,N_12762);
or UO_1875 (O_1875,N_14240,N_13484);
and UO_1876 (O_1876,N_14833,N_12883);
and UO_1877 (O_1877,N_13308,N_13538);
nor UO_1878 (O_1878,N_12442,N_12838);
nand UO_1879 (O_1879,N_13282,N_14820);
nand UO_1880 (O_1880,N_12071,N_14818);
or UO_1881 (O_1881,N_14763,N_13104);
or UO_1882 (O_1882,N_14030,N_14196);
or UO_1883 (O_1883,N_13173,N_14496);
or UO_1884 (O_1884,N_13343,N_12828);
or UO_1885 (O_1885,N_13862,N_12706);
or UO_1886 (O_1886,N_12200,N_12174);
nand UO_1887 (O_1887,N_14735,N_14167);
or UO_1888 (O_1888,N_13577,N_14880);
and UO_1889 (O_1889,N_14952,N_12689);
and UO_1890 (O_1890,N_14904,N_13349);
nand UO_1891 (O_1891,N_12479,N_12539);
nor UO_1892 (O_1892,N_14656,N_13543);
and UO_1893 (O_1893,N_14983,N_13874);
nand UO_1894 (O_1894,N_13302,N_12725);
and UO_1895 (O_1895,N_13728,N_13271);
nor UO_1896 (O_1896,N_12339,N_12063);
nor UO_1897 (O_1897,N_13597,N_12541);
or UO_1898 (O_1898,N_14650,N_12160);
and UO_1899 (O_1899,N_14751,N_13581);
nor UO_1900 (O_1900,N_14297,N_12268);
nor UO_1901 (O_1901,N_12788,N_14081);
nand UO_1902 (O_1902,N_14825,N_14739);
or UO_1903 (O_1903,N_13378,N_12078);
or UO_1904 (O_1904,N_13149,N_12832);
nor UO_1905 (O_1905,N_13294,N_14593);
nand UO_1906 (O_1906,N_12302,N_14105);
or UO_1907 (O_1907,N_13515,N_14495);
and UO_1908 (O_1908,N_13831,N_14738);
and UO_1909 (O_1909,N_13450,N_12901);
and UO_1910 (O_1910,N_14236,N_14230);
nor UO_1911 (O_1911,N_14485,N_13152);
nand UO_1912 (O_1912,N_14915,N_13870);
and UO_1913 (O_1913,N_13684,N_13045);
nand UO_1914 (O_1914,N_12931,N_12421);
or UO_1915 (O_1915,N_14340,N_13076);
and UO_1916 (O_1916,N_13596,N_12003);
or UO_1917 (O_1917,N_12224,N_14670);
nand UO_1918 (O_1918,N_13420,N_13652);
nor UO_1919 (O_1919,N_14656,N_12315);
or UO_1920 (O_1920,N_14491,N_12272);
nand UO_1921 (O_1921,N_13458,N_14081);
nor UO_1922 (O_1922,N_14829,N_12602);
and UO_1923 (O_1923,N_13648,N_12839);
nor UO_1924 (O_1924,N_12925,N_13831);
or UO_1925 (O_1925,N_12393,N_12741);
nand UO_1926 (O_1926,N_13444,N_12265);
nand UO_1927 (O_1927,N_14943,N_13776);
nand UO_1928 (O_1928,N_14564,N_12473);
nand UO_1929 (O_1929,N_14824,N_12393);
nor UO_1930 (O_1930,N_12528,N_14632);
or UO_1931 (O_1931,N_12170,N_13980);
nand UO_1932 (O_1932,N_14923,N_13917);
nand UO_1933 (O_1933,N_13330,N_14298);
and UO_1934 (O_1934,N_12094,N_14447);
nor UO_1935 (O_1935,N_12344,N_13332);
nand UO_1936 (O_1936,N_12001,N_13528);
and UO_1937 (O_1937,N_13337,N_12962);
nor UO_1938 (O_1938,N_13009,N_14639);
and UO_1939 (O_1939,N_14419,N_13329);
nor UO_1940 (O_1940,N_13044,N_12966);
and UO_1941 (O_1941,N_12748,N_14756);
and UO_1942 (O_1942,N_12581,N_12959);
nand UO_1943 (O_1943,N_14298,N_13425);
nand UO_1944 (O_1944,N_14181,N_14461);
and UO_1945 (O_1945,N_13646,N_14245);
and UO_1946 (O_1946,N_14014,N_13523);
nor UO_1947 (O_1947,N_13486,N_14218);
nor UO_1948 (O_1948,N_14153,N_14587);
nor UO_1949 (O_1949,N_12563,N_14706);
and UO_1950 (O_1950,N_12679,N_14770);
nand UO_1951 (O_1951,N_12123,N_13394);
and UO_1952 (O_1952,N_14901,N_12782);
nand UO_1953 (O_1953,N_12546,N_14135);
or UO_1954 (O_1954,N_14142,N_12244);
nand UO_1955 (O_1955,N_12176,N_14786);
and UO_1956 (O_1956,N_12827,N_14907);
or UO_1957 (O_1957,N_12053,N_13909);
or UO_1958 (O_1958,N_14091,N_12429);
nor UO_1959 (O_1959,N_13459,N_12177);
nand UO_1960 (O_1960,N_12887,N_14676);
nor UO_1961 (O_1961,N_12630,N_13884);
nor UO_1962 (O_1962,N_12384,N_12713);
nor UO_1963 (O_1963,N_12684,N_14415);
or UO_1964 (O_1964,N_14590,N_13230);
nand UO_1965 (O_1965,N_13054,N_12894);
and UO_1966 (O_1966,N_14509,N_13370);
nor UO_1967 (O_1967,N_13642,N_14523);
or UO_1968 (O_1968,N_12120,N_12589);
nor UO_1969 (O_1969,N_13863,N_14008);
nor UO_1970 (O_1970,N_14925,N_13764);
nand UO_1971 (O_1971,N_12255,N_12712);
nor UO_1972 (O_1972,N_12494,N_14259);
and UO_1973 (O_1973,N_13233,N_14844);
nor UO_1974 (O_1974,N_13635,N_12785);
nand UO_1975 (O_1975,N_12570,N_13987);
or UO_1976 (O_1976,N_12173,N_12532);
or UO_1977 (O_1977,N_12931,N_12381);
nand UO_1978 (O_1978,N_13541,N_12032);
nand UO_1979 (O_1979,N_14900,N_13518);
and UO_1980 (O_1980,N_14633,N_13528);
nand UO_1981 (O_1981,N_12728,N_12367);
and UO_1982 (O_1982,N_14206,N_12869);
and UO_1983 (O_1983,N_13185,N_14653);
nand UO_1984 (O_1984,N_12343,N_12350);
nand UO_1985 (O_1985,N_12062,N_13082);
nor UO_1986 (O_1986,N_13244,N_12793);
or UO_1987 (O_1987,N_13818,N_12719);
or UO_1988 (O_1988,N_14198,N_13546);
nor UO_1989 (O_1989,N_14873,N_14664);
or UO_1990 (O_1990,N_13094,N_12656);
nor UO_1991 (O_1991,N_14528,N_14097);
and UO_1992 (O_1992,N_13072,N_13904);
nand UO_1993 (O_1993,N_14126,N_13626);
and UO_1994 (O_1994,N_14428,N_14317);
and UO_1995 (O_1995,N_12670,N_14302);
and UO_1996 (O_1996,N_13373,N_12084);
nor UO_1997 (O_1997,N_13617,N_14997);
or UO_1998 (O_1998,N_14406,N_12270);
and UO_1999 (O_1999,N_14551,N_12553);
endmodule