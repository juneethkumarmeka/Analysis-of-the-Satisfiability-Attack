module basic_500_3000_500_30_levels_2xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_108,In_23);
nand U1 (N_1,In_131,In_235);
or U2 (N_2,In_269,In_15);
xor U3 (N_3,In_326,In_316);
and U4 (N_4,In_340,In_221);
nand U5 (N_5,In_29,In_163);
nor U6 (N_6,In_72,In_452);
or U7 (N_7,In_404,In_483);
or U8 (N_8,In_164,In_265);
nor U9 (N_9,In_142,In_188);
nor U10 (N_10,In_320,In_226);
nand U11 (N_11,In_247,In_484);
nand U12 (N_12,In_26,In_444);
and U13 (N_13,In_127,In_300);
nand U14 (N_14,In_465,In_437);
nor U15 (N_15,In_302,In_412);
or U16 (N_16,In_372,In_330);
nand U17 (N_17,In_84,In_449);
nor U18 (N_18,In_463,In_18);
and U19 (N_19,In_357,In_301);
nand U20 (N_20,In_224,In_119);
and U21 (N_21,In_85,In_332);
and U22 (N_22,In_289,In_7);
nor U23 (N_23,In_443,In_432);
nand U24 (N_24,In_71,In_280);
nor U25 (N_25,In_175,In_42);
and U26 (N_26,In_322,In_485);
nor U27 (N_27,In_376,In_91);
or U28 (N_28,In_161,In_136);
or U29 (N_29,In_475,In_411);
or U30 (N_30,In_88,In_130);
or U31 (N_31,In_474,In_408);
and U32 (N_32,In_407,In_450);
and U33 (N_33,In_364,In_219);
nand U34 (N_34,In_342,In_196);
and U35 (N_35,In_422,In_214);
or U36 (N_36,In_410,In_370);
nand U37 (N_37,In_109,In_406);
nand U38 (N_38,In_191,In_95);
or U39 (N_39,In_166,In_321);
nand U40 (N_40,In_67,In_327);
nor U41 (N_41,In_305,In_436);
nor U42 (N_42,In_377,In_120);
or U43 (N_43,In_49,In_202);
nand U44 (N_44,In_152,In_464);
and U45 (N_45,In_156,In_424);
nor U46 (N_46,In_295,In_11);
and U47 (N_47,In_126,In_276);
nand U48 (N_48,In_386,In_54);
and U49 (N_49,In_24,In_21);
nor U50 (N_50,In_70,In_168);
nand U51 (N_51,In_180,In_195);
nand U52 (N_52,In_471,In_60);
nand U53 (N_53,In_293,In_256);
or U54 (N_54,In_129,In_204);
nand U55 (N_55,In_241,In_262);
nor U56 (N_56,In_368,In_251);
nor U57 (N_57,In_104,In_27);
and U58 (N_58,In_493,In_283);
or U59 (N_59,In_213,In_299);
nor U60 (N_60,In_296,In_157);
or U61 (N_61,In_499,In_413);
nor U62 (N_62,In_43,In_466);
nand U63 (N_63,In_110,In_16);
or U64 (N_64,In_239,In_496);
or U65 (N_65,In_121,In_456);
nor U66 (N_66,In_143,In_480);
nand U67 (N_67,In_440,In_97);
nor U68 (N_68,In_489,In_186);
nand U69 (N_69,In_417,In_55);
or U70 (N_70,In_113,In_341);
nor U71 (N_71,In_47,In_260);
and U72 (N_72,In_201,In_114);
or U73 (N_73,In_392,In_420);
nand U74 (N_74,In_249,In_398);
nand U75 (N_75,In_277,In_61);
nor U76 (N_76,In_315,In_428);
nand U77 (N_77,In_2,In_292);
nand U78 (N_78,In_179,In_137);
nor U79 (N_79,In_101,In_73);
and U80 (N_80,In_310,In_461);
and U81 (N_81,In_323,In_405);
nand U82 (N_82,In_116,In_8);
or U83 (N_83,In_150,In_497);
or U84 (N_84,In_100,In_438);
nor U85 (N_85,In_76,In_154);
nor U86 (N_86,In_379,In_375);
or U87 (N_87,In_185,In_355);
or U88 (N_88,In_259,In_177);
and U89 (N_89,In_271,In_106);
nand U90 (N_90,In_267,In_275);
or U91 (N_91,In_374,In_181);
nand U92 (N_92,In_288,In_335);
nand U93 (N_93,In_176,In_402);
or U94 (N_94,In_3,In_442);
nor U95 (N_95,In_381,In_380);
or U96 (N_96,In_365,In_98);
nor U97 (N_97,In_90,In_74);
and U98 (N_98,In_286,In_146);
or U99 (N_99,In_20,In_318);
and U100 (N_100,In_347,In_486);
nor U101 (N_101,In_273,N_99);
and U102 (N_102,In_345,In_385);
and U103 (N_103,In_190,In_348);
or U104 (N_104,N_88,In_139);
or U105 (N_105,N_25,N_14);
nor U106 (N_106,In_240,In_434);
nand U107 (N_107,N_75,In_314);
or U108 (N_108,In_215,In_93);
and U109 (N_109,In_56,N_49);
or U110 (N_110,N_68,In_83);
or U111 (N_111,In_22,In_457);
or U112 (N_112,In_94,In_263);
and U113 (N_113,In_253,In_37);
nor U114 (N_114,In_31,N_9);
and U115 (N_115,In_250,In_306);
or U116 (N_116,In_311,N_98);
nand U117 (N_117,In_401,N_64);
nand U118 (N_118,In_81,In_282);
nand U119 (N_119,In_303,In_68);
or U120 (N_120,N_10,In_89);
nand U121 (N_121,In_173,N_22);
and U122 (N_122,N_20,In_135);
and U123 (N_123,N_23,In_171);
xor U124 (N_124,In_133,In_445);
and U125 (N_125,In_414,In_298);
nor U126 (N_126,N_18,In_361);
and U127 (N_127,In_193,In_159);
and U128 (N_128,N_83,In_231);
nand U129 (N_129,N_70,In_459);
and U130 (N_130,In_418,N_90);
nor U131 (N_131,In_59,N_29);
and U132 (N_132,In_165,N_94);
nand U133 (N_133,In_170,In_75);
nand U134 (N_134,In_352,In_237);
and U135 (N_135,In_25,In_52);
nand U136 (N_136,N_73,In_132);
or U137 (N_137,In_158,In_236);
and U138 (N_138,In_328,In_384);
and U139 (N_139,In_454,N_71);
or U140 (N_140,N_67,In_426);
xor U141 (N_141,N_39,In_346);
nor U142 (N_142,In_210,In_439);
and U143 (N_143,N_19,In_387);
nand U144 (N_144,In_107,In_391);
nand U145 (N_145,N_2,In_495);
nand U146 (N_146,In_488,In_69);
or U147 (N_147,N_50,N_41);
xnor U148 (N_148,In_467,In_13);
or U149 (N_149,N_78,In_350);
or U150 (N_150,In_230,In_285);
and U151 (N_151,In_344,In_393);
and U152 (N_152,In_212,In_460);
and U153 (N_153,In_366,In_334);
and U154 (N_154,In_220,In_112);
and U155 (N_155,In_478,In_32);
or U156 (N_156,N_72,In_206);
and U157 (N_157,In_498,In_198);
nand U158 (N_158,In_244,In_6);
nand U159 (N_159,N_60,In_308);
or U160 (N_160,In_144,In_10);
and U161 (N_161,In_338,In_360);
nor U162 (N_162,N_63,N_26);
and U163 (N_163,In_45,In_272);
and U164 (N_164,N_1,N_15);
and U165 (N_165,In_397,In_469);
nor U166 (N_166,In_278,In_205);
and U167 (N_167,In_359,N_6);
nand U168 (N_168,In_229,In_87);
or U169 (N_169,In_30,N_37);
or U170 (N_170,N_89,In_4);
and U171 (N_171,In_363,In_390);
nor U172 (N_172,In_153,In_228);
or U173 (N_173,In_351,In_431);
and U174 (N_174,In_79,In_403);
nand U175 (N_175,N_51,In_243);
nor U176 (N_176,In_35,In_383);
or U177 (N_177,N_42,In_184);
nor U178 (N_178,N_57,In_33);
nand U179 (N_179,N_33,In_50);
and U180 (N_180,In_105,In_473);
nand U181 (N_181,N_82,In_118);
or U182 (N_182,N_8,In_297);
nand U183 (N_183,In_138,In_476);
or U184 (N_184,N_40,N_31);
or U185 (N_185,In_468,In_223);
or U186 (N_186,In_266,N_46);
or U187 (N_187,In_458,N_84);
nand U188 (N_188,In_416,In_233);
or U189 (N_189,In_58,In_446);
and U190 (N_190,N_34,In_246);
or U191 (N_191,In_167,In_234);
and U192 (N_192,In_304,N_38);
nor U193 (N_193,In_382,N_81);
and U194 (N_194,In_312,In_255);
and U195 (N_195,In_399,In_189);
nor U196 (N_196,In_423,In_441);
xor U197 (N_197,In_287,In_169);
nand U198 (N_198,In_86,In_435);
nor U199 (N_199,In_325,In_279);
or U200 (N_200,In_38,N_111);
and U201 (N_201,N_24,N_114);
or U202 (N_202,In_261,N_109);
or U203 (N_203,In_19,In_477);
xnor U204 (N_204,In_151,In_462);
nor U205 (N_205,In_80,In_281);
nand U206 (N_206,In_394,In_183);
or U207 (N_207,In_41,N_115);
nor U208 (N_208,In_17,In_472);
nand U209 (N_209,N_145,N_151);
nand U210 (N_210,In_122,In_140);
and U211 (N_211,N_188,In_470);
nor U212 (N_212,In_57,N_119);
nand U213 (N_213,In_82,N_80);
nand U214 (N_214,N_170,N_152);
nand U215 (N_215,In_14,In_217);
and U216 (N_216,In_232,In_174);
and U217 (N_217,In_258,In_369);
xnor U218 (N_218,N_69,N_138);
or U219 (N_219,N_143,In_78);
and U220 (N_220,In_200,N_139);
or U221 (N_221,In_389,N_169);
nand U222 (N_222,N_96,In_182);
or U223 (N_223,In_66,In_487);
or U224 (N_224,In_162,In_36);
nor U225 (N_225,In_395,In_194);
nand U226 (N_226,In_216,N_191);
nor U227 (N_227,In_491,N_192);
nor U228 (N_228,N_155,In_451);
nand U229 (N_229,In_203,In_155);
nand U230 (N_230,In_453,N_59);
nor U231 (N_231,N_161,N_86);
nand U232 (N_232,In_252,In_329);
and U233 (N_233,N_184,In_362);
and U234 (N_234,In_447,N_54);
nor U235 (N_235,In_494,N_124);
or U236 (N_236,In_337,N_56);
nand U237 (N_237,In_433,In_53);
nor U238 (N_238,N_32,In_63);
nor U239 (N_239,In_343,N_0);
xor U240 (N_240,In_429,In_147);
or U241 (N_241,In_207,In_160);
or U242 (N_242,In_294,In_141);
or U243 (N_243,N_171,N_194);
or U244 (N_244,N_61,In_92);
nand U245 (N_245,N_44,In_425);
nor U246 (N_246,N_122,In_28);
nand U247 (N_247,N_12,N_43);
or U248 (N_248,N_93,N_167);
nor U249 (N_249,In_111,In_248);
nor U250 (N_250,In_358,In_307);
nor U251 (N_251,N_150,N_162);
nor U252 (N_252,N_164,In_96);
nor U253 (N_253,N_183,In_481);
or U254 (N_254,N_95,In_245);
or U255 (N_255,N_45,In_218);
or U256 (N_256,N_128,In_339);
or U257 (N_257,In_192,N_117);
nor U258 (N_258,In_427,In_254);
or U259 (N_259,In_371,N_105);
or U260 (N_260,N_153,N_66);
and U261 (N_261,In_115,N_157);
nand U262 (N_262,N_113,N_126);
nor U263 (N_263,In_64,In_356);
nor U264 (N_264,In_145,In_5);
nor U265 (N_265,N_197,N_17);
nand U266 (N_266,In_396,N_121);
or U267 (N_267,In_187,N_100);
nor U268 (N_268,N_3,N_97);
or U269 (N_269,N_134,N_92);
nor U270 (N_270,N_16,In_40);
nor U271 (N_271,In_128,In_336);
nand U272 (N_272,N_140,N_185);
or U273 (N_273,In_290,N_27);
nor U274 (N_274,N_166,N_149);
or U275 (N_275,In_291,In_373);
nor U276 (N_276,N_106,N_13);
and U277 (N_277,N_129,N_62);
or U278 (N_278,N_137,N_146);
or U279 (N_279,In_222,N_176);
or U280 (N_280,In_238,In_482);
nor U281 (N_281,N_160,In_172);
or U282 (N_282,N_55,In_0);
or U283 (N_283,In_313,N_172);
and U284 (N_284,In_39,N_159);
or U285 (N_285,In_333,N_168);
or U286 (N_286,N_120,In_117);
nand U287 (N_287,In_134,N_180);
nor U288 (N_288,In_242,In_309);
and U289 (N_289,N_116,N_165);
nor U290 (N_290,N_48,In_378);
nor U291 (N_291,N_130,N_189);
and U292 (N_292,In_208,In_415);
or U293 (N_293,N_125,N_133);
or U294 (N_294,In_349,N_147);
or U295 (N_295,In_51,In_34);
nand U296 (N_296,N_11,In_149);
nor U297 (N_297,In_479,N_107);
or U298 (N_298,N_4,N_77);
nor U299 (N_299,N_79,In_44);
nor U300 (N_300,N_265,N_212);
or U301 (N_301,N_246,N_298);
nor U302 (N_302,N_216,N_276);
and U303 (N_303,N_235,N_76);
nor U304 (N_304,N_7,N_21);
or U305 (N_305,N_214,N_173);
xor U306 (N_306,N_205,N_277);
nor U307 (N_307,N_253,N_209);
nand U308 (N_308,N_179,N_263);
or U309 (N_309,N_175,N_47);
nor U310 (N_310,N_28,N_177);
nand U311 (N_311,N_297,N_231);
nor U312 (N_312,In_48,In_331);
nor U313 (N_313,N_221,N_230);
nor U314 (N_314,N_36,N_201);
nand U315 (N_315,N_206,In_409);
or U316 (N_316,N_200,N_144);
nand U317 (N_317,In_65,N_275);
nand U318 (N_318,N_190,N_252);
nor U319 (N_319,N_279,N_136);
xnor U320 (N_320,N_284,In_400);
and U321 (N_321,N_53,N_178);
or U322 (N_322,In_225,N_248);
and U323 (N_323,N_283,In_46);
or U324 (N_324,N_181,N_196);
or U325 (N_325,N_102,In_1);
nor U326 (N_326,N_245,In_284);
nand U327 (N_327,N_232,N_154);
and U328 (N_328,N_255,In_448);
nor U329 (N_329,N_259,In_9);
or U330 (N_330,N_272,N_226);
nor U331 (N_331,N_187,In_148);
nand U332 (N_332,In_324,In_274);
nor U333 (N_333,In_270,In_102);
or U334 (N_334,N_236,N_224);
and U335 (N_335,N_261,N_285);
nand U336 (N_336,N_241,N_290);
nand U337 (N_337,In_492,N_103);
xnor U338 (N_338,N_132,In_123);
and U339 (N_339,N_233,N_158);
and U340 (N_340,In_257,In_77);
nand U341 (N_341,In_124,N_219);
or U342 (N_342,N_267,N_174);
nor U343 (N_343,In_12,N_273);
xnor U344 (N_344,N_286,N_289);
or U345 (N_345,N_249,In_99);
nor U346 (N_346,N_30,N_110);
xnor U347 (N_347,N_215,N_156);
or U348 (N_348,In_209,N_199);
nand U349 (N_349,N_186,N_198);
or U350 (N_350,In_353,In_319);
and U351 (N_351,N_244,In_227);
xnor U352 (N_352,In_419,N_207);
and U353 (N_353,N_251,N_195);
nor U354 (N_354,In_421,N_218);
nor U355 (N_355,N_296,N_268);
and U356 (N_356,In_211,In_103);
or U357 (N_357,N_5,N_229);
nor U358 (N_358,N_292,N_141);
nor U359 (N_359,N_250,In_268);
or U360 (N_360,N_208,N_280);
and U361 (N_361,N_266,N_257);
or U362 (N_362,N_211,N_243);
or U363 (N_363,N_223,In_367);
and U364 (N_364,N_287,N_274);
nor U365 (N_365,N_203,N_217);
and U366 (N_366,N_123,N_58);
or U367 (N_367,N_256,N_85);
or U368 (N_368,N_127,N_278);
nand U369 (N_369,N_87,N_293);
and U370 (N_370,In_354,In_199);
or U371 (N_371,N_291,N_288);
or U372 (N_372,N_299,N_225);
and U373 (N_373,N_271,N_239);
xnor U374 (N_374,N_108,N_240);
nand U375 (N_375,N_193,N_202);
nor U376 (N_376,N_52,N_204);
nand U377 (N_377,N_227,N_112);
nand U378 (N_378,N_269,N_131);
nand U379 (N_379,N_182,N_238);
nor U380 (N_380,N_247,In_125);
nor U381 (N_381,In_62,In_388);
and U382 (N_382,N_254,N_220);
and U383 (N_383,N_163,N_91);
nand U384 (N_384,N_228,N_104);
or U385 (N_385,N_270,N_118);
nand U386 (N_386,N_101,N_142);
and U387 (N_387,N_264,In_264);
nor U388 (N_388,N_74,In_490);
xnor U389 (N_389,In_317,N_242);
nand U390 (N_390,N_294,In_178);
or U391 (N_391,N_260,N_148);
or U392 (N_392,In_430,N_282);
nor U393 (N_393,In_197,N_237);
or U394 (N_394,N_135,N_210);
nand U395 (N_395,N_258,N_262);
nor U396 (N_396,N_65,N_234);
nand U397 (N_397,In_455,N_213);
nand U398 (N_398,N_295,N_281);
and U399 (N_399,N_35,N_222);
nor U400 (N_400,N_335,N_327);
nor U401 (N_401,N_319,N_313);
nand U402 (N_402,N_324,N_315);
nand U403 (N_403,N_320,N_358);
nor U404 (N_404,N_378,N_340);
nor U405 (N_405,N_317,N_373);
nor U406 (N_406,N_351,N_354);
xnor U407 (N_407,N_381,N_308);
nand U408 (N_408,N_300,N_388);
nand U409 (N_409,N_359,N_383);
and U410 (N_410,N_370,N_312);
or U411 (N_411,N_323,N_379);
or U412 (N_412,N_366,N_303);
and U413 (N_413,N_380,N_399);
and U414 (N_414,N_334,N_342);
nand U415 (N_415,N_352,N_325);
or U416 (N_416,N_360,N_329);
nor U417 (N_417,N_392,N_328);
nor U418 (N_418,N_356,N_332);
nor U419 (N_419,N_384,N_367);
or U420 (N_420,N_353,N_348);
nor U421 (N_421,N_344,N_387);
nor U422 (N_422,N_385,N_371);
and U423 (N_423,N_389,N_337);
or U424 (N_424,N_304,N_322);
and U425 (N_425,N_316,N_333);
nor U426 (N_426,N_311,N_369);
and U427 (N_427,N_345,N_394);
xnor U428 (N_428,N_355,N_302);
or U429 (N_429,N_363,N_364);
or U430 (N_430,N_314,N_339);
or U431 (N_431,N_330,N_395);
nor U432 (N_432,N_307,N_372);
nor U433 (N_433,N_398,N_326);
and U434 (N_434,N_343,N_331);
nand U435 (N_435,N_349,N_362);
nor U436 (N_436,N_357,N_318);
nor U437 (N_437,N_350,N_361);
nor U438 (N_438,N_305,N_336);
xor U439 (N_439,N_374,N_365);
nor U440 (N_440,N_306,N_368);
nor U441 (N_441,N_321,N_391);
xor U442 (N_442,N_376,N_386);
nor U443 (N_443,N_375,N_346);
or U444 (N_444,N_309,N_338);
nand U445 (N_445,N_341,N_382);
or U446 (N_446,N_377,N_396);
and U447 (N_447,N_393,N_301);
and U448 (N_448,N_390,N_397);
nand U449 (N_449,N_347,N_310);
and U450 (N_450,N_387,N_330);
and U451 (N_451,N_339,N_323);
and U452 (N_452,N_393,N_324);
or U453 (N_453,N_307,N_388);
nor U454 (N_454,N_367,N_323);
or U455 (N_455,N_382,N_320);
or U456 (N_456,N_325,N_312);
or U457 (N_457,N_319,N_352);
or U458 (N_458,N_330,N_393);
or U459 (N_459,N_370,N_339);
nor U460 (N_460,N_310,N_344);
and U461 (N_461,N_303,N_314);
or U462 (N_462,N_357,N_375);
nand U463 (N_463,N_344,N_353);
xnor U464 (N_464,N_302,N_361);
and U465 (N_465,N_330,N_333);
nand U466 (N_466,N_387,N_319);
or U467 (N_467,N_395,N_373);
and U468 (N_468,N_376,N_389);
and U469 (N_469,N_370,N_385);
or U470 (N_470,N_345,N_384);
nor U471 (N_471,N_399,N_387);
nand U472 (N_472,N_308,N_396);
or U473 (N_473,N_346,N_373);
and U474 (N_474,N_338,N_396);
and U475 (N_475,N_399,N_355);
nand U476 (N_476,N_330,N_319);
or U477 (N_477,N_356,N_375);
nor U478 (N_478,N_329,N_388);
or U479 (N_479,N_355,N_380);
nor U480 (N_480,N_355,N_397);
nor U481 (N_481,N_327,N_348);
nand U482 (N_482,N_303,N_393);
nor U483 (N_483,N_362,N_322);
and U484 (N_484,N_354,N_308);
nor U485 (N_485,N_398,N_394);
nand U486 (N_486,N_302,N_362);
and U487 (N_487,N_325,N_318);
nand U488 (N_488,N_396,N_300);
or U489 (N_489,N_360,N_306);
or U490 (N_490,N_348,N_358);
nand U491 (N_491,N_383,N_394);
or U492 (N_492,N_396,N_395);
and U493 (N_493,N_395,N_314);
and U494 (N_494,N_358,N_315);
nand U495 (N_495,N_354,N_345);
nand U496 (N_496,N_333,N_382);
nand U497 (N_497,N_318,N_355);
nand U498 (N_498,N_348,N_374);
or U499 (N_499,N_380,N_352);
nand U500 (N_500,N_447,N_425);
and U501 (N_501,N_492,N_408);
nor U502 (N_502,N_430,N_483);
or U503 (N_503,N_401,N_427);
and U504 (N_504,N_493,N_467);
nand U505 (N_505,N_404,N_458);
nand U506 (N_506,N_475,N_417);
nor U507 (N_507,N_451,N_484);
nand U508 (N_508,N_466,N_409);
and U509 (N_509,N_410,N_459);
nand U510 (N_510,N_428,N_464);
nand U511 (N_511,N_479,N_485);
xnor U512 (N_512,N_443,N_489);
nand U513 (N_513,N_446,N_480);
nor U514 (N_514,N_476,N_433);
and U515 (N_515,N_416,N_407);
nor U516 (N_516,N_461,N_495);
or U517 (N_517,N_400,N_405);
and U518 (N_518,N_486,N_435);
or U519 (N_519,N_403,N_444);
nand U520 (N_520,N_421,N_473);
and U521 (N_521,N_432,N_429);
nor U522 (N_522,N_497,N_437);
nor U523 (N_523,N_414,N_431);
or U524 (N_524,N_487,N_456);
nand U525 (N_525,N_415,N_445);
nand U526 (N_526,N_442,N_452);
or U527 (N_527,N_426,N_465);
nor U528 (N_528,N_406,N_482);
nand U529 (N_529,N_420,N_412);
nor U530 (N_530,N_468,N_453);
or U531 (N_531,N_424,N_494);
and U532 (N_532,N_499,N_474);
nor U533 (N_533,N_490,N_488);
or U534 (N_534,N_481,N_441);
nand U535 (N_535,N_440,N_454);
nor U536 (N_536,N_439,N_463);
nand U537 (N_537,N_457,N_472);
nor U538 (N_538,N_471,N_455);
and U539 (N_539,N_448,N_462);
or U540 (N_540,N_470,N_496);
or U541 (N_541,N_491,N_450);
nand U542 (N_542,N_469,N_498);
nor U543 (N_543,N_478,N_419);
nor U544 (N_544,N_460,N_418);
or U545 (N_545,N_402,N_422);
and U546 (N_546,N_411,N_436);
xnor U547 (N_547,N_438,N_449);
and U548 (N_548,N_413,N_423);
nand U549 (N_549,N_477,N_434);
or U550 (N_550,N_480,N_490);
nor U551 (N_551,N_481,N_490);
or U552 (N_552,N_423,N_467);
nand U553 (N_553,N_427,N_490);
nor U554 (N_554,N_493,N_413);
nand U555 (N_555,N_403,N_404);
nand U556 (N_556,N_437,N_479);
nand U557 (N_557,N_476,N_471);
nand U558 (N_558,N_478,N_430);
nand U559 (N_559,N_419,N_497);
nand U560 (N_560,N_472,N_430);
and U561 (N_561,N_456,N_471);
nand U562 (N_562,N_402,N_426);
nand U563 (N_563,N_419,N_470);
and U564 (N_564,N_407,N_437);
nand U565 (N_565,N_429,N_477);
nand U566 (N_566,N_455,N_419);
nor U567 (N_567,N_405,N_461);
nand U568 (N_568,N_478,N_405);
and U569 (N_569,N_455,N_417);
and U570 (N_570,N_427,N_489);
nand U571 (N_571,N_409,N_419);
nand U572 (N_572,N_470,N_427);
nor U573 (N_573,N_412,N_497);
nor U574 (N_574,N_469,N_439);
nor U575 (N_575,N_468,N_459);
and U576 (N_576,N_420,N_404);
and U577 (N_577,N_443,N_474);
nor U578 (N_578,N_405,N_462);
and U579 (N_579,N_475,N_496);
and U580 (N_580,N_408,N_481);
nand U581 (N_581,N_470,N_406);
and U582 (N_582,N_478,N_409);
and U583 (N_583,N_443,N_421);
nor U584 (N_584,N_488,N_429);
nor U585 (N_585,N_477,N_464);
or U586 (N_586,N_415,N_426);
and U587 (N_587,N_471,N_415);
or U588 (N_588,N_465,N_407);
xor U589 (N_589,N_432,N_453);
and U590 (N_590,N_441,N_461);
and U591 (N_591,N_415,N_400);
nand U592 (N_592,N_418,N_408);
nor U593 (N_593,N_488,N_443);
or U594 (N_594,N_408,N_404);
and U595 (N_595,N_491,N_478);
nand U596 (N_596,N_488,N_414);
nor U597 (N_597,N_424,N_464);
nand U598 (N_598,N_408,N_425);
nand U599 (N_599,N_470,N_416);
or U600 (N_600,N_521,N_573);
nand U601 (N_601,N_579,N_599);
or U602 (N_602,N_572,N_560);
and U603 (N_603,N_546,N_528);
or U604 (N_604,N_552,N_517);
and U605 (N_605,N_537,N_544);
nor U606 (N_606,N_509,N_501);
nor U607 (N_607,N_542,N_578);
nand U608 (N_608,N_590,N_567);
nor U609 (N_609,N_586,N_574);
nor U610 (N_610,N_536,N_562);
or U611 (N_611,N_504,N_502);
nor U612 (N_612,N_520,N_549);
or U613 (N_613,N_527,N_551);
and U614 (N_614,N_550,N_540);
and U615 (N_615,N_569,N_559);
and U616 (N_616,N_503,N_524);
and U617 (N_617,N_598,N_566);
or U618 (N_618,N_522,N_582);
and U619 (N_619,N_557,N_539);
or U620 (N_620,N_555,N_564);
and U621 (N_621,N_510,N_516);
or U622 (N_622,N_508,N_575);
nor U623 (N_623,N_543,N_583);
and U624 (N_624,N_532,N_512);
nor U625 (N_625,N_584,N_585);
nor U626 (N_626,N_577,N_556);
nor U627 (N_627,N_507,N_506);
nor U628 (N_628,N_526,N_513);
or U629 (N_629,N_519,N_591);
nand U630 (N_630,N_588,N_589);
nor U631 (N_631,N_545,N_580);
nand U632 (N_632,N_592,N_511);
nor U633 (N_633,N_505,N_596);
or U634 (N_634,N_563,N_525);
nor U635 (N_635,N_553,N_554);
and U636 (N_636,N_593,N_587);
or U637 (N_637,N_541,N_594);
and U638 (N_638,N_571,N_514);
and U639 (N_639,N_558,N_518);
nor U640 (N_640,N_534,N_500);
nor U641 (N_641,N_576,N_595);
nand U642 (N_642,N_568,N_565);
xnor U643 (N_643,N_570,N_529);
and U644 (N_644,N_515,N_548);
xor U645 (N_645,N_547,N_561);
and U646 (N_646,N_535,N_533);
and U647 (N_647,N_538,N_531);
or U648 (N_648,N_523,N_597);
and U649 (N_649,N_530,N_581);
nor U650 (N_650,N_507,N_538);
and U651 (N_651,N_568,N_538);
or U652 (N_652,N_515,N_570);
xor U653 (N_653,N_540,N_505);
nor U654 (N_654,N_530,N_592);
nand U655 (N_655,N_588,N_579);
or U656 (N_656,N_522,N_587);
nand U657 (N_657,N_510,N_544);
nand U658 (N_658,N_529,N_528);
nand U659 (N_659,N_581,N_562);
nor U660 (N_660,N_517,N_568);
and U661 (N_661,N_595,N_516);
or U662 (N_662,N_568,N_589);
nand U663 (N_663,N_562,N_595);
or U664 (N_664,N_503,N_572);
or U665 (N_665,N_559,N_521);
or U666 (N_666,N_561,N_510);
nor U667 (N_667,N_568,N_529);
nand U668 (N_668,N_548,N_582);
or U669 (N_669,N_583,N_549);
nand U670 (N_670,N_511,N_595);
nand U671 (N_671,N_539,N_533);
and U672 (N_672,N_579,N_568);
or U673 (N_673,N_583,N_534);
and U674 (N_674,N_506,N_550);
and U675 (N_675,N_508,N_569);
nand U676 (N_676,N_586,N_551);
nand U677 (N_677,N_525,N_541);
and U678 (N_678,N_549,N_510);
or U679 (N_679,N_564,N_546);
and U680 (N_680,N_516,N_557);
and U681 (N_681,N_540,N_519);
nand U682 (N_682,N_594,N_551);
xor U683 (N_683,N_542,N_573);
and U684 (N_684,N_529,N_541);
or U685 (N_685,N_529,N_518);
or U686 (N_686,N_501,N_567);
nand U687 (N_687,N_548,N_565);
nand U688 (N_688,N_504,N_535);
or U689 (N_689,N_582,N_578);
or U690 (N_690,N_526,N_581);
nand U691 (N_691,N_517,N_575);
and U692 (N_692,N_503,N_519);
nand U693 (N_693,N_554,N_586);
or U694 (N_694,N_595,N_578);
nand U695 (N_695,N_582,N_595);
nor U696 (N_696,N_598,N_567);
nor U697 (N_697,N_544,N_560);
nor U698 (N_698,N_521,N_579);
and U699 (N_699,N_565,N_586);
and U700 (N_700,N_607,N_668);
nor U701 (N_701,N_688,N_626);
nor U702 (N_702,N_658,N_686);
nand U703 (N_703,N_655,N_609);
or U704 (N_704,N_671,N_647);
or U705 (N_705,N_675,N_682);
or U706 (N_706,N_691,N_672);
xor U707 (N_707,N_602,N_615);
and U708 (N_708,N_627,N_618);
nor U709 (N_709,N_640,N_670);
and U710 (N_710,N_608,N_614);
or U711 (N_711,N_683,N_687);
nand U712 (N_712,N_645,N_689);
nor U713 (N_713,N_660,N_622);
nor U714 (N_714,N_659,N_657);
nor U715 (N_715,N_620,N_692);
or U716 (N_716,N_662,N_639);
and U717 (N_717,N_665,N_680);
nand U718 (N_718,N_695,N_616);
or U719 (N_719,N_603,N_648);
nand U720 (N_720,N_699,N_623);
xor U721 (N_721,N_690,N_651);
and U722 (N_722,N_697,N_600);
xor U723 (N_723,N_619,N_631);
or U724 (N_724,N_654,N_621);
or U725 (N_725,N_633,N_669);
nor U726 (N_726,N_638,N_666);
and U727 (N_727,N_643,N_642);
and U728 (N_728,N_641,N_653);
or U729 (N_729,N_628,N_629);
and U730 (N_730,N_696,N_661);
and U731 (N_731,N_674,N_612);
nor U732 (N_732,N_663,N_652);
nand U733 (N_733,N_637,N_636);
or U734 (N_734,N_625,N_644);
nand U735 (N_735,N_635,N_685);
nor U736 (N_736,N_634,N_656);
and U737 (N_737,N_677,N_646);
nor U738 (N_738,N_693,N_610);
and U739 (N_739,N_676,N_684);
or U740 (N_740,N_667,N_605);
and U741 (N_741,N_650,N_664);
nor U742 (N_742,N_698,N_604);
or U743 (N_743,N_673,N_630);
nor U744 (N_744,N_624,N_632);
nand U745 (N_745,N_601,N_611);
nand U746 (N_746,N_617,N_694);
nor U747 (N_747,N_681,N_679);
xnor U748 (N_748,N_606,N_678);
nor U749 (N_749,N_649,N_613);
nand U750 (N_750,N_649,N_672);
and U751 (N_751,N_601,N_688);
and U752 (N_752,N_649,N_667);
and U753 (N_753,N_627,N_625);
or U754 (N_754,N_662,N_623);
nand U755 (N_755,N_609,N_613);
and U756 (N_756,N_653,N_631);
nor U757 (N_757,N_623,N_626);
nor U758 (N_758,N_661,N_687);
or U759 (N_759,N_685,N_699);
nor U760 (N_760,N_612,N_671);
nand U761 (N_761,N_665,N_636);
and U762 (N_762,N_643,N_690);
or U763 (N_763,N_641,N_644);
nand U764 (N_764,N_622,N_638);
nor U765 (N_765,N_661,N_686);
or U766 (N_766,N_670,N_634);
nor U767 (N_767,N_600,N_618);
or U768 (N_768,N_643,N_602);
nor U769 (N_769,N_618,N_664);
or U770 (N_770,N_690,N_695);
nor U771 (N_771,N_685,N_633);
nand U772 (N_772,N_676,N_612);
xor U773 (N_773,N_657,N_658);
and U774 (N_774,N_654,N_696);
and U775 (N_775,N_645,N_675);
nand U776 (N_776,N_647,N_632);
and U777 (N_777,N_603,N_690);
or U778 (N_778,N_664,N_612);
xnor U779 (N_779,N_683,N_612);
or U780 (N_780,N_622,N_679);
xor U781 (N_781,N_606,N_683);
nor U782 (N_782,N_643,N_624);
nor U783 (N_783,N_675,N_616);
nor U784 (N_784,N_667,N_614);
nor U785 (N_785,N_677,N_687);
nand U786 (N_786,N_619,N_645);
nor U787 (N_787,N_611,N_669);
nor U788 (N_788,N_632,N_610);
nand U789 (N_789,N_637,N_659);
or U790 (N_790,N_601,N_663);
nand U791 (N_791,N_677,N_605);
or U792 (N_792,N_685,N_667);
nor U793 (N_793,N_662,N_615);
and U794 (N_794,N_617,N_652);
and U795 (N_795,N_620,N_607);
nor U796 (N_796,N_654,N_664);
and U797 (N_797,N_625,N_667);
and U798 (N_798,N_695,N_669);
nor U799 (N_799,N_671,N_652);
nor U800 (N_800,N_764,N_726);
nor U801 (N_801,N_718,N_735);
and U802 (N_802,N_774,N_736);
nand U803 (N_803,N_783,N_734);
nor U804 (N_804,N_730,N_766);
and U805 (N_805,N_779,N_784);
and U806 (N_806,N_714,N_741);
nand U807 (N_807,N_765,N_742);
and U808 (N_808,N_787,N_758);
or U809 (N_809,N_708,N_748);
or U810 (N_810,N_711,N_778);
nor U811 (N_811,N_793,N_712);
nand U812 (N_812,N_780,N_781);
and U813 (N_813,N_750,N_771);
nor U814 (N_814,N_706,N_775);
nor U815 (N_815,N_723,N_707);
nor U816 (N_816,N_786,N_744);
and U817 (N_817,N_739,N_770);
or U818 (N_818,N_769,N_761);
nor U819 (N_819,N_768,N_715);
and U820 (N_820,N_755,N_705);
nor U821 (N_821,N_760,N_738);
nor U822 (N_822,N_792,N_746);
xor U823 (N_823,N_731,N_751);
xnor U824 (N_824,N_782,N_700);
or U825 (N_825,N_767,N_756);
nor U826 (N_826,N_704,N_717);
or U827 (N_827,N_747,N_772);
nor U828 (N_828,N_776,N_789);
nand U829 (N_829,N_790,N_719);
nor U830 (N_830,N_724,N_722);
or U831 (N_831,N_713,N_791);
nand U832 (N_832,N_773,N_725);
nand U833 (N_833,N_710,N_729);
nor U834 (N_834,N_703,N_798);
nand U835 (N_835,N_796,N_752);
nand U836 (N_836,N_728,N_788);
xnor U837 (N_837,N_762,N_733);
nand U838 (N_838,N_777,N_732);
nor U839 (N_839,N_743,N_754);
nand U840 (N_840,N_749,N_795);
nand U841 (N_841,N_701,N_720);
nor U842 (N_842,N_727,N_709);
and U843 (N_843,N_745,N_797);
nor U844 (N_844,N_753,N_702);
or U845 (N_845,N_759,N_785);
nor U846 (N_846,N_737,N_716);
or U847 (N_847,N_721,N_757);
nor U848 (N_848,N_799,N_763);
nand U849 (N_849,N_794,N_740);
nand U850 (N_850,N_754,N_798);
nor U851 (N_851,N_740,N_769);
xor U852 (N_852,N_732,N_736);
or U853 (N_853,N_764,N_796);
xnor U854 (N_854,N_753,N_701);
and U855 (N_855,N_736,N_700);
nor U856 (N_856,N_724,N_770);
xnor U857 (N_857,N_782,N_706);
or U858 (N_858,N_767,N_717);
or U859 (N_859,N_795,N_794);
nand U860 (N_860,N_730,N_786);
or U861 (N_861,N_753,N_786);
or U862 (N_862,N_718,N_771);
nand U863 (N_863,N_778,N_726);
or U864 (N_864,N_770,N_781);
nor U865 (N_865,N_755,N_773);
and U866 (N_866,N_721,N_709);
nand U867 (N_867,N_786,N_775);
or U868 (N_868,N_717,N_787);
or U869 (N_869,N_769,N_759);
nand U870 (N_870,N_701,N_738);
nor U871 (N_871,N_771,N_793);
or U872 (N_872,N_756,N_772);
or U873 (N_873,N_775,N_768);
nor U874 (N_874,N_725,N_780);
and U875 (N_875,N_721,N_759);
nand U876 (N_876,N_735,N_752);
nor U877 (N_877,N_722,N_769);
nand U878 (N_878,N_790,N_776);
and U879 (N_879,N_794,N_743);
and U880 (N_880,N_755,N_793);
nor U881 (N_881,N_771,N_775);
nor U882 (N_882,N_798,N_719);
xnor U883 (N_883,N_752,N_791);
nor U884 (N_884,N_728,N_776);
xor U885 (N_885,N_748,N_795);
or U886 (N_886,N_759,N_736);
nand U887 (N_887,N_750,N_792);
nor U888 (N_888,N_751,N_798);
nor U889 (N_889,N_794,N_798);
and U890 (N_890,N_797,N_773);
nand U891 (N_891,N_773,N_700);
nor U892 (N_892,N_752,N_753);
nor U893 (N_893,N_774,N_756);
xnor U894 (N_894,N_714,N_777);
nand U895 (N_895,N_786,N_789);
and U896 (N_896,N_707,N_790);
and U897 (N_897,N_764,N_706);
or U898 (N_898,N_767,N_710);
or U899 (N_899,N_788,N_749);
and U900 (N_900,N_883,N_842);
nand U901 (N_901,N_805,N_815);
nand U902 (N_902,N_855,N_864);
or U903 (N_903,N_831,N_866);
or U904 (N_904,N_878,N_812);
nor U905 (N_905,N_847,N_894);
nor U906 (N_906,N_839,N_822);
nor U907 (N_907,N_868,N_862);
or U908 (N_908,N_859,N_882);
and U909 (N_909,N_845,N_818);
or U910 (N_910,N_844,N_816);
or U911 (N_911,N_891,N_806);
nor U912 (N_912,N_876,N_872);
nand U913 (N_913,N_879,N_838);
nand U914 (N_914,N_863,N_800);
and U915 (N_915,N_808,N_804);
nand U916 (N_916,N_858,N_821);
nor U917 (N_917,N_835,N_884);
and U918 (N_918,N_857,N_877);
and U919 (N_919,N_870,N_888);
nor U920 (N_920,N_825,N_819);
nand U921 (N_921,N_837,N_846);
or U922 (N_922,N_873,N_865);
and U923 (N_923,N_843,N_851);
and U924 (N_924,N_829,N_814);
nor U925 (N_925,N_820,N_898);
and U926 (N_926,N_890,N_871);
nor U927 (N_927,N_801,N_874);
and U928 (N_928,N_869,N_830);
or U929 (N_929,N_895,N_833);
and U930 (N_930,N_856,N_849);
and U931 (N_931,N_828,N_886);
and U932 (N_932,N_896,N_840);
nand U933 (N_933,N_824,N_897);
or U934 (N_934,N_880,N_826);
nor U935 (N_935,N_827,N_860);
or U936 (N_936,N_817,N_803);
nor U937 (N_937,N_850,N_807);
nor U938 (N_938,N_854,N_823);
nand U939 (N_939,N_809,N_875);
nand U940 (N_940,N_832,N_853);
or U941 (N_941,N_867,N_852);
nor U942 (N_942,N_885,N_836);
nor U943 (N_943,N_881,N_810);
nand U944 (N_944,N_892,N_811);
or U945 (N_945,N_834,N_887);
nand U946 (N_946,N_841,N_802);
nor U947 (N_947,N_861,N_893);
xnor U948 (N_948,N_889,N_899);
xor U949 (N_949,N_813,N_848);
nand U950 (N_950,N_854,N_815);
or U951 (N_951,N_831,N_886);
nand U952 (N_952,N_834,N_845);
and U953 (N_953,N_869,N_895);
or U954 (N_954,N_835,N_876);
nor U955 (N_955,N_861,N_833);
or U956 (N_956,N_874,N_899);
nor U957 (N_957,N_802,N_876);
or U958 (N_958,N_863,N_831);
and U959 (N_959,N_833,N_830);
nand U960 (N_960,N_827,N_868);
nor U961 (N_961,N_804,N_844);
nor U962 (N_962,N_861,N_896);
nand U963 (N_963,N_846,N_871);
and U964 (N_964,N_813,N_837);
and U965 (N_965,N_854,N_888);
nor U966 (N_966,N_823,N_870);
and U967 (N_967,N_828,N_829);
or U968 (N_968,N_812,N_804);
or U969 (N_969,N_891,N_846);
and U970 (N_970,N_876,N_869);
or U971 (N_971,N_824,N_842);
and U972 (N_972,N_810,N_840);
nand U973 (N_973,N_889,N_865);
nand U974 (N_974,N_875,N_827);
nor U975 (N_975,N_860,N_854);
nand U976 (N_976,N_826,N_817);
nor U977 (N_977,N_803,N_833);
nand U978 (N_978,N_867,N_893);
nor U979 (N_979,N_859,N_830);
nand U980 (N_980,N_890,N_876);
nor U981 (N_981,N_832,N_803);
or U982 (N_982,N_847,N_848);
nand U983 (N_983,N_852,N_837);
and U984 (N_984,N_869,N_819);
or U985 (N_985,N_883,N_820);
nor U986 (N_986,N_872,N_813);
nor U987 (N_987,N_862,N_838);
nor U988 (N_988,N_823,N_825);
nor U989 (N_989,N_811,N_814);
nor U990 (N_990,N_831,N_873);
nand U991 (N_991,N_889,N_887);
nand U992 (N_992,N_849,N_850);
nor U993 (N_993,N_823,N_830);
nand U994 (N_994,N_816,N_811);
and U995 (N_995,N_895,N_884);
and U996 (N_996,N_878,N_848);
nor U997 (N_997,N_825,N_800);
nand U998 (N_998,N_843,N_812);
nor U999 (N_999,N_822,N_898);
or U1000 (N_1000,N_919,N_903);
xor U1001 (N_1001,N_913,N_951);
and U1002 (N_1002,N_979,N_933);
nor U1003 (N_1003,N_943,N_937);
nor U1004 (N_1004,N_900,N_989);
or U1005 (N_1005,N_956,N_948);
or U1006 (N_1006,N_993,N_930);
nor U1007 (N_1007,N_983,N_910);
nor U1008 (N_1008,N_907,N_964);
nand U1009 (N_1009,N_942,N_908);
xor U1010 (N_1010,N_967,N_997);
or U1011 (N_1011,N_952,N_957);
and U1012 (N_1012,N_914,N_959);
or U1013 (N_1013,N_915,N_970);
nand U1014 (N_1014,N_985,N_986);
nor U1015 (N_1015,N_954,N_971);
or U1016 (N_1016,N_911,N_931);
or U1017 (N_1017,N_917,N_947);
nand U1018 (N_1018,N_955,N_998);
or U1019 (N_1019,N_977,N_901);
or U1020 (N_1020,N_984,N_934);
nor U1021 (N_1021,N_958,N_996);
or U1022 (N_1022,N_965,N_906);
nor U1023 (N_1023,N_995,N_999);
or U1024 (N_1024,N_963,N_973);
nor U1025 (N_1025,N_940,N_976);
and U1026 (N_1026,N_988,N_960);
xor U1027 (N_1027,N_981,N_992);
or U1028 (N_1028,N_990,N_962);
nand U1029 (N_1029,N_953,N_902);
or U1030 (N_1030,N_949,N_950);
xor U1031 (N_1031,N_924,N_923);
nand U1032 (N_1032,N_904,N_935);
and U1033 (N_1033,N_972,N_941);
or U1034 (N_1034,N_939,N_905);
or U1035 (N_1035,N_926,N_982);
nor U1036 (N_1036,N_987,N_968);
nor U1037 (N_1037,N_916,N_946);
and U1038 (N_1038,N_928,N_945);
nor U1039 (N_1039,N_944,N_925);
nand U1040 (N_1040,N_920,N_980);
nand U1041 (N_1041,N_932,N_974);
and U1042 (N_1042,N_975,N_921);
or U1043 (N_1043,N_994,N_922);
or U1044 (N_1044,N_909,N_938);
or U1045 (N_1045,N_927,N_918);
nor U1046 (N_1046,N_936,N_991);
nor U1047 (N_1047,N_969,N_961);
and U1048 (N_1048,N_912,N_966);
and U1049 (N_1049,N_929,N_978);
or U1050 (N_1050,N_996,N_955);
nand U1051 (N_1051,N_917,N_911);
xnor U1052 (N_1052,N_948,N_926);
nand U1053 (N_1053,N_999,N_943);
and U1054 (N_1054,N_965,N_969);
or U1055 (N_1055,N_928,N_927);
nand U1056 (N_1056,N_907,N_957);
and U1057 (N_1057,N_964,N_973);
and U1058 (N_1058,N_939,N_951);
and U1059 (N_1059,N_932,N_965);
nand U1060 (N_1060,N_977,N_967);
nor U1061 (N_1061,N_924,N_965);
nand U1062 (N_1062,N_947,N_948);
or U1063 (N_1063,N_911,N_932);
nor U1064 (N_1064,N_982,N_918);
and U1065 (N_1065,N_974,N_971);
nand U1066 (N_1066,N_930,N_904);
and U1067 (N_1067,N_987,N_917);
nand U1068 (N_1068,N_983,N_949);
or U1069 (N_1069,N_933,N_983);
and U1070 (N_1070,N_940,N_956);
or U1071 (N_1071,N_926,N_925);
and U1072 (N_1072,N_920,N_938);
and U1073 (N_1073,N_968,N_962);
nor U1074 (N_1074,N_958,N_927);
or U1075 (N_1075,N_968,N_989);
nand U1076 (N_1076,N_938,N_978);
nor U1077 (N_1077,N_973,N_904);
nor U1078 (N_1078,N_953,N_903);
nor U1079 (N_1079,N_918,N_920);
nor U1080 (N_1080,N_935,N_924);
nand U1081 (N_1081,N_984,N_944);
or U1082 (N_1082,N_908,N_904);
or U1083 (N_1083,N_962,N_907);
and U1084 (N_1084,N_906,N_917);
nand U1085 (N_1085,N_961,N_962);
nor U1086 (N_1086,N_981,N_931);
nor U1087 (N_1087,N_995,N_943);
nor U1088 (N_1088,N_965,N_997);
or U1089 (N_1089,N_982,N_908);
nand U1090 (N_1090,N_944,N_956);
or U1091 (N_1091,N_932,N_929);
xnor U1092 (N_1092,N_919,N_993);
nand U1093 (N_1093,N_915,N_907);
or U1094 (N_1094,N_975,N_943);
nor U1095 (N_1095,N_943,N_906);
and U1096 (N_1096,N_922,N_997);
and U1097 (N_1097,N_951,N_941);
nor U1098 (N_1098,N_923,N_925);
nor U1099 (N_1099,N_918,N_995);
or U1100 (N_1100,N_1087,N_1061);
and U1101 (N_1101,N_1012,N_1066);
or U1102 (N_1102,N_1045,N_1060);
or U1103 (N_1103,N_1064,N_1023);
nand U1104 (N_1104,N_1067,N_1038);
or U1105 (N_1105,N_1036,N_1089);
nor U1106 (N_1106,N_1051,N_1028);
and U1107 (N_1107,N_1072,N_1080);
nor U1108 (N_1108,N_1070,N_1011);
nor U1109 (N_1109,N_1069,N_1027);
or U1110 (N_1110,N_1058,N_1004);
and U1111 (N_1111,N_1056,N_1007);
or U1112 (N_1112,N_1016,N_1014);
nand U1113 (N_1113,N_1044,N_1026);
nor U1114 (N_1114,N_1030,N_1017);
or U1115 (N_1115,N_1094,N_1034);
and U1116 (N_1116,N_1062,N_1029);
nor U1117 (N_1117,N_1009,N_1090);
or U1118 (N_1118,N_1092,N_1093);
or U1119 (N_1119,N_1097,N_1019);
and U1120 (N_1120,N_1033,N_1039);
or U1121 (N_1121,N_1075,N_1071);
nor U1122 (N_1122,N_1001,N_1046);
and U1123 (N_1123,N_1088,N_1025);
and U1124 (N_1124,N_1037,N_1013);
or U1125 (N_1125,N_1096,N_1077);
nor U1126 (N_1126,N_1018,N_1055);
or U1127 (N_1127,N_1057,N_1086);
xnor U1128 (N_1128,N_1020,N_1043);
and U1129 (N_1129,N_1078,N_1091);
and U1130 (N_1130,N_1052,N_1054);
nand U1131 (N_1131,N_1059,N_1015);
and U1132 (N_1132,N_1063,N_1047);
or U1133 (N_1133,N_1098,N_1000);
nand U1134 (N_1134,N_1048,N_1003);
and U1135 (N_1135,N_1081,N_1006);
xnor U1136 (N_1136,N_1010,N_1022);
and U1137 (N_1137,N_1042,N_1074);
nor U1138 (N_1138,N_1035,N_1002);
or U1139 (N_1139,N_1041,N_1076);
nor U1140 (N_1140,N_1049,N_1053);
and U1141 (N_1141,N_1099,N_1040);
and U1142 (N_1142,N_1050,N_1095);
xnor U1143 (N_1143,N_1082,N_1021);
nor U1144 (N_1144,N_1079,N_1031);
and U1145 (N_1145,N_1073,N_1065);
nor U1146 (N_1146,N_1024,N_1032);
nor U1147 (N_1147,N_1084,N_1068);
xnor U1148 (N_1148,N_1005,N_1083);
nand U1149 (N_1149,N_1085,N_1008);
or U1150 (N_1150,N_1026,N_1041);
and U1151 (N_1151,N_1017,N_1022);
or U1152 (N_1152,N_1030,N_1016);
and U1153 (N_1153,N_1034,N_1073);
nand U1154 (N_1154,N_1035,N_1037);
nand U1155 (N_1155,N_1069,N_1097);
or U1156 (N_1156,N_1017,N_1099);
nand U1157 (N_1157,N_1037,N_1048);
nand U1158 (N_1158,N_1016,N_1005);
nor U1159 (N_1159,N_1070,N_1068);
nor U1160 (N_1160,N_1001,N_1037);
and U1161 (N_1161,N_1061,N_1051);
or U1162 (N_1162,N_1091,N_1088);
and U1163 (N_1163,N_1053,N_1067);
nand U1164 (N_1164,N_1039,N_1051);
or U1165 (N_1165,N_1006,N_1011);
nand U1166 (N_1166,N_1042,N_1057);
nand U1167 (N_1167,N_1040,N_1023);
nand U1168 (N_1168,N_1093,N_1067);
nor U1169 (N_1169,N_1089,N_1091);
and U1170 (N_1170,N_1017,N_1061);
nand U1171 (N_1171,N_1013,N_1051);
or U1172 (N_1172,N_1065,N_1093);
xor U1173 (N_1173,N_1080,N_1006);
and U1174 (N_1174,N_1050,N_1091);
nand U1175 (N_1175,N_1075,N_1038);
and U1176 (N_1176,N_1083,N_1089);
and U1177 (N_1177,N_1049,N_1039);
and U1178 (N_1178,N_1099,N_1059);
or U1179 (N_1179,N_1038,N_1000);
or U1180 (N_1180,N_1050,N_1042);
and U1181 (N_1181,N_1064,N_1006);
nor U1182 (N_1182,N_1031,N_1029);
or U1183 (N_1183,N_1088,N_1051);
and U1184 (N_1184,N_1010,N_1004);
or U1185 (N_1185,N_1062,N_1013);
nand U1186 (N_1186,N_1024,N_1078);
nand U1187 (N_1187,N_1059,N_1087);
or U1188 (N_1188,N_1082,N_1070);
nand U1189 (N_1189,N_1084,N_1028);
nand U1190 (N_1190,N_1039,N_1095);
and U1191 (N_1191,N_1072,N_1004);
nand U1192 (N_1192,N_1027,N_1058);
nor U1193 (N_1193,N_1051,N_1003);
nor U1194 (N_1194,N_1057,N_1031);
or U1195 (N_1195,N_1028,N_1069);
and U1196 (N_1196,N_1052,N_1031);
and U1197 (N_1197,N_1000,N_1025);
and U1198 (N_1198,N_1065,N_1045);
nor U1199 (N_1199,N_1095,N_1004);
nand U1200 (N_1200,N_1168,N_1138);
and U1201 (N_1201,N_1106,N_1170);
and U1202 (N_1202,N_1150,N_1148);
and U1203 (N_1203,N_1118,N_1136);
nand U1204 (N_1204,N_1173,N_1145);
nand U1205 (N_1205,N_1182,N_1177);
nor U1206 (N_1206,N_1153,N_1104);
nand U1207 (N_1207,N_1166,N_1193);
or U1208 (N_1208,N_1142,N_1101);
nand U1209 (N_1209,N_1163,N_1107);
nand U1210 (N_1210,N_1188,N_1144);
nor U1211 (N_1211,N_1149,N_1161);
or U1212 (N_1212,N_1151,N_1176);
nor U1213 (N_1213,N_1195,N_1115);
nand U1214 (N_1214,N_1121,N_1156);
and U1215 (N_1215,N_1105,N_1184);
or U1216 (N_1216,N_1146,N_1190);
or U1217 (N_1217,N_1102,N_1183);
xor U1218 (N_1218,N_1127,N_1172);
nor U1219 (N_1219,N_1162,N_1179);
and U1220 (N_1220,N_1171,N_1152);
nor U1221 (N_1221,N_1160,N_1111);
and U1222 (N_1222,N_1180,N_1119);
nor U1223 (N_1223,N_1181,N_1100);
and U1224 (N_1224,N_1120,N_1174);
nor U1225 (N_1225,N_1122,N_1187);
and U1226 (N_1226,N_1141,N_1155);
or U1227 (N_1227,N_1169,N_1124);
and U1228 (N_1228,N_1129,N_1189);
and U1229 (N_1229,N_1194,N_1157);
nand U1230 (N_1230,N_1139,N_1192);
nor U1231 (N_1231,N_1164,N_1114);
nor U1232 (N_1232,N_1191,N_1199);
nand U1233 (N_1233,N_1178,N_1113);
or U1234 (N_1234,N_1110,N_1137);
and U1235 (N_1235,N_1165,N_1159);
nor U1236 (N_1236,N_1103,N_1140);
nor U1237 (N_1237,N_1131,N_1135);
xnor U1238 (N_1238,N_1109,N_1147);
nand U1239 (N_1239,N_1112,N_1154);
nor U1240 (N_1240,N_1158,N_1117);
nor U1241 (N_1241,N_1143,N_1186);
nand U1242 (N_1242,N_1132,N_1198);
nand U1243 (N_1243,N_1123,N_1196);
xnor U1244 (N_1244,N_1125,N_1116);
nand U1245 (N_1245,N_1133,N_1134);
and U1246 (N_1246,N_1185,N_1130);
nand U1247 (N_1247,N_1167,N_1197);
nor U1248 (N_1248,N_1175,N_1126);
nor U1249 (N_1249,N_1128,N_1108);
nand U1250 (N_1250,N_1135,N_1156);
nor U1251 (N_1251,N_1160,N_1179);
or U1252 (N_1252,N_1127,N_1160);
nand U1253 (N_1253,N_1175,N_1112);
and U1254 (N_1254,N_1158,N_1164);
nand U1255 (N_1255,N_1158,N_1146);
or U1256 (N_1256,N_1171,N_1158);
nand U1257 (N_1257,N_1109,N_1139);
nor U1258 (N_1258,N_1154,N_1166);
and U1259 (N_1259,N_1111,N_1148);
or U1260 (N_1260,N_1190,N_1136);
and U1261 (N_1261,N_1194,N_1145);
nand U1262 (N_1262,N_1110,N_1178);
or U1263 (N_1263,N_1154,N_1187);
and U1264 (N_1264,N_1134,N_1188);
nand U1265 (N_1265,N_1103,N_1167);
and U1266 (N_1266,N_1152,N_1123);
and U1267 (N_1267,N_1195,N_1162);
or U1268 (N_1268,N_1149,N_1101);
xor U1269 (N_1269,N_1186,N_1199);
nand U1270 (N_1270,N_1155,N_1145);
nor U1271 (N_1271,N_1117,N_1168);
or U1272 (N_1272,N_1171,N_1160);
nor U1273 (N_1273,N_1163,N_1168);
and U1274 (N_1274,N_1171,N_1119);
and U1275 (N_1275,N_1156,N_1198);
nand U1276 (N_1276,N_1161,N_1118);
and U1277 (N_1277,N_1111,N_1151);
nor U1278 (N_1278,N_1158,N_1159);
and U1279 (N_1279,N_1131,N_1181);
nand U1280 (N_1280,N_1133,N_1156);
or U1281 (N_1281,N_1171,N_1115);
or U1282 (N_1282,N_1171,N_1108);
nor U1283 (N_1283,N_1191,N_1139);
or U1284 (N_1284,N_1162,N_1175);
nand U1285 (N_1285,N_1112,N_1113);
or U1286 (N_1286,N_1108,N_1188);
and U1287 (N_1287,N_1110,N_1179);
and U1288 (N_1288,N_1185,N_1184);
or U1289 (N_1289,N_1133,N_1109);
nor U1290 (N_1290,N_1118,N_1102);
nand U1291 (N_1291,N_1112,N_1148);
nand U1292 (N_1292,N_1157,N_1155);
and U1293 (N_1293,N_1155,N_1129);
and U1294 (N_1294,N_1191,N_1159);
nor U1295 (N_1295,N_1191,N_1162);
nor U1296 (N_1296,N_1195,N_1198);
and U1297 (N_1297,N_1114,N_1144);
or U1298 (N_1298,N_1101,N_1118);
and U1299 (N_1299,N_1181,N_1107);
nand U1300 (N_1300,N_1253,N_1236);
nand U1301 (N_1301,N_1245,N_1203);
nor U1302 (N_1302,N_1262,N_1246);
or U1303 (N_1303,N_1277,N_1211);
nand U1304 (N_1304,N_1256,N_1249);
nand U1305 (N_1305,N_1289,N_1267);
nor U1306 (N_1306,N_1264,N_1284);
nor U1307 (N_1307,N_1271,N_1263);
xnor U1308 (N_1308,N_1234,N_1280);
nor U1309 (N_1309,N_1270,N_1272);
nand U1310 (N_1310,N_1298,N_1227);
or U1311 (N_1311,N_1202,N_1220);
nand U1312 (N_1312,N_1299,N_1215);
xor U1313 (N_1313,N_1250,N_1226);
nor U1314 (N_1314,N_1231,N_1240);
or U1315 (N_1315,N_1200,N_1286);
nand U1316 (N_1316,N_1241,N_1257);
nand U1317 (N_1317,N_1291,N_1237);
or U1318 (N_1318,N_1293,N_1212);
or U1319 (N_1319,N_1239,N_1279);
nor U1320 (N_1320,N_1274,N_1260);
nand U1321 (N_1321,N_1209,N_1248);
nand U1322 (N_1322,N_1295,N_1254);
nand U1323 (N_1323,N_1214,N_1204);
xnor U1324 (N_1324,N_1252,N_1208);
and U1325 (N_1325,N_1297,N_1210);
nand U1326 (N_1326,N_1218,N_1285);
and U1327 (N_1327,N_1233,N_1219);
nand U1328 (N_1328,N_1281,N_1261);
nor U1329 (N_1329,N_1213,N_1242);
or U1330 (N_1330,N_1276,N_1223);
and U1331 (N_1331,N_1258,N_1221);
xnor U1332 (N_1332,N_1216,N_1290);
nor U1333 (N_1333,N_1259,N_1296);
and U1334 (N_1334,N_1275,N_1228);
nand U1335 (N_1335,N_1225,N_1201);
nand U1336 (N_1336,N_1232,N_1243);
nand U1337 (N_1337,N_1269,N_1222);
or U1338 (N_1338,N_1282,N_1265);
and U1339 (N_1339,N_1224,N_1251);
or U1340 (N_1340,N_1230,N_1294);
and U1341 (N_1341,N_1206,N_1235);
and U1342 (N_1342,N_1247,N_1238);
nor U1343 (N_1343,N_1229,N_1255);
and U1344 (N_1344,N_1283,N_1287);
nand U1345 (N_1345,N_1244,N_1268);
nand U1346 (N_1346,N_1266,N_1217);
or U1347 (N_1347,N_1205,N_1278);
or U1348 (N_1348,N_1207,N_1292);
nand U1349 (N_1349,N_1273,N_1288);
or U1350 (N_1350,N_1295,N_1217);
or U1351 (N_1351,N_1258,N_1204);
and U1352 (N_1352,N_1210,N_1239);
and U1353 (N_1353,N_1279,N_1256);
nand U1354 (N_1354,N_1282,N_1280);
or U1355 (N_1355,N_1204,N_1292);
nor U1356 (N_1356,N_1282,N_1234);
and U1357 (N_1357,N_1242,N_1232);
or U1358 (N_1358,N_1243,N_1291);
or U1359 (N_1359,N_1224,N_1220);
nand U1360 (N_1360,N_1295,N_1206);
or U1361 (N_1361,N_1240,N_1295);
nand U1362 (N_1362,N_1251,N_1218);
nor U1363 (N_1363,N_1294,N_1291);
nor U1364 (N_1364,N_1207,N_1253);
or U1365 (N_1365,N_1202,N_1257);
nand U1366 (N_1366,N_1283,N_1214);
or U1367 (N_1367,N_1297,N_1208);
nor U1368 (N_1368,N_1264,N_1269);
xnor U1369 (N_1369,N_1236,N_1214);
nor U1370 (N_1370,N_1201,N_1259);
and U1371 (N_1371,N_1257,N_1221);
or U1372 (N_1372,N_1299,N_1246);
nor U1373 (N_1373,N_1289,N_1256);
or U1374 (N_1374,N_1205,N_1218);
nor U1375 (N_1375,N_1243,N_1279);
and U1376 (N_1376,N_1215,N_1216);
nand U1377 (N_1377,N_1295,N_1255);
nand U1378 (N_1378,N_1212,N_1222);
and U1379 (N_1379,N_1290,N_1247);
nand U1380 (N_1380,N_1290,N_1275);
or U1381 (N_1381,N_1201,N_1242);
nand U1382 (N_1382,N_1250,N_1256);
xnor U1383 (N_1383,N_1239,N_1263);
nand U1384 (N_1384,N_1218,N_1223);
nand U1385 (N_1385,N_1226,N_1263);
or U1386 (N_1386,N_1200,N_1276);
nand U1387 (N_1387,N_1260,N_1291);
and U1388 (N_1388,N_1233,N_1231);
nand U1389 (N_1389,N_1225,N_1211);
nand U1390 (N_1390,N_1261,N_1275);
or U1391 (N_1391,N_1241,N_1231);
or U1392 (N_1392,N_1233,N_1239);
and U1393 (N_1393,N_1295,N_1266);
or U1394 (N_1394,N_1281,N_1248);
nor U1395 (N_1395,N_1261,N_1233);
nor U1396 (N_1396,N_1281,N_1283);
and U1397 (N_1397,N_1225,N_1258);
nand U1398 (N_1398,N_1240,N_1204);
or U1399 (N_1399,N_1294,N_1265);
nand U1400 (N_1400,N_1323,N_1347);
nand U1401 (N_1401,N_1300,N_1328);
and U1402 (N_1402,N_1359,N_1365);
nor U1403 (N_1403,N_1302,N_1397);
nor U1404 (N_1404,N_1316,N_1393);
nand U1405 (N_1405,N_1353,N_1398);
or U1406 (N_1406,N_1392,N_1321);
and U1407 (N_1407,N_1379,N_1334);
and U1408 (N_1408,N_1336,N_1335);
and U1409 (N_1409,N_1363,N_1345);
nor U1410 (N_1410,N_1331,N_1317);
or U1411 (N_1411,N_1343,N_1367);
and U1412 (N_1412,N_1304,N_1320);
xnor U1413 (N_1413,N_1309,N_1346);
nand U1414 (N_1414,N_1352,N_1387);
nor U1415 (N_1415,N_1313,N_1314);
nor U1416 (N_1416,N_1389,N_1356);
nand U1417 (N_1417,N_1325,N_1342);
or U1418 (N_1418,N_1383,N_1370);
nand U1419 (N_1419,N_1394,N_1322);
nor U1420 (N_1420,N_1382,N_1315);
xnor U1421 (N_1421,N_1327,N_1376);
and U1422 (N_1422,N_1337,N_1357);
nor U1423 (N_1423,N_1354,N_1339);
nor U1424 (N_1424,N_1366,N_1360);
nor U1425 (N_1425,N_1318,N_1332);
and U1426 (N_1426,N_1390,N_1388);
nand U1427 (N_1427,N_1396,N_1306);
nor U1428 (N_1428,N_1324,N_1329);
nor U1429 (N_1429,N_1377,N_1319);
or U1430 (N_1430,N_1348,N_1364);
or U1431 (N_1431,N_1311,N_1395);
and U1432 (N_1432,N_1384,N_1307);
and U1433 (N_1433,N_1330,N_1399);
nor U1434 (N_1434,N_1373,N_1312);
nor U1435 (N_1435,N_1326,N_1310);
or U1436 (N_1436,N_1391,N_1351);
and U1437 (N_1437,N_1308,N_1372);
nand U1438 (N_1438,N_1369,N_1378);
and U1439 (N_1439,N_1375,N_1386);
or U1440 (N_1440,N_1362,N_1301);
nand U1441 (N_1441,N_1385,N_1350);
or U1442 (N_1442,N_1303,N_1358);
or U1443 (N_1443,N_1380,N_1381);
nor U1444 (N_1444,N_1338,N_1340);
and U1445 (N_1445,N_1368,N_1349);
nor U1446 (N_1446,N_1371,N_1355);
nand U1447 (N_1447,N_1344,N_1361);
and U1448 (N_1448,N_1374,N_1341);
nor U1449 (N_1449,N_1305,N_1333);
nor U1450 (N_1450,N_1371,N_1349);
nand U1451 (N_1451,N_1362,N_1313);
or U1452 (N_1452,N_1376,N_1358);
nor U1453 (N_1453,N_1308,N_1377);
and U1454 (N_1454,N_1324,N_1377);
and U1455 (N_1455,N_1373,N_1357);
nor U1456 (N_1456,N_1399,N_1303);
nor U1457 (N_1457,N_1315,N_1384);
and U1458 (N_1458,N_1303,N_1345);
xor U1459 (N_1459,N_1322,N_1314);
nor U1460 (N_1460,N_1395,N_1348);
nor U1461 (N_1461,N_1351,N_1390);
nor U1462 (N_1462,N_1315,N_1357);
nand U1463 (N_1463,N_1384,N_1342);
or U1464 (N_1464,N_1305,N_1309);
and U1465 (N_1465,N_1316,N_1345);
or U1466 (N_1466,N_1394,N_1309);
or U1467 (N_1467,N_1352,N_1385);
or U1468 (N_1468,N_1391,N_1396);
or U1469 (N_1469,N_1332,N_1313);
nand U1470 (N_1470,N_1317,N_1327);
and U1471 (N_1471,N_1323,N_1328);
nand U1472 (N_1472,N_1351,N_1350);
nor U1473 (N_1473,N_1359,N_1301);
and U1474 (N_1474,N_1356,N_1305);
nand U1475 (N_1475,N_1349,N_1307);
nor U1476 (N_1476,N_1367,N_1360);
nand U1477 (N_1477,N_1390,N_1315);
or U1478 (N_1478,N_1316,N_1350);
nor U1479 (N_1479,N_1327,N_1379);
nor U1480 (N_1480,N_1396,N_1332);
or U1481 (N_1481,N_1380,N_1366);
and U1482 (N_1482,N_1302,N_1310);
or U1483 (N_1483,N_1396,N_1374);
nand U1484 (N_1484,N_1316,N_1372);
nand U1485 (N_1485,N_1365,N_1380);
or U1486 (N_1486,N_1343,N_1301);
and U1487 (N_1487,N_1390,N_1363);
nand U1488 (N_1488,N_1333,N_1307);
and U1489 (N_1489,N_1386,N_1389);
or U1490 (N_1490,N_1317,N_1347);
and U1491 (N_1491,N_1352,N_1303);
nand U1492 (N_1492,N_1364,N_1357);
nor U1493 (N_1493,N_1390,N_1337);
nand U1494 (N_1494,N_1306,N_1354);
nand U1495 (N_1495,N_1385,N_1390);
or U1496 (N_1496,N_1328,N_1308);
nor U1497 (N_1497,N_1369,N_1328);
or U1498 (N_1498,N_1387,N_1381);
nand U1499 (N_1499,N_1371,N_1359);
and U1500 (N_1500,N_1452,N_1436);
nor U1501 (N_1501,N_1475,N_1400);
nor U1502 (N_1502,N_1431,N_1435);
and U1503 (N_1503,N_1447,N_1428);
nor U1504 (N_1504,N_1404,N_1403);
nand U1505 (N_1505,N_1408,N_1429);
nor U1506 (N_1506,N_1486,N_1454);
and U1507 (N_1507,N_1450,N_1425);
or U1508 (N_1508,N_1409,N_1451);
and U1509 (N_1509,N_1488,N_1439);
and U1510 (N_1510,N_1410,N_1418);
and U1511 (N_1511,N_1459,N_1477);
and U1512 (N_1512,N_1494,N_1487);
and U1513 (N_1513,N_1497,N_1442);
or U1514 (N_1514,N_1446,N_1405);
nand U1515 (N_1515,N_1498,N_1419);
nand U1516 (N_1516,N_1402,N_1417);
and U1517 (N_1517,N_1413,N_1443);
or U1518 (N_1518,N_1481,N_1423);
or U1519 (N_1519,N_1476,N_1479);
nand U1520 (N_1520,N_1463,N_1427);
nor U1521 (N_1521,N_1466,N_1483);
and U1522 (N_1522,N_1482,N_1438);
nor U1523 (N_1523,N_1440,N_1480);
nand U1524 (N_1524,N_1467,N_1401);
nor U1525 (N_1525,N_1422,N_1414);
nor U1526 (N_1526,N_1407,N_1415);
or U1527 (N_1527,N_1471,N_1445);
or U1528 (N_1528,N_1426,N_1411);
or U1529 (N_1529,N_1468,N_1434);
or U1530 (N_1530,N_1473,N_1478);
nand U1531 (N_1531,N_1484,N_1461);
nand U1532 (N_1532,N_1455,N_1424);
or U1533 (N_1533,N_1491,N_1495);
or U1534 (N_1534,N_1465,N_1412);
or U1535 (N_1535,N_1456,N_1460);
nand U1536 (N_1536,N_1464,N_1421);
or U1537 (N_1537,N_1499,N_1485);
and U1538 (N_1538,N_1420,N_1493);
or U1539 (N_1539,N_1490,N_1453);
and U1540 (N_1540,N_1469,N_1457);
and U1541 (N_1541,N_1492,N_1472);
nor U1542 (N_1542,N_1448,N_1449);
nand U1543 (N_1543,N_1437,N_1406);
and U1544 (N_1544,N_1474,N_1458);
nand U1545 (N_1545,N_1416,N_1496);
nand U1546 (N_1546,N_1433,N_1462);
and U1547 (N_1547,N_1430,N_1444);
or U1548 (N_1548,N_1441,N_1432);
nor U1549 (N_1549,N_1489,N_1470);
and U1550 (N_1550,N_1451,N_1459);
nand U1551 (N_1551,N_1476,N_1454);
and U1552 (N_1552,N_1472,N_1444);
or U1553 (N_1553,N_1404,N_1469);
nand U1554 (N_1554,N_1420,N_1471);
and U1555 (N_1555,N_1494,N_1484);
nor U1556 (N_1556,N_1472,N_1441);
xor U1557 (N_1557,N_1404,N_1482);
nand U1558 (N_1558,N_1437,N_1470);
nand U1559 (N_1559,N_1403,N_1437);
nand U1560 (N_1560,N_1412,N_1415);
nor U1561 (N_1561,N_1469,N_1413);
nor U1562 (N_1562,N_1478,N_1463);
nand U1563 (N_1563,N_1497,N_1405);
nor U1564 (N_1564,N_1495,N_1437);
or U1565 (N_1565,N_1423,N_1480);
or U1566 (N_1566,N_1476,N_1427);
or U1567 (N_1567,N_1490,N_1455);
and U1568 (N_1568,N_1419,N_1488);
nor U1569 (N_1569,N_1492,N_1475);
or U1570 (N_1570,N_1424,N_1437);
nand U1571 (N_1571,N_1489,N_1436);
and U1572 (N_1572,N_1411,N_1498);
nor U1573 (N_1573,N_1426,N_1413);
nor U1574 (N_1574,N_1457,N_1498);
nand U1575 (N_1575,N_1462,N_1477);
xor U1576 (N_1576,N_1442,N_1454);
nand U1577 (N_1577,N_1456,N_1471);
or U1578 (N_1578,N_1441,N_1455);
or U1579 (N_1579,N_1412,N_1456);
and U1580 (N_1580,N_1484,N_1497);
and U1581 (N_1581,N_1468,N_1449);
or U1582 (N_1582,N_1465,N_1439);
and U1583 (N_1583,N_1492,N_1479);
nand U1584 (N_1584,N_1489,N_1455);
and U1585 (N_1585,N_1479,N_1429);
nor U1586 (N_1586,N_1447,N_1418);
nor U1587 (N_1587,N_1407,N_1448);
nand U1588 (N_1588,N_1465,N_1483);
nor U1589 (N_1589,N_1430,N_1409);
nor U1590 (N_1590,N_1479,N_1419);
and U1591 (N_1591,N_1447,N_1488);
nand U1592 (N_1592,N_1470,N_1450);
and U1593 (N_1593,N_1445,N_1475);
and U1594 (N_1594,N_1452,N_1432);
nor U1595 (N_1595,N_1496,N_1489);
or U1596 (N_1596,N_1454,N_1431);
or U1597 (N_1597,N_1473,N_1488);
nand U1598 (N_1598,N_1421,N_1403);
nor U1599 (N_1599,N_1467,N_1408);
nor U1600 (N_1600,N_1507,N_1599);
nand U1601 (N_1601,N_1526,N_1545);
or U1602 (N_1602,N_1565,N_1589);
and U1603 (N_1603,N_1559,N_1591);
nand U1604 (N_1604,N_1557,N_1514);
nand U1605 (N_1605,N_1536,N_1580);
or U1606 (N_1606,N_1571,N_1590);
or U1607 (N_1607,N_1511,N_1517);
or U1608 (N_1608,N_1518,N_1544);
nand U1609 (N_1609,N_1563,N_1584);
and U1610 (N_1610,N_1572,N_1504);
nand U1611 (N_1611,N_1510,N_1564);
nor U1612 (N_1612,N_1566,N_1596);
nand U1613 (N_1613,N_1529,N_1512);
and U1614 (N_1614,N_1534,N_1549);
or U1615 (N_1615,N_1509,N_1508);
nand U1616 (N_1616,N_1528,N_1521);
nand U1617 (N_1617,N_1522,N_1525);
and U1618 (N_1618,N_1516,N_1502);
and U1619 (N_1619,N_1593,N_1515);
nand U1620 (N_1620,N_1531,N_1538);
and U1621 (N_1621,N_1547,N_1527);
or U1622 (N_1622,N_1576,N_1595);
nor U1623 (N_1623,N_1583,N_1500);
nor U1624 (N_1624,N_1598,N_1524);
and U1625 (N_1625,N_1588,N_1585);
and U1626 (N_1626,N_1586,N_1573);
and U1627 (N_1627,N_1579,N_1555);
or U1628 (N_1628,N_1537,N_1597);
and U1629 (N_1629,N_1561,N_1570);
nand U1630 (N_1630,N_1581,N_1505);
nor U1631 (N_1631,N_1501,N_1578);
and U1632 (N_1632,N_1554,N_1587);
nor U1633 (N_1633,N_1520,N_1506);
or U1634 (N_1634,N_1562,N_1556);
nor U1635 (N_1635,N_1551,N_1574);
nand U1636 (N_1636,N_1543,N_1513);
and U1637 (N_1637,N_1575,N_1519);
nor U1638 (N_1638,N_1541,N_1503);
and U1639 (N_1639,N_1582,N_1568);
or U1640 (N_1640,N_1535,N_1532);
xor U1641 (N_1641,N_1550,N_1567);
or U1642 (N_1642,N_1523,N_1569);
nand U1643 (N_1643,N_1594,N_1546);
nor U1644 (N_1644,N_1539,N_1577);
and U1645 (N_1645,N_1592,N_1530);
nand U1646 (N_1646,N_1542,N_1548);
nor U1647 (N_1647,N_1540,N_1553);
and U1648 (N_1648,N_1558,N_1552);
and U1649 (N_1649,N_1533,N_1560);
and U1650 (N_1650,N_1501,N_1537);
and U1651 (N_1651,N_1503,N_1564);
nand U1652 (N_1652,N_1553,N_1558);
nor U1653 (N_1653,N_1571,N_1547);
xnor U1654 (N_1654,N_1538,N_1530);
or U1655 (N_1655,N_1548,N_1512);
or U1656 (N_1656,N_1570,N_1567);
nand U1657 (N_1657,N_1554,N_1562);
nand U1658 (N_1658,N_1507,N_1508);
and U1659 (N_1659,N_1533,N_1500);
nand U1660 (N_1660,N_1549,N_1595);
or U1661 (N_1661,N_1577,N_1523);
nand U1662 (N_1662,N_1562,N_1584);
and U1663 (N_1663,N_1557,N_1587);
nor U1664 (N_1664,N_1546,N_1510);
nand U1665 (N_1665,N_1500,N_1535);
nor U1666 (N_1666,N_1503,N_1547);
or U1667 (N_1667,N_1595,N_1523);
nor U1668 (N_1668,N_1560,N_1592);
or U1669 (N_1669,N_1535,N_1527);
and U1670 (N_1670,N_1572,N_1507);
and U1671 (N_1671,N_1521,N_1501);
and U1672 (N_1672,N_1596,N_1594);
nand U1673 (N_1673,N_1501,N_1516);
or U1674 (N_1674,N_1525,N_1517);
and U1675 (N_1675,N_1507,N_1534);
nand U1676 (N_1676,N_1590,N_1518);
and U1677 (N_1677,N_1536,N_1549);
and U1678 (N_1678,N_1594,N_1585);
and U1679 (N_1679,N_1559,N_1589);
or U1680 (N_1680,N_1538,N_1501);
and U1681 (N_1681,N_1529,N_1539);
or U1682 (N_1682,N_1508,N_1598);
and U1683 (N_1683,N_1500,N_1576);
nand U1684 (N_1684,N_1527,N_1591);
nand U1685 (N_1685,N_1551,N_1546);
or U1686 (N_1686,N_1507,N_1527);
and U1687 (N_1687,N_1535,N_1561);
or U1688 (N_1688,N_1544,N_1539);
nand U1689 (N_1689,N_1506,N_1529);
nand U1690 (N_1690,N_1522,N_1576);
or U1691 (N_1691,N_1518,N_1538);
nor U1692 (N_1692,N_1543,N_1502);
and U1693 (N_1693,N_1593,N_1508);
and U1694 (N_1694,N_1579,N_1548);
nand U1695 (N_1695,N_1536,N_1512);
and U1696 (N_1696,N_1509,N_1565);
and U1697 (N_1697,N_1504,N_1527);
nor U1698 (N_1698,N_1571,N_1572);
nand U1699 (N_1699,N_1548,N_1593);
and U1700 (N_1700,N_1622,N_1632);
or U1701 (N_1701,N_1607,N_1612);
nor U1702 (N_1702,N_1628,N_1630);
or U1703 (N_1703,N_1683,N_1641);
and U1704 (N_1704,N_1631,N_1650);
or U1705 (N_1705,N_1687,N_1620);
or U1706 (N_1706,N_1668,N_1663);
nand U1707 (N_1707,N_1633,N_1629);
nor U1708 (N_1708,N_1609,N_1666);
nor U1709 (N_1709,N_1655,N_1677);
nand U1710 (N_1710,N_1669,N_1670);
nand U1711 (N_1711,N_1610,N_1685);
and U1712 (N_1712,N_1693,N_1667);
nor U1713 (N_1713,N_1657,N_1605);
and U1714 (N_1714,N_1682,N_1603);
nor U1715 (N_1715,N_1688,N_1676);
or U1716 (N_1716,N_1621,N_1640);
nand U1717 (N_1717,N_1615,N_1619);
nand U1718 (N_1718,N_1606,N_1646);
or U1719 (N_1719,N_1699,N_1673);
nor U1720 (N_1720,N_1664,N_1692);
or U1721 (N_1721,N_1680,N_1651);
nand U1722 (N_1722,N_1636,N_1645);
and U1723 (N_1723,N_1681,N_1635);
or U1724 (N_1724,N_1686,N_1626);
or U1725 (N_1725,N_1665,N_1601);
and U1726 (N_1726,N_1694,N_1614);
and U1727 (N_1727,N_1600,N_1678);
and U1728 (N_1728,N_1644,N_1624);
nor U1729 (N_1729,N_1638,N_1660);
nand U1730 (N_1730,N_1653,N_1654);
nand U1731 (N_1731,N_1604,N_1698);
nor U1732 (N_1732,N_1679,N_1616);
or U1733 (N_1733,N_1671,N_1647);
or U1734 (N_1734,N_1613,N_1662);
and U1735 (N_1735,N_1674,N_1672);
nand U1736 (N_1736,N_1652,N_1634);
nor U1737 (N_1737,N_1618,N_1690);
nor U1738 (N_1738,N_1611,N_1675);
nor U1739 (N_1739,N_1617,N_1625);
nor U1740 (N_1740,N_1656,N_1608);
and U1741 (N_1741,N_1623,N_1695);
nand U1742 (N_1742,N_1639,N_1696);
and U1743 (N_1743,N_1642,N_1658);
nor U1744 (N_1744,N_1691,N_1648);
xnor U1745 (N_1745,N_1627,N_1643);
or U1746 (N_1746,N_1684,N_1649);
nor U1747 (N_1747,N_1689,N_1659);
or U1748 (N_1748,N_1661,N_1697);
and U1749 (N_1749,N_1602,N_1637);
xnor U1750 (N_1750,N_1643,N_1624);
nand U1751 (N_1751,N_1602,N_1668);
nor U1752 (N_1752,N_1608,N_1602);
nand U1753 (N_1753,N_1694,N_1630);
nor U1754 (N_1754,N_1635,N_1652);
and U1755 (N_1755,N_1659,N_1634);
nand U1756 (N_1756,N_1631,N_1641);
nor U1757 (N_1757,N_1648,N_1622);
nor U1758 (N_1758,N_1641,N_1624);
nand U1759 (N_1759,N_1612,N_1620);
and U1760 (N_1760,N_1676,N_1686);
nor U1761 (N_1761,N_1696,N_1684);
nand U1762 (N_1762,N_1618,N_1624);
or U1763 (N_1763,N_1667,N_1614);
nor U1764 (N_1764,N_1636,N_1693);
nand U1765 (N_1765,N_1661,N_1607);
and U1766 (N_1766,N_1676,N_1650);
or U1767 (N_1767,N_1615,N_1636);
or U1768 (N_1768,N_1670,N_1638);
or U1769 (N_1769,N_1695,N_1666);
nand U1770 (N_1770,N_1631,N_1645);
or U1771 (N_1771,N_1663,N_1654);
or U1772 (N_1772,N_1662,N_1699);
and U1773 (N_1773,N_1628,N_1642);
nand U1774 (N_1774,N_1652,N_1679);
nand U1775 (N_1775,N_1669,N_1630);
or U1776 (N_1776,N_1698,N_1662);
or U1777 (N_1777,N_1671,N_1626);
nor U1778 (N_1778,N_1612,N_1664);
and U1779 (N_1779,N_1617,N_1687);
nor U1780 (N_1780,N_1634,N_1604);
and U1781 (N_1781,N_1672,N_1691);
or U1782 (N_1782,N_1682,N_1647);
nand U1783 (N_1783,N_1625,N_1656);
nand U1784 (N_1784,N_1660,N_1649);
and U1785 (N_1785,N_1646,N_1686);
nor U1786 (N_1786,N_1690,N_1683);
nand U1787 (N_1787,N_1661,N_1658);
nor U1788 (N_1788,N_1685,N_1612);
nor U1789 (N_1789,N_1668,N_1665);
and U1790 (N_1790,N_1612,N_1695);
nand U1791 (N_1791,N_1683,N_1605);
and U1792 (N_1792,N_1605,N_1660);
and U1793 (N_1793,N_1686,N_1680);
or U1794 (N_1794,N_1647,N_1649);
nor U1795 (N_1795,N_1661,N_1663);
and U1796 (N_1796,N_1649,N_1612);
nand U1797 (N_1797,N_1628,N_1610);
nor U1798 (N_1798,N_1647,N_1604);
nor U1799 (N_1799,N_1689,N_1664);
nor U1800 (N_1800,N_1717,N_1786);
nand U1801 (N_1801,N_1706,N_1701);
nor U1802 (N_1802,N_1719,N_1758);
nor U1803 (N_1803,N_1788,N_1745);
nand U1804 (N_1804,N_1757,N_1760);
nor U1805 (N_1805,N_1724,N_1785);
nand U1806 (N_1806,N_1734,N_1744);
and U1807 (N_1807,N_1771,N_1714);
nand U1808 (N_1808,N_1783,N_1755);
and U1809 (N_1809,N_1732,N_1720);
and U1810 (N_1810,N_1794,N_1778);
and U1811 (N_1811,N_1723,N_1751);
and U1812 (N_1812,N_1774,N_1704);
nor U1813 (N_1813,N_1787,N_1707);
and U1814 (N_1814,N_1705,N_1782);
xnor U1815 (N_1815,N_1749,N_1743);
nor U1816 (N_1816,N_1799,N_1772);
or U1817 (N_1817,N_1746,N_1796);
nor U1818 (N_1818,N_1726,N_1798);
nor U1819 (N_1819,N_1750,N_1777);
or U1820 (N_1820,N_1752,N_1776);
or U1821 (N_1821,N_1735,N_1733);
or U1822 (N_1822,N_1767,N_1731);
or U1823 (N_1823,N_1741,N_1793);
nor U1824 (N_1824,N_1754,N_1721);
and U1825 (N_1825,N_1738,N_1722);
and U1826 (N_1826,N_1784,N_1740);
nand U1827 (N_1827,N_1713,N_1725);
or U1828 (N_1828,N_1775,N_1715);
nor U1829 (N_1829,N_1730,N_1728);
or U1830 (N_1830,N_1761,N_1702);
nand U1831 (N_1831,N_1766,N_1716);
nor U1832 (N_1832,N_1759,N_1765);
nor U1833 (N_1833,N_1768,N_1792);
nand U1834 (N_1834,N_1737,N_1797);
or U1835 (N_1835,N_1762,N_1742);
nor U1836 (N_1836,N_1709,N_1729);
nor U1837 (N_1837,N_1748,N_1795);
nand U1838 (N_1838,N_1756,N_1770);
nand U1839 (N_1839,N_1710,N_1712);
nor U1840 (N_1840,N_1763,N_1703);
and U1841 (N_1841,N_1781,N_1789);
or U1842 (N_1842,N_1764,N_1711);
xnor U1843 (N_1843,N_1747,N_1791);
nor U1844 (N_1844,N_1780,N_1753);
and U1845 (N_1845,N_1736,N_1718);
and U1846 (N_1846,N_1708,N_1769);
and U1847 (N_1847,N_1779,N_1790);
and U1848 (N_1848,N_1739,N_1700);
and U1849 (N_1849,N_1773,N_1727);
nor U1850 (N_1850,N_1739,N_1791);
nand U1851 (N_1851,N_1759,N_1745);
and U1852 (N_1852,N_1706,N_1784);
or U1853 (N_1853,N_1738,N_1702);
and U1854 (N_1854,N_1766,N_1772);
nand U1855 (N_1855,N_1751,N_1722);
nor U1856 (N_1856,N_1729,N_1775);
nand U1857 (N_1857,N_1758,N_1725);
or U1858 (N_1858,N_1732,N_1737);
nand U1859 (N_1859,N_1702,N_1743);
or U1860 (N_1860,N_1772,N_1768);
nand U1861 (N_1861,N_1759,N_1744);
or U1862 (N_1862,N_1705,N_1703);
or U1863 (N_1863,N_1799,N_1771);
xor U1864 (N_1864,N_1736,N_1757);
or U1865 (N_1865,N_1729,N_1794);
nor U1866 (N_1866,N_1709,N_1733);
nand U1867 (N_1867,N_1775,N_1765);
nand U1868 (N_1868,N_1705,N_1708);
and U1869 (N_1869,N_1745,N_1738);
nand U1870 (N_1870,N_1741,N_1754);
and U1871 (N_1871,N_1761,N_1711);
nand U1872 (N_1872,N_1753,N_1734);
nor U1873 (N_1873,N_1708,N_1702);
or U1874 (N_1874,N_1766,N_1759);
nand U1875 (N_1875,N_1729,N_1732);
nor U1876 (N_1876,N_1788,N_1743);
or U1877 (N_1877,N_1786,N_1723);
nor U1878 (N_1878,N_1716,N_1709);
nor U1879 (N_1879,N_1747,N_1709);
nor U1880 (N_1880,N_1757,N_1773);
or U1881 (N_1881,N_1751,N_1736);
or U1882 (N_1882,N_1721,N_1731);
or U1883 (N_1883,N_1723,N_1793);
and U1884 (N_1884,N_1758,N_1703);
nor U1885 (N_1885,N_1754,N_1727);
and U1886 (N_1886,N_1727,N_1723);
and U1887 (N_1887,N_1709,N_1787);
or U1888 (N_1888,N_1731,N_1739);
or U1889 (N_1889,N_1746,N_1704);
or U1890 (N_1890,N_1767,N_1759);
and U1891 (N_1891,N_1749,N_1744);
xnor U1892 (N_1892,N_1701,N_1779);
and U1893 (N_1893,N_1753,N_1764);
nor U1894 (N_1894,N_1768,N_1710);
nand U1895 (N_1895,N_1766,N_1705);
nand U1896 (N_1896,N_1734,N_1717);
and U1897 (N_1897,N_1766,N_1735);
or U1898 (N_1898,N_1761,N_1767);
and U1899 (N_1899,N_1797,N_1787);
nor U1900 (N_1900,N_1860,N_1890);
or U1901 (N_1901,N_1836,N_1849);
nor U1902 (N_1902,N_1829,N_1831);
and U1903 (N_1903,N_1822,N_1823);
and U1904 (N_1904,N_1856,N_1862);
and U1905 (N_1905,N_1839,N_1807);
nor U1906 (N_1906,N_1809,N_1870);
or U1907 (N_1907,N_1857,N_1848);
nand U1908 (N_1908,N_1816,N_1877);
nor U1909 (N_1909,N_1878,N_1893);
or U1910 (N_1910,N_1866,N_1815);
nor U1911 (N_1911,N_1887,N_1825);
nor U1912 (N_1912,N_1845,N_1882);
nand U1913 (N_1913,N_1879,N_1873);
and U1914 (N_1914,N_1837,N_1865);
nand U1915 (N_1915,N_1853,N_1827);
nand U1916 (N_1916,N_1864,N_1898);
nor U1917 (N_1917,N_1896,N_1812);
nand U1918 (N_1918,N_1844,N_1884);
and U1919 (N_1919,N_1820,N_1803);
or U1920 (N_1920,N_1892,N_1869);
nand U1921 (N_1921,N_1805,N_1880);
nand U1922 (N_1922,N_1824,N_1854);
and U1923 (N_1923,N_1881,N_1843);
nand U1924 (N_1924,N_1850,N_1886);
and U1925 (N_1925,N_1885,N_1863);
and U1926 (N_1926,N_1847,N_1851);
nor U1927 (N_1927,N_1874,N_1830);
nor U1928 (N_1928,N_1895,N_1800);
or U1929 (N_1929,N_1834,N_1833);
or U1930 (N_1930,N_1894,N_1813);
or U1931 (N_1931,N_1841,N_1835);
nand U1932 (N_1932,N_1808,N_1819);
nor U1933 (N_1933,N_1891,N_1868);
nand U1934 (N_1934,N_1840,N_1897);
nand U1935 (N_1935,N_1802,N_1861);
and U1936 (N_1936,N_1826,N_1888);
nand U1937 (N_1937,N_1806,N_1852);
nor U1938 (N_1938,N_1838,N_1858);
nor U1939 (N_1939,N_1871,N_1875);
nor U1940 (N_1940,N_1876,N_1810);
nor U1941 (N_1941,N_1855,N_1842);
and U1942 (N_1942,N_1846,N_1828);
and U1943 (N_1943,N_1899,N_1821);
nand U1944 (N_1944,N_1889,N_1883);
nand U1945 (N_1945,N_1817,N_1801);
nor U1946 (N_1946,N_1804,N_1818);
and U1947 (N_1947,N_1814,N_1872);
or U1948 (N_1948,N_1867,N_1832);
nor U1949 (N_1949,N_1811,N_1859);
nand U1950 (N_1950,N_1817,N_1861);
xnor U1951 (N_1951,N_1889,N_1832);
and U1952 (N_1952,N_1820,N_1897);
nor U1953 (N_1953,N_1896,N_1813);
nor U1954 (N_1954,N_1829,N_1810);
or U1955 (N_1955,N_1876,N_1855);
or U1956 (N_1956,N_1811,N_1850);
or U1957 (N_1957,N_1818,N_1899);
or U1958 (N_1958,N_1896,N_1880);
nand U1959 (N_1959,N_1893,N_1824);
or U1960 (N_1960,N_1852,N_1821);
or U1961 (N_1961,N_1837,N_1885);
and U1962 (N_1962,N_1845,N_1836);
nand U1963 (N_1963,N_1866,N_1873);
or U1964 (N_1964,N_1843,N_1838);
nor U1965 (N_1965,N_1868,N_1851);
nand U1966 (N_1966,N_1878,N_1846);
xor U1967 (N_1967,N_1804,N_1892);
xnor U1968 (N_1968,N_1862,N_1897);
nor U1969 (N_1969,N_1899,N_1898);
nand U1970 (N_1970,N_1849,N_1892);
or U1971 (N_1971,N_1844,N_1887);
nor U1972 (N_1972,N_1863,N_1899);
nor U1973 (N_1973,N_1840,N_1888);
and U1974 (N_1974,N_1882,N_1831);
or U1975 (N_1975,N_1824,N_1861);
or U1976 (N_1976,N_1830,N_1853);
or U1977 (N_1977,N_1847,N_1849);
or U1978 (N_1978,N_1885,N_1808);
nand U1979 (N_1979,N_1881,N_1894);
and U1980 (N_1980,N_1804,N_1852);
nand U1981 (N_1981,N_1823,N_1802);
and U1982 (N_1982,N_1888,N_1803);
nand U1983 (N_1983,N_1817,N_1869);
nand U1984 (N_1984,N_1806,N_1853);
nand U1985 (N_1985,N_1803,N_1813);
and U1986 (N_1986,N_1882,N_1895);
nor U1987 (N_1987,N_1868,N_1846);
and U1988 (N_1988,N_1873,N_1862);
or U1989 (N_1989,N_1816,N_1869);
nor U1990 (N_1990,N_1855,N_1834);
or U1991 (N_1991,N_1835,N_1872);
nor U1992 (N_1992,N_1838,N_1819);
nor U1993 (N_1993,N_1810,N_1820);
nand U1994 (N_1994,N_1850,N_1866);
nor U1995 (N_1995,N_1844,N_1804);
nor U1996 (N_1996,N_1854,N_1876);
nand U1997 (N_1997,N_1842,N_1883);
nand U1998 (N_1998,N_1867,N_1846);
nor U1999 (N_1999,N_1833,N_1836);
nand U2000 (N_2000,N_1991,N_1900);
nand U2001 (N_2001,N_1966,N_1984);
nor U2002 (N_2002,N_1989,N_1997);
or U2003 (N_2003,N_1957,N_1983);
xnor U2004 (N_2004,N_1978,N_1995);
or U2005 (N_2005,N_1905,N_1904);
or U2006 (N_2006,N_1926,N_1936);
or U2007 (N_2007,N_1986,N_1976);
and U2008 (N_2008,N_1999,N_1933);
nand U2009 (N_2009,N_1974,N_1911);
or U2010 (N_2010,N_1958,N_1918);
nor U2011 (N_2011,N_1964,N_1939);
and U2012 (N_2012,N_1955,N_1920);
or U2013 (N_2013,N_1975,N_1963);
and U2014 (N_2014,N_1944,N_1940);
and U2015 (N_2015,N_1993,N_1931);
nand U2016 (N_2016,N_1953,N_1951);
xnor U2017 (N_2017,N_1973,N_1987);
nand U2018 (N_2018,N_1956,N_1934);
or U2019 (N_2019,N_1927,N_1924);
nand U2020 (N_2020,N_1946,N_1945);
or U2021 (N_2021,N_1968,N_1922);
nand U2022 (N_2022,N_1943,N_1979);
or U2023 (N_2023,N_1948,N_1906);
or U2024 (N_2024,N_1954,N_1967);
xor U2025 (N_2025,N_1994,N_1932);
nand U2026 (N_2026,N_1941,N_1960);
and U2027 (N_2027,N_1950,N_1977);
nand U2028 (N_2028,N_1914,N_1902);
and U2029 (N_2029,N_1909,N_1928);
nand U2030 (N_2030,N_1969,N_1901);
and U2031 (N_2031,N_1972,N_1952);
nor U2032 (N_2032,N_1910,N_1985);
and U2033 (N_2033,N_1937,N_1970);
nor U2034 (N_2034,N_1988,N_1930);
nor U2035 (N_2035,N_1980,N_1935);
nand U2036 (N_2036,N_1961,N_1908);
xnor U2037 (N_2037,N_1919,N_1959);
or U2038 (N_2038,N_1962,N_1925);
nand U2039 (N_2039,N_1923,N_1971);
nand U2040 (N_2040,N_1982,N_1912);
nor U2041 (N_2041,N_1949,N_1981);
or U2042 (N_2042,N_1938,N_1915);
nor U2043 (N_2043,N_1907,N_1992);
and U2044 (N_2044,N_1921,N_1916);
nand U2045 (N_2045,N_1947,N_1913);
and U2046 (N_2046,N_1996,N_1942);
or U2047 (N_2047,N_1917,N_1965);
nand U2048 (N_2048,N_1929,N_1998);
nand U2049 (N_2049,N_1903,N_1990);
nor U2050 (N_2050,N_1976,N_1906);
nor U2051 (N_2051,N_1948,N_1988);
nand U2052 (N_2052,N_1948,N_1930);
nor U2053 (N_2053,N_1998,N_1980);
or U2054 (N_2054,N_1977,N_1979);
nor U2055 (N_2055,N_1962,N_1999);
or U2056 (N_2056,N_1921,N_1901);
nand U2057 (N_2057,N_1979,N_1926);
nor U2058 (N_2058,N_1952,N_1994);
nand U2059 (N_2059,N_1997,N_1981);
nor U2060 (N_2060,N_1990,N_1992);
nand U2061 (N_2061,N_1942,N_1958);
nand U2062 (N_2062,N_1900,N_1911);
xor U2063 (N_2063,N_1939,N_1923);
and U2064 (N_2064,N_1961,N_1937);
and U2065 (N_2065,N_1984,N_1929);
xnor U2066 (N_2066,N_1918,N_1952);
and U2067 (N_2067,N_1917,N_1968);
and U2068 (N_2068,N_1968,N_1996);
nor U2069 (N_2069,N_1988,N_1916);
or U2070 (N_2070,N_1906,N_1937);
nor U2071 (N_2071,N_1956,N_1947);
nor U2072 (N_2072,N_1981,N_1970);
or U2073 (N_2073,N_1978,N_1979);
xnor U2074 (N_2074,N_1982,N_1956);
and U2075 (N_2075,N_1925,N_1991);
xnor U2076 (N_2076,N_1916,N_1906);
nor U2077 (N_2077,N_1991,N_1955);
or U2078 (N_2078,N_1980,N_1921);
or U2079 (N_2079,N_1986,N_1933);
or U2080 (N_2080,N_1963,N_1962);
and U2081 (N_2081,N_1955,N_1954);
nor U2082 (N_2082,N_1967,N_1924);
and U2083 (N_2083,N_1911,N_1973);
nor U2084 (N_2084,N_1902,N_1923);
nand U2085 (N_2085,N_1902,N_1925);
nand U2086 (N_2086,N_1921,N_1902);
nand U2087 (N_2087,N_1901,N_1925);
and U2088 (N_2088,N_1932,N_1966);
and U2089 (N_2089,N_1984,N_1964);
and U2090 (N_2090,N_1960,N_1900);
nand U2091 (N_2091,N_1900,N_1952);
nand U2092 (N_2092,N_1913,N_1927);
xor U2093 (N_2093,N_1961,N_1955);
nand U2094 (N_2094,N_1971,N_1920);
and U2095 (N_2095,N_1974,N_1954);
and U2096 (N_2096,N_1944,N_1943);
nand U2097 (N_2097,N_1902,N_1985);
xnor U2098 (N_2098,N_1905,N_1921);
or U2099 (N_2099,N_1952,N_1912);
nand U2100 (N_2100,N_2083,N_2098);
or U2101 (N_2101,N_2056,N_2036);
and U2102 (N_2102,N_2007,N_2019);
and U2103 (N_2103,N_2079,N_2040);
nand U2104 (N_2104,N_2068,N_2086);
nor U2105 (N_2105,N_2064,N_2050);
nand U2106 (N_2106,N_2002,N_2067);
and U2107 (N_2107,N_2087,N_2058);
and U2108 (N_2108,N_2014,N_2015);
nor U2109 (N_2109,N_2065,N_2054);
nand U2110 (N_2110,N_2055,N_2011);
or U2111 (N_2111,N_2038,N_2071);
nor U2112 (N_2112,N_2006,N_2059);
or U2113 (N_2113,N_2082,N_2018);
nor U2114 (N_2114,N_2013,N_2045);
or U2115 (N_2115,N_2076,N_2037);
or U2116 (N_2116,N_2075,N_2093);
nor U2117 (N_2117,N_2091,N_2032);
and U2118 (N_2118,N_2001,N_2090);
and U2119 (N_2119,N_2053,N_2063);
and U2120 (N_2120,N_2051,N_2052);
and U2121 (N_2121,N_2042,N_2028);
nand U2122 (N_2122,N_2012,N_2030);
nor U2123 (N_2123,N_2048,N_2004);
and U2124 (N_2124,N_2074,N_2072);
or U2125 (N_2125,N_2069,N_2039);
nor U2126 (N_2126,N_2026,N_2073);
or U2127 (N_2127,N_2027,N_2005);
and U2128 (N_2128,N_2003,N_2000);
or U2129 (N_2129,N_2044,N_2099);
nand U2130 (N_2130,N_2025,N_2023);
or U2131 (N_2131,N_2094,N_2009);
nand U2132 (N_2132,N_2046,N_2070);
nor U2133 (N_2133,N_2088,N_2017);
nor U2134 (N_2134,N_2043,N_2035);
or U2135 (N_2135,N_2031,N_2057);
and U2136 (N_2136,N_2041,N_2084);
and U2137 (N_2137,N_2078,N_2024);
nor U2138 (N_2138,N_2077,N_2085);
nand U2139 (N_2139,N_2047,N_2029);
and U2140 (N_2140,N_2096,N_2016);
or U2141 (N_2141,N_2061,N_2080);
or U2142 (N_2142,N_2060,N_2020);
or U2143 (N_2143,N_2089,N_2097);
and U2144 (N_2144,N_2095,N_2066);
and U2145 (N_2145,N_2062,N_2008);
nor U2146 (N_2146,N_2081,N_2034);
and U2147 (N_2147,N_2021,N_2049);
nor U2148 (N_2148,N_2022,N_2010);
or U2149 (N_2149,N_2092,N_2033);
nand U2150 (N_2150,N_2088,N_2009);
and U2151 (N_2151,N_2007,N_2002);
or U2152 (N_2152,N_2005,N_2033);
nand U2153 (N_2153,N_2082,N_2002);
and U2154 (N_2154,N_2009,N_2041);
or U2155 (N_2155,N_2074,N_2070);
nand U2156 (N_2156,N_2060,N_2005);
and U2157 (N_2157,N_2042,N_2073);
or U2158 (N_2158,N_2067,N_2036);
or U2159 (N_2159,N_2032,N_2074);
nor U2160 (N_2160,N_2091,N_2089);
or U2161 (N_2161,N_2040,N_2016);
nand U2162 (N_2162,N_2097,N_2024);
and U2163 (N_2163,N_2051,N_2037);
or U2164 (N_2164,N_2037,N_2077);
nor U2165 (N_2165,N_2081,N_2033);
nand U2166 (N_2166,N_2066,N_2002);
and U2167 (N_2167,N_2065,N_2073);
nand U2168 (N_2168,N_2061,N_2086);
nor U2169 (N_2169,N_2062,N_2079);
nand U2170 (N_2170,N_2000,N_2033);
and U2171 (N_2171,N_2025,N_2005);
nand U2172 (N_2172,N_2063,N_2033);
or U2173 (N_2173,N_2000,N_2069);
xnor U2174 (N_2174,N_2012,N_2001);
nand U2175 (N_2175,N_2013,N_2063);
xor U2176 (N_2176,N_2044,N_2025);
or U2177 (N_2177,N_2010,N_2091);
nor U2178 (N_2178,N_2095,N_2063);
and U2179 (N_2179,N_2057,N_2017);
and U2180 (N_2180,N_2002,N_2076);
nor U2181 (N_2181,N_2008,N_2002);
nand U2182 (N_2182,N_2073,N_2017);
nand U2183 (N_2183,N_2088,N_2033);
nor U2184 (N_2184,N_2046,N_2005);
nor U2185 (N_2185,N_2054,N_2026);
and U2186 (N_2186,N_2053,N_2067);
nand U2187 (N_2187,N_2068,N_2051);
or U2188 (N_2188,N_2063,N_2024);
or U2189 (N_2189,N_2042,N_2012);
nand U2190 (N_2190,N_2092,N_2034);
and U2191 (N_2191,N_2097,N_2087);
or U2192 (N_2192,N_2012,N_2035);
or U2193 (N_2193,N_2080,N_2098);
or U2194 (N_2194,N_2030,N_2069);
or U2195 (N_2195,N_2084,N_2091);
nand U2196 (N_2196,N_2009,N_2085);
and U2197 (N_2197,N_2054,N_2096);
nand U2198 (N_2198,N_2068,N_2085);
or U2199 (N_2199,N_2062,N_2033);
nor U2200 (N_2200,N_2178,N_2130);
and U2201 (N_2201,N_2193,N_2123);
nor U2202 (N_2202,N_2139,N_2156);
or U2203 (N_2203,N_2142,N_2164);
and U2204 (N_2204,N_2152,N_2122);
nor U2205 (N_2205,N_2118,N_2159);
nand U2206 (N_2206,N_2185,N_2143);
or U2207 (N_2207,N_2182,N_2137);
or U2208 (N_2208,N_2187,N_2188);
or U2209 (N_2209,N_2138,N_2183);
and U2210 (N_2210,N_2150,N_2116);
and U2211 (N_2211,N_2100,N_2196);
nand U2212 (N_2212,N_2136,N_2110);
nand U2213 (N_2213,N_2162,N_2154);
nor U2214 (N_2214,N_2160,N_2135);
nor U2215 (N_2215,N_2144,N_2126);
and U2216 (N_2216,N_2168,N_2125);
nand U2217 (N_2217,N_2117,N_2170);
and U2218 (N_2218,N_2106,N_2119);
or U2219 (N_2219,N_2157,N_2189);
nand U2220 (N_2220,N_2171,N_2174);
and U2221 (N_2221,N_2102,N_2197);
nand U2222 (N_2222,N_2191,N_2105);
and U2223 (N_2223,N_2131,N_2108);
and U2224 (N_2224,N_2128,N_2111);
nand U2225 (N_2225,N_2127,N_2192);
nor U2226 (N_2226,N_2140,N_2175);
nand U2227 (N_2227,N_2186,N_2163);
and U2228 (N_2228,N_2199,N_2115);
or U2229 (N_2229,N_2166,N_2165);
and U2230 (N_2230,N_2177,N_2149);
or U2231 (N_2231,N_2181,N_2190);
and U2232 (N_2232,N_2129,N_2151);
or U2233 (N_2233,N_2146,N_2107);
nor U2234 (N_2234,N_2161,N_2109);
nand U2235 (N_2235,N_2145,N_2104);
nor U2236 (N_2236,N_2120,N_2195);
and U2237 (N_2237,N_2112,N_2113);
or U2238 (N_2238,N_2179,N_2133);
or U2239 (N_2239,N_2180,N_2169);
nand U2240 (N_2240,N_2173,N_2172);
xor U2241 (N_2241,N_2141,N_2167);
and U2242 (N_2242,N_2194,N_2176);
nor U2243 (N_2243,N_2158,N_2103);
nor U2244 (N_2244,N_2155,N_2101);
nand U2245 (N_2245,N_2114,N_2132);
nor U2246 (N_2246,N_2134,N_2153);
nor U2247 (N_2247,N_2148,N_2147);
xor U2248 (N_2248,N_2198,N_2184);
and U2249 (N_2249,N_2121,N_2124);
or U2250 (N_2250,N_2122,N_2178);
nand U2251 (N_2251,N_2169,N_2168);
nor U2252 (N_2252,N_2191,N_2166);
and U2253 (N_2253,N_2129,N_2188);
or U2254 (N_2254,N_2151,N_2101);
nor U2255 (N_2255,N_2169,N_2171);
or U2256 (N_2256,N_2152,N_2138);
nor U2257 (N_2257,N_2162,N_2140);
nor U2258 (N_2258,N_2147,N_2162);
and U2259 (N_2259,N_2122,N_2137);
nand U2260 (N_2260,N_2195,N_2197);
and U2261 (N_2261,N_2198,N_2133);
nand U2262 (N_2262,N_2108,N_2194);
nor U2263 (N_2263,N_2136,N_2100);
nor U2264 (N_2264,N_2104,N_2173);
nor U2265 (N_2265,N_2129,N_2166);
nor U2266 (N_2266,N_2173,N_2129);
nor U2267 (N_2267,N_2197,N_2109);
or U2268 (N_2268,N_2110,N_2159);
and U2269 (N_2269,N_2124,N_2151);
and U2270 (N_2270,N_2142,N_2171);
or U2271 (N_2271,N_2136,N_2164);
and U2272 (N_2272,N_2170,N_2155);
and U2273 (N_2273,N_2147,N_2179);
nand U2274 (N_2274,N_2156,N_2192);
or U2275 (N_2275,N_2188,N_2119);
or U2276 (N_2276,N_2104,N_2129);
nand U2277 (N_2277,N_2194,N_2163);
or U2278 (N_2278,N_2165,N_2134);
or U2279 (N_2279,N_2187,N_2174);
and U2280 (N_2280,N_2174,N_2146);
nor U2281 (N_2281,N_2137,N_2120);
and U2282 (N_2282,N_2139,N_2171);
nand U2283 (N_2283,N_2186,N_2128);
or U2284 (N_2284,N_2135,N_2107);
nand U2285 (N_2285,N_2136,N_2195);
nand U2286 (N_2286,N_2107,N_2170);
or U2287 (N_2287,N_2108,N_2168);
or U2288 (N_2288,N_2182,N_2156);
nor U2289 (N_2289,N_2101,N_2108);
and U2290 (N_2290,N_2171,N_2136);
nor U2291 (N_2291,N_2160,N_2113);
or U2292 (N_2292,N_2117,N_2104);
nand U2293 (N_2293,N_2109,N_2148);
xor U2294 (N_2294,N_2119,N_2138);
and U2295 (N_2295,N_2154,N_2117);
or U2296 (N_2296,N_2161,N_2191);
nor U2297 (N_2297,N_2143,N_2112);
nand U2298 (N_2298,N_2197,N_2183);
or U2299 (N_2299,N_2125,N_2115);
nand U2300 (N_2300,N_2238,N_2290);
or U2301 (N_2301,N_2237,N_2272);
nand U2302 (N_2302,N_2268,N_2298);
or U2303 (N_2303,N_2262,N_2299);
and U2304 (N_2304,N_2235,N_2294);
nor U2305 (N_2305,N_2270,N_2249);
or U2306 (N_2306,N_2211,N_2253);
and U2307 (N_2307,N_2274,N_2226);
and U2308 (N_2308,N_2263,N_2287);
and U2309 (N_2309,N_2250,N_2257);
or U2310 (N_2310,N_2256,N_2241);
nand U2311 (N_2311,N_2251,N_2276);
and U2312 (N_2312,N_2203,N_2229);
nand U2313 (N_2313,N_2205,N_2254);
or U2314 (N_2314,N_2281,N_2215);
nor U2315 (N_2315,N_2240,N_2239);
and U2316 (N_2316,N_2224,N_2209);
nand U2317 (N_2317,N_2282,N_2234);
nor U2318 (N_2318,N_2291,N_2265);
nor U2319 (N_2319,N_2207,N_2228);
nor U2320 (N_2320,N_2288,N_2217);
and U2321 (N_2321,N_2216,N_2236);
or U2322 (N_2322,N_2273,N_2201);
xor U2323 (N_2323,N_2231,N_2283);
or U2324 (N_2324,N_2200,N_2206);
or U2325 (N_2325,N_2225,N_2233);
and U2326 (N_2326,N_2204,N_2260);
nand U2327 (N_2327,N_2213,N_2223);
nand U2328 (N_2328,N_2292,N_2230);
or U2329 (N_2329,N_2208,N_2259);
and U2330 (N_2330,N_2261,N_2212);
xor U2331 (N_2331,N_2242,N_2284);
and U2332 (N_2332,N_2269,N_2258);
or U2333 (N_2333,N_2214,N_2279);
nand U2334 (N_2334,N_2246,N_2266);
nor U2335 (N_2335,N_2220,N_2267);
and U2336 (N_2336,N_2297,N_2202);
nor U2337 (N_2337,N_2245,N_2271);
nor U2338 (N_2338,N_2255,N_2278);
xor U2339 (N_2339,N_2227,N_2243);
xor U2340 (N_2340,N_2248,N_2285);
nor U2341 (N_2341,N_2286,N_2280);
and U2342 (N_2342,N_2210,N_2296);
or U2343 (N_2343,N_2293,N_2275);
or U2344 (N_2344,N_2252,N_2264);
and U2345 (N_2345,N_2222,N_2219);
nand U2346 (N_2346,N_2277,N_2295);
and U2347 (N_2347,N_2232,N_2218);
nor U2348 (N_2348,N_2289,N_2221);
nor U2349 (N_2349,N_2247,N_2244);
and U2350 (N_2350,N_2212,N_2259);
nand U2351 (N_2351,N_2284,N_2271);
nand U2352 (N_2352,N_2284,N_2236);
xor U2353 (N_2353,N_2223,N_2266);
and U2354 (N_2354,N_2229,N_2245);
nand U2355 (N_2355,N_2228,N_2258);
and U2356 (N_2356,N_2263,N_2252);
or U2357 (N_2357,N_2295,N_2239);
or U2358 (N_2358,N_2279,N_2243);
and U2359 (N_2359,N_2208,N_2251);
and U2360 (N_2360,N_2269,N_2267);
and U2361 (N_2361,N_2247,N_2291);
nor U2362 (N_2362,N_2230,N_2299);
nand U2363 (N_2363,N_2240,N_2292);
nor U2364 (N_2364,N_2241,N_2263);
or U2365 (N_2365,N_2290,N_2237);
nand U2366 (N_2366,N_2224,N_2223);
and U2367 (N_2367,N_2270,N_2204);
nor U2368 (N_2368,N_2273,N_2284);
nor U2369 (N_2369,N_2256,N_2200);
nand U2370 (N_2370,N_2216,N_2267);
xnor U2371 (N_2371,N_2298,N_2204);
or U2372 (N_2372,N_2272,N_2256);
or U2373 (N_2373,N_2234,N_2208);
nor U2374 (N_2374,N_2232,N_2212);
nor U2375 (N_2375,N_2233,N_2273);
nand U2376 (N_2376,N_2230,N_2239);
or U2377 (N_2377,N_2299,N_2205);
nor U2378 (N_2378,N_2275,N_2284);
xnor U2379 (N_2379,N_2259,N_2200);
or U2380 (N_2380,N_2243,N_2297);
and U2381 (N_2381,N_2235,N_2246);
nor U2382 (N_2382,N_2224,N_2261);
or U2383 (N_2383,N_2252,N_2297);
and U2384 (N_2384,N_2281,N_2239);
nor U2385 (N_2385,N_2255,N_2273);
nor U2386 (N_2386,N_2213,N_2220);
or U2387 (N_2387,N_2202,N_2281);
nand U2388 (N_2388,N_2203,N_2295);
nor U2389 (N_2389,N_2270,N_2223);
and U2390 (N_2390,N_2263,N_2217);
and U2391 (N_2391,N_2287,N_2214);
and U2392 (N_2392,N_2248,N_2273);
nand U2393 (N_2393,N_2269,N_2226);
or U2394 (N_2394,N_2271,N_2239);
and U2395 (N_2395,N_2246,N_2280);
nand U2396 (N_2396,N_2292,N_2211);
and U2397 (N_2397,N_2284,N_2232);
or U2398 (N_2398,N_2288,N_2259);
and U2399 (N_2399,N_2293,N_2214);
nand U2400 (N_2400,N_2310,N_2301);
nor U2401 (N_2401,N_2340,N_2336);
or U2402 (N_2402,N_2304,N_2392);
nand U2403 (N_2403,N_2343,N_2338);
or U2404 (N_2404,N_2370,N_2351);
nand U2405 (N_2405,N_2346,N_2321);
or U2406 (N_2406,N_2345,N_2371);
nand U2407 (N_2407,N_2305,N_2333);
nor U2408 (N_2408,N_2363,N_2360);
xor U2409 (N_2409,N_2359,N_2332);
nand U2410 (N_2410,N_2314,N_2367);
nor U2411 (N_2411,N_2390,N_2365);
nand U2412 (N_2412,N_2357,N_2373);
or U2413 (N_2413,N_2307,N_2318);
and U2414 (N_2414,N_2308,N_2328);
or U2415 (N_2415,N_2303,N_2323);
nor U2416 (N_2416,N_2383,N_2350);
nand U2417 (N_2417,N_2302,N_2382);
or U2418 (N_2418,N_2313,N_2316);
and U2419 (N_2419,N_2312,N_2355);
and U2420 (N_2420,N_2387,N_2388);
nor U2421 (N_2421,N_2342,N_2374);
nor U2422 (N_2422,N_2369,N_2368);
and U2423 (N_2423,N_2320,N_2306);
nand U2424 (N_2424,N_2389,N_2325);
nand U2425 (N_2425,N_2347,N_2330);
nor U2426 (N_2426,N_2300,N_2311);
and U2427 (N_2427,N_2394,N_2372);
and U2428 (N_2428,N_2391,N_2364);
nand U2429 (N_2429,N_2379,N_2324);
nand U2430 (N_2430,N_2358,N_2398);
nor U2431 (N_2431,N_2329,N_2376);
xor U2432 (N_2432,N_2397,N_2381);
and U2433 (N_2433,N_2326,N_2385);
nand U2434 (N_2434,N_2349,N_2366);
nand U2435 (N_2435,N_2322,N_2341);
or U2436 (N_2436,N_2309,N_2377);
and U2437 (N_2437,N_2384,N_2319);
and U2438 (N_2438,N_2378,N_2356);
nor U2439 (N_2439,N_2335,N_2327);
and U2440 (N_2440,N_2317,N_2339);
and U2441 (N_2441,N_2315,N_2354);
xor U2442 (N_2442,N_2399,N_2344);
and U2443 (N_2443,N_2353,N_2393);
nand U2444 (N_2444,N_2380,N_2352);
xnor U2445 (N_2445,N_2395,N_2361);
nor U2446 (N_2446,N_2331,N_2396);
nor U2447 (N_2447,N_2375,N_2337);
or U2448 (N_2448,N_2334,N_2362);
and U2449 (N_2449,N_2348,N_2386);
nor U2450 (N_2450,N_2320,N_2392);
and U2451 (N_2451,N_2304,N_2331);
and U2452 (N_2452,N_2324,N_2338);
and U2453 (N_2453,N_2353,N_2387);
nand U2454 (N_2454,N_2344,N_2303);
nor U2455 (N_2455,N_2387,N_2363);
nor U2456 (N_2456,N_2338,N_2333);
nand U2457 (N_2457,N_2396,N_2375);
and U2458 (N_2458,N_2314,N_2386);
and U2459 (N_2459,N_2310,N_2313);
nand U2460 (N_2460,N_2334,N_2357);
or U2461 (N_2461,N_2399,N_2333);
nor U2462 (N_2462,N_2385,N_2360);
nand U2463 (N_2463,N_2337,N_2302);
nor U2464 (N_2464,N_2370,N_2362);
and U2465 (N_2465,N_2320,N_2384);
xnor U2466 (N_2466,N_2326,N_2374);
and U2467 (N_2467,N_2317,N_2392);
and U2468 (N_2468,N_2348,N_2325);
nand U2469 (N_2469,N_2388,N_2350);
or U2470 (N_2470,N_2301,N_2355);
and U2471 (N_2471,N_2317,N_2380);
nand U2472 (N_2472,N_2384,N_2356);
nand U2473 (N_2473,N_2333,N_2349);
or U2474 (N_2474,N_2351,N_2367);
nand U2475 (N_2475,N_2398,N_2371);
and U2476 (N_2476,N_2362,N_2311);
nand U2477 (N_2477,N_2357,N_2303);
and U2478 (N_2478,N_2346,N_2309);
xnor U2479 (N_2479,N_2393,N_2392);
and U2480 (N_2480,N_2379,N_2375);
or U2481 (N_2481,N_2359,N_2346);
nand U2482 (N_2482,N_2378,N_2309);
nand U2483 (N_2483,N_2395,N_2393);
and U2484 (N_2484,N_2370,N_2322);
or U2485 (N_2485,N_2314,N_2375);
and U2486 (N_2486,N_2382,N_2315);
nor U2487 (N_2487,N_2315,N_2350);
or U2488 (N_2488,N_2382,N_2310);
and U2489 (N_2489,N_2344,N_2355);
or U2490 (N_2490,N_2397,N_2338);
and U2491 (N_2491,N_2356,N_2324);
nand U2492 (N_2492,N_2349,N_2330);
or U2493 (N_2493,N_2330,N_2365);
nand U2494 (N_2494,N_2328,N_2304);
nand U2495 (N_2495,N_2328,N_2342);
nand U2496 (N_2496,N_2390,N_2355);
or U2497 (N_2497,N_2328,N_2390);
or U2498 (N_2498,N_2326,N_2383);
nor U2499 (N_2499,N_2313,N_2339);
and U2500 (N_2500,N_2458,N_2495);
or U2501 (N_2501,N_2448,N_2498);
xor U2502 (N_2502,N_2480,N_2477);
nand U2503 (N_2503,N_2457,N_2417);
nor U2504 (N_2504,N_2465,N_2456);
nand U2505 (N_2505,N_2470,N_2413);
nor U2506 (N_2506,N_2403,N_2415);
and U2507 (N_2507,N_2410,N_2490);
or U2508 (N_2508,N_2430,N_2473);
nor U2509 (N_2509,N_2466,N_2497);
or U2510 (N_2510,N_2452,N_2454);
nand U2511 (N_2511,N_2488,N_2442);
and U2512 (N_2512,N_2444,N_2412);
or U2513 (N_2513,N_2482,N_2475);
and U2514 (N_2514,N_2418,N_2414);
nor U2515 (N_2515,N_2446,N_2440);
or U2516 (N_2516,N_2461,N_2432);
nand U2517 (N_2517,N_2424,N_2437);
and U2518 (N_2518,N_2464,N_2493);
xor U2519 (N_2519,N_2409,N_2460);
nor U2520 (N_2520,N_2489,N_2469);
nand U2521 (N_2521,N_2427,N_2425);
nand U2522 (N_2522,N_2499,N_2416);
or U2523 (N_2523,N_2435,N_2463);
nand U2524 (N_2524,N_2496,N_2478);
or U2525 (N_2525,N_2434,N_2449);
nor U2526 (N_2526,N_2402,N_2474);
or U2527 (N_2527,N_2428,N_2492);
or U2528 (N_2528,N_2467,N_2401);
or U2529 (N_2529,N_2407,N_2438);
xnor U2530 (N_2530,N_2421,N_2420);
nand U2531 (N_2531,N_2423,N_2447);
and U2532 (N_2532,N_2422,N_2436);
nor U2533 (N_2533,N_2431,N_2441);
nor U2534 (N_2534,N_2472,N_2443);
nand U2535 (N_2535,N_2451,N_2485);
nand U2536 (N_2536,N_2476,N_2419);
nand U2537 (N_2537,N_2453,N_2471);
and U2538 (N_2538,N_2406,N_2468);
and U2539 (N_2539,N_2400,N_2411);
or U2540 (N_2540,N_2426,N_2429);
and U2541 (N_2541,N_2486,N_2487);
or U2542 (N_2542,N_2404,N_2483);
nor U2543 (N_2543,N_2479,N_2433);
and U2544 (N_2544,N_2481,N_2450);
nand U2545 (N_2545,N_2445,N_2491);
or U2546 (N_2546,N_2455,N_2408);
nor U2547 (N_2547,N_2484,N_2494);
or U2548 (N_2548,N_2459,N_2405);
or U2549 (N_2549,N_2462,N_2439);
nor U2550 (N_2550,N_2441,N_2443);
nand U2551 (N_2551,N_2488,N_2426);
nand U2552 (N_2552,N_2418,N_2407);
nor U2553 (N_2553,N_2453,N_2462);
or U2554 (N_2554,N_2477,N_2475);
nand U2555 (N_2555,N_2429,N_2436);
or U2556 (N_2556,N_2421,N_2467);
xor U2557 (N_2557,N_2422,N_2464);
or U2558 (N_2558,N_2400,N_2478);
nor U2559 (N_2559,N_2451,N_2463);
nor U2560 (N_2560,N_2434,N_2408);
and U2561 (N_2561,N_2463,N_2441);
or U2562 (N_2562,N_2490,N_2477);
nor U2563 (N_2563,N_2449,N_2487);
or U2564 (N_2564,N_2407,N_2455);
and U2565 (N_2565,N_2494,N_2465);
or U2566 (N_2566,N_2420,N_2443);
or U2567 (N_2567,N_2497,N_2465);
and U2568 (N_2568,N_2459,N_2456);
and U2569 (N_2569,N_2452,N_2419);
nor U2570 (N_2570,N_2457,N_2412);
nand U2571 (N_2571,N_2490,N_2414);
nor U2572 (N_2572,N_2422,N_2463);
nor U2573 (N_2573,N_2435,N_2406);
nor U2574 (N_2574,N_2439,N_2490);
nor U2575 (N_2575,N_2465,N_2403);
or U2576 (N_2576,N_2470,N_2492);
and U2577 (N_2577,N_2440,N_2403);
nor U2578 (N_2578,N_2402,N_2459);
nor U2579 (N_2579,N_2476,N_2459);
nand U2580 (N_2580,N_2410,N_2487);
or U2581 (N_2581,N_2460,N_2425);
nor U2582 (N_2582,N_2402,N_2457);
and U2583 (N_2583,N_2492,N_2471);
and U2584 (N_2584,N_2450,N_2469);
nand U2585 (N_2585,N_2413,N_2484);
nand U2586 (N_2586,N_2472,N_2462);
and U2587 (N_2587,N_2437,N_2469);
nand U2588 (N_2588,N_2417,N_2458);
and U2589 (N_2589,N_2471,N_2417);
nor U2590 (N_2590,N_2456,N_2494);
xor U2591 (N_2591,N_2446,N_2403);
and U2592 (N_2592,N_2422,N_2404);
and U2593 (N_2593,N_2406,N_2450);
and U2594 (N_2594,N_2484,N_2455);
or U2595 (N_2595,N_2437,N_2446);
nor U2596 (N_2596,N_2413,N_2427);
or U2597 (N_2597,N_2489,N_2410);
nor U2598 (N_2598,N_2433,N_2402);
nor U2599 (N_2599,N_2477,N_2497);
nor U2600 (N_2600,N_2505,N_2531);
nor U2601 (N_2601,N_2574,N_2580);
nor U2602 (N_2602,N_2561,N_2565);
nand U2603 (N_2603,N_2530,N_2528);
and U2604 (N_2604,N_2548,N_2526);
nor U2605 (N_2605,N_2562,N_2571);
nor U2606 (N_2606,N_2522,N_2576);
and U2607 (N_2607,N_2547,N_2519);
nand U2608 (N_2608,N_2517,N_2536);
or U2609 (N_2609,N_2557,N_2523);
nand U2610 (N_2610,N_2567,N_2549);
nand U2611 (N_2611,N_2533,N_2573);
or U2612 (N_2612,N_2577,N_2556);
nand U2613 (N_2613,N_2501,N_2598);
and U2614 (N_2614,N_2541,N_2569);
and U2615 (N_2615,N_2550,N_2507);
nor U2616 (N_2616,N_2510,N_2546);
nand U2617 (N_2617,N_2570,N_2585);
nor U2618 (N_2618,N_2539,N_2583);
and U2619 (N_2619,N_2592,N_2588);
and U2620 (N_2620,N_2589,N_2511);
nand U2621 (N_2621,N_2540,N_2527);
and U2622 (N_2622,N_2599,N_2566);
or U2623 (N_2623,N_2534,N_2537);
nand U2624 (N_2624,N_2538,N_2553);
and U2625 (N_2625,N_2525,N_2514);
or U2626 (N_2626,N_2595,N_2529);
and U2627 (N_2627,N_2551,N_2543);
nor U2628 (N_2628,N_2503,N_2502);
and U2629 (N_2629,N_2559,N_2590);
nand U2630 (N_2630,N_2512,N_2575);
or U2631 (N_2631,N_2564,N_2532);
or U2632 (N_2632,N_2594,N_2500);
or U2633 (N_2633,N_2579,N_2587);
and U2634 (N_2634,N_2563,N_2568);
and U2635 (N_2635,N_2524,N_2508);
nand U2636 (N_2636,N_2535,N_2552);
nand U2637 (N_2637,N_2521,N_2596);
nor U2638 (N_2638,N_2518,N_2584);
nor U2639 (N_2639,N_2509,N_2558);
nor U2640 (N_2640,N_2555,N_2572);
or U2641 (N_2641,N_2597,N_2586);
nor U2642 (N_2642,N_2582,N_2506);
nand U2643 (N_2643,N_2560,N_2544);
nor U2644 (N_2644,N_2515,N_2504);
nand U2645 (N_2645,N_2520,N_2554);
and U2646 (N_2646,N_2545,N_2591);
nor U2647 (N_2647,N_2593,N_2513);
nor U2648 (N_2648,N_2581,N_2542);
or U2649 (N_2649,N_2578,N_2516);
and U2650 (N_2650,N_2569,N_2525);
and U2651 (N_2651,N_2596,N_2518);
and U2652 (N_2652,N_2586,N_2583);
nor U2653 (N_2653,N_2501,N_2510);
and U2654 (N_2654,N_2524,N_2594);
nor U2655 (N_2655,N_2511,N_2524);
nor U2656 (N_2656,N_2583,N_2533);
nor U2657 (N_2657,N_2528,N_2549);
nor U2658 (N_2658,N_2519,N_2557);
and U2659 (N_2659,N_2580,N_2504);
and U2660 (N_2660,N_2564,N_2574);
or U2661 (N_2661,N_2598,N_2532);
or U2662 (N_2662,N_2587,N_2539);
nand U2663 (N_2663,N_2501,N_2552);
xor U2664 (N_2664,N_2563,N_2500);
and U2665 (N_2665,N_2562,N_2514);
and U2666 (N_2666,N_2534,N_2503);
or U2667 (N_2667,N_2588,N_2516);
or U2668 (N_2668,N_2544,N_2551);
and U2669 (N_2669,N_2504,N_2564);
or U2670 (N_2670,N_2589,N_2537);
nor U2671 (N_2671,N_2557,N_2501);
nand U2672 (N_2672,N_2556,N_2554);
or U2673 (N_2673,N_2510,N_2506);
and U2674 (N_2674,N_2544,N_2527);
nor U2675 (N_2675,N_2578,N_2518);
and U2676 (N_2676,N_2575,N_2510);
and U2677 (N_2677,N_2595,N_2560);
and U2678 (N_2678,N_2542,N_2500);
nand U2679 (N_2679,N_2510,N_2526);
nor U2680 (N_2680,N_2509,N_2564);
or U2681 (N_2681,N_2535,N_2546);
and U2682 (N_2682,N_2595,N_2512);
nor U2683 (N_2683,N_2540,N_2531);
nor U2684 (N_2684,N_2571,N_2500);
nand U2685 (N_2685,N_2541,N_2585);
and U2686 (N_2686,N_2530,N_2569);
nand U2687 (N_2687,N_2570,N_2528);
nor U2688 (N_2688,N_2587,N_2585);
and U2689 (N_2689,N_2559,N_2566);
or U2690 (N_2690,N_2504,N_2585);
nand U2691 (N_2691,N_2568,N_2512);
nor U2692 (N_2692,N_2509,N_2591);
nor U2693 (N_2693,N_2597,N_2566);
and U2694 (N_2694,N_2574,N_2577);
or U2695 (N_2695,N_2593,N_2576);
xor U2696 (N_2696,N_2504,N_2588);
or U2697 (N_2697,N_2556,N_2513);
nor U2698 (N_2698,N_2541,N_2557);
nand U2699 (N_2699,N_2557,N_2514);
and U2700 (N_2700,N_2606,N_2676);
nor U2701 (N_2701,N_2610,N_2614);
and U2702 (N_2702,N_2634,N_2664);
nand U2703 (N_2703,N_2695,N_2690);
and U2704 (N_2704,N_2618,N_2620);
nand U2705 (N_2705,N_2678,N_2656);
or U2706 (N_2706,N_2612,N_2673);
nor U2707 (N_2707,N_2674,N_2652);
nand U2708 (N_2708,N_2669,N_2636);
and U2709 (N_2709,N_2686,N_2685);
nor U2710 (N_2710,N_2688,N_2611);
nor U2711 (N_2711,N_2662,N_2689);
nor U2712 (N_2712,N_2681,N_2672);
or U2713 (N_2713,N_2699,N_2613);
nand U2714 (N_2714,N_2645,N_2677);
nor U2715 (N_2715,N_2661,N_2698);
nand U2716 (N_2716,N_2658,N_2600);
and U2717 (N_2717,N_2670,N_2627);
or U2718 (N_2718,N_2629,N_2657);
or U2719 (N_2719,N_2609,N_2619);
and U2720 (N_2720,N_2647,N_2679);
nor U2721 (N_2721,N_2655,N_2607);
nand U2722 (N_2722,N_2666,N_2697);
nor U2723 (N_2723,N_2696,N_2640);
and U2724 (N_2724,N_2622,N_2649);
or U2725 (N_2725,N_2642,N_2683);
or U2726 (N_2726,N_2684,N_2601);
and U2727 (N_2727,N_2682,N_2631);
nor U2728 (N_2728,N_2687,N_2643);
or U2729 (N_2729,N_2660,N_2635);
nand U2730 (N_2730,N_2621,N_2632);
and U2731 (N_2731,N_2639,N_2671);
xor U2732 (N_2732,N_2659,N_2650);
nand U2733 (N_2733,N_2626,N_2608);
or U2734 (N_2734,N_2680,N_2653);
nand U2735 (N_2735,N_2604,N_2641);
nor U2736 (N_2736,N_2691,N_2667);
or U2737 (N_2737,N_2624,N_2603);
and U2738 (N_2738,N_2654,N_2648);
or U2739 (N_2739,N_2694,N_2605);
nor U2740 (N_2740,N_2651,N_2644);
nor U2741 (N_2741,N_2692,N_2615);
or U2742 (N_2742,N_2637,N_2693);
nand U2743 (N_2743,N_2616,N_2630);
xnor U2744 (N_2744,N_2623,N_2617);
and U2745 (N_2745,N_2628,N_2602);
or U2746 (N_2746,N_2646,N_2638);
nor U2747 (N_2747,N_2665,N_2633);
or U2748 (N_2748,N_2675,N_2668);
xnor U2749 (N_2749,N_2625,N_2663);
nor U2750 (N_2750,N_2693,N_2671);
or U2751 (N_2751,N_2695,N_2652);
and U2752 (N_2752,N_2684,N_2651);
nand U2753 (N_2753,N_2614,N_2615);
nand U2754 (N_2754,N_2639,N_2618);
nor U2755 (N_2755,N_2684,N_2677);
nand U2756 (N_2756,N_2658,N_2654);
or U2757 (N_2757,N_2664,N_2673);
or U2758 (N_2758,N_2679,N_2680);
nor U2759 (N_2759,N_2603,N_2658);
or U2760 (N_2760,N_2684,N_2676);
or U2761 (N_2761,N_2675,N_2626);
and U2762 (N_2762,N_2604,N_2688);
and U2763 (N_2763,N_2645,N_2629);
nor U2764 (N_2764,N_2636,N_2625);
and U2765 (N_2765,N_2676,N_2695);
nand U2766 (N_2766,N_2666,N_2601);
and U2767 (N_2767,N_2601,N_2698);
nor U2768 (N_2768,N_2695,N_2613);
nand U2769 (N_2769,N_2636,N_2664);
nor U2770 (N_2770,N_2656,N_2661);
and U2771 (N_2771,N_2686,N_2683);
or U2772 (N_2772,N_2622,N_2603);
or U2773 (N_2773,N_2669,N_2642);
nand U2774 (N_2774,N_2682,N_2692);
and U2775 (N_2775,N_2630,N_2692);
nand U2776 (N_2776,N_2653,N_2614);
and U2777 (N_2777,N_2699,N_2650);
or U2778 (N_2778,N_2630,N_2679);
or U2779 (N_2779,N_2626,N_2678);
nand U2780 (N_2780,N_2643,N_2600);
and U2781 (N_2781,N_2656,N_2695);
nand U2782 (N_2782,N_2632,N_2666);
or U2783 (N_2783,N_2648,N_2673);
and U2784 (N_2784,N_2636,N_2637);
nand U2785 (N_2785,N_2642,N_2659);
nand U2786 (N_2786,N_2620,N_2600);
nor U2787 (N_2787,N_2611,N_2619);
nor U2788 (N_2788,N_2609,N_2635);
nor U2789 (N_2789,N_2635,N_2657);
nor U2790 (N_2790,N_2654,N_2611);
nor U2791 (N_2791,N_2699,N_2654);
or U2792 (N_2792,N_2674,N_2644);
or U2793 (N_2793,N_2676,N_2623);
nand U2794 (N_2794,N_2661,N_2605);
and U2795 (N_2795,N_2665,N_2646);
nor U2796 (N_2796,N_2611,N_2658);
and U2797 (N_2797,N_2698,N_2662);
and U2798 (N_2798,N_2682,N_2622);
nand U2799 (N_2799,N_2617,N_2646);
or U2800 (N_2800,N_2764,N_2721);
or U2801 (N_2801,N_2782,N_2766);
nor U2802 (N_2802,N_2799,N_2737);
or U2803 (N_2803,N_2726,N_2772);
nand U2804 (N_2804,N_2769,N_2708);
or U2805 (N_2805,N_2732,N_2784);
nand U2806 (N_2806,N_2765,N_2701);
nand U2807 (N_2807,N_2750,N_2776);
or U2808 (N_2808,N_2709,N_2792);
nor U2809 (N_2809,N_2735,N_2786);
nand U2810 (N_2810,N_2759,N_2716);
nor U2811 (N_2811,N_2724,N_2717);
nand U2812 (N_2812,N_2727,N_2790);
and U2813 (N_2813,N_2719,N_2731);
nand U2814 (N_2814,N_2728,N_2730);
or U2815 (N_2815,N_2711,N_2720);
nand U2816 (N_2816,N_2788,N_2748);
and U2817 (N_2817,N_2729,N_2798);
nand U2818 (N_2818,N_2747,N_2794);
nor U2819 (N_2819,N_2751,N_2704);
nor U2820 (N_2820,N_2738,N_2779);
nand U2821 (N_2821,N_2725,N_2783);
nor U2822 (N_2822,N_2758,N_2700);
nor U2823 (N_2823,N_2778,N_2796);
or U2824 (N_2824,N_2793,N_2710);
nand U2825 (N_2825,N_2740,N_2718);
or U2826 (N_2826,N_2757,N_2762);
nor U2827 (N_2827,N_2703,N_2791);
and U2828 (N_2828,N_2797,N_2713);
and U2829 (N_2829,N_2745,N_2746);
nand U2830 (N_2830,N_2723,N_2763);
nor U2831 (N_2831,N_2787,N_2705);
nor U2832 (N_2832,N_2760,N_2753);
xnor U2833 (N_2833,N_2739,N_2702);
nor U2834 (N_2834,N_2755,N_2742);
and U2835 (N_2835,N_2771,N_2774);
or U2836 (N_2836,N_2773,N_2722);
nor U2837 (N_2837,N_2781,N_2734);
and U2838 (N_2838,N_2749,N_2736);
xnor U2839 (N_2839,N_2770,N_2733);
or U2840 (N_2840,N_2752,N_2761);
or U2841 (N_2841,N_2768,N_2706);
or U2842 (N_2842,N_2714,N_2744);
nand U2843 (N_2843,N_2785,N_2767);
or U2844 (N_2844,N_2780,N_2754);
and U2845 (N_2845,N_2777,N_2743);
or U2846 (N_2846,N_2715,N_2775);
nand U2847 (N_2847,N_2789,N_2795);
nand U2848 (N_2848,N_2756,N_2707);
and U2849 (N_2849,N_2712,N_2741);
and U2850 (N_2850,N_2763,N_2733);
or U2851 (N_2851,N_2703,N_2700);
nand U2852 (N_2852,N_2751,N_2750);
or U2853 (N_2853,N_2794,N_2716);
nand U2854 (N_2854,N_2758,N_2792);
or U2855 (N_2855,N_2747,N_2755);
or U2856 (N_2856,N_2700,N_2775);
and U2857 (N_2857,N_2771,N_2702);
xor U2858 (N_2858,N_2715,N_2735);
nor U2859 (N_2859,N_2798,N_2749);
or U2860 (N_2860,N_2733,N_2771);
and U2861 (N_2861,N_2718,N_2785);
and U2862 (N_2862,N_2766,N_2719);
nand U2863 (N_2863,N_2764,N_2749);
nor U2864 (N_2864,N_2744,N_2780);
nand U2865 (N_2865,N_2789,N_2752);
nand U2866 (N_2866,N_2723,N_2784);
nand U2867 (N_2867,N_2703,N_2715);
nand U2868 (N_2868,N_2793,N_2728);
nor U2869 (N_2869,N_2783,N_2758);
nor U2870 (N_2870,N_2790,N_2798);
nor U2871 (N_2871,N_2721,N_2706);
or U2872 (N_2872,N_2741,N_2718);
nand U2873 (N_2873,N_2756,N_2792);
and U2874 (N_2874,N_2759,N_2731);
and U2875 (N_2875,N_2705,N_2777);
nand U2876 (N_2876,N_2742,N_2751);
and U2877 (N_2877,N_2773,N_2707);
and U2878 (N_2878,N_2784,N_2729);
and U2879 (N_2879,N_2736,N_2723);
nor U2880 (N_2880,N_2724,N_2796);
or U2881 (N_2881,N_2763,N_2761);
and U2882 (N_2882,N_2708,N_2752);
or U2883 (N_2883,N_2730,N_2708);
nor U2884 (N_2884,N_2757,N_2780);
nand U2885 (N_2885,N_2738,N_2791);
nor U2886 (N_2886,N_2773,N_2787);
and U2887 (N_2887,N_2795,N_2785);
and U2888 (N_2888,N_2706,N_2795);
and U2889 (N_2889,N_2737,N_2726);
and U2890 (N_2890,N_2706,N_2775);
or U2891 (N_2891,N_2725,N_2723);
and U2892 (N_2892,N_2739,N_2745);
and U2893 (N_2893,N_2711,N_2741);
nand U2894 (N_2894,N_2742,N_2790);
xnor U2895 (N_2895,N_2762,N_2777);
nor U2896 (N_2896,N_2798,N_2714);
and U2897 (N_2897,N_2703,N_2764);
nor U2898 (N_2898,N_2715,N_2746);
and U2899 (N_2899,N_2748,N_2725);
and U2900 (N_2900,N_2860,N_2876);
and U2901 (N_2901,N_2867,N_2844);
and U2902 (N_2902,N_2800,N_2846);
nor U2903 (N_2903,N_2834,N_2858);
nand U2904 (N_2904,N_2828,N_2893);
nand U2905 (N_2905,N_2880,N_2855);
or U2906 (N_2906,N_2814,N_2856);
nand U2907 (N_2907,N_2833,N_2820);
nand U2908 (N_2908,N_2879,N_2850);
nor U2909 (N_2909,N_2889,N_2872);
nand U2910 (N_2910,N_2835,N_2857);
nand U2911 (N_2911,N_2881,N_2815);
and U2912 (N_2912,N_2830,N_2866);
nand U2913 (N_2913,N_2808,N_2892);
nor U2914 (N_2914,N_2803,N_2832);
nand U2915 (N_2915,N_2852,N_2824);
and U2916 (N_2916,N_2812,N_2851);
nor U2917 (N_2917,N_2826,N_2806);
nor U2918 (N_2918,N_2805,N_2877);
nor U2919 (N_2919,N_2891,N_2807);
nor U2920 (N_2920,N_2825,N_2888);
nor U2921 (N_2921,N_2809,N_2890);
nand U2922 (N_2922,N_2818,N_2887);
or U2923 (N_2923,N_2865,N_2804);
nor U2924 (N_2924,N_2895,N_2816);
nand U2925 (N_2925,N_2854,N_2839);
nor U2926 (N_2926,N_2841,N_2864);
xnor U2927 (N_2927,N_2821,N_2875);
nand U2928 (N_2928,N_2817,N_2896);
nor U2929 (N_2929,N_2870,N_2899);
nand U2930 (N_2930,N_2894,N_2897);
or U2931 (N_2931,N_2882,N_2869);
nor U2932 (N_2932,N_2885,N_2843);
and U2933 (N_2933,N_2801,N_2831);
and U2934 (N_2934,N_2847,N_2823);
nor U2935 (N_2935,N_2884,N_2898);
or U2936 (N_2936,N_2838,N_2861);
or U2937 (N_2937,N_2829,N_2848);
nand U2938 (N_2938,N_2883,N_2868);
nand U2939 (N_2939,N_2849,N_2886);
or U2940 (N_2940,N_2874,N_2837);
nand U2941 (N_2941,N_2840,N_2871);
nor U2942 (N_2942,N_2853,N_2842);
or U2943 (N_2943,N_2863,N_2802);
nand U2944 (N_2944,N_2859,N_2822);
xnor U2945 (N_2945,N_2862,N_2819);
nor U2946 (N_2946,N_2873,N_2811);
and U2947 (N_2947,N_2878,N_2845);
or U2948 (N_2948,N_2810,N_2836);
and U2949 (N_2949,N_2827,N_2813);
and U2950 (N_2950,N_2824,N_2867);
and U2951 (N_2951,N_2821,N_2884);
nand U2952 (N_2952,N_2853,N_2834);
or U2953 (N_2953,N_2863,N_2893);
nor U2954 (N_2954,N_2889,N_2800);
nor U2955 (N_2955,N_2885,N_2830);
nand U2956 (N_2956,N_2847,N_2842);
or U2957 (N_2957,N_2842,N_2815);
or U2958 (N_2958,N_2856,N_2862);
nand U2959 (N_2959,N_2823,N_2895);
nor U2960 (N_2960,N_2818,N_2880);
and U2961 (N_2961,N_2873,N_2857);
nor U2962 (N_2962,N_2841,N_2898);
nand U2963 (N_2963,N_2898,N_2887);
nor U2964 (N_2964,N_2849,N_2890);
or U2965 (N_2965,N_2810,N_2858);
nand U2966 (N_2966,N_2848,N_2857);
nand U2967 (N_2967,N_2803,N_2808);
or U2968 (N_2968,N_2897,N_2812);
nor U2969 (N_2969,N_2887,N_2813);
xor U2970 (N_2970,N_2848,N_2855);
xnor U2971 (N_2971,N_2883,N_2827);
and U2972 (N_2972,N_2863,N_2827);
or U2973 (N_2973,N_2822,N_2820);
and U2974 (N_2974,N_2811,N_2820);
nand U2975 (N_2975,N_2807,N_2897);
and U2976 (N_2976,N_2807,N_2870);
and U2977 (N_2977,N_2824,N_2811);
nand U2978 (N_2978,N_2819,N_2853);
nand U2979 (N_2979,N_2804,N_2840);
nor U2980 (N_2980,N_2803,N_2899);
nand U2981 (N_2981,N_2871,N_2853);
and U2982 (N_2982,N_2856,N_2888);
nand U2983 (N_2983,N_2893,N_2896);
nand U2984 (N_2984,N_2849,N_2869);
or U2985 (N_2985,N_2897,N_2815);
nand U2986 (N_2986,N_2881,N_2869);
nand U2987 (N_2987,N_2808,N_2881);
and U2988 (N_2988,N_2820,N_2807);
nor U2989 (N_2989,N_2889,N_2829);
and U2990 (N_2990,N_2823,N_2846);
nand U2991 (N_2991,N_2838,N_2818);
nor U2992 (N_2992,N_2889,N_2898);
nand U2993 (N_2993,N_2830,N_2809);
or U2994 (N_2994,N_2887,N_2810);
nand U2995 (N_2995,N_2837,N_2847);
or U2996 (N_2996,N_2808,N_2883);
nand U2997 (N_2997,N_2888,N_2839);
or U2998 (N_2998,N_2804,N_2800);
nand U2999 (N_2999,N_2892,N_2844);
nand UO_0 (O_0,N_2967,N_2940);
or UO_1 (O_1,N_2983,N_2912);
nor UO_2 (O_2,N_2937,N_2941);
or UO_3 (O_3,N_2905,N_2945);
or UO_4 (O_4,N_2908,N_2953);
or UO_5 (O_5,N_2947,N_2963);
nand UO_6 (O_6,N_2911,N_2920);
or UO_7 (O_7,N_2999,N_2927);
xnor UO_8 (O_8,N_2902,N_2921);
or UO_9 (O_9,N_2933,N_2982);
and UO_10 (O_10,N_2959,N_2992);
nor UO_11 (O_11,N_2900,N_2932);
nor UO_12 (O_12,N_2976,N_2934);
or UO_13 (O_13,N_2994,N_2951);
nor UO_14 (O_14,N_2962,N_2975);
or UO_15 (O_15,N_2977,N_2989);
and UO_16 (O_16,N_2942,N_2922);
and UO_17 (O_17,N_2923,N_2987);
and UO_18 (O_18,N_2960,N_2926);
nand UO_19 (O_19,N_2996,N_2991);
and UO_20 (O_20,N_2979,N_2970);
nor UO_21 (O_21,N_2997,N_2950);
nand UO_22 (O_22,N_2981,N_2931);
and UO_23 (O_23,N_2910,N_2915);
and UO_24 (O_24,N_2924,N_2939);
and UO_25 (O_25,N_2954,N_2901);
nand UO_26 (O_26,N_2944,N_2974);
or UO_27 (O_27,N_2966,N_2909);
nor UO_28 (O_28,N_2984,N_2957);
nor UO_29 (O_29,N_2973,N_2980);
nand UO_30 (O_30,N_2956,N_2938);
nor UO_31 (O_31,N_2961,N_2917);
and UO_32 (O_32,N_2985,N_2969);
nand UO_33 (O_33,N_2972,N_2929);
or UO_34 (O_34,N_2993,N_2918);
nand UO_35 (O_35,N_2971,N_2928);
nand UO_36 (O_36,N_2968,N_2930);
nor UO_37 (O_37,N_2935,N_2986);
nor UO_38 (O_38,N_2907,N_2988);
nor UO_39 (O_39,N_2936,N_2925);
and UO_40 (O_40,N_2955,N_2998);
and UO_41 (O_41,N_2952,N_2914);
xnor UO_42 (O_42,N_2946,N_2903);
nand UO_43 (O_43,N_2990,N_2958);
nor UO_44 (O_44,N_2965,N_2904);
nor UO_45 (O_45,N_2978,N_2949);
nand UO_46 (O_46,N_2948,N_2995);
nor UO_47 (O_47,N_2916,N_2964);
nor UO_48 (O_48,N_2913,N_2943);
or UO_49 (O_49,N_2906,N_2919);
or UO_50 (O_50,N_2982,N_2911);
nor UO_51 (O_51,N_2942,N_2975);
and UO_52 (O_52,N_2984,N_2983);
nand UO_53 (O_53,N_2951,N_2908);
nand UO_54 (O_54,N_2928,N_2951);
and UO_55 (O_55,N_2966,N_2950);
or UO_56 (O_56,N_2916,N_2948);
xnor UO_57 (O_57,N_2996,N_2960);
or UO_58 (O_58,N_2917,N_2954);
nor UO_59 (O_59,N_2949,N_2965);
nor UO_60 (O_60,N_2994,N_2981);
or UO_61 (O_61,N_2995,N_2924);
nand UO_62 (O_62,N_2993,N_2951);
or UO_63 (O_63,N_2941,N_2979);
and UO_64 (O_64,N_2967,N_2997);
and UO_65 (O_65,N_2918,N_2976);
nor UO_66 (O_66,N_2923,N_2979);
nand UO_67 (O_67,N_2930,N_2997);
nor UO_68 (O_68,N_2967,N_2984);
nor UO_69 (O_69,N_2948,N_2974);
xnor UO_70 (O_70,N_2913,N_2949);
and UO_71 (O_71,N_2992,N_2955);
nor UO_72 (O_72,N_2938,N_2997);
and UO_73 (O_73,N_2928,N_2958);
nand UO_74 (O_74,N_2928,N_2912);
and UO_75 (O_75,N_2936,N_2969);
nor UO_76 (O_76,N_2967,N_2992);
nor UO_77 (O_77,N_2992,N_2976);
nor UO_78 (O_78,N_2924,N_2979);
nand UO_79 (O_79,N_2920,N_2997);
and UO_80 (O_80,N_2963,N_2907);
or UO_81 (O_81,N_2930,N_2952);
and UO_82 (O_82,N_2923,N_2958);
or UO_83 (O_83,N_2936,N_2980);
nor UO_84 (O_84,N_2955,N_2995);
and UO_85 (O_85,N_2975,N_2995);
and UO_86 (O_86,N_2902,N_2905);
nor UO_87 (O_87,N_2918,N_2977);
or UO_88 (O_88,N_2915,N_2924);
and UO_89 (O_89,N_2972,N_2946);
or UO_90 (O_90,N_2950,N_2965);
or UO_91 (O_91,N_2982,N_2960);
nor UO_92 (O_92,N_2956,N_2953);
xor UO_93 (O_93,N_2908,N_2986);
or UO_94 (O_94,N_2912,N_2927);
nor UO_95 (O_95,N_2903,N_2938);
nand UO_96 (O_96,N_2909,N_2968);
or UO_97 (O_97,N_2992,N_2914);
nor UO_98 (O_98,N_2916,N_2926);
or UO_99 (O_99,N_2907,N_2940);
nand UO_100 (O_100,N_2963,N_2910);
or UO_101 (O_101,N_2925,N_2921);
nor UO_102 (O_102,N_2949,N_2904);
and UO_103 (O_103,N_2915,N_2998);
or UO_104 (O_104,N_2970,N_2981);
or UO_105 (O_105,N_2928,N_2954);
or UO_106 (O_106,N_2958,N_2934);
or UO_107 (O_107,N_2964,N_2979);
and UO_108 (O_108,N_2939,N_2945);
nand UO_109 (O_109,N_2955,N_2910);
nand UO_110 (O_110,N_2962,N_2903);
nor UO_111 (O_111,N_2991,N_2915);
nor UO_112 (O_112,N_2942,N_2925);
nand UO_113 (O_113,N_2914,N_2962);
or UO_114 (O_114,N_2970,N_2917);
nand UO_115 (O_115,N_2989,N_2975);
nand UO_116 (O_116,N_2926,N_2998);
nand UO_117 (O_117,N_2952,N_2944);
nand UO_118 (O_118,N_2922,N_2956);
nand UO_119 (O_119,N_2981,N_2979);
nand UO_120 (O_120,N_2937,N_2963);
or UO_121 (O_121,N_2955,N_2903);
nor UO_122 (O_122,N_2997,N_2913);
xor UO_123 (O_123,N_2939,N_2915);
nand UO_124 (O_124,N_2952,N_2991);
nand UO_125 (O_125,N_2903,N_2927);
nor UO_126 (O_126,N_2948,N_2967);
nand UO_127 (O_127,N_2976,N_2997);
nor UO_128 (O_128,N_2937,N_2934);
nor UO_129 (O_129,N_2992,N_2966);
or UO_130 (O_130,N_2913,N_2932);
and UO_131 (O_131,N_2974,N_2934);
and UO_132 (O_132,N_2982,N_2968);
nor UO_133 (O_133,N_2984,N_2959);
nand UO_134 (O_134,N_2907,N_2999);
and UO_135 (O_135,N_2900,N_2943);
nor UO_136 (O_136,N_2917,N_2907);
and UO_137 (O_137,N_2902,N_2979);
or UO_138 (O_138,N_2964,N_2960);
or UO_139 (O_139,N_2939,N_2968);
and UO_140 (O_140,N_2954,N_2950);
and UO_141 (O_141,N_2975,N_2902);
nor UO_142 (O_142,N_2948,N_2960);
nand UO_143 (O_143,N_2925,N_2911);
nand UO_144 (O_144,N_2902,N_2911);
nand UO_145 (O_145,N_2930,N_2940);
nand UO_146 (O_146,N_2915,N_2959);
or UO_147 (O_147,N_2925,N_2907);
nand UO_148 (O_148,N_2954,N_2999);
or UO_149 (O_149,N_2977,N_2947);
or UO_150 (O_150,N_2938,N_2902);
nand UO_151 (O_151,N_2983,N_2934);
nor UO_152 (O_152,N_2910,N_2918);
and UO_153 (O_153,N_2960,N_2937);
nor UO_154 (O_154,N_2912,N_2913);
or UO_155 (O_155,N_2981,N_2903);
or UO_156 (O_156,N_2969,N_2924);
and UO_157 (O_157,N_2970,N_2901);
and UO_158 (O_158,N_2986,N_2905);
nand UO_159 (O_159,N_2985,N_2987);
or UO_160 (O_160,N_2998,N_2937);
or UO_161 (O_161,N_2972,N_2986);
xnor UO_162 (O_162,N_2940,N_2955);
or UO_163 (O_163,N_2988,N_2937);
nand UO_164 (O_164,N_2917,N_2931);
nor UO_165 (O_165,N_2948,N_2915);
nand UO_166 (O_166,N_2952,N_2939);
nand UO_167 (O_167,N_2922,N_2906);
nor UO_168 (O_168,N_2987,N_2964);
and UO_169 (O_169,N_2961,N_2905);
nor UO_170 (O_170,N_2962,N_2906);
or UO_171 (O_171,N_2917,N_2926);
and UO_172 (O_172,N_2938,N_2993);
and UO_173 (O_173,N_2995,N_2903);
nand UO_174 (O_174,N_2984,N_2931);
nor UO_175 (O_175,N_2910,N_2924);
nand UO_176 (O_176,N_2925,N_2951);
or UO_177 (O_177,N_2926,N_2931);
nor UO_178 (O_178,N_2919,N_2989);
nor UO_179 (O_179,N_2961,N_2985);
nor UO_180 (O_180,N_2912,N_2923);
nand UO_181 (O_181,N_2952,N_2937);
and UO_182 (O_182,N_2974,N_2924);
and UO_183 (O_183,N_2970,N_2903);
nor UO_184 (O_184,N_2994,N_2944);
nand UO_185 (O_185,N_2996,N_2922);
nor UO_186 (O_186,N_2939,N_2917);
and UO_187 (O_187,N_2997,N_2983);
and UO_188 (O_188,N_2972,N_2969);
and UO_189 (O_189,N_2906,N_2944);
and UO_190 (O_190,N_2902,N_2958);
or UO_191 (O_191,N_2996,N_2914);
nand UO_192 (O_192,N_2986,N_2981);
and UO_193 (O_193,N_2957,N_2923);
nand UO_194 (O_194,N_2948,N_2939);
or UO_195 (O_195,N_2940,N_2986);
nand UO_196 (O_196,N_2979,N_2993);
or UO_197 (O_197,N_2958,N_2910);
nor UO_198 (O_198,N_2977,N_2969);
nand UO_199 (O_199,N_2909,N_2970);
nand UO_200 (O_200,N_2921,N_2928);
and UO_201 (O_201,N_2926,N_2905);
and UO_202 (O_202,N_2936,N_2979);
nor UO_203 (O_203,N_2944,N_2977);
nor UO_204 (O_204,N_2971,N_2926);
nor UO_205 (O_205,N_2944,N_2985);
or UO_206 (O_206,N_2977,N_2911);
nor UO_207 (O_207,N_2933,N_2915);
and UO_208 (O_208,N_2982,N_2910);
and UO_209 (O_209,N_2966,N_2970);
nor UO_210 (O_210,N_2929,N_2915);
nor UO_211 (O_211,N_2976,N_2943);
and UO_212 (O_212,N_2959,N_2932);
and UO_213 (O_213,N_2907,N_2953);
or UO_214 (O_214,N_2963,N_2985);
or UO_215 (O_215,N_2913,N_2916);
or UO_216 (O_216,N_2914,N_2913);
nor UO_217 (O_217,N_2950,N_2946);
nand UO_218 (O_218,N_2960,N_2976);
xor UO_219 (O_219,N_2945,N_2947);
and UO_220 (O_220,N_2928,N_2950);
xor UO_221 (O_221,N_2953,N_2992);
and UO_222 (O_222,N_2912,N_2920);
and UO_223 (O_223,N_2920,N_2967);
and UO_224 (O_224,N_2950,N_2969);
nor UO_225 (O_225,N_2971,N_2999);
and UO_226 (O_226,N_2961,N_2950);
or UO_227 (O_227,N_2945,N_2902);
and UO_228 (O_228,N_2986,N_2909);
nor UO_229 (O_229,N_2907,N_2967);
or UO_230 (O_230,N_2977,N_2925);
and UO_231 (O_231,N_2918,N_2908);
nand UO_232 (O_232,N_2965,N_2936);
or UO_233 (O_233,N_2971,N_2938);
nand UO_234 (O_234,N_2944,N_2948);
nand UO_235 (O_235,N_2923,N_2965);
or UO_236 (O_236,N_2906,N_2927);
nor UO_237 (O_237,N_2955,N_2958);
nor UO_238 (O_238,N_2960,N_2989);
or UO_239 (O_239,N_2975,N_2970);
nor UO_240 (O_240,N_2924,N_2903);
and UO_241 (O_241,N_2942,N_2993);
nor UO_242 (O_242,N_2950,N_2984);
and UO_243 (O_243,N_2905,N_2985);
and UO_244 (O_244,N_2905,N_2979);
nor UO_245 (O_245,N_2941,N_2976);
and UO_246 (O_246,N_2926,N_2962);
nor UO_247 (O_247,N_2923,N_2971);
and UO_248 (O_248,N_2921,N_2904);
and UO_249 (O_249,N_2988,N_2942);
xor UO_250 (O_250,N_2963,N_2905);
nor UO_251 (O_251,N_2903,N_2933);
and UO_252 (O_252,N_2951,N_2959);
and UO_253 (O_253,N_2912,N_2966);
nand UO_254 (O_254,N_2998,N_2992);
nand UO_255 (O_255,N_2905,N_2988);
nor UO_256 (O_256,N_2983,N_2910);
nor UO_257 (O_257,N_2916,N_2988);
or UO_258 (O_258,N_2915,N_2935);
or UO_259 (O_259,N_2995,N_2939);
and UO_260 (O_260,N_2952,N_2904);
or UO_261 (O_261,N_2963,N_2951);
or UO_262 (O_262,N_2915,N_2960);
nor UO_263 (O_263,N_2957,N_2997);
and UO_264 (O_264,N_2909,N_2950);
nand UO_265 (O_265,N_2955,N_2964);
xnor UO_266 (O_266,N_2987,N_2933);
nor UO_267 (O_267,N_2980,N_2954);
and UO_268 (O_268,N_2946,N_2998);
and UO_269 (O_269,N_2968,N_2924);
and UO_270 (O_270,N_2903,N_2989);
and UO_271 (O_271,N_2944,N_2915);
nand UO_272 (O_272,N_2993,N_2972);
and UO_273 (O_273,N_2941,N_2977);
and UO_274 (O_274,N_2900,N_2979);
nand UO_275 (O_275,N_2991,N_2906);
or UO_276 (O_276,N_2970,N_2952);
nand UO_277 (O_277,N_2987,N_2968);
or UO_278 (O_278,N_2936,N_2912);
nand UO_279 (O_279,N_2964,N_2908);
nand UO_280 (O_280,N_2927,N_2952);
nand UO_281 (O_281,N_2927,N_2918);
or UO_282 (O_282,N_2935,N_2944);
or UO_283 (O_283,N_2902,N_2964);
nor UO_284 (O_284,N_2971,N_2991);
nand UO_285 (O_285,N_2995,N_2965);
or UO_286 (O_286,N_2901,N_2949);
nand UO_287 (O_287,N_2962,N_2970);
nand UO_288 (O_288,N_2902,N_2955);
and UO_289 (O_289,N_2923,N_2933);
and UO_290 (O_290,N_2911,N_2972);
nand UO_291 (O_291,N_2920,N_2943);
or UO_292 (O_292,N_2938,N_2984);
or UO_293 (O_293,N_2965,N_2986);
or UO_294 (O_294,N_2980,N_2956);
and UO_295 (O_295,N_2942,N_2999);
and UO_296 (O_296,N_2942,N_2907);
or UO_297 (O_297,N_2922,N_2948);
nor UO_298 (O_298,N_2987,N_2937);
or UO_299 (O_299,N_2916,N_2901);
or UO_300 (O_300,N_2911,N_2917);
nor UO_301 (O_301,N_2969,N_2995);
and UO_302 (O_302,N_2979,N_2949);
nor UO_303 (O_303,N_2949,N_2948);
nor UO_304 (O_304,N_2936,N_2988);
nor UO_305 (O_305,N_2982,N_2990);
nand UO_306 (O_306,N_2964,N_2978);
nor UO_307 (O_307,N_2925,N_2961);
nand UO_308 (O_308,N_2939,N_2971);
and UO_309 (O_309,N_2914,N_2903);
and UO_310 (O_310,N_2981,N_2988);
and UO_311 (O_311,N_2947,N_2927);
or UO_312 (O_312,N_2961,N_2973);
nand UO_313 (O_313,N_2943,N_2940);
nand UO_314 (O_314,N_2972,N_2926);
nor UO_315 (O_315,N_2936,N_2916);
or UO_316 (O_316,N_2971,N_2901);
nor UO_317 (O_317,N_2966,N_2933);
nor UO_318 (O_318,N_2983,N_2939);
nor UO_319 (O_319,N_2997,N_2960);
nor UO_320 (O_320,N_2997,N_2953);
nand UO_321 (O_321,N_2951,N_2996);
and UO_322 (O_322,N_2960,N_2984);
nor UO_323 (O_323,N_2961,N_2986);
nand UO_324 (O_324,N_2948,N_2990);
nor UO_325 (O_325,N_2906,N_2992);
nor UO_326 (O_326,N_2974,N_2982);
nand UO_327 (O_327,N_2979,N_2992);
nor UO_328 (O_328,N_2953,N_2986);
nand UO_329 (O_329,N_2939,N_2970);
nand UO_330 (O_330,N_2928,N_2940);
or UO_331 (O_331,N_2992,N_2946);
nand UO_332 (O_332,N_2935,N_2922);
and UO_333 (O_333,N_2976,N_2928);
or UO_334 (O_334,N_2969,N_2940);
and UO_335 (O_335,N_2971,N_2930);
nand UO_336 (O_336,N_2982,N_2996);
nor UO_337 (O_337,N_2972,N_2919);
nor UO_338 (O_338,N_2988,N_2913);
xor UO_339 (O_339,N_2906,N_2935);
nor UO_340 (O_340,N_2913,N_2975);
and UO_341 (O_341,N_2972,N_2987);
or UO_342 (O_342,N_2967,N_2923);
or UO_343 (O_343,N_2934,N_2948);
and UO_344 (O_344,N_2902,N_2959);
nand UO_345 (O_345,N_2918,N_2992);
nand UO_346 (O_346,N_2904,N_2931);
and UO_347 (O_347,N_2914,N_2921);
and UO_348 (O_348,N_2901,N_2953);
and UO_349 (O_349,N_2910,N_2992);
or UO_350 (O_350,N_2962,N_2930);
nor UO_351 (O_351,N_2908,N_2917);
nor UO_352 (O_352,N_2941,N_2907);
and UO_353 (O_353,N_2950,N_2953);
nand UO_354 (O_354,N_2907,N_2919);
xnor UO_355 (O_355,N_2916,N_2934);
nor UO_356 (O_356,N_2947,N_2957);
and UO_357 (O_357,N_2958,N_2936);
or UO_358 (O_358,N_2916,N_2957);
and UO_359 (O_359,N_2991,N_2936);
or UO_360 (O_360,N_2904,N_2914);
and UO_361 (O_361,N_2960,N_2931);
nand UO_362 (O_362,N_2944,N_2932);
or UO_363 (O_363,N_2951,N_2924);
nand UO_364 (O_364,N_2994,N_2961);
nand UO_365 (O_365,N_2964,N_2925);
nor UO_366 (O_366,N_2917,N_2921);
nor UO_367 (O_367,N_2976,N_2945);
and UO_368 (O_368,N_2912,N_2918);
nand UO_369 (O_369,N_2949,N_2954);
nand UO_370 (O_370,N_2947,N_2991);
and UO_371 (O_371,N_2963,N_2960);
nor UO_372 (O_372,N_2991,N_2961);
xnor UO_373 (O_373,N_2999,N_2972);
or UO_374 (O_374,N_2909,N_2919);
and UO_375 (O_375,N_2930,N_2956);
nand UO_376 (O_376,N_2931,N_2985);
nor UO_377 (O_377,N_2929,N_2955);
and UO_378 (O_378,N_2942,N_2984);
nand UO_379 (O_379,N_2986,N_2941);
or UO_380 (O_380,N_2962,N_2923);
nand UO_381 (O_381,N_2953,N_2944);
xor UO_382 (O_382,N_2949,N_2908);
or UO_383 (O_383,N_2942,N_2977);
or UO_384 (O_384,N_2941,N_2910);
and UO_385 (O_385,N_2913,N_2968);
nand UO_386 (O_386,N_2943,N_2949);
nand UO_387 (O_387,N_2935,N_2983);
nor UO_388 (O_388,N_2937,N_2917);
nor UO_389 (O_389,N_2909,N_2906);
nand UO_390 (O_390,N_2943,N_2955);
and UO_391 (O_391,N_2921,N_2938);
and UO_392 (O_392,N_2986,N_2914);
nand UO_393 (O_393,N_2920,N_2909);
nand UO_394 (O_394,N_2993,N_2999);
nand UO_395 (O_395,N_2946,N_2918);
nor UO_396 (O_396,N_2968,N_2911);
or UO_397 (O_397,N_2959,N_2906);
nor UO_398 (O_398,N_2931,N_2993);
and UO_399 (O_399,N_2945,N_2952);
and UO_400 (O_400,N_2956,N_2990);
and UO_401 (O_401,N_2982,N_2925);
nor UO_402 (O_402,N_2935,N_2911);
nor UO_403 (O_403,N_2954,N_2972);
xor UO_404 (O_404,N_2947,N_2914);
nor UO_405 (O_405,N_2994,N_2934);
and UO_406 (O_406,N_2969,N_2937);
or UO_407 (O_407,N_2905,N_2933);
nand UO_408 (O_408,N_2905,N_2970);
nor UO_409 (O_409,N_2990,N_2980);
nor UO_410 (O_410,N_2980,N_2987);
and UO_411 (O_411,N_2901,N_2961);
and UO_412 (O_412,N_2980,N_2967);
nand UO_413 (O_413,N_2947,N_2943);
nor UO_414 (O_414,N_2924,N_2997);
nand UO_415 (O_415,N_2904,N_2960);
and UO_416 (O_416,N_2953,N_2930);
and UO_417 (O_417,N_2926,N_2938);
xnor UO_418 (O_418,N_2921,N_2966);
nor UO_419 (O_419,N_2985,N_2960);
nor UO_420 (O_420,N_2954,N_2985);
and UO_421 (O_421,N_2904,N_2986);
and UO_422 (O_422,N_2901,N_2910);
nand UO_423 (O_423,N_2953,N_2942);
xor UO_424 (O_424,N_2906,N_2917);
nand UO_425 (O_425,N_2995,N_2920);
nand UO_426 (O_426,N_2960,N_2927);
nor UO_427 (O_427,N_2903,N_2998);
nand UO_428 (O_428,N_2907,N_2982);
xnor UO_429 (O_429,N_2993,N_2983);
nand UO_430 (O_430,N_2940,N_2938);
or UO_431 (O_431,N_2979,N_2971);
nor UO_432 (O_432,N_2921,N_2954);
and UO_433 (O_433,N_2996,N_2948);
xnor UO_434 (O_434,N_2984,N_2997);
or UO_435 (O_435,N_2955,N_2945);
and UO_436 (O_436,N_2920,N_2921);
nor UO_437 (O_437,N_2956,N_2929);
nor UO_438 (O_438,N_2949,N_2938);
nand UO_439 (O_439,N_2954,N_2968);
xnor UO_440 (O_440,N_2962,N_2969);
or UO_441 (O_441,N_2903,N_2907);
nand UO_442 (O_442,N_2927,N_2983);
nand UO_443 (O_443,N_2987,N_2988);
and UO_444 (O_444,N_2928,N_2977);
nor UO_445 (O_445,N_2967,N_2903);
nor UO_446 (O_446,N_2920,N_2981);
nand UO_447 (O_447,N_2995,N_2985);
nand UO_448 (O_448,N_2944,N_2991);
and UO_449 (O_449,N_2967,N_2941);
nor UO_450 (O_450,N_2971,N_2905);
nor UO_451 (O_451,N_2977,N_2974);
nor UO_452 (O_452,N_2905,N_2972);
nor UO_453 (O_453,N_2985,N_2986);
or UO_454 (O_454,N_2986,N_2921);
or UO_455 (O_455,N_2931,N_2987);
nor UO_456 (O_456,N_2976,N_2921);
nand UO_457 (O_457,N_2906,N_2933);
and UO_458 (O_458,N_2929,N_2911);
or UO_459 (O_459,N_2965,N_2932);
nand UO_460 (O_460,N_2977,N_2988);
or UO_461 (O_461,N_2995,N_2973);
nor UO_462 (O_462,N_2959,N_2910);
nor UO_463 (O_463,N_2988,N_2966);
nor UO_464 (O_464,N_2990,N_2910);
nand UO_465 (O_465,N_2936,N_2996);
nand UO_466 (O_466,N_2903,N_2978);
nor UO_467 (O_467,N_2956,N_2910);
nor UO_468 (O_468,N_2923,N_2973);
nand UO_469 (O_469,N_2972,N_2922);
or UO_470 (O_470,N_2985,N_2932);
or UO_471 (O_471,N_2958,N_2957);
or UO_472 (O_472,N_2935,N_2954);
and UO_473 (O_473,N_2975,N_2934);
and UO_474 (O_474,N_2921,N_2949);
or UO_475 (O_475,N_2980,N_2902);
nand UO_476 (O_476,N_2992,N_2965);
or UO_477 (O_477,N_2936,N_2998);
and UO_478 (O_478,N_2919,N_2952);
or UO_479 (O_479,N_2988,N_2927);
nand UO_480 (O_480,N_2946,N_2932);
or UO_481 (O_481,N_2988,N_2990);
nand UO_482 (O_482,N_2910,N_2900);
nand UO_483 (O_483,N_2912,N_2999);
or UO_484 (O_484,N_2930,N_2937);
nor UO_485 (O_485,N_2911,N_2901);
nand UO_486 (O_486,N_2946,N_2928);
nand UO_487 (O_487,N_2982,N_2956);
and UO_488 (O_488,N_2933,N_2907);
nor UO_489 (O_489,N_2901,N_2992);
or UO_490 (O_490,N_2918,N_2961);
or UO_491 (O_491,N_2905,N_2937);
and UO_492 (O_492,N_2955,N_2907);
and UO_493 (O_493,N_2962,N_2951);
nand UO_494 (O_494,N_2982,N_2927);
or UO_495 (O_495,N_2975,N_2993);
or UO_496 (O_496,N_2987,N_2990);
nand UO_497 (O_497,N_2984,N_2961);
xnor UO_498 (O_498,N_2991,N_2910);
nand UO_499 (O_499,N_2940,N_2916);
endmodule