module basic_2000_20000_2500_4_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_1829,In_27);
or U1 (N_1,In_423,In_1180);
or U2 (N_2,In_1363,In_1735);
xor U3 (N_3,In_1774,In_64);
xor U4 (N_4,In_1654,In_1628);
nor U5 (N_5,In_1604,In_116);
xor U6 (N_6,In_1087,In_145);
and U7 (N_7,In_672,In_899);
xor U8 (N_8,In_1513,In_987);
or U9 (N_9,In_382,In_763);
or U10 (N_10,In_1530,In_1570);
nand U11 (N_11,In_1995,In_1270);
nor U12 (N_12,In_607,In_246);
nand U13 (N_13,In_1635,In_1780);
and U14 (N_14,In_451,In_66);
or U15 (N_15,In_1069,In_1719);
nand U16 (N_16,In_1267,In_1406);
nand U17 (N_17,In_749,In_1494);
xnor U18 (N_18,In_1967,In_715);
nor U19 (N_19,In_240,In_253);
nor U20 (N_20,In_661,In_162);
xor U21 (N_21,In_72,In_1279);
nand U22 (N_22,In_1788,In_479);
or U23 (N_23,In_366,In_202);
nand U24 (N_24,In_1748,In_1445);
or U25 (N_25,In_1928,In_105);
xor U26 (N_26,In_1534,In_480);
xor U27 (N_27,In_986,In_1629);
or U28 (N_28,In_1986,In_1124);
xor U29 (N_29,In_1236,In_1471);
xnor U30 (N_30,In_900,In_223);
nor U31 (N_31,In_130,In_941);
and U32 (N_32,In_503,In_853);
xnor U33 (N_33,In_723,In_669);
nor U34 (N_34,In_1386,In_292);
or U35 (N_35,In_1883,In_1500);
and U36 (N_36,In_412,In_3);
and U37 (N_37,In_1999,In_1097);
nand U38 (N_38,In_319,In_1094);
or U39 (N_39,In_422,In_1099);
xnor U40 (N_40,In_426,In_1259);
or U41 (N_41,In_991,In_946);
nand U42 (N_42,In_609,In_415);
and U43 (N_43,In_67,In_1324);
and U44 (N_44,In_1410,In_1474);
nand U45 (N_45,In_729,In_1865);
xor U46 (N_46,In_981,In_1765);
and U47 (N_47,In_1061,In_926);
or U48 (N_48,In_239,In_1319);
or U49 (N_49,In_784,In_1238);
xor U50 (N_50,In_1264,In_196);
xor U51 (N_51,In_1975,In_572);
xnor U52 (N_52,In_653,In_1804);
or U53 (N_53,In_1427,In_831);
or U54 (N_54,In_49,In_1593);
and U55 (N_55,In_1462,In_1492);
xor U56 (N_56,In_1280,In_1630);
and U57 (N_57,In_864,In_1390);
nor U58 (N_58,In_534,In_685);
nor U59 (N_59,In_1939,In_978);
xnor U60 (N_60,In_772,In_1556);
nand U61 (N_61,In_213,In_13);
and U62 (N_62,In_309,In_1712);
nand U63 (N_63,In_808,In_513);
nor U64 (N_64,In_1508,In_1090);
nand U65 (N_65,In_1218,In_378);
and U66 (N_66,In_172,In_1875);
or U67 (N_67,In_262,In_948);
nand U68 (N_68,In_1466,In_1373);
or U69 (N_69,In_1882,In_1920);
xnor U70 (N_70,In_1913,In_81);
xnor U71 (N_71,In_1790,In_376);
or U72 (N_72,In_102,In_1666);
or U73 (N_73,In_6,In_19);
and U74 (N_74,In_1917,In_320);
nor U75 (N_75,In_146,In_333);
or U76 (N_76,In_217,In_905);
or U77 (N_77,In_815,In_838);
and U78 (N_78,In_1538,In_577);
nand U79 (N_79,In_501,In_956);
xnor U80 (N_80,In_1825,In_1495);
xnor U81 (N_81,In_326,In_1045);
nand U82 (N_82,In_1395,In_457);
nor U83 (N_83,In_1950,In_256);
and U84 (N_84,In_1115,In_1755);
and U85 (N_85,In_1348,In_341);
nand U86 (N_86,In_716,In_757);
xor U87 (N_87,In_1844,In_1532);
nand U88 (N_88,In_1299,In_635);
nand U89 (N_89,In_1050,In_1442);
nor U90 (N_90,In_1220,In_1132);
nor U91 (N_91,In_335,In_231);
nand U92 (N_92,In_1961,In_1745);
and U93 (N_93,In_1842,In_1643);
and U94 (N_94,In_1232,In_1905);
xnor U95 (N_95,In_1853,In_869);
xor U96 (N_96,In_1358,In_295);
nor U97 (N_97,In_34,In_1794);
xor U98 (N_98,In_1268,In_390);
or U99 (N_99,In_1867,In_88);
or U100 (N_100,In_1980,In_1447);
or U101 (N_101,In_1426,In_446);
nand U102 (N_102,In_1720,In_1958);
and U103 (N_103,In_521,In_1199);
xnor U104 (N_104,In_346,In_252);
xnor U105 (N_105,In_682,In_1384);
nor U106 (N_106,In_797,In_1070);
nor U107 (N_107,In_1339,In_1903);
and U108 (N_108,In_884,In_238);
and U109 (N_109,In_505,In_478);
nand U110 (N_110,In_1891,In_135);
nand U111 (N_111,In_1775,In_1896);
xor U112 (N_112,In_325,In_929);
or U113 (N_113,In_149,In_187);
nor U114 (N_114,In_1456,In_1375);
nand U115 (N_115,In_1713,In_1658);
xnor U116 (N_116,In_278,In_1707);
nor U117 (N_117,In_488,In_1681);
or U118 (N_118,In_212,In_518);
xnor U119 (N_119,In_449,In_337);
or U120 (N_120,In_355,In_1607);
nor U121 (N_121,In_1443,In_1831);
or U122 (N_122,In_1371,In_1816);
or U123 (N_123,In_758,In_975);
and U124 (N_124,In_1152,In_1849);
xor U125 (N_125,In_1465,In_448);
nor U126 (N_126,In_621,In_1838);
and U127 (N_127,In_1457,In_874);
nor U128 (N_128,In_526,In_1473);
or U129 (N_129,In_314,In_51);
and U130 (N_130,In_143,In_110);
or U131 (N_131,In_509,In_357);
nor U132 (N_132,In_1893,In_1388);
and U133 (N_133,In_552,In_730);
or U134 (N_134,In_396,In_1423);
nor U135 (N_135,In_1496,In_1901);
or U136 (N_136,In_80,In_680);
or U137 (N_137,In_9,In_1082);
and U138 (N_138,In_544,In_454);
or U139 (N_139,In_507,In_988);
or U140 (N_140,In_768,In_1540);
nand U141 (N_141,In_1753,In_912);
or U142 (N_142,In_304,In_1313);
xor U143 (N_143,In_1291,In_1321);
or U144 (N_144,In_566,In_1800);
nor U145 (N_145,In_1285,In_351);
or U146 (N_146,In_1524,In_1173);
nand U147 (N_147,In_1618,In_1596);
nand U148 (N_148,In_1506,In_261);
nand U149 (N_149,In_127,In_628);
and U150 (N_150,In_101,In_134);
nor U151 (N_151,In_1481,In_1163);
or U152 (N_152,In_1702,In_484);
xnor U153 (N_153,In_637,In_430);
or U154 (N_154,In_1143,In_828);
nor U155 (N_155,In_1779,In_1963);
and U156 (N_156,In_235,In_475);
nor U157 (N_157,In_183,In_54);
nand U158 (N_158,In_55,In_192);
nand U159 (N_159,In_342,In_1729);
or U160 (N_160,In_1365,In_236);
and U161 (N_161,In_474,In_1158);
xor U162 (N_162,In_1409,In_995);
nand U163 (N_163,In_303,In_1847);
nor U164 (N_164,In_1294,In_736);
and U165 (N_165,In_1919,In_1974);
and U166 (N_166,In_321,In_617);
and U167 (N_167,In_955,In_1212);
xor U168 (N_168,In_1142,In_530);
or U169 (N_169,In_750,In_1942);
or U170 (N_170,In_1116,In_1487);
or U171 (N_171,In_1167,In_892);
nor U172 (N_172,In_490,In_582);
xor U173 (N_173,In_1472,In_129);
and U174 (N_174,In_767,In_463);
nand U175 (N_175,In_1572,In_845);
nand U176 (N_176,In_1726,In_1554);
xnor U177 (N_177,In_1664,In_456);
and U178 (N_178,In_322,In_1505);
or U179 (N_179,In_695,In_234);
or U180 (N_180,In_1455,In_860);
and U181 (N_181,In_197,In_691);
xor U182 (N_182,In_1960,In_1764);
or U183 (N_183,In_22,In_570);
xor U184 (N_184,In_812,In_734);
and U185 (N_185,In_1971,In_622);
and U186 (N_186,In_1636,In_1183);
nand U187 (N_187,In_316,In_43);
nor U188 (N_188,In_26,In_1811);
nor U189 (N_189,In_397,In_520);
xnor U190 (N_190,In_408,In_1823);
xor U191 (N_191,In_1200,In_1688);
and U192 (N_192,In_20,In_1172);
and U193 (N_193,In_1906,In_1965);
or U194 (N_194,In_1011,In_180);
and U195 (N_195,In_282,In_458);
xnor U196 (N_196,In_837,In_1044);
or U197 (N_197,In_1955,In_538);
or U198 (N_198,In_1957,In_330);
or U199 (N_199,In_392,In_910);
and U200 (N_200,In_1073,In_1036);
nor U201 (N_201,In_755,In_189);
xor U202 (N_202,In_1921,In_1425);
nand U203 (N_203,In_1485,In_895);
xor U204 (N_204,In_574,In_851);
xnor U205 (N_205,In_1542,In_265);
and U206 (N_206,In_1568,In_207);
or U207 (N_207,In_612,In_1504);
or U208 (N_208,In_1668,In_2);
nor U209 (N_209,In_754,In_1626);
nand U210 (N_210,In_643,In_965);
xnor U211 (N_211,In_1886,In_191);
xnor U212 (N_212,In_760,In_1146);
xnor U213 (N_213,In_377,In_546);
nor U214 (N_214,In_391,In_1047);
or U215 (N_215,In_1298,In_1791);
nand U216 (N_216,In_1512,In_1012);
xor U217 (N_217,In_30,In_1102);
xnor U218 (N_218,In_935,In_636);
nor U219 (N_219,In_1761,In_1897);
xnor U220 (N_220,In_863,In_1461);
nand U221 (N_221,In_111,In_1213);
and U222 (N_222,In_218,In_746);
nor U223 (N_223,In_268,In_85);
nand U224 (N_224,In_1598,In_1413);
xnor U225 (N_225,In_571,In_388);
or U226 (N_226,In_974,In_1938);
nor U227 (N_227,In_891,In_1229);
nor U228 (N_228,In_1340,In_1994);
xnor U229 (N_229,In_249,In_692);
and U230 (N_230,In_1223,In_568);
nand U231 (N_231,In_561,In_533);
and U232 (N_232,In_1907,In_1450);
and U233 (N_233,In_620,In_798);
xor U234 (N_234,In_1813,In_1689);
and U235 (N_235,In_244,In_1981);
nor U236 (N_236,In_290,In_704);
and U237 (N_237,In_1149,In_293);
and U238 (N_238,In_927,In_250);
or U239 (N_239,In_283,In_558);
and U240 (N_240,In_1076,In_1065);
and U241 (N_241,In_318,In_1013);
and U242 (N_242,In_676,In_447);
and U243 (N_243,In_1641,In_1184);
nand U244 (N_244,In_597,In_1204);
xnor U245 (N_245,In_1262,In_1990);
xnor U246 (N_246,In_587,In_69);
nand U247 (N_247,In_997,In_1064);
and U248 (N_248,In_897,In_1943);
nand U249 (N_249,In_940,In_1966);
or U250 (N_250,In_1600,In_59);
xor U251 (N_251,In_1347,In_839);
and U252 (N_252,In_159,In_462);
nand U253 (N_253,In_114,In_1731);
and U254 (N_254,In_1118,In_1736);
xor U255 (N_255,In_1412,In_1873);
nor U256 (N_256,In_1150,In_302);
and U257 (N_257,In_164,In_1468);
or U258 (N_258,In_1746,In_1756);
and U259 (N_259,In_1710,In_737);
nor U260 (N_260,In_1740,In_194);
nand U261 (N_261,In_1916,In_1095);
nand U262 (N_262,In_1329,In_32);
xor U263 (N_263,In_324,In_1718);
or U264 (N_264,In_73,In_1252);
and U265 (N_265,In_1805,In_800);
nor U266 (N_266,In_764,In_923);
nand U267 (N_267,In_151,In_259);
or U268 (N_268,In_1130,In_274);
xnor U269 (N_269,In_1246,In_1098);
nand U270 (N_270,In_108,In_858);
nor U271 (N_271,In_1219,In_1429);
and U272 (N_272,In_1161,In_854);
nor U273 (N_273,In_7,In_1871);
xor U274 (N_274,In_1595,In_565);
and U275 (N_275,In_793,In_272);
and U276 (N_276,In_1640,In_386);
nor U277 (N_277,In_1562,In_1430);
nor U278 (N_278,In_226,In_1162);
nor U279 (N_279,In_525,In_799);
xor U280 (N_280,In_623,In_467);
and U281 (N_281,In_352,In_1028);
nand U282 (N_282,In_1603,In_1970);
or U283 (N_283,In_395,In_1422);
xor U284 (N_284,In_701,In_1139);
nor U285 (N_285,In_1634,In_1516);
or U286 (N_286,In_1803,In_762);
or U287 (N_287,In_1749,In_407);
nor U288 (N_288,In_411,In_563);
nand U289 (N_289,In_611,In_169);
and U290 (N_290,In_1397,In_747);
xnor U291 (N_291,In_911,In_204);
xnor U292 (N_292,In_470,In_1205);
and U293 (N_293,In_270,In_638);
and U294 (N_294,In_1079,In_1850);
and U295 (N_295,In_751,In_971);
or U296 (N_296,In_924,In_708);
xnor U297 (N_297,In_340,In_1863);
nand U298 (N_298,In_728,In_1032);
or U299 (N_299,In_489,In_1667);
nand U300 (N_300,In_588,In_1711);
or U301 (N_301,In_1052,In_631);
or U302 (N_302,In_976,In_1208);
and U303 (N_303,In_285,In_90);
and U304 (N_304,In_1002,In_684);
nor U305 (N_305,In_1314,In_1704);
nand U306 (N_306,In_158,In_1334);
xor U307 (N_307,In_1344,In_1039);
xnor U308 (N_308,In_1864,In_1801);
nand U309 (N_309,In_1698,In_1117);
and U310 (N_310,In_1337,In_429);
nand U311 (N_311,In_967,In_527);
and U312 (N_312,In_1126,In_1523);
and U313 (N_313,In_57,In_286);
and U314 (N_314,In_1378,In_1571);
xnor U315 (N_315,In_1781,In_649);
nand U316 (N_316,In_1787,In_508);
xnor U317 (N_317,In_78,In_725);
nand U318 (N_318,In_1341,In_868);
or U319 (N_319,In_1522,In_549);
nand U320 (N_320,In_1066,In_913);
and U321 (N_321,In_1936,In_908);
and U322 (N_322,In_1545,In_1862);
or U323 (N_323,In_267,In_774);
nor U324 (N_324,In_724,In_296);
or U325 (N_325,In_1660,In_95);
or U326 (N_326,In_1946,In_671);
or U327 (N_327,In_444,In_1945);
and U328 (N_328,In_44,In_1125);
nand U329 (N_329,In_175,In_979);
nand U330 (N_330,In_771,In_539);
or U331 (N_331,In_880,In_14);
or U332 (N_332,In_156,In_354);
xnor U333 (N_333,In_707,In_1541);
or U334 (N_334,In_792,In_883);
nor U335 (N_335,In_742,In_632);
nand U336 (N_336,In_990,In_1777);
xor U337 (N_337,In_495,In_220);
nand U338 (N_338,In_210,In_1501);
nor U339 (N_339,In_94,In_807);
and U340 (N_340,In_1843,In_994);
nand U341 (N_341,In_1049,In_1295);
nand U342 (N_342,In_1104,In_1573);
nor U343 (N_343,In_1215,In_548);
and U344 (N_344,In_846,In_616);
xor U345 (N_345,In_1996,In_23);
nor U346 (N_346,In_497,In_1464);
xor U347 (N_347,In_1349,In_1296);
xnor U348 (N_348,In_711,In_600);
xnor U349 (N_349,In_1679,In_405);
or U350 (N_350,In_1058,In_1156);
and U351 (N_351,In_810,In_1927);
nor U352 (N_352,In_1467,In_190);
nor U353 (N_353,In_1354,In_343);
nor U354 (N_354,In_1376,In_1237);
and U355 (N_355,In_348,In_222);
or U356 (N_356,In_882,In_1480);
nor U357 (N_357,In_1860,In_1539);
nor U358 (N_358,In_1870,In_1320);
xor U359 (N_359,In_641,In_1370);
nor U360 (N_360,In_694,In_440);
or U361 (N_361,In_977,In_1389);
nor U362 (N_362,In_424,In_410);
or U363 (N_363,In_425,In_150);
or U364 (N_364,In_604,In_1109);
nor U365 (N_365,In_954,In_1725);
or U366 (N_366,In_1866,In_1226);
and U367 (N_367,In_719,In_1317);
and U368 (N_368,In_17,In_1451);
or U369 (N_369,In_1675,In_970);
and U370 (N_370,In_1091,In_589);
nor U371 (N_371,In_1776,In_1715);
and U372 (N_372,In_1484,In_1869);
nor U373 (N_373,In_1005,In_1227);
xor U374 (N_374,In_417,In_1686);
xor U375 (N_375,In_1682,In_816);
xnor U376 (N_376,In_1806,In_416);
xor U377 (N_377,In_515,In_1954);
or U378 (N_378,In_1260,In_761);
xor U379 (N_379,In_317,In_394);
nand U380 (N_380,In_1733,In_855);
nor U381 (N_381,In_1657,In_400);
nand U382 (N_382,In_174,In_919);
nand U383 (N_383,In_1716,In_60);
and U384 (N_384,In_1851,In_713);
nor U385 (N_385,In_1855,In_1224);
or U386 (N_386,In_1263,In_1287);
xor U387 (N_387,In_1356,In_586);
nand U388 (N_388,In_119,In_1414);
nand U389 (N_389,In_46,In_567);
and U390 (N_390,In_361,In_115);
xnor U391 (N_391,In_1690,In_966);
and U392 (N_392,In_1123,In_675);
nand U393 (N_393,In_91,In_1819);
nor U394 (N_394,In_1489,In_113);
xnor U395 (N_395,In_1799,In_1385);
and U396 (N_396,In_1581,In_531);
nor U397 (N_397,In_705,In_1826);
and U398 (N_398,In_254,In_1724);
nor U399 (N_399,In_540,In_1709);
or U400 (N_400,In_275,In_1773);
or U401 (N_401,In_1821,In_1056);
xor U402 (N_402,In_1216,In_1105);
nand U403 (N_403,In_511,In_327);
or U404 (N_404,In_1998,In_155);
xor U405 (N_405,In_247,In_1792);
nand U406 (N_406,In_1408,In_494);
and U407 (N_407,In_24,In_847);
or U408 (N_408,In_442,In_1141);
nor U409 (N_409,In_471,In_1693);
xnor U410 (N_410,In_1475,In_1367);
xnor U411 (N_411,In_1828,In_124);
or U412 (N_412,In_1293,In_794);
nor U413 (N_413,In_76,In_951);
xnor U414 (N_414,In_499,In_1739);
nor U415 (N_415,In_933,In_811);
and U416 (N_416,In_125,In_315);
nand U417 (N_417,In_1976,In_1818);
or U418 (N_418,In_1222,In_1196);
nor U419 (N_419,In_419,In_1727);
xnor U420 (N_420,In_1446,In_1692);
xor U421 (N_421,In_459,In_1670);
nor U422 (N_422,In_677,In_528);
xor U423 (N_423,In_305,In_1835);
xnor U424 (N_424,In_796,In_660);
xnor U425 (N_425,In_1019,In_62);
and U426 (N_426,In_1585,In_437);
and U427 (N_427,In_364,In_1258);
nor U428 (N_428,In_1840,In_1548);
xor U429 (N_429,In_287,In_284);
and U430 (N_430,In_171,In_398);
nor U431 (N_431,In_199,In_251);
or U432 (N_432,In_1054,In_307);
and U433 (N_433,In_1926,In_178);
or U434 (N_434,In_1683,In_1059);
and U435 (N_435,In_1357,In_185);
xnor U436 (N_436,In_744,In_1529);
nor U437 (N_437,In_1274,In_992);
nor U438 (N_438,In_165,In_258);
nand U439 (N_439,In_1304,In_1964);
and U440 (N_440,In_945,In_1351);
nand U441 (N_441,In_1645,In_867);
and U442 (N_442,In_752,In_1135);
and U443 (N_443,In_117,In_380);
nand U444 (N_444,In_896,In_745);
or U445 (N_445,In_65,In_1482);
nand U446 (N_446,In_42,In_790);
nor U447 (N_447,In_1256,In_658);
nand U448 (N_448,In_1233,In_1431);
nor U449 (N_449,In_1338,In_1922);
xnor U450 (N_450,In_937,In_801);
and U451 (N_451,In_1411,In_647);
nor U452 (N_452,In_960,In_1283);
nor U453 (N_453,In_1159,In_599);
xor U454 (N_454,In_782,In_887);
nand U455 (N_455,In_242,In_1885);
nand U456 (N_456,In_575,In_128);
xnor U457 (N_457,In_1537,In_1631);
and U458 (N_458,In_1652,In_1890);
nand U459 (N_459,In_1108,In_1085);
nor U460 (N_460,In_1616,In_1269);
nor U461 (N_461,In_104,In_1372);
and U462 (N_462,In_560,In_1817);
and U463 (N_463,In_1759,In_776);
and U464 (N_464,In_1382,In_601);
or U465 (N_465,In_1507,In_674);
or U466 (N_466,In_1705,In_1837);
or U467 (N_467,In_1239,In_766);
xor U468 (N_468,In_1421,In_541);
xnor U469 (N_469,In_1766,In_1307);
nand U470 (N_470,In_922,In_626);
nand U471 (N_471,In_1323,In_112);
xnor U472 (N_472,In_789,In_1499);
nor U473 (N_473,In_806,In_931);
and U474 (N_474,In_1273,In_885);
nand U475 (N_475,In_273,In_1997);
nor U476 (N_476,In_173,In_1306);
and U477 (N_477,In_537,In_502);
or U478 (N_478,In_1836,In_512);
or U479 (N_479,In_809,In_1694);
nor U480 (N_480,In_1190,In_714);
nand U481 (N_481,In_193,In_141);
nand U482 (N_482,In_1243,In_576);
nand U483 (N_483,In_943,In_706);
and U484 (N_484,In_1379,In_1586);
nand U485 (N_485,In_876,In_871);
and U486 (N_486,In_61,In_201);
xnor U487 (N_487,In_787,In_181);
nand U488 (N_488,In_1144,In_1007);
xor U489 (N_489,In_608,In_773);
nand U490 (N_490,In_1051,In_487);
nor U491 (N_491,In_1582,In_827);
and U492 (N_492,In_1546,In_1006);
nor U493 (N_493,In_384,In_934);
and U494 (N_494,In_311,In_1723);
or U495 (N_495,In_1644,In_1732);
xnor U496 (N_496,In_1587,In_473);
and U497 (N_497,In_1272,In_1820);
or U498 (N_498,In_177,In_1650);
and U499 (N_499,In_96,In_500);
xor U500 (N_500,In_87,In_120);
xor U501 (N_501,In_1760,In_1343);
xor U502 (N_502,In_506,In_1569);
and U503 (N_503,In_1589,In_100);
xnor U504 (N_504,In_1602,In_336);
and U505 (N_505,In_1072,In_843);
xor U506 (N_506,In_1845,In_781);
nor U507 (N_507,In_1017,In_1663);
or U508 (N_508,In_1401,In_312);
xnor U509 (N_509,In_1469,In_543);
nor U510 (N_510,In_1405,In_1560);
nand U511 (N_511,In_949,In_633);
or U512 (N_512,In_418,In_1574);
nor U513 (N_513,In_849,In_906);
or U514 (N_514,In_1744,In_374);
or U515 (N_515,In_1526,In_1973);
nand U516 (N_516,In_1841,In_1174);
xnor U517 (N_517,In_1311,In_942);
and U518 (N_518,In_237,In_1784);
and U519 (N_519,In_627,In_1591);
nand U520 (N_520,In_153,In_161);
and U521 (N_521,In_1832,In_857);
and U522 (N_522,In_603,In_1248);
and U523 (N_523,In_38,In_1033);
and U524 (N_524,In_1309,In_722);
nand U525 (N_525,In_1147,In_152);
and U526 (N_526,In_852,In_1859);
and U527 (N_527,In_595,In_93);
xnor U528 (N_528,In_1661,In_1266);
nand U529 (N_529,In_230,In_1129);
or U530 (N_530,In_427,In_667);
xnor U531 (N_531,In_365,In_441);
xnor U532 (N_532,In_826,In_1428);
nand U533 (N_533,In_619,In_1665);
or U534 (N_534,In_1627,In_1361);
nand U535 (N_535,In_1415,In_1985);
xor U536 (N_536,In_532,In_1014);
or U537 (N_537,In_850,In_1368);
and U538 (N_538,In_373,In_257);
nand U539 (N_539,In_428,In_1228);
nor U540 (N_540,In_1278,In_1493);
xnor U541 (N_541,In_1121,In_1594);
nand U542 (N_542,In_276,In_1884);
xor U543 (N_543,In_1308,In_1300);
nor U544 (N_544,In_1793,In_614);
xnor U545 (N_545,In_1,In_613);
nand U546 (N_546,In_1191,In_50);
nor U547 (N_547,In_703,In_1909);
nand U548 (N_548,In_1941,In_1576);
and U549 (N_549,In_301,In_1312);
and U550 (N_550,In_759,In_1902);
nand U551 (N_551,In_435,In_413);
or U552 (N_552,In_375,In_288);
or U553 (N_553,In_1275,In_1520);
xnor U554 (N_554,In_485,In_1714);
nand U555 (N_555,In_1241,In_369);
nor U556 (N_556,In_1782,In_859);
xor U557 (N_557,In_1463,In_1947);
or U558 (N_558,In_644,In_89);
nand U559 (N_559,In_132,In_1904);
nand U560 (N_560,In_720,In_82);
or U561 (N_561,In_712,In_731);
or U562 (N_562,In_1419,In_634);
nor U563 (N_563,In_1289,In_1659);
or U564 (N_564,In_835,In_1458);
xnor U565 (N_565,In_5,In_1235);
nand U566 (N_566,In_35,In_1148);
and U567 (N_567,In_1609,In_1154);
nor U568 (N_568,In_1750,In_453);
xnor U569 (N_569,In_980,In_1741);
and U570 (N_570,In_186,In_1249);
xnor U571 (N_571,In_968,In_1555);
and U572 (N_572,In_1717,In_118);
nor U573 (N_573,In_630,In_1878);
nor U574 (N_574,In_1834,In_596);
or U575 (N_575,In_1676,In_1915);
nor U576 (N_576,In_1721,In_542);
nor U577 (N_577,In_844,In_1613);
nand U578 (N_578,In_904,In_460);
and U579 (N_579,In_280,In_1653);
or U580 (N_580,In_1952,In_700);
or U581 (N_581,In_97,In_953);
or U582 (N_582,In_1509,In_1738);
or U583 (N_583,In_1622,In_1286);
nand U584 (N_584,In_1951,In_344);
nand U585 (N_585,In_1483,In_1435);
xnor U586 (N_586,In_1684,In_1277);
nor U587 (N_587,In_1257,In_1908);
nand U588 (N_588,In_1519,In_804);
nand U589 (N_589,In_697,In_875);
nand U590 (N_590,In_1706,In_140);
nor U591 (N_591,In_522,In_947);
nor U592 (N_592,In_1550,In_890);
xor U593 (N_593,In_1424,In_1551);
nand U594 (N_594,In_819,In_1833);
or U595 (N_595,In_1175,In_998);
and U596 (N_596,In_1185,In_329);
and U597 (N_597,In_1701,In_993);
nor U598 (N_598,In_229,In_1557);
xnor U599 (N_599,In_1877,In_881);
nor U600 (N_600,In_184,In_1987);
nor U601 (N_601,In_33,In_1477);
and U602 (N_602,In_1503,In_1671);
nand U603 (N_603,In_1673,In_1528);
or U604 (N_604,In_1460,In_1977);
nand U605 (N_605,In_1225,In_227);
nor U606 (N_606,In_74,In_53);
nand U607 (N_607,In_310,In_70);
xor U608 (N_608,In_615,In_1034);
or U609 (N_609,In_1763,In_339);
and U610 (N_610,In_817,In_1742);
nor U611 (N_611,In_921,In_370);
xnor U612 (N_612,In_79,In_188);
xnor U613 (N_613,In_1402,In_648);
nor U614 (N_614,In_1768,In_245);
xor U615 (N_615,In_939,In_902);
xor U616 (N_616,In_1318,In_1984);
xor U617 (N_617,In_385,In_1606);
nand U618 (N_618,In_1610,In_916);
or U619 (N_619,In_1140,In_1083);
and U620 (N_620,In_122,In_1822);
and U621 (N_621,In_137,In_168);
nand U622 (N_622,In_862,In_216);
nand U623 (N_623,In_1876,In_1687);
and U624 (N_624,In_1400,In_469);
or U625 (N_625,In_1168,In_1394);
nor U626 (N_626,In_1305,In_1391);
xnor U627 (N_627,In_1959,In_1195);
nor U628 (N_628,In_1077,In_1531);
or U629 (N_629,In_1912,In_1448);
or U630 (N_630,In_1350,In_1814);
nand U631 (N_631,In_266,In_371);
nand U632 (N_632,In_785,In_1333);
nand U633 (N_633,In_903,In_1547);
xor U634 (N_634,In_840,In_1695);
xnor U635 (N_635,In_1944,In_1858);
or U636 (N_636,In_368,In_468);
or U637 (N_637,In_1003,In_1558);
nand U638 (N_638,In_959,In_157);
nor U639 (N_639,In_1326,In_1510);
or U640 (N_640,In_523,In_657);
or U641 (N_641,In_1881,In_1900);
nand U642 (N_642,In_0,In_248);
and U643 (N_643,In_1737,In_255);
and U644 (N_644,In_345,In_1164);
nand U645 (N_645,In_1008,In_1383);
nand U646 (N_646,In_1282,In_71);
nor U647 (N_647,In_1029,In_547);
xnor U648 (N_648,In_10,In_1231);
and U649 (N_649,In_1189,In_1166);
and U650 (N_650,In_291,In_985);
and U651 (N_651,In_461,In_779);
nand U652 (N_652,In_1001,In_401);
xnor U653 (N_653,In_1815,In_1111);
nor U654 (N_654,In_756,In_1983);
nand U655 (N_655,In_1120,In_1271);
nor U656 (N_656,In_421,In_693);
xor U657 (N_657,In_498,In_1023);
or U658 (N_658,In_1620,In_1265);
and U659 (N_659,In_431,In_1197);
xor U660 (N_660,In_289,In_663);
nand U661 (N_661,In_578,In_1808);
and U662 (N_662,In_445,In_504);
nand U663 (N_663,In_1895,In_841);
nand U664 (N_664,In_1441,In_1112);
nor U665 (N_665,In_331,In_1796);
and U666 (N_666,In_323,In_1332);
xor U667 (N_667,In_1026,In_443);
xor U668 (N_668,In_777,In_1608);
nor U669 (N_669,In_842,In_1588);
nor U670 (N_670,In_379,In_182);
and U671 (N_671,In_1580,In_709);
nand U672 (N_672,In_878,In_1566);
and U673 (N_673,In_1396,In_1353);
nor U674 (N_674,In_203,In_1734);
nand U675 (N_675,In_232,In_1060);
or U676 (N_676,In_683,In_28);
xor U677 (N_677,In_1880,In_1762);
and U678 (N_678,In_198,In_493);
nor U679 (N_679,In_1134,In_297);
nor U680 (N_680,In_1747,In_651);
nand U681 (N_681,In_372,In_1982);
nor U682 (N_682,In_687,In_778);
or U683 (N_683,In_969,In_562);
xor U684 (N_684,In_642,In_1119);
and U685 (N_685,In_1439,In_1662);
nor U686 (N_686,In_1092,In_1202);
and U687 (N_687,In_1797,In_1207);
nand U688 (N_688,In_925,In_1899);
and U689 (N_689,In_1025,In_1122);
nand U690 (N_690,In_1931,In_1217);
nand U691 (N_691,In_836,In_1632);
nor U692 (N_692,In_450,In_1057);
and U693 (N_693,In_455,In_1027);
xor U694 (N_694,In_1758,In_1244);
nand U695 (N_695,In_233,In_1533);
and U696 (N_696,In_1288,In_350);
xnor U697 (N_697,In_1230,In_733);
or U698 (N_698,In_1700,In_1128);
xnor U699 (N_699,In_1935,In_269);
or U700 (N_700,In_1261,In_1674);
or U701 (N_701,In_211,In_1898);
nand U702 (N_702,In_1639,In_11);
nor U703 (N_703,In_585,In_1543);
and U704 (N_704,In_1301,In_1993);
and U705 (N_705,In_914,In_1685);
nor U706 (N_706,In_898,In_1810);
nand U707 (N_707,In_1807,In_25);
xnor U708 (N_708,In_481,In_1176);
nand U709 (N_709,In_144,In_1434);
nor U710 (N_710,In_1444,In_1100);
xnor U711 (N_711,In_1151,In_84);
or U712 (N_712,In_1179,In_1362);
or U713 (N_713,In_1253,In_689);
nand U714 (N_714,In_1669,In_564);
or U715 (N_715,In_1086,In_825);
or U716 (N_716,In_464,In_1096);
nor U717 (N_717,In_1517,In_721);
or U718 (N_718,In_1490,In_1923);
nor U719 (N_719,In_710,In_788);
and U720 (N_720,In_136,In_358);
nand U721 (N_721,In_1868,In_1857);
xnor U722 (N_722,In_1856,In_769);
nand U723 (N_723,In_206,In_63);
xor U724 (N_724,In_243,In_1345);
xnor U725 (N_725,In_399,In_833);
nor U726 (N_726,In_735,In_264);
nor U727 (N_727,In_1038,In_1925);
and U728 (N_728,In_592,In_1284);
nand U729 (N_729,In_1182,In_1879);
or U730 (N_730,In_1080,In_805);
and U731 (N_731,In_1962,In_381);
xor U732 (N_732,In_909,In_359);
or U733 (N_733,In_918,In_1035);
and U734 (N_734,In_1088,In_1436);
xor U735 (N_735,In_686,In_1292);
and U736 (N_736,In_972,In_160);
xnor U737 (N_737,In_1316,In_294);
xor U738 (N_738,In_1042,In_1798);
or U739 (N_739,In_1479,In_983);
or U740 (N_740,In_1789,In_646);
and U741 (N_741,In_1617,In_436);
xnor U742 (N_742,In_524,In_1624);
nor U743 (N_743,In_1336,In_167);
nor U744 (N_744,In_1956,In_77);
and U745 (N_745,In_228,In_48);
nor U746 (N_746,In_907,In_681);
xnor U747 (N_747,In_1514,In_221);
nand U748 (N_748,In_1113,In_1062);
or U749 (N_749,In_1251,In_556);
nand U750 (N_750,In_18,In_1839);
and U751 (N_751,In_92,In_1331);
xor U752 (N_752,In_573,In_832);
nor U753 (N_753,In_1417,In_1178);
nor U754 (N_754,In_1459,In_1824);
and U755 (N_755,In_166,In_1638);
nand U756 (N_756,In_1452,In_1491);
or U757 (N_757,In_414,In_353);
or U758 (N_758,In_109,In_1381);
or U759 (N_759,In_477,In_466);
nand U760 (N_760,In_126,In_1953);
or U761 (N_761,In_1145,In_12);
nand U762 (N_762,In_901,In_823);
nand U763 (N_763,In_438,In_432);
and U764 (N_764,In_639,In_879);
nand U765 (N_765,In_154,In_618);
nand U766 (N_766,In_1418,In_1770);
and U767 (N_767,In_738,In_281);
nor U768 (N_768,In_121,In_1438);
and U769 (N_769,In_308,In_964);
and U770 (N_770,In_298,In_482);
and U771 (N_771,In_1979,In_1021);
nor U772 (N_772,In_624,In_1809);
or U773 (N_773,In_1192,In_271);
or U774 (N_774,In_848,In_1068);
and U775 (N_775,In_1772,In_780);
nor U776 (N_776,In_726,In_1392);
or U777 (N_777,In_409,In_1018);
nand U778 (N_778,In_1470,In_551);
and U779 (N_779,In_952,In_1171);
nor U780 (N_780,In_16,In_999);
nand U781 (N_781,In_1992,In_1355);
and U782 (N_782,In_1101,In_598);
xnor U783 (N_783,In_610,In_1785);
or U784 (N_784,In_40,In_1209);
nor U785 (N_785,In_870,In_698);
nor U786 (N_786,In_1934,In_1649);
or U787 (N_787,In_886,In_1561);
or U788 (N_788,In_1440,In_1127);
nor U789 (N_789,In_591,In_1625);
nor U790 (N_790,In_1924,In_775);
or U791 (N_791,In_496,In_1369);
xnor U792 (N_792,In_606,In_37);
xor U793 (N_793,In_1771,In_928);
nor U794 (N_794,In_629,In_741);
and U795 (N_795,In_1360,In_1812);
nor U796 (N_796,In_550,In_1453);
nand U797 (N_797,In_1187,In_1211);
or U798 (N_798,In_1699,In_200);
xor U799 (N_799,In_1188,In_1352);
and U800 (N_800,In_670,In_529);
xnor U801 (N_801,In_208,In_142);
nand U802 (N_802,In_664,In_139);
nor U803 (N_803,In_356,In_1894);
or U804 (N_804,In_861,In_590);
or U805 (N_805,In_1107,In_569);
nor U806 (N_806,In_205,In_434);
xor U807 (N_807,In_1497,In_214);
and U808 (N_808,In_1708,In_1563);
xor U809 (N_809,In_1910,In_1281);
nand U810 (N_810,In_1678,In_1578);
nor U811 (N_811,In_1240,In_510);
and U812 (N_812,In_1751,In_936);
nand U813 (N_813,In_1648,In_748);
nor U814 (N_814,In_938,In_8);
and U815 (N_815,In_103,In_1030);
and U816 (N_816,In_403,In_873);
and U817 (N_817,In_349,In_655);
or U818 (N_818,In_1322,In_1769);
xor U819 (N_819,In_1535,In_279);
and U820 (N_820,In_584,In_973);
nand U821 (N_821,In_662,In_1621);
xnor U822 (N_822,In_1991,In_1106);
nand U823 (N_823,In_1359,In_877);
and U824 (N_824,In_1567,In_1177);
or U825 (N_825,In_1553,In_679);
nor U826 (N_826,In_1046,In_1000);
and U827 (N_827,In_866,In_147);
and U828 (N_828,In_1201,In_29);
or U829 (N_829,In_1432,In_277);
nand U830 (N_830,In_1407,In_1518);
nand U831 (N_831,In_519,In_1084);
nor U832 (N_832,In_829,In_654);
xor U833 (N_833,In_1041,In_1081);
nand U834 (N_834,In_492,In_1615);
and U835 (N_835,In_215,In_1651);
nor U836 (N_836,In_920,In_1677);
xor U837 (N_837,In_465,In_1786);
nand U838 (N_838,In_814,In_360);
nand U839 (N_839,In_1137,In_1053);
and U840 (N_840,In_894,In_1290);
or U841 (N_841,In_1612,In_996);
nor U842 (N_842,In_1932,In_856);
and U843 (N_843,In_1722,In_1565);
nor U844 (N_844,In_717,In_516);
xor U845 (N_845,In_517,In_1133);
nand U846 (N_846,In_1525,In_783);
or U847 (N_847,In_1374,In_1948);
nor U848 (N_848,In_224,In_15);
or U849 (N_849,In_1861,In_1198);
and U850 (N_850,In_555,In_1752);
xnor U851 (N_851,In_1380,In_1377);
or U852 (N_852,In_813,In_472);
and U853 (N_853,In_1579,In_889);
xnor U854 (N_854,In_299,In_56);
nor U855 (N_855,In_1583,In_338);
nor U856 (N_856,In_133,In_383);
nor U857 (N_857,In_1968,In_802);
and U858 (N_858,In_241,In_31);
or U859 (N_859,In_581,In_1914);
nor U860 (N_860,In_1476,In_404);
nor U861 (N_861,In_915,In_1247);
or U862 (N_862,In_1016,In_452);
xor U863 (N_863,In_1827,In_1131);
or U864 (N_864,In_21,In_1043);
nor U865 (N_865,In_1310,In_602);
nor U866 (N_866,In_1696,In_702);
or U867 (N_867,In_179,In_1325);
xnor U868 (N_868,In_138,In_1221);
and U869 (N_869,In_1802,In_47);
and U870 (N_870,In_1703,In_1399);
nand U871 (N_871,In_1342,In_1672);
or U872 (N_872,In_1075,In_1590);
xor U873 (N_873,In_1040,In_1366);
nand U874 (N_874,In_1024,In_1155);
or U875 (N_875,In_99,In_1754);
nand U876 (N_876,In_1031,In_1605);
nand U877 (N_877,In_334,In_865);
nor U878 (N_878,In_1393,In_803);
nand U879 (N_879,In_1978,In_1093);
nand U880 (N_880,In_347,In_1346);
and U881 (N_881,In_1420,In_1063);
or U882 (N_882,In_1918,In_1564);
xor U883 (N_883,In_1892,In_98);
or U884 (N_884,In_106,In_1186);
nor U885 (N_885,In_393,In_963);
nor U886 (N_886,In_554,In_665);
nand U887 (N_887,In_483,In_1330);
nor U888 (N_888,In_387,In_406);
or U889 (N_889,In_1488,In_770);
or U890 (N_890,In_1206,In_957);
or U891 (N_891,In_1437,In_989);
and U892 (N_892,In_1642,In_1110);
and U893 (N_893,In_83,In_820);
nor U894 (N_894,In_4,In_743);
nand U895 (N_895,In_1009,In_1929);
xor U896 (N_896,In_625,In_678);
or U897 (N_897,In_559,In_1214);
nor U898 (N_898,In_944,In_1521);
or U899 (N_899,In_536,In_1181);
xor U900 (N_900,In_1730,In_1633);
or U901 (N_901,In_1210,In_690);
nor U902 (N_902,In_962,In_176);
nor U903 (N_903,In_363,In_834);
nand U904 (N_904,In_68,In_1848);
nor U905 (N_905,In_1637,In_1114);
nand U906 (N_906,In_1972,In_696);
nand U907 (N_907,In_673,In_893);
and U908 (N_908,In_1433,In_219);
and U909 (N_909,In_58,In_107);
and U910 (N_910,In_1536,In_1611);
and U911 (N_911,In_1302,In_1854);
or U912 (N_912,In_557,In_917);
or U913 (N_913,In_1930,In_1969);
or U914 (N_914,In_732,In_1646);
nor U915 (N_915,In_1949,In_1515);
or U916 (N_916,In_830,In_1136);
and U917 (N_917,In_699,In_1242);
nor U918 (N_918,In_300,In_1783);
or U919 (N_919,In_1940,In_1795);
nand U920 (N_920,In_1846,In_791);
or U921 (N_921,In_593,In_41);
nor U922 (N_922,In_1315,In_888);
nand U923 (N_923,In_389,In_1153);
or U924 (N_924,In_402,In_553);
xor U925 (N_925,In_209,In_961);
xnor U926 (N_926,In_1888,In_1303);
or U927 (N_927,In_332,In_1911);
xor U928 (N_928,In_1055,In_1619);
nor U929 (N_929,In_1478,In_1549);
xnor U930 (N_930,In_656,In_1297);
nand U931 (N_931,In_932,In_1387);
nand U932 (N_932,In_652,In_1778);
or U933 (N_933,In_1889,In_640);
nand U934 (N_934,In_579,In_958);
xor U935 (N_935,In_1697,In_1728);
nor U936 (N_936,In_514,In_1486);
xnor U937 (N_937,In_439,In_486);
nor U938 (N_938,In_1364,In_795);
nor U939 (N_939,In_367,In_740);
nand U940 (N_940,In_1328,In_86);
xnor U941 (N_941,In_718,In_1015);
xor U942 (N_942,In_1203,In_1597);
nor U943 (N_943,In_1757,In_1623);
or U944 (N_944,In_1010,In_1575);
or U945 (N_945,In_1037,In_1511);
xnor U946 (N_946,In_1502,In_1157);
or U947 (N_947,In_45,In_1614);
nor U948 (N_948,In_75,In_1416);
xnor U949 (N_949,In_753,In_1937);
nand U950 (N_950,In_1327,In_163);
nand U951 (N_951,In_1022,In_1454);
and U952 (N_952,In_1193,In_148);
nor U953 (N_953,In_1599,In_1254);
or U954 (N_954,In_950,In_263);
and U955 (N_955,In_1404,In_1194);
nand U956 (N_956,In_1067,In_1074);
nor U957 (N_957,In_605,In_1989);
xor U958 (N_958,In_1655,In_1743);
xnor U959 (N_959,In_1071,In_1103);
nor U960 (N_960,In_666,In_1577);
nor U961 (N_961,In_984,In_476);
and U962 (N_962,In_39,In_1691);
or U963 (N_963,In_1234,In_650);
xor U964 (N_964,In_583,In_1647);
xor U965 (N_965,In_1250,In_1544);
or U966 (N_966,In_1559,In_1656);
and U967 (N_967,In_1089,In_1592);
nand U968 (N_968,In_420,In_1584);
or U969 (N_969,In_1552,In_306);
and U970 (N_970,In_1169,In_1255);
nor U971 (N_971,In_1498,In_131);
nand U972 (N_972,In_433,In_1276);
nor U973 (N_973,In_1170,In_1872);
and U974 (N_974,In_328,In_1078);
or U975 (N_975,In_225,In_260);
or U976 (N_976,In_727,In_818);
xor U977 (N_977,In_982,In_659);
nand U978 (N_978,In_822,In_765);
nand U979 (N_979,In_1830,In_545);
and U980 (N_980,In_1852,In_580);
and U981 (N_981,In_170,In_739);
xnor U982 (N_982,In_313,In_824);
xor U983 (N_983,In_1245,In_1988);
nor U984 (N_984,In_1403,In_1601);
or U985 (N_985,In_1165,In_195);
and U986 (N_986,In_594,In_1335);
xnor U987 (N_987,In_491,In_1004);
or U988 (N_988,In_362,In_1680);
nand U989 (N_989,In_1887,In_1048);
xnor U990 (N_990,In_930,In_1020);
or U991 (N_991,In_1449,In_821);
or U992 (N_992,In_1767,In_1398);
and U993 (N_993,In_123,In_668);
and U994 (N_994,In_688,In_1160);
nor U995 (N_995,In_535,In_645);
nor U996 (N_996,In_872,In_1933);
and U997 (N_997,In_1874,In_1527);
xor U998 (N_998,In_1138,In_52);
and U999 (N_999,In_36,In_786);
and U1000 (N_1000,In_1676,In_942);
and U1001 (N_1001,In_748,In_1035);
or U1002 (N_1002,In_35,In_438);
xor U1003 (N_1003,In_1206,In_50);
nand U1004 (N_1004,In_1399,In_757);
and U1005 (N_1005,In_1412,In_848);
xor U1006 (N_1006,In_660,In_593);
and U1007 (N_1007,In_125,In_1531);
nor U1008 (N_1008,In_867,In_840);
or U1009 (N_1009,In_1228,In_1611);
nor U1010 (N_1010,In_1037,In_553);
nor U1011 (N_1011,In_730,In_969);
or U1012 (N_1012,In_1291,In_618);
nand U1013 (N_1013,In_1287,In_388);
or U1014 (N_1014,In_1372,In_413);
nor U1015 (N_1015,In_1676,In_1408);
xnor U1016 (N_1016,In_990,In_20);
nor U1017 (N_1017,In_1337,In_891);
nor U1018 (N_1018,In_1828,In_1985);
nand U1019 (N_1019,In_1205,In_44);
nor U1020 (N_1020,In_945,In_1566);
xnor U1021 (N_1021,In_768,In_1327);
and U1022 (N_1022,In_646,In_187);
nand U1023 (N_1023,In_1421,In_1915);
and U1024 (N_1024,In_1764,In_561);
xnor U1025 (N_1025,In_1395,In_1616);
xnor U1026 (N_1026,In_1996,In_470);
nor U1027 (N_1027,In_13,In_1027);
nand U1028 (N_1028,In_194,In_450);
nor U1029 (N_1029,In_1181,In_413);
and U1030 (N_1030,In_421,In_56);
xnor U1031 (N_1031,In_1163,In_454);
nor U1032 (N_1032,In_970,In_192);
nand U1033 (N_1033,In_618,In_1161);
nor U1034 (N_1034,In_817,In_933);
and U1035 (N_1035,In_185,In_1523);
nor U1036 (N_1036,In_484,In_1108);
or U1037 (N_1037,In_115,In_581);
or U1038 (N_1038,In_1399,In_834);
xnor U1039 (N_1039,In_875,In_1509);
nand U1040 (N_1040,In_1891,In_1378);
nor U1041 (N_1041,In_1043,In_1027);
nor U1042 (N_1042,In_646,In_1219);
xnor U1043 (N_1043,In_884,In_156);
xnor U1044 (N_1044,In_593,In_1260);
nor U1045 (N_1045,In_1160,In_592);
nand U1046 (N_1046,In_1870,In_1264);
nor U1047 (N_1047,In_698,In_1740);
or U1048 (N_1048,In_738,In_32);
or U1049 (N_1049,In_604,In_406);
nor U1050 (N_1050,In_70,In_702);
nand U1051 (N_1051,In_764,In_644);
or U1052 (N_1052,In_1805,In_1917);
or U1053 (N_1053,In_132,In_1168);
and U1054 (N_1054,In_819,In_424);
nor U1055 (N_1055,In_626,In_484);
or U1056 (N_1056,In_1029,In_1069);
and U1057 (N_1057,In_801,In_1522);
or U1058 (N_1058,In_1797,In_142);
xnor U1059 (N_1059,In_1090,In_583);
or U1060 (N_1060,In_364,In_765);
or U1061 (N_1061,In_180,In_521);
xor U1062 (N_1062,In_1565,In_659);
or U1063 (N_1063,In_1341,In_14);
and U1064 (N_1064,In_1778,In_794);
nand U1065 (N_1065,In_1261,In_505);
xor U1066 (N_1066,In_1497,In_741);
xor U1067 (N_1067,In_523,In_157);
xnor U1068 (N_1068,In_682,In_177);
and U1069 (N_1069,In_1866,In_1822);
and U1070 (N_1070,In_1576,In_309);
nor U1071 (N_1071,In_1631,In_381);
or U1072 (N_1072,In_1086,In_1035);
nand U1073 (N_1073,In_1543,In_462);
or U1074 (N_1074,In_1070,In_765);
or U1075 (N_1075,In_1545,In_201);
and U1076 (N_1076,In_1247,In_1804);
nand U1077 (N_1077,In_1087,In_397);
or U1078 (N_1078,In_1964,In_74);
nand U1079 (N_1079,In_828,In_9);
nor U1080 (N_1080,In_285,In_1180);
or U1081 (N_1081,In_298,In_329);
nand U1082 (N_1082,In_348,In_286);
or U1083 (N_1083,In_380,In_1937);
and U1084 (N_1084,In_273,In_1077);
nor U1085 (N_1085,In_523,In_1439);
nor U1086 (N_1086,In_1287,In_569);
or U1087 (N_1087,In_1152,In_107);
and U1088 (N_1088,In_999,In_1812);
or U1089 (N_1089,In_137,In_1217);
or U1090 (N_1090,In_1172,In_309);
xnor U1091 (N_1091,In_1700,In_768);
nor U1092 (N_1092,In_660,In_1940);
or U1093 (N_1093,In_438,In_1887);
or U1094 (N_1094,In_821,In_1082);
nor U1095 (N_1095,In_1532,In_386);
nand U1096 (N_1096,In_170,In_1095);
nor U1097 (N_1097,In_1109,In_1730);
or U1098 (N_1098,In_1495,In_938);
xor U1099 (N_1099,In_1591,In_1320);
and U1100 (N_1100,In_806,In_691);
or U1101 (N_1101,In_1824,In_793);
and U1102 (N_1102,In_303,In_1800);
xnor U1103 (N_1103,In_478,In_176);
or U1104 (N_1104,In_457,In_1813);
nand U1105 (N_1105,In_52,In_1093);
or U1106 (N_1106,In_1391,In_927);
xor U1107 (N_1107,In_1837,In_2);
xor U1108 (N_1108,In_1656,In_1421);
or U1109 (N_1109,In_1447,In_1610);
nor U1110 (N_1110,In_1298,In_1546);
xnor U1111 (N_1111,In_1591,In_57);
xnor U1112 (N_1112,In_135,In_284);
or U1113 (N_1113,In_66,In_324);
nand U1114 (N_1114,In_260,In_1833);
or U1115 (N_1115,In_280,In_633);
and U1116 (N_1116,In_667,In_366);
and U1117 (N_1117,In_1817,In_1666);
and U1118 (N_1118,In_1455,In_139);
xor U1119 (N_1119,In_1074,In_173);
nor U1120 (N_1120,In_15,In_558);
and U1121 (N_1121,In_710,In_1231);
xnor U1122 (N_1122,In_1948,In_536);
nor U1123 (N_1123,In_530,In_1786);
nor U1124 (N_1124,In_110,In_1364);
or U1125 (N_1125,In_1314,In_1235);
or U1126 (N_1126,In_1488,In_584);
xor U1127 (N_1127,In_1137,In_900);
or U1128 (N_1128,In_129,In_354);
or U1129 (N_1129,In_1962,In_960);
and U1130 (N_1130,In_1195,In_1141);
or U1131 (N_1131,In_229,In_988);
nor U1132 (N_1132,In_922,In_308);
xor U1133 (N_1133,In_568,In_1354);
and U1134 (N_1134,In_1355,In_1362);
or U1135 (N_1135,In_890,In_1209);
nand U1136 (N_1136,In_1335,In_1124);
or U1137 (N_1137,In_1517,In_149);
nor U1138 (N_1138,In_1247,In_926);
and U1139 (N_1139,In_648,In_449);
and U1140 (N_1140,In_1217,In_1535);
and U1141 (N_1141,In_456,In_879);
or U1142 (N_1142,In_20,In_584);
and U1143 (N_1143,In_977,In_1806);
and U1144 (N_1144,In_1176,In_273);
nand U1145 (N_1145,In_630,In_1200);
and U1146 (N_1146,In_1309,In_634);
and U1147 (N_1147,In_1351,In_1623);
nand U1148 (N_1148,In_154,In_285);
nor U1149 (N_1149,In_1016,In_653);
nor U1150 (N_1150,In_680,In_337);
xor U1151 (N_1151,In_401,In_1797);
nand U1152 (N_1152,In_1693,In_646);
nand U1153 (N_1153,In_1139,In_267);
or U1154 (N_1154,In_1785,In_96);
nor U1155 (N_1155,In_658,In_473);
and U1156 (N_1156,In_838,In_166);
or U1157 (N_1157,In_1065,In_1539);
nand U1158 (N_1158,In_777,In_638);
nand U1159 (N_1159,In_1181,In_289);
xnor U1160 (N_1160,In_683,In_1945);
nand U1161 (N_1161,In_1078,In_94);
or U1162 (N_1162,In_1905,In_1869);
or U1163 (N_1163,In_1316,In_632);
nor U1164 (N_1164,In_1468,In_1124);
and U1165 (N_1165,In_818,In_1998);
nor U1166 (N_1166,In_1462,In_245);
nand U1167 (N_1167,In_1704,In_1802);
xor U1168 (N_1168,In_926,In_1045);
and U1169 (N_1169,In_292,In_714);
nor U1170 (N_1170,In_880,In_1636);
nor U1171 (N_1171,In_1638,In_85);
nor U1172 (N_1172,In_1701,In_1339);
and U1173 (N_1173,In_452,In_1574);
and U1174 (N_1174,In_882,In_1117);
nand U1175 (N_1175,In_679,In_856);
and U1176 (N_1176,In_747,In_1857);
or U1177 (N_1177,In_1472,In_1316);
nor U1178 (N_1178,In_1078,In_886);
or U1179 (N_1179,In_582,In_770);
and U1180 (N_1180,In_101,In_806);
or U1181 (N_1181,In_1720,In_1985);
nand U1182 (N_1182,In_88,In_1953);
xnor U1183 (N_1183,In_73,In_1773);
xnor U1184 (N_1184,In_293,In_107);
and U1185 (N_1185,In_1392,In_1957);
nor U1186 (N_1186,In_1225,In_459);
or U1187 (N_1187,In_1142,In_383);
nor U1188 (N_1188,In_87,In_1224);
nand U1189 (N_1189,In_1095,In_850);
or U1190 (N_1190,In_1416,In_663);
xor U1191 (N_1191,In_1201,In_495);
nor U1192 (N_1192,In_1590,In_1343);
nor U1193 (N_1193,In_1287,In_943);
xor U1194 (N_1194,In_1119,In_1424);
xnor U1195 (N_1195,In_1461,In_503);
xnor U1196 (N_1196,In_1787,In_228);
nor U1197 (N_1197,In_506,In_629);
nor U1198 (N_1198,In_1340,In_460);
xnor U1199 (N_1199,In_164,In_637);
xnor U1200 (N_1200,In_1883,In_1428);
and U1201 (N_1201,In_1604,In_576);
or U1202 (N_1202,In_1177,In_1061);
or U1203 (N_1203,In_1311,In_639);
or U1204 (N_1204,In_1854,In_587);
nor U1205 (N_1205,In_998,In_1414);
and U1206 (N_1206,In_1589,In_887);
nor U1207 (N_1207,In_211,In_20);
xnor U1208 (N_1208,In_1374,In_1272);
or U1209 (N_1209,In_1133,In_442);
xor U1210 (N_1210,In_1096,In_1299);
nor U1211 (N_1211,In_1899,In_1554);
and U1212 (N_1212,In_1890,In_1956);
nand U1213 (N_1213,In_969,In_122);
or U1214 (N_1214,In_68,In_1279);
nor U1215 (N_1215,In_124,In_996);
xnor U1216 (N_1216,In_232,In_736);
or U1217 (N_1217,In_870,In_1191);
and U1218 (N_1218,In_1143,In_389);
or U1219 (N_1219,In_604,In_712);
nand U1220 (N_1220,In_1780,In_1894);
nor U1221 (N_1221,In_254,In_249);
and U1222 (N_1222,In_443,In_71);
nor U1223 (N_1223,In_85,In_1151);
and U1224 (N_1224,In_237,In_1397);
xor U1225 (N_1225,In_1175,In_1764);
and U1226 (N_1226,In_513,In_520);
or U1227 (N_1227,In_1244,In_1370);
nor U1228 (N_1228,In_221,In_252);
nor U1229 (N_1229,In_1681,In_1559);
nand U1230 (N_1230,In_203,In_50);
nor U1231 (N_1231,In_239,In_775);
and U1232 (N_1232,In_786,In_258);
nor U1233 (N_1233,In_1239,In_172);
nand U1234 (N_1234,In_1810,In_118);
and U1235 (N_1235,In_1622,In_880);
or U1236 (N_1236,In_272,In_1453);
or U1237 (N_1237,In_1978,In_1012);
and U1238 (N_1238,In_375,In_415);
or U1239 (N_1239,In_1472,In_1034);
and U1240 (N_1240,In_182,In_108);
or U1241 (N_1241,In_595,In_1154);
or U1242 (N_1242,In_1003,In_1352);
or U1243 (N_1243,In_1333,In_908);
nand U1244 (N_1244,In_37,In_558);
nand U1245 (N_1245,In_1156,In_457);
nor U1246 (N_1246,In_1364,In_656);
xor U1247 (N_1247,In_530,In_998);
xnor U1248 (N_1248,In_604,In_1635);
xor U1249 (N_1249,In_1576,In_462);
nand U1250 (N_1250,In_1711,In_1601);
xnor U1251 (N_1251,In_1606,In_549);
xnor U1252 (N_1252,In_1741,In_1359);
and U1253 (N_1253,In_1267,In_1321);
xnor U1254 (N_1254,In_1642,In_64);
nor U1255 (N_1255,In_1122,In_1337);
or U1256 (N_1256,In_744,In_1989);
xor U1257 (N_1257,In_381,In_1657);
nand U1258 (N_1258,In_1000,In_1455);
xnor U1259 (N_1259,In_1286,In_1198);
or U1260 (N_1260,In_1746,In_1898);
or U1261 (N_1261,In_1558,In_1309);
nor U1262 (N_1262,In_171,In_1569);
nand U1263 (N_1263,In_829,In_1688);
nand U1264 (N_1264,In_1949,In_1985);
or U1265 (N_1265,In_1474,In_331);
nor U1266 (N_1266,In_555,In_10);
xnor U1267 (N_1267,In_217,In_506);
nor U1268 (N_1268,In_1027,In_1955);
and U1269 (N_1269,In_811,In_1040);
nand U1270 (N_1270,In_1383,In_810);
or U1271 (N_1271,In_127,In_1279);
or U1272 (N_1272,In_991,In_226);
and U1273 (N_1273,In_728,In_1473);
nor U1274 (N_1274,In_729,In_1090);
nand U1275 (N_1275,In_1199,In_1617);
and U1276 (N_1276,In_1194,In_475);
and U1277 (N_1277,In_847,In_1723);
nand U1278 (N_1278,In_1015,In_926);
or U1279 (N_1279,In_75,In_601);
and U1280 (N_1280,In_838,In_477);
nand U1281 (N_1281,In_1927,In_1895);
or U1282 (N_1282,In_492,In_1454);
or U1283 (N_1283,In_1612,In_169);
and U1284 (N_1284,In_251,In_1677);
nor U1285 (N_1285,In_1760,In_944);
nand U1286 (N_1286,In_452,In_1891);
nor U1287 (N_1287,In_1325,In_1991);
and U1288 (N_1288,In_816,In_319);
nand U1289 (N_1289,In_1147,In_255);
or U1290 (N_1290,In_1210,In_511);
nand U1291 (N_1291,In_832,In_73);
xnor U1292 (N_1292,In_1266,In_1190);
xnor U1293 (N_1293,In_1616,In_140);
xnor U1294 (N_1294,In_1406,In_104);
nor U1295 (N_1295,In_290,In_761);
or U1296 (N_1296,In_1948,In_1205);
nand U1297 (N_1297,In_1143,In_770);
or U1298 (N_1298,In_592,In_259);
nand U1299 (N_1299,In_1374,In_50);
nor U1300 (N_1300,In_7,In_1895);
nand U1301 (N_1301,In_1203,In_939);
and U1302 (N_1302,In_1406,In_1176);
and U1303 (N_1303,In_1650,In_487);
nor U1304 (N_1304,In_177,In_858);
xnor U1305 (N_1305,In_213,In_749);
nand U1306 (N_1306,In_1193,In_399);
or U1307 (N_1307,In_1122,In_1668);
or U1308 (N_1308,In_568,In_760);
xor U1309 (N_1309,In_923,In_1654);
nand U1310 (N_1310,In_1797,In_609);
nor U1311 (N_1311,In_843,In_378);
nor U1312 (N_1312,In_634,In_1248);
and U1313 (N_1313,In_81,In_520);
xnor U1314 (N_1314,In_1130,In_1819);
or U1315 (N_1315,In_1335,In_1741);
and U1316 (N_1316,In_880,In_1428);
nor U1317 (N_1317,In_306,In_324);
and U1318 (N_1318,In_428,In_1288);
nand U1319 (N_1319,In_1333,In_658);
and U1320 (N_1320,In_1009,In_592);
or U1321 (N_1321,In_1710,In_634);
or U1322 (N_1322,In_1876,In_300);
nand U1323 (N_1323,In_1580,In_860);
nand U1324 (N_1324,In_126,In_120);
or U1325 (N_1325,In_1715,In_718);
nor U1326 (N_1326,In_329,In_1766);
nor U1327 (N_1327,In_1411,In_1833);
or U1328 (N_1328,In_1221,In_560);
nand U1329 (N_1329,In_370,In_1747);
xnor U1330 (N_1330,In_1850,In_205);
nor U1331 (N_1331,In_1927,In_437);
xor U1332 (N_1332,In_583,In_1608);
xor U1333 (N_1333,In_811,In_713);
or U1334 (N_1334,In_475,In_872);
nor U1335 (N_1335,In_835,In_253);
nand U1336 (N_1336,In_172,In_119);
or U1337 (N_1337,In_917,In_689);
nand U1338 (N_1338,In_410,In_1072);
xor U1339 (N_1339,In_1637,In_1515);
nor U1340 (N_1340,In_230,In_1742);
or U1341 (N_1341,In_1985,In_396);
xor U1342 (N_1342,In_1687,In_790);
nand U1343 (N_1343,In_1611,In_743);
nor U1344 (N_1344,In_372,In_1831);
nand U1345 (N_1345,In_297,In_1743);
and U1346 (N_1346,In_404,In_1031);
xor U1347 (N_1347,In_413,In_329);
and U1348 (N_1348,In_372,In_1280);
nand U1349 (N_1349,In_246,In_394);
nand U1350 (N_1350,In_336,In_1249);
xnor U1351 (N_1351,In_1355,In_1922);
xor U1352 (N_1352,In_19,In_1519);
nor U1353 (N_1353,In_1024,In_249);
and U1354 (N_1354,In_162,In_806);
xor U1355 (N_1355,In_1779,In_1134);
xnor U1356 (N_1356,In_71,In_1386);
and U1357 (N_1357,In_1181,In_1728);
nor U1358 (N_1358,In_842,In_1691);
nor U1359 (N_1359,In_964,In_243);
and U1360 (N_1360,In_1111,In_1624);
nand U1361 (N_1361,In_662,In_908);
xnor U1362 (N_1362,In_1018,In_445);
or U1363 (N_1363,In_445,In_1548);
and U1364 (N_1364,In_860,In_1998);
nor U1365 (N_1365,In_538,In_772);
and U1366 (N_1366,In_1860,In_308);
nor U1367 (N_1367,In_416,In_653);
or U1368 (N_1368,In_1303,In_353);
nand U1369 (N_1369,In_1308,In_1472);
nand U1370 (N_1370,In_716,In_1257);
nor U1371 (N_1371,In_537,In_1456);
or U1372 (N_1372,In_277,In_1097);
or U1373 (N_1373,In_411,In_920);
nor U1374 (N_1374,In_612,In_599);
nand U1375 (N_1375,In_1198,In_1868);
and U1376 (N_1376,In_1306,In_1401);
and U1377 (N_1377,In_1873,In_494);
and U1378 (N_1378,In_697,In_1427);
xnor U1379 (N_1379,In_702,In_1825);
xnor U1380 (N_1380,In_1272,In_1816);
and U1381 (N_1381,In_1888,In_4);
and U1382 (N_1382,In_1490,In_1046);
nor U1383 (N_1383,In_792,In_1607);
nand U1384 (N_1384,In_1111,In_1844);
nor U1385 (N_1385,In_1490,In_951);
or U1386 (N_1386,In_1344,In_815);
and U1387 (N_1387,In_1690,In_853);
and U1388 (N_1388,In_706,In_632);
nor U1389 (N_1389,In_1125,In_1953);
and U1390 (N_1390,In_315,In_304);
nor U1391 (N_1391,In_1907,In_298);
xor U1392 (N_1392,In_1574,In_978);
nor U1393 (N_1393,In_620,In_1128);
xnor U1394 (N_1394,In_187,In_598);
nor U1395 (N_1395,In_68,In_1149);
nor U1396 (N_1396,In_1880,In_1374);
or U1397 (N_1397,In_1348,In_534);
nand U1398 (N_1398,In_1269,In_1742);
nand U1399 (N_1399,In_1935,In_1292);
or U1400 (N_1400,In_1640,In_1502);
and U1401 (N_1401,In_1714,In_12);
nand U1402 (N_1402,In_1102,In_534);
and U1403 (N_1403,In_408,In_278);
or U1404 (N_1404,In_362,In_862);
xnor U1405 (N_1405,In_1676,In_1748);
and U1406 (N_1406,In_1801,In_1536);
and U1407 (N_1407,In_744,In_481);
xor U1408 (N_1408,In_1371,In_493);
xnor U1409 (N_1409,In_1873,In_1152);
and U1410 (N_1410,In_808,In_14);
xor U1411 (N_1411,In_440,In_1747);
or U1412 (N_1412,In_1888,In_350);
nand U1413 (N_1413,In_444,In_563);
xnor U1414 (N_1414,In_1938,In_56);
or U1415 (N_1415,In_919,In_305);
nand U1416 (N_1416,In_1845,In_110);
and U1417 (N_1417,In_1527,In_1359);
or U1418 (N_1418,In_606,In_1163);
nor U1419 (N_1419,In_1005,In_120);
or U1420 (N_1420,In_1382,In_1730);
or U1421 (N_1421,In_1764,In_577);
nor U1422 (N_1422,In_249,In_140);
and U1423 (N_1423,In_529,In_28);
xnor U1424 (N_1424,In_1805,In_1777);
or U1425 (N_1425,In_1143,In_615);
xor U1426 (N_1426,In_860,In_1897);
nor U1427 (N_1427,In_1439,In_903);
or U1428 (N_1428,In_1588,In_1831);
and U1429 (N_1429,In_145,In_577);
or U1430 (N_1430,In_160,In_219);
or U1431 (N_1431,In_215,In_1499);
xor U1432 (N_1432,In_1275,In_1601);
nor U1433 (N_1433,In_1654,In_1648);
and U1434 (N_1434,In_1814,In_1519);
nand U1435 (N_1435,In_884,In_368);
and U1436 (N_1436,In_21,In_1298);
xor U1437 (N_1437,In_1028,In_1284);
nor U1438 (N_1438,In_1723,In_1671);
nor U1439 (N_1439,In_687,In_1296);
or U1440 (N_1440,In_1096,In_1130);
nor U1441 (N_1441,In_1036,In_374);
and U1442 (N_1442,In_1894,In_970);
or U1443 (N_1443,In_243,In_1590);
nand U1444 (N_1444,In_114,In_1286);
nand U1445 (N_1445,In_773,In_235);
and U1446 (N_1446,In_672,In_1284);
or U1447 (N_1447,In_1506,In_1838);
and U1448 (N_1448,In_1761,In_1610);
nor U1449 (N_1449,In_983,In_448);
xnor U1450 (N_1450,In_1782,In_1607);
nand U1451 (N_1451,In_858,In_689);
or U1452 (N_1452,In_233,In_770);
nand U1453 (N_1453,In_1561,In_1695);
or U1454 (N_1454,In_1928,In_628);
and U1455 (N_1455,In_1933,In_1897);
and U1456 (N_1456,In_461,In_1909);
or U1457 (N_1457,In_196,In_1165);
xor U1458 (N_1458,In_14,In_1583);
nand U1459 (N_1459,In_390,In_1942);
nand U1460 (N_1460,In_766,In_1547);
xnor U1461 (N_1461,In_546,In_1489);
nor U1462 (N_1462,In_1103,In_1001);
and U1463 (N_1463,In_70,In_1362);
and U1464 (N_1464,In_456,In_567);
nor U1465 (N_1465,In_1839,In_715);
or U1466 (N_1466,In_1861,In_627);
xnor U1467 (N_1467,In_419,In_124);
nand U1468 (N_1468,In_1245,In_313);
nor U1469 (N_1469,In_1758,In_1216);
nor U1470 (N_1470,In_1380,In_1553);
nand U1471 (N_1471,In_1653,In_454);
and U1472 (N_1472,In_1356,In_1703);
and U1473 (N_1473,In_1486,In_277);
nand U1474 (N_1474,In_1486,In_1796);
nand U1475 (N_1475,In_1340,In_1946);
and U1476 (N_1476,In_1179,In_637);
or U1477 (N_1477,In_192,In_1237);
xnor U1478 (N_1478,In_1942,In_808);
nand U1479 (N_1479,In_258,In_1213);
or U1480 (N_1480,In_943,In_423);
xnor U1481 (N_1481,In_933,In_1593);
nand U1482 (N_1482,In_1918,In_454);
xnor U1483 (N_1483,In_370,In_866);
or U1484 (N_1484,In_895,In_1191);
nor U1485 (N_1485,In_1468,In_1178);
nand U1486 (N_1486,In_507,In_1777);
or U1487 (N_1487,In_1635,In_1935);
xnor U1488 (N_1488,In_1750,In_294);
nor U1489 (N_1489,In_399,In_671);
nor U1490 (N_1490,In_206,In_1323);
or U1491 (N_1491,In_441,In_1304);
nand U1492 (N_1492,In_1761,In_692);
and U1493 (N_1493,In_636,In_1756);
nor U1494 (N_1494,In_1083,In_1230);
or U1495 (N_1495,In_1990,In_1000);
or U1496 (N_1496,In_1902,In_1090);
and U1497 (N_1497,In_1587,In_919);
nand U1498 (N_1498,In_1347,In_53);
nand U1499 (N_1499,In_1043,In_1075);
nand U1500 (N_1500,In_489,In_852);
xnor U1501 (N_1501,In_546,In_1015);
or U1502 (N_1502,In_1266,In_647);
or U1503 (N_1503,In_1637,In_1360);
nand U1504 (N_1504,In_134,In_1203);
xnor U1505 (N_1505,In_1388,In_1683);
nand U1506 (N_1506,In_1657,In_1406);
or U1507 (N_1507,In_68,In_1065);
nor U1508 (N_1508,In_653,In_1220);
and U1509 (N_1509,In_683,In_1358);
xnor U1510 (N_1510,In_614,In_270);
or U1511 (N_1511,In_1638,In_1787);
nor U1512 (N_1512,In_767,In_570);
xnor U1513 (N_1513,In_1778,In_355);
xnor U1514 (N_1514,In_97,In_1159);
nand U1515 (N_1515,In_622,In_205);
nor U1516 (N_1516,In_1332,In_349);
and U1517 (N_1517,In_1831,In_1301);
xor U1518 (N_1518,In_52,In_1699);
or U1519 (N_1519,In_542,In_1387);
and U1520 (N_1520,In_108,In_1016);
nor U1521 (N_1521,In_869,In_69);
or U1522 (N_1522,In_1625,In_26);
or U1523 (N_1523,In_1175,In_869);
and U1524 (N_1524,In_1242,In_1432);
xnor U1525 (N_1525,In_25,In_1421);
nand U1526 (N_1526,In_1008,In_777);
nand U1527 (N_1527,In_1246,In_259);
nor U1528 (N_1528,In_1666,In_1311);
and U1529 (N_1529,In_1669,In_460);
and U1530 (N_1530,In_1680,In_1461);
nand U1531 (N_1531,In_1237,In_788);
and U1532 (N_1532,In_365,In_1868);
nand U1533 (N_1533,In_1745,In_951);
and U1534 (N_1534,In_1439,In_991);
nor U1535 (N_1535,In_274,In_954);
or U1536 (N_1536,In_1334,In_1895);
nand U1537 (N_1537,In_826,In_775);
xnor U1538 (N_1538,In_814,In_1096);
and U1539 (N_1539,In_810,In_936);
xnor U1540 (N_1540,In_467,In_1159);
and U1541 (N_1541,In_913,In_1129);
nand U1542 (N_1542,In_594,In_55);
and U1543 (N_1543,In_723,In_982);
or U1544 (N_1544,In_620,In_121);
xor U1545 (N_1545,In_658,In_416);
and U1546 (N_1546,In_423,In_923);
nor U1547 (N_1547,In_1681,In_168);
and U1548 (N_1548,In_743,In_1009);
xnor U1549 (N_1549,In_1546,In_1008);
or U1550 (N_1550,In_1,In_1407);
nor U1551 (N_1551,In_115,In_586);
nor U1552 (N_1552,In_147,In_1101);
nand U1553 (N_1553,In_1643,In_1758);
nor U1554 (N_1554,In_808,In_1020);
or U1555 (N_1555,In_804,In_1407);
xnor U1556 (N_1556,In_1563,In_1966);
nand U1557 (N_1557,In_1939,In_1573);
or U1558 (N_1558,In_596,In_1118);
nand U1559 (N_1559,In_1901,In_689);
or U1560 (N_1560,In_1599,In_1368);
and U1561 (N_1561,In_506,In_913);
xor U1562 (N_1562,In_1155,In_1784);
xnor U1563 (N_1563,In_18,In_780);
nor U1564 (N_1564,In_1747,In_1924);
nand U1565 (N_1565,In_992,In_1009);
and U1566 (N_1566,In_1253,In_1338);
xor U1567 (N_1567,In_439,In_113);
or U1568 (N_1568,In_213,In_1349);
and U1569 (N_1569,In_1429,In_52);
and U1570 (N_1570,In_757,In_471);
xnor U1571 (N_1571,In_1566,In_956);
or U1572 (N_1572,In_286,In_1370);
and U1573 (N_1573,In_1515,In_232);
or U1574 (N_1574,In_1313,In_51);
nor U1575 (N_1575,In_308,In_1899);
or U1576 (N_1576,In_419,In_114);
nor U1577 (N_1577,In_108,In_1668);
xor U1578 (N_1578,In_1830,In_557);
and U1579 (N_1579,In_1697,In_1995);
nor U1580 (N_1580,In_371,In_1470);
nand U1581 (N_1581,In_101,In_1714);
and U1582 (N_1582,In_1429,In_1753);
or U1583 (N_1583,In_1425,In_867);
and U1584 (N_1584,In_303,In_1797);
and U1585 (N_1585,In_414,In_589);
nor U1586 (N_1586,In_1222,In_1063);
xor U1587 (N_1587,In_1685,In_1213);
nor U1588 (N_1588,In_1277,In_1092);
nand U1589 (N_1589,In_434,In_543);
nor U1590 (N_1590,In_1951,In_747);
or U1591 (N_1591,In_137,In_1644);
and U1592 (N_1592,In_124,In_120);
nand U1593 (N_1593,In_1459,In_1529);
and U1594 (N_1594,In_1855,In_100);
xor U1595 (N_1595,In_538,In_1233);
nor U1596 (N_1596,In_1518,In_1300);
and U1597 (N_1597,In_1856,In_864);
xnor U1598 (N_1598,In_1248,In_607);
and U1599 (N_1599,In_1244,In_1438);
nand U1600 (N_1600,In_813,In_888);
or U1601 (N_1601,In_1792,In_576);
and U1602 (N_1602,In_1634,In_1745);
nor U1603 (N_1603,In_1401,In_77);
nor U1604 (N_1604,In_1587,In_300);
xnor U1605 (N_1605,In_1487,In_146);
nand U1606 (N_1606,In_913,In_1836);
nor U1607 (N_1607,In_716,In_1180);
and U1608 (N_1608,In_116,In_288);
and U1609 (N_1609,In_1807,In_923);
xor U1610 (N_1610,In_1117,In_1179);
nand U1611 (N_1611,In_1522,In_489);
nor U1612 (N_1612,In_1685,In_1144);
nand U1613 (N_1613,In_1989,In_1801);
xor U1614 (N_1614,In_347,In_1589);
xnor U1615 (N_1615,In_1709,In_181);
and U1616 (N_1616,In_590,In_356);
nand U1617 (N_1617,In_1802,In_201);
or U1618 (N_1618,In_1106,In_1328);
and U1619 (N_1619,In_1590,In_693);
xor U1620 (N_1620,In_1479,In_681);
xnor U1621 (N_1621,In_1308,In_1073);
nand U1622 (N_1622,In_654,In_638);
or U1623 (N_1623,In_1100,In_141);
or U1624 (N_1624,In_1943,In_1203);
and U1625 (N_1625,In_350,In_1015);
or U1626 (N_1626,In_893,In_924);
or U1627 (N_1627,In_1850,In_262);
nand U1628 (N_1628,In_140,In_1985);
nor U1629 (N_1629,In_1474,In_1130);
and U1630 (N_1630,In_955,In_679);
or U1631 (N_1631,In_757,In_539);
xor U1632 (N_1632,In_1825,In_1099);
nand U1633 (N_1633,In_426,In_1088);
xor U1634 (N_1634,In_710,In_781);
and U1635 (N_1635,In_658,In_697);
and U1636 (N_1636,In_31,In_813);
or U1637 (N_1637,In_342,In_626);
or U1638 (N_1638,In_1668,In_304);
and U1639 (N_1639,In_1899,In_350);
nor U1640 (N_1640,In_1223,In_159);
nand U1641 (N_1641,In_1292,In_493);
nand U1642 (N_1642,In_1680,In_311);
nand U1643 (N_1643,In_814,In_1957);
xnor U1644 (N_1644,In_1851,In_444);
nand U1645 (N_1645,In_1446,In_132);
nor U1646 (N_1646,In_1072,In_757);
nor U1647 (N_1647,In_321,In_1276);
or U1648 (N_1648,In_1100,In_1720);
or U1649 (N_1649,In_197,In_1931);
xnor U1650 (N_1650,In_542,In_1090);
xor U1651 (N_1651,In_1537,In_1270);
and U1652 (N_1652,In_1776,In_944);
and U1653 (N_1653,In_877,In_741);
nand U1654 (N_1654,In_1269,In_249);
and U1655 (N_1655,In_305,In_1987);
xor U1656 (N_1656,In_550,In_57);
nand U1657 (N_1657,In_895,In_960);
nor U1658 (N_1658,In_913,In_269);
or U1659 (N_1659,In_1801,In_1390);
nor U1660 (N_1660,In_1465,In_361);
nor U1661 (N_1661,In_1368,In_1247);
and U1662 (N_1662,In_960,In_984);
and U1663 (N_1663,In_1536,In_1973);
nor U1664 (N_1664,In_1990,In_1192);
or U1665 (N_1665,In_1010,In_1362);
and U1666 (N_1666,In_467,In_1118);
nor U1667 (N_1667,In_306,In_1065);
xor U1668 (N_1668,In_1167,In_61);
nand U1669 (N_1669,In_1919,In_1115);
nand U1670 (N_1670,In_1122,In_915);
nor U1671 (N_1671,In_527,In_885);
or U1672 (N_1672,In_685,In_1670);
xnor U1673 (N_1673,In_27,In_232);
and U1674 (N_1674,In_1767,In_551);
or U1675 (N_1675,In_859,In_1565);
xnor U1676 (N_1676,In_167,In_1994);
and U1677 (N_1677,In_55,In_554);
or U1678 (N_1678,In_878,In_1400);
or U1679 (N_1679,In_1963,In_972);
nand U1680 (N_1680,In_361,In_879);
and U1681 (N_1681,In_983,In_1318);
xnor U1682 (N_1682,In_1117,In_1636);
nor U1683 (N_1683,In_40,In_1465);
and U1684 (N_1684,In_934,In_1);
and U1685 (N_1685,In_876,In_1487);
nor U1686 (N_1686,In_1326,In_243);
xnor U1687 (N_1687,In_265,In_574);
or U1688 (N_1688,In_1216,In_1723);
xor U1689 (N_1689,In_1351,In_1595);
xor U1690 (N_1690,In_217,In_1943);
nand U1691 (N_1691,In_1005,In_1098);
nor U1692 (N_1692,In_204,In_544);
or U1693 (N_1693,In_1826,In_1951);
nor U1694 (N_1694,In_873,In_1914);
xor U1695 (N_1695,In_878,In_894);
or U1696 (N_1696,In_489,In_1817);
nand U1697 (N_1697,In_1408,In_1070);
nand U1698 (N_1698,In_555,In_552);
and U1699 (N_1699,In_626,In_1388);
xnor U1700 (N_1700,In_1106,In_418);
nand U1701 (N_1701,In_979,In_1117);
and U1702 (N_1702,In_1220,In_1920);
nand U1703 (N_1703,In_1856,In_1086);
or U1704 (N_1704,In_1457,In_290);
xor U1705 (N_1705,In_1179,In_1530);
and U1706 (N_1706,In_133,In_1782);
nand U1707 (N_1707,In_1004,In_864);
xnor U1708 (N_1708,In_618,In_887);
nor U1709 (N_1709,In_409,In_629);
xor U1710 (N_1710,In_117,In_1202);
nor U1711 (N_1711,In_1432,In_1206);
nor U1712 (N_1712,In_1112,In_1224);
nor U1713 (N_1713,In_837,In_1259);
nand U1714 (N_1714,In_1375,In_407);
xor U1715 (N_1715,In_1374,In_1354);
and U1716 (N_1716,In_354,In_635);
xor U1717 (N_1717,In_851,In_1850);
nor U1718 (N_1718,In_739,In_1517);
nor U1719 (N_1719,In_482,In_1747);
or U1720 (N_1720,In_708,In_747);
or U1721 (N_1721,In_1910,In_267);
nand U1722 (N_1722,In_1557,In_1411);
xor U1723 (N_1723,In_1473,In_967);
nor U1724 (N_1724,In_1030,In_1782);
and U1725 (N_1725,In_1654,In_1479);
nand U1726 (N_1726,In_1706,In_47);
or U1727 (N_1727,In_1691,In_854);
nand U1728 (N_1728,In_1460,In_1971);
xnor U1729 (N_1729,In_823,In_324);
nor U1730 (N_1730,In_1078,In_1529);
xnor U1731 (N_1731,In_27,In_20);
nor U1732 (N_1732,In_1944,In_272);
xor U1733 (N_1733,In_1944,In_1479);
nor U1734 (N_1734,In_924,In_791);
nor U1735 (N_1735,In_865,In_844);
xnor U1736 (N_1736,In_1460,In_157);
or U1737 (N_1737,In_1834,In_205);
xnor U1738 (N_1738,In_355,In_1840);
and U1739 (N_1739,In_535,In_362);
or U1740 (N_1740,In_45,In_1746);
and U1741 (N_1741,In_1337,In_866);
nand U1742 (N_1742,In_536,In_1867);
and U1743 (N_1743,In_340,In_1922);
nor U1744 (N_1744,In_1739,In_427);
xor U1745 (N_1745,In_320,In_403);
and U1746 (N_1746,In_1752,In_380);
xor U1747 (N_1747,In_1178,In_1563);
nor U1748 (N_1748,In_665,In_1063);
and U1749 (N_1749,In_1268,In_965);
and U1750 (N_1750,In_1259,In_1791);
or U1751 (N_1751,In_947,In_1257);
xor U1752 (N_1752,In_1825,In_1236);
nand U1753 (N_1753,In_1350,In_1760);
nor U1754 (N_1754,In_1079,In_996);
nor U1755 (N_1755,In_96,In_851);
and U1756 (N_1756,In_732,In_32);
or U1757 (N_1757,In_80,In_789);
xor U1758 (N_1758,In_1714,In_1220);
xor U1759 (N_1759,In_400,In_1977);
or U1760 (N_1760,In_1782,In_1970);
and U1761 (N_1761,In_1125,In_1511);
or U1762 (N_1762,In_1036,In_1782);
nand U1763 (N_1763,In_1676,In_646);
xnor U1764 (N_1764,In_1712,In_247);
or U1765 (N_1765,In_689,In_1857);
nand U1766 (N_1766,In_1083,In_13);
or U1767 (N_1767,In_1954,In_665);
nand U1768 (N_1768,In_1260,In_1279);
nor U1769 (N_1769,In_596,In_1097);
and U1770 (N_1770,In_1388,In_1833);
nor U1771 (N_1771,In_434,In_1919);
nand U1772 (N_1772,In_1442,In_1379);
nor U1773 (N_1773,In_1093,In_1866);
xnor U1774 (N_1774,In_297,In_1155);
xor U1775 (N_1775,In_628,In_1671);
nand U1776 (N_1776,In_1645,In_1648);
and U1777 (N_1777,In_1430,In_1264);
or U1778 (N_1778,In_920,In_1880);
or U1779 (N_1779,In_1492,In_244);
xnor U1780 (N_1780,In_1660,In_1722);
nor U1781 (N_1781,In_494,In_1132);
xor U1782 (N_1782,In_1424,In_830);
nor U1783 (N_1783,In_1238,In_444);
nand U1784 (N_1784,In_226,In_1436);
nand U1785 (N_1785,In_99,In_661);
nand U1786 (N_1786,In_104,In_1973);
xnor U1787 (N_1787,In_1329,In_1331);
nand U1788 (N_1788,In_1265,In_751);
nor U1789 (N_1789,In_1554,In_1598);
and U1790 (N_1790,In_1817,In_26);
xor U1791 (N_1791,In_130,In_1274);
nand U1792 (N_1792,In_637,In_467);
and U1793 (N_1793,In_1422,In_294);
nand U1794 (N_1794,In_1016,In_1406);
nand U1795 (N_1795,In_4,In_1756);
and U1796 (N_1796,In_389,In_87);
or U1797 (N_1797,In_919,In_1286);
nand U1798 (N_1798,In_1800,In_1378);
nand U1799 (N_1799,In_153,In_466);
nor U1800 (N_1800,In_70,In_117);
nand U1801 (N_1801,In_291,In_1356);
or U1802 (N_1802,In_1112,In_581);
xnor U1803 (N_1803,In_1515,In_1941);
nand U1804 (N_1804,In_613,In_1810);
or U1805 (N_1805,In_1384,In_284);
or U1806 (N_1806,In_1323,In_628);
xor U1807 (N_1807,In_1436,In_491);
and U1808 (N_1808,In_1970,In_637);
nand U1809 (N_1809,In_1428,In_1650);
or U1810 (N_1810,In_1082,In_11);
nand U1811 (N_1811,In_272,In_928);
and U1812 (N_1812,In_696,In_1586);
xnor U1813 (N_1813,In_634,In_1694);
or U1814 (N_1814,In_1297,In_1383);
nor U1815 (N_1815,In_1838,In_1597);
nor U1816 (N_1816,In_594,In_1943);
or U1817 (N_1817,In_1600,In_243);
and U1818 (N_1818,In_389,In_1400);
and U1819 (N_1819,In_1666,In_711);
or U1820 (N_1820,In_320,In_615);
nand U1821 (N_1821,In_1754,In_754);
xor U1822 (N_1822,In_1521,In_1015);
and U1823 (N_1823,In_324,In_58);
and U1824 (N_1824,In_443,In_739);
or U1825 (N_1825,In_56,In_105);
and U1826 (N_1826,In_1495,In_1222);
nand U1827 (N_1827,In_937,In_1732);
xnor U1828 (N_1828,In_408,In_349);
xor U1829 (N_1829,In_835,In_458);
or U1830 (N_1830,In_796,In_74);
or U1831 (N_1831,In_637,In_1153);
xor U1832 (N_1832,In_807,In_1696);
nand U1833 (N_1833,In_132,In_549);
nor U1834 (N_1834,In_1066,In_1300);
nand U1835 (N_1835,In_1928,In_1301);
nor U1836 (N_1836,In_1658,In_593);
xor U1837 (N_1837,In_1099,In_581);
nand U1838 (N_1838,In_831,In_1645);
nor U1839 (N_1839,In_1917,In_1115);
nor U1840 (N_1840,In_204,In_725);
nor U1841 (N_1841,In_925,In_1504);
or U1842 (N_1842,In_1042,In_1957);
or U1843 (N_1843,In_93,In_237);
xor U1844 (N_1844,In_1837,In_776);
or U1845 (N_1845,In_1619,In_446);
or U1846 (N_1846,In_1332,In_1814);
nand U1847 (N_1847,In_1092,In_701);
and U1848 (N_1848,In_1493,In_935);
xnor U1849 (N_1849,In_478,In_1857);
nor U1850 (N_1850,In_669,In_176);
nor U1851 (N_1851,In_771,In_841);
xor U1852 (N_1852,In_957,In_857);
or U1853 (N_1853,In_1987,In_162);
nand U1854 (N_1854,In_270,In_869);
nand U1855 (N_1855,In_653,In_859);
and U1856 (N_1856,In_1966,In_927);
or U1857 (N_1857,In_258,In_264);
or U1858 (N_1858,In_1904,In_1477);
nand U1859 (N_1859,In_402,In_1234);
nand U1860 (N_1860,In_1916,In_595);
xnor U1861 (N_1861,In_12,In_86);
nand U1862 (N_1862,In_881,In_420);
nor U1863 (N_1863,In_1569,In_1215);
xor U1864 (N_1864,In_282,In_1262);
and U1865 (N_1865,In_1511,In_19);
nand U1866 (N_1866,In_1696,In_487);
xor U1867 (N_1867,In_1429,In_1356);
or U1868 (N_1868,In_1186,In_1741);
nor U1869 (N_1869,In_398,In_1102);
and U1870 (N_1870,In_725,In_367);
and U1871 (N_1871,In_1759,In_483);
nor U1872 (N_1872,In_1921,In_1654);
xnor U1873 (N_1873,In_10,In_1144);
and U1874 (N_1874,In_236,In_1023);
and U1875 (N_1875,In_1199,In_1962);
nor U1876 (N_1876,In_679,In_526);
nor U1877 (N_1877,In_1107,In_1290);
nand U1878 (N_1878,In_1237,In_162);
nand U1879 (N_1879,In_110,In_364);
or U1880 (N_1880,In_576,In_1587);
nand U1881 (N_1881,In_73,In_836);
nand U1882 (N_1882,In_1248,In_597);
nand U1883 (N_1883,In_623,In_995);
nor U1884 (N_1884,In_178,In_1742);
and U1885 (N_1885,In_437,In_1248);
nand U1886 (N_1886,In_603,In_1170);
xnor U1887 (N_1887,In_1559,In_458);
nand U1888 (N_1888,In_890,In_462);
and U1889 (N_1889,In_745,In_1000);
nand U1890 (N_1890,In_1080,In_1447);
xnor U1891 (N_1891,In_700,In_1671);
xor U1892 (N_1892,In_185,In_1821);
and U1893 (N_1893,In_1249,In_1632);
and U1894 (N_1894,In_674,In_1323);
or U1895 (N_1895,In_849,In_124);
or U1896 (N_1896,In_1315,In_1259);
or U1897 (N_1897,In_1009,In_1296);
and U1898 (N_1898,In_1215,In_604);
and U1899 (N_1899,In_1345,In_274);
xor U1900 (N_1900,In_1589,In_1333);
or U1901 (N_1901,In_520,In_1643);
and U1902 (N_1902,In_1254,In_621);
and U1903 (N_1903,In_1239,In_397);
xnor U1904 (N_1904,In_1301,In_359);
nor U1905 (N_1905,In_356,In_1111);
nor U1906 (N_1906,In_1070,In_1321);
or U1907 (N_1907,In_807,In_1679);
nor U1908 (N_1908,In_1094,In_1680);
nor U1909 (N_1909,In_1015,In_1148);
nand U1910 (N_1910,In_962,In_663);
xnor U1911 (N_1911,In_1523,In_341);
nand U1912 (N_1912,In_347,In_90);
and U1913 (N_1913,In_288,In_1009);
or U1914 (N_1914,In_1052,In_358);
and U1915 (N_1915,In_95,In_231);
xnor U1916 (N_1916,In_1599,In_460);
xor U1917 (N_1917,In_1641,In_1726);
and U1918 (N_1918,In_692,In_1043);
xor U1919 (N_1919,In_476,In_1760);
nor U1920 (N_1920,In_1526,In_1901);
xor U1921 (N_1921,In_442,In_1454);
nand U1922 (N_1922,In_1060,In_540);
or U1923 (N_1923,In_228,In_569);
or U1924 (N_1924,In_1301,In_1946);
or U1925 (N_1925,In_558,In_646);
xnor U1926 (N_1926,In_408,In_1612);
xnor U1927 (N_1927,In_109,In_412);
and U1928 (N_1928,In_630,In_1262);
or U1929 (N_1929,In_262,In_1353);
xnor U1930 (N_1930,In_643,In_996);
nor U1931 (N_1931,In_776,In_853);
xnor U1932 (N_1932,In_303,In_1331);
xor U1933 (N_1933,In_153,In_142);
and U1934 (N_1934,In_1498,In_578);
or U1935 (N_1935,In_133,In_327);
nand U1936 (N_1936,In_1928,In_1354);
nand U1937 (N_1937,In_308,In_1475);
xor U1938 (N_1938,In_1770,In_1672);
nand U1939 (N_1939,In_753,In_707);
xnor U1940 (N_1940,In_1594,In_126);
nand U1941 (N_1941,In_664,In_1850);
nand U1942 (N_1942,In_520,In_338);
or U1943 (N_1943,In_1146,In_630);
nor U1944 (N_1944,In_705,In_45);
xor U1945 (N_1945,In_1342,In_24);
nor U1946 (N_1946,In_958,In_988);
nand U1947 (N_1947,In_1212,In_464);
or U1948 (N_1948,In_1943,In_427);
nand U1949 (N_1949,In_1160,In_1756);
xor U1950 (N_1950,In_326,In_1953);
xnor U1951 (N_1951,In_1279,In_758);
xor U1952 (N_1952,In_1305,In_1306);
nor U1953 (N_1953,In_1324,In_1891);
nor U1954 (N_1954,In_887,In_1083);
nand U1955 (N_1955,In_1087,In_1485);
nand U1956 (N_1956,In_767,In_1050);
and U1957 (N_1957,In_27,In_513);
and U1958 (N_1958,In_292,In_1241);
and U1959 (N_1959,In_1778,In_1203);
nor U1960 (N_1960,In_1109,In_1634);
xnor U1961 (N_1961,In_991,In_1280);
nor U1962 (N_1962,In_210,In_346);
nor U1963 (N_1963,In_283,In_245);
and U1964 (N_1964,In_1585,In_1355);
and U1965 (N_1965,In_86,In_755);
and U1966 (N_1966,In_1633,In_1103);
or U1967 (N_1967,In_540,In_349);
nand U1968 (N_1968,In_139,In_205);
nand U1969 (N_1969,In_1152,In_365);
nor U1970 (N_1970,In_67,In_188);
nor U1971 (N_1971,In_1476,In_1339);
nand U1972 (N_1972,In_1623,In_1408);
xor U1973 (N_1973,In_1225,In_891);
and U1974 (N_1974,In_156,In_836);
nand U1975 (N_1975,In_1575,In_556);
and U1976 (N_1976,In_69,In_927);
and U1977 (N_1977,In_1989,In_1685);
or U1978 (N_1978,In_1914,In_241);
nor U1979 (N_1979,In_182,In_368);
nand U1980 (N_1980,In_1510,In_1292);
xnor U1981 (N_1981,In_183,In_52);
or U1982 (N_1982,In_269,In_705);
nor U1983 (N_1983,In_1878,In_1912);
nand U1984 (N_1984,In_1043,In_1346);
and U1985 (N_1985,In_221,In_1879);
xnor U1986 (N_1986,In_472,In_1164);
xor U1987 (N_1987,In_377,In_1868);
and U1988 (N_1988,In_1135,In_1992);
and U1989 (N_1989,In_1763,In_873);
or U1990 (N_1990,In_399,In_1248);
or U1991 (N_1991,In_1536,In_884);
or U1992 (N_1992,In_1065,In_1447);
xor U1993 (N_1993,In_1824,In_341);
xor U1994 (N_1994,In_1427,In_1211);
or U1995 (N_1995,In_789,In_706);
nor U1996 (N_1996,In_412,In_1560);
nor U1997 (N_1997,In_1403,In_464);
and U1998 (N_1998,In_1706,In_211);
and U1999 (N_1999,In_1158,In_609);
xor U2000 (N_2000,In_441,In_803);
nor U2001 (N_2001,In_548,In_324);
xor U2002 (N_2002,In_1911,In_1307);
xor U2003 (N_2003,In_1503,In_1480);
and U2004 (N_2004,In_433,In_95);
and U2005 (N_2005,In_669,In_1964);
nor U2006 (N_2006,In_717,In_685);
nand U2007 (N_2007,In_392,In_1092);
nor U2008 (N_2008,In_1287,In_1563);
xor U2009 (N_2009,In_1935,In_1308);
or U2010 (N_2010,In_295,In_1924);
nor U2011 (N_2011,In_94,In_1275);
nand U2012 (N_2012,In_940,In_1545);
and U2013 (N_2013,In_1178,In_255);
or U2014 (N_2014,In_1968,In_498);
xor U2015 (N_2015,In_1099,In_649);
xor U2016 (N_2016,In_384,In_1817);
nand U2017 (N_2017,In_153,In_146);
xnor U2018 (N_2018,In_436,In_11);
nand U2019 (N_2019,In_69,In_21);
nand U2020 (N_2020,In_815,In_1846);
xor U2021 (N_2021,In_1734,In_1152);
xor U2022 (N_2022,In_168,In_276);
nand U2023 (N_2023,In_415,In_1242);
or U2024 (N_2024,In_1220,In_1869);
or U2025 (N_2025,In_1725,In_646);
nor U2026 (N_2026,In_589,In_966);
nand U2027 (N_2027,In_138,In_1834);
nand U2028 (N_2028,In_1950,In_109);
nand U2029 (N_2029,In_1785,In_1801);
xnor U2030 (N_2030,In_1393,In_302);
nand U2031 (N_2031,In_1230,In_1345);
xnor U2032 (N_2032,In_1873,In_440);
xnor U2033 (N_2033,In_1428,In_1655);
or U2034 (N_2034,In_327,In_519);
nand U2035 (N_2035,In_234,In_1124);
or U2036 (N_2036,In_1080,In_673);
or U2037 (N_2037,In_385,In_1572);
nor U2038 (N_2038,In_983,In_1027);
nor U2039 (N_2039,In_467,In_1274);
or U2040 (N_2040,In_1475,In_615);
nor U2041 (N_2041,In_750,In_562);
nor U2042 (N_2042,In_1468,In_1386);
nor U2043 (N_2043,In_1438,In_585);
or U2044 (N_2044,In_122,In_1801);
xor U2045 (N_2045,In_64,In_1050);
nor U2046 (N_2046,In_1087,In_1608);
xnor U2047 (N_2047,In_1408,In_1677);
nand U2048 (N_2048,In_1726,In_784);
and U2049 (N_2049,In_1168,In_315);
nand U2050 (N_2050,In_656,In_1795);
xor U2051 (N_2051,In_1460,In_791);
xor U2052 (N_2052,In_195,In_1616);
nand U2053 (N_2053,In_1934,In_1047);
or U2054 (N_2054,In_1610,In_1443);
nand U2055 (N_2055,In_733,In_134);
xor U2056 (N_2056,In_404,In_1364);
nor U2057 (N_2057,In_1209,In_1652);
or U2058 (N_2058,In_1667,In_1112);
and U2059 (N_2059,In_1034,In_1406);
nor U2060 (N_2060,In_1480,In_893);
nor U2061 (N_2061,In_87,In_1120);
xnor U2062 (N_2062,In_399,In_1938);
and U2063 (N_2063,In_1146,In_1189);
xnor U2064 (N_2064,In_1144,In_1305);
nor U2065 (N_2065,In_806,In_43);
nor U2066 (N_2066,In_5,In_583);
nor U2067 (N_2067,In_1014,In_455);
or U2068 (N_2068,In_627,In_1900);
xor U2069 (N_2069,In_1580,In_890);
or U2070 (N_2070,In_31,In_1229);
xnor U2071 (N_2071,In_458,In_113);
and U2072 (N_2072,In_872,In_1324);
and U2073 (N_2073,In_193,In_546);
nand U2074 (N_2074,In_1932,In_459);
xor U2075 (N_2075,In_1666,In_1576);
and U2076 (N_2076,In_1135,In_849);
nand U2077 (N_2077,In_373,In_694);
and U2078 (N_2078,In_926,In_842);
nand U2079 (N_2079,In_225,In_1821);
and U2080 (N_2080,In_1631,In_395);
nor U2081 (N_2081,In_32,In_1036);
nor U2082 (N_2082,In_464,In_993);
and U2083 (N_2083,In_950,In_848);
nand U2084 (N_2084,In_178,In_1658);
nor U2085 (N_2085,In_51,In_817);
or U2086 (N_2086,In_1540,In_815);
or U2087 (N_2087,In_1781,In_1507);
and U2088 (N_2088,In_336,In_1409);
nor U2089 (N_2089,In_819,In_556);
xor U2090 (N_2090,In_1297,In_1417);
and U2091 (N_2091,In_188,In_1119);
nor U2092 (N_2092,In_210,In_1192);
or U2093 (N_2093,In_1884,In_1853);
nor U2094 (N_2094,In_1825,In_1427);
nor U2095 (N_2095,In_153,In_493);
or U2096 (N_2096,In_1883,In_67);
nor U2097 (N_2097,In_467,In_1270);
and U2098 (N_2098,In_1023,In_1954);
or U2099 (N_2099,In_916,In_1268);
nor U2100 (N_2100,In_543,In_817);
nand U2101 (N_2101,In_739,In_273);
nor U2102 (N_2102,In_277,In_389);
nor U2103 (N_2103,In_1108,In_1465);
and U2104 (N_2104,In_417,In_1820);
nor U2105 (N_2105,In_257,In_1970);
or U2106 (N_2106,In_2,In_1056);
nand U2107 (N_2107,In_1435,In_1502);
and U2108 (N_2108,In_611,In_1460);
xor U2109 (N_2109,In_402,In_1138);
and U2110 (N_2110,In_1674,In_943);
xor U2111 (N_2111,In_1819,In_470);
nand U2112 (N_2112,In_897,In_22);
nor U2113 (N_2113,In_94,In_1635);
xor U2114 (N_2114,In_650,In_1636);
xor U2115 (N_2115,In_352,In_562);
nand U2116 (N_2116,In_280,In_1723);
and U2117 (N_2117,In_1240,In_1660);
nor U2118 (N_2118,In_399,In_569);
and U2119 (N_2119,In_831,In_1095);
or U2120 (N_2120,In_1646,In_1424);
xor U2121 (N_2121,In_1312,In_167);
xnor U2122 (N_2122,In_786,In_310);
and U2123 (N_2123,In_1058,In_1828);
xnor U2124 (N_2124,In_347,In_1762);
nor U2125 (N_2125,In_547,In_773);
and U2126 (N_2126,In_1936,In_1780);
and U2127 (N_2127,In_1357,In_679);
and U2128 (N_2128,In_1624,In_1066);
xnor U2129 (N_2129,In_625,In_1369);
nor U2130 (N_2130,In_973,In_1905);
and U2131 (N_2131,In_19,In_736);
nor U2132 (N_2132,In_259,In_1597);
nand U2133 (N_2133,In_1959,In_398);
and U2134 (N_2134,In_693,In_1471);
nor U2135 (N_2135,In_27,In_1273);
or U2136 (N_2136,In_84,In_1334);
nand U2137 (N_2137,In_1297,In_1752);
xor U2138 (N_2138,In_336,In_1898);
nor U2139 (N_2139,In_1687,In_1220);
nand U2140 (N_2140,In_253,In_1339);
nand U2141 (N_2141,In_340,In_613);
nor U2142 (N_2142,In_986,In_266);
nor U2143 (N_2143,In_673,In_1786);
xor U2144 (N_2144,In_137,In_856);
or U2145 (N_2145,In_1432,In_334);
nor U2146 (N_2146,In_1760,In_1965);
or U2147 (N_2147,In_957,In_1759);
nand U2148 (N_2148,In_1846,In_3);
and U2149 (N_2149,In_1216,In_1959);
nand U2150 (N_2150,In_1062,In_546);
or U2151 (N_2151,In_1770,In_1464);
or U2152 (N_2152,In_1263,In_1748);
and U2153 (N_2153,In_270,In_842);
xnor U2154 (N_2154,In_933,In_1029);
xnor U2155 (N_2155,In_583,In_1451);
nand U2156 (N_2156,In_1178,In_1052);
or U2157 (N_2157,In_519,In_1107);
nor U2158 (N_2158,In_429,In_343);
and U2159 (N_2159,In_1379,In_20);
nand U2160 (N_2160,In_1140,In_252);
nand U2161 (N_2161,In_1,In_290);
nor U2162 (N_2162,In_1066,In_164);
and U2163 (N_2163,In_1961,In_1420);
nand U2164 (N_2164,In_1168,In_1216);
nand U2165 (N_2165,In_743,In_961);
nand U2166 (N_2166,In_1955,In_924);
and U2167 (N_2167,In_911,In_794);
nor U2168 (N_2168,In_1608,In_1368);
xor U2169 (N_2169,In_1909,In_198);
or U2170 (N_2170,In_662,In_1196);
xnor U2171 (N_2171,In_1504,In_35);
nand U2172 (N_2172,In_578,In_48);
and U2173 (N_2173,In_1073,In_522);
and U2174 (N_2174,In_205,In_1433);
nand U2175 (N_2175,In_1330,In_246);
nor U2176 (N_2176,In_1909,In_869);
and U2177 (N_2177,In_112,In_444);
or U2178 (N_2178,In_379,In_812);
or U2179 (N_2179,In_1167,In_720);
or U2180 (N_2180,In_1917,In_715);
nor U2181 (N_2181,In_693,In_352);
nor U2182 (N_2182,In_445,In_1371);
and U2183 (N_2183,In_129,In_83);
and U2184 (N_2184,In_326,In_1780);
nand U2185 (N_2185,In_1778,In_1828);
and U2186 (N_2186,In_1257,In_793);
or U2187 (N_2187,In_627,In_1096);
nand U2188 (N_2188,In_803,In_1611);
nor U2189 (N_2189,In_1863,In_1203);
and U2190 (N_2190,In_1443,In_55);
or U2191 (N_2191,In_493,In_319);
nand U2192 (N_2192,In_1490,In_876);
nand U2193 (N_2193,In_652,In_751);
xnor U2194 (N_2194,In_1451,In_29);
nand U2195 (N_2195,In_1365,In_626);
nand U2196 (N_2196,In_492,In_672);
and U2197 (N_2197,In_1112,In_915);
nor U2198 (N_2198,In_881,In_1109);
and U2199 (N_2199,In_1730,In_635);
or U2200 (N_2200,In_760,In_1746);
nand U2201 (N_2201,In_1210,In_468);
xor U2202 (N_2202,In_1797,In_1825);
nand U2203 (N_2203,In_1412,In_677);
or U2204 (N_2204,In_343,In_266);
nor U2205 (N_2205,In_105,In_923);
or U2206 (N_2206,In_1601,In_421);
xnor U2207 (N_2207,In_257,In_697);
nand U2208 (N_2208,In_871,In_281);
and U2209 (N_2209,In_1982,In_886);
or U2210 (N_2210,In_1658,In_1236);
nor U2211 (N_2211,In_1533,In_1581);
nand U2212 (N_2212,In_1034,In_1366);
nor U2213 (N_2213,In_103,In_669);
nand U2214 (N_2214,In_593,In_1773);
xor U2215 (N_2215,In_139,In_1660);
nand U2216 (N_2216,In_1355,In_139);
and U2217 (N_2217,In_1951,In_1390);
and U2218 (N_2218,In_187,In_991);
or U2219 (N_2219,In_1389,In_1146);
xnor U2220 (N_2220,In_118,In_1701);
and U2221 (N_2221,In_585,In_1671);
xnor U2222 (N_2222,In_19,In_668);
or U2223 (N_2223,In_960,In_1879);
xor U2224 (N_2224,In_772,In_1091);
or U2225 (N_2225,In_1181,In_537);
or U2226 (N_2226,In_948,In_1544);
xor U2227 (N_2227,In_394,In_1660);
and U2228 (N_2228,In_1895,In_865);
or U2229 (N_2229,In_89,In_1298);
nor U2230 (N_2230,In_483,In_613);
xor U2231 (N_2231,In_1560,In_1485);
xor U2232 (N_2232,In_1290,In_1257);
xor U2233 (N_2233,In_153,In_221);
nor U2234 (N_2234,In_245,In_509);
nor U2235 (N_2235,In_56,In_637);
or U2236 (N_2236,In_615,In_1720);
and U2237 (N_2237,In_1753,In_302);
nor U2238 (N_2238,In_866,In_1915);
or U2239 (N_2239,In_852,In_788);
or U2240 (N_2240,In_1376,In_1811);
nand U2241 (N_2241,In_34,In_1474);
and U2242 (N_2242,In_142,In_568);
xnor U2243 (N_2243,In_1121,In_102);
or U2244 (N_2244,In_938,In_175);
and U2245 (N_2245,In_138,In_657);
and U2246 (N_2246,In_1290,In_942);
xnor U2247 (N_2247,In_301,In_1761);
xor U2248 (N_2248,In_1891,In_175);
or U2249 (N_2249,In_1922,In_1858);
xnor U2250 (N_2250,In_1929,In_301);
or U2251 (N_2251,In_1448,In_1085);
and U2252 (N_2252,In_1271,In_1848);
nor U2253 (N_2253,In_811,In_1598);
or U2254 (N_2254,In_408,In_18);
nand U2255 (N_2255,In_257,In_1290);
xnor U2256 (N_2256,In_1186,In_138);
and U2257 (N_2257,In_700,In_1793);
xnor U2258 (N_2258,In_493,In_1999);
and U2259 (N_2259,In_1650,In_1111);
nor U2260 (N_2260,In_1695,In_1703);
nor U2261 (N_2261,In_1476,In_444);
nand U2262 (N_2262,In_1027,In_886);
nor U2263 (N_2263,In_1570,In_712);
and U2264 (N_2264,In_921,In_1157);
nand U2265 (N_2265,In_672,In_1425);
and U2266 (N_2266,In_1309,In_1325);
or U2267 (N_2267,In_295,In_774);
nand U2268 (N_2268,In_216,In_30);
nand U2269 (N_2269,In_466,In_1488);
xor U2270 (N_2270,In_1568,In_1122);
or U2271 (N_2271,In_1935,In_772);
xnor U2272 (N_2272,In_1125,In_1029);
xnor U2273 (N_2273,In_608,In_267);
nor U2274 (N_2274,In_1859,In_851);
or U2275 (N_2275,In_1694,In_225);
nand U2276 (N_2276,In_877,In_58);
nor U2277 (N_2277,In_1291,In_1212);
nand U2278 (N_2278,In_802,In_1246);
xor U2279 (N_2279,In_152,In_34);
xnor U2280 (N_2280,In_1564,In_484);
nand U2281 (N_2281,In_1470,In_1260);
or U2282 (N_2282,In_739,In_634);
and U2283 (N_2283,In_1417,In_949);
and U2284 (N_2284,In_1695,In_1477);
nor U2285 (N_2285,In_895,In_648);
or U2286 (N_2286,In_1728,In_1453);
or U2287 (N_2287,In_1858,In_1105);
or U2288 (N_2288,In_1223,In_1931);
nor U2289 (N_2289,In_850,In_1674);
or U2290 (N_2290,In_1531,In_1579);
xnor U2291 (N_2291,In_1662,In_1704);
nor U2292 (N_2292,In_692,In_1816);
nand U2293 (N_2293,In_1940,In_73);
nand U2294 (N_2294,In_1289,In_1363);
and U2295 (N_2295,In_1639,In_491);
or U2296 (N_2296,In_1176,In_1507);
or U2297 (N_2297,In_653,In_1683);
xor U2298 (N_2298,In_1234,In_908);
nand U2299 (N_2299,In_1342,In_1695);
xnor U2300 (N_2300,In_1949,In_1415);
or U2301 (N_2301,In_1222,In_1050);
nor U2302 (N_2302,In_75,In_473);
xor U2303 (N_2303,In_1541,In_1048);
xor U2304 (N_2304,In_1832,In_666);
xnor U2305 (N_2305,In_1547,In_1060);
xor U2306 (N_2306,In_857,In_920);
nand U2307 (N_2307,In_1081,In_1628);
and U2308 (N_2308,In_1148,In_1172);
and U2309 (N_2309,In_850,In_754);
xor U2310 (N_2310,In_1215,In_873);
or U2311 (N_2311,In_1960,In_1842);
nand U2312 (N_2312,In_359,In_903);
xor U2313 (N_2313,In_1512,In_1603);
or U2314 (N_2314,In_737,In_59);
xor U2315 (N_2315,In_824,In_1617);
or U2316 (N_2316,In_1203,In_1108);
nor U2317 (N_2317,In_1057,In_683);
or U2318 (N_2318,In_1768,In_1575);
or U2319 (N_2319,In_880,In_398);
nand U2320 (N_2320,In_1358,In_987);
nand U2321 (N_2321,In_1353,In_1694);
xnor U2322 (N_2322,In_380,In_1614);
xor U2323 (N_2323,In_196,In_1834);
and U2324 (N_2324,In_1796,In_1229);
and U2325 (N_2325,In_667,In_1261);
and U2326 (N_2326,In_724,In_233);
nand U2327 (N_2327,In_1554,In_1450);
nand U2328 (N_2328,In_1898,In_678);
or U2329 (N_2329,In_1379,In_1216);
and U2330 (N_2330,In_1657,In_1435);
nand U2331 (N_2331,In_1141,In_1972);
xnor U2332 (N_2332,In_1768,In_111);
and U2333 (N_2333,In_14,In_1493);
and U2334 (N_2334,In_1466,In_1068);
and U2335 (N_2335,In_123,In_581);
nor U2336 (N_2336,In_1674,In_1688);
and U2337 (N_2337,In_135,In_1120);
nor U2338 (N_2338,In_835,In_580);
and U2339 (N_2339,In_1785,In_1712);
or U2340 (N_2340,In_1067,In_908);
or U2341 (N_2341,In_1500,In_1747);
and U2342 (N_2342,In_94,In_1446);
and U2343 (N_2343,In_1682,In_815);
xor U2344 (N_2344,In_79,In_724);
nor U2345 (N_2345,In_210,In_235);
and U2346 (N_2346,In_307,In_747);
nand U2347 (N_2347,In_1977,In_1251);
and U2348 (N_2348,In_1933,In_176);
or U2349 (N_2349,In_605,In_1206);
and U2350 (N_2350,In_1450,In_1110);
and U2351 (N_2351,In_501,In_159);
and U2352 (N_2352,In_1330,In_1575);
nor U2353 (N_2353,In_1302,In_569);
and U2354 (N_2354,In_178,In_30);
nor U2355 (N_2355,In_786,In_1482);
nor U2356 (N_2356,In_139,In_1372);
xnor U2357 (N_2357,In_1573,In_1773);
xor U2358 (N_2358,In_312,In_1801);
xnor U2359 (N_2359,In_606,In_1071);
and U2360 (N_2360,In_1430,In_1606);
and U2361 (N_2361,In_1275,In_35);
xnor U2362 (N_2362,In_453,In_821);
or U2363 (N_2363,In_1174,In_1675);
or U2364 (N_2364,In_1577,In_1552);
xor U2365 (N_2365,In_101,In_1828);
and U2366 (N_2366,In_111,In_1284);
xor U2367 (N_2367,In_673,In_1991);
nor U2368 (N_2368,In_165,In_1972);
nor U2369 (N_2369,In_1696,In_81);
nand U2370 (N_2370,In_1703,In_1737);
and U2371 (N_2371,In_1629,In_1838);
xor U2372 (N_2372,In_539,In_1171);
and U2373 (N_2373,In_826,In_1661);
or U2374 (N_2374,In_1192,In_1932);
nand U2375 (N_2375,In_890,In_1657);
and U2376 (N_2376,In_1886,In_694);
and U2377 (N_2377,In_1792,In_1723);
and U2378 (N_2378,In_887,In_840);
or U2379 (N_2379,In_496,In_1390);
xnor U2380 (N_2380,In_600,In_820);
xnor U2381 (N_2381,In_1058,In_1631);
nand U2382 (N_2382,In_572,In_1954);
or U2383 (N_2383,In_1754,In_782);
or U2384 (N_2384,In_602,In_1264);
nor U2385 (N_2385,In_1578,In_42);
nand U2386 (N_2386,In_1417,In_1941);
or U2387 (N_2387,In_585,In_413);
or U2388 (N_2388,In_997,In_1349);
nand U2389 (N_2389,In_1168,In_1228);
and U2390 (N_2390,In_1851,In_1327);
or U2391 (N_2391,In_548,In_870);
and U2392 (N_2392,In_913,In_716);
nor U2393 (N_2393,In_1390,In_528);
xor U2394 (N_2394,In_697,In_258);
or U2395 (N_2395,In_1563,In_501);
and U2396 (N_2396,In_412,In_131);
xor U2397 (N_2397,In_247,In_546);
xnor U2398 (N_2398,In_908,In_383);
and U2399 (N_2399,In_1794,In_767);
nor U2400 (N_2400,In_1468,In_87);
nand U2401 (N_2401,In_1386,In_202);
xor U2402 (N_2402,In_289,In_504);
nor U2403 (N_2403,In_287,In_936);
or U2404 (N_2404,In_132,In_1442);
xor U2405 (N_2405,In_918,In_245);
or U2406 (N_2406,In_507,In_788);
nor U2407 (N_2407,In_1420,In_628);
nand U2408 (N_2408,In_278,In_1784);
or U2409 (N_2409,In_792,In_1002);
xnor U2410 (N_2410,In_828,In_936);
or U2411 (N_2411,In_260,In_461);
and U2412 (N_2412,In_1549,In_1773);
xor U2413 (N_2413,In_1338,In_240);
and U2414 (N_2414,In_481,In_1405);
nor U2415 (N_2415,In_1004,In_418);
nand U2416 (N_2416,In_726,In_972);
or U2417 (N_2417,In_1978,In_720);
and U2418 (N_2418,In_1896,In_1796);
nor U2419 (N_2419,In_55,In_1019);
xor U2420 (N_2420,In_1795,In_208);
xor U2421 (N_2421,In_1490,In_422);
or U2422 (N_2422,In_1970,In_853);
or U2423 (N_2423,In_1337,In_1146);
or U2424 (N_2424,In_1611,In_1386);
nor U2425 (N_2425,In_1859,In_344);
xor U2426 (N_2426,In_395,In_616);
nor U2427 (N_2427,In_227,In_1398);
and U2428 (N_2428,In_1109,In_703);
xnor U2429 (N_2429,In_1669,In_798);
and U2430 (N_2430,In_9,In_1667);
nand U2431 (N_2431,In_1043,In_1460);
xnor U2432 (N_2432,In_725,In_1715);
and U2433 (N_2433,In_394,In_1130);
nor U2434 (N_2434,In_1306,In_1469);
or U2435 (N_2435,In_256,In_1942);
nor U2436 (N_2436,In_1217,In_710);
xor U2437 (N_2437,In_1063,In_282);
and U2438 (N_2438,In_215,In_539);
nand U2439 (N_2439,In_1907,In_1415);
nor U2440 (N_2440,In_534,In_1024);
xor U2441 (N_2441,In_1844,In_1939);
or U2442 (N_2442,In_1929,In_804);
or U2443 (N_2443,In_1849,In_1252);
xor U2444 (N_2444,In_533,In_1595);
or U2445 (N_2445,In_673,In_1102);
nor U2446 (N_2446,In_343,In_186);
and U2447 (N_2447,In_522,In_1833);
and U2448 (N_2448,In_629,In_1510);
or U2449 (N_2449,In_1244,In_838);
xnor U2450 (N_2450,In_1186,In_1635);
and U2451 (N_2451,In_1248,In_92);
and U2452 (N_2452,In_894,In_1568);
xnor U2453 (N_2453,In_1660,In_1568);
xnor U2454 (N_2454,In_66,In_1271);
nand U2455 (N_2455,In_1576,In_425);
nor U2456 (N_2456,In_1922,In_497);
nor U2457 (N_2457,In_305,In_325);
nor U2458 (N_2458,In_137,In_160);
or U2459 (N_2459,In_1264,In_1773);
or U2460 (N_2460,In_1258,In_34);
nand U2461 (N_2461,In_1838,In_423);
nand U2462 (N_2462,In_501,In_626);
xor U2463 (N_2463,In_1650,In_1160);
and U2464 (N_2464,In_20,In_163);
and U2465 (N_2465,In_140,In_179);
or U2466 (N_2466,In_427,In_332);
nand U2467 (N_2467,In_1508,In_1044);
nand U2468 (N_2468,In_40,In_1308);
nor U2469 (N_2469,In_1275,In_714);
nor U2470 (N_2470,In_1468,In_1510);
or U2471 (N_2471,In_1947,In_859);
and U2472 (N_2472,In_1084,In_808);
or U2473 (N_2473,In_1501,In_1253);
and U2474 (N_2474,In_927,In_464);
and U2475 (N_2475,In_886,In_708);
nor U2476 (N_2476,In_1049,In_1773);
and U2477 (N_2477,In_1805,In_638);
nand U2478 (N_2478,In_792,In_1084);
nor U2479 (N_2479,In_628,In_1486);
nor U2480 (N_2480,In_1524,In_1691);
nor U2481 (N_2481,In_211,In_1780);
or U2482 (N_2482,In_771,In_1491);
nor U2483 (N_2483,In_889,In_1895);
xor U2484 (N_2484,In_1951,In_1684);
and U2485 (N_2485,In_1958,In_71);
nor U2486 (N_2486,In_603,In_1703);
xor U2487 (N_2487,In_1602,In_483);
xor U2488 (N_2488,In_1354,In_409);
nor U2489 (N_2489,In_1385,In_257);
nand U2490 (N_2490,In_712,In_1498);
and U2491 (N_2491,In_1558,In_167);
nand U2492 (N_2492,In_1540,In_157);
and U2493 (N_2493,In_219,In_151);
nor U2494 (N_2494,In_1027,In_70);
and U2495 (N_2495,In_1189,In_675);
or U2496 (N_2496,In_1471,In_873);
nor U2497 (N_2497,In_931,In_805);
xor U2498 (N_2498,In_1746,In_172);
and U2499 (N_2499,In_1003,In_461);
nor U2500 (N_2500,In_1781,In_950);
or U2501 (N_2501,In_1470,In_1762);
nor U2502 (N_2502,In_43,In_1757);
nand U2503 (N_2503,In_1040,In_1716);
and U2504 (N_2504,In_1116,In_929);
or U2505 (N_2505,In_1536,In_448);
or U2506 (N_2506,In_534,In_732);
nor U2507 (N_2507,In_1239,In_1025);
or U2508 (N_2508,In_1153,In_1442);
xor U2509 (N_2509,In_1219,In_1935);
and U2510 (N_2510,In_1051,In_697);
xor U2511 (N_2511,In_777,In_1620);
and U2512 (N_2512,In_1998,In_1834);
and U2513 (N_2513,In_818,In_777);
or U2514 (N_2514,In_1826,In_94);
and U2515 (N_2515,In_1226,In_1633);
nor U2516 (N_2516,In_806,In_501);
nand U2517 (N_2517,In_33,In_1624);
nor U2518 (N_2518,In_1082,In_517);
nor U2519 (N_2519,In_244,In_447);
xnor U2520 (N_2520,In_988,In_1312);
nand U2521 (N_2521,In_1812,In_1791);
nor U2522 (N_2522,In_506,In_1361);
nor U2523 (N_2523,In_125,In_1639);
nand U2524 (N_2524,In_1580,In_241);
and U2525 (N_2525,In_527,In_1030);
xnor U2526 (N_2526,In_636,In_1514);
nand U2527 (N_2527,In_1730,In_425);
and U2528 (N_2528,In_536,In_638);
xor U2529 (N_2529,In_152,In_1624);
nand U2530 (N_2530,In_1490,In_687);
and U2531 (N_2531,In_1048,In_689);
or U2532 (N_2532,In_235,In_1934);
nand U2533 (N_2533,In_1494,In_48);
or U2534 (N_2534,In_727,In_699);
or U2535 (N_2535,In_1657,In_1555);
nand U2536 (N_2536,In_346,In_855);
nor U2537 (N_2537,In_219,In_1139);
or U2538 (N_2538,In_528,In_1820);
or U2539 (N_2539,In_630,In_1354);
or U2540 (N_2540,In_1239,In_1482);
and U2541 (N_2541,In_614,In_12);
or U2542 (N_2542,In_1894,In_1508);
nor U2543 (N_2543,In_1171,In_1792);
or U2544 (N_2544,In_332,In_483);
nor U2545 (N_2545,In_1199,In_1928);
or U2546 (N_2546,In_676,In_458);
or U2547 (N_2547,In_507,In_1978);
and U2548 (N_2548,In_1983,In_748);
or U2549 (N_2549,In_1798,In_1238);
xor U2550 (N_2550,In_1190,In_1488);
xnor U2551 (N_2551,In_1775,In_1569);
xor U2552 (N_2552,In_364,In_10);
xnor U2553 (N_2553,In_1482,In_1830);
nand U2554 (N_2554,In_568,In_695);
or U2555 (N_2555,In_1859,In_517);
and U2556 (N_2556,In_1110,In_1052);
or U2557 (N_2557,In_1615,In_113);
nand U2558 (N_2558,In_670,In_487);
xor U2559 (N_2559,In_661,In_894);
xor U2560 (N_2560,In_255,In_1843);
and U2561 (N_2561,In_1886,In_1325);
or U2562 (N_2562,In_1399,In_239);
nand U2563 (N_2563,In_658,In_539);
nand U2564 (N_2564,In_137,In_73);
and U2565 (N_2565,In_291,In_1867);
and U2566 (N_2566,In_1915,In_1085);
xor U2567 (N_2567,In_387,In_1674);
nor U2568 (N_2568,In_1759,In_1240);
or U2569 (N_2569,In_712,In_876);
nand U2570 (N_2570,In_72,In_1545);
nor U2571 (N_2571,In_1766,In_277);
or U2572 (N_2572,In_1696,In_673);
and U2573 (N_2573,In_1975,In_267);
or U2574 (N_2574,In_507,In_1906);
or U2575 (N_2575,In_1012,In_1046);
nor U2576 (N_2576,In_112,In_1401);
nand U2577 (N_2577,In_209,In_1435);
and U2578 (N_2578,In_1884,In_1515);
xnor U2579 (N_2579,In_1715,In_23);
xnor U2580 (N_2580,In_254,In_1794);
or U2581 (N_2581,In_206,In_1780);
nor U2582 (N_2582,In_1258,In_1091);
nor U2583 (N_2583,In_1953,In_1073);
or U2584 (N_2584,In_529,In_1166);
or U2585 (N_2585,In_1047,In_1649);
or U2586 (N_2586,In_1506,In_1846);
xor U2587 (N_2587,In_813,In_1226);
nand U2588 (N_2588,In_1480,In_1872);
and U2589 (N_2589,In_1618,In_942);
nor U2590 (N_2590,In_176,In_1426);
xor U2591 (N_2591,In_585,In_1288);
and U2592 (N_2592,In_199,In_1738);
nand U2593 (N_2593,In_1809,In_281);
nand U2594 (N_2594,In_1882,In_565);
and U2595 (N_2595,In_160,In_589);
and U2596 (N_2596,In_822,In_1506);
xnor U2597 (N_2597,In_1228,In_194);
nand U2598 (N_2598,In_1131,In_1187);
nand U2599 (N_2599,In_468,In_101);
and U2600 (N_2600,In_1296,In_1483);
and U2601 (N_2601,In_1171,In_292);
nand U2602 (N_2602,In_874,In_1382);
nor U2603 (N_2603,In_336,In_894);
nor U2604 (N_2604,In_841,In_1952);
and U2605 (N_2605,In_1747,In_292);
and U2606 (N_2606,In_608,In_129);
xnor U2607 (N_2607,In_1983,In_693);
xor U2608 (N_2608,In_550,In_1942);
and U2609 (N_2609,In_85,In_876);
nand U2610 (N_2610,In_1786,In_1516);
xor U2611 (N_2611,In_887,In_1279);
nand U2612 (N_2612,In_1987,In_1120);
nand U2613 (N_2613,In_1108,In_815);
xnor U2614 (N_2614,In_227,In_684);
xor U2615 (N_2615,In_1697,In_1849);
nor U2616 (N_2616,In_1037,In_720);
xor U2617 (N_2617,In_392,In_774);
or U2618 (N_2618,In_1180,In_1780);
xnor U2619 (N_2619,In_173,In_152);
or U2620 (N_2620,In_1692,In_788);
xor U2621 (N_2621,In_1311,In_1257);
nor U2622 (N_2622,In_1773,In_1980);
nor U2623 (N_2623,In_1610,In_1201);
and U2624 (N_2624,In_854,In_1957);
or U2625 (N_2625,In_1287,In_501);
nor U2626 (N_2626,In_574,In_1330);
or U2627 (N_2627,In_1328,In_1792);
or U2628 (N_2628,In_1455,In_1713);
nor U2629 (N_2629,In_1926,In_283);
nor U2630 (N_2630,In_420,In_494);
nand U2631 (N_2631,In_411,In_1532);
xnor U2632 (N_2632,In_477,In_1766);
nand U2633 (N_2633,In_421,In_326);
and U2634 (N_2634,In_88,In_1378);
nand U2635 (N_2635,In_1645,In_1139);
and U2636 (N_2636,In_1572,In_1494);
nor U2637 (N_2637,In_1561,In_790);
and U2638 (N_2638,In_716,In_416);
or U2639 (N_2639,In_1752,In_1467);
nand U2640 (N_2640,In_1573,In_266);
or U2641 (N_2641,In_882,In_1345);
nor U2642 (N_2642,In_824,In_224);
nand U2643 (N_2643,In_47,In_1378);
and U2644 (N_2644,In_1036,In_1026);
nand U2645 (N_2645,In_661,In_432);
xnor U2646 (N_2646,In_50,In_1719);
nand U2647 (N_2647,In_94,In_1210);
and U2648 (N_2648,In_688,In_909);
nor U2649 (N_2649,In_610,In_921);
xnor U2650 (N_2650,In_1754,In_1464);
xor U2651 (N_2651,In_1984,In_257);
and U2652 (N_2652,In_1737,In_1255);
xor U2653 (N_2653,In_770,In_883);
or U2654 (N_2654,In_796,In_1985);
xnor U2655 (N_2655,In_243,In_1585);
xor U2656 (N_2656,In_3,In_977);
xnor U2657 (N_2657,In_1597,In_124);
or U2658 (N_2658,In_471,In_1068);
nor U2659 (N_2659,In_1901,In_693);
and U2660 (N_2660,In_629,In_1174);
and U2661 (N_2661,In_1297,In_1989);
or U2662 (N_2662,In_532,In_8);
xnor U2663 (N_2663,In_790,In_535);
nor U2664 (N_2664,In_1586,In_62);
nor U2665 (N_2665,In_379,In_1047);
nand U2666 (N_2666,In_675,In_470);
nor U2667 (N_2667,In_1596,In_991);
nand U2668 (N_2668,In_590,In_381);
and U2669 (N_2669,In_960,In_566);
nor U2670 (N_2670,In_248,In_1154);
nand U2671 (N_2671,In_1789,In_1458);
nand U2672 (N_2672,In_1471,In_571);
nand U2673 (N_2673,In_1428,In_141);
nand U2674 (N_2674,In_1294,In_1345);
nand U2675 (N_2675,In_590,In_969);
or U2676 (N_2676,In_1683,In_631);
xnor U2677 (N_2677,In_1150,In_1534);
nor U2678 (N_2678,In_257,In_813);
and U2679 (N_2679,In_256,In_1382);
nor U2680 (N_2680,In_69,In_1456);
xor U2681 (N_2681,In_1175,In_905);
or U2682 (N_2682,In_1079,In_1959);
nand U2683 (N_2683,In_1865,In_1528);
and U2684 (N_2684,In_189,In_249);
xor U2685 (N_2685,In_215,In_1036);
xnor U2686 (N_2686,In_1873,In_1428);
nor U2687 (N_2687,In_1896,In_516);
or U2688 (N_2688,In_1061,In_1102);
and U2689 (N_2689,In_184,In_927);
nand U2690 (N_2690,In_169,In_772);
xnor U2691 (N_2691,In_1850,In_1302);
xnor U2692 (N_2692,In_1824,In_717);
nor U2693 (N_2693,In_1658,In_1586);
nand U2694 (N_2694,In_1578,In_1496);
nand U2695 (N_2695,In_1793,In_1231);
or U2696 (N_2696,In_642,In_298);
nand U2697 (N_2697,In_1570,In_1697);
nand U2698 (N_2698,In_1520,In_1042);
nor U2699 (N_2699,In_425,In_1804);
or U2700 (N_2700,In_1985,In_284);
nand U2701 (N_2701,In_723,In_1074);
xor U2702 (N_2702,In_835,In_1504);
or U2703 (N_2703,In_1470,In_1315);
nor U2704 (N_2704,In_213,In_1033);
and U2705 (N_2705,In_1755,In_868);
xnor U2706 (N_2706,In_54,In_1522);
xor U2707 (N_2707,In_1876,In_148);
nand U2708 (N_2708,In_764,In_930);
nand U2709 (N_2709,In_1536,In_410);
nor U2710 (N_2710,In_1936,In_543);
nand U2711 (N_2711,In_554,In_915);
nor U2712 (N_2712,In_836,In_734);
xor U2713 (N_2713,In_1469,In_95);
and U2714 (N_2714,In_1026,In_1516);
and U2715 (N_2715,In_409,In_1055);
or U2716 (N_2716,In_513,In_347);
xnor U2717 (N_2717,In_208,In_541);
and U2718 (N_2718,In_1843,In_874);
and U2719 (N_2719,In_47,In_162);
xor U2720 (N_2720,In_419,In_842);
xnor U2721 (N_2721,In_908,In_1298);
or U2722 (N_2722,In_1161,In_1353);
xor U2723 (N_2723,In_124,In_1843);
nand U2724 (N_2724,In_660,In_986);
nor U2725 (N_2725,In_214,In_570);
nor U2726 (N_2726,In_1893,In_1584);
or U2727 (N_2727,In_1487,In_456);
nand U2728 (N_2728,In_389,In_1435);
or U2729 (N_2729,In_1220,In_561);
and U2730 (N_2730,In_1016,In_48);
nor U2731 (N_2731,In_1364,In_1981);
nor U2732 (N_2732,In_1140,In_767);
nor U2733 (N_2733,In_1034,In_56);
nor U2734 (N_2734,In_1293,In_153);
or U2735 (N_2735,In_1233,In_1060);
nor U2736 (N_2736,In_768,In_107);
and U2737 (N_2737,In_569,In_1666);
xor U2738 (N_2738,In_50,In_1952);
and U2739 (N_2739,In_129,In_324);
and U2740 (N_2740,In_777,In_1550);
or U2741 (N_2741,In_1641,In_1783);
or U2742 (N_2742,In_1874,In_86);
or U2743 (N_2743,In_1630,In_1970);
and U2744 (N_2744,In_684,In_1450);
and U2745 (N_2745,In_764,In_1208);
xnor U2746 (N_2746,In_1137,In_1984);
xor U2747 (N_2747,In_1667,In_257);
nand U2748 (N_2748,In_1577,In_531);
xor U2749 (N_2749,In_1214,In_1546);
nand U2750 (N_2750,In_358,In_899);
or U2751 (N_2751,In_1749,In_1792);
xor U2752 (N_2752,In_1602,In_1856);
or U2753 (N_2753,In_1060,In_548);
and U2754 (N_2754,In_1168,In_411);
and U2755 (N_2755,In_338,In_723);
or U2756 (N_2756,In_656,In_126);
xor U2757 (N_2757,In_1445,In_765);
and U2758 (N_2758,In_841,In_1936);
or U2759 (N_2759,In_859,In_362);
nor U2760 (N_2760,In_1694,In_107);
and U2761 (N_2761,In_1633,In_237);
nand U2762 (N_2762,In_1502,In_353);
and U2763 (N_2763,In_1014,In_1833);
or U2764 (N_2764,In_1283,In_0);
or U2765 (N_2765,In_633,In_1813);
nor U2766 (N_2766,In_1565,In_546);
xnor U2767 (N_2767,In_1547,In_1446);
nand U2768 (N_2768,In_1660,In_1993);
nand U2769 (N_2769,In_742,In_1562);
xnor U2770 (N_2770,In_1684,In_827);
nand U2771 (N_2771,In_1079,In_609);
nand U2772 (N_2772,In_1337,In_200);
and U2773 (N_2773,In_1932,In_375);
xnor U2774 (N_2774,In_1787,In_404);
xnor U2775 (N_2775,In_216,In_1828);
nor U2776 (N_2776,In_297,In_1562);
or U2777 (N_2777,In_330,In_1268);
nand U2778 (N_2778,In_1142,In_1074);
xnor U2779 (N_2779,In_1434,In_1285);
nor U2780 (N_2780,In_585,In_217);
nor U2781 (N_2781,In_1147,In_524);
and U2782 (N_2782,In_875,In_262);
nor U2783 (N_2783,In_1367,In_906);
and U2784 (N_2784,In_281,In_726);
nand U2785 (N_2785,In_1055,In_872);
nand U2786 (N_2786,In_703,In_1774);
xor U2787 (N_2787,In_1872,In_735);
or U2788 (N_2788,In_1777,In_1287);
xnor U2789 (N_2789,In_605,In_1556);
xnor U2790 (N_2790,In_1882,In_130);
or U2791 (N_2791,In_1922,In_1657);
nor U2792 (N_2792,In_770,In_18);
nand U2793 (N_2793,In_946,In_1160);
or U2794 (N_2794,In_286,In_704);
xor U2795 (N_2795,In_1567,In_1981);
nor U2796 (N_2796,In_1021,In_493);
or U2797 (N_2797,In_1750,In_1316);
nor U2798 (N_2798,In_72,In_1626);
xor U2799 (N_2799,In_692,In_1983);
nor U2800 (N_2800,In_1735,In_371);
and U2801 (N_2801,In_1315,In_118);
and U2802 (N_2802,In_1734,In_1548);
nand U2803 (N_2803,In_1535,In_9);
nand U2804 (N_2804,In_1607,In_1158);
nor U2805 (N_2805,In_408,In_697);
or U2806 (N_2806,In_1456,In_1643);
or U2807 (N_2807,In_146,In_1001);
or U2808 (N_2808,In_589,In_1238);
nor U2809 (N_2809,In_1812,In_1627);
and U2810 (N_2810,In_1418,In_671);
xor U2811 (N_2811,In_1571,In_1987);
or U2812 (N_2812,In_923,In_1945);
xnor U2813 (N_2813,In_1824,In_529);
xor U2814 (N_2814,In_171,In_1870);
xor U2815 (N_2815,In_1561,In_1908);
and U2816 (N_2816,In_1967,In_705);
nand U2817 (N_2817,In_109,In_1676);
nor U2818 (N_2818,In_845,In_1218);
nand U2819 (N_2819,In_1301,In_1639);
xor U2820 (N_2820,In_557,In_881);
and U2821 (N_2821,In_54,In_1529);
nand U2822 (N_2822,In_1490,In_971);
xor U2823 (N_2823,In_1774,In_986);
nand U2824 (N_2824,In_1457,In_1921);
xor U2825 (N_2825,In_890,In_1742);
and U2826 (N_2826,In_150,In_1002);
xnor U2827 (N_2827,In_1697,In_860);
nor U2828 (N_2828,In_1761,In_686);
or U2829 (N_2829,In_377,In_1808);
nand U2830 (N_2830,In_156,In_1876);
or U2831 (N_2831,In_1492,In_687);
nor U2832 (N_2832,In_1080,In_716);
xor U2833 (N_2833,In_804,In_171);
or U2834 (N_2834,In_112,In_1364);
xnor U2835 (N_2835,In_860,In_1875);
and U2836 (N_2836,In_1314,In_1865);
and U2837 (N_2837,In_1377,In_535);
xnor U2838 (N_2838,In_35,In_828);
nand U2839 (N_2839,In_224,In_1613);
and U2840 (N_2840,In_704,In_361);
or U2841 (N_2841,In_819,In_1211);
xnor U2842 (N_2842,In_1858,In_1993);
nand U2843 (N_2843,In_819,In_1943);
xor U2844 (N_2844,In_320,In_97);
nand U2845 (N_2845,In_284,In_59);
nand U2846 (N_2846,In_1726,In_1340);
nor U2847 (N_2847,In_182,In_787);
nor U2848 (N_2848,In_1508,In_1847);
xnor U2849 (N_2849,In_1763,In_677);
or U2850 (N_2850,In_1646,In_486);
nor U2851 (N_2851,In_1696,In_1576);
and U2852 (N_2852,In_1128,In_1345);
or U2853 (N_2853,In_1736,In_454);
or U2854 (N_2854,In_1077,In_1831);
and U2855 (N_2855,In_1808,In_1409);
xor U2856 (N_2856,In_924,In_594);
xor U2857 (N_2857,In_57,In_649);
nor U2858 (N_2858,In_625,In_414);
xnor U2859 (N_2859,In_537,In_287);
and U2860 (N_2860,In_634,In_1116);
and U2861 (N_2861,In_1000,In_804);
nor U2862 (N_2862,In_447,In_210);
nor U2863 (N_2863,In_1284,In_1669);
xor U2864 (N_2864,In_577,In_345);
or U2865 (N_2865,In_839,In_259);
and U2866 (N_2866,In_849,In_1051);
and U2867 (N_2867,In_164,In_748);
nand U2868 (N_2868,In_1023,In_82);
nor U2869 (N_2869,In_1459,In_1326);
xor U2870 (N_2870,In_1418,In_349);
or U2871 (N_2871,In_1731,In_905);
xnor U2872 (N_2872,In_689,In_93);
or U2873 (N_2873,In_143,In_1436);
and U2874 (N_2874,In_488,In_521);
and U2875 (N_2875,In_536,In_1792);
nor U2876 (N_2876,In_1640,In_1190);
nor U2877 (N_2877,In_229,In_81);
xnor U2878 (N_2878,In_1788,In_648);
or U2879 (N_2879,In_1682,In_494);
or U2880 (N_2880,In_1162,In_207);
and U2881 (N_2881,In_1236,In_1582);
or U2882 (N_2882,In_89,In_1457);
and U2883 (N_2883,In_532,In_444);
or U2884 (N_2884,In_61,In_1572);
and U2885 (N_2885,In_581,In_75);
nand U2886 (N_2886,In_1782,In_774);
nand U2887 (N_2887,In_1422,In_1293);
xor U2888 (N_2888,In_1738,In_1149);
and U2889 (N_2889,In_1337,In_504);
or U2890 (N_2890,In_1146,In_469);
xor U2891 (N_2891,In_151,In_1989);
nor U2892 (N_2892,In_1125,In_435);
nor U2893 (N_2893,In_1257,In_657);
xor U2894 (N_2894,In_694,In_884);
or U2895 (N_2895,In_1437,In_146);
or U2896 (N_2896,In_1543,In_655);
and U2897 (N_2897,In_1724,In_260);
nor U2898 (N_2898,In_1302,In_1992);
xnor U2899 (N_2899,In_53,In_1763);
xor U2900 (N_2900,In_1736,In_1741);
or U2901 (N_2901,In_351,In_1853);
nand U2902 (N_2902,In_54,In_1618);
or U2903 (N_2903,In_720,In_743);
and U2904 (N_2904,In_1828,In_1374);
xnor U2905 (N_2905,In_1590,In_1798);
xnor U2906 (N_2906,In_153,In_695);
xor U2907 (N_2907,In_360,In_1412);
and U2908 (N_2908,In_482,In_1125);
xnor U2909 (N_2909,In_1234,In_121);
xor U2910 (N_2910,In_1815,In_243);
nor U2911 (N_2911,In_1780,In_1159);
xor U2912 (N_2912,In_745,In_126);
nand U2913 (N_2913,In_1896,In_1742);
or U2914 (N_2914,In_92,In_567);
nor U2915 (N_2915,In_1187,In_907);
and U2916 (N_2916,In_898,In_900);
nand U2917 (N_2917,In_1753,In_320);
xnor U2918 (N_2918,In_1500,In_1554);
and U2919 (N_2919,In_975,In_1983);
xnor U2920 (N_2920,In_1468,In_1665);
and U2921 (N_2921,In_292,In_821);
nand U2922 (N_2922,In_266,In_388);
and U2923 (N_2923,In_1253,In_1319);
xnor U2924 (N_2924,In_166,In_1924);
and U2925 (N_2925,In_428,In_1970);
xor U2926 (N_2926,In_1869,In_415);
and U2927 (N_2927,In_353,In_984);
or U2928 (N_2928,In_1830,In_1893);
and U2929 (N_2929,In_1358,In_547);
or U2930 (N_2930,In_1669,In_762);
nand U2931 (N_2931,In_1073,In_723);
xnor U2932 (N_2932,In_636,In_398);
nor U2933 (N_2933,In_1909,In_1276);
nand U2934 (N_2934,In_1038,In_1317);
nor U2935 (N_2935,In_1180,In_1181);
nand U2936 (N_2936,In_176,In_982);
or U2937 (N_2937,In_835,In_264);
xnor U2938 (N_2938,In_1711,In_1353);
nor U2939 (N_2939,In_1472,In_358);
xor U2940 (N_2940,In_493,In_684);
nor U2941 (N_2941,In_963,In_245);
nor U2942 (N_2942,In_1384,In_1070);
xor U2943 (N_2943,In_1559,In_80);
and U2944 (N_2944,In_1140,In_87);
nand U2945 (N_2945,In_1704,In_128);
nand U2946 (N_2946,In_857,In_1208);
and U2947 (N_2947,In_1902,In_2);
nand U2948 (N_2948,In_1083,In_1458);
nor U2949 (N_2949,In_1340,In_1498);
and U2950 (N_2950,In_1470,In_1397);
and U2951 (N_2951,In_479,In_77);
nor U2952 (N_2952,In_644,In_414);
xor U2953 (N_2953,In_346,In_1409);
nand U2954 (N_2954,In_445,In_1347);
xor U2955 (N_2955,In_1849,In_1718);
and U2956 (N_2956,In_930,In_369);
and U2957 (N_2957,In_1541,In_395);
and U2958 (N_2958,In_1126,In_1283);
or U2959 (N_2959,In_288,In_767);
xnor U2960 (N_2960,In_1346,In_1167);
nor U2961 (N_2961,In_90,In_1799);
nand U2962 (N_2962,In_673,In_1464);
nor U2963 (N_2963,In_1996,In_463);
nor U2964 (N_2964,In_1633,In_818);
or U2965 (N_2965,In_397,In_828);
and U2966 (N_2966,In_1207,In_324);
xnor U2967 (N_2967,In_28,In_937);
and U2968 (N_2968,In_1751,In_1836);
nand U2969 (N_2969,In_821,In_72);
xnor U2970 (N_2970,In_835,In_1789);
nor U2971 (N_2971,In_1684,In_440);
and U2972 (N_2972,In_1699,In_792);
nand U2973 (N_2973,In_1083,In_615);
and U2974 (N_2974,In_1031,In_1992);
nor U2975 (N_2975,In_1911,In_1419);
nand U2976 (N_2976,In_111,In_1090);
nand U2977 (N_2977,In_175,In_1292);
nor U2978 (N_2978,In_918,In_1406);
or U2979 (N_2979,In_1261,In_635);
or U2980 (N_2980,In_1299,In_1609);
nand U2981 (N_2981,In_33,In_1375);
nand U2982 (N_2982,In_1915,In_189);
xnor U2983 (N_2983,In_1362,In_418);
nand U2984 (N_2984,In_961,In_91);
nor U2985 (N_2985,In_808,In_234);
nand U2986 (N_2986,In_1740,In_25);
and U2987 (N_2987,In_648,In_1497);
or U2988 (N_2988,In_693,In_1803);
nor U2989 (N_2989,In_1729,In_889);
or U2990 (N_2990,In_1585,In_344);
and U2991 (N_2991,In_1372,In_947);
and U2992 (N_2992,In_1806,In_1392);
and U2993 (N_2993,In_1764,In_377);
or U2994 (N_2994,In_1531,In_41);
nor U2995 (N_2995,In_38,In_789);
and U2996 (N_2996,In_572,In_1828);
and U2997 (N_2997,In_198,In_1544);
nand U2998 (N_2998,In_1087,In_307);
or U2999 (N_2999,In_1418,In_1996);
nand U3000 (N_3000,In_1508,In_1262);
and U3001 (N_3001,In_1008,In_487);
or U3002 (N_3002,In_1844,In_1471);
or U3003 (N_3003,In_129,In_1479);
nor U3004 (N_3004,In_1555,In_1339);
or U3005 (N_3005,In_89,In_81);
nand U3006 (N_3006,In_1131,In_350);
and U3007 (N_3007,In_928,In_1082);
and U3008 (N_3008,In_654,In_593);
or U3009 (N_3009,In_1134,In_571);
and U3010 (N_3010,In_718,In_237);
or U3011 (N_3011,In_1059,In_283);
or U3012 (N_3012,In_1445,In_965);
or U3013 (N_3013,In_1404,In_320);
nor U3014 (N_3014,In_1818,In_1657);
and U3015 (N_3015,In_105,In_1768);
xor U3016 (N_3016,In_18,In_814);
and U3017 (N_3017,In_943,In_1362);
xnor U3018 (N_3018,In_121,In_1576);
or U3019 (N_3019,In_308,In_1253);
nor U3020 (N_3020,In_566,In_1617);
nand U3021 (N_3021,In_1699,In_1618);
nor U3022 (N_3022,In_893,In_729);
nor U3023 (N_3023,In_1813,In_595);
and U3024 (N_3024,In_414,In_1940);
nand U3025 (N_3025,In_1169,In_1512);
nand U3026 (N_3026,In_996,In_1934);
nor U3027 (N_3027,In_240,In_964);
or U3028 (N_3028,In_1902,In_1247);
nor U3029 (N_3029,In_1395,In_1660);
and U3030 (N_3030,In_1125,In_735);
nand U3031 (N_3031,In_1371,In_47);
nor U3032 (N_3032,In_433,In_1209);
xor U3033 (N_3033,In_1245,In_275);
nor U3034 (N_3034,In_1291,In_1957);
nor U3035 (N_3035,In_1284,In_580);
or U3036 (N_3036,In_1570,In_848);
or U3037 (N_3037,In_803,In_1515);
xor U3038 (N_3038,In_1674,In_1086);
nor U3039 (N_3039,In_1816,In_1824);
xnor U3040 (N_3040,In_255,In_338);
nand U3041 (N_3041,In_992,In_1962);
or U3042 (N_3042,In_607,In_1019);
nor U3043 (N_3043,In_1644,In_335);
nor U3044 (N_3044,In_1531,In_1940);
xnor U3045 (N_3045,In_1991,In_1720);
or U3046 (N_3046,In_669,In_637);
or U3047 (N_3047,In_801,In_439);
xor U3048 (N_3048,In_300,In_542);
xnor U3049 (N_3049,In_1131,In_28);
or U3050 (N_3050,In_1399,In_692);
and U3051 (N_3051,In_1039,In_737);
nand U3052 (N_3052,In_155,In_1902);
nor U3053 (N_3053,In_1352,In_452);
or U3054 (N_3054,In_1218,In_597);
and U3055 (N_3055,In_1735,In_845);
xor U3056 (N_3056,In_1058,In_1125);
and U3057 (N_3057,In_861,In_1272);
nand U3058 (N_3058,In_112,In_650);
xnor U3059 (N_3059,In_1390,In_383);
nor U3060 (N_3060,In_600,In_322);
xor U3061 (N_3061,In_1600,In_1926);
nor U3062 (N_3062,In_652,In_1848);
nand U3063 (N_3063,In_152,In_1135);
and U3064 (N_3064,In_840,In_316);
or U3065 (N_3065,In_601,In_811);
or U3066 (N_3066,In_470,In_483);
or U3067 (N_3067,In_302,In_1499);
and U3068 (N_3068,In_1207,In_672);
or U3069 (N_3069,In_1404,In_688);
and U3070 (N_3070,In_634,In_1962);
and U3071 (N_3071,In_548,In_1959);
nor U3072 (N_3072,In_1614,In_1959);
and U3073 (N_3073,In_1963,In_590);
nand U3074 (N_3074,In_1918,In_289);
nand U3075 (N_3075,In_1476,In_1290);
xnor U3076 (N_3076,In_1606,In_1313);
or U3077 (N_3077,In_1606,In_908);
or U3078 (N_3078,In_1381,In_334);
or U3079 (N_3079,In_757,In_822);
and U3080 (N_3080,In_1611,In_407);
or U3081 (N_3081,In_1955,In_1587);
nor U3082 (N_3082,In_488,In_721);
xor U3083 (N_3083,In_527,In_1356);
xnor U3084 (N_3084,In_1575,In_850);
xor U3085 (N_3085,In_1444,In_264);
xnor U3086 (N_3086,In_326,In_933);
nand U3087 (N_3087,In_1104,In_103);
xor U3088 (N_3088,In_1200,In_932);
nor U3089 (N_3089,In_1877,In_1725);
nor U3090 (N_3090,In_981,In_255);
or U3091 (N_3091,In_981,In_1596);
nor U3092 (N_3092,In_963,In_863);
or U3093 (N_3093,In_77,In_1749);
xnor U3094 (N_3094,In_1342,In_993);
nor U3095 (N_3095,In_108,In_1241);
and U3096 (N_3096,In_1246,In_1024);
nor U3097 (N_3097,In_910,In_1126);
or U3098 (N_3098,In_1227,In_388);
or U3099 (N_3099,In_1396,In_384);
and U3100 (N_3100,In_1827,In_1742);
or U3101 (N_3101,In_573,In_1121);
or U3102 (N_3102,In_212,In_1621);
nor U3103 (N_3103,In_218,In_645);
or U3104 (N_3104,In_181,In_80);
or U3105 (N_3105,In_1526,In_532);
or U3106 (N_3106,In_902,In_1657);
or U3107 (N_3107,In_1909,In_1487);
nor U3108 (N_3108,In_1342,In_1512);
xnor U3109 (N_3109,In_1247,In_1672);
xnor U3110 (N_3110,In_1023,In_1239);
xnor U3111 (N_3111,In_427,In_265);
and U3112 (N_3112,In_1064,In_1463);
and U3113 (N_3113,In_1208,In_1081);
xor U3114 (N_3114,In_286,In_499);
xor U3115 (N_3115,In_1025,In_41);
nand U3116 (N_3116,In_197,In_1473);
nand U3117 (N_3117,In_324,In_610);
nor U3118 (N_3118,In_277,In_952);
nor U3119 (N_3119,In_749,In_1563);
xor U3120 (N_3120,In_1599,In_1322);
nand U3121 (N_3121,In_1594,In_1210);
or U3122 (N_3122,In_814,In_499);
or U3123 (N_3123,In_1876,In_516);
and U3124 (N_3124,In_759,In_74);
xor U3125 (N_3125,In_570,In_1332);
and U3126 (N_3126,In_487,In_969);
nor U3127 (N_3127,In_1116,In_1954);
xor U3128 (N_3128,In_1004,In_1910);
or U3129 (N_3129,In_527,In_1803);
or U3130 (N_3130,In_348,In_575);
xnor U3131 (N_3131,In_809,In_316);
or U3132 (N_3132,In_870,In_105);
nor U3133 (N_3133,In_1915,In_1745);
nand U3134 (N_3134,In_1803,In_531);
or U3135 (N_3135,In_1797,In_1849);
or U3136 (N_3136,In_648,In_1138);
nor U3137 (N_3137,In_714,In_1610);
and U3138 (N_3138,In_1050,In_1017);
nand U3139 (N_3139,In_118,In_1295);
nor U3140 (N_3140,In_1085,In_197);
and U3141 (N_3141,In_962,In_1334);
nand U3142 (N_3142,In_408,In_456);
nor U3143 (N_3143,In_1153,In_1671);
nor U3144 (N_3144,In_1171,In_499);
nor U3145 (N_3145,In_1667,In_538);
or U3146 (N_3146,In_1631,In_492);
nor U3147 (N_3147,In_1890,In_1521);
or U3148 (N_3148,In_701,In_1742);
nand U3149 (N_3149,In_420,In_1254);
nor U3150 (N_3150,In_1823,In_245);
xor U3151 (N_3151,In_699,In_1949);
nand U3152 (N_3152,In_787,In_1806);
or U3153 (N_3153,In_1026,In_1723);
or U3154 (N_3154,In_788,In_1380);
nand U3155 (N_3155,In_130,In_831);
xnor U3156 (N_3156,In_189,In_1971);
or U3157 (N_3157,In_719,In_843);
xor U3158 (N_3158,In_1001,In_1716);
xnor U3159 (N_3159,In_1200,In_1466);
and U3160 (N_3160,In_304,In_949);
nor U3161 (N_3161,In_232,In_1433);
xnor U3162 (N_3162,In_210,In_1825);
nand U3163 (N_3163,In_1074,In_315);
and U3164 (N_3164,In_898,In_433);
and U3165 (N_3165,In_1875,In_1020);
nand U3166 (N_3166,In_811,In_803);
and U3167 (N_3167,In_404,In_610);
nor U3168 (N_3168,In_1434,In_104);
nand U3169 (N_3169,In_1394,In_275);
and U3170 (N_3170,In_244,In_1580);
nor U3171 (N_3171,In_1950,In_583);
and U3172 (N_3172,In_1085,In_707);
nand U3173 (N_3173,In_327,In_767);
nand U3174 (N_3174,In_1545,In_1735);
or U3175 (N_3175,In_1245,In_778);
or U3176 (N_3176,In_903,In_18);
and U3177 (N_3177,In_1975,In_1681);
xnor U3178 (N_3178,In_6,In_1550);
or U3179 (N_3179,In_57,In_1843);
and U3180 (N_3180,In_387,In_359);
xnor U3181 (N_3181,In_1433,In_833);
nand U3182 (N_3182,In_1708,In_885);
nand U3183 (N_3183,In_1816,In_916);
nor U3184 (N_3184,In_1238,In_588);
and U3185 (N_3185,In_1490,In_317);
nor U3186 (N_3186,In_354,In_1188);
nand U3187 (N_3187,In_207,In_1679);
nor U3188 (N_3188,In_1108,In_135);
nand U3189 (N_3189,In_1260,In_1886);
and U3190 (N_3190,In_252,In_738);
nor U3191 (N_3191,In_1830,In_925);
and U3192 (N_3192,In_1780,In_921);
xor U3193 (N_3193,In_1979,In_1320);
or U3194 (N_3194,In_1545,In_396);
xor U3195 (N_3195,In_203,In_818);
nor U3196 (N_3196,In_1314,In_914);
xor U3197 (N_3197,In_26,In_280);
nor U3198 (N_3198,In_1989,In_1570);
nor U3199 (N_3199,In_561,In_1753);
nor U3200 (N_3200,In_1825,In_1264);
nand U3201 (N_3201,In_1298,In_1478);
xor U3202 (N_3202,In_1004,In_1653);
nand U3203 (N_3203,In_1851,In_211);
or U3204 (N_3204,In_642,In_71);
xnor U3205 (N_3205,In_1360,In_1736);
nor U3206 (N_3206,In_1961,In_295);
or U3207 (N_3207,In_1192,In_571);
or U3208 (N_3208,In_959,In_751);
xor U3209 (N_3209,In_607,In_1551);
nor U3210 (N_3210,In_1955,In_262);
and U3211 (N_3211,In_769,In_290);
nand U3212 (N_3212,In_1125,In_1660);
or U3213 (N_3213,In_1661,In_788);
nand U3214 (N_3214,In_335,In_839);
nand U3215 (N_3215,In_1608,In_997);
nor U3216 (N_3216,In_627,In_1998);
and U3217 (N_3217,In_1589,In_67);
or U3218 (N_3218,In_149,In_1568);
xnor U3219 (N_3219,In_28,In_24);
and U3220 (N_3220,In_118,In_753);
xor U3221 (N_3221,In_1127,In_1142);
or U3222 (N_3222,In_1706,In_194);
or U3223 (N_3223,In_1904,In_772);
nor U3224 (N_3224,In_1126,In_1217);
and U3225 (N_3225,In_26,In_224);
and U3226 (N_3226,In_829,In_96);
nor U3227 (N_3227,In_523,In_355);
xnor U3228 (N_3228,In_874,In_1520);
and U3229 (N_3229,In_1795,In_1660);
nor U3230 (N_3230,In_310,In_623);
or U3231 (N_3231,In_1713,In_916);
xor U3232 (N_3232,In_1347,In_459);
nor U3233 (N_3233,In_793,In_1216);
xor U3234 (N_3234,In_641,In_1183);
xor U3235 (N_3235,In_1014,In_908);
xnor U3236 (N_3236,In_1839,In_428);
and U3237 (N_3237,In_1522,In_1961);
xor U3238 (N_3238,In_1279,In_1181);
and U3239 (N_3239,In_545,In_1984);
and U3240 (N_3240,In_1295,In_805);
xor U3241 (N_3241,In_1275,In_904);
nand U3242 (N_3242,In_792,In_1118);
nand U3243 (N_3243,In_1652,In_1);
or U3244 (N_3244,In_1932,In_1689);
or U3245 (N_3245,In_638,In_110);
or U3246 (N_3246,In_1003,In_901);
nand U3247 (N_3247,In_1644,In_893);
or U3248 (N_3248,In_975,In_557);
and U3249 (N_3249,In_820,In_1240);
nor U3250 (N_3250,In_1014,In_217);
nor U3251 (N_3251,In_620,In_601);
nor U3252 (N_3252,In_973,In_1225);
and U3253 (N_3253,In_137,In_108);
nor U3254 (N_3254,In_639,In_1180);
nor U3255 (N_3255,In_644,In_680);
or U3256 (N_3256,In_1928,In_884);
or U3257 (N_3257,In_452,In_779);
or U3258 (N_3258,In_750,In_143);
nor U3259 (N_3259,In_986,In_1882);
xor U3260 (N_3260,In_307,In_1116);
or U3261 (N_3261,In_1019,In_1931);
nor U3262 (N_3262,In_407,In_532);
or U3263 (N_3263,In_1761,In_227);
nor U3264 (N_3264,In_176,In_45);
nor U3265 (N_3265,In_1745,In_1526);
xor U3266 (N_3266,In_638,In_1005);
or U3267 (N_3267,In_982,In_1296);
or U3268 (N_3268,In_1545,In_1097);
xor U3269 (N_3269,In_848,In_195);
nor U3270 (N_3270,In_1310,In_1718);
nor U3271 (N_3271,In_1255,In_1160);
nor U3272 (N_3272,In_1556,In_1623);
xor U3273 (N_3273,In_1213,In_1331);
and U3274 (N_3274,In_1958,In_3);
or U3275 (N_3275,In_4,In_534);
and U3276 (N_3276,In_1998,In_1154);
or U3277 (N_3277,In_276,In_452);
nor U3278 (N_3278,In_610,In_902);
nand U3279 (N_3279,In_1113,In_226);
xnor U3280 (N_3280,In_1159,In_1259);
or U3281 (N_3281,In_1845,In_1049);
xnor U3282 (N_3282,In_622,In_1401);
or U3283 (N_3283,In_1587,In_918);
nor U3284 (N_3284,In_1516,In_1401);
and U3285 (N_3285,In_572,In_1188);
nand U3286 (N_3286,In_249,In_1069);
nand U3287 (N_3287,In_1028,In_749);
or U3288 (N_3288,In_1309,In_1995);
nand U3289 (N_3289,In_256,In_1517);
xnor U3290 (N_3290,In_179,In_633);
nor U3291 (N_3291,In_1229,In_1219);
nor U3292 (N_3292,In_1244,In_1586);
or U3293 (N_3293,In_1597,In_1546);
xor U3294 (N_3294,In_1577,In_751);
nand U3295 (N_3295,In_1937,In_1042);
nand U3296 (N_3296,In_361,In_376);
and U3297 (N_3297,In_94,In_697);
nor U3298 (N_3298,In_715,In_1504);
or U3299 (N_3299,In_37,In_1924);
or U3300 (N_3300,In_575,In_392);
or U3301 (N_3301,In_485,In_1439);
or U3302 (N_3302,In_154,In_338);
nand U3303 (N_3303,In_155,In_223);
and U3304 (N_3304,In_1059,In_1663);
or U3305 (N_3305,In_1280,In_735);
and U3306 (N_3306,In_1218,In_893);
xnor U3307 (N_3307,In_236,In_1285);
and U3308 (N_3308,In_279,In_625);
and U3309 (N_3309,In_902,In_407);
xnor U3310 (N_3310,In_801,In_1757);
or U3311 (N_3311,In_1274,In_415);
xnor U3312 (N_3312,In_124,In_1271);
xnor U3313 (N_3313,In_697,In_1161);
xor U3314 (N_3314,In_1460,In_782);
nand U3315 (N_3315,In_428,In_1988);
nand U3316 (N_3316,In_597,In_636);
xor U3317 (N_3317,In_778,In_952);
nand U3318 (N_3318,In_1870,In_1523);
or U3319 (N_3319,In_26,In_543);
nand U3320 (N_3320,In_1094,In_1961);
or U3321 (N_3321,In_1113,In_652);
nor U3322 (N_3322,In_635,In_69);
and U3323 (N_3323,In_1585,In_1345);
nand U3324 (N_3324,In_1411,In_282);
nor U3325 (N_3325,In_197,In_249);
and U3326 (N_3326,In_1016,In_760);
xnor U3327 (N_3327,In_1001,In_81);
and U3328 (N_3328,In_998,In_1076);
nand U3329 (N_3329,In_1348,In_1643);
nand U3330 (N_3330,In_1935,In_803);
nor U3331 (N_3331,In_1646,In_1462);
nor U3332 (N_3332,In_1302,In_1944);
and U3333 (N_3333,In_1178,In_1027);
and U3334 (N_3334,In_857,In_1562);
nand U3335 (N_3335,In_102,In_1528);
and U3336 (N_3336,In_790,In_1763);
and U3337 (N_3337,In_818,In_1565);
nand U3338 (N_3338,In_1249,In_1399);
xnor U3339 (N_3339,In_1615,In_293);
nor U3340 (N_3340,In_251,In_650);
nor U3341 (N_3341,In_600,In_287);
nand U3342 (N_3342,In_1991,In_912);
xnor U3343 (N_3343,In_726,In_1041);
and U3344 (N_3344,In_527,In_846);
xor U3345 (N_3345,In_1619,In_1940);
or U3346 (N_3346,In_874,In_1582);
xnor U3347 (N_3347,In_338,In_60);
xor U3348 (N_3348,In_225,In_78);
nor U3349 (N_3349,In_222,In_104);
xor U3350 (N_3350,In_1135,In_37);
xnor U3351 (N_3351,In_251,In_1150);
and U3352 (N_3352,In_1774,In_952);
nor U3353 (N_3353,In_1402,In_1277);
nand U3354 (N_3354,In_672,In_1978);
nand U3355 (N_3355,In_1899,In_364);
xor U3356 (N_3356,In_474,In_280);
nand U3357 (N_3357,In_1233,In_1584);
or U3358 (N_3358,In_1413,In_1101);
nand U3359 (N_3359,In_791,In_1734);
xnor U3360 (N_3360,In_1440,In_999);
nor U3361 (N_3361,In_1638,In_562);
or U3362 (N_3362,In_1643,In_1749);
nand U3363 (N_3363,In_1225,In_1323);
xnor U3364 (N_3364,In_605,In_1157);
nand U3365 (N_3365,In_1407,In_315);
nor U3366 (N_3366,In_188,In_1168);
xor U3367 (N_3367,In_1907,In_1514);
or U3368 (N_3368,In_1583,In_1274);
nor U3369 (N_3369,In_1087,In_1839);
and U3370 (N_3370,In_1132,In_1129);
nand U3371 (N_3371,In_1830,In_4);
and U3372 (N_3372,In_1125,In_1093);
nor U3373 (N_3373,In_996,In_170);
nor U3374 (N_3374,In_1173,In_1026);
or U3375 (N_3375,In_1903,In_802);
nor U3376 (N_3376,In_493,In_78);
and U3377 (N_3377,In_363,In_66);
xnor U3378 (N_3378,In_708,In_694);
nand U3379 (N_3379,In_190,In_1030);
xor U3380 (N_3380,In_1716,In_148);
and U3381 (N_3381,In_593,In_335);
xor U3382 (N_3382,In_559,In_1631);
xnor U3383 (N_3383,In_800,In_355);
and U3384 (N_3384,In_656,In_1002);
xnor U3385 (N_3385,In_420,In_609);
xor U3386 (N_3386,In_928,In_1103);
nor U3387 (N_3387,In_430,In_397);
nor U3388 (N_3388,In_1809,In_1388);
or U3389 (N_3389,In_217,In_1377);
and U3390 (N_3390,In_1476,In_1863);
nor U3391 (N_3391,In_1510,In_1571);
and U3392 (N_3392,In_174,In_26);
xor U3393 (N_3393,In_497,In_1367);
xnor U3394 (N_3394,In_124,In_1031);
xnor U3395 (N_3395,In_1784,In_81);
xnor U3396 (N_3396,In_152,In_607);
xnor U3397 (N_3397,In_1418,In_1858);
xnor U3398 (N_3398,In_958,In_92);
xor U3399 (N_3399,In_661,In_1968);
xor U3400 (N_3400,In_1414,In_168);
or U3401 (N_3401,In_646,In_1828);
nand U3402 (N_3402,In_1905,In_662);
nand U3403 (N_3403,In_1924,In_1097);
or U3404 (N_3404,In_754,In_966);
nor U3405 (N_3405,In_368,In_117);
nand U3406 (N_3406,In_1827,In_1048);
nand U3407 (N_3407,In_1871,In_1546);
xor U3408 (N_3408,In_1901,In_895);
xnor U3409 (N_3409,In_1482,In_500);
nor U3410 (N_3410,In_1411,In_411);
xnor U3411 (N_3411,In_220,In_1312);
nand U3412 (N_3412,In_1807,In_1934);
and U3413 (N_3413,In_1844,In_1040);
and U3414 (N_3414,In_843,In_1069);
nand U3415 (N_3415,In_869,In_625);
nand U3416 (N_3416,In_1231,In_1045);
and U3417 (N_3417,In_1170,In_86);
xnor U3418 (N_3418,In_104,In_513);
nand U3419 (N_3419,In_1442,In_42);
nor U3420 (N_3420,In_28,In_914);
and U3421 (N_3421,In_1925,In_733);
nor U3422 (N_3422,In_301,In_1437);
nand U3423 (N_3423,In_1684,In_1882);
and U3424 (N_3424,In_1787,In_70);
nor U3425 (N_3425,In_783,In_970);
nor U3426 (N_3426,In_1082,In_461);
xnor U3427 (N_3427,In_1003,In_46);
xor U3428 (N_3428,In_707,In_520);
nand U3429 (N_3429,In_460,In_1928);
or U3430 (N_3430,In_1612,In_541);
nand U3431 (N_3431,In_1159,In_1323);
nor U3432 (N_3432,In_1124,In_822);
nand U3433 (N_3433,In_881,In_1658);
nand U3434 (N_3434,In_927,In_1746);
nand U3435 (N_3435,In_1030,In_449);
and U3436 (N_3436,In_1761,In_229);
or U3437 (N_3437,In_1773,In_1127);
xnor U3438 (N_3438,In_1547,In_1219);
or U3439 (N_3439,In_834,In_1607);
and U3440 (N_3440,In_1826,In_1886);
nand U3441 (N_3441,In_62,In_502);
xor U3442 (N_3442,In_371,In_1195);
nor U3443 (N_3443,In_1397,In_418);
and U3444 (N_3444,In_602,In_1225);
and U3445 (N_3445,In_1997,In_592);
or U3446 (N_3446,In_261,In_417);
nand U3447 (N_3447,In_192,In_863);
or U3448 (N_3448,In_1737,In_1804);
or U3449 (N_3449,In_139,In_532);
nor U3450 (N_3450,In_1349,In_1445);
and U3451 (N_3451,In_1913,In_264);
xnor U3452 (N_3452,In_235,In_7);
and U3453 (N_3453,In_1512,In_468);
nand U3454 (N_3454,In_264,In_1879);
nor U3455 (N_3455,In_652,In_1485);
xnor U3456 (N_3456,In_62,In_981);
and U3457 (N_3457,In_1744,In_1652);
and U3458 (N_3458,In_1143,In_1164);
or U3459 (N_3459,In_1634,In_1319);
xor U3460 (N_3460,In_310,In_909);
xor U3461 (N_3461,In_355,In_1997);
or U3462 (N_3462,In_669,In_957);
and U3463 (N_3463,In_627,In_97);
xor U3464 (N_3464,In_757,In_484);
nor U3465 (N_3465,In_447,In_1681);
nor U3466 (N_3466,In_1240,In_1393);
and U3467 (N_3467,In_216,In_1937);
xor U3468 (N_3468,In_905,In_1873);
and U3469 (N_3469,In_2,In_1761);
and U3470 (N_3470,In_531,In_633);
nand U3471 (N_3471,In_469,In_1880);
and U3472 (N_3472,In_740,In_711);
or U3473 (N_3473,In_1760,In_235);
nand U3474 (N_3474,In_621,In_1854);
or U3475 (N_3475,In_1767,In_61);
nor U3476 (N_3476,In_911,In_1576);
or U3477 (N_3477,In_659,In_1713);
and U3478 (N_3478,In_1260,In_621);
nand U3479 (N_3479,In_1900,In_1144);
nor U3480 (N_3480,In_1430,In_659);
nor U3481 (N_3481,In_1132,In_1674);
and U3482 (N_3482,In_1110,In_237);
nand U3483 (N_3483,In_1972,In_898);
nand U3484 (N_3484,In_1173,In_847);
nand U3485 (N_3485,In_1439,In_1068);
or U3486 (N_3486,In_470,In_1822);
nor U3487 (N_3487,In_747,In_12);
and U3488 (N_3488,In_624,In_566);
and U3489 (N_3489,In_1901,In_1356);
nand U3490 (N_3490,In_1904,In_391);
or U3491 (N_3491,In_1751,In_966);
or U3492 (N_3492,In_1571,In_726);
or U3493 (N_3493,In_1030,In_1979);
nor U3494 (N_3494,In_751,In_433);
xnor U3495 (N_3495,In_108,In_1252);
nor U3496 (N_3496,In_1169,In_1943);
and U3497 (N_3497,In_1160,In_1614);
nand U3498 (N_3498,In_1989,In_949);
nor U3499 (N_3499,In_1704,In_1930);
and U3500 (N_3500,In_587,In_1263);
and U3501 (N_3501,In_480,In_297);
nor U3502 (N_3502,In_1043,In_356);
xnor U3503 (N_3503,In_607,In_224);
and U3504 (N_3504,In_1979,In_334);
or U3505 (N_3505,In_1711,In_1555);
nand U3506 (N_3506,In_541,In_1422);
xor U3507 (N_3507,In_1866,In_906);
nor U3508 (N_3508,In_1067,In_797);
nor U3509 (N_3509,In_635,In_608);
and U3510 (N_3510,In_578,In_196);
nor U3511 (N_3511,In_482,In_1754);
nand U3512 (N_3512,In_526,In_563);
or U3513 (N_3513,In_1888,In_1605);
or U3514 (N_3514,In_770,In_1479);
xnor U3515 (N_3515,In_1935,In_277);
or U3516 (N_3516,In_1289,In_1187);
and U3517 (N_3517,In_1242,In_1886);
nor U3518 (N_3518,In_30,In_332);
nand U3519 (N_3519,In_909,In_230);
and U3520 (N_3520,In_1466,In_1753);
nand U3521 (N_3521,In_579,In_913);
nand U3522 (N_3522,In_925,In_357);
and U3523 (N_3523,In_1713,In_263);
or U3524 (N_3524,In_791,In_798);
xnor U3525 (N_3525,In_267,In_345);
or U3526 (N_3526,In_1255,In_370);
nand U3527 (N_3527,In_1792,In_1002);
xor U3528 (N_3528,In_1547,In_777);
and U3529 (N_3529,In_302,In_888);
nor U3530 (N_3530,In_645,In_1840);
nand U3531 (N_3531,In_1173,In_1120);
and U3532 (N_3532,In_1828,In_1326);
xor U3533 (N_3533,In_1441,In_389);
nor U3534 (N_3534,In_309,In_1395);
nor U3535 (N_3535,In_1844,In_1294);
xor U3536 (N_3536,In_19,In_129);
xor U3537 (N_3537,In_1984,In_1851);
and U3538 (N_3538,In_846,In_160);
or U3539 (N_3539,In_411,In_599);
and U3540 (N_3540,In_316,In_209);
nand U3541 (N_3541,In_627,In_1792);
xnor U3542 (N_3542,In_956,In_1183);
xor U3543 (N_3543,In_713,In_1419);
nor U3544 (N_3544,In_343,In_425);
nand U3545 (N_3545,In_1077,In_1671);
nand U3546 (N_3546,In_663,In_1449);
and U3547 (N_3547,In_672,In_869);
nor U3548 (N_3548,In_848,In_472);
nand U3549 (N_3549,In_398,In_466);
or U3550 (N_3550,In_1700,In_951);
xor U3551 (N_3551,In_339,In_613);
nor U3552 (N_3552,In_396,In_381);
nor U3553 (N_3553,In_1172,In_508);
and U3554 (N_3554,In_792,In_92);
or U3555 (N_3555,In_449,In_491);
or U3556 (N_3556,In_77,In_970);
nor U3557 (N_3557,In_565,In_1113);
nand U3558 (N_3558,In_1867,In_639);
or U3559 (N_3559,In_1983,In_1835);
nand U3560 (N_3560,In_29,In_394);
xnor U3561 (N_3561,In_1188,In_1127);
or U3562 (N_3562,In_1713,In_67);
nand U3563 (N_3563,In_291,In_1394);
xor U3564 (N_3564,In_530,In_1947);
and U3565 (N_3565,In_832,In_192);
nand U3566 (N_3566,In_1212,In_701);
xor U3567 (N_3567,In_743,In_876);
nand U3568 (N_3568,In_1094,In_1262);
or U3569 (N_3569,In_1393,In_44);
xor U3570 (N_3570,In_1541,In_1339);
xnor U3571 (N_3571,In_1426,In_854);
nand U3572 (N_3572,In_1422,In_1884);
nand U3573 (N_3573,In_2,In_1524);
and U3574 (N_3574,In_922,In_1053);
and U3575 (N_3575,In_1760,In_1827);
nor U3576 (N_3576,In_1725,In_1732);
xor U3577 (N_3577,In_1492,In_386);
xnor U3578 (N_3578,In_1914,In_951);
nand U3579 (N_3579,In_960,In_558);
nor U3580 (N_3580,In_545,In_787);
or U3581 (N_3581,In_135,In_1623);
nand U3582 (N_3582,In_1284,In_1259);
nor U3583 (N_3583,In_1913,In_788);
nand U3584 (N_3584,In_987,In_883);
or U3585 (N_3585,In_1588,In_1160);
nor U3586 (N_3586,In_284,In_1631);
nor U3587 (N_3587,In_1683,In_1165);
xnor U3588 (N_3588,In_768,In_1095);
or U3589 (N_3589,In_9,In_1611);
nor U3590 (N_3590,In_551,In_830);
xnor U3591 (N_3591,In_55,In_1850);
nand U3592 (N_3592,In_797,In_1509);
nor U3593 (N_3593,In_723,In_377);
xor U3594 (N_3594,In_1985,In_1038);
xor U3595 (N_3595,In_1161,In_93);
nor U3596 (N_3596,In_1610,In_903);
and U3597 (N_3597,In_1005,In_1642);
nand U3598 (N_3598,In_678,In_1941);
xor U3599 (N_3599,In_501,In_1641);
nand U3600 (N_3600,In_938,In_934);
nor U3601 (N_3601,In_170,In_12);
nor U3602 (N_3602,In_1413,In_298);
xnor U3603 (N_3603,In_103,In_1875);
xnor U3604 (N_3604,In_1597,In_1848);
nor U3605 (N_3605,In_1580,In_1906);
nand U3606 (N_3606,In_1080,In_1508);
xnor U3607 (N_3607,In_543,In_1293);
nor U3608 (N_3608,In_1924,In_1623);
or U3609 (N_3609,In_970,In_1197);
xor U3610 (N_3610,In_240,In_768);
and U3611 (N_3611,In_1776,In_321);
nand U3612 (N_3612,In_220,In_1191);
nand U3613 (N_3613,In_1450,In_918);
and U3614 (N_3614,In_653,In_1394);
xnor U3615 (N_3615,In_1646,In_1019);
or U3616 (N_3616,In_434,In_1730);
xnor U3617 (N_3617,In_1878,In_1363);
or U3618 (N_3618,In_504,In_1513);
nor U3619 (N_3619,In_888,In_392);
nand U3620 (N_3620,In_930,In_832);
xor U3621 (N_3621,In_1101,In_654);
nor U3622 (N_3622,In_1221,In_1890);
nand U3623 (N_3623,In_860,In_1546);
xnor U3624 (N_3624,In_1592,In_1467);
xor U3625 (N_3625,In_187,In_1942);
or U3626 (N_3626,In_1481,In_1558);
nor U3627 (N_3627,In_684,In_169);
and U3628 (N_3628,In_1943,In_1065);
nor U3629 (N_3629,In_1744,In_1252);
xor U3630 (N_3630,In_1072,In_455);
nor U3631 (N_3631,In_1140,In_1845);
and U3632 (N_3632,In_1017,In_795);
nand U3633 (N_3633,In_1879,In_629);
or U3634 (N_3634,In_1844,In_1733);
xnor U3635 (N_3635,In_1981,In_454);
nand U3636 (N_3636,In_668,In_672);
and U3637 (N_3637,In_278,In_1345);
nand U3638 (N_3638,In_965,In_132);
xnor U3639 (N_3639,In_805,In_1374);
xor U3640 (N_3640,In_258,In_1911);
and U3641 (N_3641,In_1113,In_1573);
nand U3642 (N_3642,In_1302,In_975);
nand U3643 (N_3643,In_1630,In_812);
or U3644 (N_3644,In_197,In_1993);
nor U3645 (N_3645,In_1334,In_773);
and U3646 (N_3646,In_1253,In_1179);
nor U3647 (N_3647,In_1795,In_115);
xor U3648 (N_3648,In_1236,In_804);
nand U3649 (N_3649,In_840,In_1482);
xor U3650 (N_3650,In_669,In_528);
xor U3651 (N_3651,In_1834,In_854);
xor U3652 (N_3652,In_1551,In_1872);
nor U3653 (N_3653,In_213,In_1636);
nand U3654 (N_3654,In_584,In_1567);
and U3655 (N_3655,In_224,In_1125);
nor U3656 (N_3656,In_1869,In_271);
xor U3657 (N_3657,In_1331,In_372);
and U3658 (N_3658,In_161,In_1351);
nand U3659 (N_3659,In_769,In_1454);
or U3660 (N_3660,In_794,In_1916);
nor U3661 (N_3661,In_536,In_25);
and U3662 (N_3662,In_190,In_1785);
nor U3663 (N_3663,In_270,In_982);
nor U3664 (N_3664,In_1058,In_1746);
or U3665 (N_3665,In_1458,In_1876);
nor U3666 (N_3666,In_172,In_995);
xor U3667 (N_3667,In_553,In_8);
or U3668 (N_3668,In_656,In_1350);
nand U3669 (N_3669,In_1073,In_1399);
or U3670 (N_3670,In_766,In_1895);
xnor U3671 (N_3671,In_1896,In_386);
nor U3672 (N_3672,In_222,In_96);
nor U3673 (N_3673,In_1797,In_1815);
or U3674 (N_3674,In_1573,In_1145);
or U3675 (N_3675,In_1798,In_334);
and U3676 (N_3676,In_1984,In_868);
xnor U3677 (N_3677,In_1699,In_642);
nand U3678 (N_3678,In_1486,In_1438);
nand U3679 (N_3679,In_346,In_333);
xor U3680 (N_3680,In_6,In_1648);
xor U3681 (N_3681,In_73,In_1633);
or U3682 (N_3682,In_1868,In_465);
xor U3683 (N_3683,In_591,In_1618);
xnor U3684 (N_3684,In_540,In_1853);
and U3685 (N_3685,In_1132,In_1465);
nor U3686 (N_3686,In_454,In_816);
nor U3687 (N_3687,In_833,In_208);
nor U3688 (N_3688,In_757,In_915);
nand U3689 (N_3689,In_608,In_813);
and U3690 (N_3690,In_955,In_723);
xor U3691 (N_3691,In_1501,In_281);
nand U3692 (N_3692,In_923,In_236);
nor U3693 (N_3693,In_605,In_1727);
nand U3694 (N_3694,In_280,In_999);
or U3695 (N_3695,In_423,In_827);
and U3696 (N_3696,In_141,In_396);
nor U3697 (N_3697,In_446,In_622);
xor U3698 (N_3698,In_61,In_443);
xnor U3699 (N_3699,In_42,In_1905);
and U3700 (N_3700,In_1770,In_78);
xor U3701 (N_3701,In_1784,In_1930);
and U3702 (N_3702,In_16,In_192);
xor U3703 (N_3703,In_209,In_284);
xor U3704 (N_3704,In_507,In_300);
xor U3705 (N_3705,In_1236,In_1672);
and U3706 (N_3706,In_1445,In_1908);
nand U3707 (N_3707,In_1996,In_662);
xnor U3708 (N_3708,In_777,In_1956);
or U3709 (N_3709,In_117,In_1091);
or U3710 (N_3710,In_1469,In_97);
nor U3711 (N_3711,In_190,In_421);
and U3712 (N_3712,In_81,In_1460);
xnor U3713 (N_3713,In_187,In_1580);
or U3714 (N_3714,In_35,In_1459);
nand U3715 (N_3715,In_55,In_630);
or U3716 (N_3716,In_685,In_419);
xnor U3717 (N_3717,In_1079,In_100);
and U3718 (N_3718,In_1836,In_82);
nand U3719 (N_3719,In_1512,In_22);
nor U3720 (N_3720,In_974,In_1281);
nand U3721 (N_3721,In_1804,In_436);
or U3722 (N_3722,In_719,In_801);
and U3723 (N_3723,In_150,In_644);
xnor U3724 (N_3724,In_1101,In_548);
xor U3725 (N_3725,In_1930,In_1065);
xor U3726 (N_3726,In_1968,In_1265);
nor U3727 (N_3727,In_434,In_1827);
or U3728 (N_3728,In_1792,In_677);
and U3729 (N_3729,In_1711,In_88);
nor U3730 (N_3730,In_498,In_1111);
and U3731 (N_3731,In_674,In_1355);
or U3732 (N_3732,In_1090,In_1725);
nor U3733 (N_3733,In_1036,In_1354);
nor U3734 (N_3734,In_1739,In_1417);
nor U3735 (N_3735,In_538,In_1978);
or U3736 (N_3736,In_1810,In_1469);
xnor U3737 (N_3737,In_771,In_587);
nor U3738 (N_3738,In_281,In_1664);
nand U3739 (N_3739,In_1240,In_1259);
nand U3740 (N_3740,In_1724,In_262);
and U3741 (N_3741,In_862,In_724);
and U3742 (N_3742,In_93,In_1323);
xor U3743 (N_3743,In_902,In_1724);
nor U3744 (N_3744,In_1086,In_183);
and U3745 (N_3745,In_668,In_957);
xnor U3746 (N_3746,In_1678,In_75);
or U3747 (N_3747,In_401,In_1170);
xor U3748 (N_3748,In_664,In_1340);
and U3749 (N_3749,In_1964,In_1758);
and U3750 (N_3750,In_949,In_1234);
and U3751 (N_3751,In_899,In_100);
xor U3752 (N_3752,In_115,In_515);
nand U3753 (N_3753,In_762,In_1916);
nand U3754 (N_3754,In_1934,In_1160);
nand U3755 (N_3755,In_1784,In_510);
nand U3756 (N_3756,In_735,In_581);
nor U3757 (N_3757,In_149,In_914);
or U3758 (N_3758,In_1360,In_1398);
nand U3759 (N_3759,In_1367,In_967);
and U3760 (N_3760,In_48,In_566);
nand U3761 (N_3761,In_254,In_407);
nand U3762 (N_3762,In_729,In_553);
and U3763 (N_3763,In_1790,In_632);
nand U3764 (N_3764,In_231,In_770);
and U3765 (N_3765,In_1657,In_1999);
xnor U3766 (N_3766,In_521,In_1356);
xnor U3767 (N_3767,In_1821,In_1798);
nor U3768 (N_3768,In_1116,In_690);
xor U3769 (N_3769,In_1674,In_1291);
xor U3770 (N_3770,In_203,In_1982);
nand U3771 (N_3771,In_335,In_81);
xnor U3772 (N_3772,In_407,In_815);
xor U3773 (N_3773,In_560,In_1229);
nor U3774 (N_3774,In_1206,In_1633);
or U3775 (N_3775,In_924,In_1257);
nor U3776 (N_3776,In_1614,In_125);
nor U3777 (N_3777,In_1032,In_1508);
nand U3778 (N_3778,In_1372,In_308);
nand U3779 (N_3779,In_1912,In_332);
or U3780 (N_3780,In_677,In_1270);
or U3781 (N_3781,In_709,In_1472);
and U3782 (N_3782,In_1672,In_46);
nand U3783 (N_3783,In_713,In_1376);
or U3784 (N_3784,In_1924,In_1318);
nand U3785 (N_3785,In_12,In_1511);
nor U3786 (N_3786,In_86,In_862);
nor U3787 (N_3787,In_873,In_1721);
or U3788 (N_3788,In_1798,In_762);
nand U3789 (N_3789,In_1198,In_1602);
nor U3790 (N_3790,In_1771,In_608);
and U3791 (N_3791,In_1999,In_1384);
xor U3792 (N_3792,In_1256,In_1898);
and U3793 (N_3793,In_1551,In_22);
nand U3794 (N_3794,In_137,In_1466);
nor U3795 (N_3795,In_1254,In_618);
nor U3796 (N_3796,In_1334,In_437);
nand U3797 (N_3797,In_60,In_1445);
or U3798 (N_3798,In_1288,In_772);
nand U3799 (N_3799,In_1263,In_173);
nand U3800 (N_3800,In_1988,In_677);
or U3801 (N_3801,In_373,In_1293);
or U3802 (N_3802,In_306,In_1513);
xor U3803 (N_3803,In_1529,In_1203);
nand U3804 (N_3804,In_1545,In_1912);
nand U3805 (N_3805,In_1833,In_1752);
nand U3806 (N_3806,In_555,In_1672);
nor U3807 (N_3807,In_322,In_566);
xor U3808 (N_3808,In_912,In_1170);
xnor U3809 (N_3809,In_711,In_535);
and U3810 (N_3810,In_227,In_583);
xnor U3811 (N_3811,In_1016,In_1898);
and U3812 (N_3812,In_1280,In_156);
and U3813 (N_3813,In_1540,In_203);
or U3814 (N_3814,In_1859,In_200);
and U3815 (N_3815,In_1296,In_101);
or U3816 (N_3816,In_1837,In_1052);
or U3817 (N_3817,In_730,In_23);
nand U3818 (N_3818,In_778,In_1695);
nand U3819 (N_3819,In_465,In_474);
and U3820 (N_3820,In_1214,In_353);
or U3821 (N_3821,In_1315,In_1096);
nor U3822 (N_3822,In_1751,In_1375);
xnor U3823 (N_3823,In_504,In_1143);
xnor U3824 (N_3824,In_213,In_287);
or U3825 (N_3825,In_965,In_1706);
nor U3826 (N_3826,In_925,In_1243);
and U3827 (N_3827,In_1399,In_134);
or U3828 (N_3828,In_120,In_1393);
and U3829 (N_3829,In_1107,In_1149);
nand U3830 (N_3830,In_1249,In_1866);
or U3831 (N_3831,In_78,In_30);
and U3832 (N_3832,In_1354,In_1555);
xnor U3833 (N_3833,In_1218,In_588);
and U3834 (N_3834,In_1426,In_795);
nand U3835 (N_3835,In_1859,In_1777);
xnor U3836 (N_3836,In_1247,In_253);
and U3837 (N_3837,In_1683,In_56);
nor U3838 (N_3838,In_1916,In_149);
or U3839 (N_3839,In_1979,In_1968);
xor U3840 (N_3840,In_1421,In_1819);
xnor U3841 (N_3841,In_1795,In_1103);
nor U3842 (N_3842,In_1295,In_733);
xor U3843 (N_3843,In_246,In_1860);
and U3844 (N_3844,In_511,In_1278);
xnor U3845 (N_3845,In_1928,In_259);
xnor U3846 (N_3846,In_1172,In_95);
or U3847 (N_3847,In_39,In_540);
or U3848 (N_3848,In_1582,In_1089);
and U3849 (N_3849,In_1718,In_1696);
or U3850 (N_3850,In_432,In_1120);
xor U3851 (N_3851,In_958,In_1705);
nand U3852 (N_3852,In_1978,In_940);
or U3853 (N_3853,In_90,In_1401);
and U3854 (N_3854,In_844,In_1144);
xnor U3855 (N_3855,In_226,In_668);
nand U3856 (N_3856,In_412,In_727);
nor U3857 (N_3857,In_441,In_1825);
and U3858 (N_3858,In_970,In_857);
or U3859 (N_3859,In_975,In_916);
xnor U3860 (N_3860,In_142,In_1620);
nor U3861 (N_3861,In_254,In_775);
and U3862 (N_3862,In_6,In_573);
or U3863 (N_3863,In_528,In_1101);
nand U3864 (N_3864,In_1719,In_1500);
and U3865 (N_3865,In_1530,In_987);
and U3866 (N_3866,In_964,In_1451);
nand U3867 (N_3867,In_1402,In_1451);
and U3868 (N_3868,In_1750,In_26);
xor U3869 (N_3869,In_285,In_1629);
nor U3870 (N_3870,In_985,In_1174);
xor U3871 (N_3871,In_1589,In_209);
or U3872 (N_3872,In_1022,In_505);
nor U3873 (N_3873,In_1743,In_223);
xor U3874 (N_3874,In_1493,In_1398);
nor U3875 (N_3875,In_659,In_550);
xnor U3876 (N_3876,In_474,In_1505);
nand U3877 (N_3877,In_1232,In_555);
xnor U3878 (N_3878,In_1150,In_1204);
or U3879 (N_3879,In_100,In_734);
nand U3880 (N_3880,In_1836,In_1718);
xor U3881 (N_3881,In_516,In_240);
or U3882 (N_3882,In_42,In_816);
or U3883 (N_3883,In_799,In_1344);
nand U3884 (N_3884,In_1840,In_538);
or U3885 (N_3885,In_1648,In_775);
nor U3886 (N_3886,In_998,In_351);
xnor U3887 (N_3887,In_155,In_1750);
nor U3888 (N_3888,In_788,In_1828);
nand U3889 (N_3889,In_170,In_1646);
nand U3890 (N_3890,In_118,In_1540);
or U3891 (N_3891,In_291,In_1058);
xnor U3892 (N_3892,In_1864,In_286);
xor U3893 (N_3893,In_1275,In_1912);
nor U3894 (N_3894,In_716,In_241);
xor U3895 (N_3895,In_545,In_346);
nand U3896 (N_3896,In_1377,In_340);
nand U3897 (N_3897,In_1899,In_896);
or U3898 (N_3898,In_825,In_1577);
xor U3899 (N_3899,In_670,In_52);
xor U3900 (N_3900,In_331,In_455);
and U3901 (N_3901,In_1573,In_1852);
or U3902 (N_3902,In_1479,In_160);
and U3903 (N_3903,In_846,In_1902);
and U3904 (N_3904,In_854,In_1008);
and U3905 (N_3905,In_1319,In_756);
and U3906 (N_3906,In_958,In_1517);
nand U3907 (N_3907,In_1231,In_51);
or U3908 (N_3908,In_850,In_1717);
or U3909 (N_3909,In_60,In_433);
nor U3910 (N_3910,In_1833,In_1315);
nand U3911 (N_3911,In_59,In_803);
nand U3912 (N_3912,In_1259,In_141);
and U3913 (N_3913,In_328,In_1579);
xor U3914 (N_3914,In_1721,In_810);
or U3915 (N_3915,In_1019,In_1398);
and U3916 (N_3916,In_637,In_1394);
nor U3917 (N_3917,In_299,In_1772);
and U3918 (N_3918,In_597,In_1194);
or U3919 (N_3919,In_496,In_30);
or U3920 (N_3920,In_1643,In_1780);
xor U3921 (N_3921,In_629,In_1764);
xor U3922 (N_3922,In_1599,In_1612);
or U3923 (N_3923,In_1661,In_1108);
or U3924 (N_3924,In_1272,In_541);
nand U3925 (N_3925,In_536,In_929);
nand U3926 (N_3926,In_1572,In_823);
nor U3927 (N_3927,In_896,In_996);
nand U3928 (N_3928,In_123,In_317);
and U3929 (N_3929,In_438,In_220);
xor U3930 (N_3930,In_1755,In_1780);
nor U3931 (N_3931,In_1393,In_1144);
nor U3932 (N_3932,In_1736,In_340);
xnor U3933 (N_3933,In_428,In_1381);
xnor U3934 (N_3934,In_1286,In_1889);
nor U3935 (N_3935,In_1553,In_828);
nor U3936 (N_3936,In_134,In_140);
nor U3937 (N_3937,In_1603,In_203);
and U3938 (N_3938,In_1539,In_929);
nor U3939 (N_3939,In_320,In_1029);
and U3940 (N_3940,In_245,In_1611);
or U3941 (N_3941,In_245,In_1894);
and U3942 (N_3942,In_570,In_1942);
xor U3943 (N_3943,In_1711,In_597);
xnor U3944 (N_3944,In_660,In_200);
nand U3945 (N_3945,In_1195,In_1692);
nor U3946 (N_3946,In_1089,In_930);
nor U3947 (N_3947,In_123,In_1481);
or U3948 (N_3948,In_1299,In_425);
xnor U3949 (N_3949,In_390,In_357);
and U3950 (N_3950,In_1296,In_58);
nor U3951 (N_3951,In_1812,In_24);
and U3952 (N_3952,In_1293,In_1381);
and U3953 (N_3953,In_1162,In_714);
or U3954 (N_3954,In_1978,In_1258);
nand U3955 (N_3955,In_843,In_1085);
and U3956 (N_3956,In_762,In_567);
or U3957 (N_3957,In_118,In_8);
nand U3958 (N_3958,In_1544,In_767);
nor U3959 (N_3959,In_804,In_1092);
nand U3960 (N_3960,In_211,In_1321);
nor U3961 (N_3961,In_746,In_1405);
and U3962 (N_3962,In_1252,In_1630);
xnor U3963 (N_3963,In_923,In_552);
nand U3964 (N_3964,In_1297,In_69);
and U3965 (N_3965,In_41,In_1471);
and U3966 (N_3966,In_155,In_1961);
nor U3967 (N_3967,In_539,In_1846);
nor U3968 (N_3968,In_1713,In_357);
or U3969 (N_3969,In_658,In_1026);
or U3970 (N_3970,In_321,In_1855);
and U3971 (N_3971,In_1661,In_1399);
and U3972 (N_3972,In_1924,In_1606);
and U3973 (N_3973,In_19,In_1246);
xnor U3974 (N_3974,In_1054,In_248);
nor U3975 (N_3975,In_347,In_108);
nor U3976 (N_3976,In_404,In_963);
nand U3977 (N_3977,In_1859,In_933);
or U3978 (N_3978,In_732,In_425);
nand U3979 (N_3979,In_698,In_1618);
and U3980 (N_3980,In_1885,In_1149);
xnor U3981 (N_3981,In_750,In_327);
xor U3982 (N_3982,In_1697,In_967);
or U3983 (N_3983,In_651,In_1603);
nor U3984 (N_3984,In_709,In_629);
and U3985 (N_3985,In_403,In_937);
and U3986 (N_3986,In_334,In_465);
or U3987 (N_3987,In_93,In_160);
xnor U3988 (N_3988,In_378,In_161);
xor U3989 (N_3989,In_1900,In_391);
nor U3990 (N_3990,In_1733,In_1719);
nand U3991 (N_3991,In_1372,In_53);
nor U3992 (N_3992,In_1511,In_1630);
nand U3993 (N_3993,In_1636,In_1448);
nor U3994 (N_3994,In_618,In_1958);
xor U3995 (N_3995,In_1793,In_1341);
nor U3996 (N_3996,In_1437,In_331);
nor U3997 (N_3997,In_1361,In_976);
and U3998 (N_3998,In_490,In_954);
nand U3999 (N_3999,In_1006,In_1127);
nand U4000 (N_4000,In_1286,In_91);
and U4001 (N_4001,In_381,In_810);
xnor U4002 (N_4002,In_1871,In_709);
or U4003 (N_4003,In_997,In_940);
nor U4004 (N_4004,In_1431,In_1803);
or U4005 (N_4005,In_77,In_1771);
nor U4006 (N_4006,In_338,In_243);
and U4007 (N_4007,In_916,In_1708);
xor U4008 (N_4008,In_382,In_1787);
or U4009 (N_4009,In_487,In_1435);
nor U4010 (N_4010,In_1786,In_322);
xor U4011 (N_4011,In_1752,In_1401);
xnor U4012 (N_4012,In_1023,In_1715);
nand U4013 (N_4013,In_1726,In_1865);
nor U4014 (N_4014,In_4,In_942);
or U4015 (N_4015,In_1171,In_1238);
nor U4016 (N_4016,In_1270,In_535);
nand U4017 (N_4017,In_878,In_1937);
nor U4018 (N_4018,In_1011,In_1102);
nor U4019 (N_4019,In_1306,In_833);
and U4020 (N_4020,In_376,In_1617);
or U4021 (N_4021,In_653,In_1306);
and U4022 (N_4022,In_1448,In_19);
xnor U4023 (N_4023,In_136,In_1429);
and U4024 (N_4024,In_934,In_1387);
nand U4025 (N_4025,In_1666,In_540);
nor U4026 (N_4026,In_550,In_1174);
nand U4027 (N_4027,In_270,In_911);
and U4028 (N_4028,In_1387,In_242);
and U4029 (N_4029,In_617,In_981);
or U4030 (N_4030,In_1537,In_1041);
xor U4031 (N_4031,In_1884,In_490);
and U4032 (N_4032,In_554,In_1856);
and U4033 (N_4033,In_1699,In_1086);
nor U4034 (N_4034,In_812,In_1899);
and U4035 (N_4035,In_1496,In_1923);
or U4036 (N_4036,In_1344,In_681);
and U4037 (N_4037,In_1912,In_1794);
xor U4038 (N_4038,In_838,In_1611);
and U4039 (N_4039,In_1241,In_61);
xor U4040 (N_4040,In_1970,In_18);
or U4041 (N_4041,In_834,In_1057);
or U4042 (N_4042,In_911,In_1653);
or U4043 (N_4043,In_1378,In_1988);
nor U4044 (N_4044,In_1682,In_804);
nor U4045 (N_4045,In_1531,In_533);
or U4046 (N_4046,In_717,In_499);
or U4047 (N_4047,In_1855,In_810);
nand U4048 (N_4048,In_402,In_1451);
xnor U4049 (N_4049,In_1081,In_980);
nor U4050 (N_4050,In_112,In_583);
and U4051 (N_4051,In_449,In_917);
and U4052 (N_4052,In_995,In_1903);
nor U4053 (N_4053,In_887,In_388);
or U4054 (N_4054,In_808,In_730);
or U4055 (N_4055,In_1721,In_1494);
xor U4056 (N_4056,In_43,In_1204);
and U4057 (N_4057,In_85,In_722);
nor U4058 (N_4058,In_35,In_753);
and U4059 (N_4059,In_272,In_42);
and U4060 (N_4060,In_1252,In_872);
and U4061 (N_4061,In_917,In_1095);
nand U4062 (N_4062,In_1580,In_633);
or U4063 (N_4063,In_803,In_1805);
or U4064 (N_4064,In_511,In_1571);
or U4065 (N_4065,In_1057,In_764);
or U4066 (N_4066,In_1956,In_556);
nand U4067 (N_4067,In_1075,In_1684);
nor U4068 (N_4068,In_1940,In_156);
or U4069 (N_4069,In_1778,In_53);
nand U4070 (N_4070,In_871,In_246);
nand U4071 (N_4071,In_989,In_745);
nor U4072 (N_4072,In_585,In_1029);
nor U4073 (N_4073,In_423,In_1099);
nor U4074 (N_4074,In_1414,In_1966);
nor U4075 (N_4075,In_115,In_835);
or U4076 (N_4076,In_318,In_1132);
xnor U4077 (N_4077,In_1874,In_1656);
and U4078 (N_4078,In_641,In_1075);
or U4079 (N_4079,In_286,In_1919);
or U4080 (N_4080,In_1527,In_408);
nand U4081 (N_4081,In_604,In_999);
nand U4082 (N_4082,In_1001,In_1480);
or U4083 (N_4083,In_1892,In_948);
nand U4084 (N_4084,In_304,In_683);
and U4085 (N_4085,In_1664,In_1871);
and U4086 (N_4086,In_544,In_1357);
nor U4087 (N_4087,In_1096,In_664);
or U4088 (N_4088,In_733,In_1600);
and U4089 (N_4089,In_1014,In_1749);
nand U4090 (N_4090,In_126,In_395);
or U4091 (N_4091,In_672,In_777);
and U4092 (N_4092,In_1322,In_419);
nor U4093 (N_4093,In_1708,In_627);
nand U4094 (N_4094,In_216,In_1365);
nand U4095 (N_4095,In_969,In_1519);
nor U4096 (N_4096,In_847,In_331);
nand U4097 (N_4097,In_601,In_929);
and U4098 (N_4098,In_202,In_1789);
and U4099 (N_4099,In_1733,In_415);
or U4100 (N_4100,In_572,In_1720);
and U4101 (N_4101,In_223,In_1875);
xnor U4102 (N_4102,In_690,In_1630);
nand U4103 (N_4103,In_1863,In_1159);
nand U4104 (N_4104,In_1242,In_1266);
nor U4105 (N_4105,In_1664,In_230);
nor U4106 (N_4106,In_1574,In_105);
and U4107 (N_4107,In_22,In_1621);
xor U4108 (N_4108,In_820,In_1379);
xor U4109 (N_4109,In_375,In_1195);
xnor U4110 (N_4110,In_186,In_1655);
or U4111 (N_4111,In_1413,In_1587);
xnor U4112 (N_4112,In_886,In_810);
or U4113 (N_4113,In_1421,In_1452);
and U4114 (N_4114,In_526,In_919);
xnor U4115 (N_4115,In_4,In_558);
or U4116 (N_4116,In_1988,In_553);
and U4117 (N_4117,In_214,In_443);
nor U4118 (N_4118,In_1226,In_802);
xor U4119 (N_4119,In_704,In_1318);
nand U4120 (N_4120,In_958,In_1666);
nor U4121 (N_4121,In_1198,In_538);
and U4122 (N_4122,In_169,In_1297);
or U4123 (N_4123,In_1472,In_1647);
nor U4124 (N_4124,In_1891,In_1231);
xnor U4125 (N_4125,In_1276,In_1896);
nor U4126 (N_4126,In_1849,In_520);
and U4127 (N_4127,In_1271,In_53);
and U4128 (N_4128,In_87,In_664);
nand U4129 (N_4129,In_1032,In_1390);
nor U4130 (N_4130,In_856,In_1427);
xor U4131 (N_4131,In_881,In_1289);
xor U4132 (N_4132,In_636,In_1585);
or U4133 (N_4133,In_1551,In_974);
xor U4134 (N_4134,In_1882,In_1252);
nand U4135 (N_4135,In_682,In_1513);
nand U4136 (N_4136,In_645,In_76);
or U4137 (N_4137,In_325,In_877);
nor U4138 (N_4138,In_1508,In_1386);
nor U4139 (N_4139,In_868,In_1435);
or U4140 (N_4140,In_486,In_1762);
xor U4141 (N_4141,In_766,In_613);
or U4142 (N_4142,In_401,In_1030);
and U4143 (N_4143,In_844,In_148);
xor U4144 (N_4144,In_1800,In_1811);
xnor U4145 (N_4145,In_414,In_1551);
or U4146 (N_4146,In_1831,In_1785);
xor U4147 (N_4147,In_218,In_1436);
xnor U4148 (N_4148,In_1079,In_1305);
and U4149 (N_4149,In_824,In_1655);
nor U4150 (N_4150,In_781,In_720);
and U4151 (N_4151,In_1568,In_1799);
xor U4152 (N_4152,In_562,In_722);
or U4153 (N_4153,In_447,In_214);
nand U4154 (N_4154,In_525,In_484);
and U4155 (N_4155,In_1353,In_1114);
nand U4156 (N_4156,In_1939,In_1834);
and U4157 (N_4157,In_921,In_1570);
nand U4158 (N_4158,In_1426,In_1470);
nand U4159 (N_4159,In_1431,In_1358);
nor U4160 (N_4160,In_1947,In_1812);
or U4161 (N_4161,In_871,In_266);
nand U4162 (N_4162,In_332,In_193);
nand U4163 (N_4163,In_1188,In_182);
and U4164 (N_4164,In_1414,In_1200);
xor U4165 (N_4165,In_530,In_335);
and U4166 (N_4166,In_1212,In_623);
nand U4167 (N_4167,In_72,In_1461);
or U4168 (N_4168,In_560,In_345);
nand U4169 (N_4169,In_561,In_1387);
or U4170 (N_4170,In_558,In_1087);
xnor U4171 (N_4171,In_1533,In_1208);
and U4172 (N_4172,In_232,In_1915);
nand U4173 (N_4173,In_1621,In_1901);
nand U4174 (N_4174,In_967,In_414);
xnor U4175 (N_4175,In_1388,In_1889);
nor U4176 (N_4176,In_560,In_415);
nor U4177 (N_4177,In_134,In_1261);
nor U4178 (N_4178,In_174,In_1228);
nand U4179 (N_4179,In_1573,In_1797);
xnor U4180 (N_4180,In_1196,In_1824);
and U4181 (N_4181,In_1727,In_76);
or U4182 (N_4182,In_1870,In_1098);
nor U4183 (N_4183,In_1148,In_294);
or U4184 (N_4184,In_1733,In_1756);
and U4185 (N_4185,In_758,In_569);
nand U4186 (N_4186,In_1626,In_695);
nand U4187 (N_4187,In_1220,In_587);
xnor U4188 (N_4188,In_323,In_1457);
nor U4189 (N_4189,In_1111,In_531);
nand U4190 (N_4190,In_1415,In_1362);
nor U4191 (N_4191,In_380,In_1533);
nand U4192 (N_4192,In_1167,In_827);
xor U4193 (N_4193,In_549,In_1179);
nor U4194 (N_4194,In_51,In_188);
nand U4195 (N_4195,In_1673,In_1694);
xor U4196 (N_4196,In_1970,In_246);
xnor U4197 (N_4197,In_1526,In_500);
xnor U4198 (N_4198,In_836,In_1103);
nand U4199 (N_4199,In_1734,In_80);
xor U4200 (N_4200,In_561,In_248);
xnor U4201 (N_4201,In_781,In_639);
or U4202 (N_4202,In_912,In_81);
nand U4203 (N_4203,In_772,In_1468);
and U4204 (N_4204,In_267,In_1005);
nand U4205 (N_4205,In_1422,In_1370);
and U4206 (N_4206,In_785,In_1780);
and U4207 (N_4207,In_327,In_1816);
nand U4208 (N_4208,In_484,In_148);
and U4209 (N_4209,In_553,In_1424);
nand U4210 (N_4210,In_338,In_541);
xor U4211 (N_4211,In_248,In_135);
xor U4212 (N_4212,In_985,In_628);
and U4213 (N_4213,In_387,In_1104);
xor U4214 (N_4214,In_751,In_1215);
nor U4215 (N_4215,In_1305,In_294);
and U4216 (N_4216,In_1,In_980);
xnor U4217 (N_4217,In_1516,In_713);
nand U4218 (N_4218,In_1727,In_1488);
or U4219 (N_4219,In_628,In_670);
nand U4220 (N_4220,In_1822,In_1204);
and U4221 (N_4221,In_365,In_1778);
nor U4222 (N_4222,In_1069,In_1471);
xnor U4223 (N_4223,In_1759,In_1977);
xor U4224 (N_4224,In_1613,In_1);
xor U4225 (N_4225,In_1209,In_771);
or U4226 (N_4226,In_1079,In_364);
or U4227 (N_4227,In_1249,In_1919);
nand U4228 (N_4228,In_339,In_1511);
xnor U4229 (N_4229,In_1741,In_432);
or U4230 (N_4230,In_1417,In_577);
and U4231 (N_4231,In_1541,In_959);
and U4232 (N_4232,In_1632,In_1757);
or U4233 (N_4233,In_1229,In_1909);
nor U4234 (N_4234,In_176,In_1459);
nand U4235 (N_4235,In_1094,In_480);
or U4236 (N_4236,In_882,In_150);
or U4237 (N_4237,In_1964,In_951);
xnor U4238 (N_4238,In_359,In_637);
nor U4239 (N_4239,In_1093,In_950);
and U4240 (N_4240,In_457,In_651);
nand U4241 (N_4241,In_287,In_196);
nand U4242 (N_4242,In_5,In_1175);
or U4243 (N_4243,In_726,In_886);
nand U4244 (N_4244,In_1969,In_794);
xor U4245 (N_4245,In_1490,In_412);
and U4246 (N_4246,In_1666,In_796);
nor U4247 (N_4247,In_741,In_1338);
nor U4248 (N_4248,In_115,In_277);
nand U4249 (N_4249,In_1206,In_561);
or U4250 (N_4250,In_1393,In_1544);
or U4251 (N_4251,In_1796,In_820);
nor U4252 (N_4252,In_568,In_1697);
and U4253 (N_4253,In_1232,In_1505);
and U4254 (N_4254,In_1024,In_1844);
xor U4255 (N_4255,In_1235,In_1848);
or U4256 (N_4256,In_1376,In_1268);
xor U4257 (N_4257,In_1679,In_999);
or U4258 (N_4258,In_1012,In_1848);
xor U4259 (N_4259,In_1842,In_152);
nor U4260 (N_4260,In_1024,In_375);
and U4261 (N_4261,In_1628,In_1175);
xor U4262 (N_4262,In_1719,In_1301);
and U4263 (N_4263,In_208,In_935);
nor U4264 (N_4264,In_1489,In_623);
or U4265 (N_4265,In_262,In_117);
xnor U4266 (N_4266,In_997,In_1888);
nand U4267 (N_4267,In_1544,In_423);
or U4268 (N_4268,In_354,In_1478);
xor U4269 (N_4269,In_582,In_1421);
nor U4270 (N_4270,In_1154,In_1156);
or U4271 (N_4271,In_673,In_1256);
xor U4272 (N_4272,In_104,In_1156);
nor U4273 (N_4273,In_1072,In_800);
or U4274 (N_4274,In_550,In_497);
and U4275 (N_4275,In_674,In_535);
nand U4276 (N_4276,In_966,In_1059);
nand U4277 (N_4277,In_976,In_1475);
nor U4278 (N_4278,In_1661,In_1412);
xnor U4279 (N_4279,In_1166,In_500);
nand U4280 (N_4280,In_1362,In_1550);
or U4281 (N_4281,In_910,In_763);
nand U4282 (N_4282,In_113,In_316);
nor U4283 (N_4283,In_379,In_470);
and U4284 (N_4284,In_1898,In_1362);
or U4285 (N_4285,In_806,In_1346);
or U4286 (N_4286,In_1149,In_1312);
xor U4287 (N_4287,In_2,In_1160);
and U4288 (N_4288,In_425,In_1475);
and U4289 (N_4289,In_1752,In_639);
nand U4290 (N_4290,In_1014,In_767);
nand U4291 (N_4291,In_124,In_422);
and U4292 (N_4292,In_24,In_843);
nor U4293 (N_4293,In_557,In_364);
nand U4294 (N_4294,In_618,In_609);
xor U4295 (N_4295,In_287,In_429);
nor U4296 (N_4296,In_1020,In_635);
xor U4297 (N_4297,In_313,In_929);
or U4298 (N_4298,In_1827,In_1515);
xor U4299 (N_4299,In_546,In_837);
and U4300 (N_4300,In_224,In_36);
nor U4301 (N_4301,In_818,In_1432);
nand U4302 (N_4302,In_1463,In_461);
or U4303 (N_4303,In_384,In_1637);
nor U4304 (N_4304,In_969,In_1476);
xnor U4305 (N_4305,In_1563,In_1272);
or U4306 (N_4306,In_1428,In_1328);
nand U4307 (N_4307,In_36,In_37);
xnor U4308 (N_4308,In_1115,In_1080);
or U4309 (N_4309,In_1836,In_1079);
nand U4310 (N_4310,In_905,In_396);
or U4311 (N_4311,In_1128,In_339);
nand U4312 (N_4312,In_640,In_1148);
and U4313 (N_4313,In_1114,In_849);
and U4314 (N_4314,In_905,In_906);
nor U4315 (N_4315,In_1040,In_69);
or U4316 (N_4316,In_1611,In_1049);
xor U4317 (N_4317,In_692,In_700);
xor U4318 (N_4318,In_1593,In_593);
and U4319 (N_4319,In_332,In_147);
or U4320 (N_4320,In_1750,In_165);
xnor U4321 (N_4321,In_872,In_565);
nand U4322 (N_4322,In_1542,In_1399);
nand U4323 (N_4323,In_1990,In_397);
nand U4324 (N_4324,In_1702,In_1593);
or U4325 (N_4325,In_891,In_776);
nor U4326 (N_4326,In_1014,In_313);
or U4327 (N_4327,In_1919,In_1838);
and U4328 (N_4328,In_1862,In_1478);
and U4329 (N_4329,In_756,In_1968);
or U4330 (N_4330,In_1498,In_483);
nor U4331 (N_4331,In_1110,In_1598);
nand U4332 (N_4332,In_1665,In_1269);
and U4333 (N_4333,In_1896,In_603);
xnor U4334 (N_4334,In_1162,In_6);
xor U4335 (N_4335,In_196,In_550);
nor U4336 (N_4336,In_1546,In_504);
and U4337 (N_4337,In_912,In_1236);
xor U4338 (N_4338,In_1203,In_457);
nor U4339 (N_4339,In_1685,In_1557);
nand U4340 (N_4340,In_92,In_185);
or U4341 (N_4341,In_1002,In_1192);
and U4342 (N_4342,In_731,In_245);
or U4343 (N_4343,In_1653,In_20);
nand U4344 (N_4344,In_1628,In_240);
xnor U4345 (N_4345,In_1174,In_1024);
nor U4346 (N_4346,In_1966,In_514);
nor U4347 (N_4347,In_425,In_487);
nand U4348 (N_4348,In_1811,In_459);
or U4349 (N_4349,In_121,In_165);
or U4350 (N_4350,In_581,In_242);
nor U4351 (N_4351,In_667,In_1916);
and U4352 (N_4352,In_1773,In_614);
nand U4353 (N_4353,In_827,In_621);
nor U4354 (N_4354,In_626,In_703);
and U4355 (N_4355,In_1041,In_1583);
or U4356 (N_4356,In_1251,In_258);
nor U4357 (N_4357,In_285,In_899);
nor U4358 (N_4358,In_1694,In_832);
nor U4359 (N_4359,In_147,In_357);
or U4360 (N_4360,In_1241,In_859);
nand U4361 (N_4361,In_1489,In_239);
nand U4362 (N_4362,In_335,In_1859);
nor U4363 (N_4363,In_1686,In_1066);
nand U4364 (N_4364,In_1130,In_351);
nand U4365 (N_4365,In_983,In_1842);
and U4366 (N_4366,In_178,In_949);
nand U4367 (N_4367,In_415,In_167);
or U4368 (N_4368,In_311,In_637);
nand U4369 (N_4369,In_395,In_1418);
xor U4370 (N_4370,In_2,In_622);
and U4371 (N_4371,In_1816,In_540);
and U4372 (N_4372,In_1737,In_40);
and U4373 (N_4373,In_1169,In_923);
xnor U4374 (N_4374,In_102,In_1068);
xor U4375 (N_4375,In_1416,In_1551);
nand U4376 (N_4376,In_700,In_1565);
nor U4377 (N_4377,In_1679,In_86);
nor U4378 (N_4378,In_1473,In_1885);
and U4379 (N_4379,In_449,In_450);
nand U4380 (N_4380,In_1973,In_1419);
or U4381 (N_4381,In_1971,In_1763);
and U4382 (N_4382,In_1089,In_89);
xor U4383 (N_4383,In_595,In_1415);
and U4384 (N_4384,In_482,In_271);
xor U4385 (N_4385,In_1489,In_704);
and U4386 (N_4386,In_335,In_240);
xnor U4387 (N_4387,In_567,In_1198);
nand U4388 (N_4388,In_271,In_1287);
xnor U4389 (N_4389,In_481,In_1729);
nor U4390 (N_4390,In_1056,In_1286);
xor U4391 (N_4391,In_1,In_1466);
nor U4392 (N_4392,In_137,In_1042);
or U4393 (N_4393,In_889,In_292);
nand U4394 (N_4394,In_141,In_1226);
nor U4395 (N_4395,In_233,In_1362);
and U4396 (N_4396,In_1662,In_1824);
and U4397 (N_4397,In_503,In_1865);
or U4398 (N_4398,In_868,In_1929);
nor U4399 (N_4399,In_1315,In_592);
and U4400 (N_4400,In_1725,In_432);
or U4401 (N_4401,In_1645,In_271);
nand U4402 (N_4402,In_786,In_1616);
or U4403 (N_4403,In_985,In_1099);
nand U4404 (N_4404,In_1874,In_1619);
and U4405 (N_4405,In_1916,In_1897);
nor U4406 (N_4406,In_515,In_346);
or U4407 (N_4407,In_1033,In_1238);
nand U4408 (N_4408,In_1479,In_677);
and U4409 (N_4409,In_788,In_1934);
or U4410 (N_4410,In_755,In_1163);
nand U4411 (N_4411,In_1982,In_1472);
nor U4412 (N_4412,In_716,In_1082);
or U4413 (N_4413,In_1682,In_41);
nor U4414 (N_4414,In_1163,In_361);
nor U4415 (N_4415,In_146,In_74);
nor U4416 (N_4416,In_1545,In_1073);
and U4417 (N_4417,In_1731,In_1776);
nor U4418 (N_4418,In_1237,In_286);
xor U4419 (N_4419,In_1093,In_1734);
nand U4420 (N_4420,In_697,In_44);
nand U4421 (N_4421,In_856,In_951);
nand U4422 (N_4422,In_888,In_406);
nand U4423 (N_4423,In_1675,In_1449);
xor U4424 (N_4424,In_1622,In_1851);
nor U4425 (N_4425,In_1502,In_540);
or U4426 (N_4426,In_1385,In_866);
xnor U4427 (N_4427,In_515,In_466);
nand U4428 (N_4428,In_834,In_1303);
xnor U4429 (N_4429,In_929,In_990);
nand U4430 (N_4430,In_1583,In_1701);
or U4431 (N_4431,In_1454,In_1670);
nand U4432 (N_4432,In_1474,In_1768);
and U4433 (N_4433,In_1349,In_1096);
nand U4434 (N_4434,In_1044,In_1042);
nor U4435 (N_4435,In_1037,In_79);
or U4436 (N_4436,In_58,In_398);
and U4437 (N_4437,In_1947,In_1635);
or U4438 (N_4438,In_338,In_1986);
and U4439 (N_4439,In_1917,In_819);
nand U4440 (N_4440,In_1388,In_241);
nor U4441 (N_4441,In_571,In_127);
or U4442 (N_4442,In_1830,In_730);
xnor U4443 (N_4443,In_1627,In_1816);
nand U4444 (N_4444,In_728,In_898);
nand U4445 (N_4445,In_1841,In_1237);
nor U4446 (N_4446,In_1049,In_14);
nor U4447 (N_4447,In_1340,In_282);
xor U4448 (N_4448,In_1238,In_1858);
and U4449 (N_4449,In_1696,In_1086);
nand U4450 (N_4450,In_1642,In_1975);
and U4451 (N_4451,In_1930,In_181);
or U4452 (N_4452,In_970,In_405);
or U4453 (N_4453,In_181,In_439);
and U4454 (N_4454,In_1715,In_24);
nand U4455 (N_4455,In_1993,In_1716);
xor U4456 (N_4456,In_66,In_1188);
or U4457 (N_4457,In_910,In_1653);
nor U4458 (N_4458,In_946,In_557);
xor U4459 (N_4459,In_1995,In_1909);
and U4460 (N_4460,In_890,In_733);
and U4461 (N_4461,In_423,In_1321);
nand U4462 (N_4462,In_1899,In_911);
nor U4463 (N_4463,In_1979,In_1608);
xnor U4464 (N_4464,In_468,In_115);
nor U4465 (N_4465,In_256,In_1044);
and U4466 (N_4466,In_562,In_1404);
or U4467 (N_4467,In_1080,In_1543);
or U4468 (N_4468,In_923,In_397);
nor U4469 (N_4469,In_1315,In_1922);
nand U4470 (N_4470,In_514,In_100);
or U4471 (N_4471,In_971,In_1215);
nand U4472 (N_4472,In_684,In_1093);
and U4473 (N_4473,In_1988,In_1390);
xnor U4474 (N_4474,In_1311,In_668);
or U4475 (N_4475,In_1999,In_1706);
xnor U4476 (N_4476,In_422,In_1961);
xnor U4477 (N_4477,In_1875,In_452);
nand U4478 (N_4478,In_730,In_728);
and U4479 (N_4479,In_1625,In_413);
nor U4480 (N_4480,In_507,In_330);
nand U4481 (N_4481,In_1721,In_865);
nor U4482 (N_4482,In_908,In_1695);
nor U4483 (N_4483,In_1697,In_914);
xor U4484 (N_4484,In_1521,In_1308);
nand U4485 (N_4485,In_252,In_306);
and U4486 (N_4486,In_475,In_676);
and U4487 (N_4487,In_237,In_1281);
nand U4488 (N_4488,In_481,In_164);
or U4489 (N_4489,In_55,In_1786);
nor U4490 (N_4490,In_1031,In_1066);
or U4491 (N_4491,In_680,In_1900);
nand U4492 (N_4492,In_1023,In_853);
and U4493 (N_4493,In_1669,In_1207);
xnor U4494 (N_4494,In_840,In_864);
nor U4495 (N_4495,In_1842,In_1391);
xor U4496 (N_4496,In_1746,In_505);
nor U4497 (N_4497,In_105,In_36);
xor U4498 (N_4498,In_211,In_1850);
and U4499 (N_4499,In_825,In_1417);
nor U4500 (N_4500,In_124,In_765);
nor U4501 (N_4501,In_692,In_434);
nand U4502 (N_4502,In_646,In_243);
nor U4503 (N_4503,In_1420,In_756);
nor U4504 (N_4504,In_735,In_1137);
or U4505 (N_4505,In_699,In_180);
nor U4506 (N_4506,In_1384,In_298);
and U4507 (N_4507,In_1018,In_1274);
nor U4508 (N_4508,In_726,In_165);
and U4509 (N_4509,In_1287,In_1315);
xnor U4510 (N_4510,In_738,In_1958);
or U4511 (N_4511,In_474,In_1464);
nand U4512 (N_4512,In_1662,In_612);
and U4513 (N_4513,In_477,In_863);
xor U4514 (N_4514,In_136,In_1940);
xnor U4515 (N_4515,In_952,In_53);
nand U4516 (N_4516,In_328,In_940);
nand U4517 (N_4517,In_357,In_527);
nor U4518 (N_4518,In_506,In_1902);
xnor U4519 (N_4519,In_1584,In_1759);
and U4520 (N_4520,In_997,In_1053);
xor U4521 (N_4521,In_575,In_1619);
nor U4522 (N_4522,In_431,In_370);
nor U4523 (N_4523,In_845,In_1644);
nand U4524 (N_4524,In_155,In_425);
xor U4525 (N_4525,In_5,In_338);
xor U4526 (N_4526,In_1486,In_1751);
xnor U4527 (N_4527,In_1055,In_1155);
xnor U4528 (N_4528,In_914,In_680);
nor U4529 (N_4529,In_1537,In_1643);
or U4530 (N_4530,In_1787,In_1881);
xnor U4531 (N_4531,In_1864,In_1911);
or U4532 (N_4532,In_1467,In_1250);
and U4533 (N_4533,In_1989,In_1547);
nand U4534 (N_4534,In_496,In_1480);
nand U4535 (N_4535,In_992,In_1724);
xnor U4536 (N_4536,In_138,In_1282);
xor U4537 (N_4537,In_501,In_1870);
xor U4538 (N_4538,In_1634,In_1293);
nor U4539 (N_4539,In_667,In_875);
or U4540 (N_4540,In_1628,In_656);
or U4541 (N_4541,In_495,In_205);
nand U4542 (N_4542,In_1356,In_1753);
nor U4543 (N_4543,In_803,In_2);
or U4544 (N_4544,In_1033,In_63);
and U4545 (N_4545,In_1874,In_1024);
nand U4546 (N_4546,In_1385,In_10);
nor U4547 (N_4547,In_636,In_313);
and U4548 (N_4548,In_944,In_1676);
nor U4549 (N_4549,In_872,In_169);
and U4550 (N_4550,In_363,In_283);
or U4551 (N_4551,In_633,In_848);
or U4552 (N_4552,In_149,In_1848);
xor U4553 (N_4553,In_1704,In_735);
or U4554 (N_4554,In_1616,In_1843);
or U4555 (N_4555,In_343,In_1969);
xor U4556 (N_4556,In_1409,In_404);
nand U4557 (N_4557,In_19,In_1191);
nor U4558 (N_4558,In_540,In_953);
or U4559 (N_4559,In_245,In_693);
or U4560 (N_4560,In_752,In_1454);
or U4561 (N_4561,In_311,In_1728);
and U4562 (N_4562,In_1076,In_1687);
or U4563 (N_4563,In_1926,In_981);
or U4564 (N_4564,In_1816,In_535);
xnor U4565 (N_4565,In_1404,In_965);
nand U4566 (N_4566,In_760,In_1396);
or U4567 (N_4567,In_1016,In_1854);
nand U4568 (N_4568,In_1376,In_1757);
or U4569 (N_4569,In_564,In_46);
and U4570 (N_4570,In_417,In_203);
nor U4571 (N_4571,In_871,In_468);
nor U4572 (N_4572,In_323,In_1723);
nand U4573 (N_4573,In_1701,In_70);
nand U4574 (N_4574,In_584,In_658);
nor U4575 (N_4575,In_574,In_373);
xnor U4576 (N_4576,In_407,In_1711);
or U4577 (N_4577,In_1123,In_293);
and U4578 (N_4578,In_259,In_376);
nor U4579 (N_4579,In_66,In_825);
or U4580 (N_4580,In_1773,In_1284);
and U4581 (N_4581,In_319,In_1833);
and U4582 (N_4582,In_1040,In_1045);
and U4583 (N_4583,In_811,In_369);
and U4584 (N_4584,In_354,In_812);
nand U4585 (N_4585,In_555,In_1627);
nor U4586 (N_4586,In_991,In_1084);
or U4587 (N_4587,In_1331,In_678);
nor U4588 (N_4588,In_877,In_405);
nand U4589 (N_4589,In_1751,In_1298);
or U4590 (N_4590,In_1941,In_352);
or U4591 (N_4591,In_1754,In_1919);
xnor U4592 (N_4592,In_383,In_1576);
and U4593 (N_4593,In_1863,In_742);
nor U4594 (N_4594,In_900,In_694);
and U4595 (N_4595,In_849,In_1450);
and U4596 (N_4596,In_1108,In_1710);
xnor U4597 (N_4597,In_287,In_1586);
nor U4598 (N_4598,In_1350,In_1644);
and U4599 (N_4599,In_152,In_421);
nand U4600 (N_4600,In_1296,In_522);
nand U4601 (N_4601,In_563,In_380);
and U4602 (N_4602,In_1706,In_949);
xor U4603 (N_4603,In_1454,In_709);
or U4604 (N_4604,In_228,In_1112);
nand U4605 (N_4605,In_1657,In_562);
nand U4606 (N_4606,In_674,In_858);
xor U4607 (N_4607,In_71,In_1204);
or U4608 (N_4608,In_369,In_1768);
and U4609 (N_4609,In_1144,In_902);
nand U4610 (N_4610,In_1086,In_1602);
nand U4611 (N_4611,In_1831,In_1496);
nand U4612 (N_4612,In_66,In_196);
nor U4613 (N_4613,In_578,In_78);
or U4614 (N_4614,In_1398,In_1632);
nand U4615 (N_4615,In_1563,In_534);
or U4616 (N_4616,In_753,In_1468);
and U4617 (N_4617,In_496,In_1949);
or U4618 (N_4618,In_608,In_1199);
and U4619 (N_4619,In_334,In_161);
nand U4620 (N_4620,In_207,In_310);
nor U4621 (N_4621,In_204,In_1328);
xor U4622 (N_4622,In_1202,In_645);
nand U4623 (N_4623,In_54,In_804);
nand U4624 (N_4624,In_1085,In_1876);
xor U4625 (N_4625,In_509,In_679);
and U4626 (N_4626,In_449,In_332);
or U4627 (N_4627,In_1269,In_1175);
nor U4628 (N_4628,In_408,In_996);
or U4629 (N_4629,In_108,In_1884);
nor U4630 (N_4630,In_1872,In_1069);
nor U4631 (N_4631,In_781,In_1752);
and U4632 (N_4632,In_762,In_1094);
or U4633 (N_4633,In_1932,In_44);
nor U4634 (N_4634,In_1562,In_266);
and U4635 (N_4635,In_657,In_573);
or U4636 (N_4636,In_1455,In_1190);
xor U4637 (N_4637,In_617,In_637);
nand U4638 (N_4638,In_288,In_1557);
or U4639 (N_4639,In_683,In_826);
nor U4640 (N_4640,In_711,In_1860);
xnor U4641 (N_4641,In_1397,In_1813);
xnor U4642 (N_4642,In_1224,In_1689);
nand U4643 (N_4643,In_1621,In_1528);
and U4644 (N_4644,In_1514,In_434);
or U4645 (N_4645,In_392,In_638);
and U4646 (N_4646,In_795,In_284);
nor U4647 (N_4647,In_728,In_58);
and U4648 (N_4648,In_1999,In_841);
nand U4649 (N_4649,In_82,In_1318);
and U4650 (N_4650,In_270,In_1467);
xor U4651 (N_4651,In_1108,In_200);
xor U4652 (N_4652,In_342,In_708);
nand U4653 (N_4653,In_1267,In_1759);
and U4654 (N_4654,In_1217,In_379);
nand U4655 (N_4655,In_1169,In_158);
and U4656 (N_4656,In_538,In_956);
or U4657 (N_4657,In_451,In_396);
and U4658 (N_4658,In_1564,In_1106);
xnor U4659 (N_4659,In_506,In_606);
nor U4660 (N_4660,In_1430,In_1414);
nand U4661 (N_4661,In_458,In_1599);
nor U4662 (N_4662,In_206,In_784);
xor U4663 (N_4663,In_1505,In_1280);
nand U4664 (N_4664,In_1770,In_824);
nor U4665 (N_4665,In_816,In_337);
or U4666 (N_4666,In_1484,In_653);
or U4667 (N_4667,In_1985,In_348);
nand U4668 (N_4668,In_1690,In_919);
nand U4669 (N_4669,In_979,In_1415);
xnor U4670 (N_4670,In_1007,In_1438);
and U4671 (N_4671,In_1750,In_1926);
nor U4672 (N_4672,In_1779,In_163);
nand U4673 (N_4673,In_611,In_772);
xor U4674 (N_4674,In_370,In_1361);
nand U4675 (N_4675,In_1904,In_475);
or U4676 (N_4676,In_853,In_1171);
xnor U4677 (N_4677,In_1052,In_704);
and U4678 (N_4678,In_1464,In_1501);
nand U4679 (N_4679,In_269,In_313);
xnor U4680 (N_4680,In_873,In_172);
xor U4681 (N_4681,In_1718,In_557);
xnor U4682 (N_4682,In_61,In_1031);
and U4683 (N_4683,In_1068,In_1856);
nor U4684 (N_4684,In_1038,In_771);
xnor U4685 (N_4685,In_687,In_849);
nand U4686 (N_4686,In_1013,In_1460);
or U4687 (N_4687,In_1590,In_1743);
nand U4688 (N_4688,In_1079,In_416);
nor U4689 (N_4689,In_16,In_1125);
or U4690 (N_4690,In_1324,In_1590);
and U4691 (N_4691,In_1084,In_765);
and U4692 (N_4692,In_1663,In_979);
nand U4693 (N_4693,In_1798,In_506);
and U4694 (N_4694,In_698,In_1915);
nand U4695 (N_4695,In_604,In_1154);
or U4696 (N_4696,In_1844,In_1254);
nand U4697 (N_4697,In_1542,In_1317);
or U4698 (N_4698,In_885,In_93);
nand U4699 (N_4699,In_19,In_402);
or U4700 (N_4700,In_1029,In_1567);
or U4701 (N_4701,In_1710,In_1273);
and U4702 (N_4702,In_805,In_586);
or U4703 (N_4703,In_1322,In_1693);
xor U4704 (N_4704,In_605,In_563);
or U4705 (N_4705,In_1138,In_796);
and U4706 (N_4706,In_1246,In_1107);
xor U4707 (N_4707,In_1067,In_1619);
nand U4708 (N_4708,In_330,In_1510);
or U4709 (N_4709,In_1021,In_1967);
and U4710 (N_4710,In_1882,In_814);
nand U4711 (N_4711,In_1668,In_351);
xnor U4712 (N_4712,In_877,In_773);
and U4713 (N_4713,In_1547,In_915);
and U4714 (N_4714,In_807,In_1158);
or U4715 (N_4715,In_752,In_1949);
or U4716 (N_4716,In_814,In_145);
xor U4717 (N_4717,In_22,In_212);
xor U4718 (N_4718,In_864,In_158);
or U4719 (N_4719,In_1111,In_1363);
nor U4720 (N_4720,In_1151,In_780);
xor U4721 (N_4721,In_512,In_826);
nand U4722 (N_4722,In_119,In_1445);
nand U4723 (N_4723,In_1248,In_1745);
nor U4724 (N_4724,In_1848,In_758);
or U4725 (N_4725,In_838,In_657);
nand U4726 (N_4726,In_638,In_279);
xnor U4727 (N_4727,In_146,In_81);
nor U4728 (N_4728,In_1224,In_1014);
nand U4729 (N_4729,In_1077,In_650);
xnor U4730 (N_4730,In_106,In_38);
xor U4731 (N_4731,In_602,In_1669);
and U4732 (N_4732,In_1817,In_1657);
and U4733 (N_4733,In_1004,In_787);
and U4734 (N_4734,In_1220,In_1282);
or U4735 (N_4735,In_632,In_1871);
xor U4736 (N_4736,In_1668,In_652);
nand U4737 (N_4737,In_525,In_1476);
or U4738 (N_4738,In_1146,In_271);
nand U4739 (N_4739,In_672,In_481);
nor U4740 (N_4740,In_1089,In_341);
or U4741 (N_4741,In_843,In_1681);
or U4742 (N_4742,In_360,In_399);
and U4743 (N_4743,In_1311,In_451);
nand U4744 (N_4744,In_524,In_1548);
nor U4745 (N_4745,In_978,In_607);
xor U4746 (N_4746,In_1305,In_1288);
nand U4747 (N_4747,In_1280,In_486);
or U4748 (N_4748,In_574,In_37);
and U4749 (N_4749,In_1213,In_1017);
nor U4750 (N_4750,In_1991,In_220);
or U4751 (N_4751,In_335,In_1940);
xnor U4752 (N_4752,In_1143,In_270);
or U4753 (N_4753,In_1235,In_1893);
and U4754 (N_4754,In_836,In_1072);
nand U4755 (N_4755,In_253,In_1183);
and U4756 (N_4756,In_1068,In_908);
and U4757 (N_4757,In_54,In_1615);
xor U4758 (N_4758,In_1006,In_1290);
nor U4759 (N_4759,In_760,In_1363);
or U4760 (N_4760,In_1734,In_992);
nand U4761 (N_4761,In_245,In_1705);
nor U4762 (N_4762,In_1328,In_1057);
xor U4763 (N_4763,In_1460,In_1897);
and U4764 (N_4764,In_1654,In_1151);
and U4765 (N_4765,In_1479,In_1275);
or U4766 (N_4766,In_55,In_1121);
nand U4767 (N_4767,In_1121,In_846);
xnor U4768 (N_4768,In_695,In_790);
xnor U4769 (N_4769,In_453,In_911);
or U4770 (N_4770,In_247,In_1900);
nand U4771 (N_4771,In_1225,In_470);
nand U4772 (N_4772,In_576,In_1594);
or U4773 (N_4773,In_1653,In_1840);
and U4774 (N_4774,In_914,In_1387);
nand U4775 (N_4775,In_833,In_217);
nand U4776 (N_4776,In_1962,In_498);
and U4777 (N_4777,In_1371,In_1252);
and U4778 (N_4778,In_339,In_1988);
xor U4779 (N_4779,In_715,In_1895);
or U4780 (N_4780,In_1057,In_646);
nand U4781 (N_4781,In_228,In_214);
or U4782 (N_4782,In_1904,In_176);
nor U4783 (N_4783,In_1530,In_565);
xor U4784 (N_4784,In_250,In_1691);
nand U4785 (N_4785,In_395,In_1967);
nor U4786 (N_4786,In_1310,In_78);
and U4787 (N_4787,In_377,In_1042);
nor U4788 (N_4788,In_744,In_170);
nand U4789 (N_4789,In_1967,In_831);
nor U4790 (N_4790,In_571,In_1447);
and U4791 (N_4791,In_1774,In_1910);
nor U4792 (N_4792,In_1227,In_1310);
or U4793 (N_4793,In_285,In_1553);
nor U4794 (N_4794,In_29,In_660);
nand U4795 (N_4795,In_588,In_961);
and U4796 (N_4796,In_1561,In_1118);
or U4797 (N_4797,In_133,In_600);
and U4798 (N_4798,In_1224,In_141);
nor U4799 (N_4799,In_752,In_279);
nand U4800 (N_4800,In_788,In_1580);
nor U4801 (N_4801,In_68,In_968);
and U4802 (N_4802,In_243,In_966);
xnor U4803 (N_4803,In_502,In_956);
nor U4804 (N_4804,In_1966,In_1894);
nand U4805 (N_4805,In_1075,In_1313);
nand U4806 (N_4806,In_1766,In_908);
xor U4807 (N_4807,In_1745,In_1900);
xor U4808 (N_4808,In_513,In_1884);
nor U4809 (N_4809,In_1636,In_194);
and U4810 (N_4810,In_1669,In_401);
and U4811 (N_4811,In_1646,In_278);
or U4812 (N_4812,In_170,In_1279);
and U4813 (N_4813,In_152,In_579);
nand U4814 (N_4814,In_1782,In_1696);
nor U4815 (N_4815,In_476,In_1582);
or U4816 (N_4816,In_457,In_233);
and U4817 (N_4817,In_1763,In_676);
and U4818 (N_4818,In_1564,In_207);
xnor U4819 (N_4819,In_873,In_1879);
and U4820 (N_4820,In_1099,In_358);
or U4821 (N_4821,In_1197,In_1717);
xor U4822 (N_4822,In_1918,In_1127);
and U4823 (N_4823,In_1186,In_1244);
or U4824 (N_4824,In_814,In_676);
nand U4825 (N_4825,In_1990,In_1509);
or U4826 (N_4826,In_1957,In_1244);
nor U4827 (N_4827,In_547,In_1130);
xnor U4828 (N_4828,In_610,In_629);
and U4829 (N_4829,In_1581,In_1959);
nor U4830 (N_4830,In_1351,In_1528);
nor U4831 (N_4831,In_960,In_1991);
xor U4832 (N_4832,In_1813,In_1711);
and U4833 (N_4833,In_729,In_614);
and U4834 (N_4834,In_1095,In_293);
or U4835 (N_4835,In_870,In_1085);
and U4836 (N_4836,In_1422,In_234);
or U4837 (N_4837,In_133,In_1391);
and U4838 (N_4838,In_124,In_1885);
xnor U4839 (N_4839,In_1831,In_592);
or U4840 (N_4840,In_59,In_553);
xnor U4841 (N_4841,In_1538,In_1032);
xor U4842 (N_4842,In_246,In_1697);
nand U4843 (N_4843,In_1108,In_1030);
or U4844 (N_4844,In_215,In_897);
xor U4845 (N_4845,In_1954,In_1807);
nor U4846 (N_4846,In_712,In_1317);
nor U4847 (N_4847,In_590,In_733);
nand U4848 (N_4848,In_719,In_454);
or U4849 (N_4849,In_1150,In_591);
nor U4850 (N_4850,In_1919,In_407);
or U4851 (N_4851,In_234,In_1238);
or U4852 (N_4852,In_1083,In_1242);
xnor U4853 (N_4853,In_19,In_127);
xor U4854 (N_4854,In_723,In_1362);
and U4855 (N_4855,In_325,In_633);
nand U4856 (N_4856,In_451,In_885);
nor U4857 (N_4857,In_1604,In_1556);
xnor U4858 (N_4858,In_773,In_1300);
nand U4859 (N_4859,In_547,In_676);
nor U4860 (N_4860,In_1715,In_1206);
or U4861 (N_4861,In_1692,In_216);
or U4862 (N_4862,In_886,In_1302);
and U4863 (N_4863,In_1570,In_47);
or U4864 (N_4864,In_689,In_581);
or U4865 (N_4865,In_877,In_414);
and U4866 (N_4866,In_1068,In_1556);
and U4867 (N_4867,In_1695,In_1649);
and U4868 (N_4868,In_160,In_404);
xor U4869 (N_4869,In_63,In_1765);
xor U4870 (N_4870,In_1751,In_1547);
and U4871 (N_4871,In_1694,In_1759);
and U4872 (N_4872,In_1183,In_1818);
nand U4873 (N_4873,In_465,In_863);
and U4874 (N_4874,In_25,In_881);
or U4875 (N_4875,In_210,In_915);
or U4876 (N_4876,In_552,In_1032);
nand U4877 (N_4877,In_313,In_752);
and U4878 (N_4878,In_1401,In_1429);
nor U4879 (N_4879,In_86,In_1132);
and U4880 (N_4880,In_1718,In_1557);
or U4881 (N_4881,In_1586,In_335);
and U4882 (N_4882,In_938,In_1622);
or U4883 (N_4883,In_1812,In_1941);
nand U4884 (N_4884,In_279,In_924);
and U4885 (N_4885,In_1345,In_1531);
nor U4886 (N_4886,In_1711,In_232);
and U4887 (N_4887,In_404,In_1125);
xnor U4888 (N_4888,In_1562,In_1487);
or U4889 (N_4889,In_1794,In_814);
xor U4890 (N_4890,In_964,In_1609);
and U4891 (N_4891,In_414,In_1803);
or U4892 (N_4892,In_1414,In_776);
or U4893 (N_4893,In_1391,In_1885);
xor U4894 (N_4894,In_1420,In_1663);
nand U4895 (N_4895,In_1151,In_1973);
or U4896 (N_4896,In_1544,In_587);
or U4897 (N_4897,In_1260,In_1147);
and U4898 (N_4898,In_388,In_938);
nor U4899 (N_4899,In_1734,In_717);
and U4900 (N_4900,In_251,In_632);
nor U4901 (N_4901,In_865,In_1200);
xnor U4902 (N_4902,In_1993,In_591);
and U4903 (N_4903,In_1321,In_1554);
xnor U4904 (N_4904,In_972,In_281);
nor U4905 (N_4905,In_514,In_633);
xnor U4906 (N_4906,In_132,In_1278);
or U4907 (N_4907,In_1973,In_1472);
xor U4908 (N_4908,In_1584,In_1776);
xnor U4909 (N_4909,In_971,In_684);
and U4910 (N_4910,In_990,In_1396);
nand U4911 (N_4911,In_872,In_998);
nand U4912 (N_4912,In_840,In_108);
nor U4913 (N_4913,In_1377,In_293);
nor U4914 (N_4914,In_1968,In_1367);
nor U4915 (N_4915,In_90,In_1755);
xnor U4916 (N_4916,In_707,In_199);
or U4917 (N_4917,In_1280,In_1789);
xnor U4918 (N_4918,In_831,In_1320);
nand U4919 (N_4919,In_1250,In_715);
nor U4920 (N_4920,In_1005,In_1295);
nand U4921 (N_4921,In_1545,In_1030);
or U4922 (N_4922,In_1884,In_833);
nor U4923 (N_4923,In_1676,In_1942);
and U4924 (N_4924,In_81,In_1891);
or U4925 (N_4925,In_1419,In_1405);
and U4926 (N_4926,In_507,In_1337);
or U4927 (N_4927,In_1068,In_309);
or U4928 (N_4928,In_1162,In_569);
nor U4929 (N_4929,In_253,In_607);
and U4930 (N_4930,In_1422,In_1675);
nand U4931 (N_4931,In_1910,In_1747);
nor U4932 (N_4932,In_428,In_502);
or U4933 (N_4933,In_1344,In_1347);
nor U4934 (N_4934,In_1252,In_1087);
or U4935 (N_4935,In_1619,In_75);
nand U4936 (N_4936,In_938,In_1167);
or U4937 (N_4937,In_285,In_1176);
xnor U4938 (N_4938,In_179,In_752);
or U4939 (N_4939,In_886,In_1110);
or U4940 (N_4940,In_1940,In_154);
nor U4941 (N_4941,In_737,In_18);
xor U4942 (N_4942,In_577,In_1034);
nand U4943 (N_4943,In_639,In_862);
nor U4944 (N_4944,In_1428,In_1589);
and U4945 (N_4945,In_1951,In_1174);
and U4946 (N_4946,In_1494,In_226);
nor U4947 (N_4947,In_1429,In_1163);
and U4948 (N_4948,In_203,In_329);
nor U4949 (N_4949,In_1542,In_1318);
nand U4950 (N_4950,In_255,In_1015);
xnor U4951 (N_4951,In_1748,In_1656);
xor U4952 (N_4952,In_142,In_1361);
and U4953 (N_4953,In_1784,In_1537);
or U4954 (N_4954,In_481,In_1942);
and U4955 (N_4955,In_600,In_1280);
or U4956 (N_4956,In_882,In_496);
nor U4957 (N_4957,In_1286,In_1563);
nand U4958 (N_4958,In_1254,In_727);
nor U4959 (N_4959,In_446,In_873);
nand U4960 (N_4960,In_309,In_1078);
and U4961 (N_4961,In_1858,In_1374);
xor U4962 (N_4962,In_557,In_1041);
nand U4963 (N_4963,In_1081,In_1483);
nand U4964 (N_4964,In_1762,In_231);
and U4965 (N_4965,In_732,In_1116);
nor U4966 (N_4966,In_2,In_1825);
and U4967 (N_4967,In_491,In_74);
xnor U4968 (N_4968,In_1043,In_1219);
nand U4969 (N_4969,In_1785,In_660);
nand U4970 (N_4970,In_1841,In_995);
nor U4971 (N_4971,In_1859,In_1776);
nand U4972 (N_4972,In_1632,In_1899);
nand U4973 (N_4973,In_543,In_1218);
xor U4974 (N_4974,In_163,In_571);
nor U4975 (N_4975,In_386,In_1367);
or U4976 (N_4976,In_158,In_1991);
nor U4977 (N_4977,In_676,In_1183);
nor U4978 (N_4978,In_369,In_1505);
xor U4979 (N_4979,In_737,In_1906);
nor U4980 (N_4980,In_146,In_1598);
nor U4981 (N_4981,In_437,In_1304);
xor U4982 (N_4982,In_862,In_301);
or U4983 (N_4983,In_162,In_1381);
nor U4984 (N_4984,In_603,In_571);
and U4985 (N_4985,In_1872,In_1840);
or U4986 (N_4986,In_804,In_1907);
nand U4987 (N_4987,In_1937,In_1541);
or U4988 (N_4988,In_1017,In_988);
nor U4989 (N_4989,In_1156,In_403);
or U4990 (N_4990,In_1524,In_1741);
and U4991 (N_4991,In_670,In_1766);
or U4992 (N_4992,In_699,In_104);
xor U4993 (N_4993,In_1355,In_997);
or U4994 (N_4994,In_506,In_540);
xnor U4995 (N_4995,In_126,In_1362);
nor U4996 (N_4996,In_174,In_1754);
nand U4997 (N_4997,In_1937,In_1574);
and U4998 (N_4998,In_567,In_1053);
xnor U4999 (N_4999,In_158,In_769);
and U5000 (N_5000,N_131,N_2824);
or U5001 (N_5001,N_1314,N_3483);
nand U5002 (N_5002,N_3945,N_16);
or U5003 (N_5003,N_3665,N_702);
xor U5004 (N_5004,N_2160,N_90);
nand U5005 (N_5005,N_3768,N_2471);
nor U5006 (N_5006,N_4716,N_1418);
and U5007 (N_5007,N_966,N_2939);
or U5008 (N_5008,N_1184,N_183);
nor U5009 (N_5009,N_2379,N_1895);
nand U5010 (N_5010,N_4123,N_1166);
xor U5011 (N_5011,N_810,N_4974);
xor U5012 (N_5012,N_4564,N_520);
xnor U5013 (N_5013,N_219,N_1967);
nand U5014 (N_5014,N_715,N_2860);
and U5015 (N_5015,N_3480,N_3792);
nor U5016 (N_5016,N_3967,N_3084);
nor U5017 (N_5017,N_1701,N_2745);
nand U5018 (N_5018,N_4815,N_3740);
or U5019 (N_5019,N_4534,N_2317);
or U5020 (N_5020,N_2342,N_4688);
nor U5021 (N_5021,N_1082,N_3338);
and U5022 (N_5022,N_828,N_2215);
xor U5023 (N_5023,N_4099,N_2113);
and U5024 (N_5024,N_3572,N_2734);
nand U5025 (N_5025,N_2040,N_4195);
nor U5026 (N_5026,N_1815,N_3699);
xor U5027 (N_5027,N_4991,N_1442);
nand U5028 (N_5028,N_4738,N_3948);
xor U5029 (N_5029,N_491,N_2462);
and U5030 (N_5030,N_3456,N_4510);
or U5031 (N_5031,N_2224,N_4206);
xnor U5032 (N_5032,N_859,N_2764);
or U5033 (N_5033,N_3309,N_4545);
xor U5034 (N_5034,N_3494,N_1186);
and U5035 (N_5035,N_3303,N_1987);
or U5036 (N_5036,N_4365,N_4438);
nor U5037 (N_5037,N_1041,N_1250);
xor U5038 (N_5038,N_1127,N_891);
nand U5039 (N_5039,N_2509,N_4236);
xor U5040 (N_5040,N_3368,N_2136);
and U5041 (N_5041,N_714,N_3019);
or U5042 (N_5042,N_3342,N_3474);
and U5043 (N_5043,N_2754,N_2085);
or U5044 (N_5044,N_4388,N_963);
or U5045 (N_5045,N_4211,N_4913);
and U5046 (N_5046,N_2870,N_2432);
nor U5047 (N_5047,N_2909,N_2408);
xnor U5048 (N_5048,N_2024,N_140);
or U5049 (N_5049,N_2896,N_1215);
or U5050 (N_5050,N_2826,N_141);
nor U5051 (N_5051,N_2715,N_2535);
and U5052 (N_5052,N_3607,N_2131);
nand U5053 (N_5053,N_1173,N_236);
nor U5054 (N_5054,N_433,N_4932);
nor U5055 (N_5055,N_3915,N_592);
nor U5056 (N_5056,N_4647,N_1447);
nand U5057 (N_5057,N_1934,N_92);
nand U5058 (N_5058,N_575,N_154);
nor U5059 (N_5059,N_3934,N_1950);
and U5060 (N_5060,N_1362,N_2485);
nand U5061 (N_5061,N_3476,N_1993);
xnor U5062 (N_5062,N_4850,N_1309);
and U5063 (N_5063,N_3179,N_1274);
xor U5064 (N_5064,N_3714,N_4531);
and U5065 (N_5065,N_4418,N_3761);
nand U5066 (N_5066,N_3955,N_1241);
or U5067 (N_5067,N_4501,N_1907);
nor U5068 (N_5068,N_4275,N_3029);
and U5069 (N_5069,N_1552,N_685);
or U5070 (N_5070,N_1292,N_4020);
nand U5071 (N_5071,N_4617,N_4081);
nor U5072 (N_5072,N_1549,N_560);
nor U5073 (N_5073,N_3207,N_1631);
or U5074 (N_5074,N_2563,N_1461);
or U5075 (N_5075,N_4451,N_2256);
nand U5076 (N_5076,N_4906,N_1608);
nand U5077 (N_5077,N_4638,N_4892);
or U5078 (N_5078,N_3448,N_4273);
nor U5079 (N_5079,N_1755,N_264);
or U5080 (N_5080,N_3721,N_768);
and U5081 (N_5081,N_1900,N_1172);
nor U5082 (N_5082,N_1026,N_2114);
or U5083 (N_5083,N_375,N_1556);
or U5084 (N_5084,N_3775,N_3887);
and U5085 (N_5085,N_4577,N_4225);
or U5086 (N_5086,N_1330,N_2003);
nand U5087 (N_5087,N_589,N_2547);
nand U5088 (N_5088,N_3956,N_2956);
or U5089 (N_5089,N_690,N_2167);
nor U5090 (N_5090,N_2526,N_3249);
and U5091 (N_5091,N_4166,N_1405);
or U5092 (N_5092,N_4216,N_1092);
nor U5093 (N_5093,N_2900,N_1199);
and U5094 (N_5094,N_4299,N_477);
nand U5095 (N_5095,N_4823,N_280);
xor U5096 (N_5096,N_688,N_3575);
xor U5097 (N_5097,N_4477,N_3914);
nor U5098 (N_5098,N_306,N_3904);
and U5099 (N_5099,N_2952,N_1159);
nand U5100 (N_5100,N_788,N_1270);
and U5101 (N_5101,N_1410,N_1775);
xor U5102 (N_5102,N_4804,N_4491);
and U5103 (N_5103,N_3757,N_3841);
or U5104 (N_5104,N_3522,N_4851);
and U5105 (N_5105,N_510,N_4046);
nand U5106 (N_5106,N_4979,N_4652);
nor U5107 (N_5107,N_2857,N_4915);
and U5108 (N_5108,N_635,N_3534);
or U5109 (N_5109,N_2498,N_4471);
nand U5110 (N_5110,N_3846,N_1167);
or U5111 (N_5111,N_1034,N_1211);
or U5112 (N_5112,N_1102,N_2912);
or U5113 (N_5113,N_1668,N_4818);
xor U5114 (N_5114,N_3178,N_4393);
nand U5115 (N_5115,N_1814,N_3781);
nor U5116 (N_5116,N_3739,N_2991);
and U5117 (N_5117,N_826,N_350);
nand U5118 (N_5118,N_1196,N_4654);
and U5119 (N_5119,N_578,N_4676);
and U5120 (N_5120,N_2274,N_2959);
nand U5121 (N_5121,N_1933,N_1391);
nand U5122 (N_5122,N_1408,N_351);
nand U5123 (N_5123,N_1536,N_118);
nor U5124 (N_5124,N_1426,N_3732);
or U5125 (N_5125,N_921,N_1770);
and U5126 (N_5126,N_2493,N_3300);
and U5127 (N_5127,N_3095,N_3795);
nor U5128 (N_5128,N_4893,N_3843);
xor U5129 (N_5129,N_4542,N_3911);
and U5130 (N_5130,N_656,N_2648);
xor U5131 (N_5131,N_4726,N_2640);
xor U5132 (N_5132,N_3229,N_2564);
xor U5133 (N_5133,N_2869,N_2825);
or U5134 (N_5134,N_1918,N_823);
nand U5135 (N_5135,N_1020,N_3692);
nor U5136 (N_5136,N_627,N_1229);
nor U5137 (N_5137,N_2793,N_3439);
nor U5138 (N_5138,N_907,N_2183);
and U5139 (N_5139,N_2657,N_431);
nor U5140 (N_5140,N_3579,N_2185);
or U5141 (N_5141,N_3743,N_3432);
and U5142 (N_5142,N_1928,N_4172);
and U5143 (N_5143,N_298,N_4694);
and U5144 (N_5144,N_465,N_3723);
nor U5145 (N_5145,N_1824,N_1339);
xor U5146 (N_5146,N_1619,N_300);
nand U5147 (N_5147,N_2496,N_106);
and U5148 (N_5148,N_240,N_205);
or U5149 (N_5149,N_109,N_1085);
xor U5150 (N_5150,N_792,N_4079);
nand U5151 (N_5151,N_3312,N_2931);
xnor U5152 (N_5152,N_2922,N_3899);
nand U5153 (N_5153,N_4343,N_533);
xor U5154 (N_5154,N_3282,N_3489);
nor U5155 (N_5155,N_1525,N_3141);
nand U5156 (N_5156,N_3298,N_912);
xor U5157 (N_5157,N_1198,N_2382);
nor U5158 (N_5158,N_945,N_213);
and U5159 (N_5159,N_2277,N_2302);
or U5160 (N_5160,N_4740,N_3582);
xor U5161 (N_5161,N_2771,N_2550);
or U5162 (N_5162,N_732,N_939);
nor U5163 (N_5163,N_2512,N_4762);
or U5164 (N_5164,N_3852,N_4621);
nor U5165 (N_5165,N_3160,N_1296);
nand U5166 (N_5166,N_932,N_1960);
nand U5167 (N_5167,N_588,N_1839);
or U5168 (N_5168,N_2133,N_4845);
or U5169 (N_5169,N_3422,N_1913);
xnor U5170 (N_5170,N_4659,N_3398);
xor U5171 (N_5171,N_3203,N_584);
xnor U5172 (N_5172,N_2990,N_508);
nand U5173 (N_5173,N_1610,N_3814);
and U5174 (N_5174,N_755,N_609);
nand U5175 (N_5175,N_4771,N_4028);
and U5176 (N_5176,N_4870,N_4951);
xnor U5177 (N_5177,N_4095,N_763);
nand U5178 (N_5178,N_4744,N_2731);
or U5179 (N_5179,N_2806,N_1972);
nand U5180 (N_5180,N_4960,N_1040);
and U5181 (N_5181,N_1276,N_948);
nor U5182 (N_5182,N_1845,N_1580);
or U5183 (N_5183,N_865,N_2109);
or U5184 (N_5184,N_1996,N_2940);
xor U5185 (N_5185,N_349,N_1194);
nand U5186 (N_5186,N_4398,N_3774);
and U5187 (N_5187,N_1832,N_2031);
nand U5188 (N_5188,N_3230,N_2243);
and U5189 (N_5189,N_1587,N_232);
and U5190 (N_5190,N_1574,N_2315);
or U5191 (N_5191,N_2845,N_3464);
xnor U5192 (N_5192,N_3962,N_577);
xnor U5193 (N_5193,N_2589,N_3099);
and U5194 (N_5194,N_3010,N_2560);
nor U5195 (N_5195,N_4733,N_677);
nand U5196 (N_5196,N_1593,N_2582);
or U5197 (N_5197,N_1929,N_3983);
and U5198 (N_5198,N_4658,N_4780);
nor U5199 (N_5199,N_3888,N_2662);
or U5200 (N_5200,N_1476,N_4153);
nor U5201 (N_5201,N_554,N_2527);
or U5202 (N_5202,N_1660,N_2409);
or U5203 (N_5203,N_2816,N_4664);
and U5204 (N_5204,N_2448,N_3285);
nand U5205 (N_5205,N_3541,N_1393);
nand U5206 (N_5206,N_4167,N_2281);
and U5207 (N_5207,N_4389,N_2337);
nor U5208 (N_5208,N_4527,N_1334);
nand U5209 (N_5209,N_4500,N_4288);
and U5210 (N_5210,N_4433,N_666);
nor U5211 (N_5211,N_4947,N_4089);
and U5212 (N_5212,N_3715,N_4935);
nand U5213 (N_5213,N_317,N_1783);
nand U5214 (N_5214,N_2692,N_4412);
xnor U5215 (N_5215,N_2011,N_2257);
nand U5216 (N_5216,N_2981,N_1299);
and U5217 (N_5217,N_17,N_4021);
and U5218 (N_5218,N_3613,N_4778);
nor U5219 (N_5219,N_2782,N_1038);
nor U5220 (N_5220,N_1046,N_3242);
nor U5221 (N_5221,N_581,N_4916);
nor U5222 (N_5222,N_2200,N_4404);
nand U5223 (N_5223,N_1705,N_1);
xnor U5224 (N_5224,N_1699,N_2846);
xnor U5225 (N_5225,N_3198,N_3626);
or U5226 (N_5226,N_3632,N_1563);
and U5227 (N_5227,N_3266,N_4666);
xor U5228 (N_5228,N_3262,N_2331);
and U5229 (N_5229,N_2856,N_1773);
xnor U5230 (N_5230,N_3644,N_1226);
nand U5231 (N_5231,N_1336,N_1365);
and U5232 (N_5232,N_3815,N_2977);
or U5233 (N_5233,N_439,N_3656);
xor U5234 (N_5234,N_1959,N_2210);
nor U5235 (N_5235,N_370,N_1308);
or U5236 (N_5236,N_4481,N_3920);
nor U5237 (N_5237,N_1126,N_3610);
and U5238 (N_5238,N_2837,N_1949);
nand U5239 (N_5239,N_169,N_3080);
nor U5240 (N_5240,N_4769,N_3146);
nor U5241 (N_5241,N_1965,N_1140);
xnor U5242 (N_5242,N_1506,N_709);
or U5243 (N_5243,N_2893,N_3731);
nand U5244 (N_5244,N_32,N_2607);
nor U5245 (N_5245,N_626,N_981);
or U5246 (N_5246,N_1369,N_3217);
xor U5247 (N_5247,N_91,N_4923);
xnor U5248 (N_5248,N_3592,N_3202);
nand U5249 (N_5249,N_2821,N_201);
xor U5250 (N_5250,N_3561,N_150);
or U5251 (N_5251,N_1612,N_1018);
and U5252 (N_5252,N_2338,N_4461);
or U5253 (N_5253,N_3938,N_2094);
nand U5254 (N_5254,N_3462,N_4753);
xnor U5255 (N_5255,N_1953,N_3087);
xnor U5256 (N_5256,N_1661,N_2367);
nand U5257 (N_5257,N_1690,N_2012);
and U5258 (N_5258,N_1053,N_1331);
nand U5259 (N_5259,N_4297,N_978);
nand U5260 (N_5260,N_2249,N_2457);
and U5261 (N_5261,N_2310,N_4981);
nand U5262 (N_5262,N_2199,N_51);
xnor U5263 (N_5263,N_440,N_260);
nor U5264 (N_5264,N_4948,N_372);
nor U5265 (N_5265,N_521,N_1370);
and U5266 (N_5266,N_4482,N_4302);
and U5267 (N_5267,N_3053,N_846);
and U5268 (N_5268,N_234,N_733);
nand U5269 (N_5269,N_2687,N_2017);
or U5270 (N_5270,N_4293,N_3501);
or U5271 (N_5271,N_2101,N_3848);
nor U5272 (N_5272,N_2062,N_3134);
xnor U5273 (N_5273,N_2141,N_1873);
or U5274 (N_5274,N_929,N_1952);
xnor U5275 (N_5275,N_3782,N_4492);
nand U5276 (N_5276,N_4309,N_3580);
and U5277 (N_5277,N_4961,N_4570);
xor U5278 (N_5278,N_4683,N_899);
or U5279 (N_5279,N_815,N_2374);
nand U5280 (N_5280,N_3678,N_1509);
or U5281 (N_5281,N_1607,N_708);
nor U5282 (N_5282,N_1323,N_3256);
or U5283 (N_5283,N_4316,N_2320);
nand U5284 (N_5284,N_2253,N_4630);
nor U5285 (N_5285,N_444,N_4336);
nand U5286 (N_5286,N_220,N_2610);
nand U5287 (N_5287,N_1758,N_2255);
nand U5288 (N_5288,N_4591,N_4874);
and U5289 (N_5289,N_2000,N_3824);
nand U5290 (N_5290,N_1843,N_571);
xnor U5291 (N_5291,N_3313,N_2478);
nand U5292 (N_5292,N_4005,N_1135);
xor U5293 (N_5293,N_1910,N_2086);
nor U5294 (N_5294,N_4754,N_1766);
nand U5295 (N_5295,N_2352,N_3209);
nand U5296 (N_5296,N_2713,N_1313);
or U5297 (N_5297,N_4525,N_4413);
xnor U5298 (N_5298,N_4092,N_4969);
and U5299 (N_5299,N_3927,N_3059);
and U5300 (N_5300,N_3009,N_3024);
nand U5301 (N_5301,N_2862,N_4377);
xnor U5302 (N_5302,N_1079,N_808);
or U5303 (N_5303,N_4854,N_989);
xor U5304 (N_5304,N_1064,N_849);
and U5305 (N_5305,N_4468,N_2676);
nand U5306 (N_5306,N_2609,N_1677);
xor U5307 (N_5307,N_2154,N_1029);
nand U5308 (N_5308,N_619,N_4308);
xor U5309 (N_5309,N_1381,N_3026);
xor U5310 (N_5310,N_4764,N_2823);
xor U5311 (N_5311,N_4201,N_225);
and U5312 (N_5312,N_3241,N_148);
and U5313 (N_5313,N_4814,N_1961);
or U5314 (N_5314,N_4653,N_4391);
nor U5315 (N_5315,N_3508,N_3532);
nand U5316 (N_5316,N_3420,N_3314);
nand U5317 (N_5317,N_1864,N_3737);
nand U5318 (N_5318,N_2828,N_2817);
nand U5319 (N_5319,N_4171,N_4159);
nor U5320 (N_5320,N_1402,N_696);
nand U5321 (N_5321,N_4575,N_4452);
nand U5322 (N_5322,N_4997,N_4989);
nor U5323 (N_5323,N_1988,N_2882);
nor U5324 (N_5324,N_2150,N_629);
xor U5325 (N_5325,N_2838,N_4919);
and U5326 (N_5326,N_1539,N_2217);
and U5327 (N_5327,N_346,N_4485);
xor U5328 (N_5328,N_3457,N_1479);
xor U5329 (N_5329,N_4865,N_4728);
and U5330 (N_5330,N_1919,N_1582);
or U5331 (N_5331,N_612,N_2158);
nor U5332 (N_5332,N_4817,N_4258);
nor U5333 (N_5333,N_4368,N_4766);
xor U5334 (N_5334,N_1598,N_2330);
nand U5335 (N_5335,N_2791,N_559);
or U5336 (N_5336,N_3341,N_1892);
xor U5337 (N_5337,N_4295,N_1460);
nor U5338 (N_5338,N_4927,N_4498);
nor U5339 (N_5339,N_3460,N_3094);
nor U5340 (N_5340,N_1449,N_3710);
or U5341 (N_5341,N_10,N_3995);
or U5342 (N_5342,N_1317,N_395);
nor U5343 (N_5343,N_2538,N_2124);
nor U5344 (N_5344,N_229,N_2805);
or U5345 (N_5345,N_1557,N_1995);
nand U5346 (N_5346,N_2392,N_746);
nand U5347 (N_5347,N_3681,N_105);
nand U5348 (N_5348,N_1264,N_553);
nor U5349 (N_5349,N_4812,N_3400);
or U5350 (N_5350,N_4765,N_312);
nand U5351 (N_5351,N_530,N_1834);
and U5352 (N_5352,N_1616,N_2088);
xnor U5353 (N_5353,N_207,N_172);
nand U5354 (N_5354,N_1277,N_3144);
nor U5355 (N_5355,N_2997,N_4192);
nor U5356 (N_5356,N_2597,N_480);
nand U5357 (N_5357,N_4912,N_3542);
xor U5358 (N_5358,N_1114,N_3652);
and U5359 (N_5359,N_2226,N_2670);
xnor U5360 (N_5360,N_2811,N_979);
nand U5361 (N_5361,N_3576,N_455);
and U5362 (N_5362,N_2612,N_1147);
and U5363 (N_5363,N_2858,N_4361);
nand U5364 (N_5364,N_2522,N_3821);
nand U5365 (N_5365,N_4042,N_875);
and U5366 (N_5366,N_2216,N_986);
nand U5367 (N_5367,N_4731,N_1472);
and U5368 (N_5368,N_3935,N_3497);
xor U5369 (N_5369,N_4982,N_959);
nand U5370 (N_5370,N_866,N_680);
or U5371 (N_5371,N_2947,N_3868);
nor U5372 (N_5372,N_3150,N_2327);
and U5373 (N_5373,N_2357,N_4576);
xor U5374 (N_5374,N_860,N_843);
nor U5375 (N_5375,N_1981,N_4143);
or U5376 (N_5376,N_2110,N_622);
nor U5377 (N_5377,N_1028,N_3157);
or U5378 (N_5378,N_4987,N_1171);
xor U5379 (N_5379,N_2102,N_143);
and U5380 (N_5380,N_2889,N_2486);
nand U5381 (N_5381,N_1672,N_4424);
nor U5382 (N_5382,N_4941,N_4622);
and U5383 (N_5383,N_4606,N_1831);
xor U5384 (N_5384,N_889,N_2298);
nand U5385 (N_5385,N_2218,N_4553);
or U5386 (N_5386,N_500,N_3065);
or U5387 (N_5387,N_1268,N_1400);
or U5388 (N_5388,N_3212,N_3536);
xor U5389 (N_5389,N_3261,N_3905);
nand U5390 (N_5390,N_1403,N_3609);
xnor U5391 (N_5391,N_3671,N_1714);
or U5392 (N_5392,N_1122,N_1355);
nand U5393 (N_5393,N_185,N_4164);
xnor U5394 (N_5394,N_120,N_2083);
nor U5395 (N_5395,N_358,N_2426);
nand U5396 (N_5396,N_824,N_3620);
nand U5397 (N_5397,N_2312,N_3316);
xnor U5398 (N_5398,N_3655,N_4749);
nand U5399 (N_5399,N_3043,N_1951);
and U5400 (N_5400,N_4090,N_1246);
xnor U5401 (N_5401,N_4035,N_2813);
or U5402 (N_5402,N_2070,N_999);
or U5403 (N_5403,N_58,N_1465);
nand U5404 (N_5404,N_65,N_916);
nand U5405 (N_5405,N_897,N_1247);
and U5406 (N_5406,N_2859,N_4734);
and U5407 (N_5407,N_1139,N_4233);
nor U5408 (N_5408,N_2264,N_2308);
xor U5409 (N_5409,N_1170,N_385);
and U5410 (N_5410,N_1100,N_649);
xnor U5411 (N_5411,N_50,N_4029);
nor U5412 (N_5412,N_906,N_494);
nor U5413 (N_5413,N_499,N_653);
or U5414 (N_5414,N_3993,N_664);
or U5415 (N_5415,N_1665,N_1807);
or U5416 (N_5416,N_4673,N_4458);
nor U5417 (N_5417,N_3357,N_4324);
or U5418 (N_5418,N_4025,N_4601);
xnor U5419 (N_5419,N_3539,N_408);
xnor U5420 (N_5420,N_2008,N_549);
and U5421 (N_5421,N_4956,N_3593);
xor U5422 (N_5422,N_8,N_3697);
or U5423 (N_5423,N_4735,N_3549);
or U5424 (N_5424,N_3552,N_827);
and U5425 (N_5425,N_3818,N_1243);
xnor U5426 (N_5426,N_2116,N_950);
or U5427 (N_5427,N_1964,N_391);
nor U5428 (N_5428,N_1084,N_4599);
xnor U5429 (N_5429,N_4810,N_2405);
nand U5430 (N_5430,N_1611,N_2683);
nand U5431 (N_5431,N_389,N_3598);
xor U5432 (N_5432,N_4643,N_268);
nor U5433 (N_5433,N_3659,N_4745);
or U5434 (N_5434,N_1358,N_124);
nor U5435 (N_5435,N_1659,N_1434);
or U5436 (N_5436,N_748,N_104);
xnor U5437 (N_5437,N_2920,N_687);
nor U5438 (N_5438,N_1433,N_4357);
or U5439 (N_5439,N_651,N_565);
and U5440 (N_5440,N_2096,N_3327);
xnor U5441 (N_5441,N_1821,N_4221);
nand U5442 (N_5442,N_407,N_4739);
xnor U5443 (N_5443,N_1924,N_2784);
nand U5444 (N_5444,N_975,N_2853);
nor U5445 (N_5445,N_3872,N_3222);
nand U5446 (N_5446,N_4414,N_3511);
nand U5447 (N_5447,N_1419,N_1245);
nand U5448 (N_5448,N_4627,N_838);
nor U5449 (N_5449,N_829,N_1475);
nor U5450 (N_5450,N_4118,N_478);
nand U5451 (N_5451,N_4169,N_2299);
or U5452 (N_5452,N_443,N_2792);
or U5453 (N_5453,N_1177,N_2087);
or U5454 (N_5454,N_3566,N_1679);
nor U5455 (N_5455,N_2887,N_3533);
and U5456 (N_5456,N_4847,N_4871);
nor U5457 (N_5457,N_998,N_1511);
and U5458 (N_5458,N_3089,N_712);
nand U5459 (N_5459,N_3559,N_2362);
or U5460 (N_5460,N_2184,N_3925);
nor U5461 (N_5461,N_4930,N_655);
xnor U5462 (N_5462,N_3226,N_3426);
or U5463 (N_5463,N_1605,N_457);
nand U5464 (N_5464,N_3390,N_1366);
nand U5465 (N_5465,N_3132,N_1888);
nand U5466 (N_5466,N_191,N_2913);
nand U5467 (N_5467,N_4439,N_228);
nand U5468 (N_5468,N_955,N_682);
or U5469 (N_5469,N_551,N_2334);
nor U5470 (N_5470,N_4405,N_255);
nor U5471 (N_5471,N_920,N_1716);
or U5472 (N_5472,N_729,N_2556);
and U5473 (N_5473,N_2463,N_4347);
or U5474 (N_5474,N_956,N_2149);
xnor U5475 (N_5475,N_334,N_2473);
and U5476 (N_5476,N_1474,N_2779);
nor U5477 (N_5477,N_4036,N_876);
nor U5478 (N_5478,N_1573,N_1653);
xnor U5479 (N_5479,N_3081,N_1061);
nor U5480 (N_5480,N_1445,N_4061);
nand U5481 (N_5481,N_1999,N_988);
xnor U5482 (N_5482,N_2557,N_2531);
or U5483 (N_5483,N_187,N_1291);
nor U5484 (N_5484,N_4942,N_1836);
and U5485 (N_5485,N_841,N_4729);
nand U5486 (N_5486,N_2063,N_2090);
nor U5487 (N_5487,N_1176,N_821);
nand U5488 (N_5488,N_657,N_4369);
nor U5489 (N_5489,N_4878,N_304);
nor U5490 (N_5490,N_4047,N_679);
nor U5491 (N_5491,N_4348,N_515);
xnor U5492 (N_5492,N_2065,N_243);
xnor U5493 (N_5493,N_4094,N_1376);
xnor U5494 (N_5494,N_1835,N_3329);
nand U5495 (N_5495,N_3076,N_2363);
xor U5496 (N_5496,N_1164,N_2574);
nand U5497 (N_5497,N_3286,N_4589);
nor U5498 (N_5498,N_1380,N_2810);
nor U5499 (N_5499,N_2830,N_1979);
xor U5500 (N_5500,N_4808,N_1145);
or U5501 (N_5501,N_3414,N_2737);
nand U5502 (N_5502,N_1732,N_1601);
or U5503 (N_5503,N_2937,N_753);
nor U5504 (N_5504,N_2107,N_3388);
nand U5505 (N_5505,N_3588,N_3236);
nand U5506 (N_5506,N_3666,N_3964);
or U5507 (N_5507,N_2412,N_2246);
nor U5508 (N_5508,N_3802,N_607);
xor U5509 (N_5509,N_3355,N_2795);
nand U5510 (N_5510,N_1802,N_2559);
xnor U5511 (N_5511,N_2286,N_1671);
or U5512 (N_5512,N_4401,N_3811);
xor U5513 (N_5513,N_4978,N_3748);
nor U5514 (N_5514,N_4128,N_663);
xnor U5515 (N_5515,N_4681,N_2588);
or U5516 (N_5516,N_3419,N_529);
nand U5517 (N_5517,N_3900,N_4018);
nor U5518 (N_5518,N_536,N_3161);
xnor U5519 (N_5519,N_2984,N_2749);
or U5520 (N_5520,N_888,N_4528);
and U5521 (N_5521,N_3686,N_2010);
nor U5522 (N_5522,N_4039,N_2431);
nor U5523 (N_5523,N_486,N_4367);
nand U5524 (N_5524,N_757,N_1352);
or U5525 (N_5525,N_4072,N_1862);
nor U5526 (N_5526,N_2685,N_1956);
nand U5527 (N_5527,N_4826,N_879);
and U5528 (N_5528,N_245,N_2682);
and U5529 (N_5529,N_3958,N_4214);
and U5530 (N_5530,N_4472,N_4396);
or U5531 (N_5531,N_3011,N_1722);
nor U5532 (N_5532,N_1070,N_384);
and U5533 (N_5533,N_2796,N_24);
nor U5534 (N_5534,N_3208,N_2906);
and U5535 (N_5535,N_1958,N_196);
nand U5536 (N_5536,N_701,N_1353);
and U5537 (N_5537,N_1454,N_820);
nand U5538 (N_5538,N_3077,N_3548);
xnor U5539 (N_5539,N_1735,N_3658);
or U5540 (N_5540,N_4125,N_3972);
xnor U5541 (N_5541,N_3362,N_1617);
or U5542 (N_5542,N_1856,N_870);
and U5543 (N_5543,N_807,N_3859);
and U5544 (N_5544,N_2228,N_1980);
nand U5545 (N_5545,N_3614,N_1340);
nand U5546 (N_5546,N_4884,N_1760);
nand U5547 (N_5547,N_3705,N_4238);
or U5548 (N_5548,N_3786,N_2339);
nor U5549 (N_5549,N_995,N_1567);
or U5550 (N_5550,N_637,N_2595);
or U5551 (N_5551,N_2391,N_2929);
xor U5552 (N_5552,N_2122,N_4489);
nand U5553 (N_5553,N_4582,N_1940);
nor U5554 (N_5554,N_2995,N_164);
or U5555 (N_5555,N_2305,N_272);
or U5556 (N_5556,N_4184,N_2476);
and U5557 (N_5557,N_2287,N_2636);
and U5558 (N_5558,N_3219,N_4885);
xor U5559 (N_5559,N_2899,N_4946);
nand U5560 (N_5560,N_20,N_3107);
and U5561 (N_5561,N_4107,N_273);
nand U5562 (N_5562,N_4776,N_3727);
nand U5563 (N_5563,N_991,N_1427);
nand U5564 (N_5564,N_1098,N_3383);
xnor U5565 (N_5565,N_4251,N_335);
or U5566 (N_5566,N_231,N_2839);
and U5567 (N_5567,N_2415,N_738);
nor U5568 (N_5568,N_1943,N_1424);
nor U5569 (N_5569,N_1281,N_1517);
and U5570 (N_5570,N_216,N_3703);
and U5571 (N_5571,N_881,N_4152);
xnor U5572 (N_5572,N_4503,N_1106);
nor U5573 (N_5573,N_3041,N_3675);
nor U5574 (N_5574,N_4949,N_692);
or U5575 (N_5575,N_126,N_3147);
nand U5576 (N_5576,N_2701,N_4286);
and U5577 (N_5577,N_825,N_1751);
and U5578 (N_5578,N_3535,N_1535);
xor U5579 (N_5579,N_2675,N_1450);
nor U5580 (N_5580,N_117,N_3734);
xnor U5581 (N_5581,N_3038,N_2976);
nor U5582 (N_5582,N_4098,N_1397);
nand U5583 (N_5583,N_3936,N_4165);
or U5584 (N_5584,N_2306,N_3127);
nand U5585 (N_5585,N_2949,N_3006);
or U5586 (N_5586,N_3717,N_1710);
and U5587 (N_5587,N_4009,N_2963);
nor U5588 (N_5588,N_3765,N_3827);
nor U5589 (N_5589,N_430,N_2235);
nor U5590 (N_5590,N_4702,N_3429);
xnor U5591 (N_5591,N_47,N_4497);
nor U5592 (N_5592,N_1481,N_678);
and U5593 (N_5593,N_2807,N_947);
nand U5594 (N_5594,N_2074,N_1712);
nand U5595 (N_5595,N_3430,N_3284);
nand U5596 (N_5596,N_832,N_1398);
nor U5597 (N_5597,N_1878,N_558);
nor U5598 (N_5598,N_1666,N_4811);
xor U5599 (N_5599,N_4651,N_3897);
and U5600 (N_5600,N_4253,N_450);
or U5601 (N_5601,N_3917,N_3636);
xnor U5602 (N_5602,N_2414,N_4773);
nand U5603 (N_5603,N_4848,N_424);
or U5604 (N_5604,N_1507,N_902);
and U5605 (N_5605,N_636,N_2454);
or U5606 (N_5606,N_3530,N_2105);
xor U5607 (N_5607,N_14,N_3664);
xnor U5608 (N_5608,N_3417,N_4837);
and U5609 (N_5609,N_4554,N_110);
nor U5610 (N_5610,N_458,N_3154);
xnor U5611 (N_5611,N_2465,N_3869);
nand U5612 (N_5612,N_1939,N_1201);
xor U5613 (N_5613,N_2935,N_71);
and U5614 (N_5614,N_1287,N_2971);
or U5615 (N_5615,N_4971,N_4859);
or U5616 (N_5616,N_1524,N_661);
nor U5617 (N_5617,N_3250,N_3083);
and U5618 (N_5618,N_1008,N_3370);
nand U5619 (N_5619,N_2703,N_4518);
xor U5620 (N_5620,N_2245,N_4567);
or U5621 (N_5621,N_2603,N_1922);
or U5622 (N_5622,N_1795,N_4077);
nor U5623 (N_5623,N_2144,N_3597);
xnor U5624 (N_5624,N_4448,N_894);
nand U5625 (N_5625,N_2179,N_4703);
nor U5626 (N_5626,N_2626,N_1635);
and U5627 (N_5627,N_684,N_4839);
nand U5628 (N_5628,N_421,N_1588);
nand U5629 (N_5629,N_938,N_3415);
and U5630 (N_5630,N_4929,N_2435);
or U5631 (N_5631,N_883,N_4218);
xor U5632 (N_5632,N_1869,N_4717);
or U5633 (N_5633,N_2601,N_2871);
or U5634 (N_5634,N_2369,N_159);
and U5635 (N_5635,N_4852,N_2967);
nand U5636 (N_5636,N_844,N_3331);
nand U5637 (N_5637,N_2034,N_3343);
nor U5638 (N_5638,N_1487,N_1197);
nand U5639 (N_5639,N_4282,N_3528);
and U5640 (N_5640,N_2340,N_394);
nand U5641 (N_5641,N_4071,N_1223);
nand U5642 (N_5642,N_84,N_1991);
and U5643 (N_5643,N_1804,N_1853);
or U5644 (N_5644,N_745,N_4782);
xor U5645 (N_5645,N_1335,N_4894);
nor U5646 (N_5646,N_326,N_354);
xnor U5647 (N_5647,N_4511,N_4767);
xor U5648 (N_5648,N_1575,N_3604);
or U5649 (N_5649,N_3201,N_4085);
nand U5650 (N_5650,N_2525,N_1094);
or U5651 (N_5651,N_3892,N_2767);
nor U5652 (N_5652,N_1657,N_4574);
xnor U5653 (N_5653,N_4170,N_2145);
and U5654 (N_5654,N_2233,N_4318);
and U5655 (N_5655,N_2103,N_598);
nand U5656 (N_5656,N_2602,N_2766);
nor U5657 (N_5657,N_2137,N_1267);
or U5658 (N_5658,N_2790,N_1946);
nand U5659 (N_5659,N_39,N_2238);
nand U5660 (N_5660,N_2986,N_3270);
and U5661 (N_5661,N_2259,N_1590);
nor U5662 (N_5662,N_3992,N_4239);
nand U5663 (N_5663,N_1851,N_315);
or U5664 (N_5664,N_1448,N_1847);
nand U5665 (N_5665,N_1645,N_1036);
or U5666 (N_5666,N_4208,N_3619);
nor U5667 (N_5667,N_4996,N_4605);
nand U5668 (N_5668,N_3591,N_509);
or U5669 (N_5669,N_762,N_4242);
xor U5670 (N_5670,N_463,N_502);
and U5671 (N_5671,N_1883,N_546);
and U5672 (N_5672,N_614,N_4311);
and U5673 (N_5673,N_55,N_4266);
nand U5674 (N_5674,N_2057,N_1801);
nand U5675 (N_5675,N_2366,N_383);
or U5676 (N_5676,N_4720,N_3683);
or U5677 (N_5677,N_4614,N_1962);
and U5678 (N_5678,N_582,N_1974);
nand U5679 (N_5679,N_2523,N_3701);
nor U5680 (N_5680,N_4616,N_872);
or U5681 (N_5681,N_3337,N_3351);
and U5682 (N_5682,N_586,N_3729);
nor U5683 (N_5683,N_4936,N_1254);
nor U5684 (N_5684,N_4339,N_2642);
nand U5685 (N_5685,N_761,N_1520);
or U5686 (N_5686,N_419,N_1295);
nor U5687 (N_5687,N_4342,N_3758);
xor U5688 (N_5688,N_4644,N_4442);
nor U5689 (N_5689,N_3942,N_332);
xor U5690 (N_5690,N_2285,N_2332);
xor U5691 (N_5691,N_974,N_3858);
nand U5692 (N_5692,N_4725,N_3166);
and U5693 (N_5693,N_4066,N_142);
and U5694 (N_5694,N_2777,N_3086);
xor U5695 (N_5695,N_4132,N_3770);
nand U5696 (N_5696,N_2265,N_3131);
nor U5697 (N_5697,N_3386,N_703);
or U5698 (N_5698,N_1280,N_4136);
and U5699 (N_5699,N_2271,N_22);
or U5700 (N_5700,N_2630,N_4112);
and U5701 (N_5701,N_704,N_4395);
and U5702 (N_5702,N_1113,N_941);
or U5703 (N_5703,N_1203,N_4646);
xor U5704 (N_5704,N_4120,N_1150);
xnor U5705 (N_5705,N_767,N_2840);
xnor U5706 (N_5706,N_2278,N_2744);
or U5707 (N_5707,N_3272,N_2176);
nand U5708 (N_5708,N_2621,N_3793);
and U5709 (N_5709,N_1010,N_2725);
and U5710 (N_5710,N_2248,N_4134);
xnor U5711 (N_5711,N_279,N_2798);
nand U5712 (N_5712,N_1576,N_2750);
xnor U5713 (N_5713,N_1222,N_1304);
and U5714 (N_5714,N_4561,N_3634);
nand U5715 (N_5715,N_610,N_3199);
or U5716 (N_5716,N_2117,N_157);
nand U5717 (N_5717,N_3631,N_1768);
xor U5718 (N_5718,N_1111,N_4904);
or U5719 (N_5719,N_2428,N_1187);
and U5720 (N_5720,N_60,N_2521);
or U5721 (N_5721,N_1592,N_1221);
or U5722 (N_5722,N_432,N_3064);
nand U5723 (N_5723,N_4097,N_3228);
xnor U5724 (N_5724,N_2918,N_3565);
nor U5725 (N_5725,N_2741,N_73);
and U5726 (N_5726,N_4900,N_3120);
nor U5727 (N_5727,N_3344,N_683);
nor U5728 (N_5728,N_4447,N_2193);
nor U5729 (N_5729,N_160,N_2652);
or U5730 (N_5730,N_1876,N_2508);
nand U5731 (N_5731,N_4707,N_4150);
or U5732 (N_5732,N_3999,N_2038);
or U5733 (N_5733,N_3629,N_1478);
xor U5734 (N_5734,N_4478,N_3477);
and U5735 (N_5735,N_1004,N_4853);
or U5736 (N_5736,N_1546,N_2273);
and U5737 (N_5737,N_2656,N_3507);
nor U5738 (N_5738,N_2968,N_3036);
or U5739 (N_5739,N_2430,N_3953);
xnor U5740 (N_5740,N_2119,N_2742);
nand U5741 (N_5741,N_3854,N_180);
nand U5742 (N_5742,N_1319,N_1097);
and U5743 (N_5743,N_934,N_915);
nand U5744 (N_5744,N_56,N_3886);
nor U5745 (N_5745,N_4259,N_4873);
xnor U5746 (N_5746,N_4030,N_318);
xnor U5747 (N_5747,N_2211,N_640);
nor U5748 (N_5748,N_993,N_3606);
nor U5749 (N_5749,N_1387,N_3876);
xnor U5750 (N_5750,N_556,N_3449);
and U5751 (N_5751,N_2655,N_1009);
nor U5752 (N_5752,N_3673,N_3142);
and U5753 (N_5753,N_1318,N_2033);
nor U5754 (N_5754,N_2562,N_1747);
nand U5755 (N_5755,N_1662,N_204);
nor U5756 (N_5756,N_2474,N_1915);
or U5757 (N_5757,N_2515,N_1642);
nand U5758 (N_5758,N_2854,N_2025);
or U5759 (N_5759,N_111,N_2698);
nand U5760 (N_5760,N_3487,N_4139);
or U5761 (N_5761,N_4455,N_811);
nand U5762 (N_5762,N_1898,N_1589);
nor U5763 (N_5763,N_833,N_3653);
nand U5764 (N_5764,N_1630,N_1388);
nand U5765 (N_5765,N_461,N_3034);
nor U5766 (N_5766,N_1428,N_3479);
or U5767 (N_5767,N_864,N_2460);
or U5768 (N_5768,N_1500,N_482);
nor U5769 (N_5769,N_2156,N_1109);
nor U5770 (N_5770,N_1480,N_2099);
and U5771 (N_5771,N_2258,N_4538);
nand U5772 (N_5772,N_4833,N_4080);
nand U5773 (N_5773,N_263,N_1648);
and U5774 (N_5774,N_796,N_337);
xnor U5775 (N_5775,N_215,N_1361);
and U5776 (N_5776,N_3349,N_4940);
xnor U5777 (N_5777,N_3495,N_1469);
nand U5778 (N_5778,N_1235,N_1413);
or U5779 (N_5779,N_246,N_1356);
nor U5780 (N_5780,N_2047,N_1193);
xor U5781 (N_5781,N_2307,N_2436);
xnor U5782 (N_5782,N_4270,N_603);
and U5783 (N_5783,N_1547,N_4376);
xnor U5784 (N_5784,N_3267,N_4287);
nand U5785 (N_5785,N_2098,N_3519);
or U5786 (N_5786,N_4243,N_3100);
xor U5787 (N_5787,N_4310,N_3339);
nor U5788 (N_5788,N_76,N_3883);
or U5789 (N_5789,N_660,N_2765);
nand U5790 (N_5790,N_3778,N_1820);
xnor U5791 (N_5791,N_2492,N_2728);
or U5792 (N_5792,N_4199,N_3279);
and U5793 (N_5793,N_96,N_4380);
nand U5794 (N_5794,N_2148,N_903);
nand U5795 (N_5795,N_711,N_2573);
xnor U5796 (N_5796,N_3015,N_1510);
xor U5797 (N_5797,N_4406,N_4354);
nand U5798 (N_5798,N_4116,N_2876);
xor U5799 (N_5799,N_4604,N_4670);
and U5800 (N_5800,N_1259,N_1963);
nand U5801 (N_5801,N_4157,N_1137);
nor U5802 (N_5802,N_1805,N_1884);
xor U5803 (N_5803,N_931,N_248);
and U5804 (N_5804,N_2410,N_672);
and U5805 (N_5805,N_4857,N_3825);
xor U5806 (N_5806,N_2445,N_1623);
nand U5807 (N_5807,N_1297,N_1970);
nand U5808 (N_5808,N_2639,N_3902);
nor U5809 (N_5809,N_1644,N_668);
and U5810 (N_5810,N_1785,N_3171);
and U5811 (N_5811,N_813,N_4319);
nand U5812 (N_5812,N_3306,N_206);
or U5813 (N_5813,N_1416,N_3394);
and U5814 (N_5814,N_303,N_4352);
nand U5815 (N_5815,N_1759,N_4137);
nand U5816 (N_5816,N_2528,N_1872);
xor U5817 (N_5817,N_2472,N_2590);
or U5818 (N_5818,N_1708,N_3584);
xor U5819 (N_5819,N_1942,N_1501);
nor U5820 (N_5820,N_2724,N_4560);
and U5821 (N_5821,N_3694,N_4806);
nand U5822 (N_5822,N_297,N_3097);
and U5823 (N_5823,N_1882,N_628);
nand U5824 (N_5824,N_3165,N_3763);
and U5825 (N_5825,N_1089,N_3360);
and U5826 (N_5826,N_1155,N_4578);
or U5827 (N_5827,N_1282,N_1656);
and U5828 (N_5828,N_971,N_3068);
nand U5829 (N_5829,N_4712,N_2014);
xnor U5830 (N_5830,N_4333,N_3977);
nor U5831 (N_5831,N_4547,N_3986);
nand U5832 (N_5832,N_1930,N_2894);
and U5833 (N_5833,N_877,N_874);
and U5834 (N_5834,N_3742,N_2394);
nor U5835 (N_5835,N_3410,N_3976);
nand U5836 (N_5836,N_1531,N_3571);
nor U5837 (N_5837,N_514,N_1185);
nand U5838 (N_5838,N_1726,N_3882);
or U5839 (N_5839,N_2118,N_2604);
or U5840 (N_5840,N_1600,N_942);
and U5841 (N_5841,N_4609,N_3377);
nand U5842 (N_5842,N_3633,N_1077);
nand U5843 (N_5843,N_3122,N_1065);
and U5844 (N_5844,N_1146,N_4057);
nor U5845 (N_5845,N_97,N_340);
nor U5846 (N_5846,N_3513,N_3159);
nand U5847 (N_5847,N_540,N_2789);
nor U5848 (N_5848,N_2738,N_2873);
nand U5849 (N_5849,N_4684,N_28);
or U5850 (N_5850,N_2907,N_3022);
nor U5851 (N_5851,N_1571,N_2916);
nor U5852 (N_5852,N_4995,N_780);
and U5853 (N_5853,N_2351,N_1700);
or U5854 (N_5854,N_3505,N_3767);
xnor U5855 (N_5855,N_3943,N_2829);
and U5856 (N_5856,N_2309,N_1899);
or U5857 (N_5857,N_4408,N_2938);
and U5858 (N_5858,N_1440,N_36);
or U5859 (N_5859,N_4555,N_511);
nor U5860 (N_5860,N_2157,N_3720);
nor U5861 (N_5861,N_3685,N_3175);
or U5862 (N_5862,N_259,N_2455);
or U5863 (N_5863,N_2501,N_1558);
nand U5864 (N_5864,N_2513,N_4191);
or U5865 (N_5865,N_1810,N_2733);
nand U5866 (N_5866,N_4003,N_1787);
xnor U5867 (N_5867,N_83,N_1136);
nor U5868 (N_5868,N_3870,N_2762);
nand U5869 (N_5869,N_3003,N_1778);
nand U5870 (N_5870,N_4469,N_398);
nor U5871 (N_5871,N_1051,N_4068);
nor U5872 (N_5872,N_2721,N_2664);
and U5873 (N_5873,N_913,N_3416);
or U5874 (N_5874,N_2757,N_1781);
nand U5875 (N_5875,N_737,N_3156);
or U5876 (N_5876,N_2735,N_1652);
xnor U5877 (N_5877,N_522,N_2970);
or U5878 (N_5878,N_3372,N_2071);
or U5879 (N_5879,N_3784,N_4571);
and U5880 (N_5880,N_12,N_3587);
nor U5881 (N_5881,N_2468,N_4235);
and U5882 (N_5882,N_2453,N_4836);
and U5883 (N_5883,N_3243,N_1818);
nor U5884 (N_5884,N_2801,N_1926);
or U5885 (N_5885,N_2543,N_4867);
nand U5886 (N_5886,N_4802,N_922);
or U5887 (N_5887,N_1771,N_3961);
nor U5888 (N_5888,N_4454,N_4907);
and U5889 (N_5889,N_766,N_3929);
nand U5890 (N_5890,N_1684,N_3577);
or U5891 (N_5891,N_2175,N_4194);
nand U5892 (N_5892,N_2181,N_728);
nor U5893 (N_5893,N_2053,N_1932);
and U5894 (N_5894,N_1614,N_1584);
nor U5895 (N_5895,N_3974,N_2776);
nor U5896 (N_5896,N_4325,N_3862);
nor U5897 (N_5897,N_4708,N_518);
or U5898 (N_5898,N_3969,N_1149);
nor U5899 (N_5899,N_2423,N_2406);
or U5900 (N_5900,N_1636,N_2794);
or U5901 (N_5901,N_4789,N_4330);
or U5902 (N_5902,N_4840,N_2021);
and U5903 (N_5903,N_1564,N_3049);
or U5904 (N_5904,N_4831,N_2290);
xor U5905 (N_5905,N_1188,N_784);
nand U5906 (N_5906,N_1152,N_1464);
xnor U5907 (N_5907,N_1189,N_4535);
xnor U5908 (N_5908,N_1125,N_834);
and U5909 (N_5909,N_3326,N_3791);
nor U5910 (N_5910,N_3260,N_3347);
or U5911 (N_5911,N_3137,N_2292);
nor U5912 (N_5912,N_2885,N_698);
or U5913 (N_5913,N_3465,N_3008);
and U5914 (N_5914,N_3585,N_3881);
and U5915 (N_5915,N_2202,N_2780);
xnor U5916 (N_5916,N_3780,N_3278);
nand U5917 (N_5917,N_3062,N_3842);
or U5918 (N_5918,N_1776,N_1875);
and U5919 (N_5919,N_4314,N_4096);
and U5920 (N_5920,N_2985,N_2718);
and U5921 (N_5921,N_1484,N_3789);
and U5922 (N_5922,N_1303,N_3702);
nand U5923 (N_5923,N_2404,N_348);
or U5924 (N_5924,N_310,N_4111);
or U5925 (N_5925,N_4679,N_1368);
or U5926 (N_5926,N_1687,N_1997);
xnor U5927 (N_5927,N_266,N_1158);
xnor U5928 (N_5928,N_779,N_1841);
or U5929 (N_5929,N_4937,N_2570);
or U5930 (N_5930,N_926,N_3225);
xnor U5931 (N_5931,N_1311,N_3557);
and U5932 (N_5932,N_3247,N_4862);
xor U5933 (N_5933,N_4667,N_2244);
or U5934 (N_5934,N_773,N_882);
xor U5935 (N_5935,N_1060,N_2126);
nor U5936 (N_5936,N_525,N_2230);
or U5937 (N_5937,N_996,N_4899);
nand U5938 (N_5938,N_2284,N_4642);
nand U5939 (N_5939,N_3695,N_30);
xor U5940 (N_5940,N_448,N_1129);
xor U5941 (N_5941,N_3813,N_3288);
xnor U5942 (N_5942,N_2370,N_2842);
xor U5943 (N_5943,N_1249,N_654);
and U5944 (N_5944,N_3829,N_3605);
nor U5945 (N_5945,N_836,N_727);
or U5946 (N_5946,N_4743,N_1024);
nor U5947 (N_5947,N_3612,N_4154);
nor U5948 (N_5948,N_78,N_48);
nand U5949 (N_5949,N_2164,N_754);
nor U5950 (N_5950,N_1497,N_4231);
or U5951 (N_5951,N_2177,N_910);
nor U5952 (N_5952,N_542,N_1774);
nor U5953 (N_5953,N_4761,N_1733);
xor U5954 (N_5954,N_770,N_3046);
nand U5955 (N_5955,N_689,N_1389);
or U5956 (N_5956,N_4280,N_4422);
nor U5957 (N_5957,N_896,N_1502);
or U5958 (N_5958,N_880,N_3832);
and U5959 (N_5959,N_1707,N_4590);
xnor U5960 (N_5960,N_601,N_1483);
xnor U5961 (N_5961,N_791,N_479);
and U5962 (N_5962,N_3020,N_4868);
and U5963 (N_5963,N_4151,N_1780);
nand U5964 (N_5964,N_3103,N_426);
nor U5965 (N_5965,N_95,N_3406);
xor U5966 (N_5966,N_1486,N_4842);
xnor U5967 (N_5967,N_3259,N_2833);
and U5968 (N_5968,N_3353,N_1225);
or U5969 (N_5969,N_4901,N_751);
xor U5970 (N_5970,N_794,N_1941);
xnor U5971 (N_5971,N_4174,N_3589);
nor U5972 (N_5972,N_2196,N_2549);
nand U5973 (N_5973,N_1969,N_2143);
or U5974 (N_5974,N_307,N_3129);
nor U5975 (N_5975,N_4690,N_3376);
nand U5976 (N_5976,N_4705,N_371);
xnor U5977 (N_5977,N_1174,N_309);
or U5978 (N_5978,N_4048,N_2568);
nand U5979 (N_5979,N_919,N_2171);
xnor U5980 (N_5980,N_1741,N_1689);
nand U5981 (N_5981,N_3990,N_1013);
or U5982 (N_5982,N_2055,N_133);
nor U5983 (N_5983,N_599,N_1947);
and U5984 (N_5984,N_1639,N_2524);
nand U5985 (N_5985,N_1374,N_1817);
nor U5986 (N_5986,N_2710,N_156);
nand U5987 (N_5987,N_428,N_2611);
and U5988 (N_5988,N_2540,N_66);
nand U5989 (N_5989,N_3244,N_4119);
or U5990 (N_5990,N_1242,N_2872);
xor U5991 (N_5991,N_2398,N_3847);
nand U5992 (N_5992,N_122,N_53);
and U5993 (N_5993,N_3276,N_1470);
nand U5994 (N_5994,N_2542,N_552);
or U5995 (N_5995,N_1633,N_70);
xnor U5996 (N_5996,N_3173,N_2250);
or U5997 (N_5997,N_3670,N_3624);
or U5998 (N_5998,N_4687,N_2809);
nand U5999 (N_5999,N_4480,N_2295);
and U6000 (N_6000,N_3445,N_2417);
and U6001 (N_6001,N_412,N_107);
and U6002 (N_6002,N_2446,N_734);
nor U6003 (N_6003,N_1027,N_1599);
nand U6004 (N_6004,N_3485,N_3512);
and U6005 (N_6005,N_295,N_4440);
nand U6006 (N_6006,N_3567,N_3603);
or U6007 (N_6007,N_1161,N_758);
xnor U6008 (N_6008,N_1239,N_4602);
or U6009 (N_6009,N_3939,N_339);
nand U6010 (N_6010,N_2705,N_2022);
nor U6011 (N_6011,N_1828,N_3650);
nor U6012 (N_6012,N_731,N_1534);
nand U6013 (N_6013,N_3,N_241);
nor U6014 (N_6014,N_1762,N_9);
xor U6015 (N_6015,N_4278,N_5);
xnor U6016 (N_6016,N_4986,N_3894);
xor U6017 (N_6017,N_1180,N_1076);
or U6018 (N_6018,N_2998,N_4943);
and U6019 (N_6019,N_405,N_2641);
xnor U6020 (N_6020,N_4880,N_2673);
xnor U6021 (N_6021,N_1315,N_3317);
or U6022 (N_6022,N_3525,N_3361);
nor U6023 (N_6023,N_2030,N_760);
xor U6024 (N_6024,N_3073,N_1702);
nor U6025 (N_6025,N_3984,N_853);
xnor U6026 (N_6026,N_4384,N_1263);
or U6027 (N_6027,N_178,N_3845);
and U6028 (N_6028,N_3039,N_2665);
nand U6029 (N_6029,N_103,N_3251);
xor U6030 (N_6030,N_4285,N_4962);
xor U6031 (N_6031,N_1504,N_4715);
or U6032 (N_6032,N_928,N_396);
and U6033 (N_6033,N_1069,N_3423);
nor U6034 (N_6034,N_4109,N_4268);
and U6035 (N_6035,N_699,N_1439);
nand U6036 (N_6036,N_4411,N_2620);
nand U6037 (N_6037,N_1905,N_1627);
or U6038 (N_6038,N_21,N_4598);
xnor U6039 (N_6039,N_1968,N_2660);
nor U6040 (N_6040,N_3674,N_2263);
xor U6041 (N_6041,N_2711,N_641);
xor U6042 (N_6042,N_2232,N_776);
or U6043 (N_6043,N_2925,N_4891);
nor U6044 (N_6044,N_3452,N_3776);
or U6045 (N_6045,N_4523,N_3941);
and U6046 (N_6046,N_341,N_214);
nand U6047 (N_6047,N_4301,N_3325);
or U6048 (N_6048,N_3569,N_2153);
or U6049 (N_6049,N_4124,N_2719);
and U6050 (N_6050,N_2974,N_1717);
and U6051 (N_6051,N_2411,N_503);
nand U6052 (N_6052,N_3551,N_2318);
and U6053 (N_6053,N_1157,N_1544);
nand U6054 (N_6054,N_2945,N_4678);
xnor U6055 (N_6055,N_4133,N_908);
nor U6056 (N_6056,N_3113,N_4710);
nor U6057 (N_6057,N_4835,N_1704);
nor U6058 (N_6058,N_2624,N_854);
nand U6059 (N_6059,N_2895,N_3299);
nor U6060 (N_6060,N_2499,N_2923);
nand U6061 (N_6061,N_1692,N_3965);
or U6062 (N_6062,N_4313,N_35);
or U6063 (N_6063,N_1016,N_4600);
nand U6064 (N_6064,N_3745,N_1337);
nor U6065 (N_6065,N_2910,N_4772);
nand U6066 (N_6066,N_2419,N_1071);
and U6067 (N_6067,N_4450,N_3408);
or U6068 (N_6068,N_3274,N_749);
or U6069 (N_6069,N_1333,N_2395);
or U6070 (N_6070,N_534,N_1789);
xor U6071 (N_6071,N_2763,N_4476);
or U6072 (N_6072,N_1550,N_1007);
nand U6073 (N_6073,N_3047,N_4719);
and U6074 (N_6074,N_476,N_2695);
or U6075 (N_6075,N_968,N_2294);
nand U6076 (N_6076,N_4758,N_1591);
nand U6077 (N_6077,N_3169,N_2581);
or U6078 (N_6078,N_261,N_3516);
xnor U6079 (N_6079,N_1819,N_3538);
xnor U6080 (N_6080,N_4718,N_1798);
and U6081 (N_6081,N_1463,N_1830);
xnor U6082 (N_6082,N_4787,N_4586);
and U6083 (N_6083,N_275,N_400);
nor U6084 (N_6084,N_723,N_4950);
and U6085 (N_6085,N_3139,N_1435);
or U6086 (N_6086,N_2891,N_3194);
nand U6087 (N_6087,N_416,N_2355);
nand U6088 (N_6088,N_244,N_2155);
and U6089 (N_6089,N_3002,N_1492);
nand U6090 (N_6090,N_1846,N_3928);
nor U6091 (N_6091,N_2697,N_1925);
nand U6092 (N_6092,N_4307,N_3707);
and U6093 (N_6093,N_1718,N_3724);
and U6094 (N_6094,N_437,N_2954);
or U6095 (N_6095,N_4537,N_365);
nor U6096 (N_6096,N_1746,N_862);
and U6097 (N_6097,N_752,N_4618);
nor U6098 (N_6098,N_177,N_4552);
nand U6099 (N_6099,N_2194,N_4350);
nand U6100 (N_6100,N_4846,N_1425);
nand U6101 (N_6101,N_281,N_1694);
nand U6102 (N_6102,N_953,N_4403);
xnor U6103 (N_6103,N_2347,N_591);
or U6104 (N_6104,N_1737,N_4843);
nand U6105 (N_6105,N_3145,N_4637);
or U6106 (N_6106,N_1540,N_2932);
and U6107 (N_6107,N_611,N_1667);
and U6108 (N_6108,N_1285,N_1686);
and U6109 (N_6109,N_3031,N_3451);
xor U6110 (N_6110,N_2159,N_3718);
or U6111 (N_6111,N_1647,N_4775);
and U6112 (N_6112,N_2586,N_2911);
and U6113 (N_6113,N_4431,N_2848);
xor U6114 (N_6114,N_1537,N_4540);
and U6115 (N_6115,N_606,N_4198);
nand U6116 (N_6116,N_3980,N_2672);
or U6117 (N_6117,N_2615,N_3182);
and U6118 (N_6118,N_4329,N_2503);
or U6119 (N_6119,N_4514,N_1754);
nand U6120 (N_6120,N_3545,N_2333);
nand U6121 (N_6121,N_3296,N_2403);
and U6122 (N_6122,N_2048,N_676);
nand U6123 (N_6123,N_819,N_2052);
or U6124 (N_6124,N_4539,N_504);
nand U6125 (N_6125,N_633,N_2469);
and U6126 (N_6126,N_3215,N_2361);
nor U6127 (N_6127,N_857,N_1378);
xnor U6128 (N_6128,N_193,N_4114);
nand U6129 (N_6129,N_4631,N_3434);
xnor U6130 (N_6130,N_4711,N_3085);
nor U6131 (N_6131,N_4327,N_3879);
and U6132 (N_6132,N_4248,N_1326);
or U6133 (N_6133,N_3621,N_951);
and U6134 (N_6134,N_4784,N_2489);
nor U6135 (N_6135,N_774,N_1058);
nor U6136 (N_6136,N_3798,N_961);
or U6137 (N_6137,N_3615,N_4828);
nor U6138 (N_6138,N_700,N_2897);
nand U6139 (N_6139,N_3224,N_182);
and U6140 (N_6140,N_293,N_3427);
or U6141 (N_6141,N_1401,N_257);
nand U6142 (N_6142,N_3891,N_4402);
or U6143 (N_6143,N_3856,N_3264);
nand U6144 (N_6144,N_4058,N_265);
nand U6145 (N_6145,N_2554,N_4967);
nand U6146 (N_6146,N_4062,N_2722);
nand U6147 (N_6147,N_4041,N_1075);
xor U6148 (N_6148,N_1799,N_4382);
xnor U6149 (N_6149,N_740,N_1021);
nor U6150 (N_6150,N_81,N_1971);
xnor U6151 (N_6151,N_2168,N_4562);
and U6152 (N_6152,N_4038,N_2480);
nor U6153 (N_6153,N_4855,N_4756);
nand U6154 (N_6154,N_2802,N_217);
or U6155 (N_6155,N_1377,N_4633);
nor U6156 (N_6156,N_3779,N_4024);
nand U6157 (N_6157,N_3484,N_2);
and U6158 (N_6158,N_1202,N_2300);
or U6159 (N_6159,N_624,N_804);
nor U6160 (N_6160,N_3304,N_1057);
xor U6161 (N_6161,N_2464,N_1998);
nand U6162 (N_6162,N_287,N_2585);
xnor U6163 (N_6163,N_3425,N_2924);
nand U6164 (N_6164,N_4277,N_3437);
and U6165 (N_6165,N_4043,N_1458);
and U6166 (N_6166,N_4959,N_2835);
or U6167 (N_6167,N_2678,N_625);
nor U6168 (N_6168,N_1966,N_2965);
nor U6169 (N_6169,N_3321,N_1142);
nor U6170 (N_6170,N_2407,N_3502);
or U6171 (N_6171,N_2946,N_4611);
nand U6172 (N_6172,N_2658,N_4519);
nor U6173 (N_6173,N_3750,N_4569);
nor U6174 (N_6174,N_151,N_1039);
xnor U6175 (N_6175,N_1585,N_573);
and U6176 (N_6176,N_3949,N_718);
nand U6177 (N_6177,N_4662,N_4181);
or U6178 (N_6178,N_4122,N_459);
xnor U6179 (N_6179,N_3772,N_2726);
or U6180 (N_6180,N_532,N_1430);
nor U6181 (N_6181,N_2461,N_1945);
nor U6182 (N_6182,N_308,N_3809);
or U6183 (N_6183,N_1901,N_4457);
nor U6184 (N_6184,N_3359,N_99);
or U6185 (N_6185,N_4695,N_4187);
or U6186 (N_6186,N_3997,N_2020);
nor U6187 (N_6187,N_4957,N_3573);
and U6188 (N_6188,N_1286,N_3265);
or U6189 (N_6189,N_2834,N_3922);
nand U6190 (N_6190,N_2494,N_946);
or U6191 (N_6191,N_2353,N_453);
nand U6192 (N_6192,N_686,N_1553);
and U6193 (N_6193,N_1603,N_1861);
nand U6194 (N_6194,N_4883,N_596);
nand U6195 (N_6195,N_667,N_4721);
xor U6196 (N_6196,N_4732,N_901);
and U6197 (N_6197,N_2376,N_2402);
xnor U6198 (N_6198,N_2545,N_593);
and U6199 (N_6199,N_4760,N_314);
and U6200 (N_6200,N_2594,N_2686);
xnor U6201 (N_6201,N_2962,N_1081);
or U6202 (N_6202,N_175,N_4227);
or U6203 (N_6203,N_1086,N_2739);
xnor U6204 (N_6204,N_1493,N_561);
xor U6205 (N_6205,N_4475,N_4359);
nand U6206 (N_6206,N_4044,N_3504);
or U6207 (N_6207,N_713,N_2272);
xnor U6208 (N_6208,N_4232,N_3910);
and U6209 (N_6209,N_2066,N_4341);
and U6210 (N_6210,N_4383,N_4786);
nand U6211 (N_6211,N_2926,N_3968);
xor U6212 (N_6212,N_4700,N_87);
xnor U6213 (N_6213,N_3810,N_4663);
and U6214 (N_6214,N_3688,N_4668);
nor U6215 (N_6215,N_2747,N_374);
or U6216 (N_6216,N_3543,N_579);
and U6217 (N_6217,N_327,N_2653);
or U6218 (N_6218,N_4054,N_288);
xnor U6219 (N_6219,N_1023,N_1406);
or U6220 (N_6220,N_4530,N_3849);
nand U6221 (N_6221,N_4254,N_2892);
or U6222 (N_6222,N_4105,N_112);
xnor U6223 (N_6223,N_4289,N_2843);
and U6224 (N_6224,N_1068,N_230);
nor U6225 (N_6225,N_4102,N_3393);
xnor U6226 (N_6226,N_390,N_1169);
and U6227 (N_6227,N_2467,N_1871);
nand U6228 (N_6228,N_147,N_324);
nor U6229 (N_6229,N_4496,N_2026);
or U6230 (N_6230,N_4777,N_4636);
and U6231 (N_6231,N_74,N_299);
nor U6232 (N_6232,N_3560,N_4958);
and U6233 (N_6233,N_4619,N_1628);
nand U6234 (N_6234,N_1118,N_4677);
and U6235 (N_6235,N_2668,N_1417);
and U6236 (N_6236,N_3755,N_1148);
nor U6237 (N_6237,N_3118,N_595);
and U6238 (N_6238,N_2343,N_271);
and U6239 (N_6239,N_3106,N_57);
and U6240 (N_6240,N_4362,N_4017);
nand U6241 (N_6241,N_969,N_269);
xnor U6242 (N_6242,N_2166,N_1489);
xnor U6243 (N_6243,N_2296,N_3352);
and U6244 (N_6244,N_171,N_2770);
and U6245 (N_6245,N_4346,N_3751);
nor U6246 (N_6246,N_1880,N_3473);
xor U6247 (N_6247,N_3816,N_4464);
or U6248 (N_6248,N_3155,N_3957);
nor U6249 (N_6249,N_4551,N_4399);
and U6250 (N_6250,N_4219,N_2511);
xnor U6251 (N_6251,N_2680,N_2064);
and U6252 (N_6252,N_3662,N_2016);
nand U6253 (N_6253,N_52,N_1192);
nor U6254 (N_6254,N_4381,N_1011);
nand U6255 (N_6255,N_1328,N_3676);
xor U6256 (N_6256,N_1626,N_2089);
or U6257 (N_6257,N_524,N_1538);
or U6258 (N_6258,N_3181,N_4816);
or U6259 (N_6259,N_1850,N_527);
xnor U6260 (N_6260,N_1459,N_1703);
nand U6261 (N_6261,N_2208,N_1372);
and U6262 (N_6262,N_3063,N_181);
or U6263 (N_6263,N_174,N_85);
and U6264 (N_6264,N_1396,N_1518);
nor U6265 (N_6265,N_936,N_4645);
nand U6266 (N_6266,N_772,N_1638);
and U6267 (N_6267,N_3152,N_1275);
or U6268 (N_6268,N_4487,N_270);
and U6269 (N_6269,N_2884,N_4423);
xnor U6270 (N_6270,N_4699,N_254);
or U6271 (N_6271,N_1214,N_3117);
nand U6272 (N_6272,N_3153,N_2378);
and U6273 (N_6273,N_1273,N_1272);
or U6274 (N_6274,N_742,N_1618);
or U6275 (N_6275,N_1503,N_1914);
nor U6276 (N_6276,N_4737,N_775);
nand U6277 (N_6277,N_101,N_4443);
and U6278 (N_6278,N_4064,N_4742);
xor U6279 (N_6279,N_3395,N_839);
and U6280 (N_6280,N_125,N_4006);
nand U6281 (N_6281,N_1891,N_2704);
or U6282 (N_6282,N_2879,N_3471);
nand U6283 (N_6283,N_992,N_2651);
and U6284 (N_6284,N_1213,N_4007);
xnor U6285 (N_6285,N_1513,N_4888);
nor U6286 (N_6286,N_1902,N_3544);
or U6287 (N_6287,N_4397,N_2818);
or U6288 (N_6288,N_2039,N_4015);
and U6289 (N_6289,N_3435,N_294);
nand U6290 (N_6290,N_369,N_2625);
nand U6291 (N_6291,N_1854,N_285);
nor U6292 (N_6292,N_852,N_1399);
xnor U6293 (N_6293,N_2239,N_1634);
xnor U6294 (N_6294,N_3524,N_4955);
nand U6295 (N_6295,N_4303,N_4660);
or U6296 (N_6296,N_4887,N_4490);
xnor U6297 (N_6297,N_3453,N_4000);
nand U6298 (N_6298,N_3923,N_4257);
xnor U6299 (N_6299,N_2487,N_3210);
xor U6300 (N_6300,N_3389,N_3496);
or U6301 (N_6301,N_4909,N_2262);
nor U6302 (N_6302,N_4215,N_809);
xnor U6303 (N_6303,N_2078,N_59);
nand U6304 (N_6304,N_4549,N_2730);
or U6305 (N_6305,N_3269,N_1383);
nand U6306 (N_6306,N_441,N_2988);
xnor U6307 (N_6307,N_4759,N_2994);
or U6308 (N_6308,N_1436,N_4056);
xnor U6309 (N_6309,N_3878,N_2169);
or U6310 (N_6310,N_1054,N_2241);
nor U6311 (N_6311,N_203,N_4985);
nand U6312 (N_6312,N_1438,N_3190);
xor U6313 (N_6313,N_604,N_4603);
nor U6314 (N_6314,N_1983,N_2349);
xnor U6315 (N_6315,N_1033,N_4895);
and U6316 (N_6316,N_1527,N_302);
xnor U6317 (N_6317,N_3088,N_4474);
and U6318 (N_6318,N_1123,N_1530);
xor U6319 (N_6319,N_1826,N_1554);
nand U6320 (N_6320,N_3292,N_423);
nand U6321 (N_6321,N_2424,N_1107);
xnor U6322 (N_6322,N_2130,N_1047);
nor U6323 (N_6323,N_3301,N_2934);
xor U6324 (N_6324,N_2861,N_2616);
and U6325 (N_6325,N_4331,N_2234);
or U6326 (N_6326,N_4881,N_4245);
or U6327 (N_6327,N_994,N_134);
nor U6328 (N_6328,N_3149,N_4429);
or U6329 (N_6329,N_1091,N_2803);
or U6330 (N_6330,N_856,N_2958);
nor U6331 (N_6331,N_3239,N_3564);
and U6332 (N_6332,N_4724,N_2051);
xor U6333 (N_6333,N_2080,N_152);
or U6334 (N_6334,N_2565,N_4750);
nand U6335 (N_6335,N_442,N_1228);
nand U6336 (N_6336,N_2267,N_362);
nor U6337 (N_6337,N_3109,N_1052);
nand U6338 (N_6338,N_1840,N_954);
nand U6339 (N_6339,N_1491,N_397);
nor U6340 (N_6340,N_4332,N_2497);
nand U6341 (N_6341,N_3442,N_3071);
nor U6342 (N_6342,N_2079,N_1108);
nand U6343 (N_6343,N_2375,N_778);
or U6344 (N_6344,N_3796,N_1752);
nand U6345 (N_6345,N_3379,N_3204);
and U6346 (N_6346,N_2212,N_3853);
or U6347 (N_6347,N_1394,N_4755);
xor U6348 (N_6348,N_1731,N_218);
nand U6349 (N_6349,N_3654,N_1893);
nand U6350 (N_6350,N_1175,N_726);
nand U6351 (N_6351,N_2688,N_2580);
and U6352 (N_6352,N_4022,N_179);
nor U6353 (N_6353,N_4910,N_645);
or U6354 (N_6354,N_3277,N_2219);
xnor U6355 (N_6355,N_3336,N_2152);
and U6356 (N_6356,N_3617,N_1128);
nor U6357 (N_6357,N_3421,N_2969);
or U6358 (N_6358,N_4141,N_2440);
and U6359 (N_6359,N_782,N_2785);
or U6360 (N_6360,N_1842,N_1812);
nand U6361 (N_6361,N_3017,N_1332);
xor U6362 (N_6362,N_4903,N_2714);
xor U6363 (N_6363,N_2637,N_108);
xor U6364 (N_6364,N_3407,N_1837);
nor U6365 (N_6365,N_858,N_2579);
and U6366 (N_6366,N_4189,N_406);
nor U6367 (N_6367,N_1736,N_2915);
and U6368 (N_6368,N_3091,N_4113);
nand U6369 (N_6369,N_3411,N_3828);
or U6370 (N_6370,N_3646,N_925);
xor U6371 (N_6371,N_2354,N_2666);
and U6372 (N_6372,N_2418,N_4059);
nand U6373 (N_6373,N_1711,N_3563);
xor U6374 (N_6374,N_4086,N_2874);
nand U6375 (N_6375,N_3562,N_1412);
and U6376 (N_6376,N_1063,N_638);
xor U6377 (N_6377,N_1165,N_4441);
nor U6378 (N_6378,N_2447,N_4876);
xor U6379 (N_6379,N_1230,N_1043);
or U6380 (N_6380,N_4312,N_741);
or U6381 (N_6381,N_319,N_4417);
nand U6382 (N_6382,N_1030,N_4512);
xor U6383 (N_6383,N_2470,N_2510);
nand U6384 (N_6384,N_356,N_1682);
nand U6385 (N_6385,N_3164,N_789);
or U6386 (N_6386,N_4353,N_274);
and U6387 (N_6387,N_2112,N_4291);
and U6388 (N_6388,N_2768,N_2254);
nand U6389 (N_6389,N_4436,N_949);
xor U6390 (N_6390,N_4748,N_506);
nor U6391 (N_6391,N_1124,N_2778);
or U6392 (N_6392,N_800,N_1104);
nor U6393 (N_6393,N_1022,N_2622);
xnor U6394 (N_6394,N_1265,N_2684);
nand U6395 (N_6395,N_960,N_1849);
nor U6396 (N_6396,N_691,N_4998);
nor U6397 (N_6397,N_1112,N_647);
xnor U6398 (N_6398,N_1103,N_2304);
nand U6399 (N_6399,N_884,N_4121);
nor U6400 (N_6400,N_1669,N_4938);
nand U6401 (N_6401,N_3315,N_4696);
xor U6402 (N_6402,N_3193,N_1248);
xor U6403 (N_6403,N_1823,N_121);
xor U6404 (N_6404,N_4509,N_3752);
nand U6405 (N_6405,N_1443,N_850);
nand U6406 (N_6406,N_4173,N_42);
nand U6407 (N_6407,N_513,N_2227);
xnor U6408 (N_6408,N_3500,N_744);
nor U6409 (N_6409,N_3013,N_2433);
nand U6410 (N_6410,N_3987,N_3590);
nor U6411 (N_6411,N_1917,N_3310);
xnor U6412 (N_6412,N_3258,N_648);
and U6413 (N_6413,N_1138,N_4803);
nand U6414 (N_6414,N_4010,N_267);
and U6415 (N_6415,N_3237,N_2037);
xor U6416 (N_6416,N_1764,N_4693);
or U6417 (N_6417,N_1080,N_190);
nand U6418 (N_6418,N_1067,N_3332);
nor U6419 (N_6419,N_3540,N_2775);
nand U6420 (N_6420,N_3616,N_2886);
xnor U6421 (N_6421,N_1360,N_4914);
xor U6422 (N_6422,N_3635,N_1879);
or U6423 (N_6423,N_4045,N_1739);
xnor U6424 (N_6424,N_4568,N_0);
and U6425 (N_6425,N_2056,N_4588);
and U6426 (N_6426,N_399,N_952);
xnor U6427 (N_6427,N_1110,N_4800);
nor U6428 (N_6428,N_1698,N_1559);
xnor U6429 (N_6429,N_4493,N_997);
xnor U6430 (N_6430,N_3871,N_3140);
nor U6431 (N_6431,N_2880,N_3023);
nor U6432 (N_6432,N_3254,N_1364);
nor U6433 (N_6433,N_79,N_878);
or U6434 (N_6434,N_4520,N_4178);
nor U6435 (N_6435,N_2632,N_2979);
nor U6436 (N_6436,N_4544,N_1482);
and U6437 (N_6437,N_3839,N_4008);
and U6438 (N_6438,N_3079,N_4548);
nor U6439 (N_6439,N_188,N_2944);
nor U6440 (N_6440,N_495,N_1791);
or U6441 (N_6441,N_3728,N_1090);
and U6442 (N_6442,N_136,N_1579);
nor U6443 (N_6443,N_2650,N_2788);
nor U6444 (N_6444,N_1032,N_2452);
nor U6445 (N_6445,N_3509,N_4524);
nand U6446 (N_6446,N_3640,N_3104);
nor U6447 (N_6447,N_2170,N_2558);
and U6448 (N_6448,N_4533,N_4558);
and U6449 (N_6449,N_3861,N_1813);
xnor U6450 (N_6450,N_2890,N_2506);
and U6451 (N_6451,N_1865,N_4016);
nand U6452 (N_6452,N_3553,N_4805);
nor U6453 (N_6453,N_4415,N_2696);
nor U6454 (N_6454,N_2820,N_2577);
nor U6455 (N_6455,N_2439,N_756);
or U6456 (N_6456,N_3812,N_3240);
or U6457 (N_6457,N_2204,N_3446);
nand U6458 (N_6458,N_82,N_1327);
and U6459 (N_6459,N_2706,N_1994);
and U6460 (N_6460,N_3384,N_4049);
and U6461 (N_6461,N_119,N_100);
and U6462 (N_6462,N_3554,N_1806);
nand U6463 (N_6463,N_381,N_3280);
or U6464 (N_6464,N_671,N_1723);
and U6465 (N_6465,N_4115,N_2634);
nor U6466 (N_6466,N_1279,N_4751);
or U6467 (N_6467,N_3918,N_585);
nand U6468 (N_6468,N_313,N_1498);
xor U6469 (N_6469,N_4222,N_1144);
nand U6470 (N_6470,N_4241,N_2192);
and U6471 (N_6471,N_985,N_4212);
xnor U6472 (N_6472,N_3608,N_4752);
nor U6473 (N_6473,N_2186,N_2814);
and U6474 (N_6474,N_1793,N_1858);
nand U6475 (N_6475,N_1455,N_1715);
nor U6476 (N_6476,N_129,N_3637);
nor U6477 (N_6477,N_517,N_2291);
nor U6478 (N_6478,N_3790,N_4033);
and U6479 (N_6479,N_2755,N_2760);
or U6480 (N_6480,N_1742,N_4410);
or U6481 (N_6481,N_1191,N_277);
nor U6482 (N_6482,N_2180,N_3985);
nor U6483 (N_6483,N_4140,N_1838);
or U6484 (N_6484,N_2280,N_1683);
and U6485 (N_6485,N_1986,N_2567);
or U6486 (N_6486,N_325,N_3148);
xnor U6487 (N_6487,N_2787,N_608);
xor U6488 (N_6488,N_4990,N_1643);
xor U6489 (N_6489,N_600,N_543);
nor U6490 (N_6490,N_574,N_4704);
or U6491 (N_6491,N_886,N_2434);
nand U6492 (N_6492,N_3115,N_2209);
or U6493 (N_6493,N_3367,N_4304);
or U6494 (N_6494,N_2504,N_116);
or U6495 (N_6495,N_3108,N_1923);
and U6496 (N_6496,N_2146,N_377);
or U6497 (N_6497,N_675,N_4692);
nand U6498 (N_6498,N_2371,N_3238);
nor U6499 (N_6499,N_2799,N_1325);
and U6500 (N_6500,N_320,N_3069);
and U6501 (N_6501,N_3399,N_1822);
or U6502 (N_6502,N_4073,N_1728);
or U6503 (N_6503,N_417,N_2383);
nand U6504 (N_6504,N_4161,N_2812);
or U6505 (N_6505,N_4879,N_4205);
nor U6506 (N_6506,N_235,N_898);
xor U6507 (N_6507,N_2999,N_803);
nor U6508 (N_6508,N_3322,N_4963);
xor U6509 (N_6509,N_924,N_3510);
and U6510 (N_6510,N_1407,N_3170);
nor U6511 (N_6511,N_2681,N_2329);
xnor U6512 (N_6512,N_330,N_4050);
xnor U6513 (N_6513,N_145,N_2623);
nand U6514 (N_6514,N_3136,N_2268);
nor U6515 (N_6515,N_4437,N_2841);
and U6516 (N_6516,N_3391,N_77);
nand U6517 (N_6517,N_2720,N_1035);
and U6518 (N_6518,N_674,N_2247);
xnor U6519 (N_6519,N_4841,N_3402);
xor U6520 (N_6520,N_1989,N_1641);
or U6521 (N_6521,N_4499,N_2127);
xnor U6522 (N_6522,N_1827,N_2993);
or U6523 (N_6523,N_1251,N_990);
nor U6524 (N_6524,N_3116,N_2282);
xor U6525 (N_6525,N_4246,N_292);
or U6526 (N_6526,N_3788,N_382);
nand U6527 (N_6527,N_4334,N_545);
and U6528 (N_6528,N_2518,N_1116);
nand U6529 (N_6529,N_1649,N_2225);
and U6530 (N_6530,N_3760,N_2400);
nand U6531 (N_6531,N_3762,N_3817);
or U6532 (N_6532,N_2348,N_2575);
nand U6533 (N_6533,N_2451,N_422);
xnor U6534 (N_6534,N_3527,N_197);
nand U6535 (N_6535,N_34,N_3499);
or U6536 (N_6536,N_4741,N_4669);
or U6537 (N_6537,N_830,N_2516);
nor U6538 (N_6538,N_3982,N_1473);
or U6539 (N_6539,N_781,N_2619);
or U6540 (N_6540,N_415,N_4587);
or U6541 (N_6541,N_2027,N_2279);
xor U6542 (N_6542,N_3185,N_2536);
and U6543 (N_6543,N_29,N_501);
and U6544 (N_6544,N_2647,N_1056);
nand U6545 (N_6545,N_3066,N_2237);
nand U6546 (N_6546,N_3409,N_3302);
nor U6547 (N_6547,N_4546,N_2188);
nand U6548 (N_6548,N_4400,N_3959);
or U6549 (N_6549,N_2190,N_3021);
or U6550 (N_6550,N_2908,N_4337);
and U6551 (N_6551,N_4639,N_2121);
nand U6552 (N_6552,N_4180,N_89);
or U6553 (N_6553,N_252,N_1375);
or U6554 (N_6554,N_4565,N_4897);
or U6555 (N_6555,N_736,N_4088);
nor U6556 (N_6556,N_1373,N_2502);
xor U6557 (N_6557,N_3834,N_3975);
or U6558 (N_6558,N_184,N_4040);
xor U6559 (N_6559,N_562,N_3121);
or U6560 (N_6560,N_3380,N_623);
or U6561 (N_6561,N_3963,N_2883);
nor U6562 (N_6562,N_1674,N_4387);
and U6563 (N_6563,N_4252,N_1522);
nor U6564 (N_6564,N_816,N_2663);
or U6565 (N_6565,N_4593,N_114);
or U6566 (N_6566,N_1654,N_1696);
or U6567 (N_6567,N_1121,N_512);
nor U6568 (N_6568,N_1597,N_4529);
xor U6569 (N_6569,N_1183,N_283);
xor U6570 (N_6570,N_4640,N_376);
and U6571 (N_6571,N_4305,N_2450);
nand U6572 (N_6572,N_1208,N_4592);
and U6573 (N_6573,N_208,N_3855);
nor U6574 (N_6574,N_3596,N_4244);
nand U6575 (N_6575,N_1609,N_3889);
xnor U6576 (N_6576,N_1320,N_918);
nand U6577 (N_6577,N_1048,N_357);
nand U6578 (N_6578,N_4933,N_851);
nand U6579 (N_6579,N_2443,N_2544);
nand U6580 (N_6580,N_1130,N_3657);
nand U6581 (N_6581,N_4366,N_3660);
or U6582 (N_6582,N_3052,N_4019);
and U6583 (N_6583,N_845,N_3672);
nand U6584 (N_6584,N_1253,N_4583);
or U6585 (N_6585,N_3248,N_4177);
nor U6586 (N_6586,N_4931,N_4860);
and U6587 (N_6587,N_3649,N_801);
nand U6588 (N_6588,N_4117,N_4147);
and U6589 (N_6589,N_639,N_4924);
nor U6590 (N_6590,N_2427,N_3055);
nor U6591 (N_6591,N_670,N_1606);
nand U6592 (N_6592,N_471,N_2223);
nor U6593 (N_6593,N_4918,N_3058);
nor U6594 (N_6594,N_2541,N_199);
nand U6595 (N_6595,N_4260,N_3187);
or U6596 (N_6596,N_2075,N_2855);
xor U6597 (N_6597,N_1284,N_1066);
and U6598 (N_6598,N_2009,N_233);
nand U6599 (N_6599,N_2927,N_3875);
and U6600 (N_6600,N_3123,N_3954);
nand U6601 (N_6601,N_3800,N_2019);
and U6602 (N_6602,N_1329,N_2569);
nor U6603 (N_6603,N_464,N_3746);
or U6604 (N_6604,N_1346,N_474);
or U6605 (N_6605,N_3216,N_4922);
or U6606 (N_6606,N_3396,N_4466);
nor U6607 (N_6607,N_4237,N_2572);
xnor U6608 (N_6608,N_4785,N_1514);
xor U6609 (N_6609,N_467,N_620);
xor U6610 (N_6610,N_2441,N_1338);
nand U6611 (N_6611,N_4902,N_1119);
nand U6612 (N_6612,N_4106,N_4209);
and U6613 (N_6613,N_4390,N_693);
or U6614 (N_6614,N_242,N_4964);
and U6615 (N_6615,N_1719,N_548);
nor U6616 (N_6616,N_4103,N_3600);
and U6617 (N_6617,N_831,N_2996);
xnor U6618 (N_6618,N_2054,N_3004);
nor U6619 (N_6619,N_3381,N_3218);
nor U6620 (N_6620,N_4364,N_2100);
nor U6621 (N_6621,N_2761,N_1258);
or U6622 (N_6622,N_4968,N_3874);
xnor U6623 (N_6623,N_4698,N_1906);
or U6624 (N_6624,N_3075,N_3517);
nand U6625 (N_6625,N_18,N_3412);
nor U6626 (N_6626,N_166,N_2628);
xnor U6627 (N_6627,N_4300,N_933);
or U6628 (N_6628,N_4697,N_3112);
xnor U6629 (N_6629,N_4486,N_4193);
nand U6630 (N_6630,N_739,N_2270);
nand U6631 (N_6631,N_379,N_2319);
nand U6632 (N_6632,N_1990,N_2727);
xor U6633 (N_6633,N_2617,N_2163);
nand U6634 (N_6634,N_1678,N_194);
nor U6635 (N_6635,N_2629,N_3012);
nor U6636 (N_6636,N_937,N_4580);
and U6637 (N_6637,N_4446,N_3667);
or U6638 (N_6638,N_2551,N_1006);
and U6639 (N_6639,N_210,N_2482);
or U6640 (N_6640,N_2004,N_2712);
xnor U6641 (N_6641,N_1863,N_1468);
nand U6642 (N_6642,N_1896,N_3919);
or U6643 (N_6643,N_3001,N_3105);
and U6644 (N_6644,N_2905,N_3711);
and U6645 (N_6645,N_3863,N_4261);
or U6646 (N_6646,N_3061,N_1911);
nor U6647 (N_6647,N_887,N_3135);
or U6648 (N_6648,N_1693,N_1957);
or U6649 (N_6649,N_3819,N_176);
or U6650 (N_6650,N_3933,N_4954);
nand U6651 (N_6651,N_2365,N_4449);
nand U6652 (N_6652,N_1782,N_4768);
and U6653 (N_6653,N_3158,N_3555);
and U6654 (N_6654,N_460,N_4801);
xor U6655 (N_6655,N_2069,N_1446);
or U6656 (N_6656,N_162,N_2106);
nand U6657 (N_6657,N_4101,N_4788);
nor U6658 (N_6658,N_2490,N_2283);
xnor U6659 (N_6659,N_4355,N_4084);
xor U6660 (N_6660,N_345,N_144);
xnor U6661 (N_6661,N_2593,N_410);
nor U6662 (N_6662,N_2950,N_1931);
nand U6663 (N_6663,N_1797,N_2928);
xor U6664 (N_6664,N_1404,N_2214);
and U6665 (N_6665,N_3623,N_342);
and U6666 (N_6666,N_695,N_27);
xnor U6667 (N_6667,N_1809,N_2989);
or U6668 (N_6668,N_1730,N_4797);
or U6669 (N_6669,N_1566,N_2633);
nand U6670 (N_6670,N_4067,N_3273);
and U6671 (N_6671,N_4655,N_402);
nor U6672 (N_6672,N_2229,N_3382);
nand U6673 (N_6673,N_3890,N_1816);
xor U6674 (N_6674,N_23,N_2314);
nor U6675 (N_6675,N_1059,N_4866);
xnor U6676 (N_6676,N_1808,N_1725);
and U6677 (N_6677,N_1451,N_4274);
nor U6678 (N_6678,N_2005,N_2002);
nor U6679 (N_6679,N_3698,N_1695);
nor U6680 (N_6680,N_2018,N_195);
or U6681 (N_6681,N_1569,N_665);
xor U6682 (N_6682,N_2384,N_2301);
nor U6683 (N_6683,N_535,N_885);
or U6684 (N_6684,N_15,N_3042);
xnor U6685 (N_6685,N_3067,N_3163);
nand U6686 (N_6686,N_2608,N_86);
and U6687 (N_6687,N_3951,N_1210);
xnor U6688 (N_6688,N_4650,N_3196);
nor U6689 (N_6689,N_4685,N_2659);
and U6690 (N_6690,N_98,N_4774);
nor U6691 (N_6691,N_420,N_1289);
xnor U6692 (N_6692,N_3447,N_797);
nand U6693 (N_6693,N_3830,N_1278);
or U6694 (N_6694,N_3098,N_497);
nand U6695 (N_6695,N_1740,N_3916);
or U6696 (N_6696,N_2373,N_3628);
nor U6697 (N_6697,N_1935,N_296);
or U6698 (N_6698,N_1354,N_3893);
xnor U6699 (N_6699,N_3801,N_3268);
and U6700 (N_6700,N_1685,N_88);
xor U6701 (N_6701,N_730,N_3719);
nand U6702 (N_6702,N_4026,N_1543);
nand U6703 (N_6703,N_3550,N_3213);
and U6704 (N_6704,N_4532,N_411);
or U6705 (N_6705,N_1310,N_505);
and U6706 (N_6706,N_2596,N_2961);
or U6707 (N_6707,N_3749,N_2919);
or U6708 (N_6708,N_1640,N_3126);
and U6709 (N_6709,N_2592,N_1288);
nand U6710 (N_6710,N_2045,N_3491);
and U6711 (N_6711,N_4634,N_2139);
nand U6712 (N_6712,N_155,N_3689);
or U6713 (N_6713,N_904,N_488);
nor U6714 (N_6714,N_61,N_4344);
xnor U6715 (N_6715,N_1095,N_2129);
nor U6716 (N_6716,N_387,N_2865);
or U6717 (N_6717,N_1675,N_3835);
nand U6718 (N_6718,N_1488,N_2752);
or U6719 (N_6719,N_4186,N_3289);
and U6720 (N_6720,N_2396,N_4110);
nand U6721 (N_6721,N_873,N_855);
and U6722 (N_6722,N_1903,N_2276);
and U6723 (N_6723,N_3877,N_1860);
or U6724 (N_6724,N_4370,N_211);
nor U6725 (N_6725,N_2832,N_80);
or U6726 (N_6726,N_2387,N_425);
xnor U6727 (N_6727,N_3290,N_707);
and U6728 (N_6728,N_2269,N_3836);
nor U6729 (N_6729,N_485,N_2421);
xor U6730 (N_6730,N_2534,N_4146);
nand U6731 (N_6731,N_2708,N_1825);
or U6732 (N_6732,N_2645,N_3773);
or U6733 (N_6733,N_3570,N_4830);
and U6734 (N_6734,N_139,N_1767);
or U6735 (N_6735,N_4250,N_3436);
and U6736 (N_6736,N_4188,N_3255);
nand U6737 (N_6737,N_602,N_3741);
or U6738 (N_6738,N_3214,N_3625);
nor U6739 (N_6739,N_1181,N_7);
and U6740 (N_6740,N_3515,N_2389);
nand U6741 (N_6741,N_2533,N_3794);
xnor U6742 (N_6742,N_2484,N_301);
and U6743 (N_6743,N_1790,N_4944);
or U6744 (N_6744,N_799,N_3696);
nand U6745 (N_6745,N_3865,N_4953);
and U6746 (N_6746,N_4952,N_4834);
xor U6747 (N_6747,N_1001,N_3639);
xnor U6748 (N_6748,N_1833,N_4430);
nand U6749 (N_6749,N_4256,N_539);
xnor U6750 (N_6750,N_4861,N_1586);
and U6751 (N_6751,N_2266,N_4055);
and U6752 (N_6752,N_102,N_4829);
or U6753 (N_6753,N_1359,N_1796);
nand U6754 (N_6754,N_1595,N_2132);
and U6755 (N_6755,N_2350,N_1182);
xnor U6756 (N_6756,N_380,N_4183);
or U6757 (N_6757,N_2743,N_3970);
and U6758 (N_6758,N_3498,N_1392);
nor U6759 (N_6759,N_3233,N_3857);
nand U6760 (N_6760,N_3805,N_3735);
xnor U6761 (N_6761,N_4108,N_3281);
and U6762 (N_6762,N_4483,N_2393);
and U6763 (N_6763,N_4462,N_2466);
or U6764 (N_6764,N_418,N_2483);
nand U6765 (N_6765,N_3461,N_2953);
or U6766 (N_6766,N_321,N_940);
xnor U6767 (N_6767,N_137,N_605);
nand U6768 (N_6768,N_1533,N_4516);
and U6769 (N_6769,N_642,N_4641);
nand U6770 (N_6770,N_1545,N_3991);
or U6771 (N_6771,N_3340,N_368);
xor U6772 (N_6772,N_4746,N_3521);
nand U6773 (N_6773,N_1944,N_4351);
nand U6774 (N_6774,N_1622,N_615);
and U6775 (N_6775,N_2442,N_1153);
or U6776 (N_6776,N_1490,N_3366);
nor U6777 (N_6777,N_3028,N_54);
xor U6778 (N_6778,N_717,N_69);
nor U6779 (N_6779,N_3378,N_3950);
nand U6780 (N_6780,N_173,N_2800);
and U6781 (N_6781,N_286,N_4156);
nor U6782 (N_6782,N_572,N_2322);
nor U6783 (N_6783,N_4196,N_3090);
or U6784 (N_6784,N_2289,N_2326);
nor U6785 (N_6785,N_3045,N_4557);
nand U6786 (N_6786,N_4298,N_2128);
nor U6787 (N_6787,N_1244,N_793);
or U6788 (N_6788,N_1312,N_1568);
or U6789 (N_6789,N_2032,N_3365);
nor U6790 (N_6790,N_4813,N_2093);
and U6791 (N_6791,N_1283,N_2236);
xor U6792 (N_6792,N_2425,N_3648);
or U6793 (N_6793,N_3971,N_72);
xnor U6794 (N_6794,N_1014,N_3611);
nand U6795 (N_6795,N_38,N_4269);
nand U6796 (N_6796,N_3733,N_4340);
nand U6797 (N_6797,N_4023,N_2475);
nor U6798 (N_6798,N_1779,N_4736);
or U6799 (N_6799,N_3574,N_1386);
and U6800 (N_6800,N_1093,N_1002);
nand U6801 (N_6801,N_429,N_4294);
nand U6802 (N_6802,N_3428,N_31);
nor U6803 (N_6803,N_4176,N_3472);
and U6804 (N_6804,N_2972,N_1017);
and U6805 (N_6805,N_2372,N_64);
nand U6806 (N_6806,N_1877,N_2198);
nand U6807 (N_6807,N_469,N_4247);
or U6808 (N_6808,N_1955,N_2700);
nor U6809 (N_6809,N_3392,N_132);
xnor U6810 (N_6810,N_2036,N_3252);
nand U6811 (N_6811,N_2797,N_2313);
or U6812 (N_6812,N_3369,N_209);
and U6813 (N_6813,N_4328,N_724);
nor U6814 (N_6814,N_1207,N_4155);
nand U6815 (N_6815,N_719,N_311);
or U6816 (N_6816,N_202,N_2978);
nor U6817 (N_6817,N_3906,N_19);
and U6818 (N_6818,N_1765,N_2050);
nand U6819 (N_6819,N_2941,N_4934);
nor U6820 (N_6820,N_2381,N_555);
nor U6821 (N_6821,N_3931,N_3307);
nor U6822 (N_6822,N_3176,N_1042);
or U6823 (N_6823,N_2385,N_4612);
or U6824 (N_6824,N_3397,N_1266);
xnor U6825 (N_6825,N_1794,N_3978);
nor U6826 (N_6826,N_352,N_835);
nor U6827 (N_6827,N_3691,N_2677);
and U6828 (N_6828,N_3459,N_923);
xnor U6829 (N_6829,N_2943,N_3102);
or U6830 (N_6830,N_2783,N_4661);
nor U6831 (N_6831,N_930,N_3808);
and U6832 (N_6832,N_2902,N_2599);
nor U6833 (N_6833,N_1848,N_977);
xor U6834 (N_6834,N_2058,N_4680);
and U6835 (N_6835,N_2532,N_2948);
and U6836 (N_6836,N_2481,N_4856);
nor U6837 (N_6837,N_616,N_1897);
xnor U6838 (N_6838,N_1908,N_650);
nand U6839 (N_6839,N_3807,N_847);
nor U6840 (N_6840,N_3172,N_3488);
or U6841 (N_6841,N_4425,N_681);
and U6842 (N_6842,N_4444,N_3463);
or U6843 (N_6843,N_3469,N_4521);
nand U6844 (N_6844,N_4428,N_4713);
or U6845 (N_6845,N_644,N_3283);
nor U6846 (N_6846,N_3016,N_4999);
or U6847 (N_6847,N_3481,N_4526);
nor U6848 (N_6848,N_4556,N_3263);
and U6849 (N_6849,N_3973,N_2380);
xnor U6850 (N_6850,N_4358,N_4127);
xnor U6851 (N_6851,N_2983,N_3663);
nand U6852 (N_6852,N_3908,N_3330);
nand U6853 (N_6853,N_2042,N_3680);
and U6854 (N_6854,N_3405,N_4596);
xor U6855 (N_6855,N_4460,N_984);
nand U6856 (N_6856,N_537,N_3583);
nand U6857 (N_6857,N_3470,N_3235);
and U6858 (N_6858,N_1350,N_2195);
xnor U6859 (N_6859,N_2073,N_2115);
xnor U6860 (N_6860,N_911,N_6);
xnor U6861 (N_6861,N_2444,N_291);
nand U6862 (N_6862,N_3996,N_492);
and U6863 (N_6863,N_4264,N_3769);
or U6864 (N_6864,N_4502,N_4925);
xor U6865 (N_6865,N_221,N_4613);
or U6866 (N_6866,N_747,N_3642);
nand U6867 (N_6867,N_2213,N_2942);
xnor U6868 (N_6868,N_3677,N_1120);
xor U6869 (N_6869,N_2717,N_445);
and U6870 (N_6870,N_2240,N_2709);
nand U6871 (N_6871,N_427,N_3684);
nand U6872 (N_6872,N_3844,N_964);
and U6873 (N_6873,N_1978,N_2571);
xnor U6874 (N_6874,N_4794,N_3907);
nand U6875 (N_6875,N_3060,N_3221);
or U6876 (N_6876,N_3180,N_3526);
xor U6877 (N_6877,N_404,N_4970);
nor U6878 (N_6878,N_2643,N_4584);
xor U6879 (N_6879,N_2992,N_2546);
or U6880 (N_6880,N_1218,N_1477);
or U6881 (N_6881,N_3725,N_130);
or U6882 (N_6882,N_250,N_613);
xor U6883 (N_6883,N_4220,N_3125);
xnor U6884 (N_6884,N_1664,N_4229);
nand U6885 (N_6885,N_697,N_3706);
and U6886 (N_6886,N_331,N_4386);
and U6887 (N_6887,N_13,N_2973);
nor U6888 (N_6888,N_4129,N_435);
or U6889 (N_6889,N_867,N_2921);
xor U6890 (N_6890,N_1134,N_1885);
or U6891 (N_6891,N_3030,N_4869);
xor U6892 (N_6892,N_3594,N_238);
xnor U6893 (N_6893,N_787,N_2863);
nor U6894 (N_6894,N_818,N_1132);
xnor U6895 (N_6895,N_364,N_3231);
and U6896 (N_6896,N_2966,N_3364);
xor U6897 (N_6897,N_1734,N_3601);
nor U6898 (N_6898,N_4078,N_1670);
and U6899 (N_6899,N_3759,N_4628);
xor U6900 (N_6900,N_1156,N_4230);
nor U6901 (N_6901,N_3921,N_1322);
nand U6902 (N_6902,N_3988,N_2108);
xor U6903 (N_6903,N_4507,N_3909);
nand U6904 (N_6904,N_1432,N_4572);
nand U6905 (N_6905,N_4306,N_4262);
nand U6906 (N_6906,N_3885,N_3478);
or U6907 (N_6907,N_1975,N_2359);
or U6908 (N_6908,N_4722,N_2646);
and U6909 (N_6909,N_3822,N_1305);
nand U6910 (N_6910,N_2044,N_468);
or U6911 (N_6911,N_2553,N_26);
and U6912 (N_6912,N_3913,N_725);
nor U6913 (N_6913,N_3726,N_893);
xnor U6914 (N_6914,N_4065,N_2661);
and U6915 (N_6915,N_484,N_3690);
and U6916 (N_6916,N_594,N_388);
xnor U6917 (N_6917,N_1485,N_771);
xor U6918 (N_6918,N_3884,N_1422);
or U6919 (N_6919,N_4770,N_970);
or U6920 (N_6920,N_1909,N_2084);
xor U6921 (N_6921,N_3206,N_972);
and U6922 (N_6922,N_4296,N_2878);
nor U6923 (N_6923,N_4051,N_1321);
xor U6924 (N_6924,N_67,N_3826);
nor U6925 (N_6925,N_3643,N_3151);
nand U6926 (N_6926,N_802,N_842);
nor U6927 (N_6927,N_4144,N_2029);
or U6928 (N_6928,N_4488,N_531);
and U6929 (N_6929,N_4632,N_4807);
and U6930 (N_6930,N_4975,N_3294);
nor U6931 (N_6931,N_4083,N_863);
nor U6932 (N_6932,N_1894,N_716);
xnor U6933 (N_6933,N_4349,N_4204);
and U6934 (N_6934,N_764,N_2191);
nor U6935 (N_6935,N_3401,N_2013);
nor U6936 (N_6936,N_4100,N_2773);
or U6937 (N_6937,N_765,N_2324);
xor U6938 (N_6938,N_2043,N_1342);
and U6939 (N_6939,N_113,N_519);
nand U6940 (N_6940,N_1209,N_1870);
or U6941 (N_6941,N_3901,N_1973);
nor U6942 (N_6942,N_1788,N_1055);
nand U6943 (N_6943,N_1025,N_2346);
xnor U6944 (N_6944,N_2135,N_4706);
nand U6945 (N_6945,N_438,N_3096);
nor U6946 (N_6946,N_1515,N_1444);
nand U6947 (N_6947,N_516,N_1143);
xnor U6948 (N_6948,N_4723,N_1570);
nor U6949 (N_6949,N_1857,N_2552);
nand U6950 (N_6950,N_4626,N_3468);
xor U6951 (N_6951,N_4822,N_4360);
nand U6952 (N_6952,N_783,N_590);
and U6953 (N_6953,N_4326,N_3232);
nand U6954 (N_6954,N_4292,N_4781);
or U6955 (N_6955,N_4559,N_1324);
xor U6956 (N_6956,N_2980,N_2046);
nor U6957 (N_6957,N_669,N_3018);
nor U6958 (N_6958,N_2614,N_4747);
nor U6959 (N_6959,N_4921,N_1256);
nand U6960 (N_6960,N_1528,N_3627);
xor U6961 (N_6961,N_4372,N_2187);
and U6962 (N_6962,N_2707,N_3622);
nor U6963 (N_6963,N_1495,N_1555);
or U6964 (N_6964,N_2723,N_2097);
or U6965 (N_6965,N_1298,N_1293);
nor U6966 (N_6966,N_812,N_3162);
nor U6967 (N_6967,N_4031,N_987);
xnor U6968 (N_6968,N_170,N_3764);
or U6969 (N_6969,N_1561,N_2669);
or U6970 (N_6970,N_3523,N_837);
and U6971 (N_6971,N_4763,N_3050);
and U6972 (N_6972,N_2104,N_4898);
xor U6973 (N_6973,N_2386,N_1562);
xor U6974 (N_6974,N_1866,N_4779);
or U6975 (N_6975,N_1441,N_4179);
xor U6976 (N_6976,N_3234,N_4824);
or U6977 (N_6977,N_2491,N_4004);
nand U6978 (N_6978,N_1874,N_1395);
nor U6979 (N_6979,N_2649,N_4130);
nor U6980 (N_6980,N_2699,N_434);
nor U6981 (N_6981,N_3998,N_1756);
and U6982 (N_6982,N_4579,N_4465);
or U6983 (N_6983,N_4037,N_982);
nor U6984 (N_6984,N_2930,N_3722);
nor U6985 (N_6985,N_4104,N_4799);
nor U6986 (N_6986,N_454,N_3275);
nor U6987 (N_6987,N_3493,N_1231);
and U6988 (N_6988,N_3048,N_4002);
and U6989 (N_6989,N_3455,N_1829);
or U6990 (N_6990,N_4335,N_1912);
nand U6991 (N_6991,N_135,N_3467);
and U6992 (N_6992,N_2356,N_3981);
xor U6993 (N_6993,N_2082,N_1560);
xnor U6994 (N_6994,N_3195,N_568);
and U6995 (N_6995,N_2123,N_3245);
and U6996 (N_6996,N_1803,N_4175);
nor U6997 (N_6997,N_631,N_40);
nor U6998 (N_6998,N_962,N_1306);
xor U6999 (N_6999,N_4034,N_980);
or U7000 (N_7000,N_2303,N_587);
or U7001 (N_7001,N_1748,N_1236);
or U7002 (N_7002,N_3529,N_4882);
nand U7003 (N_7003,N_3937,N_1753);
nand U7004 (N_7004,N_2500,N_3756);
and U7005 (N_7005,N_3246,N_4032);
and U7006 (N_7006,N_4014,N_4886);
and U7007 (N_7007,N_1750,N_4290);
nor U7008 (N_7008,N_4983,N_3101);
xor U7009 (N_7009,N_4543,N_328);
nand U7010 (N_7010,N_359,N_795);
nor U7011 (N_7011,N_2769,N_1738);
or U7012 (N_7012,N_278,N_2007);
xnor U7013 (N_7013,N_4792,N_3454);
or U7014 (N_7014,N_4730,N_3375);
xnor U7015 (N_7015,N_2732,N_2172);
or U7016 (N_7016,N_3177,N_710);
nor U7017 (N_7017,N_1516,N_1049);
nor U7018 (N_7018,N_1261,N_226);
or U7019 (N_7019,N_1163,N_168);
or U7020 (N_7020,N_3200,N_3033);
or U7021 (N_7021,N_965,N_2644);
xnor U7022 (N_7022,N_4473,N_1680);
or U7023 (N_7023,N_3783,N_3424);
nand U7024 (N_7024,N_4394,N_1615);
and U7025 (N_7025,N_2388,N_200);
nor U7026 (N_7026,N_344,N_4864);
or U7027 (N_7027,N_2438,N_4163);
or U7028 (N_7028,N_1456,N_2772);
and U7029 (N_7029,N_1844,N_1019);
nand U7030 (N_7030,N_3404,N_161);
nand U7031 (N_7031,N_1005,N_353);
nand U7032 (N_7032,N_470,N_2068);
nand U7033 (N_7033,N_3947,N_2495);
nand U7034 (N_7034,N_493,N_1745);
xnor U7035 (N_7035,N_2702,N_2851);
or U7036 (N_7036,N_4484,N_1706);
and U7037 (N_7037,N_2061,N_4821);
xnor U7038 (N_7038,N_1596,N_1045);
xor U7039 (N_7039,N_4467,N_1749);
nor U7040 (N_7040,N_1269,N_3450);
and U7041 (N_7041,N_2401,N_3668);
nand U7042 (N_7042,N_3356,N_1096);
xor U7043 (N_7043,N_33,N_1976);
and U7044 (N_7044,N_4615,N_4585);
nand U7045 (N_7045,N_4945,N_4629);
or U7046 (N_7046,N_3082,N_1357);
nor U7047 (N_7047,N_1044,N_1521);
nor U7048 (N_7048,N_2674,N_4844);
and U7049 (N_7049,N_1548,N_538);
nand U7050 (N_7050,N_618,N_806);
xnor U7051 (N_7051,N_4689,N_2520);
nand U7052 (N_7052,N_2716,N_4624);
nand U7053 (N_7053,N_2774,N_2864);
and U7054 (N_7054,N_4052,N_1141);
and U7055 (N_7055,N_3880,N_2072);
or U7056 (N_7056,N_4508,N_3647);
or U7057 (N_7057,N_1341,N_4419);
or U7058 (N_7058,N_892,N_2933);
and U7059 (N_7059,N_1655,N_2600);
or U7060 (N_7060,N_4928,N_4281);
nand U7061 (N_7061,N_905,N_528);
nor U7062 (N_7062,N_1037,N_658);
and U7063 (N_7063,N_2399,N_1859);
and U7064 (N_7064,N_958,N_3335);
xor U7065 (N_7065,N_917,N_2325);
nand U7066 (N_7066,N_4976,N_4965);
nor U7067 (N_7067,N_4563,N_2914);
xor U7068 (N_7068,N_4973,N_4093);
nor U7069 (N_7069,N_2297,N_1088);
nand U7070 (N_7070,N_2850,N_2877);
and U7071 (N_7071,N_3630,N_4648);
xor U7072 (N_7072,N_523,N_456);
and U7073 (N_7073,N_1420,N_3005);
nand U7074 (N_7074,N_1099,N_2197);
and U7075 (N_7075,N_473,N_4345);
nor U7076 (N_7076,N_1457,N_2151);
nor U7077 (N_7077,N_4905,N_1105);
and U7078 (N_7078,N_1190,N_3736);
nand U7079 (N_7079,N_2201,N_4069);
xnor U7080 (N_7080,N_4162,N_3850);
or U7081 (N_7081,N_1131,N_4338);
and U7082 (N_7082,N_11,N_4148);
nand U7083 (N_7083,N_3374,N_4504);
and U7084 (N_7084,N_3413,N_146);
and U7085 (N_7085,N_4378,N_1583);
nor U7086 (N_7086,N_475,N_3197);
or U7087 (N_7087,N_3932,N_289);
or U7088 (N_7088,N_1867,N_976);
or U7089 (N_7089,N_4820,N_4224);
nand U7090 (N_7090,N_1602,N_253);
xnor U7091 (N_7091,N_1948,N_914);
nand U7092 (N_7092,N_4566,N_1031);
or U7093 (N_7093,N_4076,N_983);
or U7094 (N_7094,N_2598,N_3700);
nand U7095 (N_7095,N_2957,N_550);
and U7096 (N_7096,N_4371,N_1072);
xor U7097 (N_7097,N_2689,N_3860);
xor U7098 (N_7098,N_4255,N_3837);
or U7099 (N_7099,N_3323,N_4087);
nand U7100 (N_7100,N_4263,N_1937);
and U7101 (N_7101,N_3546,N_1721);
nor U7102 (N_7102,N_186,N_3433);
or U7103 (N_7103,N_4672,N_1565);
or U7104 (N_7104,N_871,N_1390);
nor U7105 (N_7105,N_547,N_3466);
and U7106 (N_7106,N_363,N_786);
or U7107 (N_7107,N_2437,N_4158);
xor U7108 (N_7108,N_322,N_1453);
and U7109 (N_7109,N_583,N_2092);
and U7110 (N_7110,N_2095,N_4063);
or U7111 (N_7111,N_158,N_1260);
and U7112 (N_7112,N_2222,N_2077);
nor U7113 (N_7113,N_4573,N_2955);
nand U7114 (N_7114,N_2288,N_2120);
xnor U7115 (N_7115,N_2587,N_1421);
xnor U7116 (N_7116,N_4379,N_75);
xnor U7117 (N_7117,N_2311,N_705);
nor U7118 (N_7118,N_2904,N_4217);
nor U7119 (N_7119,N_1625,N_759);
and U7120 (N_7120,N_3712,N_2111);
or U7121 (N_7121,N_2060,N_1529);
xnor U7122 (N_7122,N_1050,N_4908);
xor U7123 (N_7123,N_544,N_128);
and U7124 (N_7124,N_3054,N_4202);
nor U7125 (N_7125,N_4686,N_2693);
or U7126 (N_7126,N_3873,N_3651);
nor U7127 (N_7127,N_487,N_1577);
nand U7128 (N_7128,N_4082,N_3840);
xor U7129 (N_7129,N_2275,N_2189);
and U7130 (N_7130,N_4917,N_1216);
or U7131 (N_7131,N_2537,N_3183);
and U7132 (N_7132,N_4142,N_1632);
and U7133 (N_7133,N_3025,N_223);
xor U7134 (N_7134,N_3032,N_1154);
xnor U7135 (N_7135,N_3578,N_3070);
or U7136 (N_7136,N_1133,N_4623);
nor U7137 (N_7137,N_1206,N_646);
nor U7138 (N_7138,N_1800,N_68);
xor U7139 (N_7139,N_360,N_249);
and U7140 (N_7140,N_1921,N_1205);
xnor U7141 (N_7141,N_2477,N_4701);
nor U7142 (N_7142,N_2827,N_3638);
nand U7143 (N_7143,N_4581,N_3787);
nand U7144 (N_7144,N_4432,N_3661);
or U7145 (N_7145,N_4012,N_2844);
nor U7146 (N_7146,N_4363,N_2822);
xor U7147 (N_7147,N_2165,N_3458);
xnor U7148 (N_7148,N_3475,N_4226);
xor U7149 (N_7149,N_570,N_822);
xnor U7150 (N_7150,N_1290,N_41);
nor U7151 (N_7151,N_3348,N_1179);
nor U7152 (N_7152,N_3754,N_1578);
and U7153 (N_7153,N_2831,N_4060);
nor U7154 (N_7154,N_735,N_4276);
and U7155 (N_7155,N_1604,N_4607);
nor U7156 (N_7156,N_1379,N_4283);
xnor U7157 (N_7157,N_329,N_4200);
xor U7158 (N_7158,N_4635,N_483);
nor U7159 (N_7159,N_1572,N_2001);
or U7160 (N_7160,N_4284,N_1532);
and U7161 (N_7161,N_2578,N_2529);
or U7162 (N_7162,N_3358,N_449);
nor U7163 (N_7163,N_3035,N_1868);
and U7164 (N_7164,N_1168,N_489);
and U7165 (N_7165,N_3324,N_4074);
and U7166 (N_7166,N_446,N_1594);
or U7167 (N_7167,N_4517,N_785);
and U7168 (N_7168,N_1219,N_722);
nor U7169 (N_7169,N_4597,N_1744);
nand U7170 (N_7170,N_1232,N_814);
xnor U7171 (N_7171,N_4727,N_3443);
nor U7172 (N_7172,N_2566,N_3940);
and U7173 (N_7173,N_115,N_3431);
or U7174 (N_7174,N_1727,N_3363);
nor U7175 (N_7175,N_1985,N_490);
nand U7176 (N_7176,N_895,N_1729);
or U7177 (N_7177,N_2091,N_3693);
or U7178 (N_7178,N_1307,N_37);
or U7179 (N_7179,N_2868,N_3803);
nor U7180 (N_7180,N_1709,N_1784);
xnor U7181 (N_7181,N_2583,N_3898);
and U7182 (N_7182,N_1761,N_3709);
or U7183 (N_7183,N_4426,N_3168);
nand U7184 (N_7184,N_3867,N_373);
and U7185 (N_7185,N_4988,N_1496);
and U7186 (N_7186,N_3014,N_3057);
nand U7187 (N_7187,N_3000,N_1697);
xnor U7188 (N_7188,N_4671,N_1551);
and U7189 (N_7189,N_3114,N_957);
or U7190 (N_7190,N_62,N_662);
nand U7191 (N_7191,N_1437,N_3771);
nand U7192 (N_7192,N_63,N_366);
nor U7193 (N_7193,N_4832,N_1078);
xnor U7194 (N_7194,N_4374,N_413);
nand U7195 (N_7195,N_805,N_262);
or U7196 (N_7196,N_563,N_2360);
xor U7197 (N_7197,N_1904,N_1411);
nand U7198 (N_7198,N_3682,N_2203);
and U7199 (N_7199,N_2125,N_2015);
nor U7200 (N_7200,N_2429,N_2917);
nor U7201 (N_7201,N_1101,N_4791);
nor U7202 (N_7202,N_4682,N_4926);
and U7203 (N_7203,N_1343,N_935);
and U7204 (N_7204,N_3186,N_347);
xor U7205 (N_7205,N_1620,N_2076);
or U7206 (N_7206,N_3716,N_4131);
nor U7207 (N_7207,N_4793,N_4783);
nor U7208 (N_7208,N_3318,N_436);
nor U7209 (N_7209,N_2519,N_4513);
or U7210 (N_7210,N_2758,N_4505);
or U7211 (N_7211,N_4479,N_1673);
nor U7212 (N_7212,N_4796,N_4890);
nor U7213 (N_7213,N_4434,N_526);
nand U7214 (N_7214,N_4190,N_3167);
or U7215 (N_7215,N_507,N_138);
or U7216 (N_7216,N_239,N_4267);
and U7217 (N_7217,N_1855,N_1195);
or U7218 (N_7218,N_3799,N_3602);
or U7219 (N_7219,N_1887,N_2059);
nor U7220 (N_7220,N_4203,N_632);
nor U7221 (N_7221,N_3618,N_659);
nand U7222 (N_7222,N_224,N_1160);
nand U7223 (N_7223,N_1920,N_2804);
nand U7224 (N_7224,N_2671,N_817);
and U7225 (N_7225,N_1220,N_4409);
nand U7226 (N_7226,N_4279,N_3514);
nand U7227 (N_7227,N_3056,N_1262);
nor U7228 (N_7228,N_3308,N_3418);
xor U7229 (N_7229,N_943,N_1000);
nor U7230 (N_7230,N_336,N_3371);
nor U7231 (N_7231,N_2336,N_3211);
xor U7232 (N_7232,N_3027,N_1237);
or U7233 (N_7233,N_2627,N_2690);
nand U7234 (N_7234,N_1367,N_305);
nor U7235 (N_7235,N_2178,N_1763);
xnor U7236 (N_7236,N_4691,N_4213);
xnor U7237 (N_7237,N_3311,N_3492);
nor U7238 (N_7238,N_3687,N_3271);
and U7239 (N_7239,N_1792,N_3333);
nor U7240 (N_7240,N_2618,N_1519);
nand U7241 (N_7241,N_3184,N_4373);
xnor U7242 (N_7242,N_247,N_2220);
or U7243 (N_7243,N_1347,N_1233);
and U7244 (N_7244,N_3518,N_3994);
nor U7245 (N_7245,N_4070,N_3777);
nand U7246 (N_7246,N_3946,N_4984);
nor U7247 (N_7247,N_2951,N_3291);
and U7248 (N_7248,N_1471,N_3804);
nand U7249 (N_7249,N_3189,N_237);
nor U7250 (N_7250,N_3679,N_1115);
or U7251 (N_7251,N_4920,N_256);
and U7252 (N_7252,N_3403,N_1743);
and U7253 (N_7253,N_3074,N_3895);
xor U7254 (N_7254,N_4470,N_4459);
nor U7255 (N_7255,N_2635,N_4234);
nor U7256 (N_7256,N_848,N_1073);
and U7257 (N_7257,N_2740,N_4091);
xor U7258 (N_7258,N_401,N_3486);
nand U7259 (N_7259,N_4541,N_4798);
nor U7260 (N_7260,N_967,N_25);
nand U7261 (N_7261,N_597,N_1954);
xnor U7262 (N_7262,N_4356,N_1212);
or U7263 (N_7263,N_496,N_652);
nor U7264 (N_7264,N_2161,N_1252);
nand U7265 (N_7265,N_3440,N_4595);
nor U7266 (N_7266,N_743,N_2866);
and U7267 (N_7267,N_3738,N_1462);
nor U7268 (N_7268,N_2756,N_3174);
nor U7269 (N_7269,N_3785,N_3558);
or U7270 (N_7270,N_3833,N_973);
and U7271 (N_7271,N_4993,N_49);
or U7272 (N_7272,N_3989,N_2836);
and U7273 (N_7273,N_1363,N_3223);
nor U7274 (N_7274,N_2293,N_4494);
xnor U7275 (N_7275,N_4138,N_3704);
nor U7276 (N_7276,N_3581,N_1691);
and U7277 (N_7277,N_1720,N_392);
and U7278 (N_7278,N_2328,N_2694);
xor U7279 (N_7279,N_4210,N_163);
nor U7280 (N_7280,N_3944,N_4149);
or U7281 (N_7281,N_1523,N_2147);
or U7282 (N_7282,N_2140,N_4790);
xnor U7283 (N_7283,N_2960,N_3093);
nor U7284 (N_7284,N_4249,N_1890);
or U7285 (N_7285,N_1351,N_3441);
or U7286 (N_7286,N_3866,N_1371);
nor U7287 (N_7287,N_4240,N_1977);
nand U7288 (N_7288,N_1663,N_462);
or U7289 (N_7289,N_1344,N_355);
and U7290 (N_7290,N_4315,N_3385);
and U7291 (N_7291,N_4375,N_557);
nor U7292 (N_7292,N_3138,N_1178);
or U7293 (N_7293,N_466,N_2456);
nand U7294 (N_7294,N_4506,N_2134);
nor U7295 (N_7295,N_367,N_498);
nor U7296 (N_7296,N_4872,N_2539);
or U7297 (N_7297,N_861,N_4875);
or U7298 (N_7298,N_2759,N_2548);
or U7299 (N_7299,N_944,N_227);
or U7300 (N_7300,N_4013,N_2081);
xnor U7301 (N_7301,N_1302,N_1452);
and U7302 (N_7302,N_3044,N_4);
nand U7303 (N_7303,N_4939,N_630);
xor U7304 (N_7304,N_3568,N_4317);
xnor U7305 (N_7305,N_481,N_2488);
and U7306 (N_7306,N_386,N_3797);
nand U7307 (N_7307,N_4135,N_4265);
nand U7308 (N_7308,N_4197,N_2173);
nand U7309 (N_7309,N_3072,N_721);
nand U7310 (N_7310,N_3111,N_4649);
and U7311 (N_7311,N_2252,N_4819);
nor U7312 (N_7312,N_1772,N_1936);
nor U7313 (N_7313,N_1224,N_3227);
and U7314 (N_7314,N_1255,N_4994);
xnor U7315 (N_7315,N_564,N_4675);
or U7316 (N_7316,N_3924,N_3133);
and U7317 (N_7317,N_3896,N_2815);
nand U7318 (N_7318,N_1982,N_890);
xor U7319 (N_7319,N_2781,N_3531);
nor U7320 (N_7320,N_1613,N_4550);
xnor U7321 (N_7321,N_43,N_4456);
and U7322 (N_7322,N_3952,N_4271);
or U7323 (N_7323,N_1257,N_4126);
nand U7324 (N_7324,N_2041,N_576);
nor U7325 (N_7325,N_1015,N_720);
xor U7326 (N_7326,N_290,N_2345);
nor U7327 (N_7327,N_4435,N_4608);
or U7328 (N_7328,N_4536,N_2530);
nor U7329 (N_7329,N_673,N_2420);
and U7330 (N_7330,N_541,N_2422);
nor U7331 (N_7331,N_566,N_1658);
nand U7332 (N_7332,N_1624,N_1162);
or U7333 (N_7333,N_414,N_1526);
or U7334 (N_7334,N_4322,N_4182);
xor U7335 (N_7335,N_2667,N_45);
xnor U7336 (N_7336,N_4966,N_3438);
nand U7337 (N_7337,N_4223,N_2936);
nor U7338 (N_7338,N_3930,N_2748);
and U7339 (N_7339,N_3556,N_3903);
nor U7340 (N_7340,N_1688,N_3503);
and U7341 (N_7341,N_3293,N_2591);
or U7342 (N_7342,N_4053,N_4709);
or U7343 (N_7343,N_2397,N_123);
nand U7344 (N_7344,N_4416,N_2231);
or U7345 (N_7345,N_4445,N_3595);
or U7346 (N_7346,N_3547,N_3979);
xor U7347 (N_7347,N_4889,N_3130);
and U7348 (N_7348,N_3744,N_4320);
nand U7349 (N_7349,N_3766,N_165);
and U7350 (N_7350,N_2691,N_2746);
and U7351 (N_7351,N_1889,N_1200);
or U7352 (N_7352,N_1724,N_2819);
or U7353 (N_7353,N_1916,N_3319);
nand U7354 (N_7354,N_2638,N_1217);
xor U7355 (N_7355,N_2390,N_1646);
nand U7356 (N_7356,N_2613,N_4896);
nand U7357 (N_7357,N_3191,N_4972);
xnor U7358 (N_7358,N_3806,N_4185);
xor U7359 (N_7359,N_580,N_4145);
xnor U7360 (N_7360,N_569,N_127);
nor U7361 (N_7361,N_4827,N_1415);
nand U7362 (N_7362,N_3490,N_378);
xor U7363 (N_7363,N_2323,N_189);
nor U7364 (N_7364,N_4427,N_3520);
xor U7365 (N_7365,N_3912,N_1886);
nand U7366 (N_7366,N_1238,N_3119);
or U7367 (N_7367,N_1757,N_2416);
nand U7368 (N_7368,N_840,N_4795);
nand U7369 (N_7369,N_1651,N_2067);
nand U7370 (N_7370,N_790,N_1581);
nand U7371 (N_7371,N_4207,N_4594);
and U7372 (N_7372,N_4228,N_1637);
xor U7373 (N_7373,N_4620,N_621);
and U7374 (N_7374,N_798,N_198);
xor U7375 (N_7375,N_44,N_1467);
or U7376 (N_7376,N_1541,N_2221);
nor U7377 (N_7377,N_4714,N_3747);
xor U7378 (N_7378,N_900,N_2786);
nor U7379 (N_7379,N_1984,N_3334);
or U7380 (N_7380,N_447,N_2413);
xnor U7381 (N_7381,N_1382,N_1881);
xnor U7382 (N_7382,N_93,N_2606);
nor U7383 (N_7383,N_1384,N_3287);
nand U7384 (N_7384,N_2753,N_2881);
or U7385 (N_7385,N_2028,N_2847);
or U7386 (N_7386,N_4001,N_2561);
nand U7387 (N_7387,N_4515,N_4321);
xor U7388 (N_7388,N_1227,N_1204);
and U7389 (N_7389,N_403,N_316);
or U7390 (N_7390,N_3188,N_2205);
xnor U7391 (N_7391,N_2505,N_2006);
xnor U7392 (N_7392,N_212,N_1713);
nand U7393 (N_7393,N_4665,N_2751);
and U7394 (N_7394,N_2849,N_1769);
xnor U7395 (N_7395,N_46,N_3482);
nand U7396 (N_7396,N_2736,N_282);
and U7397 (N_7397,N_4825,N_3645);
xnor U7398 (N_7398,N_2901,N_4877);
or U7399 (N_7399,N_2867,N_2364);
xor U7400 (N_7400,N_3586,N_3354);
xor U7401 (N_7401,N_2260,N_4674);
xor U7402 (N_7402,N_4392,N_4168);
xnor U7403 (N_7403,N_3320,N_4027);
xnor U7404 (N_7404,N_2449,N_1414);
xnor U7405 (N_7405,N_338,N_3205);
nor U7406 (N_7406,N_167,N_4656);
and U7407 (N_7407,N_3037,N_1271);
xnor U7408 (N_7408,N_3966,N_3537);
or U7409 (N_7409,N_2514,N_4657);
or U7410 (N_7410,N_1621,N_192);
nor U7411 (N_7411,N_1062,N_3831);
or U7412 (N_7412,N_4757,N_3345);
and U7413 (N_7413,N_3669,N_222);
and U7414 (N_7414,N_4522,N_3373);
nor U7415 (N_7415,N_769,N_2316);
nand U7416 (N_7416,N_3960,N_1423);
xor U7417 (N_7417,N_2459,N_1345);
nand U7418 (N_7418,N_3350,N_3820);
nor U7419 (N_7419,N_4858,N_1316);
or U7420 (N_7420,N_3110,N_777);
nor U7421 (N_7421,N_2903,N_3305);
xor U7422 (N_7422,N_2875,N_2517);
xnor U7423 (N_7423,N_2162,N_1240);
and U7424 (N_7424,N_1429,N_3297);
or U7425 (N_7425,N_4610,N_869);
nand U7426 (N_7426,N_3713,N_4385);
xnor U7427 (N_7427,N_4992,N_1512);
or U7428 (N_7428,N_251,N_2142);
xnor U7429 (N_7429,N_1927,N_1681);
nand U7430 (N_7430,N_750,N_323);
and U7431 (N_7431,N_4495,N_2242);
nand U7432 (N_7432,N_4453,N_1499);
or U7433 (N_7433,N_1348,N_2729);
nand U7434 (N_7434,N_2584,N_3753);
or U7435 (N_7435,N_4980,N_2182);
or U7436 (N_7436,N_153,N_2377);
and U7437 (N_7437,N_4160,N_343);
and U7438 (N_7438,N_2982,N_2987);
or U7439 (N_7439,N_2888,N_1003);
and U7440 (N_7440,N_4911,N_1786);
or U7441 (N_7441,N_2251,N_3708);
and U7442 (N_7442,N_284,N_1301);
or U7443 (N_7443,N_3506,N_2174);
nand U7444 (N_7444,N_1300,N_1151);
nor U7445 (N_7445,N_1234,N_2335);
nor U7446 (N_7446,N_2321,N_452);
nand U7447 (N_7447,N_3143,N_706);
or U7448 (N_7448,N_3730,N_3253);
or U7449 (N_7449,N_1294,N_4977);
or U7450 (N_7450,N_1992,N_4272);
nand U7451 (N_7451,N_1494,N_2458);
and U7452 (N_7452,N_258,N_3864);
and U7453 (N_7453,N_2631,N_409);
nor U7454 (N_7454,N_3926,N_451);
nand U7455 (N_7455,N_1676,N_3387);
nor U7456 (N_7456,N_2808,N_472);
nand U7457 (N_7457,N_2479,N_4323);
xnor U7458 (N_7458,N_634,N_2555);
or U7459 (N_7459,N_3444,N_4838);
xnor U7460 (N_7460,N_4075,N_361);
nor U7461 (N_7461,N_4421,N_3220);
nand U7462 (N_7462,N_1777,N_1385);
nor U7463 (N_7463,N_3192,N_3295);
xor U7464 (N_7464,N_567,N_3040);
nand U7465 (N_7465,N_1466,N_333);
nor U7466 (N_7466,N_1083,N_2207);
nand U7467 (N_7467,N_3051,N_694);
xor U7468 (N_7468,N_2344,N_2654);
and U7469 (N_7469,N_617,N_2975);
and U7470 (N_7470,N_3092,N_2605);
and U7471 (N_7471,N_2138,N_4420);
nor U7472 (N_7472,N_4863,N_1938);
or U7473 (N_7473,N_1650,N_1629);
nor U7474 (N_7474,N_4849,N_3328);
or U7475 (N_7475,N_3641,N_3124);
nand U7476 (N_7476,N_1542,N_1811);
nor U7477 (N_7477,N_3257,N_4463);
nand U7478 (N_7478,N_1349,N_1087);
nand U7479 (N_7479,N_868,N_3823);
or U7480 (N_7480,N_1852,N_1431);
or U7481 (N_7481,N_4625,N_2576);
nor U7482 (N_7482,N_1409,N_2358);
xor U7483 (N_7483,N_909,N_4011);
and U7484 (N_7484,N_2261,N_2035);
nand U7485 (N_7485,N_2368,N_2964);
nand U7486 (N_7486,N_276,N_2023);
nand U7487 (N_7487,N_3128,N_3838);
or U7488 (N_7488,N_2898,N_1012);
or U7489 (N_7489,N_94,N_3599);
or U7490 (N_7490,N_1117,N_1505);
and U7491 (N_7491,N_643,N_927);
nor U7492 (N_7492,N_3007,N_3851);
or U7493 (N_7493,N_4407,N_2049);
nand U7494 (N_7494,N_2852,N_149);
and U7495 (N_7495,N_3078,N_1074);
or U7496 (N_7496,N_4809,N_1508);
nor U7497 (N_7497,N_2507,N_2341);
nor U7498 (N_7498,N_393,N_3346);
nor U7499 (N_7499,N_2679,N_2206);
xor U7500 (N_7500,N_3486,N_415);
and U7501 (N_7501,N_2374,N_380);
nor U7502 (N_7502,N_420,N_3538);
and U7503 (N_7503,N_3790,N_4111);
nor U7504 (N_7504,N_3042,N_3779);
or U7505 (N_7505,N_2599,N_879);
nand U7506 (N_7506,N_1149,N_1816);
nand U7507 (N_7507,N_1251,N_2058);
xor U7508 (N_7508,N_2210,N_2814);
xor U7509 (N_7509,N_2583,N_4503);
xnor U7510 (N_7510,N_2868,N_3109);
nand U7511 (N_7511,N_122,N_1996);
xnor U7512 (N_7512,N_4228,N_510);
xor U7513 (N_7513,N_1350,N_2827);
xnor U7514 (N_7514,N_2187,N_3347);
nor U7515 (N_7515,N_3477,N_3913);
nor U7516 (N_7516,N_110,N_2837);
or U7517 (N_7517,N_249,N_631);
nand U7518 (N_7518,N_1939,N_4619);
nor U7519 (N_7519,N_946,N_4634);
xnor U7520 (N_7520,N_1942,N_1232);
nor U7521 (N_7521,N_4967,N_2386);
or U7522 (N_7522,N_505,N_3012);
and U7523 (N_7523,N_3631,N_2007);
or U7524 (N_7524,N_2006,N_4848);
nor U7525 (N_7525,N_3343,N_130);
xor U7526 (N_7526,N_466,N_4279);
nor U7527 (N_7527,N_4688,N_1523);
nor U7528 (N_7528,N_3177,N_1896);
nor U7529 (N_7529,N_1151,N_9);
nand U7530 (N_7530,N_2551,N_1030);
nor U7531 (N_7531,N_881,N_380);
and U7532 (N_7532,N_4348,N_1828);
nand U7533 (N_7533,N_705,N_1291);
or U7534 (N_7534,N_2775,N_4289);
nor U7535 (N_7535,N_4792,N_4398);
xnor U7536 (N_7536,N_3900,N_1638);
or U7537 (N_7537,N_3317,N_4546);
nand U7538 (N_7538,N_3720,N_2121);
nor U7539 (N_7539,N_2959,N_68);
xor U7540 (N_7540,N_3919,N_730);
and U7541 (N_7541,N_4824,N_3806);
nor U7542 (N_7542,N_1790,N_2447);
nand U7543 (N_7543,N_3511,N_2528);
nor U7544 (N_7544,N_1700,N_2847);
nand U7545 (N_7545,N_1257,N_1460);
and U7546 (N_7546,N_1763,N_2822);
nand U7547 (N_7547,N_3947,N_1403);
or U7548 (N_7548,N_2905,N_882);
and U7549 (N_7549,N_301,N_2025);
or U7550 (N_7550,N_1724,N_1737);
xor U7551 (N_7551,N_211,N_3745);
nor U7552 (N_7552,N_833,N_2604);
and U7553 (N_7553,N_936,N_3497);
xor U7554 (N_7554,N_1053,N_1983);
nand U7555 (N_7555,N_540,N_1976);
or U7556 (N_7556,N_243,N_2499);
nand U7557 (N_7557,N_4426,N_164);
nor U7558 (N_7558,N_3479,N_1731);
nand U7559 (N_7559,N_1764,N_1968);
nor U7560 (N_7560,N_649,N_392);
or U7561 (N_7561,N_278,N_112);
nor U7562 (N_7562,N_196,N_2721);
or U7563 (N_7563,N_1428,N_2860);
or U7564 (N_7564,N_1928,N_863);
and U7565 (N_7565,N_1696,N_518);
xnor U7566 (N_7566,N_4050,N_1009);
nor U7567 (N_7567,N_3802,N_2491);
nor U7568 (N_7568,N_4866,N_3966);
nor U7569 (N_7569,N_3161,N_4291);
or U7570 (N_7570,N_4373,N_4675);
and U7571 (N_7571,N_483,N_3332);
nor U7572 (N_7572,N_4602,N_3255);
xnor U7573 (N_7573,N_2907,N_3740);
nor U7574 (N_7574,N_1914,N_4806);
and U7575 (N_7575,N_1165,N_2650);
or U7576 (N_7576,N_1860,N_3207);
nand U7577 (N_7577,N_2354,N_3278);
and U7578 (N_7578,N_967,N_3312);
nand U7579 (N_7579,N_817,N_2059);
nand U7580 (N_7580,N_4380,N_1813);
or U7581 (N_7581,N_385,N_1263);
nand U7582 (N_7582,N_3733,N_1368);
xnor U7583 (N_7583,N_853,N_4303);
nand U7584 (N_7584,N_4912,N_456);
nand U7585 (N_7585,N_1253,N_4374);
and U7586 (N_7586,N_2164,N_3703);
nor U7587 (N_7587,N_4033,N_4607);
xnor U7588 (N_7588,N_3560,N_2021);
xor U7589 (N_7589,N_2939,N_2797);
nand U7590 (N_7590,N_4126,N_4251);
nand U7591 (N_7591,N_1588,N_856);
and U7592 (N_7592,N_882,N_1318);
xor U7593 (N_7593,N_197,N_4332);
nor U7594 (N_7594,N_629,N_2954);
or U7595 (N_7595,N_2881,N_4233);
or U7596 (N_7596,N_2767,N_4227);
xnor U7597 (N_7597,N_2902,N_3364);
nor U7598 (N_7598,N_872,N_2860);
xor U7599 (N_7599,N_1023,N_4501);
xnor U7600 (N_7600,N_4116,N_3050);
nor U7601 (N_7601,N_1624,N_2445);
and U7602 (N_7602,N_1560,N_267);
xor U7603 (N_7603,N_4874,N_3518);
nand U7604 (N_7604,N_215,N_4321);
or U7605 (N_7605,N_3894,N_3706);
nor U7606 (N_7606,N_3154,N_2789);
nor U7607 (N_7607,N_3433,N_4696);
and U7608 (N_7608,N_2569,N_400);
xnor U7609 (N_7609,N_3245,N_1360);
nor U7610 (N_7610,N_2762,N_690);
nor U7611 (N_7611,N_311,N_568);
nor U7612 (N_7612,N_812,N_3092);
or U7613 (N_7613,N_3742,N_4329);
nand U7614 (N_7614,N_1658,N_2981);
nand U7615 (N_7615,N_2698,N_1248);
nand U7616 (N_7616,N_3222,N_1174);
or U7617 (N_7617,N_2804,N_1696);
and U7618 (N_7618,N_4768,N_676);
xor U7619 (N_7619,N_2332,N_2637);
or U7620 (N_7620,N_239,N_1657);
and U7621 (N_7621,N_289,N_2543);
nor U7622 (N_7622,N_2330,N_979);
nor U7623 (N_7623,N_2292,N_4475);
nor U7624 (N_7624,N_3168,N_2801);
nor U7625 (N_7625,N_2723,N_3147);
or U7626 (N_7626,N_2492,N_1809);
xor U7627 (N_7627,N_327,N_797);
xor U7628 (N_7628,N_3056,N_3671);
nor U7629 (N_7629,N_4368,N_2624);
and U7630 (N_7630,N_4414,N_308);
and U7631 (N_7631,N_2179,N_959);
nor U7632 (N_7632,N_2470,N_2565);
nor U7633 (N_7633,N_1945,N_3160);
xor U7634 (N_7634,N_2324,N_2604);
nand U7635 (N_7635,N_4498,N_4389);
xnor U7636 (N_7636,N_2487,N_1659);
xor U7637 (N_7637,N_47,N_1310);
and U7638 (N_7638,N_1873,N_2876);
and U7639 (N_7639,N_2379,N_1034);
xnor U7640 (N_7640,N_120,N_158);
nor U7641 (N_7641,N_3565,N_3427);
nand U7642 (N_7642,N_2889,N_1336);
or U7643 (N_7643,N_1695,N_3820);
and U7644 (N_7644,N_2488,N_1719);
or U7645 (N_7645,N_3880,N_3710);
nand U7646 (N_7646,N_2355,N_3887);
nand U7647 (N_7647,N_110,N_1922);
or U7648 (N_7648,N_4179,N_4984);
xnor U7649 (N_7649,N_3380,N_2456);
nor U7650 (N_7650,N_1210,N_4526);
nor U7651 (N_7651,N_1404,N_674);
and U7652 (N_7652,N_2140,N_1905);
nor U7653 (N_7653,N_1554,N_2203);
xnor U7654 (N_7654,N_1143,N_3372);
or U7655 (N_7655,N_2387,N_866);
xnor U7656 (N_7656,N_2588,N_2416);
or U7657 (N_7657,N_1790,N_4448);
nor U7658 (N_7658,N_2027,N_3508);
and U7659 (N_7659,N_2019,N_93);
and U7660 (N_7660,N_1211,N_806);
or U7661 (N_7661,N_3214,N_2802);
or U7662 (N_7662,N_63,N_2395);
nor U7663 (N_7663,N_4068,N_211);
nor U7664 (N_7664,N_3870,N_3315);
nand U7665 (N_7665,N_3946,N_2485);
nor U7666 (N_7666,N_504,N_2048);
nor U7667 (N_7667,N_4098,N_1045);
nor U7668 (N_7668,N_4095,N_2684);
nor U7669 (N_7669,N_1997,N_1852);
xnor U7670 (N_7670,N_4856,N_1549);
xnor U7671 (N_7671,N_4576,N_3155);
xnor U7672 (N_7672,N_3555,N_268);
nor U7673 (N_7673,N_1462,N_2940);
or U7674 (N_7674,N_4470,N_368);
nor U7675 (N_7675,N_3770,N_4718);
and U7676 (N_7676,N_3685,N_4786);
xnor U7677 (N_7677,N_1158,N_798);
nor U7678 (N_7678,N_914,N_3017);
nor U7679 (N_7679,N_1612,N_2298);
nand U7680 (N_7680,N_4358,N_4149);
nand U7681 (N_7681,N_1133,N_1476);
and U7682 (N_7682,N_3810,N_3931);
or U7683 (N_7683,N_2879,N_967);
nor U7684 (N_7684,N_4724,N_4734);
nand U7685 (N_7685,N_4445,N_3864);
nand U7686 (N_7686,N_2200,N_4437);
nand U7687 (N_7687,N_2164,N_4802);
and U7688 (N_7688,N_3395,N_2091);
and U7689 (N_7689,N_79,N_4792);
nor U7690 (N_7690,N_4323,N_3496);
or U7691 (N_7691,N_2357,N_2780);
and U7692 (N_7692,N_3469,N_1732);
or U7693 (N_7693,N_4582,N_3702);
or U7694 (N_7694,N_2118,N_455);
or U7695 (N_7695,N_4978,N_2311);
nor U7696 (N_7696,N_4703,N_1024);
nor U7697 (N_7697,N_1349,N_4474);
nand U7698 (N_7698,N_4984,N_4471);
nor U7699 (N_7699,N_3802,N_906);
nand U7700 (N_7700,N_4008,N_3992);
xnor U7701 (N_7701,N_3720,N_943);
nor U7702 (N_7702,N_3325,N_1325);
xnor U7703 (N_7703,N_369,N_97);
nor U7704 (N_7704,N_1409,N_3879);
or U7705 (N_7705,N_3797,N_1861);
xor U7706 (N_7706,N_2639,N_3746);
nand U7707 (N_7707,N_1094,N_1475);
or U7708 (N_7708,N_127,N_540);
or U7709 (N_7709,N_4158,N_580);
or U7710 (N_7710,N_4206,N_4196);
xnor U7711 (N_7711,N_4339,N_709);
or U7712 (N_7712,N_1267,N_4389);
or U7713 (N_7713,N_2905,N_2194);
nand U7714 (N_7714,N_4646,N_233);
xnor U7715 (N_7715,N_243,N_3702);
nand U7716 (N_7716,N_1175,N_3136);
xor U7717 (N_7717,N_4389,N_4690);
nand U7718 (N_7718,N_3708,N_3629);
and U7719 (N_7719,N_655,N_4532);
nor U7720 (N_7720,N_4972,N_2889);
nand U7721 (N_7721,N_2149,N_3642);
nand U7722 (N_7722,N_4025,N_862);
nand U7723 (N_7723,N_26,N_3606);
and U7724 (N_7724,N_1166,N_1048);
nor U7725 (N_7725,N_1438,N_4414);
or U7726 (N_7726,N_3065,N_2071);
xnor U7727 (N_7727,N_980,N_1445);
nor U7728 (N_7728,N_1261,N_113);
xnor U7729 (N_7729,N_2214,N_1286);
and U7730 (N_7730,N_614,N_79);
nand U7731 (N_7731,N_4395,N_3189);
xor U7732 (N_7732,N_3756,N_1040);
and U7733 (N_7733,N_4304,N_1935);
nor U7734 (N_7734,N_145,N_2219);
xnor U7735 (N_7735,N_4722,N_4962);
or U7736 (N_7736,N_1825,N_108);
nor U7737 (N_7737,N_3645,N_3276);
nand U7738 (N_7738,N_2602,N_3254);
or U7739 (N_7739,N_1334,N_1993);
or U7740 (N_7740,N_4912,N_2531);
and U7741 (N_7741,N_597,N_2824);
nor U7742 (N_7742,N_1366,N_734);
and U7743 (N_7743,N_1026,N_2322);
nor U7744 (N_7744,N_504,N_1276);
and U7745 (N_7745,N_4258,N_4208);
nor U7746 (N_7746,N_637,N_4857);
nor U7747 (N_7747,N_701,N_3341);
nand U7748 (N_7748,N_69,N_509);
xor U7749 (N_7749,N_4981,N_2116);
nand U7750 (N_7750,N_933,N_1874);
and U7751 (N_7751,N_2973,N_3337);
xor U7752 (N_7752,N_3638,N_514);
or U7753 (N_7753,N_2460,N_4579);
xor U7754 (N_7754,N_4906,N_4451);
xnor U7755 (N_7755,N_4862,N_1062);
or U7756 (N_7756,N_1606,N_1759);
or U7757 (N_7757,N_3147,N_1758);
nor U7758 (N_7758,N_1676,N_1130);
nand U7759 (N_7759,N_1400,N_2299);
nand U7760 (N_7760,N_2351,N_4337);
xnor U7761 (N_7761,N_1111,N_4781);
and U7762 (N_7762,N_2005,N_3381);
and U7763 (N_7763,N_2150,N_2984);
or U7764 (N_7764,N_3322,N_2486);
xor U7765 (N_7765,N_2196,N_1921);
nor U7766 (N_7766,N_400,N_4449);
xnor U7767 (N_7767,N_3849,N_2648);
xnor U7768 (N_7768,N_2940,N_4793);
and U7769 (N_7769,N_3752,N_1977);
or U7770 (N_7770,N_3784,N_8);
and U7771 (N_7771,N_3520,N_2083);
nand U7772 (N_7772,N_3920,N_1268);
and U7773 (N_7773,N_4252,N_4599);
or U7774 (N_7774,N_4724,N_2938);
nor U7775 (N_7775,N_3631,N_2047);
and U7776 (N_7776,N_3729,N_976);
nand U7777 (N_7777,N_423,N_3037);
and U7778 (N_7778,N_4225,N_124);
nor U7779 (N_7779,N_2154,N_2177);
and U7780 (N_7780,N_1289,N_2849);
or U7781 (N_7781,N_4692,N_2633);
xor U7782 (N_7782,N_127,N_4177);
or U7783 (N_7783,N_3859,N_1373);
nor U7784 (N_7784,N_3465,N_4005);
or U7785 (N_7785,N_4979,N_3882);
or U7786 (N_7786,N_1934,N_3207);
or U7787 (N_7787,N_3520,N_1213);
xor U7788 (N_7788,N_789,N_636);
xor U7789 (N_7789,N_4699,N_709);
xnor U7790 (N_7790,N_525,N_169);
and U7791 (N_7791,N_1896,N_4568);
nand U7792 (N_7792,N_1435,N_4879);
xor U7793 (N_7793,N_2477,N_2145);
nor U7794 (N_7794,N_4259,N_3504);
nor U7795 (N_7795,N_3768,N_3626);
nand U7796 (N_7796,N_1150,N_208);
nor U7797 (N_7797,N_4877,N_172);
xor U7798 (N_7798,N_2276,N_2996);
or U7799 (N_7799,N_4882,N_3227);
nand U7800 (N_7800,N_2625,N_2397);
nor U7801 (N_7801,N_1985,N_3644);
nor U7802 (N_7802,N_4995,N_1722);
nor U7803 (N_7803,N_631,N_1254);
and U7804 (N_7804,N_4105,N_3726);
and U7805 (N_7805,N_111,N_4495);
and U7806 (N_7806,N_1972,N_1105);
and U7807 (N_7807,N_1051,N_1925);
nand U7808 (N_7808,N_1179,N_2106);
nor U7809 (N_7809,N_4747,N_1730);
xor U7810 (N_7810,N_1829,N_13);
nand U7811 (N_7811,N_3531,N_4004);
xnor U7812 (N_7812,N_4355,N_1961);
nand U7813 (N_7813,N_3076,N_1917);
or U7814 (N_7814,N_3412,N_1735);
and U7815 (N_7815,N_3870,N_1707);
nand U7816 (N_7816,N_1414,N_1849);
xor U7817 (N_7817,N_3841,N_3678);
nor U7818 (N_7818,N_3337,N_2370);
nand U7819 (N_7819,N_2736,N_2298);
nand U7820 (N_7820,N_1436,N_1893);
and U7821 (N_7821,N_1018,N_76);
and U7822 (N_7822,N_2076,N_2923);
nor U7823 (N_7823,N_799,N_4961);
or U7824 (N_7824,N_628,N_2934);
nand U7825 (N_7825,N_3873,N_1290);
and U7826 (N_7826,N_371,N_461);
nor U7827 (N_7827,N_4233,N_244);
or U7828 (N_7828,N_3779,N_2128);
xor U7829 (N_7829,N_2183,N_4822);
xnor U7830 (N_7830,N_4114,N_3344);
or U7831 (N_7831,N_3413,N_2424);
and U7832 (N_7832,N_4646,N_470);
and U7833 (N_7833,N_1429,N_1407);
and U7834 (N_7834,N_727,N_1302);
nand U7835 (N_7835,N_3765,N_2741);
xnor U7836 (N_7836,N_1491,N_1270);
or U7837 (N_7837,N_2213,N_2024);
and U7838 (N_7838,N_691,N_2963);
nand U7839 (N_7839,N_3257,N_869);
nor U7840 (N_7840,N_4469,N_432);
xor U7841 (N_7841,N_2368,N_4499);
xnor U7842 (N_7842,N_1551,N_2717);
nor U7843 (N_7843,N_1407,N_130);
and U7844 (N_7844,N_1942,N_3194);
xor U7845 (N_7845,N_3206,N_48);
nor U7846 (N_7846,N_652,N_2944);
or U7847 (N_7847,N_2360,N_317);
xnor U7848 (N_7848,N_582,N_1150);
xnor U7849 (N_7849,N_428,N_2340);
and U7850 (N_7850,N_3851,N_4021);
xor U7851 (N_7851,N_1593,N_3860);
or U7852 (N_7852,N_2115,N_2685);
nor U7853 (N_7853,N_860,N_571);
nand U7854 (N_7854,N_4180,N_3578);
xor U7855 (N_7855,N_1938,N_3149);
or U7856 (N_7856,N_446,N_2776);
nor U7857 (N_7857,N_3498,N_943);
nor U7858 (N_7858,N_3607,N_3455);
and U7859 (N_7859,N_4491,N_2834);
nand U7860 (N_7860,N_4222,N_2258);
nor U7861 (N_7861,N_1910,N_942);
nor U7862 (N_7862,N_555,N_1376);
nand U7863 (N_7863,N_1901,N_3510);
or U7864 (N_7864,N_3262,N_4876);
xor U7865 (N_7865,N_2553,N_4444);
and U7866 (N_7866,N_3831,N_3752);
or U7867 (N_7867,N_3928,N_1179);
and U7868 (N_7868,N_153,N_1726);
and U7869 (N_7869,N_4702,N_4729);
nor U7870 (N_7870,N_351,N_3054);
nand U7871 (N_7871,N_1395,N_1151);
or U7872 (N_7872,N_2631,N_1449);
or U7873 (N_7873,N_1686,N_4103);
and U7874 (N_7874,N_3040,N_2272);
xnor U7875 (N_7875,N_3385,N_27);
nand U7876 (N_7876,N_1334,N_1951);
nand U7877 (N_7877,N_3970,N_81);
nand U7878 (N_7878,N_348,N_2361);
or U7879 (N_7879,N_2241,N_3839);
or U7880 (N_7880,N_3478,N_687);
and U7881 (N_7881,N_1022,N_2257);
xor U7882 (N_7882,N_2843,N_3026);
nand U7883 (N_7883,N_3990,N_305);
nor U7884 (N_7884,N_2871,N_2088);
or U7885 (N_7885,N_3075,N_4863);
and U7886 (N_7886,N_1590,N_106);
nand U7887 (N_7887,N_2771,N_4153);
or U7888 (N_7888,N_1229,N_1623);
and U7889 (N_7889,N_2400,N_3136);
or U7890 (N_7890,N_2921,N_2974);
nand U7891 (N_7891,N_882,N_247);
nor U7892 (N_7892,N_2933,N_1531);
or U7893 (N_7893,N_4101,N_1620);
nor U7894 (N_7894,N_1509,N_1914);
and U7895 (N_7895,N_1375,N_4450);
nor U7896 (N_7896,N_2096,N_4103);
nor U7897 (N_7897,N_2735,N_1923);
or U7898 (N_7898,N_1046,N_4518);
nand U7899 (N_7899,N_2663,N_3733);
nor U7900 (N_7900,N_1408,N_3577);
or U7901 (N_7901,N_3414,N_4720);
and U7902 (N_7902,N_537,N_215);
nor U7903 (N_7903,N_2613,N_2552);
and U7904 (N_7904,N_1901,N_3918);
xnor U7905 (N_7905,N_746,N_3005);
xnor U7906 (N_7906,N_3721,N_4008);
and U7907 (N_7907,N_2042,N_2379);
or U7908 (N_7908,N_2821,N_1727);
or U7909 (N_7909,N_980,N_3907);
nor U7910 (N_7910,N_2092,N_1288);
xnor U7911 (N_7911,N_2820,N_4485);
xnor U7912 (N_7912,N_1555,N_3);
or U7913 (N_7913,N_4253,N_1342);
or U7914 (N_7914,N_4270,N_2938);
xor U7915 (N_7915,N_4191,N_3642);
nor U7916 (N_7916,N_1568,N_1358);
nor U7917 (N_7917,N_1907,N_2849);
or U7918 (N_7918,N_1058,N_2945);
nand U7919 (N_7919,N_4917,N_4725);
nand U7920 (N_7920,N_1805,N_299);
or U7921 (N_7921,N_2879,N_3696);
and U7922 (N_7922,N_3089,N_1654);
nand U7923 (N_7923,N_4370,N_4667);
and U7924 (N_7924,N_3102,N_4733);
or U7925 (N_7925,N_973,N_2007);
xnor U7926 (N_7926,N_4242,N_2838);
nor U7927 (N_7927,N_780,N_709);
or U7928 (N_7928,N_2614,N_1139);
nor U7929 (N_7929,N_3855,N_4547);
and U7930 (N_7930,N_1544,N_3745);
xor U7931 (N_7931,N_1118,N_2820);
nor U7932 (N_7932,N_3509,N_298);
nand U7933 (N_7933,N_864,N_2261);
nand U7934 (N_7934,N_701,N_3566);
nor U7935 (N_7935,N_1014,N_2544);
nand U7936 (N_7936,N_1399,N_3405);
or U7937 (N_7937,N_4475,N_120);
or U7938 (N_7938,N_3732,N_4479);
xor U7939 (N_7939,N_4820,N_4936);
and U7940 (N_7940,N_4639,N_1694);
or U7941 (N_7941,N_1564,N_3808);
nor U7942 (N_7942,N_4892,N_2020);
and U7943 (N_7943,N_1191,N_1271);
xor U7944 (N_7944,N_3255,N_4049);
and U7945 (N_7945,N_887,N_2246);
xnor U7946 (N_7946,N_1464,N_2137);
nand U7947 (N_7947,N_2393,N_1213);
nor U7948 (N_7948,N_4904,N_3504);
nand U7949 (N_7949,N_1409,N_2089);
xor U7950 (N_7950,N_54,N_4104);
and U7951 (N_7951,N_3441,N_2293);
nand U7952 (N_7952,N_2726,N_3588);
nor U7953 (N_7953,N_3676,N_2030);
or U7954 (N_7954,N_1335,N_2550);
nor U7955 (N_7955,N_1337,N_4049);
nor U7956 (N_7956,N_2235,N_629);
nand U7957 (N_7957,N_2579,N_4591);
nand U7958 (N_7958,N_2465,N_1036);
nand U7959 (N_7959,N_3465,N_2086);
xor U7960 (N_7960,N_2490,N_3121);
and U7961 (N_7961,N_4989,N_4150);
nand U7962 (N_7962,N_3135,N_2549);
nor U7963 (N_7963,N_165,N_3054);
or U7964 (N_7964,N_599,N_2917);
xnor U7965 (N_7965,N_4045,N_4036);
or U7966 (N_7966,N_1900,N_2430);
and U7967 (N_7967,N_4532,N_1400);
nor U7968 (N_7968,N_3097,N_488);
and U7969 (N_7969,N_2549,N_4837);
and U7970 (N_7970,N_1062,N_482);
nand U7971 (N_7971,N_3838,N_20);
or U7972 (N_7972,N_2053,N_3614);
and U7973 (N_7973,N_706,N_3699);
nand U7974 (N_7974,N_3120,N_3490);
xnor U7975 (N_7975,N_1237,N_4935);
and U7976 (N_7976,N_2069,N_3677);
nor U7977 (N_7977,N_1564,N_1687);
and U7978 (N_7978,N_705,N_3275);
or U7979 (N_7979,N_3258,N_1046);
nand U7980 (N_7980,N_2639,N_2074);
nand U7981 (N_7981,N_4407,N_17);
xor U7982 (N_7982,N_1783,N_2462);
nor U7983 (N_7983,N_2611,N_3522);
nor U7984 (N_7984,N_1561,N_98);
or U7985 (N_7985,N_3471,N_1769);
xor U7986 (N_7986,N_2251,N_3172);
or U7987 (N_7987,N_4562,N_2090);
xor U7988 (N_7988,N_1778,N_2306);
xor U7989 (N_7989,N_889,N_497);
xor U7990 (N_7990,N_482,N_3842);
nor U7991 (N_7991,N_2979,N_760);
nor U7992 (N_7992,N_1881,N_3832);
or U7993 (N_7993,N_2463,N_208);
and U7994 (N_7994,N_201,N_2754);
and U7995 (N_7995,N_3983,N_1326);
and U7996 (N_7996,N_4009,N_1812);
and U7997 (N_7997,N_2223,N_3564);
xor U7998 (N_7998,N_2416,N_1322);
nand U7999 (N_7999,N_2128,N_901);
xnor U8000 (N_8000,N_4633,N_2662);
xor U8001 (N_8001,N_1317,N_4105);
and U8002 (N_8002,N_2929,N_91);
and U8003 (N_8003,N_1393,N_735);
and U8004 (N_8004,N_4841,N_3168);
nand U8005 (N_8005,N_2598,N_2180);
nand U8006 (N_8006,N_3495,N_546);
nand U8007 (N_8007,N_1958,N_3809);
or U8008 (N_8008,N_2023,N_1843);
or U8009 (N_8009,N_418,N_3374);
xor U8010 (N_8010,N_3100,N_2063);
or U8011 (N_8011,N_4099,N_314);
nand U8012 (N_8012,N_1868,N_1960);
nand U8013 (N_8013,N_1353,N_4914);
nor U8014 (N_8014,N_4745,N_3415);
nand U8015 (N_8015,N_2741,N_4498);
nor U8016 (N_8016,N_4743,N_1675);
nor U8017 (N_8017,N_4845,N_998);
and U8018 (N_8018,N_1447,N_2315);
or U8019 (N_8019,N_4028,N_4778);
and U8020 (N_8020,N_3537,N_4480);
xnor U8021 (N_8021,N_1594,N_1903);
nor U8022 (N_8022,N_530,N_4648);
and U8023 (N_8023,N_862,N_1347);
xor U8024 (N_8024,N_4054,N_2312);
nor U8025 (N_8025,N_2461,N_475);
or U8026 (N_8026,N_1844,N_1477);
nor U8027 (N_8027,N_3950,N_3024);
and U8028 (N_8028,N_435,N_4049);
nand U8029 (N_8029,N_3912,N_4467);
xor U8030 (N_8030,N_943,N_1736);
nand U8031 (N_8031,N_202,N_3860);
and U8032 (N_8032,N_4545,N_4371);
xor U8033 (N_8033,N_3053,N_4032);
or U8034 (N_8034,N_4384,N_1545);
and U8035 (N_8035,N_4126,N_703);
xor U8036 (N_8036,N_3344,N_4121);
or U8037 (N_8037,N_142,N_841);
and U8038 (N_8038,N_3125,N_2706);
and U8039 (N_8039,N_4460,N_4507);
and U8040 (N_8040,N_2146,N_2092);
nor U8041 (N_8041,N_3990,N_1463);
and U8042 (N_8042,N_442,N_631);
nand U8043 (N_8043,N_1270,N_2607);
nand U8044 (N_8044,N_1800,N_984);
nor U8045 (N_8045,N_148,N_4153);
xnor U8046 (N_8046,N_2755,N_238);
nor U8047 (N_8047,N_1809,N_3049);
nand U8048 (N_8048,N_1240,N_4207);
or U8049 (N_8049,N_1713,N_4672);
xor U8050 (N_8050,N_4952,N_1130);
nor U8051 (N_8051,N_2523,N_767);
or U8052 (N_8052,N_3556,N_3200);
nand U8053 (N_8053,N_740,N_2629);
and U8054 (N_8054,N_346,N_2640);
xor U8055 (N_8055,N_3206,N_3106);
and U8056 (N_8056,N_1798,N_1376);
nand U8057 (N_8057,N_734,N_3185);
and U8058 (N_8058,N_1993,N_660);
nand U8059 (N_8059,N_2949,N_2485);
and U8060 (N_8060,N_2472,N_3112);
and U8061 (N_8061,N_322,N_3253);
or U8062 (N_8062,N_36,N_4457);
nand U8063 (N_8063,N_2454,N_1988);
and U8064 (N_8064,N_2680,N_3637);
xor U8065 (N_8065,N_4398,N_1649);
and U8066 (N_8066,N_3632,N_3369);
or U8067 (N_8067,N_2187,N_3152);
nand U8068 (N_8068,N_3889,N_4286);
nor U8069 (N_8069,N_1370,N_3890);
xnor U8070 (N_8070,N_1830,N_2883);
xnor U8071 (N_8071,N_2420,N_3439);
nor U8072 (N_8072,N_934,N_1288);
and U8073 (N_8073,N_4813,N_2268);
nand U8074 (N_8074,N_4933,N_4282);
xor U8075 (N_8075,N_2378,N_2542);
nand U8076 (N_8076,N_4139,N_2936);
or U8077 (N_8077,N_1141,N_4850);
xor U8078 (N_8078,N_698,N_3202);
or U8079 (N_8079,N_873,N_1824);
nor U8080 (N_8080,N_3723,N_3487);
and U8081 (N_8081,N_881,N_1800);
nor U8082 (N_8082,N_1607,N_2405);
xor U8083 (N_8083,N_2636,N_2607);
nor U8084 (N_8084,N_2848,N_1563);
xor U8085 (N_8085,N_4873,N_710);
and U8086 (N_8086,N_4119,N_4201);
and U8087 (N_8087,N_2932,N_3947);
nor U8088 (N_8088,N_3641,N_4362);
and U8089 (N_8089,N_3545,N_1966);
or U8090 (N_8090,N_2821,N_4170);
and U8091 (N_8091,N_3642,N_4121);
and U8092 (N_8092,N_3015,N_519);
xor U8093 (N_8093,N_3776,N_3796);
and U8094 (N_8094,N_4434,N_4305);
or U8095 (N_8095,N_2546,N_2159);
xnor U8096 (N_8096,N_658,N_2370);
or U8097 (N_8097,N_1254,N_1846);
nor U8098 (N_8098,N_3822,N_4036);
or U8099 (N_8099,N_680,N_1557);
nor U8100 (N_8100,N_1658,N_3468);
and U8101 (N_8101,N_4611,N_1235);
or U8102 (N_8102,N_1873,N_3483);
nor U8103 (N_8103,N_4956,N_1606);
or U8104 (N_8104,N_2861,N_2214);
or U8105 (N_8105,N_1052,N_168);
xnor U8106 (N_8106,N_1447,N_1165);
nor U8107 (N_8107,N_1454,N_404);
xnor U8108 (N_8108,N_1302,N_305);
nor U8109 (N_8109,N_1816,N_2322);
xnor U8110 (N_8110,N_1627,N_3358);
nand U8111 (N_8111,N_4308,N_2542);
nor U8112 (N_8112,N_2184,N_3696);
nand U8113 (N_8113,N_721,N_1378);
nor U8114 (N_8114,N_2921,N_4126);
xnor U8115 (N_8115,N_2378,N_4045);
nor U8116 (N_8116,N_2700,N_4956);
and U8117 (N_8117,N_3123,N_1687);
xor U8118 (N_8118,N_1803,N_3565);
and U8119 (N_8119,N_2406,N_970);
xnor U8120 (N_8120,N_2134,N_60);
or U8121 (N_8121,N_4865,N_4610);
or U8122 (N_8122,N_1445,N_2048);
xnor U8123 (N_8123,N_1440,N_4156);
and U8124 (N_8124,N_3506,N_3005);
nor U8125 (N_8125,N_2357,N_1050);
nand U8126 (N_8126,N_3181,N_1077);
nor U8127 (N_8127,N_2870,N_3008);
xor U8128 (N_8128,N_4907,N_4932);
nand U8129 (N_8129,N_3208,N_844);
xor U8130 (N_8130,N_1218,N_4282);
xor U8131 (N_8131,N_299,N_3759);
or U8132 (N_8132,N_4382,N_2172);
or U8133 (N_8133,N_2207,N_1647);
or U8134 (N_8134,N_2296,N_3098);
xor U8135 (N_8135,N_430,N_984);
nand U8136 (N_8136,N_56,N_4776);
nand U8137 (N_8137,N_3660,N_3328);
nand U8138 (N_8138,N_4075,N_3556);
or U8139 (N_8139,N_4077,N_4447);
nor U8140 (N_8140,N_2167,N_1343);
and U8141 (N_8141,N_4546,N_4271);
nand U8142 (N_8142,N_2766,N_4161);
nand U8143 (N_8143,N_2396,N_2931);
xnor U8144 (N_8144,N_4304,N_1331);
and U8145 (N_8145,N_2770,N_1108);
xor U8146 (N_8146,N_1413,N_568);
or U8147 (N_8147,N_2440,N_4634);
and U8148 (N_8148,N_4792,N_1237);
and U8149 (N_8149,N_2243,N_1315);
nand U8150 (N_8150,N_2845,N_3410);
xor U8151 (N_8151,N_3738,N_532);
xnor U8152 (N_8152,N_735,N_2180);
nor U8153 (N_8153,N_1226,N_4420);
and U8154 (N_8154,N_1500,N_593);
xor U8155 (N_8155,N_842,N_1816);
xor U8156 (N_8156,N_1016,N_4357);
nand U8157 (N_8157,N_496,N_1065);
nor U8158 (N_8158,N_1011,N_1107);
and U8159 (N_8159,N_4295,N_652);
nor U8160 (N_8160,N_1578,N_3776);
and U8161 (N_8161,N_1986,N_1039);
and U8162 (N_8162,N_500,N_4167);
or U8163 (N_8163,N_4313,N_2744);
nand U8164 (N_8164,N_1869,N_4702);
or U8165 (N_8165,N_4515,N_798);
and U8166 (N_8166,N_3362,N_1421);
or U8167 (N_8167,N_514,N_1430);
or U8168 (N_8168,N_1512,N_724);
xor U8169 (N_8169,N_717,N_2456);
nor U8170 (N_8170,N_2467,N_556);
nand U8171 (N_8171,N_3433,N_369);
or U8172 (N_8172,N_3488,N_2804);
nor U8173 (N_8173,N_4871,N_2997);
nor U8174 (N_8174,N_224,N_3449);
nand U8175 (N_8175,N_3530,N_2698);
or U8176 (N_8176,N_432,N_538);
nand U8177 (N_8177,N_3790,N_252);
or U8178 (N_8178,N_1561,N_387);
nor U8179 (N_8179,N_497,N_1948);
and U8180 (N_8180,N_397,N_2464);
xnor U8181 (N_8181,N_3732,N_2512);
nor U8182 (N_8182,N_2977,N_4303);
nand U8183 (N_8183,N_1438,N_3052);
and U8184 (N_8184,N_3158,N_2060);
nand U8185 (N_8185,N_1117,N_3336);
nor U8186 (N_8186,N_4000,N_2433);
and U8187 (N_8187,N_2734,N_1312);
or U8188 (N_8188,N_3168,N_302);
xnor U8189 (N_8189,N_1246,N_2523);
nand U8190 (N_8190,N_959,N_2395);
or U8191 (N_8191,N_1185,N_4430);
xnor U8192 (N_8192,N_4227,N_3488);
nand U8193 (N_8193,N_2297,N_1423);
nand U8194 (N_8194,N_322,N_693);
or U8195 (N_8195,N_177,N_1858);
or U8196 (N_8196,N_3128,N_3005);
xor U8197 (N_8197,N_337,N_4663);
nand U8198 (N_8198,N_1189,N_159);
xor U8199 (N_8199,N_4450,N_3565);
xnor U8200 (N_8200,N_4410,N_2789);
nor U8201 (N_8201,N_3547,N_1649);
xor U8202 (N_8202,N_3203,N_2452);
nor U8203 (N_8203,N_1275,N_1193);
nor U8204 (N_8204,N_937,N_2183);
nand U8205 (N_8205,N_600,N_2553);
xnor U8206 (N_8206,N_3398,N_3192);
and U8207 (N_8207,N_325,N_4945);
nand U8208 (N_8208,N_3239,N_1796);
or U8209 (N_8209,N_1681,N_3406);
and U8210 (N_8210,N_4414,N_723);
nor U8211 (N_8211,N_3317,N_1837);
xnor U8212 (N_8212,N_2782,N_2200);
xor U8213 (N_8213,N_913,N_4128);
or U8214 (N_8214,N_2070,N_253);
and U8215 (N_8215,N_2468,N_4354);
and U8216 (N_8216,N_4095,N_1948);
nor U8217 (N_8217,N_56,N_340);
or U8218 (N_8218,N_2005,N_3484);
nand U8219 (N_8219,N_1775,N_3040);
nand U8220 (N_8220,N_1215,N_4310);
and U8221 (N_8221,N_3764,N_3119);
xnor U8222 (N_8222,N_3398,N_3025);
or U8223 (N_8223,N_1776,N_374);
xor U8224 (N_8224,N_3445,N_3181);
xor U8225 (N_8225,N_273,N_802);
or U8226 (N_8226,N_2372,N_605);
nand U8227 (N_8227,N_3424,N_3850);
nor U8228 (N_8228,N_1063,N_4259);
and U8229 (N_8229,N_3987,N_115);
xor U8230 (N_8230,N_1213,N_2305);
and U8231 (N_8231,N_3940,N_3337);
and U8232 (N_8232,N_1324,N_319);
xnor U8233 (N_8233,N_4125,N_4831);
xor U8234 (N_8234,N_927,N_2257);
xor U8235 (N_8235,N_3024,N_2143);
nor U8236 (N_8236,N_1736,N_4631);
or U8237 (N_8237,N_3617,N_4614);
or U8238 (N_8238,N_2653,N_2741);
and U8239 (N_8239,N_4255,N_4614);
nor U8240 (N_8240,N_2549,N_2868);
nand U8241 (N_8241,N_2035,N_4324);
nor U8242 (N_8242,N_2728,N_2812);
xor U8243 (N_8243,N_2745,N_4147);
or U8244 (N_8244,N_3439,N_2445);
and U8245 (N_8245,N_1681,N_3887);
or U8246 (N_8246,N_2636,N_4695);
nand U8247 (N_8247,N_1984,N_1472);
xor U8248 (N_8248,N_958,N_4477);
xor U8249 (N_8249,N_2970,N_3107);
xnor U8250 (N_8250,N_4927,N_4663);
and U8251 (N_8251,N_4406,N_1340);
or U8252 (N_8252,N_1458,N_4203);
nor U8253 (N_8253,N_4520,N_2593);
xor U8254 (N_8254,N_3681,N_4911);
nor U8255 (N_8255,N_3593,N_1851);
nand U8256 (N_8256,N_478,N_4673);
nor U8257 (N_8257,N_4072,N_1462);
and U8258 (N_8258,N_578,N_4498);
or U8259 (N_8259,N_4550,N_3465);
xnor U8260 (N_8260,N_742,N_4349);
nand U8261 (N_8261,N_50,N_2792);
nand U8262 (N_8262,N_4943,N_1117);
nand U8263 (N_8263,N_3015,N_3797);
nand U8264 (N_8264,N_2561,N_3947);
nand U8265 (N_8265,N_2407,N_176);
or U8266 (N_8266,N_3330,N_1234);
nor U8267 (N_8267,N_3908,N_2274);
and U8268 (N_8268,N_706,N_4573);
nand U8269 (N_8269,N_3200,N_4882);
or U8270 (N_8270,N_152,N_3052);
and U8271 (N_8271,N_3400,N_1526);
nand U8272 (N_8272,N_1313,N_1385);
nand U8273 (N_8273,N_4922,N_1440);
nor U8274 (N_8274,N_3280,N_4121);
nor U8275 (N_8275,N_629,N_3848);
nand U8276 (N_8276,N_157,N_2088);
or U8277 (N_8277,N_3335,N_1097);
nor U8278 (N_8278,N_848,N_3459);
xnor U8279 (N_8279,N_1635,N_3526);
nand U8280 (N_8280,N_67,N_1455);
and U8281 (N_8281,N_1606,N_3227);
nand U8282 (N_8282,N_1862,N_2240);
nand U8283 (N_8283,N_1009,N_4711);
or U8284 (N_8284,N_2610,N_3690);
xnor U8285 (N_8285,N_2524,N_39);
nor U8286 (N_8286,N_3189,N_1560);
nor U8287 (N_8287,N_3406,N_3343);
and U8288 (N_8288,N_2819,N_2570);
or U8289 (N_8289,N_4094,N_4936);
nand U8290 (N_8290,N_1184,N_4382);
xor U8291 (N_8291,N_1072,N_3038);
and U8292 (N_8292,N_2762,N_518);
nand U8293 (N_8293,N_4059,N_2028);
xor U8294 (N_8294,N_2987,N_1902);
nand U8295 (N_8295,N_4616,N_2860);
nand U8296 (N_8296,N_3124,N_679);
xnor U8297 (N_8297,N_1382,N_442);
xor U8298 (N_8298,N_997,N_4059);
or U8299 (N_8299,N_4673,N_1211);
nor U8300 (N_8300,N_2601,N_504);
or U8301 (N_8301,N_2877,N_3271);
nor U8302 (N_8302,N_4412,N_1332);
nand U8303 (N_8303,N_1504,N_4701);
xnor U8304 (N_8304,N_4723,N_4495);
xnor U8305 (N_8305,N_2817,N_3176);
and U8306 (N_8306,N_276,N_4049);
nor U8307 (N_8307,N_2928,N_1581);
and U8308 (N_8308,N_2673,N_2722);
xnor U8309 (N_8309,N_1450,N_1745);
and U8310 (N_8310,N_2265,N_148);
nand U8311 (N_8311,N_4565,N_4934);
and U8312 (N_8312,N_1208,N_3199);
xnor U8313 (N_8313,N_3377,N_373);
or U8314 (N_8314,N_4196,N_1962);
xor U8315 (N_8315,N_2675,N_3884);
or U8316 (N_8316,N_4642,N_920);
and U8317 (N_8317,N_3059,N_4253);
or U8318 (N_8318,N_4883,N_3545);
and U8319 (N_8319,N_3933,N_667);
xnor U8320 (N_8320,N_3327,N_241);
nand U8321 (N_8321,N_2865,N_306);
and U8322 (N_8322,N_4921,N_1514);
xor U8323 (N_8323,N_3570,N_4421);
nor U8324 (N_8324,N_4488,N_1531);
xnor U8325 (N_8325,N_2287,N_1874);
and U8326 (N_8326,N_3504,N_2174);
nand U8327 (N_8327,N_2654,N_1414);
nand U8328 (N_8328,N_515,N_2711);
or U8329 (N_8329,N_3837,N_3656);
and U8330 (N_8330,N_955,N_3836);
xor U8331 (N_8331,N_61,N_2275);
or U8332 (N_8332,N_13,N_1027);
nor U8333 (N_8333,N_3547,N_4707);
and U8334 (N_8334,N_1892,N_4871);
or U8335 (N_8335,N_3632,N_4938);
nand U8336 (N_8336,N_3768,N_4680);
xnor U8337 (N_8337,N_519,N_3598);
nand U8338 (N_8338,N_1933,N_1882);
nand U8339 (N_8339,N_4129,N_2768);
or U8340 (N_8340,N_1798,N_2691);
xor U8341 (N_8341,N_3302,N_1910);
or U8342 (N_8342,N_4165,N_4301);
nor U8343 (N_8343,N_3024,N_2134);
nor U8344 (N_8344,N_1047,N_1539);
or U8345 (N_8345,N_1127,N_3401);
and U8346 (N_8346,N_1587,N_3189);
or U8347 (N_8347,N_1508,N_2293);
nor U8348 (N_8348,N_1401,N_3668);
nand U8349 (N_8349,N_4347,N_4067);
xor U8350 (N_8350,N_2173,N_4188);
nand U8351 (N_8351,N_2183,N_481);
nand U8352 (N_8352,N_1441,N_2020);
xor U8353 (N_8353,N_2992,N_3458);
nand U8354 (N_8354,N_176,N_1260);
nand U8355 (N_8355,N_3058,N_3666);
nand U8356 (N_8356,N_1082,N_3380);
nor U8357 (N_8357,N_1790,N_4854);
nor U8358 (N_8358,N_3582,N_1449);
nand U8359 (N_8359,N_1203,N_3446);
xor U8360 (N_8360,N_2110,N_2048);
or U8361 (N_8361,N_3609,N_4739);
xor U8362 (N_8362,N_728,N_3236);
nor U8363 (N_8363,N_3724,N_2002);
nor U8364 (N_8364,N_237,N_893);
nand U8365 (N_8365,N_1800,N_4938);
and U8366 (N_8366,N_1701,N_4551);
and U8367 (N_8367,N_3614,N_3408);
and U8368 (N_8368,N_1749,N_1447);
and U8369 (N_8369,N_2192,N_4008);
nor U8370 (N_8370,N_3300,N_338);
or U8371 (N_8371,N_4018,N_3572);
nand U8372 (N_8372,N_337,N_1492);
and U8373 (N_8373,N_4486,N_942);
nand U8374 (N_8374,N_1309,N_2558);
nand U8375 (N_8375,N_4188,N_2950);
or U8376 (N_8376,N_2701,N_1476);
nor U8377 (N_8377,N_886,N_4418);
xor U8378 (N_8378,N_1068,N_1569);
nand U8379 (N_8379,N_2826,N_4663);
xnor U8380 (N_8380,N_4106,N_4557);
nand U8381 (N_8381,N_4544,N_2747);
and U8382 (N_8382,N_1757,N_1754);
nand U8383 (N_8383,N_246,N_4510);
nand U8384 (N_8384,N_4050,N_4939);
or U8385 (N_8385,N_1230,N_3881);
and U8386 (N_8386,N_214,N_181);
and U8387 (N_8387,N_1154,N_3124);
nand U8388 (N_8388,N_3766,N_4875);
xnor U8389 (N_8389,N_4083,N_4114);
nand U8390 (N_8390,N_2546,N_3282);
nand U8391 (N_8391,N_4427,N_2152);
or U8392 (N_8392,N_4521,N_692);
nand U8393 (N_8393,N_2301,N_2185);
or U8394 (N_8394,N_3000,N_3214);
and U8395 (N_8395,N_271,N_317);
nand U8396 (N_8396,N_4007,N_3103);
nand U8397 (N_8397,N_2748,N_4524);
and U8398 (N_8398,N_2720,N_4555);
nand U8399 (N_8399,N_3467,N_4184);
and U8400 (N_8400,N_2184,N_4322);
nand U8401 (N_8401,N_1005,N_1043);
nor U8402 (N_8402,N_3117,N_1842);
or U8403 (N_8403,N_4333,N_3382);
nor U8404 (N_8404,N_15,N_3010);
or U8405 (N_8405,N_1154,N_2266);
xnor U8406 (N_8406,N_2799,N_4539);
and U8407 (N_8407,N_170,N_1205);
nor U8408 (N_8408,N_635,N_1373);
or U8409 (N_8409,N_4576,N_2235);
and U8410 (N_8410,N_2651,N_1122);
nor U8411 (N_8411,N_188,N_1894);
and U8412 (N_8412,N_4503,N_2984);
and U8413 (N_8413,N_3375,N_4539);
nand U8414 (N_8414,N_4095,N_3709);
and U8415 (N_8415,N_612,N_2661);
or U8416 (N_8416,N_3891,N_4680);
xnor U8417 (N_8417,N_767,N_1974);
nand U8418 (N_8418,N_219,N_133);
and U8419 (N_8419,N_4766,N_4228);
nand U8420 (N_8420,N_1262,N_3513);
or U8421 (N_8421,N_4937,N_3553);
or U8422 (N_8422,N_3895,N_4870);
and U8423 (N_8423,N_1386,N_4249);
xnor U8424 (N_8424,N_498,N_4277);
or U8425 (N_8425,N_3935,N_3293);
and U8426 (N_8426,N_2661,N_4307);
and U8427 (N_8427,N_1282,N_4117);
or U8428 (N_8428,N_293,N_3560);
and U8429 (N_8429,N_2656,N_1230);
or U8430 (N_8430,N_2374,N_3464);
nor U8431 (N_8431,N_4925,N_1510);
or U8432 (N_8432,N_1617,N_2425);
or U8433 (N_8433,N_624,N_4994);
nor U8434 (N_8434,N_772,N_1948);
nor U8435 (N_8435,N_118,N_3035);
and U8436 (N_8436,N_1653,N_4189);
xnor U8437 (N_8437,N_3115,N_744);
xnor U8438 (N_8438,N_440,N_2641);
nor U8439 (N_8439,N_2471,N_711);
nand U8440 (N_8440,N_1179,N_3798);
nor U8441 (N_8441,N_2274,N_4486);
nor U8442 (N_8442,N_3757,N_2372);
or U8443 (N_8443,N_823,N_1273);
xor U8444 (N_8444,N_3111,N_4932);
nand U8445 (N_8445,N_3271,N_739);
nor U8446 (N_8446,N_4795,N_2442);
or U8447 (N_8447,N_741,N_3994);
nor U8448 (N_8448,N_3292,N_3800);
xor U8449 (N_8449,N_928,N_789);
nor U8450 (N_8450,N_4260,N_413);
or U8451 (N_8451,N_371,N_743);
nor U8452 (N_8452,N_4363,N_4898);
or U8453 (N_8453,N_4227,N_4936);
or U8454 (N_8454,N_4585,N_4318);
or U8455 (N_8455,N_2798,N_3592);
nand U8456 (N_8456,N_4857,N_3617);
or U8457 (N_8457,N_2070,N_3203);
nor U8458 (N_8458,N_1136,N_2331);
or U8459 (N_8459,N_1256,N_4708);
nor U8460 (N_8460,N_4131,N_4252);
and U8461 (N_8461,N_2930,N_4622);
or U8462 (N_8462,N_617,N_1596);
nor U8463 (N_8463,N_1514,N_3371);
xor U8464 (N_8464,N_2985,N_2070);
xor U8465 (N_8465,N_2116,N_717);
nand U8466 (N_8466,N_1534,N_2855);
or U8467 (N_8467,N_2178,N_3131);
nor U8468 (N_8468,N_875,N_1034);
and U8469 (N_8469,N_2843,N_747);
xnor U8470 (N_8470,N_4457,N_3214);
nor U8471 (N_8471,N_2742,N_4233);
xnor U8472 (N_8472,N_2371,N_1320);
and U8473 (N_8473,N_2203,N_2492);
nor U8474 (N_8474,N_2196,N_3434);
or U8475 (N_8475,N_1523,N_653);
nand U8476 (N_8476,N_4389,N_4957);
xnor U8477 (N_8477,N_3026,N_2715);
nand U8478 (N_8478,N_35,N_837);
nand U8479 (N_8479,N_1044,N_3676);
or U8480 (N_8480,N_1742,N_3504);
nor U8481 (N_8481,N_4248,N_848);
xnor U8482 (N_8482,N_2401,N_3675);
and U8483 (N_8483,N_401,N_2845);
or U8484 (N_8484,N_836,N_1600);
xor U8485 (N_8485,N_695,N_4814);
nor U8486 (N_8486,N_3633,N_2137);
nor U8487 (N_8487,N_2596,N_1762);
or U8488 (N_8488,N_3399,N_2068);
nand U8489 (N_8489,N_4813,N_2928);
and U8490 (N_8490,N_3244,N_968);
nand U8491 (N_8491,N_2113,N_4113);
and U8492 (N_8492,N_918,N_3419);
or U8493 (N_8493,N_3503,N_4041);
nand U8494 (N_8494,N_3432,N_4742);
nand U8495 (N_8495,N_1758,N_1644);
nor U8496 (N_8496,N_3906,N_4973);
nand U8497 (N_8497,N_2629,N_2910);
or U8498 (N_8498,N_1764,N_3261);
nor U8499 (N_8499,N_1917,N_2058);
nor U8500 (N_8500,N_3850,N_4123);
nand U8501 (N_8501,N_4366,N_604);
xnor U8502 (N_8502,N_881,N_4827);
xnor U8503 (N_8503,N_3015,N_4976);
and U8504 (N_8504,N_4137,N_2175);
xor U8505 (N_8505,N_1309,N_4575);
and U8506 (N_8506,N_2925,N_1405);
or U8507 (N_8507,N_2805,N_3772);
xor U8508 (N_8508,N_4711,N_3995);
nand U8509 (N_8509,N_4477,N_4531);
and U8510 (N_8510,N_3895,N_593);
and U8511 (N_8511,N_2659,N_1960);
or U8512 (N_8512,N_3865,N_3531);
nand U8513 (N_8513,N_2930,N_559);
or U8514 (N_8514,N_420,N_4145);
and U8515 (N_8515,N_59,N_480);
xor U8516 (N_8516,N_1322,N_24);
nor U8517 (N_8517,N_14,N_1361);
and U8518 (N_8518,N_4359,N_3415);
and U8519 (N_8519,N_3192,N_198);
or U8520 (N_8520,N_2579,N_1164);
nor U8521 (N_8521,N_4513,N_2276);
nor U8522 (N_8522,N_4437,N_1938);
or U8523 (N_8523,N_4438,N_3878);
and U8524 (N_8524,N_94,N_671);
nor U8525 (N_8525,N_3959,N_2628);
xnor U8526 (N_8526,N_2039,N_2383);
nand U8527 (N_8527,N_1647,N_4458);
or U8528 (N_8528,N_3378,N_1367);
or U8529 (N_8529,N_2013,N_922);
xnor U8530 (N_8530,N_4741,N_3196);
xor U8531 (N_8531,N_3236,N_3202);
or U8532 (N_8532,N_4053,N_1638);
or U8533 (N_8533,N_2269,N_4860);
or U8534 (N_8534,N_4316,N_71);
xnor U8535 (N_8535,N_4518,N_812);
or U8536 (N_8536,N_4534,N_278);
nor U8537 (N_8537,N_4262,N_219);
xnor U8538 (N_8538,N_2180,N_4042);
or U8539 (N_8539,N_2752,N_2658);
nand U8540 (N_8540,N_237,N_4547);
or U8541 (N_8541,N_2153,N_4262);
nor U8542 (N_8542,N_1302,N_29);
nor U8543 (N_8543,N_1227,N_3315);
and U8544 (N_8544,N_2215,N_2371);
and U8545 (N_8545,N_4111,N_3114);
nor U8546 (N_8546,N_432,N_2863);
or U8547 (N_8547,N_667,N_3501);
or U8548 (N_8548,N_1642,N_824);
and U8549 (N_8549,N_2069,N_1089);
nor U8550 (N_8550,N_2771,N_2249);
nand U8551 (N_8551,N_3025,N_4454);
or U8552 (N_8552,N_1670,N_907);
or U8553 (N_8553,N_1008,N_3160);
nand U8554 (N_8554,N_2843,N_113);
xor U8555 (N_8555,N_4300,N_4482);
nor U8556 (N_8556,N_1903,N_4815);
and U8557 (N_8557,N_2318,N_2200);
and U8558 (N_8558,N_1859,N_3238);
or U8559 (N_8559,N_1928,N_1490);
or U8560 (N_8560,N_983,N_4378);
or U8561 (N_8561,N_2580,N_1058);
nor U8562 (N_8562,N_1513,N_4532);
and U8563 (N_8563,N_4391,N_2873);
nand U8564 (N_8564,N_3599,N_55);
nor U8565 (N_8565,N_4472,N_3653);
or U8566 (N_8566,N_1715,N_4071);
nand U8567 (N_8567,N_4762,N_2759);
nand U8568 (N_8568,N_518,N_1807);
xnor U8569 (N_8569,N_1618,N_963);
xnor U8570 (N_8570,N_3083,N_73);
and U8571 (N_8571,N_1057,N_4286);
and U8572 (N_8572,N_4895,N_1077);
or U8573 (N_8573,N_2003,N_441);
nand U8574 (N_8574,N_1131,N_1729);
or U8575 (N_8575,N_4836,N_2141);
xor U8576 (N_8576,N_3781,N_4894);
nand U8577 (N_8577,N_4923,N_3355);
nor U8578 (N_8578,N_2756,N_956);
xnor U8579 (N_8579,N_2999,N_2470);
or U8580 (N_8580,N_4493,N_2911);
nor U8581 (N_8581,N_1272,N_3183);
xnor U8582 (N_8582,N_695,N_3449);
xnor U8583 (N_8583,N_236,N_285);
or U8584 (N_8584,N_3978,N_4945);
nor U8585 (N_8585,N_4854,N_1712);
or U8586 (N_8586,N_2638,N_3975);
and U8587 (N_8587,N_3616,N_3846);
and U8588 (N_8588,N_2387,N_816);
xnor U8589 (N_8589,N_4529,N_2775);
or U8590 (N_8590,N_4882,N_2442);
nor U8591 (N_8591,N_4561,N_2769);
and U8592 (N_8592,N_4199,N_2700);
and U8593 (N_8593,N_4324,N_4487);
or U8594 (N_8594,N_3912,N_1192);
xor U8595 (N_8595,N_4086,N_2212);
nand U8596 (N_8596,N_3,N_4521);
xor U8597 (N_8597,N_2932,N_3775);
or U8598 (N_8598,N_1673,N_691);
nand U8599 (N_8599,N_2704,N_1671);
or U8600 (N_8600,N_4024,N_547);
and U8601 (N_8601,N_1285,N_3717);
or U8602 (N_8602,N_1324,N_838);
nand U8603 (N_8603,N_443,N_2270);
xor U8604 (N_8604,N_852,N_2799);
and U8605 (N_8605,N_2514,N_488);
xor U8606 (N_8606,N_998,N_3710);
nand U8607 (N_8607,N_410,N_2446);
nor U8608 (N_8608,N_30,N_3270);
or U8609 (N_8609,N_3030,N_3523);
nor U8610 (N_8610,N_1228,N_3059);
nor U8611 (N_8611,N_4356,N_4441);
xnor U8612 (N_8612,N_3771,N_4703);
or U8613 (N_8613,N_3994,N_2365);
or U8614 (N_8614,N_1522,N_35);
and U8615 (N_8615,N_1666,N_1158);
nor U8616 (N_8616,N_548,N_2340);
xor U8617 (N_8617,N_3387,N_4757);
xnor U8618 (N_8618,N_4114,N_1347);
and U8619 (N_8619,N_1588,N_4788);
nor U8620 (N_8620,N_1518,N_3076);
nor U8621 (N_8621,N_1096,N_1333);
nor U8622 (N_8622,N_370,N_3983);
and U8623 (N_8623,N_572,N_2740);
or U8624 (N_8624,N_900,N_3592);
nor U8625 (N_8625,N_4366,N_742);
and U8626 (N_8626,N_4899,N_1028);
xnor U8627 (N_8627,N_3918,N_3898);
and U8628 (N_8628,N_3321,N_3539);
nor U8629 (N_8629,N_1730,N_3908);
or U8630 (N_8630,N_1173,N_1368);
xnor U8631 (N_8631,N_1840,N_2887);
nand U8632 (N_8632,N_1076,N_2143);
and U8633 (N_8633,N_138,N_2108);
or U8634 (N_8634,N_4199,N_2029);
or U8635 (N_8635,N_4790,N_4410);
or U8636 (N_8636,N_1296,N_459);
nand U8637 (N_8637,N_779,N_2072);
xnor U8638 (N_8638,N_4071,N_558);
or U8639 (N_8639,N_2970,N_4282);
nand U8640 (N_8640,N_3962,N_2124);
nand U8641 (N_8641,N_2092,N_4558);
xor U8642 (N_8642,N_3727,N_549);
or U8643 (N_8643,N_3481,N_2520);
nand U8644 (N_8644,N_3224,N_1730);
nand U8645 (N_8645,N_4535,N_2426);
xnor U8646 (N_8646,N_4154,N_492);
nand U8647 (N_8647,N_980,N_1293);
nor U8648 (N_8648,N_3280,N_3364);
or U8649 (N_8649,N_4600,N_79);
and U8650 (N_8650,N_4390,N_3625);
and U8651 (N_8651,N_4502,N_4534);
nor U8652 (N_8652,N_1769,N_2873);
xor U8653 (N_8653,N_4195,N_158);
and U8654 (N_8654,N_1330,N_2063);
nand U8655 (N_8655,N_2016,N_802);
xnor U8656 (N_8656,N_2044,N_239);
nor U8657 (N_8657,N_2707,N_2103);
and U8658 (N_8658,N_415,N_3556);
nand U8659 (N_8659,N_1065,N_4194);
and U8660 (N_8660,N_3541,N_1083);
or U8661 (N_8661,N_647,N_4328);
nor U8662 (N_8662,N_48,N_3863);
xnor U8663 (N_8663,N_4887,N_2916);
nor U8664 (N_8664,N_389,N_1630);
xnor U8665 (N_8665,N_1733,N_812);
xor U8666 (N_8666,N_981,N_1363);
or U8667 (N_8667,N_4638,N_904);
nor U8668 (N_8668,N_3198,N_2653);
nand U8669 (N_8669,N_1178,N_2234);
xnor U8670 (N_8670,N_547,N_238);
xnor U8671 (N_8671,N_2733,N_1841);
xnor U8672 (N_8672,N_2854,N_2032);
xor U8673 (N_8673,N_2192,N_3157);
or U8674 (N_8674,N_987,N_2231);
or U8675 (N_8675,N_1793,N_316);
xor U8676 (N_8676,N_1528,N_45);
xor U8677 (N_8677,N_4529,N_667);
or U8678 (N_8678,N_2402,N_3604);
and U8679 (N_8679,N_366,N_52);
nor U8680 (N_8680,N_4484,N_4077);
nor U8681 (N_8681,N_3086,N_3242);
and U8682 (N_8682,N_198,N_3687);
and U8683 (N_8683,N_1673,N_2090);
and U8684 (N_8684,N_1601,N_1622);
nand U8685 (N_8685,N_3172,N_1233);
nor U8686 (N_8686,N_2685,N_2412);
or U8687 (N_8687,N_1918,N_1366);
nor U8688 (N_8688,N_4939,N_3196);
nor U8689 (N_8689,N_4515,N_952);
nand U8690 (N_8690,N_2292,N_4608);
xnor U8691 (N_8691,N_3206,N_2203);
nor U8692 (N_8692,N_187,N_1450);
or U8693 (N_8693,N_3307,N_1469);
nor U8694 (N_8694,N_4095,N_2259);
xnor U8695 (N_8695,N_2879,N_2626);
nor U8696 (N_8696,N_4691,N_641);
nand U8697 (N_8697,N_3979,N_1254);
and U8698 (N_8698,N_88,N_2880);
xor U8699 (N_8699,N_2994,N_3822);
or U8700 (N_8700,N_3810,N_2727);
and U8701 (N_8701,N_2528,N_53);
nor U8702 (N_8702,N_3979,N_1693);
xnor U8703 (N_8703,N_765,N_2305);
nor U8704 (N_8704,N_1371,N_3126);
and U8705 (N_8705,N_1854,N_2492);
nand U8706 (N_8706,N_1401,N_4476);
or U8707 (N_8707,N_301,N_4197);
xnor U8708 (N_8708,N_846,N_4363);
or U8709 (N_8709,N_2628,N_1702);
nand U8710 (N_8710,N_4743,N_689);
xnor U8711 (N_8711,N_1084,N_4018);
nand U8712 (N_8712,N_1498,N_2240);
xor U8713 (N_8713,N_199,N_2073);
nand U8714 (N_8714,N_264,N_842);
nor U8715 (N_8715,N_3713,N_1251);
and U8716 (N_8716,N_788,N_283);
nand U8717 (N_8717,N_2472,N_2948);
xor U8718 (N_8718,N_400,N_2175);
nor U8719 (N_8719,N_1587,N_3188);
xnor U8720 (N_8720,N_4025,N_3220);
xnor U8721 (N_8721,N_460,N_4382);
xor U8722 (N_8722,N_3045,N_920);
nand U8723 (N_8723,N_4968,N_2964);
or U8724 (N_8724,N_3052,N_1827);
xnor U8725 (N_8725,N_4193,N_1197);
or U8726 (N_8726,N_3082,N_4214);
and U8727 (N_8727,N_3140,N_3011);
xnor U8728 (N_8728,N_4171,N_1781);
xnor U8729 (N_8729,N_3961,N_4208);
nor U8730 (N_8730,N_1767,N_2159);
and U8731 (N_8731,N_1439,N_1050);
xor U8732 (N_8732,N_1349,N_1657);
xor U8733 (N_8733,N_4372,N_660);
nor U8734 (N_8734,N_715,N_708);
or U8735 (N_8735,N_3990,N_2203);
xor U8736 (N_8736,N_115,N_1554);
xor U8737 (N_8737,N_2768,N_1092);
or U8738 (N_8738,N_4519,N_3791);
nor U8739 (N_8739,N_52,N_2792);
nand U8740 (N_8740,N_3611,N_1826);
nand U8741 (N_8741,N_3671,N_1014);
nor U8742 (N_8742,N_4187,N_4920);
nand U8743 (N_8743,N_3596,N_2339);
nand U8744 (N_8744,N_3097,N_420);
nor U8745 (N_8745,N_160,N_1934);
xor U8746 (N_8746,N_333,N_4898);
nand U8747 (N_8747,N_4111,N_105);
and U8748 (N_8748,N_3174,N_3587);
xor U8749 (N_8749,N_3089,N_3065);
or U8750 (N_8750,N_189,N_4858);
nand U8751 (N_8751,N_2359,N_214);
nor U8752 (N_8752,N_880,N_1917);
and U8753 (N_8753,N_2795,N_3926);
nand U8754 (N_8754,N_2717,N_2549);
xnor U8755 (N_8755,N_4802,N_4744);
and U8756 (N_8756,N_789,N_1399);
xor U8757 (N_8757,N_4363,N_3605);
or U8758 (N_8758,N_2392,N_3977);
xnor U8759 (N_8759,N_3392,N_2790);
and U8760 (N_8760,N_473,N_1584);
or U8761 (N_8761,N_760,N_789);
or U8762 (N_8762,N_1630,N_1247);
and U8763 (N_8763,N_1583,N_1294);
or U8764 (N_8764,N_3171,N_2016);
or U8765 (N_8765,N_1247,N_4326);
or U8766 (N_8766,N_1366,N_3879);
xor U8767 (N_8767,N_1730,N_3517);
nand U8768 (N_8768,N_4625,N_4824);
and U8769 (N_8769,N_3909,N_1577);
xor U8770 (N_8770,N_2050,N_1983);
xor U8771 (N_8771,N_1332,N_4850);
and U8772 (N_8772,N_2148,N_4348);
or U8773 (N_8773,N_3231,N_1285);
and U8774 (N_8774,N_298,N_3961);
xnor U8775 (N_8775,N_488,N_4146);
nand U8776 (N_8776,N_2755,N_4336);
xor U8777 (N_8777,N_4715,N_62);
or U8778 (N_8778,N_3049,N_3979);
xor U8779 (N_8779,N_1773,N_653);
and U8780 (N_8780,N_3017,N_398);
and U8781 (N_8781,N_4068,N_2606);
nand U8782 (N_8782,N_3673,N_3932);
nor U8783 (N_8783,N_1149,N_3814);
nand U8784 (N_8784,N_4679,N_690);
nand U8785 (N_8785,N_2837,N_2936);
nor U8786 (N_8786,N_744,N_3686);
nand U8787 (N_8787,N_2929,N_4651);
or U8788 (N_8788,N_4260,N_3075);
xnor U8789 (N_8789,N_2825,N_4758);
nand U8790 (N_8790,N_1864,N_3517);
nand U8791 (N_8791,N_3012,N_3624);
nor U8792 (N_8792,N_3928,N_4379);
or U8793 (N_8793,N_4150,N_4722);
nand U8794 (N_8794,N_2550,N_4465);
or U8795 (N_8795,N_1963,N_4375);
and U8796 (N_8796,N_1585,N_3433);
nand U8797 (N_8797,N_3757,N_3471);
xor U8798 (N_8798,N_461,N_2638);
nor U8799 (N_8799,N_3890,N_820);
or U8800 (N_8800,N_4662,N_4369);
nor U8801 (N_8801,N_2343,N_2365);
and U8802 (N_8802,N_288,N_2479);
nor U8803 (N_8803,N_2687,N_443);
and U8804 (N_8804,N_3377,N_2526);
nor U8805 (N_8805,N_547,N_700);
and U8806 (N_8806,N_3569,N_3299);
and U8807 (N_8807,N_921,N_2666);
nand U8808 (N_8808,N_372,N_4244);
and U8809 (N_8809,N_2221,N_1233);
or U8810 (N_8810,N_3089,N_3248);
and U8811 (N_8811,N_1461,N_2465);
nand U8812 (N_8812,N_1851,N_2150);
nand U8813 (N_8813,N_4818,N_975);
nand U8814 (N_8814,N_4795,N_971);
xnor U8815 (N_8815,N_3485,N_4278);
and U8816 (N_8816,N_1279,N_609);
or U8817 (N_8817,N_141,N_2992);
xor U8818 (N_8818,N_0,N_143);
and U8819 (N_8819,N_4265,N_1301);
or U8820 (N_8820,N_3347,N_4374);
nor U8821 (N_8821,N_1838,N_1448);
nor U8822 (N_8822,N_2341,N_1283);
or U8823 (N_8823,N_353,N_3450);
and U8824 (N_8824,N_4487,N_3112);
xor U8825 (N_8825,N_4873,N_462);
nor U8826 (N_8826,N_3052,N_3089);
and U8827 (N_8827,N_584,N_4697);
or U8828 (N_8828,N_2209,N_3312);
nor U8829 (N_8829,N_4090,N_2444);
nor U8830 (N_8830,N_4595,N_48);
and U8831 (N_8831,N_2936,N_887);
nand U8832 (N_8832,N_1043,N_928);
and U8833 (N_8833,N_45,N_2157);
nand U8834 (N_8834,N_1818,N_1447);
nor U8835 (N_8835,N_4267,N_3049);
xor U8836 (N_8836,N_4269,N_2109);
xor U8837 (N_8837,N_988,N_584);
xor U8838 (N_8838,N_2731,N_230);
and U8839 (N_8839,N_4083,N_3054);
nand U8840 (N_8840,N_4248,N_3452);
nor U8841 (N_8841,N_3101,N_4441);
nor U8842 (N_8842,N_2535,N_4780);
or U8843 (N_8843,N_2846,N_2403);
or U8844 (N_8844,N_3396,N_2933);
nor U8845 (N_8845,N_1498,N_1491);
and U8846 (N_8846,N_340,N_3197);
xnor U8847 (N_8847,N_4704,N_66);
xnor U8848 (N_8848,N_2759,N_727);
or U8849 (N_8849,N_3607,N_1558);
and U8850 (N_8850,N_1755,N_4195);
nor U8851 (N_8851,N_2333,N_623);
or U8852 (N_8852,N_1994,N_1749);
or U8853 (N_8853,N_3414,N_1876);
xnor U8854 (N_8854,N_3744,N_1809);
nand U8855 (N_8855,N_2872,N_393);
xnor U8856 (N_8856,N_1082,N_1915);
xnor U8857 (N_8857,N_4633,N_2936);
xor U8858 (N_8858,N_3940,N_263);
xnor U8859 (N_8859,N_2765,N_1893);
nand U8860 (N_8860,N_4824,N_2370);
nor U8861 (N_8861,N_2531,N_168);
xnor U8862 (N_8862,N_646,N_1197);
nor U8863 (N_8863,N_3038,N_602);
or U8864 (N_8864,N_2112,N_2101);
xor U8865 (N_8865,N_850,N_4063);
nor U8866 (N_8866,N_1471,N_4533);
and U8867 (N_8867,N_2262,N_3700);
or U8868 (N_8868,N_2656,N_3619);
or U8869 (N_8869,N_953,N_2564);
xnor U8870 (N_8870,N_749,N_3819);
nand U8871 (N_8871,N_1539,N_1030);
xor U8872 (N_8872,N_4776,N_2308);
xnor U8873 (N_8873,N_3736,N_4708);
nand U8874 (N_8874,N_1395,N_3973);
nor U8875 (N_8875,N_3271,N_3944);
or U8876 (N_8876,N_648,N_224);
nor U8877 (N_8877,N_2363,N_2555);
nand U8878 (N_8878,N_2240,N_537);
xnor U8879 (N_8879,N_2800,N_389);
or U8880 (N_8880,N_4417,N_3026);
and U8881 (N_8881,N_4421,N_2944);
nor U8882 (N_8882,N_454,N_2182);
xor U8883 (N_8883,N_327,N_85);
nor U8884 (N_8884,N_4397,N_3669);
and U8885 (N_8885,N_838,N_236);
nor U8886 (N_8886,N_3055,N_4149);
nand U8887 (N_8887,N_220,N_3885);
nand U8888 (N_8888,N_3720,N_807);
xnor U8889 (N_8889,N_3530,N_3984);
xnor U8890 (N_8890,N_3527,N_872);
or U8891 (N_8891,N_3428,N_973);
and U8892 (N_8892,N_1958,N_1702);
or U8893 (N_8893,N_4317,N_159);
xor U8894 (N_8894,N_2606,N_2469);
and U8895 (N_8895,N_2868,N_1457);
nor U8896 (N_8896,N_2741,N_2721);
nand U8897 (N_8897,N_2397,N_2806);
or U8898 (N_8898,N_1143,N_683);
and U8899 (N_8899,N_3296,N_2624);
or U8900 (N_8900,N_2595,N_1091);
xnor U8901 (N_8901,N_901,N_864);
nor U8902 (N_8902,N_3709,N_5);
xor U8903 (N_8903,N_1436,N_4507);
nor U8904 (N_8904,N_898,N_3786);
xnor U8905 (N_8905,N_154,N_2763);
and U8906 (N_8906,N_1645,N_1731);
xnor U8907 (N_8907,N_2932,N_2496);
or U8908 (N_8908,N_3782,N_1410);
xor U8909 (N_8909,N_4850,N_2672);
nor U8910 (N_8910,N_2178,N_425);
or U8911 (N_8911,N_1426,N_3800);
nand U8912 (N_8912,N_4778,N_402);
nand U8913 (N_8913,N_2884,N_3608);
xnor U8914 (N_8914,N_3849,N_2668);
or U8915 (N_8915,N_4597,N_4257);
nor U8916 (N_8916,N_3170,N_1324);
nand U8917 (N_8917,N_3862,N_4440);
and U8918 (N_8918,N_1638,N_2005);
nor U8919 (N_8919,N_1187,N_4537);
nand U8920 (N_8920,N_1749,N_1692);
nand U8921 (N_8921,N_151,N_2790);
nor U8922 (N_8922,N_2036,N_1739);
xor U8923 (N_8923,N_3435,N_3388);
nor U8924 (N_8924,N_220,N_4055);
and U8925 (N_8925,N_2879,N_276);
and U8926 (N_8926,N_665,N_769);
xnor U8927 (N_8927,N_2357,N_3783);
and U8928 (N_8928,N_4051,N_993);
xnor U8929 (N_8929,N_797,N_3118);
or U8930 (N_8930,N_1789,N_2112);
and U8931 (N_8931,N_4261,N_1607);
or U8932 (N_8932,N_1755,N_3333);
nand U8933 (N_8933,N_3413,N_2119);
nor U8934 (N_8934,N_1626,N_2918);
or U8935 (N_8935,N_2042,N_4762);
or U8936 (N_8936,N_981,N_4008);
or U8937 (N_8937,N_3260,N_2576);
nor U8938 (N_8938,N_3427,N_3147);
nor U8939 (N_8939,N_611,N_4479);
or U8940 (N_8940,N_4787,N_3222);
nand U8941 (N_8941,N_3566,N_179);
or U8942 (N_8942,N_3094,N_495);
and U8943 (N_8943,N_1321,N_2951);
and U8944 (N_8944,N_754,N_2941);
nand U8945 (N_8945,N_4240,N_560);
or U8946 (N_8946,N_911,N_4915);
and U8947 (N_8947,N_3445,N_3411);
xor U8948 (N_8948,N_2757,N_3276);
nand U8949 (N_8949,N_3684,N_2690);
nand U8950 (N_8950,N_2788,N_1755);
nand U8951 (N_8951,N_1242,N_3608);
or U8952 (N_8952,N_3572,N_1795);
and U8953 (N_8953,N_3614,N_3826);
nor U8954 (N_8954,N_1137,N_3166);
nand U8955 (N_8955,N_1374,N_4939);
nand U8956 (N_8956,N_3271,N_3433);
nor U8957 (N_8957,N_4119,N_2903);
xnor U8958 (N_8958,N_3123,N_2241);
or U8959 (N_8959,N_269,N_256);
or U8960 (N_8960,N_183,N_3064);
xor U8961 (N_8961,N_748,N_40);
nor U8962 (N_8962,N_4958,N_76);
xor U8963 (N_8963,N_1637,N_3302);
xor U8964 (N_8964,N_4994,N_2475);
nor U8965 (N_8965,N_955,N_811);
and U8966 (N_8966,N_666,N_2702);
nor U8967 (N_8967,N_1295,N_3848);
xnor U8968 (N_8968,N_4434,N_427);
nor U8969 (N_8969,N_3834,N_2354);
xor U8970 (N_8970,N_30,N_3684);
and U8971 (N_8971,N_2687,N_1009);
nand U8972 (N_8972,N_2113,N_3591);
xor U8973 (N_8973,N_43,N_605);
nor U8974 (N_8974,N_1510,N_1221);
and U8975 (N_8975,N_1863,N_2582);
nor U8976 (N_8976,N_4084,N_1143);
or U8977 (N_8977,N_4020,N_3714);
or U8978 (N_8978,N_4968,N_4087);
nor U8979 (N_8979,N_270,N_3401);
nor U8980 (N_8980,N_1655,N_2422);
nand U8981 (N_8981,N_573,N_4651);
nor U8982 (N_8982,N_4195,N_995);
or U8983 (N_8983,N_2995,N_2648);
and U8984 (N_8984,N_131,N_3268);
xnor U8985 (N_8985,N_2405,N_4445);
nand U8986 (N_8986,N_1801,N_2178);
xnor U8987 (N_8987,N_715,N_4037);
or U8988 (N_8988,N_3751,N_69);
or U8989 (N_8989,N_3578,N_3845);
and U8990 (N_8990,N_159,N_1606);
or U8991 (N_8991,N_4442,N_1353);
and U8992 (N_8992,N_2377,N_4573);
nor U8993 (N_8993,N_4995,N_3324);
nand U8994 (N_8994,N_3391,N_3821);
and U8995 (N_8995,N_2264,N_4058);
xnor U8996 (N_8996,N_267,N_531);
nand U8997 (N_8997,N_2528,N_2781);
and U8998 (N_8998,N_1524,N_2222);
nand U8999 (N_8999,N_2671,N_2185);
xnor U9000 (N_9000,N_410,N_4886);
or U9001 (N_9001,N_111,N_924);
xnor U9002 (N_9002,N_4311,N_4389);
or U9003 (N_9003,N_2714,N_4698);
nand U9004 (N_9004,N_1168,N_2601);
nand U9005 (N_9005,N_779,N_2024);
nand U9006 (N_9006,N_4749,N_868);
nor U9007 (N_9007,N_499,N_2274);
nor U9008 (N_9008,N_4874,N_4007);
or U9009 (N_9009,N_472,N_2775);
nor U9010 (N_9010,N_135,N_2125);
nor U9011 (N_9011,N_656,N_2870);
nor U9012 (N_9012,N_4252,N_722);
nand U9013 (N_9013,N_4019,N_4540);
and U9014 (N_9014,N_804,N_2738);
or U9015 (N_9015,N_2307,N_2774);
xor U9016 (N_9016,N_1322,N_3411);
nor U9017 (N_9017,N_4035,N_1979);
xor U9018 (N_9018,N_2337,N_4518);
or U9019 (N_9019,N_3038,N_1297);
or U9020 (N_9020,N_2376,N_1247);
nand U9021 (N_9021,N_4260,N_283);
xnor U9022 (N_9022,N_3917,N_2739);
or U9023 (N_9023,N_2989,N_3444);
or U9024 (N_9024,N_269,N_2995);
or U9025 (N_9025,N_1859,N_4151);
and U9026 (N_9026,N_1685,N_4495);
and U9027 (N_9027,N_1417,N_3730);
xnor U9028 (N_9028,N_3092,N_4248);
nor U9029 (N_9029,N_4108,N_1198);
nor U9030 (N_9030,N_3187,N_4815);
and U9031 (N_9031,N_2947,N_2499);
nand U9032 (N_9032,N_2877,N_1103);
nor U9033 (N_9033,N_4550,N_2819);
and U9034 (N_9034,N_624,N_2524);
nor U9035 (N_9035,N_3016,N_1295);
nand U9036 (N_9036,N_446,N_2764);
or U9037 (N_9037,N_607,N_914);
nand U9038 (N_9038,N_4429,N_3272);
xor U9039 (N_9039,N_1918,N_3018);
xor U9040 (N_9040,N_3884,N_1803);
or U9041 (N_9041,N_2381,N_999);
xnor U9042 (N_9042,N_4491,N_3467);
or U9043 (N_9043,N_4370,N_3447);
nand U9044 (N_9044,N_4216,N_180);
or U9045 (N_9045,N_1255,N_3131);
nand U9046 (N_9046,N_1045,N_4271);
nand U9047 (N_9047,N_1849,N_265);
and U9048 (N_9048,N_4353,N_4449);
xor U9049 (N_9049,N_668,N_3564);
and U9050 (N_9050,N_2421,N_3351);
or U9051 (N_9051,N_3710,N_697);
nor U9052 (N_9052,N_1991,N_3468);
xor U9053 (N_9053,N_4860,N_1028);
and U9054 (N_9054,N_2456,N_4376);
nor U9055 (N_9055,N_4417,N_4190);
or U9056 (N_9056,N_1862,N_2651);
xnor U9057 (N_9057,N_4887,N_329);
nor U9058 (N_9058,N_3341,N_4297);
nor U9059 (N_9059,N_1658,N_1551);
or U9060 (N_9060,N_2965,N_2348);
or U9061 (N_9061,N_3105,N_1335);
nor U9062 (N_9062,N_4867,N_1343);
and U9063 (N_9063,N_3861,N_4385);
nand U9064 (N_9064,N_4518,N_2401);
and U9065 (N_9065,N_3885,N_431);
and U9066 (N_9066,N_1353,N_3450);
nor U9067 (N_9067,N_432,N_3514);
xor U9068 (N_9068,N_46,N_3834);
nand U9069 (N_9069,N_2611,N_1204);
xnor U9070 (N_9070,N_1560,N_3279);
nor U9071 (N_9071,N_1027,N_245);
and U9072 (N_9072,N_4459,N_1589);
or U9073 (N_9073,N_3046,N_1418);
xnor U9074 (N_9074,N_3141,N_1109);
nand U9075 (N_9075,N_1455,N_3697);
and U9076 (N_9076,N_1015,N_3790);
xor U9077 (N_9077,N_1580,N_2850);
or U9078 (N_9078,N_1148,N_4501);
nand U9079 (N_9079,N_708,N_4505);
nand U9080 (N_9080,N_3678,N_2042);
nand U9081 (N_9081,N_2988,N_3596);
nor U9082 (N_9082,N_3786,N_831);
nor U9083 (N_9083,N_1111,N_2988);
and U9084 (N_9084,N_4447,N_2164);
and U9085 (N_9085,N_4724,N_3434);
xor U9086 (N_9086,N_1187,N_1911);
xor U9087 (N_9087,N_2266,N_3050);
nor U9088 (N_9088,N_2705,N_3955);
or U9089 (N_9089,N_2318,N_2412);
and U9090 (N_9090,N_2755,N_2495);
or U9091 (N_9091,N_1182,N_1056);
xor U9092 (N_9092,N_4672,N_2480);
and U9093 (N_9093,N_2629,N_3464);
or U9094 (N_9094,N_1691,N_4028);
and U9095 (N_9095,N_2966,N_1485);
xor U9096 (N_9096,N_2201,N_807);
nor U9097 (N_9097,N_730,N_259);
or U9098 (N_9098,N_4620,N_3113);
and U9099 (N_9099,N_528,N_2949);
nor U9100 (N_9100,N_2844,N_4445);
or U9101 (N_9101,N_496,N_1445);
xor U9102 (N_9102,N_3553,N_3672);
and U9103 (N_9103,N_415,N_2381);
nand U9104 (N_9104,N_3725,N_3337);
xnor U9105 (N_9105,N_1507,N_4017);
and U9106 (N_9106,N_876,N_3096);
nor U9107 (N_9107,N_3017,N_4531);
nor U9108 (N_9108,N_4831,N_3513);
nand U9109 (N_9109,N_2889,N_792);
xor U9110 (N_9110,N_3745,N_1100);
or U9111 (N_9111,N_4857,N_1698);
nor U9112 (N_9112,N_911,N_1143);
or U9113 (N_9113,N_3600,N_580);
and U9114 (N_9114,N_1132,N_715);
nor U9115 (N_9115,N_2549,N_4639);
xnor U9116 (N_9116,N_2206,N_3996);
and U9117 (N_9117,N_1170,N_3485);
nand U9118 (N_9118,N_1607,N_3922);
nor U9119 (N_9119,N_1427,N_3933);
and U9120 (N_9120,N_3451,N_4729);
nand U9121 (N_9121,N_1674,N_3210);
and U9122 (N_9122,N_3966,N_4791);
and U9123 (N_9123,N_649,N_3704);
or U9124 (N_9124,N_300,N_3493);
nand U9125 (N_9125,N_3431,N_4236);
nand U9126 (N_9126,N_3128,N_234);
nor U9127 (N_9127,N_139,N_1418);
and U9128 (N_9128,N_1512,N_2532);
nand U9129 (N_9129,N_2105,N_768);
nor U9130 (N_9130,N_2407,N_4910);
nand U9131 (N_9131,N_1356,N_1241);
nand U9132 (N_9132,N_4469,N_4574);
nand U9133 (N_9133,N_4951,N_1943);
xor U9134 (N_9134,N_3982,N_334);
nand U9135 (N_9135,N_1047,N_777);
and U9136 (N_9136,N_1779,N_177);
xnor U9137 (N_9137,N_2333,N_3475);
and U9138 (N_9138,N_126,N_334);
and U9139 (N_9139,N_3669,N_4447);
xnor U9140 (N_9140,N_4841,N_3192);
nand U9141 (N_9141,N_4912,N_3486);
and U9142 (N_9142,N_3847,N_4219);
or U9143 (N_9143,N_1018,N_3424);
and U9144 (N_9144,N_4071,N_1707);
xor U9145 (N_9145,N_3328,N_2247);
or U9146 (N_9146,N_1712,N_63);
and U9147 (N_9147,N_2540,N_3968);
nor U9148 (N_9148,N_230,N_1613);
nand U9149 (N_9149,N_3464,N_1480);
and U9150 (N_9150,N_148,N_4955);
nor U9151 (N_9151,N_1629,N_3591);
nor U9152 (N_9152,N_2933,N_2861);
nand U9153 (N_9153,N_2717,N_2859);
and U9154 (N_9154,N_3677,N_4005);
and U9155 (N_9155,N_58,N_2765);
xor U9156 (N_9156,N_3080,N_448);
xor U9157 (N_9157,N_354,N_642);
and U9158 (N_9158,N_415,N_1102);
nor U9159 (N_9159,N_4539,N_551);
nand U9160 (N_9160,N_4492,N_4698);
nor U9161 (N_9161,N_3078,N_4782);
and U9162 (N_9162,N_181,N_4022);
and U9163 (N_9163,N_4235,N_2965);
or U9164 (N_9164,N_2464,N_1840);
nor U9165 (N_9165,N_4139,N_3312);
nor U9166 (N_9166,N_2240,N_4303);
or U9167 (N_9167,N_4674,N_1498);
xor U9168 (N_9168,N_130,N_724);
nand U9169 (N_9169,N_2596,N_526);
or U9170 (N_9170,N_4163,N_3845);
nand U9171 (N_9171,N_936,N_1764);
xor U9172 (N_9172,N_1832,N_2974);
nand U9173 (N_9173,N_562,N_1294);
nand U9174 (N_9174,N_4818,N_1333);
nor U9175 (N_9175,N_2812,N_2993);
and U9176 (N_9176,N_2880,N_2867);
and U9177 (N_9177,N_1881,N_4060);
nor U9178 (N_9178,N_613,N_3600);
and U9179 (N_9179,N_2350,N_2824);
or U9180 (N_9180,N_4255,N_4437);
or U9181 (N_9181,N_926,N_917);
nor U9182 (N_9182,N_261,N_1378);
and U9183 (N_9183,N_3502,N_669);
xor U9184 (N_9184,N_3204,N_4808);
xnor U9185 (N_9185,N_1755,N_3265);
nor U9186 (N_9186,N_460,N_2955);
or U9187 (N_9187,N_4863,N_149);
xor U9188 (N_9188,N_168,N_2091);
xor U9189 (N_9189,N_4706,N_566);
nand U9190 (N_9190,N_2144,N_4881);
xnor U9191 (N_9191,N_762,N_4976);
or U9192 (N_9192,N_2727,N_4859);
xor U9193 (N_9193,N_827,N_4764);
xnor U9194 (N_9194,N_872,N_463);
nor U9195 (N_9195,N_1242,N_4682);
xor U9196 (N_9196,N_4399,N_1832);
nor U9197 (N_9197,N_1917,N_4363);
xor U9198 (N_9198,N_657,N_3481);
nor U9199 (N_9199,N_3104,N_4715);
xor U9200 (N_9200,N_1788,N_522);
nand U9201 (N_9201,N_794,N_3016);
nand U9202 (N_9202,N_955,N_3988);
xor U9203 (N_9203,N_2094,N_4300);
xnor U9204 (N_9204,N_2617,N_4997);
nor U9205 (N_9205,N_4619,N_4547);
and U9206 (N_9206,N_3,N_3497);
xor U9207 (N_9207,N_2763,N_1895);
nor U9208 (N_9208,N_4876,N_2795);
or U9209 (N_9209,N_2697,N_2660);
or U9210 (N_9210,N_1254,N_3703);
nor U9211 (N_9211,N_4944,N_621);
nand U9212 (N_9212,N_1883,N_4637);
nor U9213 (N_9213,N_857,N_281);
nand U9214 (N_9214,N_380,N_2422);
xor U9215 (N_9215,N_1458,N_2171);
xnor U9216 (N_9216,N_784,N_2930);
or U9217 (N_9217,N_2604,N_2464);
xnor U9218 (N_9218,N_4530,N_1685);
or U9219 (N_9219,N_1277,N_2029);
and U9220 (N_9220,N_3476,N_727);
xor U9221 (N_9221,N_375,N_3228);
xor U9222 (N_9222,N_4332,N_3204);
or U9223 (N_9223,N_713,N_982);
nor U9224 (N_9224,N_3397,N_124);
nand U9225 (N_9225,N_3614,N_185);
xor U9226 (N_9226,N_1758,N_2031);
nor U9227 (N_9227,N_1953,N_1472);
xnor U9228 (N_9228,N_2088,N_3792);
xnor U9229 (N_9229,N_3549,N_4389);
nor U9230 (N_9230,N_3432,N_969);
xor U9231 (N_9231,N_2556,N_4353);
xor U9232 (N_9232,N_3678,N_666);
or U9233 (N_9233,N_3514,N_711);
or U9234 (N_9234,N_2038,N_768);
or U9235 (N_9235,N_2690,N_4057);
nand U9236 (N_9236,N_4934,N_2043);
and U9237 (N_9237,N_4489,N_2511);
nand U9238 (N_9238,N_2651,N_4251);
or U9239 (N_9239,N_1708,N_3650);
xor U9240 (N_9240,N_3980,N_4656);
and U9241 (N_9241,N_2633,N_1476);
nand U9242 (N_9242,N_4728,N_2375);
nor U9243 (N_9243,N_1324,N_3248);
xor U9244 (N_9244,N_4463,N_3942);
and U9245 (N_9245,N_4181,N_687);
nand U9246 (N_9246,N_3105,N_4677);
nor U9247 (N_9247,N_2102,N_95);
xnor U9248 (N_9248,N_4726,N_2863);
nand U9249 (N_9249,N_4300,N_4287);
or U9250 (N_9250,N_2846,N_695);
and U9251 (N_9251,N_2583,N_484);
nand U9252 (N_9252,N_1043,N_2927);
or U9253 (N_9253,N_1495,N_4508);
or U9254 (N_9254,N_1868,N_3172);
or U9255 (N_9255,N_3282,N_4182);
or U9256 (N_9256,N_2974,N_181);
xnor U9257 (N_9257,N_3492,N_1580);
nor U9258 (N_9258,N_4762,N_642);
xnor U9259 (N_9259,N_3678,N_3133);
nand U9260 (N_9260,N_1409,N_708);
nand U9261 (N_9261,N_1939,N_673);
xnor U9262 (N_9262,N_4023,N_2095);
nand U9263 (N_9263,N_2977,N_1225);
nor U9264 (N_9264,N_3901,N_3244);
xor U9265 (N_9265,N_2844,N_182);
xnor U9266 (N_9266,N_2960,N_258);
or U9267 (N_9267,N_4971,N_2724);
and U9268 (N_9268,N_3994,N_434);
xnor U9269 (N_9269,N_219,N_3024);
xnor U9270 (N_9270,N_61,N_3639);
and U9271 (N_9271,N_4931,N_4908);
nand U9272 (N_9272,N_3449,N_3051);
and U9273 (N_9273,N_2253,N_4573);
nand U9274 (N_9274,N_4056,N_1089);
xnor U9275 (N_9275,N_4875,N_243);
and U9276 (N_9276,N_2498,N_872);
nand U9277 (N_9277,N_753,N_3723);
xnor U9278 (N_9278,N_1557,N_1798);
nand U9279 (N_9279,N_4126,N_1982);
and U9280 (N_9280,N_1562,N_1862);
nor U9281 (N_9281,N_3967,N_2794);
and U9282 (N_9282,N_1457,N_4522);
nand U9283 (N_9283,N_2739,N_1118);
nor U9284 (N_9284,N_3170,N_2161);
and U9285 (N_9285,N_4759,N_1589);
or U9286 (N_9286,N_945,N_3961);
and U9287 (N_9287,N_817,N_2931);
or U9288 (N_9288,N_1524,N_3925);
or U9289 (N_9289,N_4964,N_1050);
or U9290 (N_9290,N_127,N_4589);
and U9291 (N_9291,N_612,N_1367);
xnor U9292 (N_9292,N_1447,N_2002);
and U9293 (N_9293,N_1927,N_3956);
and U9294 (N_9294,N_495,N_2005);
nand U9295 (N_9295,N_4217,N_2056);
or U9296 (N_9296,N_3087,N_1137);
nor U9297 (N_9297,N_1829,N_617);
or U9298 (N_9298,N_1308,N_1883);
xor U9299 (N_9299,N_4390,N_506);
or U9300 (N_9300,N_4083,N_3610);
nor U9301 (N_9301,N_4480,N_3592);
nor U9302 (N_9302,N_1565,N_2748);
xor U9303 (N_9303,N_3379,N_704);
nor U9304 (N_9304,N_2744,N_3129);
nor U9305 (N_9305,N_3510,N_1324);
nor U9306 (N_9306,N_2053,N_3702);
nand U9307 (N_9307,N_1304,N_4449);
nor U9308 (N_9308,N_3856,N_1956);
and U9309 (N_9309,N_3705,N_326);
xnor U9310 (N_9310,N_1022,N_2667);
nor U9311 (N_9311,N_543,N_1481);
and U9312 (N_9312,N_3723,N_824);
nand U9313 (N_9313,N_4628,N_1961);
and U9314 (N_9314,N_1975,N_2536);
xnor U9315 (N_9315,N_1921,N_2592);
and U9316 (N_9316,N_490,N_1314);
or U9317 (N_9317,N_583,N_2711);
and U9318 (N_9318,N_4048,N_3001);
nand U9319 (N_9319,N_4055,N_227);
nor U9320 (N_9320,N_1910,N_3623);
or U9321 (N_9321,N_1185,N_1331);
and U9322 (N_9322,N_4564,N_2230);
or U9323 (N_9323,N_3157,N_4133);
and U9324 (N_9324,N_1488,N_3878);
nor U9325 (N_9325,N_1773,N_3369);
xor U9326 (N_9326,N_4104,N_2501);
xor U9327 (N_9327,N_3714,N_2492);
nand U9328 (N_9328,N_754,N_2600);
xnor U9329 (N_9329,N_1933,N_4507);
and U9330 (N_9330,N_4694,N_164);
or U9331 (N_9331,N_3855,N_2994);
nor U9332 (N_9332,N_4356,N_2048);
xor U9333 (N_9333,N_1950,N_4440);
nor U9334 (N_9334,N_2933,N_1426);
and U9335 (N_9335,N_2430,N_4364);
xor U9336 (N_9336,N_2779,N_4343);
nor U9337 (N_9337,N_4727,N_3058);
or U9338 (N_9338,N_4906,N_2119);
xnor U9339 (N_9339,N_1730,N_4270);
xor U9340 (N_9340,N_3168,N_2065);
nand U9341 (N_9341,N_2480,N_3940);
nand U9342 (N_9342,N_765,N_3407);
nand U9343 (N_9343,N_1124,N_900);
xnor U9344 (N_9344,N_2169,N_569);
xor U9345 (N_9345,N_1056,N_1321);
nor U9346 (N_9346,N_2999,N_4226);
or U9347 (N_9347,N_3092,N_839);
or U9348 (N_9348,N_3045,N_2752);
xnor U9349 (N_9349,N_980,N_4225);
nand U9350 (N_9350,N_2551,N_4608);
or U9351 (N_9351,N_1062,N_1606);
nand U9352 (N_9352,N_4632,N_147);
or U9353 (N_9353,N_2997,N_3309);
xor U9354 (N_9354,N_3093,N_3798);
nand U9355 (N_9355,N_918,N_1398);
or U9356 (N_9356,N_3280,N_3379);
and U9357 (N_9357,N_1023,N_3074);
nor U9358 (N_9358,N_3868,N_2259);
nand U9359 (N_9359,N_654,N_3904);
nand U9360 (N_9360,N_2508,N_4079);
and U9361 (N_9361,N_808,N_4751);
and U9362 (N_9362,N_2930,N_650);
or U9363 (N_9363,N_597,N_1802);
nor U9364 (N_9364,N_929,N_3436);
and U9365 (N_9365,N_4617,N_2118);
or U9366 (N_9366,N_2777,N_4235);
xnor U9367 (N_9367,N_4038,N_4563);
xnor U9368 (N_9368,N_2582,N_2403);
or U9369 (N_9369,N_4429,N_3579);
and U9370 (N_9370,N_3292,N_1370);
nor U9371 (N_9371,N_976,N_4050);
and U9372 (N_9372,N_1642,N_4848);
xor U9373 (N_9373,N_3475,N_3585);
xnor U9374 (N_9374,N_2135,N_2608);
nand U9375 (N_9375,N_1987,N_4792);
nor U9376 (N_9376,N_2712,N_2448);
nor U9377 (N_9377,N_2827,N_932);
or U9378 (N_9378,N_137,N_3270);
and U9379 (N_9379,N_3573,N_4800);
or U9380 (N_9380,N_3617,N_663);
and U9381 (N_9381,N_678,N_857);
nand U9382 (N_9382,N_4179,N_1293);
or U9383 (N_9383,N_1844,N_2684);
xor U9384 (N_9384,N_3164,N_3317);
nor U9385 (N_9385,N_1749,N_1694);
nand U9386 (N_9386,N_4716,N_686);
xor U9387 (N_9387,N_824,N_3254);
nand U9388 (N_9388,N_2815,N_3290);
and U9389 (N_9389,N_3373,N_2162);
xnor U9390 (N_9390,N_3646,N_4128);
nand U9391 (N_9391,N_2711,N_1131);
nand U9392 (N_9392,N_4163,N_3848);
and U9393 (N_9393,N_153,N_1518);
and U9394 (N_9394,N_3355,N_229);
or U9395 (N_9395,N_2556,N_2333);
or U9396 (N_9396,N_3721,N_1213);
or U9397 (N_9397,N_245,N_4698);
nor U9398 (N_9398,N_3505,N_4024);
nor U9399 (N_9399,N_3603,N_1358);
nand U9400 (N_9400,N_4308,N_3084);
and U9401 (N_9401,N_2450,N_1332);
or U9402 (N_9402,N_1550,N_1751);
and U9403 (N_9403,N_4395,N_4319);
and U9404 (N_9404,N_4086,N_4714);
and U9405 (N_9405,N_2742,N_301);
xnor U9406 (N_9406,N_4493,N_3863);
nand U9407 (N_9407,N_3941,N_2710);
xnor U9408 (N_9408,N_266,N_2293);
nor U9409 (N_9409,N_2338,N_3943);
or U9410 (N_9410,N_1433,N_3120);
or U9411 (N_9411,N_606,N_3760);
or U9412 (N_9412,N_468,N_1958);
nor U9413 (N_9413,N_1778,N_512);
or U9414 (N_9414,N_1383,N_2476);
and U9415 (N_9415,N_491,N_3541);
and U9416 (N_9416,N_116,N_3458);
or U9417 (N_9417,N_3763,N_1774);
or U9418 (N_9418,N_2814,N_3267);
or U9419 (N_9419,N_1583,N_1176);
nor U9420 (N_9420,N_3129,N_1006);
nand U9421 (N_9421,N_2072,N_2834);
or U9422 (N_9422,N_4384,N_1276);
xor U9423 (N_9423,N_1819,N_3104);
and U9424 (N_9424,N_772,N_4538);
nand U9425 (N_9425,N_2641,N_3452);
and U9426 (N_9426,N_4898,N_4664);
nor U9427 (N_9427,N_1104,N_666);
or U9428 (N_9428,N_636,N_1835);
nor U9429 (N_9429,N_954,N_563);
nor U9430 (N_9430,N_1221,N_4896);
nor U9431 (N_9431,N_488,N_184);
and U9432 (N_9432,N_1173,N_1913);
xnor U9433 (N_9433,N_2837,N_2168);
or U9434 (N_9434,N_3497,N_2433);
nor U9435 (N_9435,N_4395,N_1247);
and U9436 (N_9436,N_2246,N_1243);
and U9437 (N_9437,N_2071,N_3001);
xnor U9438 (N_9438,N_1871,N_913);
nor U9439 (N_9439,N_4642,N_1522);
and U9440 (N_9440,N_3321,N_592);
xnor U9441 (N_9441,N_1562,N_2703);
and U9442 (N_9442,N_4110,N_3249);
or U9443 (N_9443,N_1228,N_1746);
nand U9444 (N_9444,N_4682,N_298);
nand U9445 (N_9445,N_2168,N_2865);
and U9446 (N_9446,N_2327,N_2495);
and U9447 (N_9447,N_3255,N_1631);
xnor U9448 (N_9448,N_3134,N_662);
nand U9449 (N_9449,N_3172,N_3776);
nand U9450 (N_9450,N_878,N_3858);
nand U9451 (N_9451,N_178,N_3897);
and U9452 (N_9452,N_4866,N_4993);
nor U9453 (N_9453,N_499,N_1019);
xor U9454 (N_9454,N_1296,N_4304);
nand U9455 (N_9455,N_1048,N_4339);
nor U9456 (N_9456,N_3203,N_323);
xor U9457 (N_9457,N_4636,N_2461);
or U9458 (N_9458,N_2250,N_3110);
or U9459 (N_9459,N_2612,N_3300);
or U9460 (N_9460,N_2180,N_2638);
xor U9461 (N_9461,N_4549,N_3721);
or U9462 (N_9462,N_969,N_4621);
nor U9463 (N_9463,N_1965,N_2487);
nand U9464 (N_9464,N_4059,N_871);
or U9465 (N_9465,N_3178,N_2758);
or U9466 (N_9466,N_9,N_1493);
or U9467 (N_9467,N_4946,N_861);
and U9468 (N_9468,N_3449,N_4573);
nand U9469 (N_9469,N_4007,N_166);
or U9470 (N_9470,N_4908,N_3660);
nor U9471 (N_9471,N_1838,N_3458);
and U9472 (N_9472,N_1462,N_4370);
nor U9473 (N_9473,N_2645,N_2634);
and U9474 (N_9474,N_2874,N_1538);
or U9475 (N_9475,N_3656,N_4854);
nor U9476 (N_9476,N_911,N_68);
xnor U9477 (N_9477,N_4646,N_1819);
nor U9478 (N_9478,N_3083,N_3718);
xnor U9479 (N_9479,N_4378,N_3753);
or U9480 (N_9480,N_1625,N_3886);
xor U9481 (N_9481,N_124,N_3776);
and U9482 (N_9482,N_4169,N_3402);
or U9483 (N_9483,N_4754,N_979);
or U9484 (N_9484,N_113,N_1183);
nand U9485 (N_9485,N_794,N_947);
nand U9486 (N_9486,N_3230,N_4861);
xor U9487 (N_9487,N_3217,N_580);
nor U9488 (N_9488,N_1040,N_47);
or U9489 (N_9489,N_2003,N_2866);
nand U9490 (N_9490,N_3323,N_3912);
xor U9491 (N_9491,N_3687,N_1977);
xor U9492 (N_9492,N_2368,N_1362);
or U9493 (N_9493,N_2170,N_2062);
or U9494 (N_9494,N_2712,N_2268);
nor U9495 (N_9495,N_4082,N_577);
nor U9496 (N_9496,N_4037,N_4537);
and U9497 (N_9497,N_1830,N_3043);
xor U9498 (N_9498,N_1282,N_1206);
nand U9499 (N_9499,N_1541,N_2667);
and U9500 (N_9500,N_2836,N_2056);
nand U9501 (N_9501,N_3573,N_4270);
nand U9502 (N_9502,N_1868,N_596);
xor U9503 (N_9503,N_193,N_4274);
or U9504 (N_9504,N_2407,N_4381);
and U9505 (N_9505,N_1158,N_3615);
and U9506 (N_9506,N_4407,N_1124);
nand U9507 (N_9507,N_2176,N_4146);
and U9508 (N_9508,N_4266,N_1347);
or U9509 (N_9509,N_4173,N_3870);
nand U9510 (N_9510,N_1718,N_3779);
nand U9511 (N_9511,N_1540,N_2818);
nor U9512 (N_9512,N_4014,N_1915);
nor U9513 (N_9513,N_3801,N_4260);
nor U9514 (N_9514,N_1286,N_3382);
nor U9515 (N_9515,N_620,N_2646);
xnor U9516 (N_9516,N_4693,N_4380);
or U9517 (N_9517,N_321,N_1610);
and U9518 (N_9518,N_3024,N_1845);
nor U9519 (N_9519,N_2864,N_3909);
and U9520 (N_9520,N_2309,N_2824);
nor U9521 (N_9521,N_2441,N_1288);
or U9522 (N_9522,N_3235,N_3218);
or U9523 (N_9523,N_1140,N_2935);
xor U9524 (N_9524,N_1892,N_1716);
and U9525 (N_9525,N_2310,N_269);
nor U9526 (N_9526,N_3219,N_4381);
or U9527 (N_9527,N_1751,N_2266);
or U9528 (N_9528,N_2029,N_2177);
or U9529 (N_9529,N_3579,N_4642);
nor U9530 (N_9530,N_1782,N_147);
xor U9531 (N_9531,N_4511,N_4507);
xnor U9532 (N_9532,N_4840,N_1238);
nand U9533 (N_9533,N_1988,N_1229);
or U9534 (N_9534,N_2681,N_493);
or U9535 (N_9535,N_1180,N_2339);
nor U9536 (N_9536,N_3694,N_4169);
nor U9537 (N_9537,N_497,N_1493);
nor U9538 (N_9538,N_4429,N_4260);
and U9539 (N_9539,N_3125,N_2162);
or U9540 (N_9540,N_292,N_3666);
or U9541 (N_9541,N_1607,N_1673);
xor U9542 (N_9542,N_2011,N_4271);
nor U9543 (N_9543,N_2106,N_14);
nor U9544 (N_9544,N_2863,N_3011);
and U9545 (N_9545,N_1634,N_363);
or U9546 (N_9546,N_3745,N_3412);
and U9547 (N_9547,N_971,N_3256);
nand U9548 (N_9548,N_4309,N_3182);
nor U9549 (N_9549,N_765,N_1790);
nand U9550 (N_9550,N_4171,N_2845);
xor U9551 (N_9551,N_3641,N_2250);
nand U9552 (N_9552,N_3452,N_1431);
nand U9553 (N_9553,N_1766,N_2778);
or U9554 (N_9554,N_2225,N_1866);
and U9555 (N_9555,N_2922,N_1265);
nor U9556 (N_9556,N_2597,N_2114);
and U9557 (N_9557,N_392,N_4712);
nor U9558 (N_9558,N_3869,N_1640);
nand U9559 (N_9559,N_1538,N_240);
xnor U9560 (N_9560,N_2557,N_3956);
xor U9561 (N_9561,N_3125,N_3594);
nor U9562 (N_9562,N_3649,N_3212);
nor U9563 (N_9563,N_2375,N_4179);
or U9564 (N_9564,N_1007,N_1608);
and U9565 (N_9565,N_771,N_4506);
and U9566 (N_9566,N_1479,N_2882);
or U9567 (N_9567,N_3608,N_4615);
or U9568 (N_9568,N_4499,N_1438);
nand U9569 (N_9569,N_4258,N_2555);
nor U9570 (N_9570,N_2591,N_437);
nand U9571 (N_9571,N_4209,N_1160);
or U9572 (N_9572,N_4374,N_982);
xnor U9573 (N_9573,N_921,N_1901);
or U9574 (N_9574,N_1458,N_1928);
and U9575 (N_9575,N_604,N_2455);
or U9576 (N_9576,N_3729,N_3141);
nand U9577 (N_9577,N_2138,N_430);
nor U9578 (N_9578,N_4572,N_1634);
and U9579 (N_9579,N_2891,N_3526);
and U9580 (N_9580,N_2844,N_369);
nor U9581 (N_9581,N_839,N_2698);
and U9582 (N_9582,N_3767,N_3793);
or U9583 (N_9583,N_2253,N_1400);
nand U9584 (N_9584,N_2124,N_4244);
and U9585 (N_9585,N_2148,N_945);
and U9586 (N_9586,N_1835,N_1709);
xnor U9587 (N_9587,N_3096,N_118);
nor U9588 (N_9588,N_4741,N_1012);
nand U9589 (N_9589,N_1774,N_4015);
or U9590 (N_9590,N_871,N_4379);
nor U9591 (N_9591,N_2874,N_2497);
or U9592 (N_9592,N_3232,N_1207);
nand U9593 (N_9593,N_464,N_2183);
or U9594 (N_9594,N_376,N_3808);
and U9595 (N_9595,N_3078,N_2168);
and U9596 (N_9596,N_3344,N_626);
nand U9597 (N_9597,N_1230,N_3050);
nor U9598 (N_9598,N_4982,N_3664);
nor U9599 (N_9599,N_2556,N_1902);
and U9600 (N_9600,N_4091,N_3559);
and U9601 (N_9601,N_986,N_2547);
or U9602 (N_9602,N_3709,N_2533);
and U9603 (N_9603,N_4269,N_1728);
nor U9604 (N_9604,N_4800,N_1056);
nand U9605 (N_9605,N_4109,N_2368);
nand U9606 (N_9606,N_2580,N_663);
nand U9607 (N_9607,N_14,N_4142);
nor U9608 (N_9608,N_4752,N_3545);
nand U9609 (N_9609,N_3178,N_1282);
nand U9610 (N_9610,N_1383,N_3476);
nand U9611 (N_9611,N_2839,N_3387);
or U9612 (N_9612,N_86,N_2773);
nor U9613 (N_9613,N_1798,N_1300);
xor U9614 (N_9614,N_2691,N_2232);
nor U9615 (N_9615,N_1777,N_4406);
nor U9616 (N_9616,N_749,N_841);
and U9617 (N_9617,N_1442,N_710);
xnor U9618 (N_9618,N_2789,N_503);
xor U9619 (N_9619,N_3598,N_4893);
nand U9620 (N_9620,N_4207,N_539);
or U9621 (N_9621,N_909,N_1403);
nor U9622 (N_9622,N_3856,N_4757);
xor U9623 (N_9623,N_1385,N_2893);
xnor U9624 (N_9624,N_3401,N_3875);
and U9625 (N_9625,N_2090,N_479);
and U9626 (N_9626,N_2509,N_1814);
nor U9627 (N_9627,N_666,N_2073);
xor U9628 (N_9628,N_2269,N_2328);
or U9629 (N_9629,N_2075,N_2566);
xnor U9630 (N_9630,N_3339,N_834);
and U9631 (N_9631,N_2134,N_1229);
xnor U9632 (N_9632,N_1422,N_4309);
and U9633 (N_9633,N_3388,N_4140);
and U9634 (N_9634,N_1467,N_3574);
nand U9635 (N_9635,N_1640,N_2822);
and U9636 (N_9636,N_4480,N_4319);
nor U9637 (N_9637,N_443,N_4739);
and U9638 (N_9638,N_1643,N_3156);
nor U9639 (N_9639,N_717,N_3110);
nor U9640 (N_9640,N_3441,N_2375);
and U9641 (N_9641,N_2783,N_4222);
xor U9642 (N_9642,N_458,N_2918);
and U9643 (N_9643,N_2915,N_582);
xnor U9644 (N_9644,N_2203,N_2777);
nand U9645 (N_9645,N_3646,N_4617);
nand U9646 (N_9646,N_2225,N_3208);
nor U9647 (N_9647,N_2290,N_3284);
nand U9648 (N_9648,N_3598,N_4574);
or U9649 (N_9649,N_2219,N_4710);
nand U9650 (N_9650,N_1969,N_2654);
nor U9651 (N_9651,N_4459,N_2497);
or U9652 (N_9652,N_1326,N_2983);
xor U9653 (N_9653,N_2514,N_2146);
and U9654 (N_9654,N_4483,N_2346);
nand U9655 (N_9655,N_1910,N_1917);
nor U9656 (N_9656,N_3402,N_1826);
nor U9657 (N_9657,N_1183,N_1859);
nor U9658 (N_9658,N_2709,N_695);
and U9659 (N_9659,N_1660,N_2895);
nand U9660 (N_9660,N_1112,N_2699);
and U9661 (N_9661,N_4699,N_1981);
xnor U9662 (N_9662,N_2493,N_1130);
nor U9663 (N_9663,N_4770,N_3843);
nand U9664 (N_9664,N_4411,N_384);
xor U9665 (N_9665,N_1127,N_4338);
and U9666 (N_9666,N_935,N_786);
nor U9667 (N_9667,N_436,N_2767);
or U9668 (N_9668,N_4963,N_436);
and U9669 (N_9669,N_703,N_3886);
xnor U9670 (N_9670,N_1227,N_3807);
nand U9671 (N_9671,N_10,N_1147);
nor U9672 (N_9672,N_1072,N_2169);
or U9673 (N_9673,N_1810,N_2405);
or U9674 (N_9674,N_4673,N_859);
or U9675 (N_9675,N_4573,N_4005);
nand U9676 (N_9676,N_1591,N_4967);
nand U9677 (N_9677,N_3269,N_1571);
xnor U9678 (N_9678,N_796,N_691);
and U9679 (N_9679,N_418,N_3823);
and U9680 (N_9680,N_248,N_2370);
nor U9681 (N_9681,N_3869,N_4702);
nand U9682 (N_9682,N_3909,N_1389);
and U9683 (N_9683,N_2149,N_1818);
or U9684 (N_9684,N_147,N_4809);
or U9685 (N_9685,N_3395,N_4883);
xnor U9686 (N_9686,N_1140,N_4731);
nor U9687 (N_9687,N_1728,N_154);
xnor U9688 (N_9688,N_3546,N_755);
and U9689 (N_9689,N_3788,N_1789);
nor U9690 (N_9690,N_1464,N_2282);
nor U9691 (N_9691,N_1315,N_2735);
and U9692 (N_9692,N_2766,N_1056);
nor U9693 (N_9693,N_1440,N_2415);
and U9694 (N_9694,N_1949,N_4325);
or U9695 (N_9695,N_4028,N_3502);
and U9696 (N_9696,N_3838,N_2850);
xor U9697 (N_9697,N_4573,N_868);
and U9698 (N_9698,N_1959,N_751);
xor U9699 (N_9699,N_4302,N_2247);
nor U9700 (N_9700,N_1903,N_3364);
nand U9701 (N_9701,N_1822,N_2009);
xnor U9702 (N_9702,N_3295,N_1567);
and U9703 (N_9703,N_1836,N_1444);
and U9704 (N_9704,N_1876,N_3087);
xor U9705 (N_9705,N_2518,N_2176);
and U9706 (N_9706,N_3855,N_708);
nand U9707 (N_9707,N_2012,N_564);
xor U9708 (N_9708,N_3462,N_4485);
and U9709 (N_9709,N_2010,N_586);
or U9710 (N_9710,N_2584,N_4248);
nand U9711 (N_9711,N_1332,N_4535);
xnor U9712 (N_9712,N_2520,N_3779);
nor U9713 (N_9713,N_4923,N_3082);
and U9714 (N_9714,N_3307,N_1425);
or U9715 (N_9715,N_1333,N_824);
and U9716 (N_9716,N_4281,N_3835);
xor U9717 (N_9717,N_3278,N_2497);
and U9718 (N_9718,N_3823,N_3331);
and U9719 (N_9719,N_2297,N_4304);
nor U9720 (N_9720,N_4834,N_4764);
or U9721 (N_9721,N_2897,N_1647);
or U9722 (N_9722,N_2411,N_1398);
or U9723 (N_9723,N_2317,N_4226);
or U9724 (N_9724,N_2571,N_3811);
or U9725 (N_9725,N_1912,N_2956);
xnor U9726 (N_9726,N_2971,N_3535);
nor U9727 (N_9727,N_945,N_668);
and U9728 (N_9728,N_992,N_4359);
nand U9729 (N_9729,N_2209,N_4320);
xnor U9730 (N_9730,N_2083,N_954);
and U9731 (N_9731,N_915,N_3030);
and U9732 (N_9732,N_1289,N_4121);
and U9733 (N_9733,N_1147,N_2138);
nor U9734 (N_9734,N_3022,N_4987);
or U9735 (N_9735,N_1548,N_2913);
or U9736 (N_9736,N_2409,N_4519);
or U9737 (N_9737,N_1153,N_1956);
and U9738 (N_9738,N_3920,N_1923);
or U9739 (N_9739,N_586,N_233);
or U9740 (N_9740,N_644,N_935);
xnor U9741 (N_9741,N_2347,N_790);
and U9742 (N_9742,N_4237,N_689);
nand U9743 (N_9743,N_2883,N_3452);
xnor U9744 (N_9744,N_1683,N_4196);
xnor U9745 (N_9745,N_3800,N_264);
nand U9746 (N_9746,N_4717,N_3270);
xnor U9747 (N_9747,N_2139,N_4033);
or U9748 (N_9748,N_2114,N_1893);
and U9749 (N_9749,N_3789,N_4555);
nand U9750 (N_9750,N_4369,N_2704);
xnor U9751 (N_9751,N_1471,N_2524);
or U9752 (N_9752,N_797,N_2408);
and U9753 (N_9753,N_4298,N_31);
nand U9754 (N_9754,N_4890,N_2987);
and U9755 (N_9755,N_3343,N_233);
nand U9756 (N_9756,N_485,N_4794);
nor U9757 (N_9757,N_2900,N_4591);
nand U9758 (N_9758,N_540,N_1033);
nand U9759 (N_9759,N_606,N_3050);
and U9760 (N_9760,N_3994,N_1824);
nor U9761 (N_9761,N_832,N_1024);
nand U9762 (N_9762,N_456,N_1104);
xor U9763 (N_9763,N_3782,N_2215);
xnor U9764 (N_9764,N_2347,N_4227);
xor U9765 (N_9765,N_3942,N_3532);
xor U9766 (N_9766,N_2412,N_31);
xor U9767 (N_9767,N_1230,N_4112);
xnor U9768 (N_9768,N_2988,N_2057);
xnor U9769 (N_9769,N_2693,N_3890);
xor U9770 (N_9770,N_3461,N_344);
xnor U9771 (N_9771,N_1916,N_2796);
xnor U9772 (N_9772,N_4423,N_4980);
xor U9773 (N_9773,N_2740,N_3677);
and U9774 (N_9774,N_866,N_4194);
nor U9775 (N_9775,N_238,N_2815);
nand U9776 (N_9776,N_1302,N_1254);
or U9777 (N_9777,N_4180,N_3594);
xor U9778 (N_9778,N_2678,N_1900);
nand U9779 (N_9779,N_1206,N_3910);
and U9780 (N_9780,N_3124,N_3718);
nand U9781 (N_9781,N_4562,N_1798);
and U9782 (N_9782,N_3612,N_834);
nor U9783 (N_9783,N_3814,N_4371);
or U9784 (N_9784,N_3073,N_3995);
and U9785 (N_9785,N_282,N_922);
nor U9786 (N_9786,N_1365,N_4483);
nor U9787 (N_9787,N_1289,N_1534);
and U9788 (N_9788,N_4543,N_1762);
xor U9789 (N_9789,N_2673,N_659);
or U9790 (N_9790,N_2371,N_3171);
nor U9791 (N_9791,N_2681,N_2230);
or U9792 (N_9792,N_3862,N_659);
nor U9793 (N_9793,N_1241,N_622);
nand U9794 (N_9794,N_2661,N_4192);
xor U9795 (N_9795,N_1942,N_4060);
or U9796 (N_9796,N_3895,N_2823);
and U9797 (N_9797,N_252,N_2500);
or U9798 (N_9798,N_2253,N_3415);
xnor U9799 (N_9799,N_537,N_883);
and U9800 (N_9800,N_1026,N_3451);
nor U9801 (N_9801,N_3772,N_1805);
or U9802 (N_9802,N_250,N_437);
or U9803 (N_9803,N_1090,N_1598);
nor U9804 (N_9804,N_3415,N_3735);
or U9805 (N_9805,N_3921,N_923);
or U9806 (N_9806,N_1573,N_3416);
nand U9807 (N_9807,N_4645,N_3089);
and U9808 (N_9808,N_3566,N_959);
xor U9809 (N_9809,N_70,N_4847);
xnor U9810 (N_9810,N_1256,N_3497);
nor U9811 (N_9811,N_4494,N_441);
and U9812 (N_9812,N_4832,N_117);
and U9813 (N_9813,N_2992,N_1644);
xor U9814 (N_9814,N_3681,N_2932);
and U9815 (N_9815,N_958,N_1692);
nor U9816 (N_9816,N_1027,N_3915);
xor U9817 (N_9817,N_1155,N_1159);
nor U9818 (N_9818,N_2294,N_3328);
and U9819 (N_9819,N_3046,N_4583);
and U9820 (N_9820,N_3547,N_1987);
nor U9821 (N_9821,N_4990,N_2014);
or U9822 (N_9822,N_2751,N_12);
xor U9823 (N_9823,N_1152,N_889);
or U9824 (N_9824,N_4942,N_933);
nand U9825 (N_9825,N_991,N_1720);
and U9826 (N_9826,N_1717,N_51);
nand U9827 (N_9827,N_106,N_1496);
xnor U9828 (N_9828,N_3304,N_3034);
nor U9829 (N_9829,N_3501,N_4594);
nand U9830 (N_9830,N_4387,N_3237);
or U9831 (N_9831,N_200,N_2467);
nand U9832 (N_9832,N_1592,N_192);
nand U9833 (N_9833,N_1891,N_261);
nand U9834 (N_9834,N_2146,N_1683);
or U9835 (N_9835,N_3205,N_4229);
nand U9836 (N_9836,N_586,N_670);
nand U9837 (N_9837,N_3141,N_4164);
and U9838 (N_9838,N_348,N_812);
and U9839 (N_9839,N_2270,N_4132);
xnor U9840 (N_9840,N_1448,N_4516);
nand U9841 (N_9841,N_3381,N_1712);
or U9842 (N_9842,N_4704,N_940);
nor U9843 (N_9843,N_4398,N_3122);
xnor U9844 (N_9844,N_1384,N_876);
and U9845 (N_9845,N_2684,N_1508);
xor U9846 (N_9846,N_2753,N_2328);
nand U9847 (N_9847,N_1470,N_1938);
nand U9848 (N_9848,N_2347,N_1986);
xor U9849 (N_9849,N_2413,N_1514);
nor U9850 (N_9850,N_1789,N_4458);
nor U9851 (N_9851,N_4969,N_2904);
and U9852 (N_9852,N_1726,N_4489);
nand U9853 (N_9853,N_4333,N_4054);
xnor U9854 (N_9854,N_229,N_83);
and U9855 (N_9855,N_4291,N_952);
xor U9856 (N_9856,N_2725,N_4205);
nand U9857 (N_9857,N_3003,N_3317);
xnor U9858 (N_9858,N_324,N_4552);
nor U9859 (N_9859,N_3128,N_2067);
nor U9860 (N_9860,N_3746,N_809);
nor U9861 (N_9861,N_1199,N_4045);
xnor U9862 (N_9862,N_3892,N_4400);
nor U9863 (N_9863,N_4309,N_3745);
nand U9864 (N_9864,N_943,N_522);
and U9865 (N_9865,N_1969,N_4719);
nand U9866 (N_9866,N_2721,N_2033);
or U9867 (N_9867,N_4100,N_1075);
xnor U9868 (N_9868,N_3586,N_643);
nor U9869 (N_9869,N_405,N_1796);
xnor U9870 (N_9870,N_4835,N_2710);
nor U9871 (N_9871,N_1294,N_1078);
and U9872 (N_9872,N_609,N_4223);
or U9873 (N_9873,N_3979,N_1033);
nor U9874 (N_9874,N_3211,N_4521);
xnor U9875 (N_9875,N_1064,N_1145);
xnor U9876 (N_9876,N_584,N_334);
or U9877 (N_9877,N_4071,N_3563);
nor U9878 (N_9878,N_2600,N_3267);
or U9879 (N_9879,N_4726,N_3675);
xnor U9880 (N_9880,N_4270,N_1792);
xor U9881 (N_9881,N_3392,N_2461);
nor U9882 (N_9882,N_1127,N_2119);
nand U9883 (N_9883,N_180,N_4669);
nand U9884 (N_9884,N_4339,N_2836);
and U9885 (N_9885,N_3892,N_4678);
nand U9886 (N_9886,N_4024,N_1239);
and U9887 (N_9887,N_3407,N_4111);
nor U9888 (N_9888,N_2822,N_3667);
nor U9889 (N_9889,N_1108,N_173);
nand U9890 (N_9890,N_467,N_2922);
and U9891 (N_9891,N_4862,N_373);
or U9892 (N_9892,N_1543,N_4971);
nor U9893 (N_9893,N_3661,N_3383);
xor U9894 (N_9894,N_4499,N_3374);
or U9895 (N_9895,N_851,N_3813);
nor U9896 (N_9896,N_922,N_1539);
nand U9897 (N_9897,N_2631,N_3981);
nand U9898 (N_9898,N_400,N_1053);
and U9899 (N_9899,N_3164,N_4903);
nor U9900 (N_9900,N_994,N_2167);
nor U9901 (N_9901,N_1042,N_1848);
nor U9902 (N_9902,N_897,N_2365);
nor U9903 (N_9903,N_4508,N_312);
or U9904 (N_9904,N_1994,N_4777);
nor U9905 (N_9905,N_2539,N_2992);
and U9906 (N_9906,N_584,N_3894);
xor U9907 (N_9907,N_3827,N_3245);
or U9908 (N_9908,N_3507,N_4526);
nand U9909 (N_9909,N_2821,N_3157);
nand U9910 (N_9910,N_3176,N_1976);
xnor U9911 (N_9911,N_4890,N_949);
xor U9912 (N_9912,N_1023,N_1304);
nor U9913 (N_9913,N_206,N_4386);
xor U9914 (N_9914,N_136,N_454);
or U9915 (N_9915,N_3040,N_1596);
xnor U9916 (N_9916,N_3500,N_2231);
nor U9917 (N_9917,N_2447,N_1976);
nand U9918 (N_9918,N_183,N_3844);
xor U9919 (N_9919,N_4922,N_2557);
xnor U9920 (N_9920,N_654,N_4263);
nor U9921 (N_9921,N_3390,N_3190);
xor U9922 (N_9922,N_4652,N_3841);
and U9923 (N_9923,N_828,N_637);
and U9924 (N_9924,N_4592,N_1665);
xnor U9925 (N_9925,N_29,N_1424);
and U9926 (N_9926,N_4053,N_4804);
nand U9927 (N_9927,N_2662,N_3611);
or U9928 (N_9928,N_1390,N_1090);
nand U9929 (N_9929,N_3331,N_2560);
and U9930 (N_9930,N_4850,N_3855);
nor U9931 (N_9931,N_4604,N_675);
or U9932 (N_9932,N_42,N_4163);
xnor U9933 (N_9933,N_4600,N_4744);
xnor U9934 (N_9934,N_4991,N_944);
or U9935 (N_9935,N_3848,N_156);
or U9936 (N_9936,N_88,N_4603);
nand U9937 (N_9937,N_419,N_929);
xor U9938 (N_9938,N_3306,N_351);
or U9939 (N_9939,N_4782,N_525);
xnor U9940 (N_9940,N_867,N_2188);
nor U9941 (N_9941,N_355,N_1345);
xor U9942 (N_9942,N_2967,N_4495);
nand U9943 (N_9943,N_263,N_2937);
nand U9944 (N_9944,N_864,N_4087);
nor U9945 (N_9945,N_4395,N_401);
and U9946 (N_9946,N_1775,N_3199);
nor U9947 (N_9947,N_2201,N_1060);
or U9948 (N_9948,N_1510,N_4135);
or U9949 (N_9949,N_1325,N_3861);
and U9950 (N_9950,N_2301,N_3033);
nand U9951 (N_9951,N_3430,N_1735);
or U9952 (N_9952,N_2587,N_1949);
nor U9953 (N_9953,N_4016,N_966);
xnor U9954 (N_9954,N_2700,N_866);
and U9955 (N_9955,N_1848,N_1569);
xor U9956 (N_9956,N_3448,N_2452);
nor U9957 (N_9957,N_3433,N_1842);
and U9958 (N_9958,N_2816,N_729);
nand U9959 (N_9959,N_252,N_1588);
and U9960 (N_9960,N_1048,N_1540);
nor U9961 (N_9961,N_4303,N_716);
xnor U9962 (N_9962,N_3376,N_1134);
nand U9963 (N_9963,N_0,N_1451);
nand U9964 (N_9964,N_2905,N_1349);
and U9965 (N_9965,N_4113,N_2755);
xor U9966 (N_9966,N_3210,N_1553);
xnor U9967 (N_9967,N_4026,N_2878);
or U9968 (N_9968,N_3116,N_3032);
xnor U9969 (N_9969,N_292,N_6);
xnor U9970 (N_9970,N_463,N_3771);
nand U9971 (N_9971,N_4997,N_362);
nand U9972 (N_9972,N_2165,N_3179);
nand U9973 (N_9973,N_1174,N_1325);
xor U9974 (N_9974,N_2999,N_209);
nand U9975 (N_9975,N_1268,N_2798);
xnor U9976 (N_9976,N_1214,N_1563);
nor U9977 (N_9977,N_4639,N_2558);
or U9978 (N_9978,N_4275,N_1303);
or U9979 (N_9979,N_23,N_3967);
or U9980 (N_9980,N_2627,N_2497);
or U9981 (N_9981,N_4205,N_3111);
and U9982 (N_9982,N_2536,N_3748);
xnor U9983 (N_9983,N_3155,N_208);
and U9984 (N_9984,N_1885,N_1107);
nor U9985 (N_9985,N_4717,N_3786);
nor U9986 (N_9986,N_2513,N_2772);
and U9987 (N_9987,N_240,N_3140);
nor U9988 (N_9988,N_780,N_1715);
nor U9989 (N_9989,N_1235,N_2974);
nand U9990 (N_9990,N_887,N_2415);
or U9991 (N_9991,N_808,N_430);
xnor U9992 (N_9992,N_1129,N_1811);
nand U9993 (N_9993,N_2681,N_1288);
nor U9994 (N_9994,N_2392,N_42);
nand U9995 (N_9995,N_689,N_2127);
nand U9996 (N_9996,N_1008,N_1398);
xnor U9997 (N_9997,N_2365,N_3206);
xor U9998 (N_9998,N_4781,N_32);
xnor U9999 (N_9999,N_2444,N_3012);
nor U10000 (N_10000,N_8180,N_7352);
and U10001 (N_10001,N_6734,N_6906);
nand U10002 (N_10002,N_8189,N_5512);
or U10003 (N_10003,N_7984,N_8190);
nor U10004 (N_10004,N_5131,N_8476);
nor U10005 (N_10005,N_8318,N_5685);
nor U10006 (N_10006,N_5069,N_9128);
and U10007 (N_10007,N_6759,N_9503);
nor U10008 (N_10008,N_9622,N_7986);
nor U10009 (N_10009,N_6132,N_6460);
or U10010 (N_10010,N_9418,N_9449);
nand U10011 (N_10011,N_7764,N_9716);
or U10012 (N_10012,N_9342,N_5876);
nor U10013 (N_10013,N_7643,N_8134);
or U10014 (N_10014,N_8350,N_5273);
nand U10015 (N_10015,N_9647,N_5323);
xnor U10016 (N_10016,N_8677,N_9484);
nor U10017 (N_10017,N_9678,N_9407);
nor U10018 (N_10018,N_8505,N_9152);
xnor U10019 (N_10019,N_5154,N_9677);
nand U10020 (N_10020,N_7867,N_9661);
nand U10021 (N_10021,N_8570,N_9328);
xnor U10022 (N_10022,N_5983,N_6474);
and U10023 (N_10023,N_9169,N_6608);
or U10024 (N_10024,N_7271,N_6213);
or U10025 (N_10025,N_6981,N_7022);
xnor U10026 (N_10026,N_7250,N_7014);
xor U10027 (N_10027,N_9843,N_7564);
or U10028 (N_10028,N_7964,N_5484);
nor U10029 (N_10029,N_6414,N_9664);
and U10030 (N_10030,N_8874,N_5989);
or U10031 (N_10031,N_5994,N_8962);
nand U10032 (N_10032,N_6176,N_9682);
nor U10033 (N_10033,N_8515,N_5107);
xor U10034 (N_10034,N_5104,N_6985);
xor U10035 (N_10035,N_7615,N_5871);
nand U10036 (N_10036,N_6380,N_5972);
or U10037 (N_10037,N_8866,N_8520);
and U10038 (N_10038,N_6263,N_8833);
nor U10039 (N_10039,N_6136,N_7664);
nor U10040 (N_10040,N_5927,N_9931);
xnor U10041 (N_10041,N_9060,N_6877);
nor U10042 (N_10042,N_6999,N_5436);
xnor U10043 (N_10043,N_8243,N_6321);
xnor U10044 (N_10044,N_5499,N_7686);
nand U10045 (N_10045,N_8121,N_9408);
or U10046 (N_10046,N_5633,N_7012);
nand U10047 (N_10047,N_8537,N_6060);
xor U10048 (N_10048,N_6559,N_7552);
nand U10049 (N_10049,N_8383,N_9992);
nand U10050 (N_10050,N_8933,N_5072);
xnor U10051 (N_10051,N_5977,N_9132);
nor U10052 (N_10052,N_6731,N_5655);
or U10053 (N_10053,N_9954,N_9989);
and U10054 (N_10054,N_6477,N_7602);
nor U10055 (N_10055,N_5664,N_9116);
nand U10056 (N_10056,N_6776,N_6248);
xnor U10057 (N_10057,N_6643,N_5317);
nand U10058 (N_10058,N_8750,N_6536);
nand U10059 (N_10059,N_7624,N_9141);
nand U10060 (N_10060,N_5081,N_8079);
xnor U10061 (N_10061,N_7059,N_7784);
or U10062 (N_10062,N_8917,N_6338);
and U10063 (N_10063,N_5314,N_9753);
xor U10064 (N_10064,N_9092,N_8627);
or U10065 (N_10065,N_5683,N_9430);
nand U10066 (N_10066,N_6087,N_9086);
and U10067 (N_10067,N_8393,N_6467);
xor U10068 (N_10068,N_9898,N_6539);
xnor U10069 (N_10069,N_9690,N_7662);
xor U10070 (N_10070,N_8174,N_6206);
and U10071 (N_10071,N_9631,N_9340);
or U10072 (N_10072,N_8151,N_8403);
and U10073 (N_10073,N_9040,N_7896);
nand U10074 (N_10074,N_8513,N_8111);
nand U10075 (N_10075,N_9069,N_6458);
nor U10076 (N_10076,N_9229,N_7665);
and U10077 (N_10077,N_8905,N_7902);
xnor U10078 (N_10078,N_7153,N_8078);
and U10079 (N_10079,N_9654,N_6346);
and U10080 (N_10080,N_5504,N_6145);
or U10081 (N_10081,N_6885,N_9260);
nor U10082 (N_10082,N_7337,N_9296);
and U10083 (N_10083,N_5669,N_7613);
nand U10084 (N_10084,N_8036,N_6751);
nand U10085 (N_10085,N_9115,N_5000);
and U10086 (N_10086,N_8082,N_5597);
and U10087 (N_10087,N_7502,N_6806);
xor U10088 (N_10088,N_5648,N_7150);
xor U10089 (N_10089,N_9881,N_8379);
nand U10090 (N_10090,N_8314,N_5596);
xor U10091 (N_10091,N_8132,N_5143);
nand U10092 (N_10092,N_8218,N_8658);
nand U10093 (N_10093,N_8535,N_9525);
or U10094 (N_10094,N_5352,N_5878);
and U10095 (N_10095,N_6977,N_5904);
xor U10096 (N_10096,N_8880,N_7302);
or U10097 (N_10097,N_6599,N_5568);
or U10098 (N_10098,N_8839,N_6694);
nand U10099 (N_10099,N_9043,N_6192);
xor U10100 (N_10100,N_9571,N_8568);
and U10101 (N_10101,N_7267,N_6675);
nor U10102 (N_10102,N_9318,N_6764);
nand U10103 (N_10103,N_9316,N_6855);
nor U10104 (N_10104,N_9861,N_7540);
nand U10105 (N_10105,N_8785,N_9012);
and U10106 (N_10106,N_5425,N_5213);
xor U10107 (N_10107,N_9903,N_9701);
and U10108 (N_10108,N_5838,N_7349);
or U10109 (N_10109,N_7081,N_7288);
xor U10110 (N_10110,N_5928,N_7158);
xor U10111 (N_10111,N_9470,N_6942);
nand U10112 (N_10112,N_8023,N_5916);
or U10113 (N_10113,N_7141,N_9211);
nor U10114 (N_10114,N_6691,N_7897);
nand U10115 (N_10115,N_7846,N_7528);
nand U10116 (N_10116,N_8529,N_6735);
nand U10117 (N_10117,N_8009,N_5298);
nor U10118 (N_10118,N_8137,N_7706);
xnor U10119 (N_10119,N_7497,N_6421);
xor U10120 (N_10120,N_9191,N_6221);
or U10121 (N_10121,N_5668,N_9436);
nor U10122 (N_10122,N_9594,N_5841);
or U10123 (N_10123,N_9514,N_5413);
nor U10124 (N_10124,N_8273,N_7005);
nor U10125 (N_10125,N_9944,N_7134);
nor U10126 (N_10126,N_7914,N_9447);
xnor U10127 (N_10127,N_8265,N_7123);
nand U10128 (N_10128,N_9359,N_7305);
or U10129 (N_10129,N_6296,N_7345);
xnor U10130 (N_10130,N_6898,N_9331);
xnor U10131 (N_10131,N_6696,N_9061);
and U10132 (N_10132,N_8981,N_9597);
nand U10133 (N_10133,N_8329,N_7304);
xnor U10134 (N_10134,N_9190,N_5612);
xnor U10135 (N_10135,N_7887,N_9627);
nor U10136 (N_10136,N_7608,N_6491);
nor U10137 (N_10137,N_6328,N_8032);
xor U10138 (N_10138,N_6640,N_7210);
nand U10139 (N_10139,N_5510,N_6258);
xnor U10140 (N_10140,N_6493,N_9769);
xor U10141 (N_10141,N_5300,N_8313);
and U10142 (N_10142,N_9409,N_9350);
and U10143 (N_10143,N_5952,N_9455);
xor U10144 (N_10144,N_7233,N_6378);
xor U10145 (N_10145,N_8472,N_9816);
nand U10146 (N_10146,N_6685,N_9587);
nand U10147 (N_10147,N_6451,N_6360);
or U10148 (N_10148,N_8156,N_6143);
xor U10149 (N_10149,N_9648,N_9367);
nor U10150 (N_10150,N_8085,N_7529);
nor U10151 (N_10151,N_6104,N_9228);
nand U10152 (N_10152,N_8704,N_7882);
nand U10153 (N_10153,N_8382,N_5162);
or U10154 (N_10154,N_6308,N_7946);
and U10155 (N_10155,N_5637,N_8673);
and U10156 (N_10156,N_7430,N_6719);
nand U10157 (N_10157,N_8340,N_6048);
and U10158 (N_10158,N_6201,N_5703);
and U10159 (N_10159,N_7493,N_8000);
xor U10160 (N_10160,N_6598,N_7165);
or U10161 (N_10161,N_5355,N_9310);
nor U10162 (N_10162,N_7561,N_6622);
or U10163 (N_10163,N_8187,N_8882);
nand U10164 (N_10164,N_9875,N_5270);
xnor U10165 (N_10165,N_5886,N_6121);
and U10166 (N_10166,N_5090,N_8812);
and U10167 (N_10167,N_9405,N_8021);
and U10168 (N_10168,N_6850,N_8972);
nand U10169 (N_10169,N_7184,N_9822);
xor U10170 (N_10170,N_5820,N_7104);
xnor U10171 (N_10171,N_5256,N_5457);
nand U10172 (N_10172,N_6266,N_5527);
nand U10173 (N_10173,N_8489,N_5823);
nand U10174 (N_10174,N_5106,N_7264);
and U10175 (N_10175,N_8290,N_8827);
nand U10176 (N_10176,N_8296,N_8395);
and U10177 (N_10177,N_8824,N_7135);
and U10178 (N_10178,N_9926,N_5053);
or U10179 (N_10179,N_8649,N_6285);
nand U10180 (N_10180,N_8286,N_5327);
or U10181 (N_10181,N_8978,N_5850);
xor U10182 (N_10182,N_7688,N_8266);
nand U10183 (N_10183,N_6398,N_6080);
and U10184 (N_10184,N_6573,N_6688);
nand U10185 (N_10185,N_5555,N_8510);
xnor U10186 (N_10186,N_8295,N_8714);
nand U10187 (N_10187,N_6367,N_9669);
nand U10188 (N_10188,N_5138,N_9492);
nor U10189 (N_10189,N_7173,N_7700);
and U10190 (N_10190,N_6142,N_9083);
nand U10191 (N_10191,N_6769,N_9885);
nor U10192 (N_10192,N_6124,N_8644);
and U10193 (N_10193,N_8963,N_7963);
nor U10194 (N_10194,N_9464,N_5292);
nor U10195 (N_10195,N_8847,N_7750);
xor U10196 (N_10196,N_5447,N_8059);
nor U10197 (N_10197,N_6365,N_8223);
nor U10198 (N_10198,N_9502,N_8903);
or U10199 (N_10199,N_7282,N_6409);
or U10200 (N_10200,N_5339,N_6086);
xnor U10201 (N_10201,N_7145,N_9939);
and U10202 (N_10202,N_5877,N_6819);
nor U10203 (N_10203,N_5260,N_6077);
nor U10204 (N_10204,N_6307,N_5462);
and U10205 (N_10205,N_7651,N_8779);
or U10206 (N_10206,N_6770,N_8851);
nor U10207 (N_10207,N_9650,N_7911);
or U10208 (N_10208,N_5465,N_9065);
or U10209 (N_10209,N_5266,N_6144);
nand U10210 (N_10210,N_8835,N_5584);
nand U10211 (N_10211,N_8718,N_7415);
and U10212 (N_10212,N_6200,N_5762);
or U10213 (N_10213,N_5624,N_7402);
nor U10214 (N_10214,N_6320,N_5939);
or U10215 (N_10215,N_9642,N_7572);
and U10216 (N_10216,N_7129,N_6229);
and U10217 (N_10217,N_6560,N_8752);
nor U10218 (N_10218,N_5189,N_6700);
xor U10219 (N_10219,N_8283,N_9501);
and U10220 (N_10220,N_6472,N_7072);
and U10221 (N_10221,N_7649,N_5769);
and U10222 (N_10222,N_9013,N_9022);
nor U10223 (N_10223,N_8241,N_8890);
and U10224 (N_10224,N_7108,N_9512);
and U10225 (N_10225,N_5384,N_9135);
or U10226 (N_10226,N_8317,N_6520);
nor U10227 (N_10227,N_9553,N_5564);
nand U10228 (N_10228,N_5840,N_8519);
xor U10229 (N_10229,N_7919,N_6010);
xor U10230 (N_10230,N_5716,N_5414);
or U10231 (N_10231,N_6801,N_9073);
nor U10232 (N_10232,N_6076,N_7110);
xnor U10233 (N_10233,N_8511,N_9706);
xnor U10234 (N_10234,N_9815,N_5360);
or U10235 (N_10235,N_6337,N_8264);
or U10236 (N_10236,N_7730,N_7417);
xor U10237 (N_10237,N_7853,N_9760);
and U10238 (N_10238,N_7363,N_6646);
nor U10239 (N_10239,N_5477,N_7289);
xnor U10240 (N_10240,N_6055,N_9727);
nand U10241 (N_10241,N_6616,N_5696);
and U10242 (N_10242,N_7843,N_6529);
nor U10243 (N_10243,N_7298,N_6358);
or U10244 (N_10244,N_7819,N_9304);
and U10245 (N_10245,N_8877,N_7756);
xnor U10246 (N_10246,N_9749,N_6746);
nor U10247 (N_10247,N_5613,N_6094);
nand U10248 (N_10248,N_6811,N_6817);
or U10249 (N_10249,N_6034,N_7100);
or U10250 (N_10250,N_7944,N_6941);
xnor U10251 (N_10251,N_9017,N_9240);
and U10252 (N_10252,N_8524,N_9595);
and U10253 (N_10253,N_9142,N_9231);
nor U10254 (N_10254,N_9101,N_9981);
xnor U10255 (N_10255,N_5418,N_9972);
nor U10256 (N_10256,N_7637,N_9071);
nor U10257 (N_10257,N_5007,N_5581);
nand U10258 (N_10258,N_6901,N_5306);
nand U10259 (N_10259,N_9871,N_7916);
xnor U10260 (N_10260,N_7926,N_5813);
nand U10261 (N_10261,N_8342,N_8729);
or U10262 (N_10262,N_5250,N_7742);
nor U10263 (N_10263,N_9032,N_6035);
nand U10264 (N_10264,N_9715,N_7127);
and U10265 (N_10265,N_5950,N_6293);
nand U10266 (N_10266,N_5423,N_9349);
and U10267 (N_10267,N_8456,N_6923);
xor U10268 (N_10268,N_9937,N_7391);
or U10269 (N_10269,N_8122,N_7114);
nand U10270 (N_10270,N_5417,N_8479);
or U10271 (N_10271,N_7575,N_9860);
xor U10272 (N_10272,N_7287,N_5221);
and U10273 (N_10273,N_6677,N_8607);
nor U10274 (N_10274,N_7120,N_9030);
nor U10275 (N_10275,N_7755,N_6208);
or U10276 (N_10276,N_5640,N_9672);
and U10277 (N_10277,N_6462,N_6628);
xnor U10278 (N_10278,N_8950,N_5780);
xor U10279 (N_10279,N_5526,N_9075);
nand U10280 (N_10280,N_5604,N_5434);
xor U10281 (N_10281,N_6858,N_6828);
or U10282 (N_10282,N_9508,N_5538);
xor U10283 (N_10283,N_8719,N_7315);
nand U10284 (N_10284,N_7996,N_5013);
xnor U10285 (N_10285,N_9942,N_5966);
or U10286 (N_10286,N_6260,N_6317);
nand U10287 (N_10287,N_9108,N_6908);
nor U10288 (N_10288,N_5313,N_5194);
xnor U10289 (N_10289,N_6912,N_6930);
nand U10290 (N_10290,N_9536,N_7708);
xor U10291 (N_10291,N_7702,N_8623);
nand U10292 (N_10292,N_9524,N_6499);
or U10293 (N_10293,N_9351,N_5023);
and U10294 (N_10294,N_9936,N_9561);
xor U10295 (N_10295,N_9019,N_9845);
or U10296 (N_10296,N_5231,N_5486);
nor U10297 (N_10297,N_9663,N_9037);
nor U10298 (N_10298,N_6023,N_6921);
and U10299 (N_10299,N_8365,N_7719);
or U10300 (N_10300,N_7166,N_6259);
and U10301 (N_10301,N_9439,N_7043);
nand U10302 (N_10302,N_8095,N_9431);
nor U10303 (N_10303,N_7676,N_7201);
and U10304 (N_10304,N_6235,N_6487);
xor U10305 (N_10305,N_9914,N_9879);
or U10306 (N_10306,N_7490,N_6821);
xor U10307 (N_10307,N_8744,N_9560);
and U10308 (N_10308,N_5095,N_6108);
and U10309 (N_10309,N_7235,N_9840);
nand U10310 (N_10310,N_7714,N_7310);
nand U10311 (N_10311,N_5995,N_5898);
nand U10312 (N_10312,N_5100,N_5678);
nor U10313 (N_10313,N_8894,N_6214);
nor U10314 (N_10314,N_5215,N_8388);
nand U10315 (N_10315,N_5501,N_7036);
and U10316 (N_10316,N_7217,N_7607);
xnor U10317 (N_10317,N_5918,N_5617);
and U10318 (N_10318,N_7521,N_8098);
and U10319 (N_10319,N_9835,N_6165);
nor U10320 (N_10320,N_7979,N_9705);
nand U10321 (N_10321,N_9156,N_5547);
and U10322 (N_10322,N_6045,N_8540);
or U10323 (N_10323,N_9993,N_8923);
or U10324 (N_10324,N_5570,N_6186);
and U10325 (N_10325,N_8343,N_5257);
xnor U10326 (N_10326,N_8927,N_9427);
or U10327 (N_10327,N_7594,N_5986);
nand U10328 (N_10328,N_8346,N_8352);
nand U10329 (N_10329,N_8404,N_8061);
or U10330 (N_10330,N_6809,N_9710);
nand U10331 (N_10331,N_6062,N_6410);
nor U10332 (N_10332,N_8154,N_8319);
or U10333 (N_10333,N_5505,N_8054);
nand U10334 (N_10334,N_5185,N_5748);
and U10335 (N_10335,N_7972,N_7035);
xnor U10336 (N_10336,N_6827,N_5035);
and U10337 (N_10337,N_9401,N_7457);
nand U10338 (N_10338,N_6532,N_5350);
or U10339 (N_10339,N_7186,N_8637);
xnor U10340 (N_10340,N_8942,N_5003);
xor U10341 (N_10341,N_6519,N_8982);
and U10342 (N_10342,N_6888,N_6780);
nor U10343 (N_10343,N_7617,N_7291);
nor U10344 (N_10344,N_8803,N_6925);
xnor U10345 (N_10345,N_5046,N_5021);
nor U10346 (N_10346,N_5925,N_6239);
and U10347 (N_10347,N_9222,N_5326);
nor U10348 (N_10348,N_7913,N_9528);
nor U10349 (N_10349,N_8247,N_7478);
xor U10350 (N_10350,N_9245,N_6934);
nor U10351 (N_10351,N_8349,N_6140);
nand U10352 (N_10352,N_9049,N_7346);
xnor U10353 (N_10353,N_8274,N_7499);
nand U10354 (N_10354,N_8011,N_5309);
nand U10355 (N_10355,N_6151,N_6969);
nand U10356 (N_10356,N_5150,N_8091);
xnor U10357 (N_10357,N_7246,N_7894);
nor U10358 (N_10358,N_8705,N_6386);
and U10359 (N_10359,N_6318,N_5643);
nor U10360 (N_10360,N_5663,N_9563);
nand U10361 (N_10361,N_7690,N_5011);
xor U10362 (N_10362,N_8583,N_9603);
or U10363 (N_10363,N_7074,N_5695);
and U10364 (N_10364,N_6543,N_9963);
nand U10365 (N_10365,N_9806,N_9410);
or U10366 (N_10366,N_8141,N_5151);
nor U10367 (N_10367,N_6413,N_6383);
nor U10368 (N_10368,N_6355,N_6994);
or U10369 (N_10369,N_7577,N_6336);
or U10370 (N_10370,N_5737,N_8363);
or U10371 (N_10371,N_6808,N_6298);
nor U10372 (N_10372,N_7486,N_8415);
nand U10373 (N_10373,N_9122,N_9422);
xnor U10374 (N_10374,N_9633,N_7320);
nor U10375 (N_10375,N_5688,N_8376);
and U10376 (N_10376,N_6902,N_5161);
and U10377 (N_10377,N_7510,N_9913);
or U10378 (N_10378,N_8864,N_8051);
or U10379 (N_10379,N_9919,N_5055);
and U10380 (N_10380,N_9708,N_7672);
and U10381 (N_10381,N_7898,N_7859);
or U10382 (N_10382,N_8786,N_6927);
xnor U10383 (N_10383,N_6506,N_8072);
nor U10384 (N_10384,N_8022,N_8581);
nand U10385 (N_10385,N_9140,N_8699);
nor U10386 (N_10386,N_7815,N_8634);
or U10387 (N_10387,N_8183,N_6683);
xor U10388 (N_10388,N_5768,N_9203);
or U10389 (N_10389,N_7831,N_5765);
nor U10390 (N_10390,N_9505,N_7865);
nand U10391 (N_10391,N_6130,N_9298);
nor U10392 (N_10392,N_7020,N_7342);
nand U10393 (N_10393,N_7582,N_6348);
nor U10394 (N_10394,N_5521,N_5856);
nor U10395 (N_10395,N_9036,N_6917);
nor U10396 (N_10396,N_5761,N_8696);
xnor U10397 (N_10397,N_9489,N_5404);
nand U10398 (N_10398,N_8324,N_5701);
or U10399 (N_10399,N_8660,N_7641);
and U10400 (N_10400,N_8086,N_9858);
and U10401 (N_10401,N_5537,N_6204);
or U10402 (N_10402,N_7749,N_9281);
or U10403 (N_10403,N_8780,N_5324);
and U10404 (N_10404,N_7943,N_8553);
nand U10405 (N_10405,N_7132,N_5310);
nand U10406 (N_10406,N_7469,N_7297);
nor U10407 (N_10407,N_5321,N_5195);
xor U10408 (N_10408,N_6389,N_9754);
nand U10409 (N_10409,N_9490,N_5789);
nor U10410 (N_10410,N_8038,N_5278);
xor U10411 (N_10411,N_7669,N_8574);
and U10412 (N_10412,N_8777,N_9957);
xor U10413 (N_10413,N_7160,N_6575);
and U10414 (N_10414,N_5987,N_9081);
and U10415 (N_10415,N_5660,N_9181);
xor U10416 (N_10416,N_8276,N_9784);
or U10417 (N_10417,N_7745,N_7045);
nand U10418 (N_10418,N_6310,N_8820);
nor U10419 (N_10419,N_9983,N_9168);
xnor U10420 (N_10420,N_7844,N_5357);
xnor U10421 (N_10421,N_9555,N_7174);
or U10422 (N_10422,N_5034,N_9988);
or U10423 (N_10423,N_8881,N_6601);
or U10424 (N_10424,N_5563,N_7405);
nand U10425 (N_10425,N_8397,N_5393);
nand U10426 (N_10426,N_5859,N_7195);
nand U10427 (N_10427,N_6088,N_9125);
nand U10428 (N_10428,N_9659,N_9357);
nand U10429 (N_10429,N_6558,N_7625);
nor U10430 (N_10430,N_6793,N_6212);
xnor U10431 (N_10431,N_7170,N_6388);
or U10432 (N_10432,N_8916,N_5870);
xor U10433 (N_10433,N_5790,N_7475);
nor U10434 (N_10434,N_6630,N_8443);
nand U10435 (N_10435,N_6114,N_5828);
nand U10436 (N_10436,N_6468,N_9014);
and U10437 (N_10437,N_5108,N_5620);
nor U10438 (N_10438,N_6092,N_7767);
nand U10439 (N_10439,N_6653,N_9626);
xnor U10440 (N_10440,N_9802,N_8508);
and U10441 (N_10441,N_6861,N_9208);
or U10442 (N_10442,N_9239,N_8925);
nand U10443 (N_10443,N_7748,N_9730);
nand U10444 (N_10444,N_6216,N_5059);
nor U10445 (N_10445,N_5873,N_8630);
xnor U10446 (N_10446,N_6489,N_9620);
and U10447 (N_10447,N_8661,N_6604);
xor U10448 (N_10448,N_9549,N_6971);
or U10449 (N_10449,N_6392,N_9504);
nand U10450 (N_10450,N_6119,N_9757);
and U10451 (N_10451,N_7442,N_7322);
or U10452 (N_10452,N_8944,N_8113);
or U10453 (N_10453,N_8341,N_7272);
and U10454 (N_10454,N_5671,N_8423);
nand U10455 (N_10455,N_5005,N_8772);
and U10456 (N_10456,N_6729,N_9419);
nand U10457 (N_10457,N_8019,N_5379);
nor U10458 (N_10458,N_6319,N_5800);
or U10459 (N_10459,N_8179,N_9960);
nand U10460 (N_10460,N_9438,N_6486);
xnor U10461 (N_10461,N_6129,N_9870);
xnor U10462 (N_10462,N_7149,N_6919);
and U10463 (N_10463,N_9162,N_5440);
nor U10464 (N_10464,N_7794,N_8569);
nor U10465 (N_10465,N_9366,N_7621);
nand U10466 (N_10466,N_9697,N_7107);
nand U10467 (N_10467,N_8959,N_5001);
nand U10468 (N_10468,N_5642,N_6098);
or U10469 (N_10469,N_5665,N_9067);
xnor U10470 (N_10470,N_5753,N_7878);
and U10471 (N_10471,N_9904,N_7358);
xnor U10472 (N_10472,N_8868,N_8299);
xor U10473 (N_10473,N_6050,N_8138);
nand U10474 (N_10474,N_6372,N_9801);
xnor U10475 (N_10475,N_7078,N_6122);
xnor U10476 (N_10476,N_7600,N_6101);
xor U10477 (N_10477,N_5211,N_9709);
and U10478 (N_10478,N_9666,N_8548);
nand U10479 (N_10479,N_7397,N_8966);
and U10480 (N_10480,N_8775,N_9475);
or U10481 (N_10481,N_7509,N_7087);
nand U10482 (N_10482,N_9787,N_6126);
or U10483 (N_10483,N_9901,N_7658);
or U10484 (N_10484,N_9987,N_6281);
or U10485 (N_10485,N_7194,N_9507);
nor U10486 (N_10486,N_6227,N_6693);
nor U10487 (N_10487,N_7786,N_6538);
nor U10488 (N_10488,N_8155,N_9966);
and U10489 (N_10489,N_5065,N_6311);
nand U10490 (N_10490,N_6480,N_6147);
nor U10491 (N_10491,N_7666,N_5432);
and U10492 (N_10492,N_9862,N_5057);
xor U10493 (N_10493,N_7172,N_9052);
xor U10494 (N_10494,N_6528,N_5579);
and U10495 (N_10495,N_5082,N_8328);
nand U10496 (N_10496,N_8196,N_9254);
xnor U10497 (N_10497,N_6394,N_8119);
nand U10498 (N_10498,N_5851,N_5202);
nor U10499 (N_10499,N_5825,N_5497);
nor U10500 (N_10500,N_7816,N_6368);
nand U10501 (N_10501,N_5784,N_9250);
or U10502 (N_10502,N_8207,N_7538);
and U10503 (N_10503,N_6178,N_7950);
nor U10504 (N_10504,N_5105,N_6313);
nand U10505 (N_10505,N_7880,N_5304);
or U10506 (N_10506,N_9358,N_6804);
and U10507 (N_10507,N_5865,N_8258);
or U10508 (N_10508,N_6860,N_6111);
and U10509 (N_10509,N_8904,N_7514);
or U10510 (N_10510,N_7650,N_6041);
nor U10511 (N_10511,N_8055,N_6016);
or U10512 (N_10512,N_6156,N_6024);
or U10513 (N_10513,N_7290,N_7976);
and U10514 (N_10514,N_9258,N_5732);
and U10515 (N_10515,N_7640,N_9050);
nor U10516 (N_10516,N_9442,N_5184);
nand U10517 (N_10517,N_6219,N_9147);
and U10518 (N_10518,N_9977,N_6405);
nand U10519 (N_10519,N_5187,N_5644);
nor U10520 (N_10520,N_7675,N_9117);
and U10521 (N_10521,N_5307,N_8674);
and U10522 (N_10522,N_7136,N_9632);
or U10523 (N_10523,N_9130,N_7551);
or U10524 (N_10524,N_9575,N_9703);
or U10525 (N_10525,N_8279,N_8831);
nand U10526 (N_10526,N_8702,N_5480);
nand U10527 (N_10527,N_7095,N_6865);
nor U10528 (N_10528,N_7622,N_9499);
and U10529 (N_10529,N_6028,N_7579);
and U10530 (N_10530,N_7741,N_9856);
or U10531 (N_10531,N_7323,N_9485);
and U10532 (N_10532,N_7142,N_8049);
xnor U10533 (N_10533,N_9291,N_9940);
nand U10534 (N_10534,N_6639,N_8285);
xnor U10535 (N_10535,N_8776,N_7209);
nor U10536 (N_10536,N_8206,N_9657);
and U10537 (N_10537,N_5822,N_6515);
nand U10538 (N_10538,N_5603,N_8353);
or U10539 (N_10539,N_8766,N_5729);
xnor U10540 (N_10540,N_8117,N_8210);
nor U10541 (N_10541,N_5677,N_8018);
or U10542 (N_10542,N_6956,N_7791);
xnor U10543 (N_10543,N_5836,N_6185);
and U10544 (N_10544,N_7673,N_9289);
nor U10545 (N_10545,N_6871,N_9533);
xor U10546 (N_10546,N_9255,N_8691);
nand U10547 (N_10547,N_6605,N_9339);
or U10548 (N_10548,N_8860,N_9297);
xor U10549 (N_10549,N_5196,N_6576);
nor U10550 (N_10550,N_7626,N_8861);
and U10551 (N_10551,N_9341,N_9432);
and U10552 (N_10552,N_7954,N_8976);
or U10553 (N_10553,N_9932,N_5083);
or U10554 (N_10554,N_8236,N_9839);
nor U10555 (N_10555,N_6255,N_7071);
nor U10556 (N_10556,N_9453,N_5618);
nor U10557 (N_10557,N_6051,N_9417);
and U10558 (N_10558,N_5710,N_7721);
nor U10559 (N_10559,N_6012,N_8840);
nor U10560 (N_10560,N_5387,N_7011);
or U10561 (N_10561,N_6826,N_7434);
nand U10562 (N_10562,N_5673,N_8302);
and U10563 (N_10563,N_5955,N_5899);
and U10564 (N_10564,N_9589,N_9866);
nor U10565 (N_10565,N_8763,N_6960);
and U10566 (N_10566,N_7704,N_6783);
nor U10567 (N_10567,N_5445,N_7086);
xnor U10568 (N_10568,N_6779,N_9775);
nor U10569 (N_10569,N_7835,N_7197);
nor U10570 (N_10570,N_5879,N_5903);
xnor U10571 (N_10571,N_8665,N_5777);
nor U10572 (N_10572,N_9592,N_6690);
and U10573 (N_10573,N_9540,N_7921);
nor U10574 (N_10574,N_5265,N_7424);
nand U10575 (N_10575,N_5274,N_9863);
xor U10576 (N_10576,N_8555,N_7023);
nand U10577 (N_10577,N_5862,N_9679);
and U10578 (N_10578,N_9728,N_8372);
nand U10579 (N_10579,N_6332,N_7341);
xor U10580 (N_10580,N_7870,N_9921);
and U10581 (N_10581,N_8879,N_6679);
nor U10582 (N_10582,N_9774,N_5111);
or U10583 (N_10583,N_5735,N_5830);
or U10584 (N_10584,N_6533,N_9593);
or U10585 (N_10585,N_5985,N_7606);
xor U10586 (N_10586,N_9567,N_6955);
nor U10587 (N_10587,N_9922,N_6950);
nand U10588 (N_10588,N_8960,N_6849);
xnor U10589 (N_10589,N_5364,N_5513);
nand U10590 (N_10590,N_5222,N_5429);
nor U10591 (N_10591,N_7855,N_7633);
or U10592 (N_10592,N_7953,N_8182);
and U10593 (N_10593,N_5365,N_6008);
xor U10594 (N_10594,N_6089,N_5294);
or U10595 (N_10595,N_6445,N_7049);
nand U10596 (N_10596,N_7279,N_9737);
or U10597 (N_10597,N_6947,N_5908);
and U10598 (N_10598,N_9520,N_9276);
nand U10599 (N_10599,N_9462,N_5984);
or U10600 (N_10600,N_6135,N_6090);
nand U10601 (N_10601,N_5747,N_9372);
nand U10602 (N_10602,N_5374,N_9624);
and U10603 (N_10603,N_8417,N_6015);
nand U10604 (N_10604,N_5233,N_5969);
or U10605 (N_10605,N_5667,N_6959);
nand U10606 (N_10606,N_8315,N_7037);
xor U10607 (N_10607,N_7055,N_5330);
or U10608 (N_10608,N_9274,N_5319);
nor U10609 (N_10609,N_8770,N_8126);
or U10610 (N_10610,N_8572,N_6610);
nand U10611 (N_10611,N_9739,N_5881);
or U10612 (N_10612,N_9767,N_8462);
nand U10613 (N_10613,N_5110,N_7871);
nand U10614 (N_10614,N_5889,N_8811);
nor U10615 (N_10615,N_8214,N_8509);
nand U10616 (N_10616,N_5809,N_6818);
nand U10617 (N_10617,N_5253,N_9266);
xnor U10618 (N_10618,N_7654,N_6017);
nand U10619 (N_10619,N_7709,N_5571);
and U10620 (N_10620,N_6065,N_5258);
xnor U10621 (N_10621,N_9105,N_8271);
and U10622 (N_10622,N_6949,N_6844);
nor U10623 (N_10623,N_5942,N_9267);
and U10624 (N_10624,N_9387,N_6563);
nand U10625 (N_10625,N_5277,N_7623);
and U10626 (N_10626,N_6995,N_6788);
xnor U10627 (N_10627,N_5290,N_5341);
nand U10628 (N_10628,N_8402,N_6881);
or U10629 (N_10629,N_8734,N_7125);
and U10630 (N_10630,N_8528,N_6723);
xor U10631 (N_10631,N_8862,N_6889);
nor U10632 (N_10632,N_7981,N_9927);
nand U10633 (N_10633,N_8512,N_5086);
xnor U10634 (N_10634,N_5944,N_5806);
xor U10635 (N_10635,N_6155,N_8773);
and U10636 (N_10636,N_7106,N_5435);
nand U10637 (N_10637,N_8467,N_8186);
and U10638 (N_10638,N_8810,N_6521);
and U10639 (N_10639,N_7073,N_8709);
nor U10640 (N_10640,N_9965,N_8816);
nor U10641 (N_10641,N_6264,N_7360);
nor U10642 (N_10642,N_5420,N_5645);
nand U10643 (N_10643,N_8225,N_6978);
nand U10644 (N_10644,N_8280,N_9096);
or U10645 (N_10645,N_9346,N_9039);
nor U10646 (N_10646,N_6262,N_8603);
and U10647 (N_10647,N_6325,N_9583);
nand U10648 (N_10648,N_5666,N_7332);
xnor U10649 (N_10649,N_6534,N_7772);
or U10650 (N_10650,N_8053,N_7818);
or U10651 (N_10651,N_5706,N_5731);
and U10652 (N_10652,N_8454,N_7941);
nand U10653 (N_10653,N_8544,N_6437);
xor U10654 (N_10654,N_5722,N_6411);
nor U10655 (N_10655,N_5281,N_5232);
or U10656 (N_10656,N_8902,N_7983);
and U10657 (N_10657,N_9692,N_7013);
xnor U10658 (N_10658,N_7830,N_9393);
and U10659 (N_10659,N_7119,N_7088);
and U10660 (N_10660,N_8012,N_5529);
xor U10661 (N_10661,N_8220,N_7206);
xnor U10662 (N_10662,N_7491,N_8348);
or U10663 (N_10663,N_6713,N_7413);
and U10664 (N_10664,N_8150,N_5073);
or U10665 (N_10665,N_7306,N_8045);
or U10666 (N_10666,N_7223,N_8701);
nor U10667 (N_10667,N_6148,N_8723);
and U10668 (N_10668,N_9134,N_7255);
nand U10669 (N_10669,N_9400,N_9643);
or U10670 (N_10670,N_7027,N_8631);
or U10671 (N_10671,N_7592,N_9759);
nand U10672 (N_10672,N_5817,N_9198);
nor U10673 (N_10673,N_5869,N_7477);
xnor U10674 (N_10674,N_6632,N_7262);
xnor U10675 (N_10675,N_9917,N_8610);
nor U10676 (N_10676,N_8305,N_7047);
nor U10677 (N_10677,N_7699,N_7144);
and U10678 (N_10678,N_8008,N_9195);
or U10679 (N_10679,N_5588,N_8435);
nor U10680 (N_10680,N_9416,N_7556);
or U10681 (N_10681,N_8671,N_9909);
xor U10682 (N_10682,N_5229,N_9947);
xor U10683 (N_10683,N_6803,N_5367);
and U10684 (N_10684,N_9187,N_5874);
or U10685 (N_10685,N_5242,N_9821);
nor U10686 (N_10686,N_7854,N_9557);
nor U10687 (N_10687,N_8159,N_7344);
and U10688 (N_10688,N_8988,N_5467);
or U10689 (N_10689,N_8852,N_5063);
nor U10690 (N_10690,N_5463,N_9010);
xnor U10691 (N_10691,N_6820,N_8896);
or U10692 (N_10692,N_5794,N_5426);
xor U10693 (N_10693,N_8539,N_7343);
xor U10694 (N_10694,N_7573,N_6636);
nor U10695 (N_10695,N_8197,N_5241);
nand U10696 (N_10696,N_9526,N_8848);
xnor U10697 (N_10697,N_5860,N_7467);
and U10698 (N_10698,N_7105,N_7046);
nor U10699 (N_10699,N_5142,N_8501);
or U10700 (N_10700,N_5015,N_7191);
or U10701 (N_10701,N_7082,N_6840);
and U10702 (N_10702,N_8767,N_9764);
or U10703 (N_10703,N_6434,N_5515);
or U10704 (N_10704,N_5392,N_9214);
xnor U10705 (N_10705,N_6989,N_6708);
nand U10706 (N_10706,N_5120,N_5116);
or U10707 (N_10707,N_8788,N_9009);
or U10708 (N_10708,N_7991,N_5276);
nor U10709 (N_10709,N_5844,N_5079);
and U10710 (N_10710,N_8013,N_8843);
xor U10711 (N_10711,N_7956,N_9287);
nor U10712 (N_10712,N_8062,N_7554);
nor U10713 (N_10713,N_5974,N_5749);
nand U10714 (N_10714,N_6591,N_5866);
nor U10715 (N_10715,N_8590,N_8076);
or U10716 (N_10716,N_8407,N_9800);
nor U10717 (N_10717,N_7795,N_9742);
nand U10718 (N_10718,N_8495,N_6974);
or U10719 (N_10719,N_9788,N_7801);
and U10720 (N_10720,N_8030,N_5402);
nor U10721 (N_10721,N_7507,N_8298);
nand U10722 (N_10722,N_7032,N_9205);
nand U10723 (N_10723,N_8192,N_6890);
or U10724 (N_10724,N_6761,N_9348);
nor U10725 (N_10725,N_5488,N_7451);
xnor U10726 (N_10726,N_5247,N_9024);
nand U10727 (N_10727,N_7541,N_7807);
or U10728 (N_10728,N_7912,N_6514);
or U10729 (N_10729,N_9450,N_7251);
nand U10730 (N_10730,N_8361,N_6182);
nand U10731 (N_10731,N_8558,N_7798);
or U10732 (N_10732,N_8952,N_9104);
nor U10733 (N_10733,N_8201,N_9386);
nand U10734 (N_10734,N_5799,N_9138);
xor U10735 (N_10735,N_9883,N_7308);
and U10736 (N_10736,N_8127,N_5552);
or U10737 (N_10737,N_5112,N_6478);
or U10738 (N_10738,N_6724,N_6614);
and U10739 (N_10739,N_8808,N_6209);
or U10740 (N_10740,N_7216,N_9094);
nor U10741 (N_10741,N_8108,N_6501);
nand U10742 (N_10742,N_7609,N_7674);
nor U10743 (N_10743,N_6740,N_8983);
and U10744 (N_10744,N_7627,N_8430);
or U10745 (N_10745,N_6406,N_8761);
and U10746 (N_10746,N_8834,N_9293);
xnor U10747 (N_10747,N_6864,N_8246);
xor U10748 (N_10748,N_9670,N_6131);
nor U10749 (N_10749,N_7179,N_8806);
or U10750 (N_10750,N_7379,N_6428);
nor U10751 (N_10751,N_9999,N_7542);
nand U10752 (N_10752,N_9906,N_6527);
nor U10753 (N_10753,N_7715,N_6711);
and U10754 (N_10754,N_5509,N_7256);
nand U10755 (N_10755,N_6542,N_6562);
and U10756 (N_10756,N_6580,N_5778);
and U10757 (N_10757,N_6429,N_8029);
nor U10758 (N_10758,N_9958,N_5123);
and U10759 (N_10759,N_7769,N_5125);
nand U10760 (N_10760,N_5574,N_7244);
or U10761 (N_10761,N_9253,N_8612);
xnor U10762 (N_10762,N_5814,N_6391);
nand U10763 (N_10763,N_6007,N_7026);
or U10764 (N_10764,N_5796,N_5157);
and U10765 (N_10765,N_7404,N_6261);
xnor U10766 (N_10766,N_7810,N_9262);
xnor U10767 (N_10767,N_5119,N_8725);
and U10768 (N_10768,N_6805,N_9681);
and U10769 (N_10769,N_6606,N_7163);
and U10770 (N_10770,N_9482,N_8106);
nand U10771 (N_10771,N_7313,N_9628);
and U10772 (N_10772,N_9016,N_7156);
or U10773 (N_10773,N_6004,N_5263);
and U10774 (N_10774,N_8736,N_5587);
nor U10775 (N_10775,N_9131,N_6497);
and U10776 (N_10776,N_5635,N_7416);
or U10777 (N_10777,N_6920,N_9243);
nand U10778 (N_10778,N_8792,N_5450);
nand U10779 (N_10779,N_9761,N_6327);
xor U10780 (N_10780,N_7545,N_8711);
or U10781 (N_10781,N_8270,N_7789);
and U10782 (N_10782,N_7559,N_6374);
nor U10783 (N_10783,N_7934,N_6412);
nor U10784 (N_10784,N_5159,N_9413);
and U10785 (N_10785,N_9580,N_5130);
or U10786 (N_10786,N_8234,N_5296);
nor U10787 (N_10787,N_9641,N_9740);
nor U10788 (N_10788,N_9689,N_6684);
nor U10789 (N_10789,N_9164,N_7455);
or U10790 (N_10790,N_5268,N_7681);
nand U10791 (N_10791,N_9891,N_5988);
xnor U10792 (N_10792,N_9723,N_7274);
nor U10793 (N_10793,N_9674,N_6615);
xnor U10794 (N_10794,N_7982,N_8757);
nor U10795 (N_10795,N_6704,N_8968);
xor U10796 (N_10796,N_6887,N_6846);
nor U10797 (N_10797,N_6698,N_6006);
nand U10798 (N_10798,N_7131,N_5389);
nand U10799 (N_10799,N_6737,N_9448);
nor U10800 (N_10800,N_8100,N_9952);
or U10801 (N_10801,N_5567,N_5353);
nor U10802 (N_10802,N_7175,N_8931);
nor U10803 (N_10803,N_7875,N_8964);
and U10804 (N_10804,N_6470,N_9655);
and U10805 (N_10805,N_6620,N_5022);
nand U10806 (N_10806,N_9193,N_6800);
and U10807 (N_10807,N_9380,N_5132);
or U10808 (N_10808,N_7960,N_6555);
nor U10809 (N_10809,N_7895,N_7048);
nand U10810 (N_10810,N_7969,N_9259);
nand U10811 (N_10811,N_5168,N_5804);
nand U10812 (N_10812,N_7441,N_7024);
nand U10813 (N_10813,N_5759,N_5359);
xnor U10814 (N_10814,N_6482,N_5419);
and U10815 (N_10815,N_8146,N_6666);
nor U10816 (N_10816,N_9103,N_7793);
nand U10817 (N_10817,N_9360,N_5334);
xor U10818 (N_10818,N_9235,N_9021);
and U10819 (N_10819,N_6556,N_8222);
and U10820 (N_10820,N_8422,N_6286);
nand U10821 (N_10821,N_9804,N_5433);
nand U10822 (N_10822,N_8088,N_7864);
and U10823 (N_10823,N_9089,N_6179);
nor U10824 (N_10824,N_6913,N_6931);
nand U10825 (N_10825,N_9996,N_6641);
nand U10826 (N_10826,N_5815,N_8034);
nor U10827 (N_10827,N_6899,N_6669);
xor U10828 (N_10828,N_7038,N_8482);
xnor U10829 (N_10829,N_8858,N_7717);
and U10830 (N_10830,N_5451,N_8457);
and U10831 (N_10831,N_7068,N_7225);
xnor U10832 (N_10832,N_7300,N_6965);
nand U10833 (N_10833,N_5163,N_5155);
and U10834 (N_10834,N_7678,N_8050);
xnor U10835 (N_10835,N_8195,N_5272);
nor U10836 (N_10836,N_9137,N_9412);
xnor U10837 (N_10837,N_5411,N_5245);
xor U10838 (N_10838,N_9488,N_7802);
xnor U10839 (N_10839,N_7498,N_8168);
or U10840 (N_10840,N_7164,N_6607);
and U10841 (N_10841,N_5236,N_9838);
nand U10842 (N_10842,N_7616,N_8774);
or U10843 (N_10843,N_8726,N_8096);
xnor U10844 (N_10844,N_6914,N_6670);
or U10845 (N_10845,N_6180,N_5207);
and U10846 (N_10846,N_7427,N_6807);
or U10847 (N_10847,N_7168,N_8943);
or U10848 (N_10848,N_7955,N_8370);
xor U10849 (N_10849,N_6998,N_8957);
nor U10850 (N_10850,N_8541,N_7790);
nand U10851 (N_10851,N_7995,N_9955);
nor U10852 (N_10852,N_8829,N_7463);
xor U10853 (N_10853,N_6771,N_6672);
nor U10854 (N_10854,N_6505,N_7433);
nor U10855 (N_10855,N_6446,N_5754);
and U10856 (N_10856,N_7412,N_5964);
and U10857 (N_10857,N_9607,N_8801);
nor U10858 (N_10858,N_5980,N_6425);
xor U10859 (N_10859,N_9859,N_6648);
and U10860 (N_10860,N_9846,N_7292);
xor U10861 (N_10861,N_6862,N_5863);
nand U10862 (N_10862,N_7098,N_6897);
nor U10863 (N_10863,N_7832,N_9713);
nand U10864 (N_10864,N_7436,N_6824);
xnor U10865 (N_10865,N_9599,N_6687);
or U10866 (N_10866,N_8160,N_9910);
nand U10867 (N_10867,N_7930,N_5507);
nand U10868 (N_10868,N_8549,N_5092);
and U10869 (N_10869,N_6276,N_6314);
and U10870 (N_10870,N_9300,N_8795);
or U10871 (N_10871,N_8940,N_8463);
xnor U10872 (N_10872,N_6600,N_9112);
and U10873 (N_10873,N_7004,N_6516);
nor U10874 (N_10874,N_5713,N_6456);
xnor U10875 (N_10875,N_8899,N_7411);
and U10876 (N_10876,N_5704,N_6043);
nand U10877 (N_10877,N_6561,N_7489);
xnor U10878 (N_10878,N_8685,N_6535);
nand U10879 (N_10879,N_8639,N_7778);
nor U10880 (N_10880,N_5502,N_9154);
nand U10881 (N_10881,N_9877,N_8025);
nor U10882 (N_10882,N_7260,N_5518);
nor U10883 (N_10883,N_5029,N_9015);
nor U10884 (N_10884,N_6002,N_6153);
and U10885 (N_10885,N_6652,N_7547);
nor U10886 (N_10886,N_6634,N_9129);
nand U10887 (N_10887,N_9044,N_7642);
xor U10888 (N_10888,N_6280,N_5052);
xnor U10889 (N_10889,N_9573,N_5191);
or U10890 (N_10890,N_8288,N_8419);
or U10891 (N_10891,N_7605,N_5658);
or U10892 (N_10892,N_5913,N_7971);
nand U10893 (N_10893,N_5549,N_8682);
xor U10894 (N_10894,N_9509,N_8911);
and U10895 (N_10895,N_7740,N_5622);
nor U10896 (N_10896,N_6253,N_8125);
nor U10897 (N_10897,N_7696,N_9365);
and U10898 (N_10898,N_8922,N_7667);
nand U10899 (N_10899,N_5598,N_6278);
xor U10900 (N_10900,N_6282,N_9902);
or U10901 (N_10901,N_9908,N_9773);
and U10902 (N_10902,N_7431,N_7293);
nand U10903 (N_10903,N_7655,N_8377);
and U10904 (N_10904,N_6838,N_5816);
nand U10905 (N_10905,N_8003,N_6686);
nor U10906 (N_10906,N_6000,N_7967);
or U10907 (N_10907,N_9813,N_9717);
and U10908 (N_10908,N_9941,N_7084);
nand U10909 (N_10909,N_7050,N_6175);
nand U10910 (N_10910,N_7533,N_8756);
nand U10911 (N_10911,N_7569,N_6835);
and U10912 (N_10912,N_6537,N_9660);
or U10913 (N_10913,N_8600,N_6117);
xnor U10914 (N_10914,N_8193,N_8043);
or U10915 (N_10915,N_5066,N_7827);
nor U10916 (N_10916,N_8327,N_5175);
nand U10917 (N_10917,N_5914,N_7684);
nor U10918 (N_10918,N_6404,N_5926);
or U10919 (N_10919,N_7367,N_7711);
and U10920 (N_10920,N_7638,N_5303);
and U10921 (N_10921,N_7445,N_7196);
or U10922 (N_10922,N_7639,N_6100);
and U10923 (N_10923,N_6303,N_5548);
or U10924 (N_10924,N_9207,N_5572);
or U10925 (N_10925,N_7993,N_6188);
xor U10926 (N_10926,N_7030,N_9832);
and U10927 (N_10927,N_7180,N_8074);
nand U10928 (N_10928,N_9498,N_9991);
or U10929 (N_10929,N_9830,N_6883);
and U10930 (N_10930,N_6882,N_6894);
or U10931 (N_10931,N_6095,N_6635);
or U10932 (N_10932,N_8958,N_9391);
xor U10933 (N_10933,N_6979,N_7459);
or U10934 (N_10934,N_7029,N_6550);
or U10935 (N_10935,N_5322,N_9729);
and U10936 (N_10936,N_8200,N_7326);
nand U10937 (N_10937,N_5380,N_7957);
nand U10938 (N_10938,N_7999,N_6019);
nor U10939 (N_10939,N_8099,N_7776);
and U10940 (N_10940,N_9273,N_6617);
nand U10941 (N_10941,N_8938,N_9811);
or U10942 (N_10942,N_8889,N_9673);
xnor U10943 (N_10943,N_9063,N_7922);
and U10944 (N_10944,N_7336,N_8124);
nand U10945 (N_10945,N_5812,N_8475);
nand U10946 (N_10946,N_8460,N_6510);
nor U10947 (N_10947,N_5585,N_6333);
or U10948 (N_10948,N_9457,N_9961);
xnor U10949 (N_10949,N_5376,N_6757);
nand U10950 (N_10950,N_6395,N_5228);
nor U10951 (N_10951,N_6309,N_6230);
or U10952 (N_10952,N_8420,N_6594);
and U10953 (N_10953,N_6928,N_8006);
nand U10954 (N_10954,N_9111,N_7961);
nor U10955 (N_10955,N_8656,N_7781);
nand U10956 (N_10956,N_5600,N_9810);
xor U10957 (N_10957,N_6217,N_8093);
or U10958 (N_10958,N_8926,N_7219);
and U10959 (N_10959,N_9209,N_7176);
nor U10960 (N_10960,N_6074,N_5430);
and U10961 (N_10961,N_7148,N_5682);
nand U10962 (N_10962,N_8026,N_5981);
or U10963 (N_10963,N_7208,N_7070);
xnor U10964 (N_10964,N_8507,N_9653);
xor U10965 (N_10965,N_9865,N_8058);
xnor U10966 (N_10966,N_7399,N_7691);
and U10967 (N_10967,N_9635,N_7659);
nor U10968 (N_10968,N_7614,N_9625);
nand U10969 (N_10969,N_8438,N_5386);
xnor U10970 (N_10970,N_6854,N_8335);
or U10971 (N_10971,N_6283,N_5395);
nor U10972 (N_10972,N_5727,N_5930);
or U10973 (N_10973,N_5478,N_5730);
or U10974 (N_10974,N_5101,N_6732);
xor U10975 (N_10975,N_9888,N_5139);
or U10976 (N_10976,N_6814,N_5234);
or U10977 (N_10977,N_9234,N_7891);
and U10978 (N_10978,N_7327,N_9184);
or U10979 (N_10979,N_8052,N_7645);
nor U10980 (N_10980,N_5349,N_5218);
or U10981 (N_10981,N_7154,N_6812);
nand U10982 (N_10982,N_6250,N_6895);
and U10983 (N_10983,N_7414,N_9303);
nand U10984 (N_10984,N_5399,N_6752);
and U10985 (N_10985,N_8961,N_9383);
or U10986 (N_10986,N_8065,N_5370);
nor U10987 (N_10987,N_9124,N_6483);
xor U10988 (N_10988,N_9998,N_5179);
or U10989 (N_10989,N_8629,N_9829);
nor U10990 (N_10990,N_8683,N_8888);
and U10991 (N_10991,N_9421,N_5398);
nor U10992 (N_10992,N_6364,N_9836);
nand U10993 (N_10993,N_6822,N_5594);
nor U10994 (N_10994,N_7375,N_8670);
nor U10995 (N_10995,N_8129,N_6726);
and U10996 (N_10996,N_8235,N_8869);
xnor U10997 (N_10997,N_9248,N_5750);
nor U10998 (N_10998,N_8284,N_6629);
and U10999 (N_10999,N_9600,N_9001);
xnor U11000 (N_11000,N_5442,N_7927);
and U11001 (N_11001,N_9326,N_5922);
or U11002 (N_11002,N_6133,N_5606);
nand U11003 (N_11003,N_6765,N_9064);
xnor U11004 (N_11004,N_8728,N_7092);
nand U11005 (N_11005,N_7710,N_9598);
or U11006 (N_11006,N_6433,N_5094);
and U11007 (N_11007,N_9396,N_9864);
nor U11008 (N_11008,N_5764,N_5776);
or U11009 (N_11009,N_9976,N_9849);
and U11010 (N_11010,N_6256,N_5331);
nor U11011 (N_11011,N_7237,N_9070);
and U11012 (N_11012,N_6234,N_7511);
or U11013 (N_11013,N_5708,N_7977);
and U11014 (N_11014,N_7328,N_5206);
and U11015 (N_11015,N_9463,N_7276);
and U11016 (N_11016,N_9803,N_7612);
nor U11017 (N_11017,N_7473,N_9046);
and U11018 (N_11018,N_8620,N_6106);
xor U11019 (N_11019,N_7817,N_8717);
nand U11020 (N_11020,N_6530,N_8016);
and U11021 (N_11021,N_8865,N_6892);
nand U11022 (N_11022,N_8878,N_5724);
or U11023 (N_11023,N_8057,N_8497);
nand U11024 (N_11024,N_5396,N_7025);
or U11025 (N_11025,N_8547,N_7679);
or U11026 (N_11026,N_5763,N_9435);
xnor U11027 (N_11027,N_9459,N_7268);
and U11028 (N_11028,N_8410,N_6587);
xor U11029 (N_11029,N_5975,N_6397);
nand U11030 (N_11030,N_9933,N_7758);
nor U11031 (N_11031,N_7390,N_8300);
nand U11032 (N_11032,N_7792,N_7096);
xor U11033 (N_11033,N_7663,N_5556);
nand U11034 (N_11034,N_8444,N_8892);
and U11035 (N_11035,N_8740,N_6500);
xnor U11036 (N_11036,N_8796,N_5602);
xnor U11037 (N_11037,N_7348,N_8114);
nor U11038 (N_11038,N_7813,N_6937);
nor U11039 (N_11039,N_5219,N_9651);
or U11040 (N_11040,N_7066,N_8172);
or U11041 (N_11041,N_9121,N_9093);
or U11042 (N_11042,N_7590,N_5621);
nor U11043 (N_11043,N_7845,N_7899);
or U11044 (N_11044,N_8667,N_6655);
xnor U11045 (N_11045,N_7307,N_5362);
xnor U11046 (N_11046,N_7517,N_9460);
xor U11047 (N_11047,N_6665,N_9636);
nand U11048 (N_11048,N_7693,N_9576);
nor U11049 (N_11049,N_9532,N_9066);
or U11050 (N_11050,N_6001,N_5214);
or U11051 (N_11051,N_6306,N_9746);
xnor U11052 (N_11052,N_7860,N_6381);
nor U11053 (N_11053,N_8991,N_5689);
nand U11054 (N_11054,N_8920,N_9696);
and U11055 (N_11055,N_8518,N_6167);
nand U11056 (N_11056,N_7868,N_8666);
or U11057 (N_11057,N_5193,N_8953);
xor U11058 (N_11058,N_8135,N_5494);
nor U11059 (N_11059,N_9376,N_7782);
nor U11060 (N_11060,N_7437,N_7671);
nor U11061 (N_11061,N_6330,N_9978);
xnor U11062 (N_11062,N_6013,N_9469);
nor U11063 (N_11063,N_7874,N_9275);
and U11064 (N_11064,N_8414,N_5424);
or U11065 (N_11065,N_9712,N_9777);
nor U11066 (N_11066,N_7249,N_5781);
nand U11067 (N_11067,N_8598,N_6836);
or U11068 (N_11068,N_9118,N_8854);
or U11069 (N_11069,N_7937,N_6444);
nand U11070 (N_11070,N_5038,N_9054);
nor U11071 (N_11071,N_9100,N_7851);
and U11072 (N_11072,N_7516,N_6676);
and U11073 (N_11073,N_8585,N_7396);
or U11074 (N_11074,N_9897,N_5064);
and U11075 (N_11075,N_7962,N_9946);
or U11076 (N_11076,N_6870,N_5915);
nand U11077 (N_11077,N_6848,N_8503);
or U11078 (N_11078,N_5608,N_5971);
and U11079 (N_11079,N_6569,N_7273);
xnor U11080 (N_11080,N_8751,N_7394);
and U11081 (N_11081,N_7766,N_5400);
nor U11082 (N_11082,N_8784,N_9373);
or U11083 (N_11083,N_5388,N_9294);
nand U11084 (N_11084,N_6247,N_6187);
nand U11085 (N_11085,N_8619,N_9098);
nand U11086 (N_11086,N_9618,N_9577);
or U11087 (N_11087,N_6149,N_6962);
or U11088 (N_11088,N_5474,N_8081);
nand U11089 (N_11089,N_5127,N_8613);
nand U11090 (N_11090,N_8277,N_9687);
nor U11091 (N_11091,N_6246,N_6054);
and U11092 (N_11092,N_6796,N_7823);
or U11093 (N_11093,N_7202,N_6681);
and U11094 (N_11094,N_5511,N_8198);
nor U11095 (N_11095,N_9566,N_6093);
xor U11096 (N_11096,N_6551,N_8566);
nand U11097 (N_11097,N_6787,N_9718);
nor U11098 (N_11098,N_7143,N_6291);
and U11099 (N_11099,N_8979,N_9197);
xor U11100 (N_11100,N_8814,N_8924);
or U11101 (N_11101,N_8815,N_5824);
xor U11102 (N_11102,N_5791,N_8586);
xor U11103 (N_11103,N_9915,N_5591);
xnor U11104 (N_11104,N_7128,N_9930);
and U11105 (N_11105,N_7161,N_9548);
nand U11106 (N_11106,N_9246,N_7508);
nand U11107 (N_11107,N_7800,N_5887);
and U11108 (N_11108,N_9882,N_9586);
nor U11109 (N_11109,N_9005,N_5962);
and U11110 (N_11110,N_8556,N_6673);
nor U11111 (N_11111,N_5267,N_7203);
and U11112 (N_11112,N_5715,N_8601);
xor U11113 (N_11113,N_8326,N_8655);
xnor U11114 (N_11114,N_7712,N_9812);
and U11115 (N_11115,N_7117,N_8387);
nand U11116 (N_11116,N_5868,N_6705);
or U11117 (N_11117,N_7848,N_9986);
nand U11118 (N_11118,N_7587,N_6042);
xor U11119 (N_11119,N_5212,N_9700);
nand U11120 (N_11120,N_8199,N_9114);
nor U11121 (N_11121,N_7232,N_8496);
or U11122 (N_11122,N_7599,N_8543);
and U11123 (N_11123,N_7908,N_8876);
xnor U11124 (N_11124,N_5711,N_9337);
or U11125 (N_11125,N_9370,N_8347);
and U11126 (N_11126,N_9831,N_6473);
and U11127 (N_11127,N_8999,N_6222);
nand U11128 (N_11128,N_9301,N_8176);
nand U11129 (N_11129,N_7040,N_8278);
and U11130 (N_11130,N_8359,N_5786);
and U11131 (N_11131,N_9344,N_6072);
nand U11132 (N_11132,N_9322,N_8320);
nor U11133 (N_11133,N_9148,N_9320);
xnor U11134 (N_11134,N_9959,N_8428);
xnor U11135 (N_11135,N_6157,N_5718);
and U11136 (N_11136,N_9756,N_7535);
xnor U11137 (N_11137,N_9473,N_5681);
and U11138 (N_11138,N_6872,N_7063);
or U11139 (N_11139,N_7553,N_8912);
or U11140 (N_11140,N_6018,N_6896);
nor U11141 (N_11141,N_5471,N_6795);
or U11142 (N_11142,N_8263,N_8721);
or U11143 (N_11143,N_6588,N_8738);
xor U11144 (N_11144,N_6233,N_6618);
or U11145 (N_11145,N_6236,N_9374);
xnor U11146 (N_11146,N_7557,N_8514);
nand U11147 (N_11147,N_8391,N_8449);
or U11148 (N_11148,N_6415,N_8491);
nor U11149 (N_11149,N_9519,N_9916);
or U11150 (N_11150,N_7374,N_9824);
and U11151 (N_11151,N_8056,N_6739);
nand U11152 (N_11152,N_6926,N_6033);
nand U11153 (N_11153,N_7366,N_7539);
nor U11154 (N_11154,N_5385,N_8429);
nand U11155 (N_11155,N_7915,N_9311);
nand U11156 (N_11156,N_6797,N_5489);
or U11157 (N_11157,N_7829,N_7989);
xnor U11158 (N_11158,N_6322,N_8097);
and U11159 (N_11159,N_6929,N_5967);
nor U11160 (N_11160,N_7505,N_6011);
xnor U11161 (N_11161,N_6706,N_7788);
and U11162 (N_11162,N_7465,N_6511);
and U11163 (N_11163,N_9765,N_7102);
xnor U11164 (N_11164,N_5740,N_5134);
nand U11165 (N_11165,N_8219,N_9027);
nand U11166 (N_11166,N_7732,N_7400);
nor U11167 (N_11167,N_7949,N_9637);
xnor U11168 (N_11168,N_6275,N_5849);
nand U11169 (N_11169,N_7889,N_8886);
nand U11170 (N_11170,N_7483,N_9194);
or U11171 (N_11171,N_6349,N_5238);
nor U11172 (N_11172,N_7277,N_5473);
nor U11173 (N_11173,N_5672,N_8828);
and U11174 (N_11174,N_8771,N_7670);
nor U11175 (N_11175,N_7112,N_8031);
and U11176 (N_11176,N_9220,N_8232);
nor U11177 (N_11177,N_8048,N_9151);
nand U11178 (N_11178,N_8487,N_7735);
and U11179 (N_11179,N_7785,N_5959);
and U11180 (N_11180,N_6701,N_9934);
xor U11181 (N_11181,N_6968,N_5767);
xnor U11182 (N_11182,N_5826,N_5550);
or U11183 (N_11183,N_8819,N_9180);
or U11184 (N_11184,N_5951,N_8727);
or U11185 (N_11185,N_9616,N_8576);
or U11186 (N_11186,N_9949,N_6798);
xnor U11187 (N_11187,N_7006,N_7470);
xor U11188 (N_11188,N_6725,N_5390);
xor U11189 (N_11189,N_5269,N_9270);
xor U11190 (N_11190,N_5283,N_8604);
nand U11191 (N_11191,N_7883,N_8805);
xor U11192 (N_11192,N_8046,N_8984);
nor U11193 (N_11193,N_7746,N_5717);
nand U11194 (N_11194,N_9176,N_9725);
nand U11195 (N_11195,N_5329,N_6891);
or U11196 (N_11196,N_9534,N_9890);
or U11197 (N_11197,N_8144,N_6703);
and U11198 (N_11198,N_8224,N_8887);
nand U11199 (N_11199,N_7387,N_8148);
xor U11200 (N_11200,N_6935,N_6884);
or U11201 (N_11201,N_9543,N_6038);
and U11202 (N_11202,N_5770,N_5935);
xnor U11203 (N_11203,N_8181,N_7464);
nand U11204 (N_11204,N_6097,N_8648);
or U11205 (N_11205,N_5496,N_7091);
and U11206 (N_11206,N_7019,N_5792);
and U11207 (N_11207,N_9355,N_6270);
and U11208 (N_11208,N_8068,N_8471);
nand U11209 (N_11209,N_8695,N_5224);
and U11210 (N_11210,N_6356,N_8650);
nor U11211 (N_11211,N_9744,N_8578);
nor U11212 (N_11212,N_9149,N_7016);
nor U11213 (N_11213,N_6037,N_7537);
nor U11214 (N_11214,N_5540,N_6986);
xor U11215 (N_11215,N_7409,N_8259);
nand U11216 (N_11216,N_9818,N_5252);
or U11217 (N_11217,N_5819,N_7932);
nand U11218 (N_11218,N_9332,N_5351);
nand U11219 (N_11219,N_6940,N_8531);
xor U11220 (N_11220,N_6290,N_9656);
nor U11221 (N_11221,N_7668,N_7198);
or U11222 (N_11222,N_6619,N_8170);
nor U11223 (N_11223,N_9758,N_7705);
and U11224 (N_11224,N_9935,N_8654);
or U11225 (N_11225,N_5773,N_5996);
nor U11226 (N_11226,N_6763,N_6345);
and U11227 (N_11227,N_6334,N_9445);
or U11228 (N_11228,N_7286,N_6557);
nor U11229 (N_11229,N_7028,N_9082);
nor U11230 (N_11230,N_6774,N_7471);
or U11231 (N_11231,N_7472,N_7384);
xor U11232 (N_11232,N_7151,N_7177);
or U11233 (N_11233,N_8625,N_8554);
nand U11234 (N_11234,N_9750,N_7604);
nor U11235 (N_11235,N_8386,N_7975);
nand U11236 (N_11236,N_7212,N_8614);
and U11237 (N_11237,N_7017,N_9389);
or U11238 (N_11238,N_5953,N_5301);
nand U11239 (N_11239,N_5328,N_6873);
nand U11240 (N_11240,N_9011,N_5626);
nand U11241 (N_11241,N_5811,N_8105);
and U11242 (N_11242,N_6403,N_8597);
and U11243 (N_11243,N_5054,N_5045);
and U11244 (N_11244,N_7856,N_5895);
xnor U11245 (N_11245,N_5519,N_5192);
xnor U11246 (N_11246,N_9072,N_8292);
xor U11247 (N_11247,N_8469,N_5476);
xor U11248 (N_11248,N_9165,N_7373);
and U11249 (N_11249,N_6335,N_5783);
xor U11250 (N_11250,N_5891,N_7532);
or U11251 (N_11251,N_8102,N_5318);
and U11252 (N_11252,N_8360,N_5288);
nand U11253 (N_11253,N_9867,N_9414);
and U11254 (N_11254,N_6020,N_5609);
and U11255 (N_11255,N_5543,N_8662);
and U11256 (N_11256,N_5166,N_7421);
and U11257 (N_11257,N_6475,N_7456);
xnor U11258 (N_11258,N_8652,N_6692);
nor U11259 (N_11259,N_8466,N_7660);
nor U11260 (N_11260,N_8692,N_7204);
nor U11261 (N_11261,N_6195,N_5039);
nand U11262 (N_11262,N_5449,N_9221);
xor U11263 (N_11263,N_8445,N_7935);
nand U11264 (N_11264,N_5285,N_6347);
nor U11265 (N_11265,N_8955,N_5675);
or U11266 (N_11266,N_8260,N_7487);
and U11267 (N_11267,N_6651,N_6758);
nor U11268 (N_11268,N_9779,N_7356);
xor U11269 (N_11269,N_7067,N_9556);
or U11270 (N_11270,N_9201,N_9572);
and U11271 (N_11271,N_7018,N_9035);
xor U11272 (N_11272,N_6422,N_8678);
nor U11273 (N_11273,N_9216,N_5558);
or U11274 (N_11274,N_5679,N_6689);
nor U11275 (N_11275,N_6073,N_7904);
nand U11276 (N_11276,N_9338,N_5382);
xnor U11277 (N_11277,N_8608,N_7576);
nand U11278 (N_11278,N_6987,N_6566);
and U11279 (N_11279,N_7543,N_7079);
xnor U11280 (N_11280,N_6938,N_7568);
xnor U11281 (N_11281,N_8123,N_9588);
or U11282 (N_11282,N_6727,N_6154);
or U11283 (N_11283,N_8212,N_9426);
or U11284 (N_11284,N_6863,N_5048);
xor U11285 (N_11285,N_7869,N_5554);
or U11286 (N_11286,N_8338,N_5625);
and U11287 (N_11287,N_6823,N_8171);
nor U11288 (N_11288,N_8312,N_8971);
xnor U11289 (N_11289,N_5997,N_5043);
nor U11290 (N_11290,N_6128,N_8077);
nand U11291 (N_11291,N_8898,N_8588);
nor U11292 (N_11292,N_6512,N_6005);
and U11293 (N_11293,N_6393,N_6083);
and U11294 (N_11294,N_8856,N_8906);
and U11295 (N_11295,N_9584,N_5297);
nor U11296 (N_11296,N_9238,N_8227);
and U11297 (N_11297,N_5172,N_8615);
or U11298 (N_11298,N_6799,N_8686);
nand U11299 (N_11299,N_9002,N_8573);
and U11300 (N_11300,N_7974,N_8389);
or U11301 (N_11301,N_9605,N_6810);
nor U11302 (N_11302,N_9617,N_9962);
nand U11303 (N_11303,N_5611,N_8737);
and U11304 (N_11304,N_6571,N_6728);
nand U11305 (N_11305,N_9321,N_5743);
nand U11306 (N_11306,N_5662,N_5968);
xor U11307 (N_11307,N_5961,N_5536);
xnor U11308 (N_11308,N_7918,N_8229);
xor U11309 (N_11309,N_8949,N_8375);
nand U11310 (N_11310,N_9639,N_5026);
xor U11311 (N_11311,N_6980,N_6027);
xnor U11312 (N_11312,N_8551,N_7265);
xnor U11313 (N_11313,N_9188,N_5676);
xnor U11314 (N_11314,N_7003,N_7007);
nand U11315 (N_11315,N_7488,N_6066);
xor U11316 (N_11316,N_5197,N_9889);
and U11317 (N_11317,N_5801,N_8748);
nor U11318 (N_11318,N_5528,N_6794);
xor U11319 (N_11319,N_9237,N_5756);
and U11320 (N_11320,N_9511,N_8798);
nor U11321 (N_11321,N_8841,N_6492);
xnor U11322 (N_11322,N_5709,N_6172);
and U11323 (N_11323,N_7812,N_9510);
and U11324 (N_11324,N_5932,N_9306);
nand U11325 (N_11325,N_5248,N_7850);
xnor U11326 (N_11326,N_9230,N_5733);
nand U11327 (N_11327,N_8208,N_8281);
nand U11328 (N_11328,N_7228,N_8090);
or U11329 (N_11329,N_9109,N_6650);
xor U11330 (N_11330,N_7171,N_7862);
nor U11331 (N_11331,N_9356,N_7311);
and U11332 (N_11332,N_9477,N_8907);
nor U11333 (N_11333,N_9327,N_5818);
nor U11334 (N_11334,N_6373,N_7109);
or U11335 (N_11335,N_9848,N_5147);
and U11336 (N_11336,N_6375,N_6625);
xor U11337 (N_11337,N_6039,N_7574);
nor U11338 (N_11338,N_9127,N_9088);
xnor U11339 (N_11339,N_7558,N_8484);
or U11340 (N_11340,N_6513,N_5311);
and U11341 (N_11341,N_9852,N_6970);
or U11342 (N_11342,N_5203,N_5405);
nor U11343 (N_11343,N_6660,N_6416);
nand U11344 (N_11344,N_8005,N_8855);
nor U11345 (N_11345,N_8230,N_8832);
xor U11346 (N_11346,N_9912,N_8799);
nand U11347 (N_11347,N_8308,N_5428);
nand U11348 (N_11348,N_9404,N_8364);
nor U11349 (N_11349,N_8645,N_9161);
nand U11350 (N_11350,N_7768,N_6816);
nor U11351 (N_11351,N_9368,N_8732);
xnor U11352 (N_11352,N_9979,N_5299);
xnor U11353 (N_11353,N_8297,N_9704);
nand U11354 (N_11354,N_7183,N_6479);
nand U11355 (N_11355,N_6420,N_5810);
nand U11356 (N_11356,N_8427,N_8118);
xor U11357 (N_11357,N_7221,N_5347);
xor U11358 (N_11358,N_5354,N_7454);
nand U11359 (N_11359,N_5149,N_9895);
xnor U11360 (N_11360,N_5051,N_7566);
nor U11361 (N_11361,N_8409,N_6160);
nand U11362 (N_11362,N_8448,N_5004);
and U11363 (N_11363,N_8080,N_9493);
xnor U11364 (N_11364,N_7479,N_5545);
nor U11365 (N_11365,N_7466,N_6667);
xor U11366 (N_11366,N_5183,N_6582);
nand U11367 (N_11367,N_9312,N_7494);
nor U11368 (N_11368,N_9964,N_8242);
xnor U11369 (N_11369,N_8228,N_9619);
xnor U11370 (N_11370,N_6664,N_5089);
xnor U11371 (N_11371,N_9394,N_9797);
or U11372 (N_11372,N_5506,N_5240);
or U11373 (N_11373,N_5264,N_6071);
or U11374 (N_11374,N_9465,N_6441);
and U11375 (N_11375,N_8724,N_5595);
or U11376 (N_11376,N_9615,N_7513);
nor U11377 (N_11377,N_9823,N_7727);
xnor U11378 (N_11378,N_8901,N_8408);
and U11379 (N_11379,N_7958,N_8883);
nand U11380 (N_11380,N_7051,N_5533);
nand U11381 (N_11381,N_6069,N_9403);
nand U11382 (N_11382,N_6712,N_7583);
nor U11383 (N_11383,N_5368,N_7884);
nand U11384 (N_11384,N_8115,N_6570);
or U11385 (N_11385,N_7440,N_6274);
nor U11386 (N_11386,N_6343,N_7350);
nand U11387 (N_11387,N_5088,N_8001);
nor U11388 (N_11388,N_7550,N_7603);
nand U11389 (N_11389,N_5437,N_6975);
xnor U11390 (N_11390,N_6944,N_7752);
and U11391 (N_11391,N_9610,N_9798);
nor U11392 (N_11392,N_7185,N_5237);
xnor U11393 (N_11393,N_5037,N_5070);
or U11394 (N_11394,N_8194,N_5535);
nor U11395 (N_11395,N_8304,N_7555);
nand U11396 (N_11396,N_8813,N_8646);
nand U11397 (N_11397,N_9621,N_9025);
xor U11398 (N_11398,N_5651,N_7763);
or U11399 (N_11399,N_8680,N_8447);
or U11400 (N_11400,N_8642,N_7220);
nor U11401 (N_11401,N_6040,N_9167);
or U11402 (N_11402,N_9494,N_8437);
nor U11403 (N_11403,N_8424,N_6436);
nand U11404 (N_11404,N_6215,N_5490);
and U11405 (N_11405,N_8325,N_9264);
nand U11406 (N_11406,N_8157,N_6856);
nand U11407 (N_11407,N_7296,N_8041);
and U11408 (N_11408,N_6762,N_6292);
nor U11409 (N_11409,N_7365,N_6166);
and U11410 (N_11410,N_5894,N_5728);
nand U11411 (N_11411,N_8973,N_9884);
nor U11412 (N_11412,N_8759,N_7041);
or U11413 (N_11413,N_6459,N_9399);
xor U11414 (N_11414,N_8087,N_7357);
xor U11415 (N_11415,N_7369,N_7940);
nand U11416 (N_11416,N_6079,N_5657);
or U11417 (N_11417,N_5947,N_9177);
nor U11418 (N_11418,N_6061,N_5062);
nand U11419 (N_11419,N_8884,N_7425);
nand U11420 (N_11420,N_8257,N_7245);
and U11421 (N_11421,N_9241,N_9087);
and U11422 (N_11422,N_5295,N_8965);
nor U11423 (N_11423,N_5707,N_9029);
or U11424 (N_11424,N_7631,N_9783);
or U11425 (N_11425,N_7316,N_8215);
xnor U11426 (N_11426,N_5834,N_7692);
nand U11427 (N_11427,N_7783,N_6067);
nand U11428 (N_11428,N_7042,N_7698);
xor U11429 (N_11429,N_9458,N_6240);
and U11430 (N_11430,N_8406,N_7181);
or U11431 (N_11431,N_7193,N_6315);
and U11432 (N_11432,N_9390,N_6496);
and U11433 (N_11433,N_6948,N_6342);
and U11434 (N_11434,N_7200,N_7834);
and U11435 (N_11435,N_5068,N_5854);
xnor U11436 (N_11436,N_5456,N_8107);
and U11437 (N_11437,N_5097,N_7419);
nor U11438 (N_11438,N_9420,N_5963);
nor U11439 (N_11439,N_8939,N_7501);
and U11440 (N_11440,N_8703,N_8781);
nor U11441 (N_11441,N_5909,N_9053);
nor U11442 (N_11442,N_7580,N_9667);
xnor U11443 (N_11443,N_9720,N_7401);
and U11444 (N_11444,N_6102,N_5061);
nor U11445 (N_11445,N_8431,N_6463);
xor U11446 (N_11446,N_9596,N_8063);
or U11447 (N_11447,N_5864,N_5024);
nand U11448 (N_11448,N_9684,N_9263);
or U11449 (N_11449,N_5475,N_5466);
and U11450 (N_11450,N_7113,N_8945);
nand U11451 (N_11451,N_6448,N_8893);
nand U11452 (N_11452,N_7103,N_7372);
and U11453 (N_11453,N_8033,N_8451);
xor U11454 (N_11454,N_6396,N_5308);
and U11455 (N_11455,N_8562,N_9731);
nor U11456 (N_11456,N_5771,N_6387);
and U11457 (N_11457,N_9968,N_5495);
or U11458 (N_11458,N_7820,N_9517);
or U11459 (N_11459,N_7248,N_9171);
nand U11460 (N_11460,N_9685,N_6789);
or U11461 (N_11461,N_8688,N_9371);
nor U11462 (N_11462,N_5469,N_9781);
nand U11463 (N_11463,N_6567,N_8697);
and U11464 (N_11464,N_5356,N_7263);
nand U11465 (N_11465,N_9719,N_6254);
or U11466 (N_11466,N_8778,N_9726);
and U11467 (N_11467,N_6029,N_6289);
nor U11468 (N_11468,N_5121,N_5397);
nand U11469 (N_11469,N_6249,N_9807);
nand U11470 (N_11470,N_6661,N_5165);
and U11471 (N_11471,N_9640,N_5010);
nor U11472 (N_11472,N_7754,N_6447);
xor U11473 (N_11473,N_8321,N_7259);
or U11474 (N_11474,N_7503,N_8261);
or U11475 (N_11475,N_8044,N_9878);
nand U11476 (N_11476,N_6755,N_6857);
nor U11477 (N_11477,N_9652,N_5372);
nand U11478 (N_11478,N_8821,N_5829);
xor U11479 (N_11479,N_5093,N_9041);
nor U11480 (N_11480,N_9074,N_8252);
nor U11481 (N_11481,N_9732,N_9305);
nand U11482 (N_11482,N_9570,N_5539);
xnor U11483 (N_11483,N_9997,N_9518);
nor U11484 (N_11484,N_7947,N_8399);
nor U11485 (N_11485,N_6851,N_8396);
nor U11486 (N_11486,N_6476,N_7877);
xor U11487 (N_11487,N_6301,N_9527);
and U11488 (N_11488,N_9630,N_8722);
xor U11489 (N_11489,N_7452,N_9206);
nor U11490 (N_11490,N_9646,N_6163);
nand U11491 (N_11491,N_9738,N_8416);
or U11492 (N_11492,N_6141,N_7618);
nor U11493 (N_11493,N_7178,N_6453);
nand U11494 (N_11494,N_9269,N_9733);
or U11495 (N_11495,N_6586,N_6009);
xnor U11496 (N_11496,N_5565,N_9721);
xnor U11497 (N_11497,N_7118,N_6773);
nand U11498 (N_11498,N_6910,N_6922);
xor U11499 (N_11499,N_6174,N_7836);
nand U11500 (N_11500,N_5210,N_6524);
or U11501 (N_11501,N_6498,N_6508);
xnor U11502 (N_11502,N_5325,N_6269);
nand U11503 (N_11503,N_8239,N_6581);
xor U11504 (N_11504,N_7716,N_6893);
or U11505 (N_11505,N_6302,N_9252);
xnor U11506 (N_11506,N_9196,N_8354);
xor U11507 (N_11507,N_8668,N_5757);
nand U11508 (N_11508,N_7657,N_9271);
nand U11509 (N_11509,N_7418,N_6370);
or U11510 (N_11510,N_5170,N_8380);
nor U11511 (N_11511,N_9748,N_8715);
or U11512 (N_11512,N_7647,N_6171);
and U11513 (N_11513,N_8398,N_9911);
nand U11514 (N_11514,N_6112,N_8822);
nor U11515 (N_11515,N_7907,N_6036);
or U11516 (N_11516,N_7099,N_6245);
or U11517 (N_11517,N_6329,N_5680);
or U11518 (N_11518,N_6638,N_9982);
nand U11519 (N_11519,N_8116,N_5255);
nor U11520 (N_11520,N_7959,N_8287);
nor U11521 (N_11521,N_5745,N_8256);
xor U11522 (N_11522,N_7847,N_5148);
or U11523 (N_11523,N_8708,N_5176);
and U11524 (N_11524,N_8989,N_7893);
xor U11525 (N_11525,N_6384,N_6831);
nor U11526 (N_11526,N_8204,N_5516);
xor U11527 (N_11527,N_9047,N_9855);
and U11528 (N_11528,N_7317,N_7644);
and U11529 (N_11529,N_7724,N_9562);
nor U11530 (N_11530,N_5239,N_8502);
nand U11531 (N_11531,N_5684,N_9377);
nand U11532 (N_11532,N_5897,N_7240);
and U11533 (N_11533,N_6158,N_9956);
xor U11534 (N_11534,N_5827,N_7760);
nor U11535 (N_11535,N_5014,N_8664);
nor U11536 (N_11536,N_8754,N_6743);
and U11537 (N_11537,N_9535,N_7596);
xor U11538 (N_11538,N_8500,N_5056);
or U11539 (N_11539,N_7448,N_8797);
xnor U11540 (N_11540,N_7089,N_8628);
xor U11541 (N_11541,N_5755,N_7814);
nand U11542 (N_11542,N_8209,N_8473);
nand U11543 (N_11543,N_6642,N_5182);
nand U11544 (N_11544,N_9578,N_6021);
nand U11545 (N_11545,N_5226,N_7214);
nand U11546 (N_11546,N_8533,N_6847);
or U11547 (N_11547,N_8103,N_8470);
nor U11548 (N_11548,N_9971,N_6964);
and U11549 (N_11549,N_7381,N_8142);
nor U11550 (N_11550,N_7439,N_7567);
nand U11551 (N_11551,N_6123,N_7211);
xnor U11552 (N_11552,N_8908,N_7218);
nand U11553 (N_11553,N_6552,N_7252);
nand U11554 (N_11554,N_9182,N_6170);
nand U11555 (N_11555,N_6326,N_9613);
nor U11556 (N_11556,N_5541,N_5699);
or U11557 (N_11557,N_6443,N_8267);
and U11558 (N_11558,N_9424,N_7444);
or U11559 (N_11559,N_5153,N_8071);
and U11560 (N_11560,N_6193,N_7324);
nand U11561 (N_11561,N_5282,N_6244);
and U11562 (N_11562,N_7822,N_9938);
xor U11563 (N_11563,N_5623,N_5693);
and U11564 (N_11564,N_7689,N_7901);
or U11565 (N_11565,N_8245,N_7354);
or U11566 (N_11566,N_7482,N_9441);
or U11567 (N_11567,N_7774,N_5335);
and U11568 (N_11568,N_5141,N_8136);
or U11569 (N_11569,N_6904,N_6105);
and U11570 (N_11570,N_8758,N_5481);
nor U11571 (N_11571,N_8400,N_9675);
xor U11572 (N_11572,N_5078,N_8185);
and U11573 (N_11573,N_7295,N_5080);
and U11574 (N_11574,N_6196,N_5118);
nor U11575 (N_11575,N_8594,N_8617);
xnor U11576 (N_11576,N_6549,N_6716);
nand U11577 (N_11577,N_5128,N_6988);
and U11578 (N_11578,N_9645,N_9953);
and U11579 (N_11579,N_9741,N_5208);
xnor U11580 (N_11580,N_7990,N_8545);
xnor U11581 (N_11581,N_7222,N_9123);
xor U11582 (N_11582,N_5230,N_9974);
nand U11583 (N_11583,N_9375,N_6350);
xor U11584 (N_11584,N_8332,N_8994);
xnor U11585 (N_11585,N_6867,N_9395);
and U11586 (N_11586,N_5805,N_8707);
or U11587 (N_11587,N_5468,N_6815);
and U11588 (N_11588,N_8745,N_5912);
nand U11589 (N_11589,N_6933,N_7097);
or U11590 (N_11590,N_6058,N_6168);
nand U11591 (N_11591,N_8040,N_6056);
or U11592 (N_11592,N_6231,N_8977);
or U11593 (N_11593,N_9491,N_5654);
and U11594 (N_11594,N_9585,N_5949);
nand U11595 (N_11595,N_6049,N_6295);
or U11596 (N_11596,N_9841,N_7085);
nand U11597 (N_11597,N_9183,N_8712);
nor U11598 (N_11598,N_6484,N_8331);
or U11599 (N_11599,N_6574,N_8439);
and U11600 (N_11600,N_9638,N_6417);
and U11601 (N_11601,N_7318,N_5171);
nand U11602 (N_11602,N_7929,N_6626);
or U11603 (N_11603,N_9918,N_5047);
nand U11604 (N_11604,N_8764,N_6967);
nor U11605 (N_11605,N_9591,N_6748);
or U11606 (N_11606,N_5958,N_5627);
nor U11607 (N_11607,N_6852,N_7619);
xnor U11608 (N_11608,N_7701,N_7728);
xor U11609 (N_11609,N_6495,N_7713);
xnor U11610 (N_11610,N_5982,N_9772);
nand U11611 (N_11611,N_8935,N_9951);
nand U11612 (N_11612,N_6695,N_7723);
and U11613 (N_11613,N_9215,N_8405);
nor U11614 (N_11614,N_6869,N_5199);
xnor U11615 (N_11615,N_9257,N_7190);
or U11616 (N_11616,N_7527,N_6294);
xnor U11617 (N_11617,N_8492,N_9174);
or U11618 (N_11618,N_5459,N_9542);
xor U11619 (N_11619,N_8152,N_5346);
or U11620 (N_11620,N_8133,N_5758);
nand U11621 (N_11621,N_7484,N_9172);
and U11622 (N_11622,N_5998,N_8875);
nand U11623 (N_11623,N_7515,N_9384);
nor U11624 (N_11624,N_6924,N_6070);
xnor U11625 (N_11625,N_9423,N_6025);
and U11626 (N_11626,N_7284,N_8985);
xor U11627 (N_11627,N_5246,N_7009);
xor U11628 (N_11628,N_5650,N_5921);
nor U11629 (N_11629,N_6085,N_8516);
or U11630 (N_11630,N_5991,N_7314);
nor U11631 (N_11631,N_5848,N_8934);
xor U11632 (N_11632,N_6624,N_9189);
nand U11633 (N_11633,N_9078,N_6613);
and U11634 (N_11634,N_8850,N_5443);
nor U11635 (N_11635,N_9538,N_6284);
and U11636 (N_11636,N_6753,N_9212);
nor U11637 (N_11637,N_5807,N_6579);
or U11638 (N_11638,N_5320,N_9752);
nor U11639 (N_11639,N_6402,N_5524);
and U11640 (N_11640,N_9411,N_8254);
nor U11641 (N_11641,N_7787,N_7147);
xnor U11642 (N_11642,N_7034,N_9058);
or U11643 (N_11643,N_7876,N_8164);
and U11644 (N_11644,N_7443,N_6781);
nand U11645 (N_11645,N_5957,N_8765);
nand U11646 (N_11646,N_7951,N_5371);
or U11647 (N_11647,N_5439,N_8789);
or U11648 (N_11648,N_8782,N_5315);
nand U11649 (N_11649,N_7275,N_8921);
nand U11650 (N_11650,N_5702,N_8980);
xor U11651 (N_11651,N_8017,N_6572);
nand U11652 (N_11652,N_8253,N_5407);
or U11653 (N_11653,N_6287,N_9280);
xnor U11654 (N_11654,N_8863,N_8316);
xor U11655 (N_11655,N_9782,N_7371);
and U11656 (N_11656,N_5578,N_5098);
xnor U11657 (N_11657,N_6031,N_7581);
nor U11658 (N_11658,N_6859,N_9219);
nand U11659 (N_11659,N_9623,N_6502);
or U11660 (N_11660,N_7446,N_9688);
nor U11661 (N_11661,N_7094,N_6205);
and U11662 (N_11662,N_8636,N_8369);
xor U11663 (N_11663,N_9113,N_9766);
nor U11664 (N_11664,N_7879,N_8830);
and U11665 (N_11665,N_5483,N_7242);
nor U11666 (N_11666,N_5025,N_8602);
nor U11667 (N_11667,N_8366,N_7718);
and U11668 (N_11668,N_7722,N_7258);
nor U11669 (N_11669,N_8488,N_6115);
and U11670 (N_11670,N_7155,N_5279);
nor U11671 (N_11671,N_7536,N_8334);
xor U11672 (N_11672,N_7886,N_9095);
xnor U11673 (N_11673,N_5614,N_5030);
and U11674 (N_11674,N_8066,N_9119);
nand U11675 (N_11675,N_7506,N_8211);
nor U11676 (N_11676,N_9751,N_6323);
nor U11677 (N_11677,N_6983,N_7936);
and U11678 (N_11678,N_9003,N_9980);
nand U11679 (N_11679,N_9887,N_9515);
xor U11680 (N_11680,N_8857,N_6177);
xnor U11681 (N_11681,N_5448,N_7329);
nor U11682 (N_11682,N_9857,N_7806);
and U11683 (N_11683,N_5590,N_8275);
xnor U11684 (N_11684,N_7319,N_7122);
and U11685 (N_11685,N_5956,N_8557);
nor U11686 (N_11686,N_6162,N_7031);
or U11687 (N_11687,N_9261,N_6504);
or U11688 (N_11688,N_9217,N_6452);
nand U11689 (N_11689,N_8871,N_5227);
nor U11690 (N_11690,N_5122,N_8735);
nor U11691 (N_11691,N_7247,N_6951);
or U11692 (N_11692,N_9000,N_8932);
or U11693 (N_11693,N_9247,N_7213);
nor U11694 (N_11694,N_7597,N_9385);
or U11695 (N_11695,N_6408,N_8309);
xnor U11696 (N_11696,N_7270,N_5580);
or U11697 (N_11697,N_5833,N_9994);
or U11698 (N_11698,N_8593,N_6057);
xnor U11699 (N_11699,N_5586,N_5948);
and U11700 (N_11700,N_5427,N_9948);
and U11701 (N_11701,N_8073,N_9042);
or U11702 (N_11702,N_7057,N_6946);
nor U11703 (N_11703,N_9795,N_7340);
and U11704 (N_11704,N_6568,N_7476);
or U11705 (N_11705,N_5040,N_6842);
nor U11706 (N_11706,N_9150,N_7726);
nor U11707 (N_11707,N_9794,N_9722);
or U11708 (N_11708,N_7707,N_9530);
nand U11709 (N_11709,N_5033,N_9683);
nor U11710 (N_11710,N_9295,N_9199);
and U11711 (N_11711,N_6107,N_5422);
nor U11712 (N_11712,N_5180,N_9309);
nor U11713 (N_11713,N_5639,N_7056);
xnor U11714 (N_11714,N_7945,N_9724);
xor U11715 (N_11715,N_6407,N_7646);
and U11716 (N_11716,N_7269,N_7560);
nand U11717 (N_11717,N_5002,N_9175);
xor U11718 (N_11718,N_5775,N_5852);
nand U11719 (N_11719,N_8559,N_7888);
or U11720 (N_11720,N_6744,N_9145);
and U11721 (N_11721,N_8687,N_5933);
and U11722 (N_11722,N_6649,N_5670);
xor U11723 (N_11723,N_6340,N_6351);
or U11724 (N_11724,N_6426,N_8303);
and U11725 (N_11725,N_7656,N_9995);
xnor U11726 (N_11726,N_5410,N_8464);
and U11727 (N_11727,N_9649,N_5342);
and U11728 (N_11728,N_6627,N_7952);
and U11729 (N_11729,N_6139,N_9232);
xnor U11730 (N_11730,N_9905,N_5772);
xor U11731 (N_11731,N_8580,N_8825);
nor U11732 (N_11732,N_6197,N_7751);
xnor U11733 (N_11733,N_5720,N_5902);
xnor U11734 (N_11734,N_8493,N_7239);
and U11735 (N_11735,N_6369,N_8755);
xnor U11736 (N_11736,N_5638,N_5444);
nor U11737 (N_11737,N_5525,N_8306);
nand U11738 (N_11738,N_5936,N_9819);
xnor U11739 (N_11739,N_5782,N_8378);
and U11740 (N_11740,N_8560,N_8165);
nand U11741 (N_11741,N_9006,N_9153);
nand U11742 (N_11742,N_5464,N_9056);
and U11743 (N_11743,N_9382,N_8746);
or U11744 (N_11744,N_9158,N_5945);
nand U11745 (N_11745,N_7460,N_6190);
and U11746 (N_11746,N_7909,N_8885);
and U11747 (N_11747,N_7861,N_5345);
or U11748 (N_11748,N_7685,N_9236);
nor U11749 (N_11749,N_5940,N_9302);
nor U11750 (N_11750,N_5628,N_6022);
nor U11751 (N_11751,N_8635,N_9792);
and U11752 (N_11752,N_7281,N_8244);
xor U11753 (N_11753,N_5140,N_9392);
nor U11754 (N_11754,N_6401,N_6423);
or U11755 (N_11755,N_9552,N_7858);
xnor U11756 (N_11756,N_9406,N_6503);
or U11757 (N_11757,N_7852,N_5291);
nand U11758 (N_11758,N_8640,N_7101);
nor U11759 (N_11759,N_5251,N_8891);
xor U11760 (N_11760,N_9200,N_9091);
or U11761 (N_11761,N_6341,N_8184);
nor U11762 (N_11762,N_8552,N_9693);
nor U11763 (N_11763,N_5559,N_7146);
and U11764 (N_11764,N_5551,N_9826);
nor U11765 (N_11765,N_7939,N_7331);
or U11766 (N_11766,N_6481,N_8975);
or U11767 (N_11767,N_6602,N_5503);
or U11768 (N_11768,N_6091,N_7522);
and U11769 (N_11769,N_8301,N_9018);
nand U11770 (N_11770,N_7492,N_6745);
and U11771 (N_11771,N_5492,N_8339);
or U11772 (N_11772,N_6777,N_5117);
and U11773 (N_11773,N_9500,N_8532);
and U11774 (N_11774,N_8237,N_7426);
and U11775 (N_11775,N_5917,N_5634);
xnor U11776 (N_11776,N_7496,N_7584);
or U11777 (N_11777,N_9920,N_8659);
xor U11778 (N_11778,N_5803,N_6709);
or U11779 (N_11779,N_7438,N_9218);
and U11780 (N_11780,N_9068,N_7432);
nor U11781 (N_11781,N_7731,N_9268);
nor U11782 (N_11782,N_7138,N_5746);
nor U11783 (N_11783,N_5831,N_6438);
xnor U11784 (N_11784,N_7229,N_7518);
and U11785 (N_11785,N_8632,N_6120);
xor U11786 (N_11786,N_9425,N_8432);
nor U11787 (N_11787,N_7054,N_6954);
xor U11788 (N_11788,N_8217,N_6210);
or U11789 (N_11789,N_9256,N_5383);
or U11790 (N_11790,N_6361,N_5893);
nand U11791 (N_11791,N_8238,N_6717);
or U11792 (N_11792,N_5592,N_5249);
nand U11793 (N_11793,N_5583,N_9658);
nand U11794 (N_11794,N_9451,N_5659);
or U11795 (N_11795,N_9612,N_5017);
xnor U11796 (N_11796,N_6832,N_8368);
nand U11797 (N_11797,N_6053,N_8595);
or U11798 (N_11798,N_7069,N_8870);
xor U11799 (N_11799,N_9085,N_5557);
and U11800 (N_11800,N_9325,N_5378);
xor U11801 (N_11801,N_9456,N_5607);
and U11802 (N_11802,N_6760,N_8684);
nor U11803 (N_11803,N_6399,N_7060);
and U11804 (N_11804,N_8546,N_6597);
or U11805 (N_11805,N_5576,N_7403);
nor U11806 (N_11806,N_8128,N_5452);
or U11807 (N_11807,N_5144,N_7111);
xor U11808 (N_11808,N_5631,N_7182);
or U11809 (N_11809,N_5358,N_8269);
xnor U11810 (N_11810,N_9186,N_8838);
and U11811 (N_11811,N_7450,N_5332);
xor U11812 (N_11812,N_9581,N_9224);
xnor U11813 (N_11813,N_8233,N_5712);
nand U11814 (N_11814,N_5177,N_7809);
and U11815 (N_11815,N_7420,N_7254);
and U11816 (N_11816,N_5853,N_7610);
and U11817 (N_11817,N_5135,N_8498);
and U11818 (N_11818,N_7080,N_8433);
or U11819 (N_11819,N_9437,N_5275);
xor U11820 (N_11820,N_6525,N_8706);
nor U11821 (N_11821,N_8035,N_7797);
and U11822 (N_11822,N_8158,N_5431);
nor U11823 (N_11823,N_6875,N_6109);
or U11824 (N_11824,N_6915,N_9292);
xnor U11825 (N_11825,N_8794,N_6541);
and U11826 (N_11826,N_7157,N_7571);
nand U11827 (N_11827,N_7429,N_6802);
nor U11828 (N_11828,N_5653,N_5741);
or U11829 (N_11829,N_6526,N_5542);
nor U11830 (N_11830,N_5152,N_7512);
nor U11831 (N_11831,N_8845,N_7162);
and U11832 (N_11832,N_7002,N_6238);
xor U11833 (N_11833,N_9084,N_8561);
and U11834 (N_11834,N_6900,N_5508);
nand U11835 (N_11835,N_7765,N_8996);
and U11836 (N_11836,N_9506,N_7187);
and U11837 (N_11837,N_5178,N_5312);
nor U11838 (N_11838,N_5714,N_8458);
xor U11839 (N_11839,N_5169,N_8565);
or U11840 (N_11840,N_5647,N_8523);
nand U11841 (N_11841,N_6288,N_7093);
or U11842 (N_11842,N_5978,N_9080);
xnor U11843 (N_11843,N_8672,N_5629);
and U11844 (N_11844,N_7588,N_7863);
nor U11845 (N_11845,N_8823,N_6611);
and U11846 (N_11846,N_9665,N_6466);
nor U11847 (N_11847,N_7333,N_5158);
and U11848 (N_11848,N_7410,N_6137);
nor U11849 (N_11849,N_8282,N_9166);
nand U11850 (N_11850,N_5858,N_6297);
xnor U11851 (N_11851,N_5752,N_6522);
nor U11852 (N_11852,N_9662,N_9227);
and U11853 (N_11853,N_9545,N_8853);
or U11854 (N_11854,N_5646,N_9031);
nand U11855 (N_11855,N_6772,N_8248);
or U11856 (N_11856,N_7630,N_9694);
and U11857 (N_11857,N_5872,N_9793);
xor U11858 (N_11858,N_8490,N_6659);
nor U11859 (N_11859,N_5369,N_8937);
xor U11860 (N_11860,N_6146,N_9402);
nand U11861 (N_11861,N_5553,N_6366);
and U11862 (N_11862,N_8249,N_8536);
and U11863 (N_11863,N_9428,N_7231);
nor U11864 (N_11864,N_9668,N_8166);
nor U11865 (N_11865,N_7077,N_9539);
nand U11866 (N_11866,N_7720,N_5028);
and U11867 (N_11867,N_7841,N_5605);
nand U11868 (N_11868,N_6223,N_6044);
nand U11869 (N_11869,N_7942,N_5084);
or U11870 (N_11870,N_6742,N_6362);
or U11871 (N_11871,N_5500,N_7738);
or U11872 (N_11872,N_5905,N_7207);
and U11873 (N_11873,N_6026,N_9474);
nand U11874 (N_11874,N_9984,N_9059);
nand U11875 (N_11875,N_8915,N_5129);
xor U11876 (N_11876,N_7130,N_6996);
and U11877 (N_11877,N_5133,N_5616);
and U11878 (N_11878,N_5883,N_5641);
nand U11879 (N_11879,N_9873,N_6747);
nand U11880 (N_11880,N_6718,N_8542);
and U11881 (N_11881,N_9471,N_7389);
xor U11882 (N_11882,N_5835,N_5798);
and U11883 (N_11883,N_9483,N_6047);
nor U11884 (N_11884,N_6202,N_8844);
nor U11885 (N_11885,N_8669,N_8356);
and U11886 (N_11886,N_9226,N_6992);
nand U11887 (N_11887,N_6682,N_5394);
xor U11888 (N_11888,N_5779,N_8817);
and U11889 (N_11889,N_6722,N_7771);
or U11890 (N_11890,N_8465,N_7236);
nand U11891 (N_11891,N_8351,N_6707);
or U11892 (N_11892,N_6075,N_6064);
xnor U11893 (N_11893,N_5286,N_7458);
xor U11894 (N_11894,N_8571,N_8434);
nand U11895 (N_11895,N_9611,N_7628);
xnor U11896 (N_11896,N_7992,N_7544);
nor U11897 (N_11897,N_9077,N_5223);
or U11898 (N_11898,N_8657,N_9487);
nand U11899 (N_11899,N_6966,N_6540);
xor U11900 (N_11900,N_9353,N_9454);
xor U11901 (N_11901,N_6654,N_6243);
xor U11902 (N_11902,N_8240,N_8624);
nand U11903 (N_11903,N_6357,N_5577);
and U11904 (N_11904,N_9159,N_8618);
and U11905 (N_11905,N_6879,N_6430);
nand U11906 (N_11906,N_7824,N_8345);
nor U11907 (N_11907,N_8846,N_8730);
nor U11908 (N_11908,N_6880,N_8783);
xnor U11909 (N_11909,N_9315,N_5031);
nand U11910 (N_11910,N_7192,N_9574);
nand U11911 (N_11911,N_5843,N_9569);
or U11912 (N_11912,N_5700,N_6768);
nor U11913 (N_11913,N_9381,N_5103);
xor U11914 (N_11914,N_7435,N_7677);
and U11915 (N_11915,N_6749,N_5482);
nand U11916 (N_11916,N_8441,N_7126);
nor U11917 (N_11917,N_9565,N_8584);
xnor U11918 (N_11918,N_9893,N_5340);
and U11919 (N_11919,N_5698,N_5027);
xnor U11920 (N_11920,N_7021,N_7840);
xnor U11921 (N_11921,N_9899,N_5561);
or U11922 (N_11922,N_6633,N_5019);
xnor U11923 (N_11923,N_5774,N_5041);
nor U11924 (N_11924,N_7362,N_9602);
xor U11925 (N_11925,N_6471,N_8358);
or U11926 (N_11926,N_5575,N_8681);
and U11927 (N_11927,N_6267,N_5493);
and U11928 (N_11928,N_7762,N_7044);
nor U11929 (N_11929,N_6825,N_7890);
or U11930 (N_11930,N_6194,N_8760);
xor U11931 (N_11931,N_9076,N_7734);
nand U11932 (N_11932,N_8527,N_5687);
xnor U11933 (N_11933,N_9834,N_6982);
xor U11934 (N_11934,N_9055,N_9361);
or U11935 (N_11935,N_5839,N_5167);
xnor U11936 (N_11936,N_9544,N_8836);
or U11937 (N_11937,N_8936,N_9833);
xnor U11938 (N_11938,N_6767,N_8675);
xnor U11939 (N_11939,N_7997,N_9967);
and U11940 (N_11940,N_7462,N_6993);
or U11941 (N_11941,N_5632,N_6671);
xor U11942 (N_11942,N_6138,N_6518);
nand U11943 (N_11943,N_9314,N_6548);
or U11944 (N_11944,N_7453,N_7837);
xor U11945 (N_11945,N_8075,N_7407);
xnor U11946 (N_11946,N_5204,N_7116);
or U11947 (N_11947,N_6678,N_9876);
nor U11948 (N_11948,N_5619,N_6454);
or U11949 (N_11949,N_5137,N_7480);
nand U11950 (N_11950,N_9415,N_7010);
and U11951 (N_11951,N_8700,N_5910);
xnor U11952 (N_11952,N_9851,N_6909);
and U11953 (N_11953,N_5907,N_9157);
nor U11954 (N_11954,N_6577,N_5979);
or U11955 (N_11955,N_9680,N_9329);
nor U11956 (N_11956,N_9825,N_9160);
xnor U11957 (N_11957,N_9481,N_6152);
nor U11958 (N_11958,N_7224,N_9521);
xor U11959 (N_11959,N_7680,N_7234);
and U11960 (N_11960,N_5261,N_5821);
nand U11961 (N_11961,N_7062,N_8064);
and U11962 (N_11962,N_9513,N_5412);
and U11963 (N_11963,N_7115,N_6778);
and U11964 (N_11964,N_8579,N_9286);
nor U11965 (N_11965,N_9842,N_5460);
xor U11966 (N_11966,N_7653,N_6963);
and U11967 (N_11967,N_7090,N_6449);
nor U11968 (N_11968,N_6593,N_5785);
and U11969 (N_11969,N_9468,N_8418);
and U11970 (N_11970,N_9345,N_9277);
xor U11971 (N_11971,N_9079,N_7301);
nand U11972 (N_11972,N_5487,N_6945);
nor U11973 (N_11973,N_7866,N_5406);
xnor U11974 (N_11974,N_9973,N_6439);
xnor U11975 (N_11975,N_7199,N_8787);
or U11976 (N_11976,N_9629,N_9969);
nor U11977 (N_11977,N_7998,N_7167);
nor U11978 (N_11978,N_9970,N_7076);
nand U11979 (N_11979,N_5403,N_8526);
xnor U11980 (N_11980,N_7406,N_9558);
and U11981 (N_11981,N_7033,N_5337);
xor U11982 (N_11982,N_5289,N_9479);
xor U11983 (N_11983,N_5941,N_9466);
or U11984 (N_11984,N_7743,N_7739);
xor U11985 (N_11985,N_5656,N_9062);
nand U11986 (N_11986,N_8826,N_5220);
or U11987 (N_11987,N_7382,N_6431);
and U11988 (N_11988,N_9699,N_8455);
or U11989 (N_11989,N_5401,N_5164);
xnor U11990 (N_11990,N_7353,N_6207);
nand U11991 (N_11991,N_8143,N_8506);
or U11992 (N_11992,N_5857,N_8178);
xnor U11993 (N_11993,N_5361,N_9923);
and U11994 (N_11994,N_9446,N_7770);
xnor U11995 (N_11995,N_6030,N_6738);
nor U11996 (N_11996,N_8525,N_7461);
or U11997 (N_11997,N_6837,N_7398);
and U11998 (N_11998,N_6424,N_9388);
and U11999 (N_11999,N_7703,N_7570);
nand U12000 (N_12000,N_8530,N_6554);
nor U12001 (N_12001,N_7520,N_9975);
nor U12002 (N_12002,N_6741,N_5674);
nor U12003 (N_12003,N_8411,N_9155);
nand U12004 (N_12004,N_5209,N_8039);
and U12005 (N_12005,N_5381,N_5077);
xor U12006 (N_12006,N_7910,N_5919);
and U12007 (N_12007,N_6592,N_9546);
nand U12008 (N_12008,N_5855,N_6916);
or U12009 (N_12009,N_9850,N_6305);
or U12010 (N_12010,N_7347,N_6485);
nor U12011 (N_12011,N_5691,N_8413);
and U12012 (N_12012,N_9478,N_8336);
or U12013 (N_12013,N_5960,N_5884);
and U12014 (N_12014,N_5479,N_9698);
or U12015 (N_12015,N_8747,N_6595);
and U12016 (N_12016,N_9925,N_5589);
xor U12017 (N_12017,N_8069,N_6203);
nand U12018 (N_12018,N_5534,N_8089);
xor U12019 (N_12019,N_5113,N_8027);
nor U12020 (N_12020,N_9786,N_6081);
and U12021 (N_12021,N_5408,N_7523);
nor U12022 (N_12022,N_8250,N_5348);
or U12023 (N_12023,N_9170,N_9143);
and U12024 (N_12024,N_6457,N_6339);
or U12025 (N_12025,N_8690,N_8651);
nand U12026 (N_12026,N_8452,N_6189);
or U12027 (N_12027,N_6211,N_8698);
and U12028 (N_12028,N_9735,N_6531);
or U12029 (N_12029,N_5259,N_7133);
xnor U12030 (N_12030,N_8739,N_9107);
nand U12031 (N_12031,N_7380,N_8169);
or U12032 (N_12032,N_9837,N_8596);
xor U12033 (N_12033,N_7064,N_5697);
xnor U12034 (N_12034,N_5096,N_5976);
nor U12035 (N_12035,N_9579,N_5946);
nand U12036 (N_12036,N_7593,N_6766);
nor U12037 (N_12037,N_6225,N_9763);
nor U12038 (N_12038,N_5225,N_8385);
or U12039 (N_12039,N_5649,N_5008);
or U12040 (N_12040,N_8567,N_8716);
and U12041 (N_12041,N_5523,N_9202);
or U12042 (N_12042,N_8262,N_7747);
nand U12043 (N_12043,N_9924,N_9686);
xor U12044 (N_12044,N_9745,N_9048);
and U12045 (N_12045,N_5498,N_9547);
nand U12046 (N_12046,N_6656,N_5305);
nor U12047 (N_12047,N_6833,N_8589);
nor U12048 (N_12048,N_9434,N_5924);
and U12049 (N_12049,N_6961,N_9283);
xor U12050 (N_12050,N_8162,N_9691);
or U12051 (N_12051,N_9242,N_9173);
nand U12052 (N_12052,N_5892,N_6868);
and U12053 (N_12053,N_8145,N_5216);
and U12054 (N_12054,N_6733,N_9791);
nor U12055 (N_12055,N_7052,N_7924);
xnor U12056 (N_12056,N_8251,N_5694);
and U12057 (N_12057,N_7053,N_6096);
and U12058 (N_12058,N_8918,N_9480);
or U12059 (N_12059,N_6164,N_8859);
xor U12060 (N_12060,N_7075,N_5287);
xnor U12061 (N_12061,N_8947,N_6918);
nand U12062 (N_12062,N_5491,N_5911);
or U12063 (N_12063,N_8809,N_8440);
and U12064 (N_12064,N_7188,N_9288);
nor U12065 (N_12065,N_5145,N_9023);
or U12066 (N_12066,N_9808,N_8550);
and U12067 (N_12067,N_8517,N_5890);
or U12068 (N_12068,N_9853,N_6169);
xnor U12069 (N_12069,N_7759,N_5560);
xor U12070 (N_12070,N_6547,N_9319);
nor U12071 (N_12071,N_7481,N_8401);
nand U12072 (N_12072,N_7799,N_7423);
xnor U12073 (N_12073,N_7083,N_5880);
nor U12074 (N_12074,N_8837,N_7325);
nand U12075 (N_12075,N_6464,N_9768);
nand U12076 (N_12076,N_5923,N_6564);
xnor U12077 (N_12077,N_9106,N_9020);
xor U12078 (N_12078,N_8768,N_6237);
nand U12079 (N_12079,N_6316,N_5882);
and U12080 (N_12080,N_6003,N_8373);
nor U12081 (N_12081,N_8606,N_8323);
nor U12082 (N_12082,N_7629,N_6127);
nor U12083 (N_12083,N_8002,N_6377);
xor U12084 (N_12084,N_8897,N_6232);
nor U12085 (N_12085,N_9780,N_8913);
xor U12086 (N_12086,N_7504,N_7261);
or U12087 (N_12087,N_5205,N_7733);
nor U12088 (N_12088,N_8307,N_8641);
nor U12089 (N_12089,N_9496,N_8946);
nand U12090 (N_12090,N_6268,N_8997);
nor U12091 (N_12091,N_8140,N_9136);
nor U12092 (N_12092,N_7725,N_7376);
xnor U12093 (N_12093,N_7368,N_8272);
and U12094 (N_12094,N_7796,N_5336);
xnor U12095 (N_12095,N_9443,N_6710);
nor U12096 (N_12096,N_8849,N_9461);
and U12097 (N_12097,N_5787,N_7744);
or U12098 (N_12098,N_5875,N_8070);
nor U12099 (N_12099,N_5124,N_9847);
nand U12100 (N_12100,N_7000,N_8954);
or U12101 (N_12101,N_8873,N_5937);
nor U12102 (N_12102,N_5901,N_7243);
and U12103 (N_12103,N_8175,N_5421);
nand U12104 (N_12104,N_7449,N_6544);
nand U12105 (N_12105,N_6674,N_6791);
and U12106 (N_12106,N_8394,N_5736);
or U12107 (N_12107,N_6046,N_7280);
or U12108 (N_12108,N_7428,N_5517);
nand U12109 (N_12109,N_7928,N_5532);
or U12110 (N_12110,N_8060,N_6786);
xor U12111 (N_12111,N_7980,N_9894);
and U12112 (N_12112,N_9714,N_9204);
xnor U12113 (N_12113,N_5453,N_5615);
or U12114 (N_12114,N_7215,N_5744);
or U12115 (N_12115,N_7238,N_6450);
xor U12116 (N_12116,N_7903,N_9045);
nand U12117 (N_12117,N_7591,N_6991);
and U12118 (N_12118,N_8867,N_9907);
and U12119 (N_12119,N_6952,N_7393);
xor U12120 (N_12120,N_9324,N_6545);
or U12121 (N_12121,N_7383,N_6078);
and U12122 (N_12122,N_8733,N_9609);
nand U12123 (N_12123,N_6183,N_6304);
or U12124 (N_12124,N_8895,N_7524);
nand U12125 (N_12125,N_5652,N_6657);
xor U12126 (N_12126,N_5293,N_9057);
nand U12127 (N_12127,N_9644,N_5271);
or U12128 (N_12128,N_5114,N_7988);
xor U12129 (N_12129,N_6631,N_9523);
nand U12130 (N_12130,N_5391,N_8067);
nand U12131 (N_12131,N_6662,N_6874);
nand U12132 (N_12132,N_7001,N_7546);
and U12133 (N_12133,N_5900,N_6623);
xnor U12134 (N_12134,N_8450,N_9285);
and U12135 (N_12135,N_6583,N_7838);
nor U12136 (N_12136,N_8663,N_7978);
nand U12137 (N_12137,N_6363,N_9634);
or U12138 (N_12138,N_9827,N_9743);
or U12139 (N_12139,N_9608,N_6150);
nand U12140 (N_12140,N_5173,N_5472);
nor U12141 (N_12141,N_7364,N_5174);
xnor U12142 (N_12142,N_8599,N_8390);
nand U12143 (N_12143,N_8161,N_9433);
nor U12144 (N_12144,N_8311,N_8047);
xnor U12145 (N_12145,N_8494,N_9099);
and U12146 (N_12146,N_5366,N_8268);
xor U12147 (N_12147,N_8384,N_5186);
nand U12148 (N_12148,N_5018,N_5837);
and U12149 (N_12149,N_6714,N_6059);
and U12150 (N_12150,N_9790,N_7683);
xnor U12151 (N_12151,N_5970,N_5569);
and U12152 (N_12152,N_9497,N_6376);
xor U12153 (N_12153,N_6644,N_8969);
and U12154 (N_12154,N_5217,N_6905);
nand U12155 (N_12155,N_6866,N_7519);
nor U12156 (N_12156,N_6277,N_6972);
xor U12157 (N_12157,N_8083,N_5846);
xor U12158 (N_12158,N_6647,N_6936);
and U12159 (N_12159,N_6509,N_7808);
or U12160 (N_12160,N_8992,N_9522);
or U12161 (N_12161,N_8621,N_8967);
nand U12162 (N_12162,N_8791,N_5006);
or U12163 (N_12163,N_8205,N_5091);
nand U12164 (N_12164,N_6181,N_5725);
nand U12165 (N_12165,N_5333,N_9308);
xor U12166 (N_12166,N_8355,N_5415);
and U12167 (N_12167,N_5721,N_6242);
nand U12168 (N_12168,N_9278,N_5190);
or U12169 (N_12169,N_7395,N_7773);
nand U12170 (N_12170,N_6546,N_7385);
or U12171 (N_12171,N_5049,N_7682);
or U12172 (N_12172,N_6990,N_9284);
nand U12173 (N_12173,N_9444,N_6251);
and U12174 (N_12174,N_5280,N_8990);
xor U12175 (N_12175,N_6637,N_6082);
or U12176 (N_12176,N_5954,N_5076);
nor U12177 (N_12177,N_7386,N_5044);
nand U12178 (N_12178,N_9452,N_6159);
nand U12179 (N_12179,N_8374,N_9550);
xor U12180 (N_12180,N_6224,N_6775);
or U12181 (N_12181,N_8486,N_9828);
and U12182 (N_12182,N_9223,N_7828);
nor U12183 (N_12183,N_6957,N_5734);
nand U12184 (N_12184,N_9809,N_6645);
and U12185 (N_12185,N_9945,N_9531);
nor U12186 (N_12186,N_9868,N_6353);
nor U12187 (N_12187,N_5416,N_9869);
xnor U12188 (N_12188,N_9007,N_7598);
nor U12189 (N_12189,N_8622,N_7652);
or U12190 (N_12190,N_7189,N_7039);
or U12191 (N_12191,N_6721,N_5243);
nor U12192 (N_12192,N_5931,N_5920);
or U12193 (N_12193,N_8042,N_9541);
and U12194 (N_12194,N_6494,N_6876);
and U12195 (N_12195,N_6084,N_9799);
and U12196 (N_12196,N_8112,N_6324);
nor U12197 (N_12197,N_7695,N_5751);
nor U12198 (N_12198,N_8974,N_5075);
xnor U12199 (N_12199,N_5036,N_5032);
and U12200 (N_12200,N_8577,N_9244);
nand U12201 (N_12201,N_7635,N_8477);
xor U12202 (N_12202,N_5742,N_7753);
nor U12203 (N_12203,N_8446,N_6032);
nand U12204 (N_12204,N_8481,N_9352);
or U12205 (N_12205,N_7253,N_5016);
nor U12206 (N_12206,N_9604,N_6756);
nor U12207 (N_12207,N_8188,N_5087);
and U12208 (N_12208,N_6331,N_7920);
and U12209 (N_12209,N_6279,N_9102);
nor U12210 (N_12210,N_8294,N_7205);
or U12211 (N_12211,N_8310,N_9251);
or U12212 (N_12212,N_8592,N_8769);
or U12213 (N_12213,N_6790,N_6843);
or U12214 (N_12214,N_8930,N_5058);
or U12215 (N_12215,N_7065,N_9590);
nor U12216 (N_12216,N_9163,N_7388);
nor U12217 (N_12217,N_8226,N_8412);
or U12218 (N_12218,N_5485,N_7905);
or U12219 (N_12219,N_7139,N_7803);
and U12220 (N_12220,N_8998,N_8255);
nor U12221 (N_12221,N_5690,N_9378);
or U12222 (N_12222,N_7804,N_5719);
and U12223 (N_12223,N_5544,N_8948);
or U12224 (N_12224,N_6841,N_9671);
and U12225 (N_12225,N_9369,N_5343);
xnor U12226 (N_12226,N_8173,N_6469);
nand U12227 (N_12227,N_7495,N_8609);
nand U12228 (N_12228,N_9299,N_8333);
xor U12229 (N_12229,N_7968,N_7578);
nand U12230 (N_12230,N_6523,N_5566);
nand U12231 (N_12231,N_9347,N_6161);
nor U12232 (N_12232,N_7370,N_7825);
nand U12233 (N_12233,N_7872,N_9789);
nand U12234 (N_12234,N_8900,N_9814);
or U12235 (N_12235,N_6257,N_8582);
or U12236 (N_12236,N_7777,N_7565);
xnor U12237 (N_12237,N_8362,N_5235);
or U12238 (N_12238,N_5993,N_9778);
nand U12239 (N_12239,N_9362,N_6418);
xor U12240 (N_12240,N_9785,N_5514);
and U12241 (N_12241,N_9554,N_5375);
or U12242 (N_12242,N_7257,N_8459);
nor U12243 (N_12243,N_9770,N_7632);
nand U12244 (N_12244,N_9213,N_8993);
xor U12245 (N_12245,N_7873,N_6603);
and U12246 (N_12246,N_6312,N_8149);
and U12247 (N_12247,N_8221,N_8104);
xor U12248 (N_12248,N_6052,N_7241);
and U12249 (N_12249,N_8587,N_7805);
xnor U12250 (N_12250,N_8956,N_8231);
or U12251 (N_12251,N_6461,N_8499);
or U12252 (N_12252,N_8367,N_8522);
nand U12253 (N_12253,N_7283,N_5896);
xor U12254 (N_12254,N_8371,N_6344);
and U12255 (N_12255,N_9796,N_5085);
nand U12256 (N_12256,N_6782,N_6272);
or U12257 (N_12257,N_8929,N_8647);
and U12258 (N_12258,N_8793,N_8084);
xnor U12259 (N_12259,N_5845,N_9440);
or U12260 (N_12260,N_6553,N_9943);
or U12261 (N_12261,N_8110,N_6273);
and U12262 (N_12262,N_9233,N_6517);
or U12263 (N_12263,N_6658,N_7285);
nor U12264 (N_12264,N_6014,N_7994);
xor U12265 (N_12265,N_8293,N_9335);
or U12266 (N_12266,N_6932,N_5847);
nor U12267 (N_12267,N_5562,N_9192);
and U12268 (N_12268,N_7634,N_9467);
xor U12269 (N_12269,N_7923,N_8330);
xor U12270 (N_12270,N_8807,N_6134);
nor U12271 (N_12271,N_8842,N_7526);
and U12272 (N_12272,N_9336,N_6385);
xnor U12273 (N_12273,N_7531,N_8014);
nor U12274 (N_12274,N_8203,N_6465);
and U12275 (N_12275,N_8872,N_9755);
nand U12276 (N_12276,N_7586,N_7309);
xor U12277 (N_12277,N_5377,N_5573);
and U12278 (N_12278,N_5198,N_8028);
or U12279 (N_12279,N_6400,N_8694);
or U12280 (N_12280,N_9707,N_6663);
and U12281 (N_12281,N_9139,N_8337);
nand U12282 (N_12282,N_7737,N_8563);
nor U12283 (N_12283,N_5582,N_5861);
xor U12284 (N_12284,N_7525,N_8914);
xnor U12285 (N_12285,N_7687,N_5520);
nand U12286 (N_12286,N_5808,N_6068);
or U12287 (N_12287,N_5074,N_9097);
xor U12288 (N_12288,N_8591,N_6750);
nor U12289 (N_12289,N_7549,N_9179);
nand U12290 (N_12290,N_6907,N_7885);
or U12291 (N_12291,N_7169,N_6785);
xor U12292 (N_12292,N_5254,N_6754);
or U12293 (N_12293,N_9568,N_6792);
xor U12294 (N_12294,N_6590,N_8800);
and U12295 (N_12295,N_5042,N_6697);
or U12296 (N_12296,N_5842,N_7378);
nor U12297 (N_12297,N_8575,N_9820);
nand U12298 (N_12298,N_9495,N_8120);
and U12299 (N_12299,N_8004,N_5060);
and U12300 (N_12300,N_7965,N_8020);
and U12301 (N_12301,N_7780,N_6488);
or U12302 (N_12302,N_6939,N_5470);
nand U12303 (N_12303,N_9317,N_8611);
or U12304 (N_12304,N_5795,N_7361);
xor U12305 (N_12305,N_8024,N_9928);
or U12306 (N_12306,N_5522,N_7973);
nand U12307 (N_12307,N_6359,N_6427);
nand U12308 (N_12308,N_5438,N_9537);
and U12309 (N_12309,N_7757,N_9606);
nor U12310 (N_12310,N_6300,N_7339);
nand U12311 (N_12311,N_8995,N_7589);
or U12312 (N_12312,N_6565,N_7334);
nor U12313 (N_12313,N_9476,N_6265);
and U12314 (N_12314,N_6173,N_5705);
nand U12315 (N_12315,N_7121,N_7779);
xor U12316 (N_12316,N_7636,N_5344);
or U12317 (N_12317,N_8504,N_5454);
nor U12318 (N_12318,N_6442,N_9817);
xor U12319 (N_12319,N_6584,N_5262);
and U12320 (N_12320,N_5455,N_6730);
and U12321 (N_12321,N_9144,N_9398);
and U12322 (N_12322,N_9028,N_8731);
xor U12323 (N_12323,N_9033,N_6699);
nor U12324 (N_12324,N_7849,N_8010);
nor U12325 (N_12325,N_6911,N_7948);
or U12326 (N_12326,N_9529,N_7422);
and U12327 (N_12327,N_5102,N_8202);
xor U12328 (N_12328,N_6720,N_8392);
xnor U12329 (N_12329,N_9290,N_7392);
nor U12330 (N_12330,N_9178,N_9307);
nand U12331 (N_12331,N_8753,N_9330);
nand U12332 (N_12332,N_7159,N_9008);
nor U12333 (N_12333,N_7563,N_9133);
nor U12334 (N_12334,N_9985,N_5244);
xor U12335 (N_12335,N_6252,N_9844);
or U12336 (N_12336,N_5973,N_7266);
nand U12337 (N_12337,N_6118,N_5793);
nand U12338 (N_12338,N_9026,N_9551);
nor U12339 (N_12339,N_6668,N_6596);
or U12340 (N_12340,N_7447,N_8638);
nor U12341 (N_12341,N_9472,N_8442);
nor U12342 (N_12342,N_6878,N_7648);
and U12343 (N_12343,N_6507,N_5885);
or U12344 (N_12344,N_5461,N_8616);
and U12345 (N_12345,N_6578,N_9120);
xor U12346 (N_12346,N_8676,N_9126);
or U12347 (N_12347,N_6455,N_9265);
nand U12348 (N_12348,N_6354,N_7933);
nand U12349 (N_12349,N_9051,N_5126);
nor U12350 (N_12350,N_8163,N_6110);
nand U12351 (N_12351,N_9874,N_6943);
or U12352 (N_12352,N_5739,N_7987);
nor U12353 (N_12353,N_6379,N_5965);
xnor U12354 (N_12354,N_6419,N_5593);
or U12355 (N_12355,N_6715,N_9711);
xnor U12356 (N_12356,N_9334,N_9695);
nor U12357 (N_12357,N_7338,N_5109);
and U12358 (N_12358,N_7485,N_5115);
xor U12359 (N_12359,N_9892,N_6220);
nor U12360 (N_12360,N_6680,N_9676);
xnor U12361 (N_12361,N_9249,N_9771);
nand U12362 (N_12362,N_7970,N_8007);
nand U12363 (N_12363,N_8421,N_8483);
xnor U12364 (N_12364,N_7140,N_5020);
xor U12365 (N_12365,N_8015,N_8987);
nor U12366 (N_12366,N_6853,N_5181);
nand U12367 (N_12367,N_7226,N_8191);
or U12368 (N_12368,N_9363,N_7500);
nand U12369 (N_12369,N_8213,N_8919);
xnor U12370 (N_12370,N_8564,N_5726);
nor U12371 (N_12371,N_8131,N_5338);
and U12372 (N_12372,N_6784,N_5692);
or U12373 (N_12373,N_7548,N_5938);
xnor U12374 (N_12374,N_9110,N_8344);
xor U12375 (N_12375,N_5867,N_8426);
and U12376 (N_12376,N_8909,N_6440);
nand U12377 (N_12377,N_8743,N_7881);
and U12378 (N_12378,N_5599,N_8037);
and U12379 (N_12379,N_9185,N_6191);
and U12380 (N_12380,N_6621,N_6953);
nand U12381 (N_12381,N_8679,N_9582);
nand U12382 (N_12382,N_6199,N_7925);
or U12383 (N_12383,N_8804,N_7694);
or U12384 (N_12384,N_9872,N_8928);
and U12385 (N_12385,N_5797,N_8710);
or U12386 (N_12386,N_6958,N_7312);
nor U12387 (N_12387,N_7833,N_8951);
nand U12388 (N_12388,N_9805,N_7335);
and U12389 (N_12389,N_6432,N_5630);
nor U12390 (N_12390,N_9225,N_7294);
xor U12391 (N_12391,N_6609,N_7534);
nor U12392 (N_12392,N_7931,N_8910);
xor U12393 (N_12393,N_5067,N_6099);
or U12394 (N_12394,N_5302,N_9354);
or U12395 (N_12395,N_9333,N_9886);
nor U12396 (N_12396,N_5906,N_7058);
xor U12397 (N_12397,N_7061,N_8139);
nand U12398 (N_12398,N_6390,N_8693);
and U12399 (N_12399,N_8742,N_5788);
and U12400 (N_12400,N_8633,N_5546);
or U12401 (N_12401,N_9343,N_5071);
or U12402 (N_12402,N_6839,N_8689);
and U12403 (N_12403,N_8970,N_7278);
and U12404 (N_12404,N_5050,N_8790);
nor U12405 (N_12405,N_9323,N_6984);
nor U12406 (N_12406,N_8521,N_7137);
nor U12407 (N_12407,N_7620,N_9854);
xnor U12408 (N_12408,N_5661,N_7008);
and U12409 (N_12409,N_5316,N_8425);
or U12410 (N_12410,N_8357,N_8453);
and U12411 (N_12411,N_5723,N_9734);
or U12412 (N_12412,N_6113,N_6299);
or U12413 (N_12413,N_6125,N_8818);
nand U12414 (N_12414,N_7355,N_6973);
nor U12415 (N_12415,N_8101,N_6198);
xnor U12416 (N_12416,N_5160,N_5802);
or U12417 (N_12417,N_5284,N_7227);
xor U12418 (N_12418,N_7736,N_9559);
and U12419 (N_12419,N_7377,N_5992);
nor U12420 (N_12420,N_7015,N_9747);
or U12421 (N_12421,N_7530,N_9950);
and U12422 (N_12422,N_5832,N_8167);
and U12423 (N_12423,N_6435,N_6813);
xor U12424 (N_12424,N_7321,N_9516);
or U12425 (N_12425,N_9090,N_5990);
xor U12426 (N_12426,N_9929,N_5363);
or U12427 (N_12427,N_6271,N_7468);
and U12428 (N_12428,N_6845,N_5373);
xor U12429 (N_12429,N_5610,N_5738);
nand U12430 (N_12430,N_6702,N_6228);
nor U12431 (N_12431,N_8177,N_5999);
nor U12432 (N_12432,N_7917,N_7585);
or U12433 (N_12433,N_8626,N_5943);
nand U12434 (N_12434,N_6589,N_8381);
nor U12435 (N_12435,N_9486,N_9614);
and U12436 (N_12436,N_5146,N_6834);
nand U12437 (N_12437,N_6371,N_9900);
xor U12438 (N_12438,N_6226,N_9397);
nand U12439 (N_12439,N_5446,N_9004);
nor U12440 (N_12440,N_7330,N_6490);
nand U12441 (N_12441,N_7595,N_5200);
nand U12442 (N_12442,N_6184,N_6103);
xnor U12443 (N_12443,N_7697,N_6585);
nand U12444 (N_12444,N_7826,N_7359);
nor U12445 (N_12445,N_5012,N_5929);
and U12446 (N_12446,N_6116,N_9429);
nand U12447 (N_12447,N_5099,N_7985);
nand U12448 (N_12448,N_8643,N_5686);
xnor U12449 (N_12449,N_8534,N_5888);
nand U12450 (N_12450,N_8749,N_8322);
nor U12451 (N_12451,N_8291,N_6241);
xnor U12452 (N_12452,N_6997,N_9313);
nand U12453 (N_12453,N_7938,N_7611);
xnor U12454 (N_12454,N_5531,N_8941);
nand U12455 (N_12455,N_9034,N_8474);
and U12456 (N_12456,N_8216,N_8436);
nand U12457 (N_12457,N_7966,N_7811);
nor U12458 (N_12458,N_8153,N_9896);
and U12459 (N_12459,N_6382,N_7408);
nor U12460 (N_12460,N_7857,N_8762);
xor U12461 (N_12461,N_6886,N_7906);
or U12462 (N_12462,N_9762,N_9702);
xnor U12463 (N_12463,N_6976,N_6830);
and U12464 (N_12464,N_7661,N_5760);
xnor U12465 (N_12465,N_8720,N_5601);
or U12466 (N_12466,N_6903,N_6063);
xor U12467 (N_12467,N_7775,N_6218);
nand U12468 (N_12468,N_5766,N_5156);
nor U12469 (N_12469,N_6352,N_8485);
nor U12470 (N_12470,N_5201,N_8653);
nor U12471 (N_12471,N_5136,N_8480);
and U12472 (N_12472,N_8802,N_9279);
and U12473 (N_12473,N_7892,N_9364);
nor U12474 (N_12474,N_9990,N_9736);
and U12475 (N_12475,N_7562,N_8605);
nand U12476 (N_12476,N_6829,N_8468);
and U12477 (N_12477,N_8130,N_8094);
and U12478 (N_12478,N_7299,N_7124);
xnor U12479 (N_12479,N_7230,N_5458);
and U12480 (N_12480,N_8109,N_9282);
and U12481 (N_12481,N_5934,N_7601);
nor U12482 (N_12482,N_5188,N_9601);
xor U12483 (N_12483,N_9038,N_7761);
nor U12484 (N_12484,N_7152,N_7842);
nand U12485 (N_12485,N_7821,N_6612);
xor U12486 (N_12486,N_8147,N_5530);
nand U12487 (N_12487,N_5441,N_8478);
nand U12488 (N_12488,N_9210,N_9272);
or U12489 (N_12489,N_7900,N_8986);
nor U12490 (N_12490,N_8289,N_7474);
xor U12491 (N_12491,N_9146,N_5409);
and U12492 (N_12492,N_8538,N_7729);
nand U12493 (N_12493,N_8092,N_8713);
and U12494 (N_12494,N_6736,N_7839);
nor U12495 (N_12495,N_9564,N_5009);
nand U12496 (N_12496,N_9776,N_8461);
and U12497 (N_12497,N_5636,N_9880);
or U12498 (N_12498,N_9379,N_7351);
nor U12499 (N_12499,N_8741,N_7303);
nand U12500 (N_12500,N_8694,N_9345);
and U12501 (N_12501,N_7396,N_8256);
or U12502 (N_12502,N_5556,N_8409);
nand U12503 (N_12503,N_9375,N_6612);
xnor U12504 (N_12504,N_7590,N_5839);
xnor U12505 (N_12505,N_8322,N_9251);
nor U12506 (N_12506,N_6160,N_8137);
nand U12507 (N_12507,N_8751,N_5051);
nand U12508 (N_12508,N_6486,N_5800);
nor U12509 (N_12509,N_6844,N_5892);
and U12510 (N_12510,N_8671,N_9459);
or U12511 (N_12511,N_7908,N_7612);
xnor U12512 (N_12512,N_9327,N_5084);
or U12513 (N_12513,N_6918,N_7054);
xor U12514 (N_12514,N_7805,N_8699);
nand U12515 (N_12515,N_6048,N_6688);
and U12516 (N_12516,N_6766,N_6439);
and U12517 (N_12517,N_5866,N_5586);
nor U12518 (N_12518,N_7290,N_9114);
xnor U12519 (N_12519,N_8396,N_6541);
or U12520 (N_12520,N_9384,N_5190);
nor U12521 (N_12521,N_8111,N_8103);
nor U12522 (N_12522,N_8112,N_6749);
xor U12523 (N_12523,N_6853,N_9394);
nand U12524 (N_12524,N_8608,N_9610);
nand U12525 (N_12525,N_8112,N_7559);
nor U12526 (N_12526,N_8174,N_7420);
or U12527 (N_12527,N_5330,N_6236);
or U12528 (N_12528,N_5325,N_6041);
nand U12529 (N_12529,N_5383,N_5911);
or U12530 (N_12530,N_8686,N_6048);
and U12531 (N_12531,N_6571,N_8667);
xnor U12532 (N_12532,N_8339,N_8362);
nand U12533 (N_12533,N_6732,N_7547);
nor U12534 (N_12534,N_7243,N_6524);
or U12535 (N_12535,N_8382,N_9115);
or U12536 (N_12536,N_5684,N_7432);
xor U12537 (N_12537,N_5073,N_7158);
xnor U12538 (N_12538,N_8988,N_6602);
nor U12539 (N_12539,N_9174,N_5433);
and U12540 (N_12540,N_5996,N_9216);
nand U12541 (N_12541,N_9120,N_8978);
or U12542 (N_12542,N_5668,N_9704);
xnor U12543 (N_12543,N_9845,N_7717);
xnor U12544 (N_12544,N_9442,N_8417);
xor U12545 (N_12545,N_6161,N_9186);
nor U12546 (N_12546,N_7122,N_5185);
nor U12547 (N_12547,N_8842,N_9279);
nor U12548 (N_12548,N_8917,N_5129);
or U12549 (N_12549,N_9785,N_8960);
and U12550 (N_12550,N_8725,N_9311);
nor U12551 (N_12551,N_7295,N_5162);
nand U12552 (N_12552,N_8873,N_9375);
nor U12553 (N_12553,N_6356,N_9669);
nand U12554 (N_12554,N_6184,N_6538);
or U12555 (N_12555,N_6891,N_8378);
and U12556 (N_12556,N_8573,N_8169);
nand U12557 (N_12557,N_9968,N_9834);
nand U12558 (N_12558,N_8095,N_8604);
and U12559 (N_12559,N_8499,N_6894);
nor U12560 (N_12560,N_8976,N_5964);
nor U12561 (N_12561,N_5544,N_7677);
xor U12562 (N_12562,N_9264,N_8703);
or U12563 (N_12563,N_6192,N_8726);
nor U12564 (N_12564,N_7448,N_9396);
and U12565 (N_12565,N_7301,N_6697);
and U12566 (N_12566,N_5318,N_5511);
and U12567 (N_12567,N_9929,N_9430);
or U12568 (N_12568,N_5732,N_7247);
xor U12569 (N_12569,N_7170,N_5172);
and U12570 (N_12570,N_5901,N_7898);
or U12571 (N_12571,N_6290,N_6946);
xor U12572 (N_12572,N_7541,N_8908);
nor U12573 (N_12573,N_5898,N_6476);
and U12574 (N_12574,N_7353,N_7857);
xor U12575 (N_12575,N_5051,N_9313);
and U12576 (N_12576,N_7225,N_6196);
and U12577 (N_12577,N_7114,N_7604);
xor U12578 (N_12578,N_9232,N_8478);
xnor U12579 (N_12579,N_7296,N_6824);
or U12580 (N_12580,N_9896,N_5296);
nor U12581 (N_12581,N_8940,N_7504);
nor U12582 (N_12582,N_8950,N_7600);
xor U12583 (N_12583,N_5022,N_6970);
nand U12584 (N_12584,N_9099,N_5551);
nand U12585 (N_12585,N_8895,N_6353);
xnor U12586 (N_12586,N_5700,N_7007);
xor U12587 (N_12587,N_6250,N_6901);
nand U12588 (N_12588,N_5606,N_6158);
nor U12589 (N_12589,N_6709,N_5150);
nor U12590 (N_12590,N_5395,N_6803);
or U12591 (N_12591,N_8542,N_8433);
nand U12592 (N_12592,N_8655,N_9433);
and U12593 (N_12593,N_6553,N_9702);
xnor U12594 (N_12594,N_7232,N_5192);
nor U12595 (N_12595,N_9738,N_7810);
or U12596 (N_12596,N_8218,N_7288);
and U12597 (N_12597,N_9214,N_8722);
nor U12598 (N_12598,N_8409,N_8206);
xnor U12599 (N_12599,N_9732,N_9194);
and U12600 (N_12600,N_5260,N_9426);
nor U12601 (N_12601,N_8980,N_7788);
or U12602 (N_12602,N_9905,N_6667);
xnor U12603 (N_12603,N_5894,N_7079);
nand U12604 (N_12604,N_6471,N_6761);
or U12605 (N_12605,N_9387,N_7225);
and U12606 (N_12606,N_7111,N_5387);
nor U12607 (N_12607,N_6668,N_9443);
and U12608 (N_12608,N_5405,N_6516);
nand U12609 (N_12609,N_6208,N_7661);
or U12610 (N_12610,N_7173,N_5918);
nand U12611 (N_12611,N_6166,N_5205);
nor U12612 (N_12612,N_7464,N_9663);
and U12613 (N_12613,N_9512,N_7172);
nand U12614 (N_12614,N_8981,N_9432);
and U12615 (N_12615,N_9860,N_6763);
or U12616 (N_12616,N_8289,N_8444);
nand U12617 (N_12617,N_7754,N_9328);
nand U12618 (N_12618,N_9585,N_5512);
xnor U12619 (N_12619,N_8557,N_5755);
or U12620 (N_12620,N_9082,N_8972);
nand U12621 (N_12621,N_6155,N_5351);
or U12622 (N_12622,N_6092,N_6728);
xor U12623 (N_12623,N_6597,N_8513);
xnor U12624 (N_12624,N_8676,N_9593);
or U12625 (N_12625,N_7815,N_7467);
nor U12626 (N_12626,N_7140,N_5970);
and U12627 (N_12627,N_9518,N_7545);
or U12628 (N_12628,N_5431,N_6378);
nand U12629 (N_12629,N_7855,N_8958);
and U12630 (N_12630,N_8290,N_7334);
nand U12631 (N_12631,N_6981,N_7328);
and U12632 (N_12632,N_8626,N_6785);
nand U12633 (N_12633,N_9874,N_7987);
nand U12634 (N_12634,N_7948,N_5701);
nor U12635 (N_12635,N_5285,N_5693);
nor U12636 (N_12636,N_5640,N_8992);
and U12637 (N_12637,N_9668,N_7564);
nor U12638 (N_12638,N_5770,N_7275);
or U12639 (N_12639,N_8574,N_8822);
nand U12640 (N_12640,N_7535,N_9763);
nor U12641 (N_12641,N_6494,N_8323);
nand U12642 (N_12642,N_8307,N_8911);
and U12643 (N_12643,N_9521,N_8422);
or U12644 (N_12644,N_5404,N_7882);
or U12645 (N_12645,N_7690,N_9540);
or U12646 (N_12646,N_9743,N_5325);
and U12647 (N_12647,N_6927,N_8126);
and U12648 (N_12648,N_8566,N_7507);
nand U12649 (N_12649,N_8592,N_6917);
or U12650 (N_12650,N_7083,N_5914);
xor U12651 (N_12651,N_6180,N_7896);
nor U12652 (N_12652,N_9625,N_9946);
or U12653 (N_12653,N_7389,N_8473);
nor U12654 (N_12654,N_8869,N_7076);
and U12655 (N_12655,N_7848,N_8966);
and U12656 (N_12656,N_5142,N_6895);
nor U12657 (N_12657,N_5837,N_5285);
xor U12658 (N_12658,N_7711,N_6944);
nand U12659 (N_12659,N_9198,N_9649);
and U12660 (N_12660,N_9642,N_8180);
or U12661 (N_12661,N_9566,N_8709);
nand U12662 (N_12662,N_6460,N_5668);
xnor U12663 (N_12663,N_5479,N_9599);
xor U12664 (N_12664,N_9418,N_5338);
xor U12665 (N_12665,N_6923,N_9233);
nor U12666 (N_12666,N_7769,N_8118);
and U12667 (N_12667,N_5432,N_5399);
nand U12668 (N_12668,N_8406,N_6957);
nand U12669 (N_12669,N_6398,N_9871);
or U12670 (N_12670,N_6782,N_8353);
nor U12671 (N_12671,N_7048,N_6072);
nand U12672 (N_12672,N_6542,N_8181);
nand U12673 (N_12673,N_9371,N_9589);
and U12674 (N_12674,N_8099,N_7306);
or U12675 (N_12675,N_6275,N_7479);
and U12676 (N_12676,N_8651,N_9627);
xnor U12677 (N_12677,N_5754,N_5168);
or U12678 (N_12678,N_6733,N_9857);
and U12679 (N_12679,N_6463,N_9681);
and U12680 (N_12680,N_9045,N_7285);
nand U12681 (N_12681,N_7891,N_5038);
and U12682 (N_12682,N_7009,N_9300);
or U12683 (N_12683,N_9449,N_8813);
or U12684 (N_12684,N_7590,N_5465);
nand U12685 (N_12685,N_9640,N_6232);
or U12686 (N_12686,N_8656,N_7384);
nor U12687 (N_12687,N_8122,N_9843);
or U12688 (N_12688,N_5811,N_5338);
nand U12689 (N_12689,N_7880,N_6878);
or U12690 (N_12690,N_5441,N_5110);
or U12691 (N_12691,N_9856,N_7817);
and U12692 (N_12692,N_7888,N_8656);
nand U12693 (N_12693,N_8844,N_5228);
xnor U12694 (N_12694,N_9613,N_6418);
and U12695 (N_12695,N_5561,N_9288);
nor U12696 (N_12696,N_7719,N_6066);
nand U12697 (N_12697,N_7181,N_5884);
or U12698 (N_12698,N_5776,N_9766);
xnor U12699 (N_12699,N_7923,N_6031);
xnor U12700 (N_12700,N_6011,N_9608);
nand U12701 (N_12701,N_8896,N_5688);
and U12702 (N_12702,N_6369,N_6895);
nand U12703 (N_12703,N_9462,N_9883);
and U12704 (N_12704,N_6362,N_7413);
nand U12705 (N_12705,N_6003,N_5644);
or U12706 (N_12706,N_7408,N_5232);
or U12707 (N_12707,N_5739,N_9738);
and U12708 (N_12708,N_8310,N_8303);
nand U12709 (N_12709,N_9573,N_8192);
nor U12710 (N_12710,N_6101,N_5768);
and U12711 (N_12711,N_5874,N_5788);
nor U12712 (N_12712,N_8479,N_8424);
or U12713 (N_12713,N_9937,N_6828);
nor U12714 (N_12714,N_8010,N_7951);
xnor U12715 (N_12715,N_6747,N_9839);
nor U12716 (N_12716,N_8087,N_5430);
nor U12717 (N_12717,N_9730,N_8720);
nand U12718 (N_12718,N_5855,N_6514);
nor U12719 (N_12719,N_7384,N_7822);
nand U12720 (N_12720,N_8056,N_7036);
or U12721 (N_12721,N_5486,N_6502);
nand U12722 (N_12722,N_9237,N_9110);
nand U12723 (N_12723,N_6925,N_7096);
nor U12724 (N_12724,N_9294,N_7157);
xnor U12725 (N_12725,N_6365,N_5528);
nor U12726 (N_12726,N_5304,N_5068);
nand U12727 (N_12727,N_8569,N_9469);
nor U12728 (N_12728,N_5851,N_8482);
or U12729 (N_12729,N_5307,N_7567);
or U12730 (N_12730,N_9511,N_6782);
and U12731 (N_12731,N_9197,N_7738);
nand U12732 (N_12732,N_7611,N_9948);
nand U12733 (N_12733,N_6726,N_8238);
xor U12734 (N_12734,N_9399,N_5720);
and U12735 (N_12735,N_7103,N_9381);
and U12736 (N_12736,N_8608,N_5214);
nand U12737 (N_12737,N_7236,N_6736);
nand U12738 (N_12738,N_6692,N_9021);
nand U12739 (N_12739,N_5822,N_5012);
or U12740 (N_12740,N_7572,N_8494);
or U12741 (N_12741,N_6815,N_7813);
and U12742 (N_12742,N_9052,N_6644);
or U12743 (N_12743,N_6724,N_7981);
or U12744 (N_12744,N_5285,N_6807);
nor U12745 (N_12745,N_9936,N_8245);
nand U12746 (N_12746,N_6831,N_6149);
nand U12747 (N_12747,N_7540,N_8988);
nand U12748 (N_12748,N_6684,N_8328);
or U12749 (N_12749,N_9695,N_5309);
and U12750 (N_12750,N_7423,N_7594);
nor U12751 (N_12751,N_6395,N_9675);
nor U12752 (N_12752,N_8686,N_5615);
and U12753 (N_12753,N_9597,N_8098);
and U12754 (N_12754,N_8278,N_6756);
and U12755 (N_12755,N_9382,N_8489);
xnor U12756 (N_12756,N_6598,N_9324);
or U12757 (N_12757,N_7725,N_6280);
xnor U12758 (N_12758,N_6928,N_7190);
xnor U12759 (N_12759,N_7718,N_5342);
or U12760 (N_12760,N_7162,N_8172);
and U12761 (N_12761,N_6123,N_5125);
nand U12762 (N_12762,N_9492,N_7417);
or U12763 (N_12763,N_8622,N_5736);
nand U12764 (N_12764,N_6594,N_7737);
nor U12765 (N_12765,N_6470,N_6518);
nor U12766 (N_12766,N_6466,N_9103);
and U12767 (N_12767,N_8975,N_6669);
nand U12768 (N_12768,N_9419,N_7754);
nand U12769 (N_12769,N_9595,N_7102);
nand U12770 (N_12770,N_8791,N_5291);
and U12771 (N_12771,N_7007,N_9970);
nor U12772 (N_12772,N_9752,N_5019);
xnor U12773 (N_12773,N_7365,N_6935);
nor U12774 (N_12774,N_5177,N_9860);
or U12775 (N_12775,N_5667,N_6076);
xnor U12776 (N_12776,N_6370,N_7190);
xor U12777 (N_12777,N_8556,N_7066);
xor U12778 (N_12778,N_5725,N_8640);
nor U12779 (N_12779,N_7996,N_7347);
and U12780 (N_12780,N_7320,N_5916);
or U12781 (N_12781,N_8414,N_5783);
and U12782 (N_12782,N_7203,N_6676);
nor U12783 (N_12783,N_6192,N_7306);
nor U12784 (N_12784,N_9497,N_5272);
nor U12785 (N_12785,N_6339,N_8122);
xor U12786 (N_12786,N_9239,N_9968);
and U12787 (N_12787,N_6115,N_5491);
or U12788 (N_12788,N_7189,N_7815);
or U12789 (N_12789,N_8192,N_9875);
nand U12790 (N_12790,N_7184,N_9838);
and U12791 (N_12791,N_8733,N_5955);
nand U12792 (N_12792,N_7178,N_5869);
nand U12793 (N_12793,N_8888,N_6831);
nor U12794 (N_12794,N_9575,N_5204);
nand U12795 (N_12795,N_8736,N_8827);
or U12796 (N_12796,N_8102,N_9291);
and U12797 (N_12797,N_6729,N_7189);
nand U12798 (N_12798,N_6875,N_9924);
and U12799 (N_12799,N_6630,N_6615);
nor U12800 (N_12800,N_6267,N_5058);
and U12801 (N_12801,N_6380,N_9918);
or U12802 (N_12802,N_5921,N_5225);
xnor U12803 (N_12803,N_5365,N_6110);
nand U12804 (N_12804,N_5654,N_6538);
nand U12805 (N_12805,N_5013,N_7774);
nand U12806 (N_12806,N_9017,N_5796);
nor U12807 (N_12807,N_6464,N_6491);
nand U12808 (N_12808,N_9218,N_7793);
nand U12809 (N_12809,N_7021,N_9004);
xnor U12810 (N_12810,N_9199,N_7399);
or U12811 (N_12811,N_8267,N_6011);
nand U12812 (N_12812,N_7981,N_9707);
xor U12813 (N_12813,N_5579,N_5252);
xor U12814 (N_12814,N_8517,N_9897);
or U12815 (N_12815,N_5728,N_8388);
and U12816 (N_12816,N_8221,N_8638);
and U12817 (N_12817,N_5731,N_9008);
nor U12818 (N_12818,N_5622,N_6488);
xnor U12819 (N_12819,N_8366,N_8534);
nand U12820 (N_12820,N_7532,N_5825);
nand U12821 (N_12821,N_5474,N_9043);
xor U12822 (N_12822,N_5701,N_7882);
xnor U12823 (N_12823,N_5247,N_8939);
and U12824 (N_12824,N_6573,N_7812);
nand U12825 (N_12825,N_9978,N_5743);
and U12826 (N_12826,N_8262,N_7506);
xnor U12827 (N_12827,N_8861,N_8492);
and U12828 (N_12828,N_8770,N_8324);
nand U12829 (N_12829,N_8044,N_7480);
xor U12830 (N_12830,N_7874,N_9921);
nor U12831 (N_12831,N_5398,N_9163);
nand U12832 (N_12832,N_7229,N_7041);
and U12833 (N_12833,N_7640,N_7006);
xor U12834 (N_12834,N_8732,N_7561);
nand U12835 (N_12835,N_7895,N_7282);
and U12836 (N_12836,N_7908,N_5853);
or U12837 (N_12837,N_8200,N_6267);
xnor U12838 (N_12838,N_7165,N_9635);
nand U12839 (N_12839,N_9826,N_9835);
nand U12840 (N_12840,N_5769,N_8960);
nand U12841 (N_12841,N_5076,N_7972);
and U12842 (N_12842,N_7933,N_7078);
nand U12843 (N_12843,N_7612,N_5597);
or U12844 (N_12844,N_5061,N_9373);
nor U12845 (N_12845,N_8311,N_9867);
or U12846 (N_12846,N_8668,N_9712);
or U12847 (N_12847,N_8561,N_8000);
nand U12848 (N_12848,N_5558,N_5153);
or U12849 (N_12849,N_8055,N_8558);
and U12850 (N_12850,N_7843,N_6439);
xor U12851 (N_12851,N_6497,N_5591);
or U12852 (N_12852,N_6452,N_7558);
nor U12853 (N_12853,N_8198,N_8164);
or U12854 (N_12854,N_6322,N_8691);
and U12855 (N_12855,N_8030,N_7810);
nor U12856 (N_12856,N_5092,N_9232);
xnor U12857 (N_12857,N_9944,N_5836);
xor U12858 (N_12858,N_6622,N_9210);
nor U12859 (N_12859,N_8102,N_8097);
xnor U12860 (N_12860,N_9227,N_6099);
or U12861 (N_12861,N_6131,N_9301);
and U12862 (N_12862,N_8967,N_5471);
nor U12863 (N_12863,N_5256,N_5634);
and U12864 (N_12864,N_7283,N_8271);
xnor U12865 (N_12865,N_9686,N_7140);
and U12866 (N_12866,N_7002,N_8951);
and U12867 (N_12867,N_5649,N_8878);
and U12868 (N_12868,N_6554,N_9817);
or U12869 (N_12869,N_5012,N_7937);
xor U12870 (N_12870,N_9300,N_7257);
nand U12871 (N_12871,N_8087,N_8506);
nand U12872 (N_12872,N_8272,N_8774);
or U12873 (N_12873,N_8990,N_8793);
nor U12874 (N_12874,N_6819,N_5435);
xnor U12875 (N_12875,N_9556,N_6981);
or U12876 (N_12876,N_7821,N_5885);
or U12877 (N_12877,N_5959,N_8478);
nand U12878 (N_12878,N_7510,N_6894);
or U12879 (N_12879,N_7981,N_8320);
or U12880 (N_12880,N_6818,N_6754);
or U12881 (N_12881,N_6854,N_8484);
nor U12882 (N_12882,N_8884,N_5798);
xor U12883 (N_12883,N_5686,N_6367);
nand U12884 (N_12884,N_6870,N_5126);
xnor U12885 (N_12885,N_7741,N_7776);
and U12886 (N_12886,N_5436,N_7001);
nor U12887 (N_12887,N_5524,N_8819);
nand U12888 (N_12888,N_8852,N_9512);
nand U12889 (N_12889,N_6745,N_5745);
and U12890 (N_12890,N_8387,N_7440);
or U12891 (N_12891,N_6773,N_8066);
xnor U12892 (N_12892,N_5897,N_9483);
and U12893 (N_12893,N_6224,N_9684);
and U12894 (N_12894,N_5275,N_8117);
or U12895 (N_12895,N_8091,N_5209);
nand U12896 (N_12896,N_5862,N_8000);
or U12897 (N_12897,N_7093,N_5292);
or U12898 (N_12898,N_6195,N_5392);
nand U12899 (N_12899,N_6577,N_5406);
nand U12900 (N_12900,N_9314,N_6557);
xor U12901 (N_12901,N_5094,N_5019);
xor U12902 (N_12902,N_5969,N_7622);
xnor U12903 (N_12903,N_5178,N_5832);
nand U12904 (N_12904,N_7280,N_6246);
or U12905 (N_12905,N_5070,N_9204);
or U12906 (N_12906,N_7256,N_9070);
and U12907 (N_12907,N_7522,N_7415);
nor U12908 (N_12908,N_7897,N_7774);
or U12909 (N_12909,N_6132,N_8008);
nor U12910 (N_12910,N_9399,N_9537);
nor U12911 (N_12911,N_7703,N_6568);
or U12912 (N_12912,N_8890,N_8216);
xor U12913 (N_12913,N_5828,N_5751);
or U12914 (N_12914,N_6034,N_7390);
or U12915 (N_12915,N_6494,N_5068);
and U12916 (N_12916,N_6257,N_5405);
or U12917 (N_12917,N_5026,N_8276);
and U12918 (N_12918,N_9227,N_6586);
nor U12919 (N_12919,N_8027,N_9751);
nand U12920 (N_12920,N_5065,N_7605);
xor U12921 (N_12921,N_6395,N_8619);
nor U12922 (N_12922,N_8131,N_8566);
and U12923 (N_12923,N_6757,N_8975);
xor U12924 (N_12924,N_9144,N_5060);
nor U12925 (N_12925,N_5476,N_7300);
nor U12926 (N_12926,N_9763,N_9855);
xnor U12927 (N_12927,N_9230,N_8266);
xnor U12928 (N_12928,N_8326,N_5337);
nand U12929 (N_12929,N_6454,N_7559);
nand U12930 (N_12930,N_5510,N_6925);
xnor U12931 (N_12931,N_8894,N_8433);
nand U12932 (N_12932,N_9783,N_5001);
and U12933 (N_12933,N_8318,N_5302);
xnor U12934 (N_12934,N_6028,N_7838);
and U12935 (N_12935,N_9897,N_5724);
and U12936 (N_12936,N_7249,N_7004);
and U12937 (N_12937,N_5259,N_6965);
and U12938 (N_12938,N_8579,N_5064);
nor U12939 (N_12939,N_8092,N_5275);
and U12940 (N_12940,N_8003,N_6089);
nor U12941 (N_12941,N_7619,N_5336);
nand U12942 (N_12942,N_8616,N_7051);
nand U12943 (N_12943,N_9013,N_6558);
and U12944 (N_12944,N_8338,N_6762);
xnor U12945 (N_12945,N_9769,N_7167);
xnor U12946 (N_12946,N_9937,N_8378);
nor U12947 (N_12947,N_7989,N_8893);
or U12948 (N_12948,N_9545,N_6765);
or U12949 (N_12949,N_8887,N_9464);
xor U12950 (N_12950,N_5541,N_8840);
nor U12951 (N_12951,N_7456,N_8789);
xor U12952 (N_12952,N_5511,N_8215);
or U12953 (N_12953,N_9316,N_5941);
xnor U12954 (N_12954,N_8983,N_5182);
or U12955 (N_12955,N_9780,N_5629);
nand U12956 (N_12956,N_7681,N_9831);
or U12957 (N_12957,N_8803,N_9772);
and U12958 (N_12958,N_8364,N_8772);
nor U12959 (N_12959,N_8493,N_5579);
or U12960 (N_12960,N_9021,N_8600);
or U12961 (N_12961,N_5460,N_9316);
xnor U12962 (N_12962,N_7954,N_9464);
xnor U12963 (N_12963,N_6038,N_7155);
nand U12964 (N_12964,N_9628,N_5141);
and U12965 (N_12965,N_6265,N_6273);
nor U12966 (N_12966,N_6536,N_5886);
xor U12967 (N_12967,N_6544,N_7813);
or U12968 (N_12968,N_9666,N_5986);
xnor U12969 (N_12969,N_6668,N_9357);
nor U12970 (N_12970,N_7146,N_7014);
nand U12971 (N_12971,N_7968,N_7092);
or U12972 (N_12972,N_7431,N_7147);
nand U12973 (N_12973,N_7829,N_9003);
and U12974 (N_12974,N_6751,N_6058);
nand U12975 (N_12975,N_7401,N_5255);
and U12976 (N_12976,N_8178,N_7977);
nor U12977 (N_12977,N_9424,N_6006);
and U12978 (N_12978,N_8387,N_7202);
nand U12979 (N_12979,N_6211,N_8971);
and U12980 (N_12980,N_7197,N_5730);
or U12981 (N_12981,N_9027,N_9433);
and U12982 (N_12982,N_8318,N_9246);
nor U12983 (N_12983,N_7395,N_9768);
xor U12984 (N_12984,N_9916,N_7997);
and U12985 (N_12985,N_9332,N_7169);
or U12986 (N_12986,N_8409,N_6466);
and U12987 (N_12987,N_6218,N_8665);
xnor U12988 (N_12988,N_6370,N_5784);
and U12989 (N_12989,N_7820,N_7526);
xnor U12990 (N_12990,N_7240,N_9670);
and U12991 (N_12991,N_7583,N_5167);
xnor U12992 (N_12992,N_6440,N_7864);
and U12993 (N_12993,N_9602,N_9589);
and U12994 (N_12994,N_6600,N_6425);
or U12995 (N_12995,N_5140,N_8559);
or U12996 (N_12996,N_5507,N_8962);
nand U12997 (N_12997,N_5375,N_9100);
or U12998 (N_12998,N_6919,N_9489);
and U12999 (N_12999,N_7296,N_7793);
and U13000 (N_13000,N_6281,N_8245);
nor U13001 (N_13001,N_7774,N_8562);
and U13002 (N_13002,N_7360,N_5145);
xnor U13003 (N_13003,N_8065,N_9109);
xor U13004 (N_13004,N_7992,N_8365);
xnor U13005 (N_13005,N_7053,N_7196);
nor U13006 (N_13006,N_6299,N_9778);
nand U13007 (N_13007,N_8468,N_9844);
xnor U13008 (N_13008,N_9219,N_7270);
nor U13009 (N_13009,N_6463,N_7470);
nand U13010 (N_13010,N_5179,N_8561);
nand U13011 (N_13011,N_7127,N_7261);
or U13012 (N_13012,N_5902,N_8700);
or U13013 (N_13013,N_5588,N_5490);
nor U13014 (N_13014,N_7299,N_5599);
or U13015 (N_13015,N_8736,N_9640);
xor U13016 (N_13016,N_7164,N_5037);
or U13017 (N_13017,N_6485,N_7358);
and U13018 (N_13018,N_5374,N_8664);
or U13019 (N_13019,N_9727,N_8420);
and U13020 (N_13020,N_5401,N_6724);
xnor U13021 (N_13021,N_9682,N_5745);
nand U13022 (N_13022,N_5653,N_9905);
nor U13023 (N_13023,N_7229,N_9033);
nand U13024 (N_13024,N_6729,N_9382);
xor U13025 (N_13025,N_9490,N_8191);
nor U13026 (N_13026,N_5559,N_5336);
or U13027 (N_13027,N_6034,N_9184);
and U13028 (N_13028,N_5149,N_7074);
nor U13029 (N_13029,N_7295,N_5016);
nor U13030 (N_13030,N_9187,N_8495);
or U13031 (N_13031,N_6199,N_6825);
and U13032 (N_13032,N_8441,N_6406);
nor U13033 (N_13033,N_6931,N_5783);
or U13034 (N_13034,N_7535,N_9767);
xor U13035 (N_13035,N_8933,N_8237);
and U13036 (N_13036,N_7080,N_5415);
nor U13037 (N_13037,N_5341,N_9310);
nor U13038 (N_13038,N_9832,N_6158);
nor U13039 (N_13039,N_8740,N_7132);
nand U13040 (N_13040,N_9855,N_5916);
or U13041 (N_13041,N_5644,N_9049);
and U13042 (N_13042,N_9970,N_5372);
or U13043 (N_13043,N_6466,N_9687);
or U13044 (N_13044,N_5750,N_9321);
xnor U13045 (N_13045,N_8237,N_8871);
or U13046 (N_13046,N_7888,N_8496);
or U13047 (N_13047,N_6385,N_6625);
or U13048 (N_13048,N_8246,N_9545);
or U13049 (N_13049,N_7631,N_9551);
nor U13050 (N_13050,N_8514,N_8604);
and U13051 (N_13051,N_9595,N_9402);
and U13052 (N_13052,N_5261,N_7332);
xnor U13053 (N_13053,N_7447,N_8018);
xor U13054 (N_13054,N_8157,N_8666);
and U13055 (N_13055,N_9006,N_5508);
xnor U13056 (N_13056,N_8069,N_6225);
nor U13057 (N_13057,N_6795,N_8540);
nand U13058 (N_13058,N_8263,N_9086);
and U13059 (N_13059,N_8954,N_8541);
and U13060 (N_13060,N_8826,N_6960);
nand U13061 (N_13061,N_5986,N_5390);
nand U13062 (N_13062,N_9926,N_7342);
and U13063 (N_13063,N_7426,N_6475);
nand U13064 (N_13064,N_5566,N_9265);
xnor U13065 (N_13065,N_9904,N_6289);
xor U13066 (N_13066,N_9344,N_7947);
and U13067 (N_13067,N_5265,N_8949);
nor U13068 (N_13068,N_9960,N_6709);
nand U13069 (N_13069,N_5983,N_6868);
nand U13070 (N_13070,N_9172,N_8927);
or U13071 (N_13071,N_5936,N_6874);
and U13072 (N_13072,N_5608,N_6881);
nor U13073 (N_13073,N_5960,N_8860);
xnor U13074 (N_13074,N_7759,N_6754);
or U13075 (N_13075,N_5876,N_9494);
nand U13076 (N_13076,N_9030,N_8779);
xor U13077 (N_13077,N_7519,N_7837);
or U13078 (N_13078,N_5002,N_9919);
and U13079 (N_13079,N_6166,N_6467);
and U13080 (N_13080,N_6108,N_6782);
and U13081 (N_13081,N_9880,N_9127);
or U13082 (N_13082,N_6408,N_9836);
and U13083 (N_13083,N_5746,N_7615);
or U13084 (N_13084,N_5347,N_6667);
or U13085 (N_13085,N_6916,N_6849);
nor U13086 (N_13086,N_8510,N_9519);
or U13087 (N_13087,N_6276,N_5698);
nand U13088 (N_13088,N_6587,N_5146);
nor U13089 (N_13089,N_5463,N_6719);
and U13090 (N_13090,N_6587,N_5401);
nor U13091 (N_13091,N_5077,N_6760);
nand U13092 (N_13092,N_5644,N_9182);
or U13093 (N_13093,N_8968,N_6820);
nor U13094 (N_13094,N_9679,N_9779);
nor U13095 (N_13095,N_5927,N_9644);
or U13096 (N_13096,N_7346,N_7093);
and U13097 (N_13097,N_7447,N_6243);
and U13098 (N_13098,N_9784,N_8826);
and U13099 (N_13099,N_9687,N_6758);
or U13100 (N_13100,N_6678,N_5525);
xor U13101 (N_13101,N_7931,N_7816);
nand U13102 (N_13102,N_8309,N_5993);
nand U13103 (N_13103,N_9091,N_9955);
and U13104 (N_13104,N_6988,N_7551);
xnor U13105 (N_13105,N_5097,N_6031);
nor U13106 (N_13106,N_9441,N_6481);
nand U13107 (N_13107,N_9185,N_5079);
nor U13108 (N_13108,N_9360,N_8337);
nor U13109 (N_13109,N_6240,N_6785);
nor U13110 (N_13110,N_7477,N_6034);
and U13111 (N_13111,N_9643,N_8191);
or U13112 (N_13112,N_8146,N_5244);
nor U13113 (N_13113,N_6156,N_7929);
xnor U13114 (N_13114,N_5147,N_5030);
or U13115 (N_13115,N_6867,N_8123);
nor U13116 (N_13116,N_7478,N_5473);
xor U13117 (N_13117,N_8327,N_7103);
and U13118 (N_13118,N_5535,N_8249);
and U13119 (N_13119,N_7933,N_8577);
nor U13120 (N_13120,N_8935,N_7622);
xor U13121 (N_13121,N_8995,N_9263);
xor U13122 (N_13122,N_5298,N_6862);
or U13123 (N_13123,N_5349,N_8212);
nor U13124 (N_13124,N_9127,N_7597);
or U13125 (N_13125,N_6929,N_9895);
nor U13126 (N_13126,N_9420,N_9777);
and U13127 (N_13127,N_6986,N_8311);
and U13128 (N_13128,N_9674,N_6204);
xor U13129 (N_13129,N_7645,N_7861);
and U13130 (N_13130,N_6377,N_7506);
nand U13131 (N_13131,N_9519,N_9195);
or U13132 (N_13132,N_9667,N_7180);
xnor U13133 (N_13133,N_8487,N_5024);
xnor U13134 (N_13134,N_5596,N_5929);
or U13135 (N_13135,N_8550,N_5744);
or U13136 (N_13136,N_6758,N_9908);
or U13137 (N_13137,N_5022,N_7690);
xnor U13138 (N_13138,N_5785,N_9121);
nand U13139 (N_13139,N_7797,N_5581);
or U13140 (N_13140,N_9889,N_9031);
or U13141 (N_13141,N_9863,N_6701);
nand U13142 (N_13142,N_6189,N_9528);
nor U13143 (N_13143,N_8126,N_8035);
xnor U13144 (N_13144,N_6084,N_6533);
or U13145 (N_13145,N_9956,N_9534);
xor U13146 (N_13146,N_8832,N_9620);
or U13147 (N_13147,N_8866,N_8623);
nor U13148 (N_13148,N_9046,N_9627);
nand U13149 (N_13149,N_9427,N_6208);
nor U13150 (N_13150,N_8642,N_8649);
xor U13151 (N_13151,N_5106,N_8694);
xnor U13152 (N_13152,N_6282,N_9063);
xor U13153 (N_13153,N_6205,N_9099);
nand U13154 (N_13154,N_6185,N_8788);
or U13155 (N_13155,N_6463,N_8557);
nor U13156 (N_13156,N_8503,N_5294);
nand U13157 (N_13157,N_5436,N_7528);
or U13158 (N_13158,N_5912,N_8361);
or U13159 (N_13159,N_8694,N_5504);
or U13160 (N_13160,N_9795,N_9775);
nand U13161 (N_13161,N_5244,N_7245);
xnor U13162 (N_13162,N_6873,N_8151);
xor U13163 (N_13163,N_9799,N_6706);
and U13164 (N_13164,N_5063,N_6357);
nor U13165 (N_13165,N_6352,N_6109);
xnor U13166 (N_13166,N_8331,N_8523);
and U13167 (N_13167,N_6922,N_8768);
or U13168 (N_13168,N_7532,N_9788);
nand U13169 (N_13169,N_7985,N_7824);
and U13170 (N_13170,N_7506,N_5582);
and U13171 (N_13171,N_8565,N_6485);
nand U13172 (N_13172,N_7829,N_6688);
or U13173 (N_13173,N_5942,N_8633);
xor U13174 (N_13174,N_8797,N_7488);
xnor U13175 (N_13175,N_5284,N_5977);
nand U13176 (N_13176,N_7512,N_6349);
nor U13177 (N_13177,N_8211,N_7011);
or U13178 (N_13178,N_9517,N_7177);
xor U13179 (N_13179,N_7568,N_9710);
and U13180 (N_13180,N_8037,N_5090);
nor U13181 (N_13181,N_6232,N_5715);
nor U13182 (N_13182,N_7274,N_7663);
nand U13183 (N_13183,N_5163,N_6433);
and U13184 (N_13184,N_9887,N_8015);
and U13185 (N_13185,N_8850,N_6288);
and U13186 (N_13186,N_7289,N_9650);
or U13187 (N_13187,N_9215,N_9912);
nor U13188 (N_13188,N_6192,N_5884);
nand U13189 (N_13189,N_5159,N_5971);
nand U13190 (N_13190,N_6804,N_9807);
and U13191 (N_13191,N_5075,N_7563);
or U13192 (N_13192,N_9490,N_5190);
and U13193 (N_13193,N_7355,N_7790);
or U13194 (N_13194,N_8587,N_8016);
xnor U13195 (N_13195,N_6828,N_9810);
or U13196 (N_13196,N_7444,N_6143);
nor U13197 (N_13197,N_5565,N_9977);
or U13198 (N_13198,N_9331,N_9142);
or U13199 (N_13199,N_8088,N_9256);
or U13200 (N_13200,N_7766,N_7001);
and U13201 (N_13201,N_6310,N_5661);
nor U13202 (N_13202,N_9807,N_5111);
or U13203 (N_13203,N_6928,N_9294);
nand U13204 (N_13204,N_5111,N_9315);
nand U13205 (N_13205,N_6151,N_7183);
nand U13206 (N_13206,N_8164,N_8367);
and U13207 (N_13207,N_6161,N_6167);
or U13208 (N_13208,N_5009,N_8889);
and U13209 (N_13209,N_7740,N_5639);
nand U13210 (N_13210,N_7303,N_5477);
nor U13211 (N_13211,N_6146,N_7326);
or U13212 (N_13212,N_8765,N_8058);
nor U13213 (N_13213,N_9775,N_7933);
or U13214 (N_13214,N_7573,N_7466);
and U13215 (N_13215,N_7128,N_5080);
and U13216 (N_13216,N_5463,N_7913);
nand U13217 (N_13217,N_6390,N_5421);
and U13218 (N_13218,N_7723,N_7730);
nor U13219 (N_13219,N_7241,N_6906);
or U13220 (N_13220,N_9881,N_5608);
xor U13221 (N_13221,N_5371,N_6317);
and U13222 (N_13222,N_9377,N_6922);
xnor U13223 (N_13223,N_6560,N_6739);
nand U13224 (N_13224,N_8746,N_9109);
and U13225 (N_13225,N_8919,N_6134);
or U13226 (N_13226,N_7474,N_6207);
xor U13227 (N_13227,N_6784,N_7475);
or U13228 (N_13228,N_7088,N_8353);
nor U13229 (N_13229,N_7225,N_7205);
nand U13230 (N_13230,N_6682,N_5504);
or U13231 (N_13231,N_7858,N_9216);
nand U13232 (N_13232,N_7884,N_8222);
nand U13233 (N_13233,N_8648,N_8418);
or U13234 (N_13234,N_5186,N_6923);
nand U13235 (N_13235,N_9053,N_5360);
xnor U13236 (N_13236,N_7559,N_8903);
nor U13237 (N_13237,N_6627,N_6703);
nor U13238 (N_13238,N_8420,N_5992);
or U13239 (N_13239,N_6357,N_5703);
xor U13240 (N_13240,N_6437,N_6741);
nor U13241 (N_13241,N_9458,N_7716);
xor U13242 (N_13242,N_7296,N_9421);
xor U13243 (N_13243,N_7905,N_9177);
and U13244 (N_13244,N_5367,N_9260);
or U13245 (N_13245,N_6915,N_8531);
and U13246 (N_13246,N_8854,N_9786);
nor U13247 (N_13247,N_6208,N_5516);
nor U13248 (N_13248,N_5246,N_7972);
and U13249 (N_13249,N_7886,N_8798);
xor U13250 (N_13250,N_6649,N_9340);
xor U13251 (N_13251,N_9397,N_5105);
xnor U13252 (N_13252,N_6788,N_6253);
and U13253 (N_13253,N_7848,N_7269);
or U13254 (N_13254,N_8124,N_6341);
or U13255 (N_13255,N_6500,N_6169);
xor U13256 (N_13256,N_7827,N_5993);
xor U13257 (N_13257,N_6334,N_5414);
nand U13258 (N_13258,N_6054,N_8650);
xnor U13259 (N_13259,N_8479,N_9921);
xor U13260 (N_13260,N_9996,N_6313);
nor U13261 (N_13261,N_6517,N_9362);
nor U13262 (N_13262,N_6146,N_8637);
nor U13263 (N_13263,N_7387,N_7861);
nand U13264 (N_13264,N_8332,N_6790);
nor U13265 (N_13265,N_5499,N_6304);
or U13266 (N_13266,N_5923,N_8942);
xor U13267 (N_13267,N_6583,N_5245);
xor U13268 (N_13268,N_7915,N_9602);
xnor U13269 (N_13269,N_7754,N_7284);
xor U13270 (N_13270,N_7859,N_5894);
nor U13271 (N_13271,N_6630,N_6866);
and U13272 (N_13272,N_6424,N_8490);
or U13273 (N_13273,N_8732,N_7600);
and U13274 (N_13274,N_8853,N_6352);
xor U13275 (N_13275,N_7918,N_5407);
nor U13276 (N_13276,N_5928,N_6115);
and U13277 (N_13277,N_7839,N_8861);
and U13278 (N_13278,N_8706,N_8421);
nor U13279 (N_13279,N_8881,N_5792);
xnor U13280 (N_13280,N_5116,N_9748);
and U13281 (N_13281,N_9782,N_7213);
and U13282 (N_13282,N_7454,N_7329);
nor U13283 (N_13283,N_8831,N_7928);
xor U13284 (N_13284,N_8766,N_6193);
and U13285 (N_13285,N_5213,N_8540);
and U13286 (N_13286,N_5202,N_5256);
nand U13287 (N_13287,N_8952,N_7056);
and U13288 (N_13288,N_6649,N_9268);
nor U13289 (N_13289,N_7222,N_5578);
and U13290 (N_13290,N_5777,N_8370);
nand U13291 (N_13291,N_9648,N_7841);
nand U13292 (N_13292,N_9586,N_7828);
nor U13293 (N_13293,N_6858,N_7650);
nand U13294 (N_13294,N_8809,N_8079);
nor U13295 (N_13295,N_8008,N_9584);
xnor U13296 (N_13296,N_9504,N_5884);
nand U13297 (N_13297,N_9891,N_6970);
nor U13298 (N_13298,N_9125,N_5028);
nand U13299 (N_13299,N_6174,N_6586);
nor U13300 (N_13300,N_6233,N_6518);
nor U13301 (N_13301,N_8175,N_6570);
nor U13302 (N_13302,N_9741,N_9159);
or U13303 (N_13303,N_5952,N_5578);
nand U13304 (N_13304,N_9950,N_7367);
nand U13305 (N_13305,N_9592,N_6927);
and U13306 (N_13306,N_7288,N_8772);
nor U13307 (N_13307,N_8386,N_5065);
or U13308 (N_13308,N_6297,N_7021);
or U13309 (N_13309,N_8868,N_8378);
or U13310 (N_13310,N_7654,N_9405);
xor U13311 (N_13311,N_9942,N_6605);
or U13312 (N_13312,N_9938,N_8307);
xor U13313 (N_13313,N_7982,N_8821);
nor U13314 (N_13314,N_8575,N_7902);
and U13315 (N_13315,N_6688,N_7455);
nand U13316 (N_13316,N_9969,N_6456);
and U13317 (N_13317,N_5747,N_5455);
xnor U13318 (N_13318,N_9391,N_5307);
xnor U13319 (N_13319,N_9296,N_7066);
xor U13320 (N_13320,N_7559,N_5652);
or U13321 (N_13321,N_9999,N_6004);
xor U13322 (N_13322,N_7801,N_6841);
nand U13323 (N_13323,N_9071,N_6275);
and U13324 (N_13324,N_7944,N_7164);
and U13325 (N_13325,N_6083,N_5111);
xnor U13326 (N_13326,N_7043,N_9412);
and U13327 (N_13327,N_8591,N_6710);
and U13328 (N_13328,N_7905,N_7890);
and U13329 (N_13329,N_6609,N_5480);
or U13330 (N_13330,N_9992,N_8062);
xnor U13331 (N_13331,N_9180,N_6159);
and U13332 (N_13332,N_9986,N_5461);
or U13333 (N_13333,N_6632,N_6964);
nand U13334 (N_13334,N_8245,N_5065);
and U13335 (N_13335,N_5098,N_5255);
or U13336 (N_13336,N_8180,N_5069);
and U13337 (N_13337,N_7066,N_7519);
and U13338 (N_13338,N_5834,N_7660);
xor U13339 (N_13339,N_8592,N_7878);
or U13340 (N_13340,N_6536,N_7677);
nand U13341 (N_13341,N_7913,N_7679);
nor U13342 (N_13342,N_7970,N_5816);
and U13343 (N_13343,N_7255,N_8337);
or U13344 (N_13344,N_9145,N_5115);
nor U13345 (N_13345,N_7773,N_7177);
nor U13346 (N_13346,N_6810,N_7611);
and U13347 (N_13347,N_7664,N_6834);
xnor U13348 (N_13348,N_9809,N_8316);
or U13349 (N_13349,N_6424,N_9534);
nor U13350 (N_13350,N_5262,N_7212);
xnor U13351 (N_13351,N_9335,N_6688);
or U13352 (N_13352,N_5513,N_8938);
nor U13353 (N_13353,N_5369,N_9356);
or U13354 (N_13354,N_9566,N_6827);
nand U13355 (N_13355,N_7097,N_8673);
or U13356 (N_13356,N_6285,N_7648);
nor U13357 (N_13357,N_8718,N_8834);
nand U13358 (N_13358,N_5154,N_6256);
nor U13359 (N_13359,N_7740,N_9059);
or U13360 (N_13360,N_8156,N_8404);
nor U13361 (N_13361,N_7652,N_9056);
or U13362 (N_13362,N_6182,N_8338);
xnor U13363 (N_13363,N_8170,N_5997);
nand U13364 (N_13364,N_9597,N_5148);
nor U13365 (N_13365,N_8770,N_9361);
and U13366 (N_13366,N_6498,N_8355);
or U13367 (N_13367,N_6927,N_9423);
nand U13368 (N_13368,N_7508,N_8344);
or U13369 (N_13369,N_7364,N_8337);
nor U13370 (N_13370,N_5337,N_6147);
nand U13371 (N_13371,N_7755,N_8050);
nand U13372 (N_13372,N_9674,N_7536);
nand U13373 (N_13373,N_8344,N_9484);
or U13374 (N_13374,N_6481,N_8819);
nand U13375 (N_13375,N_6161,N_7756);
xor U13376 (N_13376,N_8814,N_7781);
nor U13377 (N_13377,N_8136,N_5436);
nor U13378 (N_13378,N_5603,N_5757);
nand U13379 (N_13379,N_8773,N_8361);
xor U13380 (N_13380,N_9566,N_5388);
nor U13381 (N_13381,N_6674,N_5233);
nor U13382 (N_13382,N_7962,N_6454);
nor U13383 (N_13383,N_5880,N_7295);
or U13384 (N_13384,N_5324,N_6701);
xor U13385 (N_13385,N_5838,N_5762);
and U13386 (N_13386,N_6681,N_9561);
nor U13387 (N_13387,N_7056,N_8136);
and U13388 (N_13388,N_8261,N_8128);
nor U13389 (N_13389,N_8296,N_7648);
nor U13390 (N_13390,N_7544,N_8071);
and U13391 (N_13391,N_7196,N_9572);
and U13392 (N_13392,N_7151,N_8750);
or U13393 (N_13393,N_8920,N_6728);
or U13394 (N_13394,N_5984,N_7098);
or U13395 (N_13395,N_6128,N_5213);
or U13396 (N_13396,N_9412,N_7669);
nor U13397 (N_13397,N_9447,N_5594);
nand U13398 (N_13398,N_7577,N_9966);
or U13399 (N_13399,N_5612,N_5721);
nor U13400 (N_13400,N_6230,N_9102);
or U13401 (N_13401,N_5114,N_5972);
nor U13402 (N_13402,N_7855,N_5232);
nor U13403 (N_13403,N_9870,N_6502);
nand U13404 (N_13404,N_7318,N_6018);
and U13405 (N_13405,N_8569,N_6379);
nor U13406 (N_13406,N_6712,N_5659);
nand U13407 (N_13407,N_9553,N_8495);
nand U13408 (N_13408,N_7748,N_8419);
nand U13409 (N_13409,N_6991,N_6752);
and U13410 (N_13410,N_6005,N_6121);
nand U13411 (N_13411,N_5997,N_5042);
xnor U13412 (N_13412,N_5210,N_8001);
and U13413 (N_13413,N_8503,N_7214);
or U13414 (N_13414,N_5061,N_9426);
or U13415 (N_13415,N_8588,N_8536);
and U13416 (N_13416,N_6567,N_6235);
xor U13417 (N_13417,N_9985,N_5126);
nand U13418 (N_13418,N_5318,N_9333);
nand U13419 (N_13419,N_7879,N_6105);
or U13420 (N_13420,N_6942,N_6499);
xnor U13421 (N_13421,N_8756,N_9309);
and U13422 (N_13422,N_5632,N_9070);
and U13423 (N_13423,N_9710,N_6940);
nor U13424 (N_13424,N_7584,N_6213);
xor U13425 (N_13425,N_8420,N_5129);
xnor U13426 (N_13426,N_8969,N_5979);
or U13427 (N_13427,N_6122,N_8312);
or U13428 (N_13428,N_8175,N_9870);
and U13429 (N_13429,N_7856,N_6540);
and U13430 (N_13430,N_8249,N_7002);
nor U13431 (N_13431,N_8869,N_5668);
and U13432 (N_13432,N_5555,N_8988);
nor U13433 (N_13433,N_5861,N_8681);
nor U13434 (N_13434,N_9874,N_8984);
or U13435 (N_13435,N_8777,N_7012);
or U13436 (N_13436,N_9309,N_9044);
or U13437 (N_13437,N_8033,N_7463);
nand U13438 (N_13438,N_8202,N_7010);
nand U13439 (N_13439,N_7352,N_8835);
nor U13440 (N_13440,N_6015,N_7820);
or U13441 (N_13441,N_9310,N_7248);
and U13442 (N_13442,N_7517,N_8973);
xor U13443 (N_13443,N_7017,N_5347);
nand U13444 (N_13444,N_8233,N_8173);
nand U13445 (N_13445,N_9337,N_5371);
xor U13446 (N_13446,N_8564,N_5809);
and U13447 (N_13447,N_6771,N_9059);
or U13448 (N_13448,N_6723,N_5710);
nor U13449 (N_13449,N_7319,N_7411);
or U13450 (N_13450,N_9001,N_8013);
xnor U13451 (N_13451,N_9940,N_7011);
xor U13452 (N_13452,N_8336,N_5765);
or U13453 (N_13453,N_5495,N_8274);
xor U13454 (N_13454,N_9096,N_9823);
and U13455 (N_13455,N_6005,N_9779);
or U13456 (N_13456,N_9627,N_6788);
or U13457 (N_13457,N_5624,N_7147);
and U13458 (N_13458,N_6743,N_7591);
or U13459 (N_13459,N_9068,N_9911);
nand U13460 (N_13460,N_8305,N_5611);
or U13461 (N_13461,N_5702,N_8338);
or U13462 (N_13462,N_9916,N_7281);
and U13463 (N_13463,N_5669,N_9283);
nor U13464 (N_13464,N_7995,N_9541);
xnor U13465 (N_13465,N_6621,N_6976);
nand U13466 (N_13466,N_6591,N_6270);
nor U13467 (N_13467,N_8033,N_8001);
nor U13468 (N_13468,N_5866,N_5225);
or U13469 (N_13469,N_5733,N_7984);
nand U13470 (N_13470,N_9446,N_5312);
nor U13471 (N_13471,N_9009,N_5765);
or U13472 (N_13472,N_6170,N_7439);
and U13473 (N_13473,N_9622,N_7080);
nor U13474 (N_13474,N_5585,N_7895);
and U13475 (N_13475,N_5015,N_6116);
nor U13476 (N_13476,N_8040,N_6448);
nor U13477 (N_13477,N_5965,N_8649);
and U13478 (N_13478,N_6801,N_8480);
xnor U13479 (N_13479,N_5066,N_6464);
or U13480 (N_13480,N_8969,N_6113);
and U13481 (N_13481,N_8082,N_6759);
or U13482 (N_13482,N_8402,N_5885);
or U13483 (N_13483,N_5659,N_6759);
and U13484 (N_13484,N_7748,N_7102);
nand U13485 (N_13485,N_8227,N_8302);
nand U13486 (N_13486,N_9477,N_9347);
nand U13487 (N_13487,N_9278,N_7649);
and U13488 (N_13488,N_9966,N_9297);
nand U13489 (N_13489,N_7746,N_7732);
xnor U13490 (N_13490,N_9870,N_8263);
or U13491 (N_13491,N_5160,N_6201);
or U13492 (N_13492,N_5725,N_9823);
xor U13493 (N_13493,N_5295,N_5996);
nor U13494 (N_13494,N_6567,N_8050);
or U13495 (N_13495,N_5499,N_6681);
xor U13496 (N_13496,N_8550,N_5321);
xor U13497 (N_13497,N_7768,N_5249);
and U13498 (N_13498,N_8280,N_7220);
xor U13499 (N_13499,N_5375,N_5366);
and U13500 (N_13500,N_6389,N_8771);
and U13501 (N_13501,N_9097,N_7739);
nand U13502 (N_13502,N_5237,N_5997);
xnor U13503 (N_13503,N_9043,N_5476);
and U13504 (N_13504,N_8515,N_7822);
xor U13505 (N_13505,N_9049,N_9375);
and U13506 (N_13506,N_6956,N_9108);
and U13507 (N_13507,N_8896,N_8084);
and U13508 (N_13508,N_7207,N_8829);
nor U13509 (N_13509,N_9982,N_9367);
or U13510 (N_13510,N_7498,N_8697);
xor U13511 (N_13511,N_8508,N_5724);
and U13512 (N_13512,N_6074,N_8613);
nor U13513 (N_13513,N_9323,N_6565);
nor U13514 (N_13514,N_9456,N_9610);
or U13515 (N_13515,N_8933,N_8761);
nor U13516 (N_13516,N_7391,N_8055);
nand U13517 (N_13517,N_6207,N_5163);
and U13518 (N_13518,N_5045,N_5368);
or U13519 (N_13519,N_8802,N_9551);
nand U13520 (N_13520,N_5056,N_5008);
nand U13521 (N_13521,N_5934,N_9140);
xor U13522 (N_13522,N_5107,N_5824);
nor U13523 (N_13523,N_7518,N_6130);
xor U13524 (N_13524,N_7267,N_7204);
nor U13525 (N_13525,N_9760,N_6190);
and U13526 (N_13526,N_6364,N_9724);
and U13527 (N_13527,N_8892,N_8531);
and U13528 (N_13528,N_6894,N_8684);
nand U13529 (N_13529,N_8655,N_7732);
and U13530 (N_13530,N_8946,N_7833);
nand U13531 (N_13531,N_6808,N_8588);
nand U13532 (N_13532,N_8632,N_8266);
or U13533 (N_13533,N_8244,N_5567);
nand U13534 (N_13534,N_7382,N_8689);
and U13535 (N_13535,N_9978,N_7424);
nor U13536 (N_13536,N_7319,N_8073);
xnor U13537 (N_13537,N_7726,N_9522);
nor U13538 (N_13538,N_7278,N_9471);
xor U13539 (N_13539,N_9998,N_5573);
xnor U13540 (N_13540,N_7606,N_7943);
and U13541 (N_13541,N_6524,N_5842);
or U13542 (N_13542,N_8356,N_7068);
and U13543 (N_13543,N_8060,N_5966);
and U13544 (N_13544,N_7791,N_5801);
nand U13545 (N_13545,N_5123,N_8131);
nor U13546 (N_13546,N_5375,N_5125);
and U13547 (N_13547,N_8949,N_9720);
nand U13548 (N_13548,N_5219,N_5759);
nor U13549 (N_13549,N_8480,N_7537);
nor U13550 (N_13550,N_8397,N_5939);
nor U13551 (N_13551,N_9553,N_6635);
nor U13552 (N_13552,N_8149,N_8179);
nor U13553 (N_13553,N_8696,N_8564);
and U13554 (N_13554,N_7587,N_6706);
xnor U13555 (N_13555,N_7764,N_5878);
xnor U13556 (N_13556,N_5164,N_7948);
and U13557 (N_13557,N_7514,N_6823);
xor U13558 (N_13558,N_5477,N_8263);
nor U13559 (N_13559,N_6118,N_5590);
nand U13560 (N_13560,N_7227,N_5315);
nor U13561 (N_13561,N_6158,N_5558);
nand U13562 (N_13562,N_7298,N_5255);
nor U13563 (N_13563,N_8664,N_5184);
nor U13564 (N_13564,N_9741,N_6041);
and U13565 (N_13565,N_8087,N_7342);
xor U13566 (N_13566,N_6804,N_9714);
nand U13567 (N_13567,N_8369,N_6366);
or U13568 (N_13568,N_6690,N_9279);
and U13569 (N_13569,N_6564,N_5172);
xnor U13570 (N_13570,N_6943,N_9381);
and U13571 (N_13571,N_9582,N_7339);
nand U13572 (N_13572,N_6997,N_9721);
and U13573 (N_13573,N_8516,N_9146);
nor U13574 (N_13574,N_5914,N_5975);
and U13575 (N_13575,N_5817,N_8534);
nand U13576 (N_13576,N_9416,N_8726);
xnor U13577 (N_13577,N_6545,N_6140);
and U13578 (N_13578,N_7850,N_9797);
and U13579 (N_13579,N_6621,N_7321);
or U13580 (N_13580,N_9742,N_6954);
nand U13581 (N_13581,N_8900,N_8870);
nand U13582 (N_13582,N_6040,N_5776);
nand U13583 (N_13583,N_8883,N_9645);
or U13584 (N_13584,N_8425,N_8220);
nand U13585 (N_13585,N_7475,N_7324);
xor U13586 (N_13586,N_8444,N_7523);
nand U13587 (N_13587,N_5496,N_6717);
xor U13588 (N_13588,N_7762,N_6050);
nor U13589 (N_13589,N_9193,N_7709);
nand U13590 (N_13590,N_8083,N_7103);
nand U13591 (N_13591,N_8704,N_7192);
nor U13592 (N_13592,N_8814,N_8795);
and U13593 (N_13593,N_8350,N_5739);
or U13594 (N_13594,N_6403,N_6909);
xor U13595 (N_13595,N_7291,N_9456);
nand U13596 (N_13596,N_9221,N_7882);
and U13597 (N_13597,N_5006,N_6311);
xor U13598 (N_13598,N_5935,N_8696);
and U13599 (N_13599,N_7737,N_5185);
or U13600 (N_13600,N_5364,N_9912);
nand U13601 (N_13601,N_5439,N_5354);
xor U13602 (N_13602,N_7932,N_8285);
and U13603 (N_13603,N_5748,N_6688);
xnor U13604 (N_13604,N_7668,N_7504);
and U13605 (N_13605,N_5262,N_8394);
or U13606 (N_13606,N_9730,N_8916);
xnor U13607 (N_13607,N_7279,N_5065);
nor U13608 (N_13608,N_7516,N_8414);
nand U13609 (N_13609,N_9340,N_6091);
or U13610 (N_13610,N_9620,N_8215);
or U13611 (N_13611,N_5782,N_9586);
xnor U13612 (N_13612,N_9318,N_5317);
nor U13613 (N_13613,N_5587,N_5875);
xor U13614 (N_13614,N_8564,N_6841);
nor U13615 (N_13615,N_9115,N_9362);
xnor U13616 (N_13616,N_5357,N_7903);
and U13617 (N_13617,N_8412,N_9128);
and U13618 (N_13618,N_6888,N_5780);
xor U13619 (N_13619,N_9975,N_5846);
nor U13620 (N_13620,N_7708,N_8790);
nand U13621 (N_13621,N_8470,N_5771);
nand U13622 (N_13622,N_9751,N_9548);
nand U13623 (N_13623,N_9998,N_5504);
and U13624 (N_13624,N_6650,N_5292);
and U13625 (N_13625,N_8306,N_6939);
and U13626 (N_13626,N_7609,N_6871);
xor U13627 (N_13627,N_8321,N_5558);
or U13628 (N_13628,N_5253,N_9087);
xnor U13629 (N_13629,N_6046,N_8210);
nand U13630 (N_13630,N_7971,N_5024);
or U13631 (N_13631,N_5889,N_9713);
or U13632 (N_13632,N_9970,N_7201);
nand U13633 (N_13633,N_6649,N_8395);
or U13634 (N_13634,N_7230,N_6449);
or U13635 (N_13635,N_9966,N_6394);
nor U13636 (N_13636,N_6280,N_8272);
nor U13637 (N_13637,N_8113,N_8731);
nor U13638 (N_13638,N_9292,N_7867);
nand U13639 (N_13639,N_5416,N_8594);
nand U13640 (N_13640,N_5037,N_9097);
xnor U13641 (N_13641,N_7470,N_5263);
or U13642 (N_13642,N_8413,N_7280);
xor U13643 (N_13643,N_7652,N_9247);
xor U13644 (N_13644,N_7296,N_8373);
xnor U13645 (N_13645,N_7842,N_5314);
or U13646 (N_13646,N_9225,N_7229);
and U13647 (N_13647,N_9810,N_6167);
nand U13648 (N_13648,N_6305,N_7104);
xnor U13649 (N_13649,N_7230,N_6622);
nand U13650 (N_13650,N_5576,N_5152);
and U13651 (N_13651,N_9652,N_5105);
nor U13652 (N_13652,N_9297,N_6930);
or U13653 (N_13653,N_9719,N_5682);
or U13654 (N_13654,N_9763,N_5679);
or U13655 (N_13655,N_6171,N_6045);
xnor U13656 (N_13656,N_8761,N_8744);
or U13657 (N_13657,N_9015,N_9017);
xnor U13658 (N_13658,N_5148,N_8336);
and U13659 (N_13659,N_9031,N_7161);
xor U13660 (N_13660,N_7531,N_8713);
xnor U13661 (N_13661,N_6577,N_7426);
xnor U13662 (N_13662,N_6849,N_9931);
nand U13663 (N_13663,N_9974,N_5780);
and U13664 (N_13664,N_8906,N_6184);
nand U13665 (N_13665,N_9731,N_6879);
and U13666 (N_13666,N_5547,N_7372);
nor U13667 (N_13667,N_5808,N_6590);
nand U13668 (N_13668,N_6640,N_6241);
or U13669 (N_13669,N_9344,N_5632);
or U13670 (N_13670,N_7442,N_7093);
xnor U13671 (N_13671,N_7029,N_5838);
and U13672 (N_13672,N_7268,N_6844);
nand U13673 (N_13673,N_9400,N_6667);
nand U13674 (N_13674,N_8667,N_6940);
nand U13675 (N_13675,N_7508,N_9844);
xnor U13676 (N_13676,N_5480,N_5339);
or U13677 (N_13677,N_7593,N_8646);
and U13678 (N_13678,N_7710,N_8374);
xor U13679 (N_13679,N_8347,N_5004);
or U13680 (N_13680,N_9060,N_7352);
nor U13681 (N_13681,N_5388,N_6725);
nand U13682 (N_13682,N_7438,N_9646);
nor U13683 (N_13683,N_9008,N_5893);
or U13684 (N_13684,N_9361,N_7937);
and U13685 (N_13685,N_9953,N_7237);
nand U13686 (N_13686,N_9534,N_9774);
xor U13687 (N_13687,N_6300,N_7997);
nor U13688 (N_13688,N_9139,N_9234);
or U13689 (N_13689,N_8898,N_6074);
or U13690 (N_13690,N_7594,N_9634);
and U13691 (N_13691,N_6878,N_8560);
or U13692 (N_13692,N_8399,N_5952);
xor U13693 (N_13693,N_6746,N_6424);
and U13694 (N_13694,N_9557,N_6983);
or U13695 (N_13695,N_6480,N_9739);
nand U13696 (N_13696,N_8026,N_8577);
or U13697 (N_13697,N_9525,N_8136);
nor U13698 (N_13698,N_5636,N_8242);
xnor U13699 (N_13699,N_7973,N_7411);
nor U13700 (N_13700,N_9262,N_8140);
and U13701 (N_13701,N_7440,N_8116);
and U13702 (N_13702,N_9965,N_8078);
and U13703 (N_13703,N_7633,N_5303);
nand U13704 (N_13704,N_7346,N_9185);
or U13705 (N_13705,N_7871,N_7875);
nor U13706 (N_13706,N_7962,N_8967);
and U13707 (N_13707,N_8224,N_6785);
and U13708 (N_13708,N_5512,N_6406);
xor U13709 (N_13709,N_9206,N_7599);
nand U13710 (N_13710,N_6202,N_9670);
nor U13711 (N_13711,N_7756,N_8082);
nor U13712 (N_13712,N_6605,N_8913);
and U13713 (N_13713,N_5156,N_5430);
nor U13714 (N_13714,N_9912,N_7463);
nand U13715 (N_13715,N_7244,N_9912);
or U13716 (N_13716,N_8626,N_7472);
nor U13717 (N_13717,N_7843,N_5214);
and U13718 (N_13718,N_8657,N_7947);
nand U13719 (N_13719,N_6428,N_7104);
nor U13720 (N_13720,N_8006,N_8610);
or U13721 (N_13721,N_6160,N_9928);
or U13722 (N_13722,N_5098,N_7176);
nor U13723 (N_13723,N_8782,N_8723);
nand U13724 (N_13724,N_6484,N_6448);
and U13725 (N_13725,N_9895,N_6976);
nand U13726 (N_13726,N_7822,N_7396);
nor U13727 (N_13727,N_8054,N_7335);
xnor U13728 (N_13728,N_6779,N_5273);
nand U13729 (N_13729,N_8457,N_5549);
nor U13730 (N_13730,N_7256,N_7200);
and U13731 (N_13731,N_5801,N_6364);
or U13732 (N_13732,N_5925,N_6257);
nand U13733 (N_13733,N_7728,N_8233);
and U13734 (N_13734,N_8695,N_9508);
nor U13735 (N_13735,N_9899,N_6904);
nand U13736 (N_13736,N_8068,N_7894);
nor U13737 (N_13737,N_6668,N_8491);
xor U13738 (N_13738,N_7683,N_9724);
and U13739 (N_13739,N_7244,N_8739);
nor U13740 (N_13740,N_7585,N_9427);
nand U13741 (N_13741,N_9240,N_7958);
xor U13742 (N_13742,N_7166,N_6196);
xor U13743 (N_13743,N_9985,N_6551);
xor U13744 (N_13744,N_8171,N_8949);
or U13745 (N_13745,N_7379,N_8408);
xnor U13746 (N_13746,N_9619,N_7362);
nand U13747 (N_13747,N_8648,N_8377);
nand U13748 (N_13748,N_5875,N_8956);
and U13749 (N_13749,N_7129,N_8762);
and U13750 (N_13750,N_8941,N_7069);
nor U13751 (N_13751,N_6771,N_6018);
nor U13752 (N_13752,N_6353,N_6703);
nand U13753 (N_13753,N_7088,N_7364);
nand U13754 (N_13754,N_5938,N_5249);
or U13755 (N_13755,N_8574,N_8804);
and U13756 (N_13756,N_7890,N_6706);
or U13757 (N_13757,N_6900,N_9058);
nand U13758 (N_13758,N_5916,N_9267);
or U13759 (N_13759,N_5698,N_9475);
nand U13760 (N_13760,N_8921,N_8665);
and U13761 (N_13761,N_8634,N_5680);
nor U13762 (N_13762,N_6527,N_5962);
nor U13763 (N_13763,N_9690,N_8681);
or U13764 (N_13764,N_7372,N_5280);
nor U13765 (N_13765,N_9093,N_5685);
xor U13766 (N_13766,N_5594,N_5833);
or U13767 (N_13767,N_6141,N_6248);
nand U13768 (N_13768,N_6564,N_7766);
or U13769 (N_13769,N_8343,N_9053);
nand U13770 (N_13770,N_7183,N_7384);
nor U13771 (N_13771,N_7908,N_8547);
and U13772 (N_13772,N_5546,N_5425);
xnor U13773 (N_13773,N_9250,N_8685);
xnor U13774 (N_13774,N_6834,N_8462);
nor U13775 (N_13775,N_7699,N_9595);
xor U13776 (N_13776,N_8558,N_8383);
xor U13777 (N_13777,N_9965,N_5041);
nor U13778 (N_13778,N_9833,N_5356);
and U13779 (N_13779,N_8453,N_9775);
xnor U13780 (N_13780,N_8395,N_8457);
nand U13781 (N_13781,N_5392,N_5138);
and U13782 (N_13782,N_8634,N_5494);
xnor U13783 (N_13783,N_8700,N_6112);
or U13784 (N_13784,N_8927,N_6102);
or U13785 (N_13785,N_6100,N_7268);
nand U13786 (N_13786,N_7193,N_6092);
and U13787 (N_13787,N_7729,N_9203);
and U13788 (N_13788,N_7073,N_5158);
nor U13789 (N_13789,N_7050,N_6129);
nor U13790 (N_13790,N_7161,N_6144);
xor U13791 (N_13791,N_6170,N_6419);
nand U13792 (N_13792,N_6466,N_7922);
nor U13793 (N_13793,N_7333,N_5066);
or U13794 (N_13794,N_9217,N_8094);
nor U13795 (N_13795,N_9434,N_9069);
nor U13796 (N_13796,N_7505,N_5026);
xnor U13797 (N_13797,N_5474,N_7072);
xnor U13798 (N_13798,N_7925,N_7146);
nor U13799 (N_13799,N_7670,N_7522);
nand U13800 (N_13800,N_8597,N_8593);
nand U13801 (N_13801,N_6781,N_6071);
or U13802 (N_13802,N_7524,N_7085);
and U13803 (N_13803,N_7207,N_6723);
nor U13804 (N_13804,N_5684,N_6547);
and U13805 (N_13805,N_5919,N_9737);
or U13806 (N_13806,N_5334,N_7393);
or U13807 (N_13807,N_5298,N_8967);
or U13808 (N_13808,N_5745,N_8413);
xor U13809 (N_13809,N_5202,N_5416);
or U13810 (N_13810,N_9373,N_5615);
nand U13811 (N_13811,N_8442,N_8490);
or U13812 (N_13812,N_9387,N_6988);
xnor U13813 (N_13813,N_8371,N_8316);
nor U13814 (N_13814,N_9973,N_5755);
and U13815 (N_13815,N_6536,N_9160);
nand U13816 (N_13816,N_5635,N_8686);
and U13817 (N_13817,N_7224,N_6055);
and U13818 (N_13818,N_5645,N_9918);
or U13819 (N_13819,N_9951,N_6291);
or U13820 (N_13820,N_8174,N_9400);
or U13821 (N_13821,N_5397,N_6058);
and U13822 (N_13822,N_8630,N_9779);
xor U13823 (N_13823,N_7980,N_5072);
xor U13824 (N_13824,N_9008,N_8461);
nand U13825 (N_13825,N_9721,N_6134);
or U13826 (N_13826,N_5231,N_5340);
xnor U13827 (N_13827,N_6018,N_7733);
nor U13828 (N_13828,N_6211,N_9617);
nor U13829 (N_13829,N_9241,N_8619);
or U13830 (N_13830,N_6338,N_5483);
or U13831 (N_13831,N_7057,N_7085);
or U13832 (N_13832,N_5068,N_8302);
and U13833 (N_13833,N_6140,N_8023);
nand U13834 (N_13834,N_6715,N_8328);
nor U13835 (N_13835,N_7454,N_6081);
xor U13836 (N_13836,N_9345,N_8611);
and U13837 (N_13837,N_5669,N_8958);
or U13838 (N_13838,N_9424,N_5773);
nand U13839 (N_13839,N_8890,N_9281);
xnor U13840 (N_13840,N_7869,N_7332);
nand U13841 (N_13841,N_9660,N_5977);
nand U13842 (N_13842,N_9614,N_9587);
and U13843 (N_13843,N_7176,N_6790);
nand U13844 (N_13844,N_7326,N_5895);
nor U13845 (N_13845,N_9317,N_9579);
and U13846 (N_13846,N_8098,N_9150);
nor U13847 (N_13847,N_7473,N_7385);
nor U13848 (N_13848,N_7298,N_7678);
nor U13849 (N_13849,N_5121,N_7821);
nor U13850 (N_13850,N_8587,N_6332);
or U13851 (N_13851,N_5529,N_8514);
nor U13852 (N_13852,N_5898,N_7522);
and U13853 (N_13853,N_6848,N_7904);
xor U13854 (N_13854,N_8024,N_9320);
nand U13855 (N_13855,N_7492,N_8790);
xor U13856 (N_13856,N_9194,N_7168);
xor U13857 (N_13857,N_8621,N_5800);
nand U13858 (N_13858,N_6989,N_9387);
xnor U13859 (N_13859,N_6906,N_6167);
nor U13860 (N_13860,N_8275,N_7753);
nand U13861 (N_13861,N_6288,N_7983);
xor U13862 (N_13862,N_9698,N_5415);
and U13863 (N_13863,N_5239,N_5139);
nor U13864 (N_13864,N_6278,N_8989);
xnor U13865 (N_13865,N_6534,N_8177);
or U13866 (N_13866,N_7536,N_8199);
xnor U13867 (N_13867,N_8421,N_9529);
and U13868 (N_13868,N_8903,N_5851);
nand U13869 (N_13869,N_5914,N_5206);
and U13870 (N_13870,N_9085,N_8150);
and U13871 (N_13871,N_8373,N_9345);
or U13872 (N_13872,N_8792,N_5940);
nor U13873 (N_13873,N_9739,N_7750);
or U13874 (N_13874,N_5784,N_7906);
nand U13875 (N_13875,N_9263,N_8972);
or U13876 (N_13876,N_8151,N_7679);
nand U13877 (N_13877,N_5616,N_7534);
xnor U13878 (N_13878,N_9329,N_7652);
nand U13879 (N_13879,N_5113,N_9223);
and U13880 (N_13880,N_8620,N_8538);
nor U13881 (N_13881,N_5893,N_8849);
xor U13882 (N_13882,N_7340,N_9717);
xor U13883 (N_13883,N_7590,N_8965);
nand U13884 (N_13884,N_5399,N_8258);
and U13885 (N_13885,N_8213,N_7530);
and U13886 (N_13886,N_9442,N_9303);
or U13887 (N_13887,N_9307,N_6280);
nand U13888 (N_13888,N_6647,N_5285);
xor U13889 (N_13889,N_6597,N_9156);
or U13890 (N_13890,N_8903,N_8990);
nand U13891 (N_13891,N_8950,N_6711);
nand U13892 (N_13892,N_8996,N_8170);
xnor U13893 (N_13893,N_5644,N_8331);
or U13894 (N_13894,N_6221,N_8778);
and U13895 (N_13895,N_7447,N_6290);
xor U13896 (N_13896,N_6380,N_9774);
xnor U13897 (N_13897,N_6428,N_8309);
or U13898 (N_13898,N_8521,N_6980);
nand U13899 (N_13899,N_5856,N_8215);
and U13900 (N_13900,N_7206,N_8892);
nor U13901 (N_13901,N_9681,N_5835);
xnor U13902 (N_13902,N_9863,N_7177);
and U13903 (N_13903,N_6833,N_8287);
nor U13904 (N_13904,N_5647,N_5085);
xnor U13905 (N_13905,N_7071,N_9570);
and U13906 (N_13906,N_5755,N_9138);
nand U13907 (N_13907,N_7452,N_5746);
or U13908 (N_13908,N_5581,N_6544);
xor U13909 (N_13909,N_6242,N_7814);
xor U13910 (N_13910,N_7775,N_5511);
nor U13911 (N_13911,N_7532,N_9417);
or U13912 (N_13912,N_7409,N_5379);
nand U13913 (N_13913,N_8209,N_9541);
and U13914 (N_13914,N_9899,N_6979);
nor U13915 (N_13915,N_7836,N_6568);
xnor U13916 (N_13916,N_5173,N_6091);
nand U13917 (N_13917,N_8618,N_6036);
nand U13918 (N_13918,N_7840,N_6733);
xor U13919 (N_13919,N_6618,N_5635);
xor U13920 (N_13920,N_7237,N_9198);
nor U13921 (N_13921,N_7683,N_8466);
xor U13922 (N_13922,N_8092,N_7100);
nor U13923 (N_13923,N_6670,N_5136);
nand U13924 (N_13924,N_6226,N_7232);
and U13925 (N_13925,N_8850,N_9079);
nand U13926 (N_13926,N_9396,N_6658);
xor U13927 (N_13927,N_5049,N_7427);
or U13928 (N_13928,N_8691,N_5480);
xor U13929 (N_13929,N_8618,N_6281);
nor U13930 (N_13930,N_6129,N_8718);
nand U13931 (N_13931,N_7375,N_8615);
xnor U13932 (N_13932,N_8184,N_7750);
xnor U13933 (N_13933,N_9552,N_9993);
or U13934 (N_13934,N_8958,N_8535);
or U13935 (N_13935,N_5710,N_8386);
nand U13936 (N_13936,N_8379,N_8192);
or U13937 (N_13937,N_8945,N_8547);
xnor U13938 (N_13938,N_8246,N_9091);
nor U13939 (N_13939,N_5846,N_9017);
nor U13940 (N_13940,N_7063,N_8050);
xnor U13941 (N_13941,N_9088,N_9425);
nand U13942 (N_13942,N_6886,N_8962);
nand U13943 (N_13943,N_9502,N_6470);
nor U13944 (N_13944,N_8710,N_6695);
xor U13945 (N_13945,N_8786,N_8156);
nor U13946 (N_13946,N_6501,N_6427);
nor U13947 (N_13947,N_5226,N_8384);
nor U13948 (N_13948,N_5866,N_8115);
or U13949 (N_13949,N_7561,N_6368);
nand U13950 (N_13950,N_7681,N_7187);
nand U13951 (N_13951,N_7389,N_5759);
nor U13952 (N_13952,N_7342,N_5865);
xnor U13953 (N_13953,N_5745,N_5323);
or U13954 (N_13954,N_7135,N_8598);
or U13955 (N_13955,N_6704,N_6068);
or U13956 (N_13956,N_8748,N_5513);
or U13957 (N_13957,N_7740,N_5719);
and U13958 (N_13958,N_8047,N_5688);
and U13959 (N_13959,N_9004,N_9840);
nor U13960 (N_13960,N_6180,N_9003);
nor U13961 (N_13961,N_8703,N_6341);
xor U13962 (N_13962,N_7400,N_6267);
and U13963 (N_13963,N_7936,N_8605);
or U13964 (N_13964,N_7792,N_9693);
nor U13965 (N_13965,N_6385,N_8802);
xor U13966 (N_13966,N_9865,N_9737);
or U13967 (N_13967,N_5754,N_7037);
and U13968 (N_13968,N_9438,N_5812);
nor U13969 (N_13969,N_5440,N_8979);
xnor U13970 (N_13970,N_8383,N_9916);
xor U13971 (N_13971,N_7374,N_6227);
and U13972 (N_13972,N_7109,N_9932);
or U13973 (N_13973,N_5996,N_9979);
xor U13974 (N_13974,N_9236,N_5720);
and U13975 (N_13975,N_9062,N_5371);
xnor U13976 (N_13976,N_9745,N_6441);
xor U13977 (N_13977,N_9118,N_7199);
xor U13978 (N_13978,N_9220,N_5374);
xor U13979 (N_13979,N_5152,N_7452);
nand U13980 (N_13980,N_7710,N_7824);
or U13981 (N_13981,N_6470,N_5762);
xor U13982 (N_13982,N_7843,N_8439);
nand U13983 (N_13983,N_8906,N_7899);
nor U13984 (N_13984,N_6199,N_9619);
or U13985 (N_13985,N_8095,N_7471);
and U13986 (N_13986,N_5749,N_7445);
nor U13987 (N_13987,N_5480,N_9685);
nand U13988 (N_13988,N_9009,N_5079);
and U13989 (N_13989,N_9788,N_8150);
nor U13990 (N_13990,N_6414,N_8915);
and U13991 (N_13991,N_7748,N_9981);
and U13992 (N_13992,N_9110,N_7528);
or U13993 (N_13993,N_6338,N_9093);
and U13994 (N_13994,N_7015,N_8249);
or U13995 (N_13995,N_8133,N_5023);
or U13996 (N_13996,N_6575,N_9261);
nand U13997 (N_13997,N_5373,N_7959);
nor U13998 (N_13998,N_7386,N_9487);
nor U13999 (N_13999,N_9277,N_8984);
xnor U14000 (N_14000,N_5558,N_7773);
xnor U14001 (N_14001,N_5188,N_6116);
and U14002 (N_14002,N_9767,N_9019);
nand U14003 (N_14003,N_9603,N_7389);
nand U14004 (N_14004,N_7565,N_7254);
nand U14005 (N_14005,N_7089,N_7077);
nand U14006 (N_14006,N_6265,N_6725);
nor U14007 (N_14007,N_9788,N_5026);
or U14008 (N_14008,N_6127,N_7254);
or U14009 (N_14009,N_8230,N_5354);
nand U14010 (N_14010,N_7465,N_5535);
nand U14011 (N_14011,N_8107,N_5434);
nor U14012 (N_14012,N_7936,N_5028);
nor U14013 (N_14013,N_5979,N_8053);
and U14014 (N_14014,N_5359,N_5280);
or U14015 (N_14015,N_7328,N_7182);
or U14016 (N_14016,N_7156,N_6322);
nor U14017 (N_14017,N_5794,N_5994);
and U14018 (N_14018,N_8791,N_6838);
xor U14019 (N_14019,N_6158,N_9686);
and U14020 (N_14020,N_9950,N_7841);
nor U14021 (N_14021,N_8430,N_6254);
nand U14022 (N_14022,N_9489,N_6363);
or U14023 (N_14023,N_7938,N_5066);
nand U14024 (N_14024,N_5310,N_8285);
or U14025 (N_14025,N_8622,N_7503);
nor U14026 (N_14026,N_8280,N_5128);
nand U14027 (N_14027,N_6201,N_9809);
nor U14028 (N_14028,N_8945,N_5832);
nor U14029 (N_14029,N_5093,N_6756);
xnor U14030 (N_14030,N_7380,N_7492);
or U14031 (N_14031,N_7502,N_9776);
and U14032 (N_14032,N_8313,N_7876);
and U14033 (N_14033,N_5717,N_6663);
and U14034 (N_14034,N_7603,N_9836);
nand U14035 (N_14035,N_6166,N_6869);
xnor U14036 (N_14036,N_8291,N_6644);
nand U14037 (N_14037,N_8467,N_6435);
xnor U14038 (N_14038,N_5517,N_8349);
nand U14039 (N_14039,N_7719,N_9576);
or U14040 (N_14040,N_9717,N_8251);
nand U14041 (N_14041,N_9975,N_6240);
or U14042 (N_14042,N_5097,N_7517);
and U14043 (N_14043,N_7688,N_9971);
nor U14044 (N_14044,N_9942,N_9199);
xnor U14045 (N_14045,N_8494,N_8049);
nand U14046 (N_14046,N_9761,N_9100);
and U14047 (N_14047,N_9974,N_9154);
nand U14048 (N_14048,N_8531,N_5668);
or U14049 (N_14049,N_5724,N_7657);
or U14050 (N_14050,N_7459,N_6507);
xnor U14051 (N_14051,N_5884,N_5018);
nor U14052 (N_14052,N_6466,N_6893);
nand U14053 (N_14053,N_7411,N_9783);
or U14054 (N_14054,N_8781,N_7261);
or U14055 (N_14055,N_6293,N_9468);
and U14056 (N_14056,N_5868,N_7198);
nor U14057 (N_14057,N_7847,N_6620);
nand U14058 (N_14058,N_6913,N_7039);
or U14059 (N_14059,N_5561,N_8965);
xnor U14060 (N_14060,N_6007,N_8354);
nand U14061 (N_14061,N_8364,N_5800);
xor U14062 (N_14062,N_9404,N_5929);
nor U14063 (N_14063,N_8197,N_8500);
or U14064 (N_14064,N_7047,N_6761);
or U14065 (N_14065,N_9549,N_5226);
or U14066 (N_14066,N_7700,N_6750);
nor U14067 (N_14067,N_5840,N_5294);
xor U14068 (N_14068,N_9173,N_7093);
nand U14069 (N_14069,N_9912,N_6442);
nor U14070 (N_14070,N_6957,N_7486);
or U14071 (N_14071,N_6944,N_8771);
xor U14072 (N_14072,N_8081,N_5231);
xor U14073 (N_14073,N_7954,N_9950);
nor U14074 (N_14074,N_5156,N_7150);
xnor U14075 (N_14075,N_8976,N_5115);
or U14076 (N_14076,N_6822,N_8294);
nand U14077 (N_14077,N_7242,N_9470);
or U14078 (N_14078,N_8337,N_7453);
and U14079 (N_14079,N_8261,N_7412);
nand U14080 (N_14080,N_7115,N_7943);
nor U14081 (N_14081,N_8656,N_6161);
nor U14082 (N_14082,N_9393,N_6719);
and U14083 (N_14083,N_8217,N_6670);
or U14084 (N_14084,N_8329,N_5633);
nor U14085 (N_14085,N_9573,N_5089);
and U14086 (N_14086,N_7238,N_9982);
nand U14087 (N_14087,N_8664,N_6722);
or U14088 (N_14088,N_8298,N_6826);
xor U14089 (N_14089,N_8530,N_9385);
nand U14090 (N_14090,N_5326,N_9941);
or U14091 (N_14091,N_5693,N_5778);
nand U14092 (N_14092,N_8352,N_5177);
or U14093 (N_14093,N_6465,N_9422);
nand U14094 (N_14094,N_7405,N_9593);
nand U14095 (N_14095,N_5692,N_9539);
nand U14096 (N_14096,N_5501,N_8305);
nor U14097 (N_14097,N_6595,N_5922);
nand U14098 (N_14098,N_9400,N_5411);
nand U14099 (N_14099,N_8778,N_8863);
nand U14100 (N_14100,N_7007,N_9664);
xor U14101 (N_14101,N_7505,N_5864);
or U14102 (N_14102,N_5627,N_8719);
nor U14103 (N_14103,N_9177,N_5033);
nand U14104 (N_14104,N_8135,N_7536);
nor U14105 (N_14105,N_6756,N_5893);
or U14106 (N_14106,N_9026,N_8170);
xnor U14107 (N_14107,N_5605,N_7771);
and U14108 (N_14108,N_9639,N_8624);
and U14109 (N_14109,N_9298,N_9569);
xnor U14110 (N_14110,N_5750,N_7937);
nor U14111 (N_14111,N_9827,N_5632);
xor U14112 (N_14112,N_7647,N_6026);
xor U14113 (N_14113,N_6498,N_9875);
nor U14114 (N_14114,N_9311,N_8964);
or U14115 (N_14115,N_8963,N_5381);
or U14116 (N_14116,N_9254,N_6191);
nand U14117 (N_14117,N_7281,N_9223);
xor U14118 (N_14118,N_6898,N_9792);
or U14119 (N_14119,N_8783,N_8631);
or U14120 (N_14120,N_7533,N_7445);
nor U14121 (N_14121,N_9181,N_9352);
and U14122 (N_14122,N_5615,N_8017);
or U14123 (N_14123,N_9750,N_7004);
nand U14124 (N_14124,N_8119,N_6096);
and U14125 (N_14125,N_9140,N_7460);
nor U14126 (N_14126,N_9017,N_6798);
nand U14127 (N_14127,N_8087,N_9036);
or U14128 (N_14128,N_6675,N_5182);
xor U14129 (N_14129,N_5236,N_5473);
nor U14130 (N_14130,N_6880,N_9497);
xnor U14131 (N_14131,N_9890,N_9619);
and U14132 (N_14132,N_9342,N_6709);
nor U14133 (N_14133,N_8061,N_8827);
xor U14134 (N_14134,N_9882,N_6310);
or U14135 (N_14135,N_6353,N_9287);
nor U14136 (N_14136,N_7763,N_7959);
and U14137 (N_14137,N_6787,N_9464);
or U14138 (N_14138,N_8424,N_6991);
xnor U14139 (N_14139,N_9421,N_9940);
and U14140 (N_14140,N_7234,N_9560);
xnor U14141 (N_14141,N_5942,N_6660);
or U14142 (N_14142,N_7570,N_5345);
or U14143 (N_14143,N_9897,N_9972);
nor U14144 (N_14144,N_8385,N_6111);
nand U14145 (N_14145,N_8465,N_5401);
nand U14146 (N_14146,N_9706,N_6297);
xor U14147 (N_14147,N_7018,N_6938);
or U14148 (N_14148,N_5158,N_5548);
nand U14149 (N_14149,N_6931,N_6549);
nand U14150 (N_14150,N_5088,N_5526);
or U14151 (N_14151,N_5971,N_7342);
xor U14152 (N_14152,N_6218,N_5690);
and U14153 (N_14153,N_8521,N_7951);
xnor U14154 (N_14154,N_7947,N_7043);
or U14155 (N_14155,N_7019,N_5400);
xnor U14156 (N_14156,N_5343,N_9210);
nor U14157 (N_14157,N_7472,N_9212);
or U14158 (N_14158,N_5713,N_6724);
nand U14159 (N_14159,N_5090,N_7298);
and U14160 (N_14160,N_5736,N_6777);
nand U14161 (N_14161,N_7909,N_5181);
xnor U14162 (N_14162,N_6125,N_9835);
nor U14163 (N_14163,N_8188,N_9490);
or U14164 (N_14164,N_9071,N_5618);
nand U14165 (N_14165,N_5392,N_8602);
or U14166 (N_14166,N_5466,N_8463);
nand U14167 (N_14167,N_9124,N_7568);
xor U14168 (N_14168,N_9001,N_7266);
xnor U14169 (N_14169,N_5561,N_9060);
nand U14170 (N_14170,N_8043,N_6809);
nor U14171 (N_14171,N_6964,N_9299);
nor U14172 (N_14172,N_5763,N_7074);
xnor U14173 (N_14173,N_6647,N_8812);
xnor U14174 (N_14174,N_8931,N_9538);
and U14175 (N_14175,N_8298,N_8840);
and U14176 (N_14176,N_6889,N_8597);
and U14177 (N_14177,N_8651,N_7198);
xor U14178 (N_14178,N_6318,N_6127);
nand U14179 (N_14179,N_9748,N_5952);
nand U14180 (N_14180,N_6225,N_8708);
xor U14181 (N_14181,N_6498,N_5227);
or U14182 (N_14182,N_8828,N_7055);
and U14183 (N_14183,N_9312,N_5684);
xnor U14184 (N_14184,N_8310,N_7967);
xor U14185 (N_14185,N_5626,N_8277);
xor U14186 (N_14186,N_7261,N_7820);
or U14187 (N_14187,N_9257,N_5350);
nor U14188 (N_14188,N_8216,N_5466);
and U14189 (N_14189,N_7554,N_8737);
xor U14190 (N_14190,N_6751,N_7584);
and U14191 (N_14191,N_8361,N_6957);
nand U14192 (N_14192,N_8279,N_8883);
or U14193 (N_14193,N_6649,N_6831);
xnor U14194 (N_14194,N_5437,N_7567);
nand U14195 (N_14195,N_6372,N_7048);
xnor U14196 (N_14196,N_6914,N_8346);
nor U14197 (N_14197,N_6535,N_7612);
xor U14198 (N_14198,N_5636,N_7466);
or U14199 (N_14199,N_9920,N_5861);
nand U14200 (N_14200,N_6478,N_7799);
nor U14201 (N_14201,N_9318,N_7924);
and U14202 (N_14202,N_8984,N_7827);
and U14203 (N_14203,N_7804,N_6920);
and U14204 (N_14204,N_7056,N_9427);
and U14205 (N_14205,N_6365,N_9816);
xor U14206 (N_14206,N_9185,N_7347);
or U14207 (N_14207,N_6427,N_6155);
and U14208 (N_14208,N_6223,N_9685);
xnor U14209 (N_14209,N_6210,N_6320);
or U14210 (N_14210,N_7830,N_7888);
nor U14211 (N_14211,N_5193,N_7417);
and U14212 (N_14212,N_7561,N_7743);
or U14213 (N_14213,N_7935,N_8568);
nand U14214 (N_14214,N_6233,N_9090);
or U14215 (N_14215,N_8886,N_6952);
xor U14216 (N_14216,N_9910,N_9874);
nor U14217 (N_14217,N_5933,N_8333);
xor U14218 (N_14218,N_8289,N_8659);
xor U14219 (N_14219,N_7322,N_5450);
xor U14220 (N_14220,N_5931,N_6697);
xor U14221 (N_14221,N_5803,N_6465);
nor U14222 (N_14222,N_5304,N_8481);
and U14223 (N_14223,N_8716,N_8797);
and U14224 (N_14224,N_5600,N_6603);
or U14225 (N_14225,N_6151,N_7319);
and U14226 (N_14226,N_6665,N_7300);
nand U14227 (N_14227,N_9722,N_6825);
nand U14228 (N_14228,N_7814,N_5347);
nor U14229 (N_14229,N_5045,N_9903);
nor U14230 (N_14230,N_8111,N_5523);
nor U14231 (N_14231,N_6134,N_8216);
xnor U14232 (N_14232,N_7145,N_9034);
and U14233 (N_14233,N_5290,N_8374);
and U14234 (N_14234,N_8030,N_7792);
nand U14235 (N_14235,N_9417,N_9542);
nor U14236 (N_14236,N_5633,N_7542);
nor U14237 (N_14237,N_7189,N_7201);
or U14238 (N_14238,N_6613,N_8705);
and U14239 (N_14239,N_9058,N_5075);
or U14240 (N_14240,N_7677,N_5235);
and U14241 (N_14241,N_5205,N_5397);
xnor U14242 (N_14242,N_5329,N_7186);
nor U14243 (N_14243,N_9270,N_9714);
nor U14244 (N_14244,N_6222,N_6113);
and U14245 (N_14245,N_9473,N_6867);
or U14246 (N_14246,N_9289,N_5664);
nor U14247 (N_14247,N_9717,N_7456);
and U14248 (N_14248,N_6016,N_7341);
nand U14249 (N_14249,N_5332,N_6249);
xnor U14250 (N_14250,N_6885,N_9867);
and U14251 (N_14251,N_8982,N_7466);
and U14252 (N_14252,N_6861,N_9651);
xnor U14253 (N_14253,N_8982,N_9643);
nand U14254 (N_14254,N_9667,N_7041);
nand U14255 (N_14255,N_5319,N_8981);
or U14256 (N_14256,N_9447,N_6126);
xor U14257 (N_14257,N_5835,N_5001);
xnor U14258 (N_14258,N_8875,N_7215);
and U14259 (N_14259,N_7127,N_6161);
xnor U14260 (N_14260,N_8956,N_5164);
nor U14261 (N_14261,N_5085,N_6274);
or U14262 (N_14262,N_7154,N_7574);
nand U14263 (N_14263,N_5628,N_6160);
nand U14264 (N_14264,N_8974,N_9769);
and U14265 (N_14265,N_8254,N_6303);
or U14266 (N_14266,N_6987,N_5114);
xor U14267 (N_14267,N_5245,N_8028);
or U14268 (N_14268,N_7183,N_5587);
nand U14269 (N_14269,N_9186,N_7785);
xor U14270 (N_14270,N_7148,N_8930);
nand U14271 (N_14271,N_7719,N_6560);
or U14272 (N_14272,N_8166,N_9615);
nor U14273 (N_14273,N_6141,N_5342);
or U14274 (N_14274,N_8489,N_9476);
nand U14275 (N_14275,N_9872,N_7525);
nor U14276 (N_14276,N_8344,N_9138);
xor U14277 (N_14277,N_5429,N_9815);
xor U14278 (N_14278,N_8685,N_7312);
and U14279 (N_14279,N_7875,N_9536);
nand U14280 (N_14280,N_5878,N_9911);
and U14281 (N_14281,N_7307,N_9340);
nand U14282 (N_14282,N_7165,N_9214);
and U14283 (N_14283,N_5333,N_6283);
xor U14284 (N_14284,N_8390,N_5089);
xnor U14285 (N_14285,N_5786,N_5297);
xnor U14286 (N_14286,N_8190,N_9777);
or U14287 (N_14287,N_9036,N_7591);
xnor U14288 (N_14288,N_8066,N_7796);
and U14289 (N_14289,N_8837,N_8993);
xor U14290 (N_14290,N_8236,N_9217);
xor U14291 (N_14291,N_8148,N_6303);
or U14292 (N_14292,N_8750,N_9332);
nand U14293 (N_14293,N_8444,N_6291);
or U14294 (N_14294,N_5567,N_7992);
or U14295 (N_14295,N_8676,N_6284);
nor U14296 (N_14296,N_8992,N_7756);
or U14297 (N_14297,N_5207,N_9175);
nor U14298 (N_14298,N_9820,N_5871);
and U14299 (N_14299,N_6485,N_6304);
nor U14300 (N_14300,N_6778,N_8885);
nand U14301 (N_14301,N_5001,N_5280);
and U14302 (N_14302,N_8617,N_5427);
or U14303 (N_14303,N_7073,N_8896);
and U14304 (N_14304,N_8212,N_5625);
nor U14305 (N_14305,N_9353,N_9196);
xnor U14306 (N_14306,N_5644,N_6562);
and U14307 (N_14307,N_6021,N_5197);
xor U14308 (N_14308,N_9594,N_9643);
nor U14309 (N_14309,N_9028,N_9105);
or U14310 (N_14310,N_6899,N_8182);
or U14311 (N_14311,N_9784,N_9649);
xor U14312 (N_14312,N_9265,N_5353);
nand U14313 (N_14313,N_9528,N_5651);
xnor U14314 (N_14314,N_9377,N_6096);
nor U14315 (N_14315,N_8923,N_9272);
and U14316 (N_14316,N_8246,N_5603);
and U14317 (N_14317,N_5865,N_6029);
nand U14318 (N_14318,N_9910,N_9576);
and U14319 (N_14319,N_8459,N_6223);
xnor U14320 (N_14320,N_7570,N_7031);
xor U14321 (N_14321,N_8362,N_7260);
or U14322 (N_14322,N_8236,N_6466);
xnor U14323 (N_14323,N_7686,N_8141);
xnor U14324 (N_14324,N_5661,N_9521);
nand U14325 (N_14325,N_6020,N_8491);
and U14326 (N_14326,N_9251,N_5252);
or U14327 (N_14327,N_8293,N_9143);
and U14328 (N_14328,N_8257,N_5482);
nor U14329 (N_14329,N_8971,N_9907);
nand U14330 (N_14330,N_8654,N_5021);
and U14331 (N_14331,N_8145,N_7143);
nor U14332 (N_14332,N_6399,N_7652);
nor U14333 (N_14333,N_8171,N_7925);
nor U14334 (N_14334,N_6880,N_7441);
or U14335 (N_14335,N_9816,N_8443);
nand U14336 (N_14336,N_9494,N_8899);
and U14337 (N_14337,N_8209,N_9304);
xor U14338 (N_14338,N_5699,N_9217);
xor U14339 (N_14339,N_9319,N_9246);
nor U14340 (N_14340,N_9060,N_8624);
and U14341 (N_14341,N_9640,N_6440);
nand U14342 (N_14342,N_6061,N_6172);
xor U14343 (N_14343,N_5605,N_8068);
nor U14344 (N_14344,N_6423,N_5544);
or U14345 (N_14345,N_5984,N_5691);
or U14346 (N_14346,N_5514,N_5201);
or U14347 (N_14347,N_5523,N_8692);
and U14348 (N_14348,N_6573,N_6729);
nor U14349 (N_14349,N_5279,N_8649);
or U14350 (N_14350,N_9967,N_5758);
nand U14351 (N_14351,N_8564,N_8088);
and U14352 (N_14352,N_5134,N_7539);
or U14353 (N_14353,N_6255,N_5199);
nand U14354 (N_14354,N_5222,N_5944);
nand U14355 (N_14355,N_8796,N_9736);
nand U14356 (N_14356,N_5388,N_6394);
nand U14357 (N_14357,N_6201,N_7989);
and U14358 (N_14358,N_8250,N_9134);
xor U14359 (N_14359,N_7554,N_6424);
nand U14360 (N_14360,N_9723,N_8953);
nand U14361 (N_14361,N_6453,N_8170);
or U14362 (N_14362,N_8555,N_5319);
and U14363 (N_14363,N_7613,N_7908);
and U14364 (N_14364,N_8633,N_6835);
or U14365 (N_14365,N_6707,N_6552);
or U14366 (N_14366,N_8419,N_6015);
nor U14367 (N_14367,N_9708,N_6225);
nand U14368 (N_14368,N_7997,N_8587);
xor U14369 (N_14369,N_6874,N_6847);
nand U14370 (N_14370,N_8552,N_7836);
nand U14371 (N_14371,N_6109,N_8154);
or U14372 (N_14372,N_6015,N_9329);
nand U14373 (N_14373,N_8570,N_6010);
or U14374 (N_14374,N_8775,N_7348);
and U14375 (N_14375,N_9478,N_7151);
xor U14376 (N_14376,N_8862,N_8174);
xor U14377 (N_14377,N_5028,N_5569);
and U14378 (N_14378,N_7058,N_5159);
or U14379 (N_14379,N_5223,N_8605);
or U14380 (N_14380,N_9518,N_8576);
nand U14381 (N_14381,N_7419,N_9356);
or U14382 (N_14382,N_5521,N_5926);
xnor U14383 (N_14383,N_8291,N_7646);
and U14384 (N_14384,N_9340,N_6760);
nand U14385 (N_14385,N_5895,N_6664);
nor U14386 (N_14386,N_5216,N_6574);
xor U14387 (N_14387,N_5051,N_5647);
xor U14388 (N_14388,N_5716,N_5102);
or U14389 (N_14389,N_9182,N_5850);
nor U14390 (N_14390,N_7361,N_8419);
or U14391 (N_14391,N_5241,N_7046);
and U14392 (N_14392,N_7903,N_7568);
or U14393 (N_14393,N_5974,N_6254);
and U14394 (N_14394,N_6752,N_9556);
and U14395 (N_14395,N_8115,N_6595);
nor U14396 (N_14396,N_9534,N_6446);
xnor U14397 (N_14397,N_9515,N_6888);
xnor U14398 (N_14398,N_8550,N_8333);
and U14399 (N_14399,N_8382,N_7699);
xor U14400 (N_14400,N_6302,N_5604);
nand U14401 (N_14401,N_8620,N_5918);
nor U14402 (N_14402,N_7529,N_5209);
xor U14403 (N_14403,N_9064,N_8829);
and U14404 (N_14404,N_8271,N_8306);
or U14405 (N_14405,N_5763,N_5994);
or U14406 (N_14406,N_5282,N_6636);
xnor U14407 (N_14407,N_6070,N_8599);
and U14408 (N_14408,N_9367,N_9979);
nand U14409 (N_14409,N_7525,N_5366);
nor U14410 (N_14410,N_7468,N_8944);
nor U14411 (N_14411,N_9247,N_5413);
and U14412 (N_14412,N_6657,N_5744);
and U14413 (N_14413,N_5121,N_5251);
and U14414 (N_14414,N_7859,N_6393);
and U14415 (N_14415,N_8809,N_5751);
xnor U14416 (N_14416,N_8188,N_9357);
xnor U14417 (N_14417,N_9359,N_7516);
nand U14418 (N_14418,N_7211,N_7597);
nand U14419 (N_14419,N_9878,N_6789);
nor U14420 (N_14420,N_6032,N_9634);
or U14421 (N_14421,N_8559,N_8921);
nor U14422 (N_14422,N_5252,N_5287);
nor U14423 (N_14423,N_6152,N_9762);
or U14424 (N_14424,N_8485,N_6383);
nand U14425 (N_14425,N_9859,N_7383);
nor U14426 (N_14426,N_5942,N_5195);
nor U14427 (N_14427,N_6202,N_9327);
xor U14428 (N_14428,N_8944,N_9745);
and U14429 (N_14429,N_6485,N_7706);
nor U14430 (N_14430,N_9933,N_9180);
or U14431 (N_14431,N_7908,N_5324);
or U14432 (N_14432,N_8114,N_7903);
and U14433 (N_14433,N_5314,N_7461);
nor U14434 (N_14434,N_6243,N_8459);
and U14435 (N_14435,N_6179,N_9654);
and U14436 (N_14436,N_7979,N_7791);
and U14437 (N_14437,N_6262,N_9948);
nor U14438 (N_14438,N_6181,N_8143);
nor U14439 (N_14439,N_9822,N_7050);
xor U14440 (N_14440,N_5160,N_9490);
nand U14441 (N_14441,N_8147,N_6223);
or U14442 (N_14442,N_5131,N_6056);
and U14443 (N_14443,N_6301,N_9867);
or U14444 (N_14444,N_9689,N_8564);
or U14445 (N_14445,N_7622,N_7235);
and U14446 (N_14446,N_8798,N_9976);
nand U14447 (N_14447,N_7002,N_8715);
nor U14448 (N_14448,N_5148,N_7717);
and U14449 (N_14449,N_6997,N_9881);
nor U14450 (N_14450,N_8192,N_6859);
nor U14451 (N_14451,N_7622,N_7608);
or U14452 (N_14452,N_6646,N_6370);
nand U14453 (N_14453,N_9744,N_5709);
nor U14454 (N_14454,N_5408,N_5739);
nand U14455 (N_14455,N_5612,N_8329);
and U14456 (N_14456,N_7692,N_7767);
and U14457 (N_14457,N_6232,N_8429);
nor U14458 (N_14458,N_8064,N_8924);
and U14459 (N_14459,N_8141,N_6207);
nand U14460 (N_14460,N_7089,N_9625);
or U14461 (N_14461,N_7268,N_5090);
xnor U14462 (N_14462,N_5920,N_5072);
and U14463 (N_14463,N_8047,N_8628);
and U14464 (N_14464,N_8547,N_5271);
and U14465 (N_14465,N_7801,N_7523);
nand U14466 (N_14466,N_6898,N_9472);
or U14467 (N_14467,N_6043,N_9297);
and U14468 (N_14468,N_5530,N_9728);
nand U14469 (N_14469,N_5076,N_9413);
xor U14470 (N_14470,N_5028,N_7746);
and U14471 (N_14471,N_7224,N_6205);
and U14472 (N_14472,N_8020,N_5095);
and U14473 (N_14473,N_5354,N_8484);
or U14474 (N_14474,N_8060,N_8647);
and U14475 (N_14475,N_6636,N_7372);
nor U14476 (N_14476,N_8214,N_6755);
or U14477 (N_14477,N_9942,N_5550);
nor U14478 (N_14478,N_8905,N_7026);
or U14479 (N_14479,N_8224,N_9853);
nand U14480 (N_14480,N_7259,N_8333);
or U14481 (N_14481,N_5468,N_9180);
xor U14482 (N_14482,N_6132,N_7408);
nor U14483 (N_14483,N_6760,N_9718);
xor U14484 (N_14484,N_8087,N_9246);
and U14485 (N_14485,N_6461,N_9550);
xnor U14486 (N_14486,N_6439,N_9136);
nand U14487 (N_14487,N_8840,N_7953);
or U14488 (N_14488,N_8102,N_8464);
xor U14489 (N_14489,N_8651,N_6962);
xor U14490 (N_14490,N_8635,N_7443);
xnor U14491 (N_14491,N_5739,N_9193);
xnor U14492 (N_14492,N_6673,N_6272);
or U14493 (N_14493,N_6481,N_6235);
nor U14494 (N_14494,N_9930,N_6233);
or U14495 (N_14495,N_5742,N_7033);
nand U14496 (N_14496,N_9839,N_7673);
and U14497 (N_14497,N_7814,N_8906);
and U14498 (N_14498,N_8051,N_6988);
xnor U14499 (N_14499,N_8389,N_8687);
and U14500 (N_14500,N_8381,N_7339);
or U14501 (N_14501,N_8286,N_9352);
nor U14502 (N_14502,N_7591,N_7924);
or U14503 (N_14503,N_8181,N_9977);
nand U14504 (N_14504,N_8133,N_9685);
and U14505 (N_14505,N_5298,N_9419);
or U14506 (N_14506,N_8407,N_7738);
nor U14507 (N_14507,N_8966,N_6701);
xnor U14508 (N_14508,N_7745,N_6370);
or U14509 (N_14509,N_8390,N_9502);
xor U14510 (N_14510,N_6510,N_9238);
xnor U14511 (N_14511,N_7064,N_9606);
and U14512 (N_14512,N_6565,N_7674);
and U14513 (N_14513,N_8961,N_9900);
or U14514 (N_14514,N_5432,N_7203);
and U14515 (N_14515,N_8636,N_5332);
nand U14516 (N_14516,N_5885,N_5966);
xor U14517 (N_14517,N_6061,N_8882);
nor U14518 (N_14518,N_8267,N_8150);
or U14519 (N_14519,N_5590,N_8190);
or U14520 (N_14520,N_6922,N_9971);
or U14521 (N_14521,N_7013,N_7722);
xnor U14522 (N_14522,N_8248,N_9057);
or U14523 (N_14523,N_5006,N_6781);
xnor U14524 (N_14524,N_5287,N_5593);
or U14525 (N_14525,N_6754,N_5690);
and U14526 (N_14526,N_7718,N_9498);
nand U14527 (N_14527,N_7273,N_6212);
or U14528 (N_14528,N_5969,N_8698);
nand U14529 (N_14529,N_9703,N_5404);
and U14530 (N_14530,N_6572,N_7613);
or U14531 (N_14531,N_5181,N_9475);
and U14532 (N_14532,N_8389,N_8101);
nor U14533 (N_14533,N_5057,N_9420);
and U14534 (N_14534,N_6451,N_6374);
or U14535 (N_14535,N_5316,N_7992);
and U14536 (N_14536,N_9293,N_7889);
nor U14537 (N_14537,N_6236,N_5395);
nand U14538 (N_14538,N_5585,N_9422);
nand U14539 (N_14539,N_5692,N_6713);
or U14540 (N_14540,N_6276,N_6104);
nand U14541 (N_14541,N_9106,N_9533);
and U14542 (N_14542,N_7669,N_8200);
xor U14543 (N_14543,N_8990,N_8921);
xor U14544 (N_14544,N_5619,N_9202);
xnor U14545 (N_14545,N_6175,N_8506);
nor U14546 (N_14546,N_6091,N_8791);
and U14547 (N_14547,N_5408,N_5875);
nor U14548 (N_14548,N_7622,N_7702);
nor U14549 (N_14549,N_5811,N_8375);
and U14550 (N_14550,N_8731,N_6345);
or U14551 (N_14551,N_8072,N_7957);
nand U14552 (N_14552,N_7604,N_6934);
nor U14553 (N_14553,N_7699,N_7964);
xor U14554 (N_14554,N_6093,N_6532);
or U14555 (N_14555,N_6630,N_6192);
nand U14556 (N_14556,N_7050,N_6230);
xnor U14557 (N_14557,N_7456,N_5028);
or U14558 (N_14558,N_6566,N_9323);
nand U14559 (N_14559,N_8845,N_5965);
or U14560 (N_14560,N_8577,N_7532);
and U14561 (N_14561,N_6228,N_6874);
nor U14562 (N_14562,N_7574,N_7215);
nand U14563 (N_14563,N_7381,N_5707);
nor U14564 (N_14564,N_8657,N_9114);
nor U14565 (N_14565,N_8294,N_6191);
xnor U14566 (N_14566,N_6848,N_5989);
nor U14567 (N_14567,N_7523,N_9525);
and U14568 (N_14568,N_9896,N_6048);
nand U14569 (N_14569,N_5459,N_8691);
xor U14570 (N_14570,N_6086,N_8210);
and U14571 (N_14571,N_5894,N_5279);
and U14572 (N_14572,N_8010,N_8398);
or U14573 (N_14573,N_9943,N_5105);
or U14574 (N_14574,N_8798,N_9479);
xnor U14575 (N_14575,N_5071,N_8364);
nor U14576 (N_14576,N_6156,N_6852);
nor U14577 (N_14577,N_9939,N_9376);
nor U14578 (N_14578,N_9775,N_6025);
or U14579 (N_14579,N_7599,N_5855);
xor U14580 (N_14580,N_6734,N_5912);
xnor U14581 (N_14581,N_6303,N_9271);
nor U14582 (N_14582,N_7621,N_8971);
nand U14583 (N_14583,N_6199,N_5018);
and U14584 (N_14584,N_6505,N_6288);
or U14585 (N_14585,N_8171,N_5836);
xnor U14586 (N_14586,N_8134,N_8580);
nor U14587 (N_14587,N_6112,N_7513);
or U14588 (N_14588,N_8121,N_6887);
nor U14589 (N_14589,N_8425,N_6532);
and U14590 (N_14590,N_7199,N_8221);
xnor U14591 (N_14591,N_6387,N_9257);
nand U14592 (N_14592,N_5060,N_9802);
xor U14593 (N_14593,N_5462,N_6896);
or U14594 (N_14594,N_7818,N_8862);
nor U14595 (N_14595,N_7522,N_6455);
nand U14596 (N_14596,N_7238,N_7683);
nand U14597 (N_14597,N_7419,N_9753);
nand U14598 (N_14598,N_8597,N_7958);
or U14599 (N_14599,N_5229,N_6020);
or U14600 (N_14600,N_5012,N_9484);
xnor U14601 (N_14601,N_6656,N_5372);
and U14602 (N_14602,N_6921,N_6266);
or U14603 (N_14603,N_7826,N_5559);
nand U14604 (N_14604,N_5831,N_8062);
or U14605 (N_14605,N_6841,N_5820);
and U14606 (N_14606,N_9375,N_5390);
or U14607 (N_14607,N_7366,N_7099);
nand U14608 (N_14608,N_7547,N_9140);
nor U14609 (N_14609,N_9768,N_7309);
or U14610 (N_14610,N_7219,N_6361);
xor U14611 (N_14611,N_8738,N_9695);
nand U14612 (N_14612,N_5984,N_5353);
nand U14613 (N_14613,N_5847,N_7826);
nor U14614 (N_14614,N_7317,N_9473);
nor U14615 (N_14615,N_5108,N_8311);
or U14616 (N_14616,N_5802,N_7515);
nor U14617 (N_14617,N_5393,N_9174);
nand U14618 (N_14618,N_5301,N_7592);
nand U14619 (N_14619,N_7588,N_6536);
xor U14620 (N_14620,N_7904,N_6279);
nor U14621 (N_14621,N_7973,N_8970);
xnor U14622 (N_14622,N_8175,N_7663);
or U14623 (N_14623,N_6256,N_9852);
nand U14624 (N_14624,N_6015,N_5690);
xor U14625 (N_14625,N_7260,N_9110);
and U14626 (N_14626,N_7717,N_8459);
nand U14627 (N_14627,N_9186,N_7755);
or U14628 (N_14628,N_5296,N_7768);
nor U14629 (N_14629,N_7328,N_7857);
nor U14630 (N_14630,N_9377,N_5041);
or U14631 (N_14631,N_6945,N_6461);
and U14632 (N_14632,N_9687,N_9026);
nand U14633 (N_14633,N_8232,N_6985);
nand U14634 (N_14634,N_7309,N_9304);
xnor U14635 (N_14635,N_6077,N_7178);
or U14636 (N_14636,N_5956,N_7487);
nand U14637 (N_14637,N_9895,N_7964);
nand U14638 (N_14638,N_9343,N_7538);
nand U14639 (N_14639,N_6710,N_5512);
or U14640 (N_14640,N_7119,N_5708);
nor U14641 (N_14641,N_5459,N_9499);
nor U14642 (N_14642,N_6903,N_8187);
and U14643 (N_14643,N_8402,N_7564);
nor U14644 (N_14644,N_7902,N_7722);
xnor U14645 (N_14645,N_6502,N_9797);
nand U14646 (N_14646,N_7124,N_9140);
or U14647 (N_14647,N_7718,N_5256);
xor U14648 (N_14648,N_8887,N_6582);
nand U14649 (N_14649,N_9197,N_5734);
nor U14650 (N_14650,N_7421,N_9800);
nor U14651 (N_14651,N_6094,N_6117);
and U14652 (N_14652,N_6062,N_9209);
or U14653 (N_14653,N_7875,N_9981);
nand U14654 (N_14654,N_8907,N_7664);
and U14655 (N_14655,N_8242,N_6905);
nand U14656 (N_14656,N_8341,N_7906);
and U14657 (N_14657,N_7446,N_5529);
and U14658 (N_14658,N_5831,N_6854);
and U14659 (N_14659,N_9381,N_7424);
or U14660 (N_14660,N_9444,N_8855);
xnor U14661 (N_14661,N_6037,N_5915);
xor U14662 (N_14662,N_8883,N_5537);
nand U14663 (N_14663,N_9534,N_8269);
nand U14664 (N_14664,N_8304,N_5490);
and U14665 (N_14665,N_8656,N_7779);
xnor U14666 (N_14666,N_8551,N_8142);
and U14667 (N_14667,N_7695,N_5486);
and U14668 (N_14668,N_6811,N_5948);
and U14669 (N_14669,N_9008,N_8459);
xnor U14670 (N_14670,N_8456,N_5187);
xnor U14671 (N_14671,N_6209,N_6287);
nand U14672 (N_14672,N_5532,N_8288);
or U14673 (N_14673,N_5646,N_7800);
nand U14674 (N_14674,N_9848,N_8369);
nand U14675 (N_14675,N_5783,N_6523);
xnor U14676 (N_14676,N_6853,N_6438);
nand U14677 (N_14677,N_7206,N_6272);
nand U14678 (N_14678,N_7819,N_9347);
nor U14679 (N_14679,N_7180,N_7621);
nand U14680 (N_14680,N_9528,N_8413);
xor U14681 (N_14681,N_7223,N_6319);
nor U14682 (N_14682,N_8934,N_5562);
or U14683 (N_14683,N_6639,N_9518);
or U14684 (N_14684,N_6519,N_6014);
or U14685 (N_14685,N_5476,N_9135);
and U14686 (N_14686,N_7885,N_5138);
nor U14687 (N_14687,N_6826,N_5827);
xnor U14688 (N_14688,N_9839,N_5187);
and U14689 (N_14689,N_5695,N_9682);
nor U14690 (N_14690,N_8794,N_7858);
nand U14691 (N_14691,N_7935,N_5676);
and U14692 (N_14692,N_8217,N_5657);
xor U14693 (N_14693,N_5260,N_6424);
nand U14694 (N_14694,N_8950,N_8649);
or U14695 (N_14695,N_5417,N_9861);
and U14696 (N_14696,N_7881,N_7130);
xor U14697 (N_14697,N_9433,N_5003);
or U14698 (N_14698,N_8623,N_9831);
and U14699 (N_14699,N_8970,N_5849);
nor U14700 (N_14700,N_5153,N_7502);
nor U14701 (N_14701,N_9848,N_6702);
nand U14702 (N_14702,N_6361,N_8276);
xor U14703 (N_14703,N_9922,N_6863);
and U14704 (N_14704,N_8451,N_5210);
nor U14705 (N_14705,N_7431,N_7995);
and U14706 (N_14706,N_7410,N_7210);
nand U14707 (N_14707,N_7969,N_9246);
nor U14708 (N_14708,N_9411,N_9309);
or U14709 (N_14709,N_9128,N_9209);
and U14710 (N_14710,N_6432,N_6372);
or U14711 (N_14711,N_9799,N_5446);
and U14712 (N_14712,N_8816,N_6210);
and U14713 (N_14713,N_8396,N_8036);
nand U14714 (N_14714,N_5557,N_9769);
xnor U14715 (N_14715,N_7013,N_8361);
xor U14716 (N_14716,N_6081,N_9313);
and U14717 (N_14717,N_8285,N_9194);
nand U14718 (N_14718,N_8711,N_9896);
nand U14719 (N_14719,N_8667,N_8780);
nor U14720 (N_14720,N_9448,N_9115);
or U14721 (N_14721,N_5621,N_8695);
xnor U14722 (N_14722,N_9783,N_5280);
nor U14723 (N_14723,N_9471,N_7650);
nor U14724 (N_14724,N_5381,N_7257);
or U14725 (N_14725,N_7923,N_8760);
and U14726 (N_14726,N_5431,N_9649);
nand U14727 (N_14727,N_5819,N_7662);
xnor U14728 (N_14728,N_7799,N_5833);
or U14729 (N_14729,N_6684,N_5876);
and U14730 (N_14730,N_9655,N_9324);
or U14731 (N_14731,N_8397,N_5745);
xor U14732 (N_14732,N_7877,N_8007);
or U14733 (N_14733,N_8212,N_9284);
and U14734 (N_14734,N_8543,N_5384);
or U14735 (N_14735,N_9722,N_9618);
or U14736 (N_14736,N_6991,N_7557);
or U14737 (N_14737,N_9139,N_5036);
or U14738 (N_14738,N_7996,N_6351);
nor U14739 (N_14739,N_5256,N_6534);
xor U14740 (N_14740,N_7083,N_8872);
and U14741 (N_14741,N_9881,N_9468);
nand U14742 (N_14742,N_8459,N_5390);
or U14743 (N_14743,N_6412,N_9310);
nor U14744 (N_14744,N_6964,N_7963);
xnor U14745 (N_14745,N_6957,N_8217);
xor U14746 (N_14746,N_6997,N_5564);
nand U14747 (N_14747,N_6369,N_6333);
or U14748 (N_14748,N_5390,N_8760);
and U14749 (N_14749,N_9009,N_7455);
nor U14750 (N_14750,N_8365,N_9576);
nor U14751 (N_14751,N_6876,N_7019);
or U14752 (N_14752,N_9225,N_8179);
xnor U14753 (N_14753,N_7468,N_7400);
nand U14754 (N_14754,N_7998,N_8690);
nand U14755 (N_14755,N_9869,N_8119);
xor U14756 (N_14756,N_5204,N_6665);
nor U14757 (N_14757,N_8241,N_6894);
or U14758 (N_14758,N_8432,N_8827);
xnor U14759 (N_14759,N_7058,N_8752);
nand U14760 (N_14760,N_7239,N_9621);
or U14761 (N_14761,N_9591,N_8478);
nor U14762 (N_14762,N_5464,N_7382);
nor U14763 (N_14763,N_6053,N_6041);
and U14764 (N_14764,N_9337,N_7494);
and U14765 (N_14765,N_9203,N_7428);
and U14766 (N_14766,N_6168,N_9034);
xor U14767 (N_14767,N_6320,N_8288);
nand U14768 (N_14768,N_6135,N_8386);
or U14769 (N_14769,N_5211,N_5787);
nand U14770 (N_14770,N_7184,N_9631);
xnor U14771 (N_14771,N_5569,N_9545);
and U14772 (N_14772,N_6441,N_5961);
or U14773 (N_14773,N_6082,N_8549);
or U14774 (N_14774,N_9039,N_8945);
nor U14775 (N_14775,N_7204,N_5570);
or U14776 (N_14776,N_6630,N_8064);
xor U14777 (N_14777,N_6230,N_6278);
or U14778 (N_14778,N_6324,N_6618);
and U14779 (N_14779,N_7990,N_9959);
nand U14780 (N_14780,N_9002,N_6443);
nor U14781 (N_14781,N_9537,N_8403);
nand U14782 (N_14782,N_8254,N_7519);
nand U14783 (N_14783,N_5740,N_9914);
or U14784 (N_14784,N_8705,N_6452);
and U14785 (N_14785,N_5431,N_8013);
or U14786 (N_14786,N_6320,N_8512);
xor U14787 (N_14787,N_7569,N_8301);
and U14788 (N_14788,N_5941,N_9282);
and U14789 (N_14789,N_7279,N_7803);
or U14790 (N_14790,N_7484,N_5437);
nor U14791 (N_14791,N_6942,N_9552);
nand U14792 (N_14792,N_6462,N_8698);
and U14793 (N_14793,N_6413,N_6202);
xor U14794 (N_14794,N_8683,N_7436);
and U14795 (N_14795,N_9972,N_9842);
or U14796 (N_14796,N_8335,N_8234);
nand U14797 (N_14797,N_7039,N_5035);
xor U14798 (N_14798,N_9928,N_5017);
xor U14799 (N_14799,N_9941,N_8922);
xnor U14800 (N_14800,N_8431,N_9601);
or U14801 (N_14801,N_8740,N_5281);
or U14802 (N_14802,N_8613,N_5873);
nand U14803 (N_14803,N_8202,N_8220);
nor U14804 (N_14804,N_6863,N_9647);
or U14805 (N_14805,N_7612,N_6105);
and U14806 (N_14806,N_8344,N_7088);
nand U14807 (N_14807,N_9045,N_9967);
and U14808 (N_14808,N_6390,N_9938);
nor U14809 (N_14809,N_5860,N_9593);
nor U14810 (N_14810,N_9142,N_7288);
nand U14811 (N_14811,N_7216,N_6352);
xor U14812 (N_14812,N_5411,N_8090);
and U14813 (N_14813,N_5014,N_5815);
nor U14814 (N_14814,N_9576,N_9964);
and U14815 (N_14815,N_9359,N_7214);
nor U14816 (N_14816,N_8261,N_6342);
nor U14817 (N_14817,N_7649,N_8609);
nand U14818 (N_14818,N_9991,N_6052);
nor U14819 (N_14819,N_6524,N_8917);
or U14820 (N_14820,N_5519,N_9000);
xnor U14821 (N_14821,N_8499,N_5744);
or U14822 (N_14822,N_7641,N_9137);
xnor U14823 (N_14823,N_7242,N_6933);
and U14824 (N_14824,N_8125,N_7100);
nand U14825 (N_14825,N_6125,N_8095);
nor U14826 (N_14826,N_6026,N_9431);
nor U14827 (N_14827,N_9591,N_8472);
and U14828 (N_14828,N_8447,N_9278);
nand U14829 (N_14829,N_5628,N_6320);
xnor U14830 (N_14830,N_7707,N_9124);
xor U14831 (N_14831,N_5859,N_9255);
xor U14832 (N_14832,N_7156,N_8252);
xnor U14833 (N_14833,N_8749,N_9147);
xnor U14834 (N_14834,N_6433,N_8917);
and U14835 (N_14835,N_6239,N_5711);
nand U14836 (N_14836,N_8697,N_9890);
xor U14837 (N_14837,N_8356,N_6234);
or U14838 (N_14838,N_9847,N_9838);
nand U14839 (N_14839,N_6569,N_7910);
nand U14840 (N_14840,N_7884,N_5978);
or U14841 (N_14841,N_5508,N_6365);
xnor U14842 (N_14842,N_7927,N_9960);
and U14843 (N_14843,N_8095,N_6447);
xnor U14844 (N_14844,N_6948,N_7555);
nor U14845 (N_14845,N_5828,N_6419);
nand U14846 (N_14846,N_5748,N_7934);
xor U14847 (N_14847,N_7609,N_9087);
nand U14848 (N_14848,N_8115,N_8182);
nor U14849 (N_14849,N_5858,N_8049);
or U14850 (N_14850,N_7161,N_7312);
nor U14851 (N_14851,N_7085,N_5145);
xor U14852 (N_14852,N_6145,N_8756);
and U14853 (N_14853,N_6275,N_7176);
xor U14854 (N_14854,N_7894,N_5041);
or U14855 (N_14855,N_8749,N_9356);
nand U14856 (N_14856,N_9248,N_8475);
or U14857 (N_14857,N_5193,N_7880);
xor U14858 (N_14858,N_6361,N_9394);
xor U14859 (N_14859,N_6180,N_7608);
nand U14860 (N_14860,N_9536,N_8360);
and U14861 (N_14861,N_8018,N_7065);
xnor U14862 (N_14862,N_6978,N_5176);
nor U14863 (N_14863,N_9465,N_5377);
xnor U14864 (N_14864,N_7078,N_8154);
nand U14865 (N_14865,N_6989,N_5397);
or U14866 (N_14866,N_7728,N_7511);
or U14867 (N_14867,N_5536,N_6887);
xnor U14868 (N_14868,N_6911,N_9666);
nand U14869 (N_14869,N_9318,N_6912);
xor U14870 (N_14870,N_9072,N_5704);
nand U14871 (N_14871,N_6469,N_9933);
nand U14872 (N_14872,N_5023,N_8004);
or U14873 (N_14873,N_7034,N_7832);
nor U14874 (N_14874,N_8282,N_9816);
xor U14875 (N_14875,N_6811,N_9494);
and U14876 (N_14876,N_7448,N_5272);
and U14877 (N_14877,N_7945,N_5607);
and U14878 (N_14878,N_7577,N_7991);
nor U14879 (N_14879,N_5835,N_7177);
or U14880 (N_14880,N_6709,N_7732);
or U14881 (N_14881,N_8027,N_5361);
nand U14882 (N_14882,N_7451,N_7442);
or U14883 (N_14883,N_9739,N_8137);
nand U14884 (N_14884,N_8666,N_7977);
xor U14885 (N_14885,N_8514,N_7144);
nand U14886 (N_14886,N_9922,N_6033);
nand U14887 (N_14887,N_8329,N_8423);
nor U14888 (N_14888,N_9193,N_9132);
xor U14889 (N_14889,N_8641,N_9821);
nor U14890 (N_14890,N_5590,N_6706);
xnor U14891 (N_14891,N_7147,N_7414);
and U14892 (N_14892,N_7394,N_8992);
and U14893 (N_14893,N_9531,N_9009);
or U14894 (N_14894,N_8830,N_8955);
nor U14895 (N_14895,N_7985,N_7461);
nor U14896 (N_14896,N_8531,N_9086);
nor U14897 (N_14897,N_5032,N_5806);
nand U14898 (N_14898,N_8346,N_9586);
nand U14899 (N_14899,N_6305,N_6647);
nor U14900 (N_14900,N_5929,N_5920);
xnor U14901 (N_14901,N_5210,N_9535);
nor U14902 (N_14902,N_9873,N_6939);
nor U14903 (N_14903,N_6058,N_8022);
or U14904 (N_14904,N_9511,N_6683);
nand U14905 (N_14905,N_7877,N_7277);
and U14906 (N_14906,N_5912,N_9998);
nand U14907 (N_14907,N_8364,N_7147);
and U14908 (N_14908,N_8134,N_8469);
nor U14909 (N_14909,N_7924,N_5061);
nor U14910 (N_14910,N_5329,N_8949);
and U14911 (N_14911,N_9392,N_6847);
xor U14912 (N_14912,N_9520,N_7221);
xnor U14913 (N_14913,N_6147,N_7814);
nor U14914 (N_14914,N_6623,N_9748);
or U14915 (N_14915,N_9993,N_6980);
or U14916 (N_14916,N_5984,N_6000);
nand U14917 (N_14917,N_7623,N_9342);
xnor U14918 (N_14918,N_6501,N_9032);
or U14919 (N_14919,N_8793,N_8903);
nand U14920 (N_14920,N_8529,N_7098);
and U14921 (N_14921,N_8372,N_6698);
xor U14922 (N_14922,N_9613,N_7358);
or U14923 (N_14923,N_7679,N_6725);
nand U14924 (N_14924,N_6751,N_5932);
or U14925 (N_14925,N_6575,N_9977);
nor U14926 (N_14926,N_5237,N_6721);
nor U14927 (N_14927,N_5872,N_9488);
xnor U14928 (N_14928,N_7540,N_9862);
xnor U14929 (N_14929,N_7016,N_5157);
nor U14930 (N_14930,N_9396,N_9333);
xor U14931 (N_14931,N_6486,N_7526);
or U14932 (N_14932,N_7559,N_6829);
or U14933 (N_14933,N_8190,N_8306);
and U14934 (N_14934,N_7906,N_5115);
xnor U14935 (N_14935,N_5609,N_5888);
and U14936 (N_14936,N_7965,N_8877);
nand U14937 (N_14937,N_9313,N_9182);
nor U14938 (N_14938,N_8305,N_7995);
nor U14939 (N_14939,N_6975,N_8972);
and U14940 (N_14940,N_5924,N_7560);
or U14941 (N_14941,N_9007,N_6746);
and U14942 (N_14942,N_8961,N_5788);
nor U14943 (N_14943,N_8382,N_5226);
nor U14944 (N_14944,N_7605,N_9502);
and U14945 (N_14945,N_7789,N_6828);
nand U14946 (N_14946,N_9020,N_5892);
or U14947 (N_14947,N_5088,N_6237);
or U14948 (N_14948,N_5777,N_8170);
or U14949 (N_14949,N_5841,N_8331);
nor U14950 (N_14950,N_5323,N_7772);
and U14951 (N_14951,N_5318,N_9115);
xnor U14952 (N_14952,N_9049,N_5608);
xnor U14953 (N_14953,N_8926,N_6317);
nand U14954 (N_14954,N_7500,N_9522);
xor U14955 (N_14955,N_6109,N_5282);
nor U14956 (N_14956,N_5049,N_6117);
and U14957 (N_14957,N_8760,N_8784);
or U14958 (N_14958,N_9844,N_7596);
nor U14959 (N_14959,N_7641,N_6148);
nor U14960 (N_14960,N_8360,N_7008);
nor U14961 (N_14961,N_8185,N_5030);
nor U14962 (N_14962,N_8302,N_7754);
and U14963 (N_14963,N_5320,N_8509);
and U14964 (N_14964,N_7957,N_5877);
and U14965 (N_14965,N_8957,N_5910);
or U14966 (N_14966,N_8481,N_8885);
and U14967 (N_14967,N_7603,N_7154);
nand U14968 (N_14968,N_9936,N_8945);
nand U14969 (N_14969,N_8089,N_7973);
and U14970 (N_14970,N_5905,N_8777);
nand U14971 (N_14971,N_5388,N_5812);
xor U14972 (N_14972,N_9726,N_5882);
nand U14973 (N_14973,N_5465,N_7041);
xor U14974 (N_14974,N_7694,N_6306);
nand U14975 (N_14975,N_9854,N_9484);
xnor U14976 (N_14976,N_6194,N_5146);
nand U14977 (N_14977,N_9292,N_7192);
nand U14978 (N_14978,N_9473,N_6183);
xor U14979 (N_14979,N_7643,N_6992);
or U14980 (N_14980,N_8702,N_7721);
nand U14981 (N_14981,N_9394,N_5994);
or U14982 (N_14982,N_5927,N_8687);
nand U14983 (N_14983,N_5914,N_7116);
and U14984 (N_14984,N_9677,N_7138);
nor U14985 (N_14985,N_5805,N_5689);
nand U14986 (N_14986,N_8301,N_5563);
and U14987 (N_14987,N_7137,N_8443);
or U14988 (N_14988,N_9289,N_5314);
xor U14989 (N_14989,N_6731,N_6546);
or U14990 (N_14990,N_8321,N_7909);
xnor U14991 (N_14991,N_7667,N_8277);
xnor U14992 (N_14992,N_6168,N_8188);
or U14993 (N_14993,N_7360,N_6394);
or U14994 (N_14994,N_9411,N_9878);
or U14995 (N_14995,N_8900,N_8004);
xor U14996 (N_14996,N_6960,N_8949);
nand U14997 (N_14997,N_6200,N_7690);
nor U14998 (N_14998,N_8112,N_8309);
xnor U14999 (N_14999,N_5640,N_6537);
nand U15000 (N_15000,N_13241,N_11135);
and U15001 (N_15001,N_14272,N_10013);
xnor U15002 (N_15002,N_13693,N_12163);
and U15003 (N_15003,N_12628,N_12148);
or U15004 (N_15004,N_11309,N_14731);
nor U15005 (N_15005,N_13244,N_11457);
or U15006 (N_15006,N_12881,N_12434);
or U15007 (N_15007,N_12005,N_11323);
nor U15008 (N_15008,N_14945,N_11688);
xor U15009 (N_15009,N_13364,N_12446);
nor U15010 (N_15010,N_12290,N_10109);
or U15011 (N_15011,N_13183,N_12355);
xor U15012 (N_15012,N_14285,N_13897);
or U15013 (N_15013,N_12926,N_10317);
or U15014 (N_15014,N_12387,N_14630);
or U15015 (N_15015,N_13626,N_14369);
nand U15016 (N_15016,N_11462,N_13367);
nand U15017 (N_15017,N_13429,N_11911);
or U15018 (N_15018,N_10507,N_14335);
nor U15019 (N_15019,N_11321,N_13227);
xnor U15020 (N_15020,N_13519,N_11423);
xor U15021 (N_15021,N_11763,N_12248);
nor U15022 (N_15022,N_12865,N_12461);
and U15023 (N_15023,N_14486,N_11343);
nor U15024 (N_15024,N_12295,N_13194);
or U15025 (N_15025,N_13205,N_14210);
and U15026 (N_15026,N_10837,N_12943);
nand U15027 (N_15027,N_10902,N_10459);
and U15028 (N_15028,N_13507,N_14629);
nand U15029 (N_15029,N_13860,N_13251);
or U15030 (N_15030,N_10191,N_12950);
and U15031 (N_15031,N_12502,N_12339);
xor U15032 (N_15032,N_11981,N_13365);
or U15033 (N_15033,N_11219,N_12345);
xor U15034 (N_15034,N_14553,N_11224);
nand U15035 (N_15035,N_13585,N_14310);
xor U15036 (N_15036,N_13830,N_12838);
xnor U15037 (N_15037,N_14941,N_11929);
and U15038 (N_15038,N_11094,N_10921);
nand U15039 (N_15039,N_13483,N_14943);
or U15040 (N_15040,N_10187,N_11318);
nand U15041 (N_15041,N_13518,N_11259);
xor U15042 (N_15042,N_11667,N_10944);
nand U15043 (N_15043,N_12520,N_10570);
nand U15044 (N_15044,N_12814,N_11511);
xor U15045 (N_15045,N_11487,N_13823);
and U15046 (N_15046,N_14376,N_10068);
and U15047 (N_15047,N_10455,N_14537);
or U15048 (N_15048,N_11339,N_14114);
and U15049 (N_15049,N_14993,N_14153);
nor U15050 (N_15050,N_12066,N_13913);
and U15051 (N_15051,N_12021,N_11658);
xnor U15052 (N_15052,N_11228,N_11359);
or U15053 (N_15053,N_11895,N_10793);
or U15054 (N_15054,N_10935,N_11937);
nor U15055 (N_15055,N_14870,N_11006);
nand U15056 (N_15056,N_11016,N_11108);
nand U15057 (N_15057,N_12670,N_12555);
or U15058 (N_15058,N_14355,N_11971);
nor U15059 (N_15059,N_10952,N_13013);
or U15060 (N_15060,N_12609,N_14811);
and U15061 (N_15061,N_10805,N_11247);
nor U15062 (N_15062,N_12548,N_13953);
or U15063 (N_15063,N_12448,N_12222);
or U15064 (N_15064,N_14039,N_11510);
or U15065 (N_15065,N_13706,N_14116);
or U15066 (N_15066,N_13970,N_10370);
and U15067 (N_15067,N_13843,N_14934);
nand U15068 (N_15068,N_13619,N_11948);
and U15069 (N_15069,N_14052,N_10544);
nand U15070 (N_15070,N_11753,N_10644);
nand U15071 (N_15071,N_13672,N_11188);
and U15072 (N_15072,N_13359,N_12253);
and U15073 (N_15073,N_13445,N_12964);
nor U15074 (N_15074,N_14835,N_13766);
and U15075 (N_15075,N_10602,N_14389);
nor U15076 (N_15076,N_11888,N_10053);
xor U15077 (N_15077,N_10090,N_11074);
or U15078 (N_15078,N_12260,N_11477);
or U15079 (N_15079,N_12293,N_12676);
nor U15080 (N_15080,N_10433,N_13661);
nand U15081 (N_15081,N_12318,N_12763);
nand U15082 (N_15082,N_14051,N_10242);
nand U15083 (N_15083,N_13924,N_10227);
xor U15084 (N_15084,N_14273,N_10583);
nor U15085 (N_15085,N_14715,N_10612);
or U15086 (N_15086,N_12381,N_14798);
and U15087 (N_15087,N_11921,N_11090);
nor U15088 (N_15088,N_11407,N_11338);
nor U15089 (N_15089,N_12279,N_10384);
nand U15090 (N_15090,N_13182,N_11443);
nor U15091 (N_15091,N_13000,N_14854);
and U15092 (N_15092,N_12100,N_10220);
xor U15093 (N_15093,N_12765,N_10763);
or U15094 (N_15094,N_10324,N_14559);
nand U15095 (N_15095,N_10820,N_10450);
nand U15096 (N_15096,N_14387,N_12149);
or U15097 (N_15097,N_13263,N_11479);
nand U15098 (N_15098,N_13360,N_10446);
xnor U15099 (N_15099,N_13224,N_10458);
or U15100 (N_15100,N_11990,N_12603);
or U15101 (N_15101,N_13887,N_10173);
or U15102 (N_15102,N_12326,N_14303);
or U15103 (N_15103,N_11137,N_12540);
and U15104 (N_15104,N_10794,N_14446);
or U15105 (N_15105,N_12683,N_10253);
and U15106 (N_15106,N_10353,N_14328);
xnor U15107 (N_15107,N_14425,N_12761);
nor U15108 (N_15108,N_10801,N_13374);
nor U15109 (N_15109,N_14097,N_10589);
and U15110 (N_15110,N_12693,N_13189);
xnor U15111 (N_15111,N_14851,N_11024);
nor U15112 (N_15112,N_14007,N_13108);
and U15113 (N_15113,N_14020,N_12323);
or U15114 (N_15114,N_14912,N_10243);
xnor U15115 (N_15115,N_13678,N_10943);
and U15116 (N_15116,N_13687,N_14248);
and U15117 (N_15117,N_11036,N_11947);
and U15118 (N_15118,N_11742,N_13392);
and U15119 (N_15119,N_14860,N_10383);
and U15120 (N_15120,N_14562,N_11060);
and U15121 (N_15121,N_12501,N_11675);
xnor U15122 (N_15122,N_13488,N_12311);
nor U15123 (N_15123,N_13298,N_10228);
nor U15124 (N_15124,N_12993,N_11608);
or U15125 (N_15125,N_13748,N_11110);
nand U15126 (N_15126,N_10356,N_13259);
xnor U15127 (N_15127,N_11186,N_12760);
nand U15128 (N_15128,N_10899,N_13001);
and U15129 (N_15129,N_10697,N_10780);
xnor U15130 (N_15130,N_12625,N_13396);
or U15131 (N_15131,N_12064,N_10181);
nor U15132 (N_15132,N_13212,N_12504);
nor U15133 (N_15133,N_10928,N_10756);
nand U15134 (N_15134,N_11441,N_11004);
xnor U15135 (N_15135,N_11159,N_11583);
xor U15136 (N_15136,N_12821,N_14233);
and U15137 (N_15137,N_12666,N_13733);
or U15138 (N_15138,N_11845,N_14972);
xnor U15139 (N_15139,N_10895,N_14596);
nand U15140 (N_15140,N_10574,N_10627);
and U15141 (N_15141,N_14761,N_10639);
xnor U15142 (N_15142,N_10638,N_10704);
nand U15143 (N_15143,N_11672,N_10841);
or U15144 (N_15144,N_12882,N_11569);
nor U15145 (N_15145,N_11011,N_10042);
xor U15146 (N_15146,N_11153,N_14624);
nor U15147 (N_15147,N_11160,N_14735);
or U15148 (N_15148,N_14284,N_10819);
and U15149 (N_15149,N_11570,N_11623);
nand U15150 (N_15150,N_12480,N_13426);
and U15151 (N_15151,N_14380,N_10776);
nand U15152 (N_15152,N_11915,N_13495);
and U15153 (N_15153,N_14040,N_12493);
nand U15154 (N_15154,N_11481,N_14235);
xnor U15155 (N_15155,N_10481,N_13540);
or U15156 (N_15156,N_12107,N_10186);
nor U15157 (N_15157,N_12807,N_12197);
xnor U15158 (N_15158,N_14695,N_12811);
xnor U15159 (N_15159,N_14691,N_11982);
or U15160 (N_15160,N_10308,N_10876);
xnor U15161 (N_15161,N_13199,N_12376);
and U15162 (N_15162,N_11243,N_14329);
or U15163 (N_15163,N_10047,N_10674);
xor U15164 (N_15164,N_14085,N_14100);
and U15165 (N_15165,N_13627,N_11255);
xnor U15166 (N_15166,N_10543,N_13612);
nand U15167 (N_15167,N_12099,N_11871);
nand U15168 (N_15168,N_13350,N_14110);
nand U15169 (N_15169,N_14460,N_13968);
or U15170 (N_15170,N_12654,N_10518);
nor U15171 (N_15171,N_14247,N_13902);
xor U15172 (N_15172,N_10008,N_12090);
nand U15173 (N_15173,N_10931,N_10504);
nand U15174 (N_15174,N_14175,N_13048);
or U15175 (N_15175,N_14191,N_11540);
nand U15176 (N_15176,N_14089,N_13728);
nor U15177 (N_15177,N_10698,N_13208);
nor U15178 (N_15178,N_11154,N_12818);
nor U15179 (N_15179,N_13643,N_11308);
or U15180 (N_15180,N_11772,N_11528);
xor U15181 (N_15181,N_13237,N_11180);
or U15182 (N_15182,N_14279,N_10023);
and U15183 (N_15183,N_11263,N_11674);
or U15184 (N_15184,N_12517,N_14086);
and U15185 (N_15185,N_11082,N_10366);
nor U15186 (N_15186,N_11722,N_14594);
or U15187 (N_15187,N_12224,N_12622);
or U15188 (N_15188,N_11714,N_10429);
xnor U15189 (N_15189,N_11965,N_14255);
and U15190 (N_15190,N_13710,N_14593);
nor U15191 (N_15191,N_13117,N_12105);
or U15192 (N_15192,N_12539,N_12492);
nor U15193 (N_15193,N_14589,N_12344);
xnor U15194 (N_15194,N_12073,N_13074);
or U15195 (N_15195,N_12857,N_14892);
or U15196 (N_15196,N_13475,N_10717);
nand U15197 (N_15197,N_12787,N_13236);
nor U15198 (N_15198,N_13677,N_14287);
or U15199 (N_15199,N_10522,N_14215);
and U15200 (N_15200,N_12677,N_13279);
nor U15201 (N_15201,N_10653,N_10272);
nor U15202 (N_15202,N_14539,N_13320);
and U15203 (N_15203,N_12391,N_14877);
or U15204 (N_15204,N_14022,N_10728);
or U15205 (N_15205,N_11710,N_10655);
xnor U15206 (N_15206,N_12259,N_10405);
nand U15207 (N_15207,N_10267,N_10001);
and U15208 (N_15208,N_12331,N_11284);
nand U15209 (N_15209,N_11408,N_14887);
xor U15210 (N_15210,N_10108,N_10302);
or U15211 (N_15211,N_13885,N_13128);
xnor U15212 (N_15212,N_13688,N_11053);
nor U15213 (N_15213,N_10321,N_10011);
or U15214 (N_15214,N_12367,N_12496);
and U15215 (N_15215,N_12371,N_11784);
or U15216 (N_15216,N_14890,N_10865);
and U15217 (N_15217,N_11397,N_12794);
or U15218 (N_15218,N_12712,N_13016);
or U15219 (N_15219,N_10877,N_14508);
nor U15220 (N_15220,N_10814,N_11310);
or U15221 (N_15221,N_10437,N_10143);
and U15222 (N_15222,N_12553,N_13462);
and U15223 (N_15223,N_11253,N_14212);
xnor U15224 (N_15224,N_11774,N_11531);
or U15225 (N_15225,N_11890,N_12365);
or U15226 (N_15226,N_11257,N_11704);
or U15227 (N_15227,N_14345,N_12396);
and U15228 (N_15228,N_14340,N_11313);
or U15229 (N_15229,N_13379,N_11316);
nand U15230 (N_15230,N_10381,N_12579);
or U15231 (N_15231,N_11934,N_14384);
or U15232 (N_15232,N_14981,N_14652);
xor U15233 (N_15233,N_12209,N_12895);
nor U15234 (N_15234,N_13916,N_12270);
or U15235 (N_15235,N_13010,N_10200);
or U15236 (N_15236,N_14036,N_13466);
nand U15237 (N_15237,N_13769,N_10447);
and U15238 (N_15238,N_13102,N_14808);
nor U15239 (N_15239,N_10270,N_13451);
nand U15240 (N_15240,N_13210,N_14172);
xnor U15241 (N_15241,N_13720,N_10597);
and U15242 (N_15242,N_10705,N_12506);
or U15243 (N_15243,N_10682,N_12437);
nor U15244 (N_15244,N_12108,N_10726);
nor U15245 (N_15245,N_13448,N_13510);
xor U15246 (N_15246,N_14777,N_11141);
and U15247 (N_15247,N_12831,N_11616);
and U15248 (N_15248,N_10314,N_11113);
and U15249 (N_15249,N_10249,N_12644);
xor U15250 (N_15250,N_14527,N_12960);
and U15251 (N_15251,N_11726,N_11376);
or U15252 (N_15252,N_10092,N_13204);
and U15253 (N_15253,N_11374,N_12944);
nand U15254 (N_15254,N_13958,N_14482);
or U15255 (N_15255,N_12261,N_10375);
and U15256 (N_15256,N_12218,N_10217);
or U15257 (N_15257,N_14737,N_11748);
xor U15258 (N_15258,N_11562,N_10991);
and U15259 (N_15259,N_14987,N_12020);
nand U15260 (N_15260,N_11269,N_13509);
nor U15261 (N_15261,N_11773,N_14184);
or U15262 (N_15262,N_14617,N_11476);
nor U15263 (N_15263,N_12321,N_10293);
or U15264 (N_15264,N_12274,N_13543);
nor U15265 (N_15265,N_12007,N_11372);
xnor U15266 (N_15266,N_14045,N_12645);
nand U15267 (N_15267,N_14230,N_13494);
and U15268 (N_15268,N_14775,N_10539);
or U15269 (N_15269,N_14792,N_12598);
xor U15270 (N_15270,N_11061,N_10983);
xnor U15271 (N_15271,N_14054,N_13004);
nand U15272 (N_15272,N_11118,N_12836);
or U15273 (N_15273,N_12982,N_12413);
nand U15274 (N_15274,N_13268,N_11070);
xor U15275 (N_15275,N_14785,N_14107);
nand U15276 (N_15276,N_10010,N_11926);
nor U15277 (N_15277,N_13595,N_10083);
nor U15278 (N_15278,N_11837,N_13141);
xnor U15279 (N_15279,N_14888,N_14543);
nand U15280 (N_15280,N_14370,N_13640);
and U15281 (N_15281,N_13473,N_12822);
xnor U15282 (N_15282,N_12386,N_11187);
xnor U15283 (N_15283,N_10125,N_10231);
or U15284 (N_15284,N_10860,N_11600);
nand U15285 (N_15285,N_11549,N_13007);
and U15286 (N_15286,N_11687,N_10858);
or U15287 (N_15287,N_11300,N_13253);
xnor U15288 (N_15288,N_10609,N_14059);
nor U15289 (N_15289,N_14049,N_13030);
nand U15290 (N_15290,N_13232,N_13427);
nor U15291 (N_15291,N_10786,N_13944);
nand U15292 (N_15292,N_14965,N_14827);
xnor U15293 (N_15293,N_14137,N_12533);
xor U15294 (N_15294,N_10721,N_13699);
or U15295 (N_15295,N_14592,N_14757);
or U15296 (N_15296,N_11301,N_12035);
xor U15297 (N_15297,N_10968,N_11832);
or U15298 (N_15298,N_13152,N_13525);
nor U15299 (N_15299,N_13425,N_12534);
nand U15300 (N_15300,N_10176,N_12947);
nor U15301 (N_15301,N_11625,N_10028);
nor U15302 (N_15302,N_14618,N_13752);
nor U15303 (N_15303,N_12884,N_14318);
nand U15304 (N_15304,N_14050,N_10387);
and U15305 (N_15305,N_14448,N_14166);
and U15306 (N_15306,N_10277,N_14568);
nand U15307 (N_15307,N_10907,N_13808);
xnor U15308 (N_15308,N_13135,N_14183);
nor U15309 (N_15309,N_12507,N_13038);
xnor U15310 (N_15310,N_12864,N_10255);
or U15311 (N_15311,N_13267,N_11765);
and U15312 (N_15312,N_10525,N_10621);
nand U15313 (N_15313,N_14497,N_11523);
nand U15314 (N_15314,N_14032,N_14587);
nand U15315 (N_15315,N_11144,N_10166);
or U15316 (N_15316,N_10617,N_11745);
and U15317 (N_15317,N_11946,N_13032);
nand U15318 (N_15318,N_12731,N_14241);
xor U15319 (N_15319,N_11401,N_13285);
and U15320 (N_15320,N_12178,N_14462);
nand U15321 (N_15321,N_10020,N_12435);
and U15322 (N_15322,N_14003,N_10218);
and U15323 (N_15323,N_11370,N_13417);
nor U15324 (N_15324,N_14732,N_11448);
or U15325 (N_15325,N_12157,N_13115);
nand U15326 (N_15326,N_11565,N_11178);
or U15327 (N_15327,N_14891,N_13883);
nor U15328 (N_15328,N_10325,N_12310);
nand U15329 (N_15329,N_14544,N_10867);
and U15330 (N_15330,N_14584,N_14698);
xor U15331 (N_15331,N_10567,N_14582);
and U15332 (N_15332,N_10340,N_14721);
nand U15333 (N_15333,N_14694,N_12175);
and U15334 (N_15334,N_14101,N_10665);
and U15335 (N_15335,N_12254,N_12244);
nand U15336 (N_15336,N_14920,N_14591);
nand U15337 (N_15337,N_11587,N_14784);
xnor U15338 (N_15338,N_12255,N_13565);
and U15339 (N_15339,N_14496,N_12692);
and U15340 (N_15340,N_12056,N_14492);
and U15341 (N_15341,N_10880,N_10226);
and U15342 (N_15342,N_11322,N_11147);
nor U15343 (N_15343,N_11951,N_14122);
xnor U15344 (N_15344,N_10791,N_10828);
nor U15345 (N_15345,N_12348,N_13018);
nor U15346 (N_15346,N_14009,N_10813);
xor U15347 (N_15347,N_13896,N_13891);
nand U15348 (N_15348,N_10175,N_14160);
nor U15349 (N_15349,N_12181,N_14232);
xor U15350 (N_15350,N_11634,N_12220);
and U15351 (N_15351,N_13381,N_10560);
xnor U15352 (N_15352,N_12408,N_12116);
xor U15353 (N_15353,N_12127,N_12941);
and U15354 (N_15354,N_11179,N_10280);
xor U15355 (N_15355,N_14555,N_10884);
or U15356 (N_15356,N_14947,N_11719);
nor U15357 (N_15357,N_14487,N_11788);
and U15358 (N_15358,N_10113,N_14410);
nand U15359 (N_15359,N_10582,N_11679);
nand U15360 (N_15360,N_13880,N_14646);
or U15361 (N_15361,N_10371,N_13546);
nor U15362 (N_15362,N_13035,N_13855);
xor U15363 (N_15363,N_11385,N_12052);
and U15364 (N_15364,N_11474,N_10720);
nand U15365 (N_15365,N_13341,N_13110);
and U15366 (N_15366,N_11707,N_12679);
and U15367 (N_15367,N_14615,N_11514);
nor U15368 (N_15368,N_14633,N_12164);
nand U15369 (N_15369,N_14664,N_11863);
nor U15370 (N_15370,N_11126,N_13616);
nand U15371 (N_15371,N_13915,N_14470);
nand U15372 (N_15372,N_12184,N_10483);
nand U15373 (N_15373,N_10916,N_12590);
and U15374 (N_15374,N_13816,N_10487);
or U15375 (N_15375,N_10287,N_10804);
or U15376 (N_15376,N_14703,N_13261);
and U15377 (N_15377,N_12003,N_14106);
nand U15378 (N_15378,N_14653,N_13216);
xnor U15379 (N_15379,N_12126,N_14087);
or U15380 (N_15380,N_10792,N_11544);
nor U15381 (N_15381,N_14275,N_12277);
or U15382 (N_15382,N_12397,N_13929);
and U15383 (N_15383,N_14707,N_10117);
nand U15384 (N_15384,N_13991,N_13870);
nor U15385 (N_15385,N_14865,N_13029);
or U15386 (N_15386,N_10771,N_11584);
nand U15387 (N_15387,N_12133,N_14845);
and U15388 (N_15388,N_11568,N_11146);
nor U15389 (N_15389,N_10557,N_12605);
or U15390 (N_15390,N_12893,N_14187);
and U15391 (N_15391,N_10470,N_13729);
nand U15392 (N_15392,N_10336,N_12119);
nor U15393 (N_15393,N_14031,N_12920);
xnor U15394 (N_15394,N_11738,N_10009);
and U15395 (N_15395,N_13220,N_13812);
nor U15396 (N_15396,N_12247,N_11215);
or U15397 (N_15397,N_11708,N_11449);
nand U15398 (N_15398,N_10427,N_13561);
nor U15399 (N_15399,N_12725,N_11655);
nand U15400 (N_15400,N_12160,N_13239);
xnor U15401 (N_15401,N_12414,N_14725);
and U15402 (N_15402,N_11498,N_13788);
xnor U15403 (N_15403,N_10767,N_13994);
or U15404 (N_15404,N_14412,N_12588);
nand U15405 (N_15405,N_11556,N_11350);
xor U15406 (N_15406,N_13139,N_11290);
and U15407 (N_15407,N_10981,N_13165);
or U15408 (N_15408,N_11030,N_10775);
or U15409 (N_15409,N_12452,N_12878);
nor U15410 (N_15410,N_13273,N_13431);
nand U15411 (N_15411,N_13322,N_10888);
and U15412 (N_15412,N_14734,N_14399);
and U15413 (N_15413,N_11384,N_11334);
and U15414 (N_15414,N_12143,N_10099);
xnor U15415 (N_15415,N_12004,N_12201);
nor U15416 (N_15416,N_11553,N_14342);
nor U15417 (N_15417,N_12694,N_13945);
or U15418 (N_15418,N_12742,N_10873);
xnor U15419 (N_15419,N_10626,N_14852);
nor U15420 (N_15420,N_11242,N_11841);
xnor U15421 (N_15421,N_14859,N_13796);
xor U15422 (N_15422,N_11749,N_14162);
nand U15423 (N_15423,N_12384,N_10743);
xor U15424 (N_15424,N_12046,N_14619);
nand U15425 (N_15425,N_13335,N_11236);
nor U15426 (N_15426,N_11876,N_14177);
or U15427 (N_15427,N_10297,N_12611);
and U15428 (N_15428,N_10471,N_13719);
xor U15429 (N_15429,N_13511,N_11274);
nor U15430 (N_15430,N_12550,N_11701);
and U15431 (N_15431,N_14752,N_14138);
nand U15432 (N_15432,N_14008,N_11039);
xor U15433 (N_15433,N_11711,N_12389);
nand U15434 (N_15434,N_11266,N_13919);
and U15435 (N_15435,N_11602,N_14484);
and U15436 (N_15436,N_14306,N_12667);
and U15437 (N_15437,N_13697,N_14842);
xor U15438 (N_15438,N_10784,N_14129);
and U15439 (N_15439,N_11013,N_11648);
or U15440 (N_15440,N_14519,N_13017);
nand U15441 (N_15441,N_14069,N_14078);
nand U15442 (N_15442,N_14992,N_10711);
nor U15443 (N_15443,N_11050,N_12350);
or U15444 (N_15444,N_13614,N_13079);
xnor U15445 (N_15445,N_10380,N_14021);
and U15446 (N_15446,N_13600,N_12736);
or U15447 (N_15447,N_14787,N_10320);
xnor U15448 (N_15448,N_13144,N_10265);
nand U15449 (N_15449,N_12196,N_10783);
nand U15450 (N_15450,N_13105,N_14976);
and U15451 (N_15451,N_11303,N_13905);
and U15452 (N_15452,N_10030,N_10689);
or U15453 (N_15453,N_10139,N_14495);
nand U15454 (N_15454,N_10661,N_13844);
or U15455 (N_15455,N_11775,N_13323);
or U15456 (N_15456,N_13784,N_11611);
nor U15457 (N_15457,N_13072,N_10652);
xor U15458 (N_15458,N_11940,N_12970);
or U15459 (N_15459,N_12952,N_11330);
or U15460 (N_15460,N_14826,N_12888);
xor U15461 (N_15461,N_14350,N_11431);
nand U15462 (N_15462,N_14265,N_11654);
and U15463 (N_15463,N_10499,N_10448);
nand U15464 (N_15464,N_12886,N_10757);
and U15465 (N_15465,N_13704,N_14856);
or U15466 (N_15466,N_12967,N_11059);
and U15467 (N_15467,N_10643,N_13131);
and U15468 (N_15468,N_14576,N_14529);
nand U15469 (N_15469,N_14383,N_12971);
xor U15470 (N_15470,N_10723,N_14352);
or U15471 (N_15471,N_12854,N_13589);
nor U15472 (N_15472,N_10256,N_14195);
nor U15473 (N_15473,N_10922,N_13457);
nand U15474 (N_15474,N_12380,N_11936);
xnor U15475 (N_15475,N_13779,N_12833);
nor U15476 (N_15476,N_13670,N_12470);
nor U15477 (N_15477,N_10729,N_13631);
or U15478 (N_15478,N_10871,N_11741);
xor U15479 (N_15479,N_12795,N_14294);
nor U15480 (N_15480,N_14211,N_11446);
xor U15481 (N_15481,N_14840,N_14505);
xor U15482 (N_15482,N_13646,N_13372);
and U15483 (N_15483,N_11567,N_10393);
and U15484 (N_15484,N_11904,N_13920);
nand U15485 (N_15485,N_12232,N_12852);
or U15486 (N_15486,N_12406,N_11452);
and U15487 (N_15487,N_11652,N_10894);
and U15488 (N_15488,N_13420,N_12708);
nor U15489 (N_15489,N_11560,N_12567);
xor U15490 (N_15490,N_11521,N_12976);
and U15491 (N_15491,N_14764,N_11289);
or U15492 (N_15492,N_11345,N_13601);
or U15493 (N_15493,N_12804,N_13230);
nor U15494 (N_15494,N_10645,N_14711);
nand U15495 (N_15495,N_10295,N_14468);
or U15496 (N_15496,N_11103,N_12718);
xnor U15497 (N_15497,N_13685,N_12648);
nor U15498 (N_15498,N_14464,N_14830);
nor U15499 (N_15499,N_13847,N_10795);
and U15500 (N_15500,N_10900,N_10736);
nand U15501 (N_15501,N_14140,N_10378);
nor U15502 (N_15502,N_11996,N_10565);
nor U15503 (N_15503,N_12101,N_13330);
and U15504 (N_15504,N_11107,N_11536);
or U15505 (N_15505,N_10351,N_11882);
nand U15506 (N_15506,N_10891,N_14702);
and U15507 (N_15507,N_14001,N_10342);
or U15508 (N_15508,N_10164,N_11896);
and U15509 (N_15509,N_11478,N_14867);
xor U15510 (N_15510,N_13097,N_13098);
nor U15511 (N_15511,N_13743,N_13336);
xnor U15512 (N_15512,N_11184,N_10078);
or U15513 (N_15513,N_11258,N_13893);
nor U15514 (N_15514,N_14402,N_13022);
xor U15515 (N_15515,N_12031,N_11196);
nand U15516 (N_15516,N_13764,N_11931);
and U15517 (N_15517,N_14848,N_10057);
and U15518 (N_15518,N_13465,N_14699);
and U15519 (N_15519,N_14581,N_10806);
or U15520 (N_15520,N_14781,N_14683);
xnor U15521 (N_15521,N_11430,N_14662);
or U15522 (N_15522,N_14929,N_10524);
nor U15523 (N_15523,N_10950,N_11163);
nand U15524 (N_15524,N_11912,N_11437);
or U15525 (N_15525,N_11532,N_13215);
and U15526 (N_15526,N_13656,N_14977);
nand U15527 (N_15527,N_10953,N_11033);
and U15528 (N_15528,N_11121,N_10541);
xnor U15529 (N_15529,N_13401,N_14291);
or U15530 (N_15530,N_11174,N_11286);
xor U15531 (N_15531,N_14281,N_14440);
or U15532 (N_15532,N_14432,N_14741);
nor U15533 (N_15533,N_11597,N_13964);
and U15534 (N_15534,N_13084,N_12442);
xnor U15535 (N_15535,N_11908,N_13442);
or U15536 (N_15536,N_14799,N_14214);
nor U15537 (N_15537,N_12092,N_14753);
nor U15538 (N_15538,N_11496,N_14261);
or U15539 (N_15539,N_12552,N_10386);
xor U15540 (N_15540,N_12051,N_14414);
xor U15541 (N_15541,N_13985,N_14134);
or U15542 (N_15542,N_14546,N_11983);
xor U15543 (N_15543,N_14286,N_13516);
nand U15544 (N_15544,N_11432,N_10158);
nor U15545 (N_15545,N_10318,N_11907);
xnor U15546 (N_15546,N_14400,N_10555);
and U15547 (N_15547,N_12851,N_10039);
nor U15548 (N_15548,N_12607,N_11893);
nor U15549 (N_15549,N_11293,N_12786);
nand U15550 (N_15550,N_13394,N_10586);
nand U15551 (N_15551,N_13768,N_11312);
and U15552 (N_15552,N_12309,N_11960);
or U15553 (N_15553,N_13802,N_13177);
xnor U15554 (N_15554,N_11974,N_12221);
nand U15555 (N_15555,N_13801,N_11251);
nor U15556 (N_15556,N_12585,N_13109);
nor U15557 (N_15557,N_14874,N_11613);
nor U15558 (N_15558,N_14911,N_13171);
or U15559 (N_15559,N_14254,N_12165);
nand U15560 (N_15560,N_11172,N_12615);
and U15561 (N_15561,N_11513,N_10512);
nand U15562 (N_15562,N_12990,N_10863);
and U15563 (N_15563,N_10063,N_11678);
or U15564 (N_15564,N_14042,N_10138);
nand U15565 (N_15565,N_11545,N_11129);
nor U15566 (N_15566,N_10355,N_10064);
xor U15567 (N_15567,N_10159,N_11601);
and U15568 (N_15568,N_10829,N_13963);
nor U15569 (N_15569,N_10365,N_11870);
and U15570 (N_15570,N_10585,N_13548);
or U15571 (N_15571,N_13515,N_14933);
nor U15572 (N_15572,N_13295,N_12252);
and U15573 (N_15573,N_14718,N_12770);
xor U15574 (N_15574,N_13649,N_12200);
nor U15575 (N_15575,N_12668,N_14361);
xor U15576 (N_15576,N_12128,N_12809);
or U15577 (N_15577,N_12315,N_12012);
and U15578 (N_15578,N_11621,N_14686);
xor U15579 (N_15579,N_13209,N_11794);
xor U15580 (N_15580,N_10937,N_10851);
nand U15581 (N_15581,N_10059,N_13965);
and U15582 (N_15582,N_11910,N_14771);
nor U15583 (N_15583,N_10424,N_12497);
or U15584 (N_15584,N_11373,N_14509);
nand U15585 (N_15585,N_14037,N_14048);
nor U15586 (N_15586,N_12307,N_11148);
nor U15587 (N_15587,N_13922,N_10908);
nor U15588 (N_15588,N_13145,N_11731);
xor U15589 (N_15589,N_11220,N_11482);
nor U15590 (N_15590,N_14712,N_12084);
nand U15591 (N_15591,N_11485,N_11364);
nand U15592 (N_15592,N_14058,N_13718);
xor U15593 (N_15593,N_14857,N_13966);
or U15594 (N_15594,N_11579,N_14219);
xor U15595 (N_15595,N_12966,N_11203);
and U15596 (N_15596,N_10392,N_11516);
xnor U15597 (N_15597,N_12575,N_11020);
xnor U15598 (N_15598,N_12241,N_10987);
nand U15599 (N_15599,N_11614,N_10917);
nor U15600 (N_15600,N_12652,N_12558);
nor U15601 (N_15601,N_14719,N_11396);
nand U15602 (N_15602,N_11697,N_12623);
nand U15603 (N_15603,N_14364,N_14564);
or U15604 (N_15604,N_13116,N_11720);
nor U15605 (N_15605,N_14608,N_12398);
and U15606 (N_15606,N_10391,N_10789);
or U15607 (N_15607,N_11038,N_10210);
nor U15608 (N_15608,N_13500,N_14843);
nor U15609 (N_15609,N_13777,N_13909);
nor U15610 (N_15610,N_13120,N_12190);
nand U15611 (N_15611,N_12812,N_10664);
nor U15612 (N_15612,N_10846,N_14371);
or U15613 (N_15613,N_10666,N_11792);
xnor U15614 (N_15614,N_13787,N_12996);
nor U15615 (N_15615,N_14236,N_14171);
or U15616 (N_15616,N_12030,N_10869);
or U15617 (N_15617,N_11306,N_10016);
and U15618 (N_15618,N_10566,N_11806);
xor U15619 (N_15619,N_11461,N_13691);
nor U15620 (N_15620,N_13571,N_12193);
or U15621 (N_15621,N_14634,N_12587);
or U15622 (N_15622,N_13762,N_11003);
and U15623 (N_15623,N_14242,N_14397);
nand U15624 (N_15624,N_14660,N_13037);
nand U15625 (N_15625,N_12901,N_12094);
nand U15626 (N_15626,N_11043,N_10531);
nor U15627 (N_15627,N_12439,N_10230);
and U15628 (N_15628,N_10316,N_13889);
nor U15629 (N_15629,N_14747,N_10752);
and U15630 (N_15630,N_14417,N_11295);
xnor U15631 (N_15631,N_13156,N_13723);
nand U15632 (N_15632,N_11217,N_10215);
nand U15633 (N_15633,N_12302,N_13231);
xnor U15634 (N_15634,N_13538,N_13542);
nor U15635 (N_15635,N_14476,N_13650);
and U15636 (N_15636,N_10939,N_13983);
nand U15637 (N_15637,N_12429,N_13137);
and U15638 (N_15638,N_10050,N_11698);
nor U15639 (N_15639,N_12716,N_12956);
or U15640 (N_15640,N_13362,N_14733);
nor U15641 (N_15641,N_14493,N_14421);
nor U15642 (N_15642,N_11770,N_12395);
nor U15643 (N_15643,N_14358,N_10633);
nor U15644 (N_15644,N_11622,N_10812);
and U15645 (N_15645,N_11811,N_14194);
nor U15646 (N_15646,N_13714,N_10760);
and U15647 (N_15647,N_11447,N_10817);
or U15648 (N_15648,N_12825,N_11469);
nand U15649 (N_15649,N_14549,N_14043);
nor U15650 (N_15650,N_13886,N_13879);
nand U15651 (N_15651,N_11703,N_10992);
nand U15652 (N_15652,N_14909,N_13011);
or U15653 (N_15653,N_13256,N_11386);
or U15654 (N_15654,N_10441,N_10296);
and U15655 (N_15655,N_14612,N_14783);
and U15656 (N_15656,N_13358,N_14490);
or U15657 (N_15657,N_14360,N_10421);
and U15658 (N_15658,N_11232,N_14551);
and U15659 (N_15659,N_10658,N_13055);
nor U15660 (N_15660,N_13836,N_13342);
or U15661 (N_15661,N_10538,N_14079);
nand U15662 (N_15662,N_13703,N_12891);
and U15663 (N_15663,N_10641,N_14435);
and U15664 (N_15664,N_11723,N_11869);
xor U15665 (N_15665,N_14899,N_14096);
or U15666 (N_15666,N_10758,N_11683);
xnor U15667 (N_15667,N_10359,N_10493);
nor U15668 (N_15668,N_11807,N_14755);
and U15669 (N_15669,N_14262,N_10106);
xor U15670 (N_15670,N_14954,N_10299);
and U15671 (N_15671,N_11953,N_13147);
nor U15672 (N_15672,N_11925,N_13636);
and U15673 (N_15673,N_12931,N_12896);
or U15674 (N_15674,N_13077,N_13567);
and U15675 (N_15675,N_10882,N_12924);
nor U15676 (N_15676,N_13170,N_12919);
nor U15677 (N_15677,N_14207,N_14343);
nor U15678 (N_15678,N_14320,N_11851);
or U15679 (N_15679,N_14502,N_13597);
or U15680 (N_15680,N_13894,N_13193);
and U15681 (N_15681,N_10298,N_12917);
or U15682 (N_15682,N_11109,N_12112);
and U15683 (N_15683,N_12580,N_11575);
nand U15684 (N_15684,N_11311,N_14165);
and U15685 (N_15685,N_10065,N_13686);
and U15686 (N_15686,N_13221,N_10307);
nor U15687 (N_15687,N_11819,N_11636);
and U15688 (N_15688,N_10498,N_13744);
and U15689 (N_15689,N_14141,N_11642);
or U15690 (N_15690,N_13642,N_13539);
xor U15691 (N_15691,N_14846,N_11283);
nor U15692 (N_15692,N_10033,N_14075);
or U15693 (N_15693,N_13573,N_14829);
nand U15694 (N_15694,N_11199,N_12217);
nor U15695 (N_15695,N_11968,N_12636);
and U15696 (N_15696,N_13770,N_10588);
and U15697 (N_15697,N_13988,N_10932);
nand U15698 (N_15698,N_13052,N_10993);
xnor U15699 (N_15699,N_10310,N_14170);
nor U15700 (N_15700,N_12280,N_11231);
xnor U15701 (N_15701,N_10986,N_14533);
xnor U15702 (N_15702,N_12981,N_14418);
nand U15703 (N_15703,N_12897,N_13063);
or U15704 (N_15704,N_12136,N_12205);
nor U15705 (N_15705,N_10629,N_12167);
nor U15706 (N_15706,N_13095,N_12159);
nor U15707 (N_15707,N_10965,N_13091);
nor U15708 (N_15708,N_11665,N_10190);
nand U15709 (N_15709,N_10426,N_11102);
and U15710 (N_15710,N_12747,N_12935);
and U15711 (N_15711,N_14246,N_10745);
nor U15712 (N_15712,N_13809,N_10348);
nand U15713 (N_15713,N_10036,N_13089);
or U15714 (N_15714,N_10076,N_10192);
and U15715 (N_15715,N_14875,N_12571);
or U15716 (N_15716,N_12298,N_14794);
and U15717 (N_15717,N_13305,N_14226);
xor U15718 (N_15718,N_11944,N_10258);
nor U15719 (N_15719,N_11943,N_10677);
xor U15720 (N_15720,N_13190,N_11048);
nand U15721 (N_15721,N_11838,N_11168);
and U15722 (N_15722,N_11134,N_10761);
or U15723 (N_15723,N_12139,N_13839);
nor U15724 (N_15724,N_14006,N_12249);
nand U15725 (N_15725,N_12478,N_10466);
xor U15726 (N_15726,N_11344,N_14914);
nor U15727 (N_15727,N_14012,N_10443);
or U15728 (N_15728,N_13537,N_14128);
nor U15729 (N_15729,N_12037,N_13850);
or U15730 (N_15730,N_13845,N_12885);
nand U15731 (N_15731,N_11265,N_10003);
and U15732 (N_15732,N_11574,N_13006);
xor U15733 (N_15733,N_13933,N_13684);
and U15734 (N_15734,N_13249,N_12460);
nor U15735 (N_15735,N_11914,N_10216);
and U15736 (N_15736,N_10372,N_14062);
nand U15737 (N_15737,N_11816,N_12843);
nor U15738 (N_15738,N_14463,N_14253);
or U15739 (N_15739,N_13666,N_12154);
or U15740 (N_15740,N_11111,N_12879);
xnor U15741 (N_15741,N_14674,N_14837);
xor U15742 (N_15742,N_11887,N_13291);
nor U15743 (N_15743,N_13545,N_10046);
and U15744 (N_15744,N_10480,N_14905);
or U15745 (N_15745,N_13663,N_10716);
or U15746 (N_15746,N_13472,N_11918);
or U15747 (N_15747,N_12002,N_13833);
or U15748 (N_15748,N_11909,N_12029);
nand U15749 (N_15749,N_13828,N_10141);
xnor U15750 (N_15750,N_12939,N_13940);
nand U15751 (N_15751,N_11072,N_13574);
or U15752 (N_15752,N_14216,N_12988);
nor U15753 (N_15753,N_10910,N_11298);
nor U15754 (N_15754,N_13343,N_14392);
nand U15755 (N_15755,N_10580,N_12511);
or U15756 (N_15756,N_14550,N_10719);
or U15757 (N_15757,N_10881,N_14896);
xor U15758 (N_15758,N_12349,N_11506);
xor U15759 (N_15759,N_12710,N_12848);
and U15760 (N_15760,N_11840,N_13689);
or U15761 (N_15761,N_13954,N_12844);
nor U15762 (N_15762,N_11635,N_10077);
xnor U15763 (N_15763,N_12388,N_14540);
nand U15764 (N_15764,N_11620,N_11977);
xnor U15765 (N_15765,N_11421,N_11668);
xor U15766 (N_15766,N_14072,N_13155);
and U15767 (N_15767,N_14994,N_13329);
nand U15768 (N_15768,N_12018,N_13068);
nor U15769 (N_15769,N_13522,N_12547);
nor U15770 (N_15770,N_13984,N_11758);
and U15771 (N_15771,N_13624,N_14227);
xnor U15772 (N_15772,N_13039,N_13041);
nor U15773 (N_15773,N_10770,N_11942);
nor U15774 (N_15774,N_13033,N_10240);
xor U15775 (N_15775,N_14186,N_14638);
or U15776 (N_15776,N_12294,N_11027);
xnor U15777 (N_15777,N_13292,N_11361);
nand U15778 (N_15778,N_13834,N_13551);
nand U15779 (N_15779,N_12207,N_11963);
or U15780 (N_15780,N_12475,N_10982);
nor U15781 (N_15781,N_10203,N_10897);
nor U15782 (N_15782,N_10482,N_14937);
and U15783 (N_15783,N_14956,N_10311);
xnor U15784 (N_15784,N_12841,N_14099);
nand U15785 (N_15785,N_14292,N_13995);
xor U15786 (N_15786,N_14828,N_13630);
and U15787 (N_15787,N_12565,N_11434);
or U15788 (N_15788,N_11624,N_14644);
or U15789 (N_15789,N_11739,N_11883);
and U15790 (N_15790,N_14322,N_14224);
or U15791 (N_15791,N_11515,N_13774);
nand U15792 (N_15792,N_14903,N_11197);
nand U15793 (N_15793,N_13976,N_13283);
and U15794 (N_15794,N_10442,N_13653);
and U15795 (N_15795,N_13406,N_11502);
nor U15796 (N_15796,N_12213,N_12183);
nor U15797 (N_15797,N_14503,N_14963);
xnor U15798 (N_15798,N_11657,N_13191);
xnor U15799 (N_15799,N_10251,N_14814);
nand U15800 (N_15800,N_14117,N_14973);
nor U15801 (N_15801,N_13529,N_12065);
and U15802 (N_15802,N_11880,N_12554);
and U15803 (N_15803,N_12468,N_12292);
nand U15804 (N_15804,N_13439,N_10958);
xnor U15805 (N_15805,N_13803,N_14333);
and U15806 (N_15806,N_14507,N_13741);
nor U15807 (N_15807,N_13749,N_12685);
or U15808 (N_15808,N_13961,N_10974);
and U15809 (N_15809,N_14763,N_11445);
xor U15810 (N_15810,N_14071,N_12505);
nand U15811 (N_15811,N_13489,N_12256);
and U15812 (N_15812,N_13093,N_13921);
and U15813 (N_15813,N_14750,N_10616);
nor U15814 (N_15814,N_13613,N_10571);
nor U15815 (N_15815,N_11826,N_13197);
or U15816 (N_15816,N_12291,N_10975);
xor U15817 (N_15817,N_11085,N_12206);
nand U15818 (N_15818,N_12991,N_10537);
nand U15819 (N_15819,N_10632,N_10836);
nand U15820 (N_15820,N_13717,N_11835);
xor U15821 (N_15821,N_11241,N_13580);
nand U15822 (N_15822,N_11399,N_13554);
nor U15823 (N_15823,N_12503,N_12500);
and U15824 (N_15824,N_12977,N_14133);
nor U15825 (N_15825,N_14574,N_11718);
nand U15826 (N_15826,N_10556,N_10332);
nand U15827 (N_15827,N_12828,N_14547);
nor U15828 (N_15828,N_11450,N_14918);
or U15829 (N_15829,N_10396,N_14144);
or U15830 (N_15830,N_14063,N_10174);
nor U15831 (N_15831,N_10315,N_12420);
nor U15832 (N_15832,N_10290,N_12357);
nor U15833 (N_15833,N_11210,N_13042);
nand U15834 (N_15834,N_11873,N_14081);
or U15835 (N_15835,N_12135,N_14480);
nand U15836 (N_15836,N_13008,N_12120);
nand U15837 (N_15837,N_10262,N_12001);
or U15838 (N_15838,N_11052,N_14679);
and U15839 (N_15839,N_11058,N_10527);
or U15840 (N_15840,N_12068,N_10419);
or U15841 (N_15841,N_11713,N_11534);
nand U15842 (N_15842,N_11256,N_13986);
or U15843 (N_15843,N_14375,N_10741);
and U15844 (N_15844,N_12690,N_14156);
nand U15845 (N_15845,N_10740,N_13724);
and U15846 (N_15846,N_13569,N_11078);
and U15847 (N_15847,N_12788,N_11151);
nor U15848 (N_15848,N_13607,N_14919);
nor U15849 (N_15849,N_12194,N_11938);
or U15850 (N_15850,N_11631,N_11073);
xnor U15851 (N_15851,N_13901,N_12535);
xor U15852 (N_15852,N_12637,N_13338);
xor U15853 (N_15853,N_14455,N_14643);
xor U15854 (N_15854,N_13560,N_10561);
xnor U15855 (N_15855,N_14245,N_13700);
xnor U15856 (N_15856,N_12000,N_10222);
nor U15857 (N_15857,N_10343,N_10984);
xor U15858 (N_15858,N_11277,N_13412);
nor U15859 (N_15859,N_14636,N_13655);
nand U15860 (N_15860,N_11681,N_13853);
or U15861 (N_15861,N_11028,N_11539);
or U15862 (N_15862,N_11402,N_14471);
or U15863 (N_15863,N_10671,N_10630);
xnor U15864 (N_15864,N_11375,N_12286);
nor U15865 (N_15865,N_12490,N_14415);
xor U15866 (N_15866,N_13544,N_12912);
nor U15867 (N_15867,N_13050,N_10649);
or U15868 (N_15868,N_10738,N_11691);
nand U15869 (N_15869,N_14251,N_11035);
and U15870 (N_15870,N_10328,N_13872);
or U15871 (N_15871,N_11733,N_10438);
nor U15872 (N_15872,N_13639,N_13172);
and U15873 (N_15873,N_10416,N_10465);
xor U15874 (N_15874,N_10273,N_11573);
and U15875 (N_15875,N_12997,N_12859);
nand U15876 (N_15876,N_10404,N_13349);
and U15877 (N_15877,N_11026,N_11173);
or U15878 (N_15878,N_13975,N_11012);
nor U15879 (N_15879,N_14997,N_13592);
or U15880 (N_15880,N_14901,N_11800);
nor U15881 (N_15881,N_11662,N_14451);
or U15882 (N_15882,N_11858,N_10211);
nor U15883 (N_15883,N_14256,N_13671);
nand U15884 (N_15884,N_12146,N_11398);
nor U15885 (N_15885,N_13015,N_10552);
or U15886 (N_15886,N_12034,N_11182);
and U15887 (N_15887,N_11696,N_11664);
nor U15888 (N_15888,N_13528,N_11092);
nor U15889 (N_15889,N_14161,N_10759);
or U15890 (N_15890,N_10322,N_11405);
nor U15891 (N_15891,N_14046,N_12842);
and U15892 (N_15892,N_10274,N_13934);
nand U15893 (N_15893,N_11319,N_10478);
and U15894 (N_15894,N_10874,N_10978);
xor U15895 (N_15895,N_12370,N_12684);
nand U15896 (N_15896,N_14295,N_14714);
nand U15897 (N_15897,N_12394,N_12779);
xnor U15898 (N_15898,N_10599,N_11299);
xor U15899 (N_15899,N_14810,N_14379);
or U15900 (N_15900,N_14651,N_10261);
and U15901 (N_15901,N_13245,N_13579);
nand U15902 (N_15902,N_11966,N_14738);
nor U15903 (N_15903,N_14678,N_11355);
nand U15904 (N_15904,N_10156,N_10559);
nor U15905 (N_15905,N_12797,N_11305);
or U15906 (N_15906,N_14609,N_14898);
nor U15907 (N_15907,N_13405,N_13250);
and U15908 (N_15908,N_13882,N_13481);
nand U15909 (N_15909,N_14267,N_11932);
nor U15910 (N_15910,N_13243,N_14289);
and U15911 (N_15911,N_11041,N_14607);
and U15912 (N_15912,N_12890,N_12096);
xnor U15913 (N_15913,N_13384,N_14923);
or U15914 (N_15914,N_14422,N_12185);
and U15915 (N_15915,N_13054,N_13402);
nor U15916 (N_15916,N_10685,N_11561);
nor U15917 (N_15917,N_10954,N_14104);
nor U15918 (N_15918,N_12145,N_13240);
nand U15919 (N_15919,N_12269,N_13385);
and U15920 (N_15920,N_14374,N_13028);
xnor U15921 (N_15921,N_13841,N_12574);
nor U15922 (N_15922,N_11169,N_12242);
nand U15923 (N_15923,N_12450,N_10911);
or U15924 (N_15924,N_10435,N_10346);
and U15925 (N_15925,N_11751,N_13637);
or U15926 (N_15926,N_11769,N_11331);
or U15927 (N_15927,N_10768,N_11503);
nand U15928 (N_15928,N_10149,N_11285);
and U15929 (N_15929,N_13593,N_13807);
or U15930 (N_15930,N_13073,N_14192);
and U15931 (N_15931,N_12449,N_13694);
and U15932 (N_15932,N_13615,N_13066);
nor U15933 (N_15933,N_12032,N_13622);
and U15934 (N_15934,N_10578,N_10966);
nand U15935 (N_15935,N_13832,N_14998);
xor U15936 (N_15936,N_14442,N_14697);
nor U15937 (N_15937,N_13226,N_11804);
and U15938 (N_15938,N_10349,N_10184);
nor U15939 (N_15939,N_10089,N_12653);
and U15940 (N_15940,N_10915,N_13036);
xor U15941 (N_15941,N_11859,N_10093);
and U15942 (N_15942,N_13418,N_14847);
xnor U15943 (N_15943,N_13166,N_13760);
and U15944 (N_15944,N_12172,N_11973);
nand U15945 (N_15945,N_14528,N_13315);
and U15946 (N_15946,N_13805,N_13819);
nor U15947 (N_15947,N_13869,N_14779);
xor U15948 (N_15948,N_11145,N_13854);
nand U15949 (N_15949,N_10815,N_10476);
nand U15950 (N_15950,N_13188,N_10204);
nand U15951 (N_15951,N_13654,N_12313);
or U15952 (N_15952,N_10642,N_11860);
nor U15953 (N_15953,N_13932,N_10657);
or U15954 (N_15954,N_11123,N_11898);
nand U15955 (N_15955,N_11279,N_10497);
or U15956 (N_15956,N_11271,N_12424);
xor U15957 (N_15957,N_10170,N_11903);
or U15958 (N_15958,N_10049,N_14013);
xor U15959 (N_15959,N_14904,N_13758);
xnor U15960 (N_15960,N_14413,N_10115);
nor U15961 (N_15961,N_14791,N_14832);
and U15962 (N_15962,N_14491,N_11167);
or U15963 (N_15963,N_10233,N_13123);
and U15964 (N_15964,N_11578,N_11088);
nand U15965 (N_15965,N_10303,N_14688);
xor U15966 (N_15966,N_10535,N_11358);
xor U15967 (N_15967,N_11854,N_12796);
nor U15968 (N_15968,N_11492,N_12515);
nand U15969 (N_15969,N_10157,N_10027);
and U15970 (N_15970,N_13133,N_12862);
nor U15971 (N_15971,N_13611,N_12418);
xor U15972 (N_15972,N_13149,N_11252);
xor U15973 (N_15973,N_14222,N_11287);
nor U15974 (N_15974,N_14606,N_11821);
and U15975 (N_15975,N_14202,N_12122);
nand U15976 (N_15976,N_11671,N_10019);
nand U15977 (N_15977,N_14960,N_14436);
nand U15978 (N_15978,N_12764,N_13851);
and U15979 (N_15979,N_14047,N_10912);
nor U15980 (N_15980,N_12613,N_11239);
nand U15981 (N_15981,N_14426,N_12085);
nor U15982 (N_15982,N_12352,N_11962);
xnor U15983 (N_15983,N_12151,N_13644);
nor U15984 (N_15984,N_13321,N_13759);
and U15985 (N_15985,N_13390,N_12987);
nor U15986 (N_15986,N_10702,N_11750);
and U15987 (N_15987,N_10672,N_11865);
nand U15988 (N_15988,N_14332,N_12033);
and U15989 (N_15989,N_14944,N_10533);
nor U15990 (N_15990,N_11978,N_13252);
xnor U15991 (N_15991,N_13361,N_12273);
nor U15992 (N_15992,N_10257,N_11975);
and U15993 (N_15993,N_12487,N_14041);
xor U15994 (N_15994,N_14252,N_14305);
nand U15995 (N_15995,N_12789,N_13712);
xor U15996 (N_15996,N_13668,N_13277);
nor U15997 (N_15997,N_12297,N_14821);
or U15998 (N_15998,N_14809,N_10017);
nand U15999 (N_15999,N_12777,N_13304);
nor U16000 (N_16000,N_11161,N_12240);
and U16001 (N_16001,N_12612,N_14406);
nand U16002 (N_16002,N_10281,N_11661);
nor U16003 (N_16003,N_12422,N_13340);
xnor U16004 (N_16004,N_13219,N_11127);
nand U16005 (N_16005,N_12268,N_11555);
nor U16006 (N_16006,N_12810,N_11416);
nand U16007 (N_16007,N_11558,N_10807);
nor U16008 (N_16008,N_13606,N_14142);
nand U16009 (N_16009,N_10850,N_11037);
xor U16010 (N_16010,N_12556,N_10508);
xor U16011 (N_16011,N_11676,N_14314);
or U16012 (N_16012,N_14266,N_13825);
nand U16013 (N_16013,N_14642,N_11415);
or U16014 (N_16014,N_11850,N_10909);
xor U16015 (N_16015,N_13761,N_14315);
nor U16016 (N_16016,N_13081,N_12784);
nor U16017 (N_16017,N_14803,N_14511);
or U16018 (N_16018,N_11550,N_13707);
xor U16019 (N_16019,N_14288,N_13866);
or U16020 (N_16020,N_13301,N_12346);
nand U16021 (N_16021,N_11737,N_13871);
xnor U16022 (N_16022,N_13303,N_12737);
nor U16023 (N_16023,N_11730,N_10764);
and U16024 (N_16024,N_13260,N_13910);
xor U16025 (N_16025,N_10494,N_14542);
nand U16026 (N_16026,N_10144,N_10734);
and U16027 (N_16027,N_10601,N_14065);
nand U16028 (N_16028,N_12756,N_13815);
or U16029 (N_16029,N_14936,N_11031);
or U16030 (N_16030,N_12341,N_14458);
and U16031 (N_16031,N_14200,N_14598);
or U16032 (N_16032,N_11822,N_11116);
xnor U16033 (N_16033,N_13366,N_12599);
and U16034 (N_16034,N_10864,N_10706);
nor U16035 (N_16035,N_14701,N_12266);
xnor U16036 (N_16036,N_13657,N_14028);
xor U16037 (N_16037,N_11019,N_12874);
xor U16038 (N_16038,N_10856,N_12188);
xor U16039 (N_16039,N_13307,N_12182);
or U16040 (N_16040,N_12817,N_13150);
and U16041 (N_16041,N_13625,N_10269);
xnor U16042 (N_16042,N_10151,N_13460);
and U16043 (N_16043,N_11762,N_11055);
and U16044 (N_16044,N_13526,N_12191);
and U16045 (N_16045,N_14535,N_11191);
nand U16046 (N_16046,N_10898,N_14149);
xnor U16047 (N_16047,N_14481,N_11412);
nor U16048 (N_16048,N_11793,N_11454);
nor U16049 (N_16049,N_10418,N_11368);
and U16050 (N_16050,N_13633,N_13344);
nand U16051 (N_16051,N_14639,N_13876);
or U16052 (N_16052,N_13463,N_10648);
nand U16053 (N_16053,N_13114,N_13408);
nand U16054 (N_16054,N_11825,N_10887);
nor U16055 (N_16055,N_14474,N_14196);
nor U16056 (N_16056,N_11106,N_13316);
and U16057 (N_16057,N_11491,N_12563);
nand U16058 (N_16058,N_13302,N_11782);
nand U16059 (N_16059,N_11844,N_10744);
nor U16060 (N_16060,N_10727,N_10526);
nand U16061 (N_16061,N_14884,N_12186);
and U16062 (N_16062,N_14323,N_13536);
or U16063 (N_16063,N_14396,N_14472);
nand U16064 (N_16064,N_12855,N_12994);
xor U16065 (N_16065,N_12664,N_12942);
and U16066 (N_16066,N_14724,N_13129);
nor U16067 (N_16067,N_10964,N_11233);
xor U16068 (N_16068,N_12306,N_12285);
or U16069 (N_16069,N_11356,N_14499);
xnor U16070 (N_16070,N_14984,N_13848);
nand U16071 (N_16071,N_14130,N_13480);
xor U16072 (N_16072,N_14433,N_10883);
nor U16073 (N_16073,N_12359,N_13459);
nand U16074 (N_16074,N_13895,N_10596);
nand U16075 (N_16075,N_14311,N_13799);
or U16076 (N_16076,N_10388,N_12691);
xnor U16077 (N_16077,N_11820,N_11157);
xnor U16078 (N_16078,N_12739,N_11409);
and U16079 (N_16079,N_12871,N_14103);
nor U16080 (N_16080,N_10631,N_11889);
nand U16081 (N_16081,N_14897,N_12604);
and U16082 (N_16082,N_12695,N_10110);
or U16083 (N_16083,N_14260,N_11853);
and U16084 (N_16084,N_13454,N_12621);
xor U16085 (N_16085,N_13949,N_13926);
nand U16086 (N_16086,N_13482,N_11867);
xnor U16087 (N_16087,N_12237,N_12746);
xnor U16088 (N_16088,N_10330,N_11685);
or U16089 (N_16089,N_13835,N_13535);
xor U16090 (N_16090,N_10444,N_12117);
or U16091 (N_16091,N_12053,N_13083);
nand U16092 (N_16092,N_12512,N_13937);
xnor U16093 (N_16093,N_12142,N_14953);
nor U16094 (N_16094,N_14978,N_11970);
nor U16095 (N_16095,N_14601,N_10037);
nand U16096 (N_16096,N_13621,N_11508);
or U16097 (N_16097,N_14831,N_12203);
nand U16098 (N_16098,N_12748,N_12702);
and U16099 (N_16099,N_14070,N_12894);
or U16100 (N_16100,N_14632,N_12845);
xnor U16101 (N_16101,N_11803,N_11225);
or U16102 (N_16102,N_12019,N_13746);
and U16103 (N_16103,N_12658,N_14922);
nand U16104 (N_16104,N_12755,N_12887);
and U16105 (N_16105,N_12516,N_10096);
xnor U16106 (N_16106,N_11181,N_12379);
xor U16107 (N_16107,N_12072,N_11989);
and U16108 (N_16108,N_14163,N_14197);
nor U16109 (N_16109,N_12459,N_13067);
xnor U16110 (N_16110,N_10132,N_14748);
and U16111 (N_16111,N_14514,N_13453);
and U16112 (N_16112,N_12366,N_11383);
nand U16113 (N_16113,N_13690,N_13867);
or U16114 (N_16114,N_13877,N_11969);
xnor U16115 (N_16115,N_10167,N_14908);
xnor U16116 (N_16116,N_13076,N_13009);
and U16117 (N_16117,N_12866,N_11420);
xor U16118 (N_16118,N_14067,N_14249);
nor U16119 (N_16119,N_11029,N_12829);
and U16120 (N_16120,N_10859,N_14760);
and U16121 (N_16121,N_12471,N_14538);
nor U16122 (N_16122,N_12696,N_12419);
and U16123 (N_16123,N_12620,N_13176);
nor U16124 (N_16124,N_12906,N_13479);
nand U16125 (N_16125,N_14173,N_12687);
and U16126 (N_16126,N_11577,N_13721);
and U16127 (N_16127,N_14483,N_12543);
nand U16128 (N_16128,N_13508,N_12227);
or U16129 (N_16129,N_14969,N_11843);
xor U16130 (N_16130,N_10352,N_13939);
or U16131 (N_16131,N_11176,N_11992);
nand U16132 (N_16132,N_10886,N_13992);
xor U16133 (N_16133,N_10094,N_11440);
nand U16134 (N_16134,N_11133,N_14208);
or U16135 (N_16135,N_11817,N_13019);
nand U16136 (N_16136,N_12106,N_13012);
and U16137 (N_16137,N_11112,N_14325);
and U16138 (N_16138,N_10785,N_10713);
xor U16139 (N_16139,N_13875,N_14655);
xnor U16140 (N_16140,N_14602,N_11326);
nand U16141 (N_16141,N_10137,N_10656);
nor U16142 (N_16142,N_10341,N_13369);
nor U16143 (N_16143,N_10568,N_11205);
or U16144 (N_16144,N_12457,N_11935);
nand U16145 (N_16145,N_11471,N_10122);
xnor U16146 (N_16146,N_14740,N_12564);
and U16147 (N_16147,N_12234,N_14768);
and U16148 (N_16148,N_11660,N_10073);
and U16149 (N_16149,N_10335,N_10350);
xor U16150 (N_16150,N_14304,N_14467);
and U16151 (N_16151,N_14296,N_12238);
nand U16152 (N_16152,N_13257,N_13917);
nand U16153 (N_16153,N_11183,N_13513);
xor U16154 (N_16154,N_11473,N_14324);
and U16155 (N_16155,N_11238,N_10607);
and U16156 (N_16156,N_12669,N_14801);
xor U16157 (N_16157,N_13187,N_10623);
or U16158 (N_16158,N_12362,N_11490);
or U16159 (N_16159,N_13727,N_11632);
xor U16160 (N_16160,N_10831,N_12928);
nor U16161 (N_16161,N_12283,N_13403);
and U16162 (N_16162,N_12156,N_12324);
or U16163 (N_16163,N_13745,N_11554);
nand U16164 (N_16164,N_13040,N_11695);
nand U16165 (N_16165,N_11580,N_11245);
nand U16166 (N_16166,N_12759,N_12049);
nand U16167 (N_16167,N_12816,N_10345);
nand U16168 (N_16168,N_10263,N_12109);
xnor U16169 (N_16169,N_13941,N_13211);
xor U16170 (N_16170,N_14336,N_13584);
nand U16171 (N_16171,N_11930,N_10781);
and U16172 (N_16172,N_13207,N_13118);
or U16173 (N_16173,N_12081,N_13377);
or U16174 (N_16174,N_14501,N_14290);
xnor U16175 (N_16175,N_11798,N_12087);
nand U16176 (N_16176,N_10363,N_13857);
or U16177 (N_16177,N_12583,N_11488);
nor U16178 (N_16178,N_10124,N_11644);
nand U16179 (N_16179,N_14108,N_13444);
xnor U16180 (N_16180,N_14824,N_12245);
xnor U16181 (N_16181,N_14611,N_11861);
and U16182 (N_16182,N_14250,N_13810);
nand U16183 (N_16183,N_13101,N_13409);
and U16184 (N_16184,N_11424,N_14940);
nand U16185 (N_16185,N_10134,N_12929);
xnor U16186 (N_16186,N_13715,N_11292);
nand U16187 (N_16187,N_11288,N_11136);
nor U16188 (N_16188,N_14015,N_10040);
nand U16189 (N_16189,N_11143,N_10548);
nor U16190 (N_16190,N_14033,N_13327);
nor U16191 (N_16191,N_14180,N_13373);
or U16192 (N_16192,N_11234,N_11273);
or U16193 (N_16193,N_11752,N_12383);
nand U16194 (N_16194,N_13092,N_11280);
and U16195 (N_16195,N_11913,N_14386);
xnor U16196 (N_16196,N_14244,N_10377);
xor U16197 (N_16197,N_11520,N_11630);
nand U16198 (N_16198,N_14494,N_14309);
nand U16199 (N_16199,N_14924,N_13928);
and U16200 (N_16200,N_12700,N_12961);
and U16201 (N_16201,N_12875,N_12953);
nand U16202 (N_16202,N_10268,N_13765);
nor U16203 (N_16203,N_13938,N_12195);
or U16204 (N_16204,N_11779,N_14530);
xnor U16205 (N_16205,N_11008,N_10445);
nor U16206 (N_16206,N_11564,N_13383);
or U16207 (N_16207,N_12340,N_11015);
and U16208 (N_16208,N_12758,N_13918);
or U16209 (N_16209,N_13414,N_14942);
and U16210 (N_16210,N_14198,N_14135);
or U16211 (N_16211,N_11988,N_14516);
nand U16212 (N_16212,N_10730,N_12723);
xor U16213 (N_16213,N_10592,N_14650);
nor U16214 (N_16214,N_14706,N_13003);
xor U16215 (N_16215,N_13888,N_10488);
nor U16216 (N_16216,N_10395,N_13206);
nand U16217 (N_16217,N_11831,N_13817);
and U16218 (N_16218,N_13552,N_12236);
nor U16219 (N_16219,N_13874,N_11189);
nand U16220 (N_16220,N_11976,N_14344);
and U16221 (N_16221,N_10135,N_10634);
and U16222 (N_16222,N_12481,N_14955);
or U16223 (N_16223,N_11638,N_11426);
nor U16224 (N_16224,N_10542,N_12121);
and U16225 (N_16225,N_13380,N_14545);
nand U16226 (N_16226,N_10127,N_14676);
nand U16227 (N_16227,N_10832,N_14689);
nor U16228 (N_16228,N_12258,N_12039);
and U16229 (N_16229,N_12642,N_11522);
nand U16230 (N_16230,N_12016,N_11581);
xnor U16231 (N_16231,N_14682,N_13603);
or U16232 (N_16232,N_14357,N_13890);
or U16233 (N_16233,N_10575,N_11065);
nor U16234 (N_16234,N_12062,N_13818);
nand U16235 (N_16235,N_14670,N_11732);
nand U16236 (N_16236,N_10133,N_11018);
nand U16237 (N_16237,N_13785,N_13328);
or U16238 (N_16238,N_11114,N_13491);
nand U16239 (N_16239,N_14671,N_10201);
nand U16240 (N_16240,N_14125,N_10737);
or U16241 (N_16241,N_10436,N_13375);
nand U16242 (N_16242,N_12219,N_14240);
nor U16243 (N_16243,N_14167,N_13950);
or U16244 (N_16244,N_11439,N_11848);
nor U16245 (N_16245,N_14583,N_11693);
nand U16246 (N_16246,N_14950,N_12113);
and U16247 (N_16247,N_13389,N_12114);
nor U16248 (N_16248,N_14280,N_10147);
or U16249 (N_16249,N_14705,N_12328);
xnor U16250 (N_16250,N_11063,N_12688);
xnor U16251 (N_16251,N_12013,N_14168);
nand U16252 (N_16252,N_13881,N_10790);
or U16253 (N_16253,N_10693,N_14159);
nor U16254 (N_16254,N_13795,N_10415);
or U16255 (N_16255,N_10066,N_14672);
and U16256 (N_16256,N_12317,N_13989);
nor U16257 (N_16257,N_13532,N_12482);
or U16258 (N_16258,N_12477,N_11756);
nor U16259 (N_16259,N_11530,N_10501);
or U16260 (N_16260,N_14921,N_12701);
or U16261 (N_16261,N_13044,N_14239);
nor U16262 (N_16262,N_14690,N_12606);
xnor U16263 (N_16263,N_13735,N_12689);
nand U16264 (N_16264,N_11080,N_10893);
xor U16265 (N_16265,N_11377,N_10323);
nand U16266 (N_16266,N_10920,N_13811);
xor U16267 (N_16267,N_14193,N_12153);
nand U16268 (N_16268,N_12189,N_10239);
or U16269 (N_16269,N_12006,N_12403);
or U16270 (N_16270,N_12559,N_11686);
or U16271 (N_16271,N_13821,N_11669);
nand U16272 (N_16272,N_14786,N_10021);
nor U16273 (N_16273,N_13662,N_14727);
xor U16274 (N_16274,N_12170,N_10223);
or U16275 (N_16275,N_14276,N_12287);
nor U16276 (N_16276,N_11572,N_10300);
nand U16277 (N_16277,N_12719,N_13395);
and U16278 (N_16278,N_13111,N_13898);
and U16279 (N_16279,N_10683,N_10197);
nand U16280 (N_16280,N_14739,N_11856);
and U16281 (N_16281,N_14708,N_14238);
nor U16282 (N_16282,N_12918,N_13682);
nand U16283 (N_16283,N_11099,N_13363);
nor U16284 (N_16284,N_12909,N_10440);
nand U16285 (N_16285,N_11761,N_14925);
and U16286 (N_16286,N_12876,N_11891);
or U16287 (N_16287,N_12682,N_14510);
or U16288 (N_16288,N_13288,N_12026);
xnor U16289 (N_16289,N_14659,N_12103);
or U16290 (N_16290,N_11444,N_10647);
or U16291 (N_16291,N_14274,N_13286);
nand U16292 (N_16292,N_14880,N_13398);
nand U16293 (N_16293,N_11314,N_13043);
and U16294 (N_16294,N_13583,N_11746);
xnor U16295 (N_16295,N_14269,N_10972);
nand U16296 (N_16296,N_12486,N_14654);
and U16297 (N_16297,N_10857,N_13826);
nand U16298 (N_16298,N_14459,N_11789);
nor U16299 (N_16299,N_14823,N_11537);
xnor U16300 (N_16300,N_11754,N_12530);
nand U16301 (N_16301,N_11304,N_13790);
xor U16302 (N_16302,N_11905,N_10651);
xor U16303 (N_16303,N_10163,N_13517);
or U16304 (N_16304,N_11075,N_10146);
nor U16305 (N_16305,N_11229,N_14201);
nor U16306 (N_16306,N_13382,N_12498);
or U16307 (N_16307,N_10213,N_12369);
nor U16308 (N_16308,N_14518,N_13271);
nand U16309 (N_16309,N_13432,N_14895);
or U16310 (N_16310,N_14237,N_14313);
or U16311 (N_16311,N_12592,N_13228);
nand U16312 (N_16312,N_13711,N_11998);
xnor U16313 (N_16313,N_11598,N_13297);
xnor U16314 (N_16314,N_10208,N_14980);
nor U16315 (N_16315,N_11248,N_12877);
or U16316 (N_16316,N_13229,N_10259);
and U16317 (N_16317,N_12965,N_12714);
xnor U16318 (N_16318,N_12570,N_10473);
xnor U16319 (N_16319,N_14988,N_14390);
nand U16320 (N_16320,N_14815,N_13180);
xor U16321 (N_16321,N_12358,N_14473);
and U16322 (N_16322,N_10402,N_14966);
xnor U16323 (N_16323,N_13258,N_14704);
nor U16324 (N_16324,N_10309,N_14886);
nand U16325 (N_16325,N_14385,N_12337);
or U16326 (N_16326,N_12697,N_11152);
or U16327 (N_16327,N_14437,N_10367);
and U16328 (N_16328,N_11725,N_13311);
xor U16329 (N_16329,N_14521,N_10990);
and U16330 (N_16330,N_12063,N_10914);
xnor U16331 (N_16331,N_11933,N_13692);
and U16332 (N_16332,N_13107,N_11795);
nor U16333 (N_16333,N_10080,N_14881);
or U16334 (N_16334,N_10995,N_14558);
or U16335 (N_16335,N_14115,N_11100);
and U16336 (N_16336,N_10746,N_14088);
nand U16337 (N_16337,N_13702,N_14569);
or U16338 (N_16338,N_13458,N_13674);
and U16339 (N_16339,N_14302,N_13667);
xnor U16340 (N_16340,N_10827,N_13376);
nor U16341 (N_16341,N_10250,N_10788);
nand U16342 (N_16342,N_10389,N_13740);
and U16343 (N_16343,N_12780,N_13100);
nand U16344 (N_16344,N_11392,N_12629);
or U16345 (N_16345,N_13861,N_13096);
or U16346 (N_16346,N_14866,N_10368);
nor U16347 (N_16347,N_12899,N_14597);
nor U16348 (N_16348,N_12775,N_12491);
or U16349 (N_16349,N_10162,N_11955);
nor U16350 (N_16350,N_12288,N_13134);
or U16351 (N_16351,N_11320,N_14541);
and U16352 (N_16352,N_12070,N_12354);
or U16353 (N_16353,N_14985,N_14263);
or U16354 (N_16354,N_13202,N_10128);
nor U16355 (N_16355,N_10818,N_13586);
or U16356 (N_16356,N_10842,N_12671);
and U16357 (N_16357,N_14585,N_11389);
or U16358 (N_16358,N_11001,N_13952);
nor U16359 (N_16359,N_12392,N_13299);
xnor U16360 (N_16360,N_12465,N_10408);
and U16361 (N_16361,N_13865,N_11617);
or U16362 (N_16362,N_10700,N_12431);
or U16363 (N_16363,N_10692,N_11902);
nor U16364 (N_16364,N_12798,N_14700);
nor U16365 (N_16365,N_10803,N_10833);
nand U16366 (N_16366,N_11493,N_10102);
nand U16367 (N_16367,N_10714,N_14869);
nor U16368 (N_16368,N_12913,N_11347);
nor U16369 (N_16369,N_14112,N_14645);
or U16370 (N_16370,N_11814,N_10095);
nand U16371 (N_16371,N_13264,N_14271);
xnor U16372 (N_16372,N_14176,N_10521);
nor U16373 (N_16373,N_14368,N_10467);
or U16374 (N_16374,N_13806,N_10400);
and U16375 (N_16375,N_11158,N_13421);
xor U16376 (N_16376,N_14053,N_14030);
nand U16377 (N_16377,N_12025,N_12634);
and U16378 (N_16378,N_14206,N_11593);
and U16379 (N_16379,N_10489,N_12743);
nand U16380 (N_16380,N_11612,N_12610);
and U16381 (N_16381,N_11780,N_14150);
xor U16382 (N_16382,N_12948,N_14641);
or U16383 (N_16383,N_14359,N_14915);
nor U16384 (N_16384,N_10994,N_11666);
and U16385 (N_16385,N_11699,N_11588);
nand U16386 (N_16386,N_12672,N_12757);
nor U16387 (N_16387,N_10189,N_10007);
and U16388 (N_16388,N_10576,N_12820);
and U16389 (N_16389,N_14282,N_14872);
nand U16390 (N_16390,N_11264,N_12271);
nand U16391 (N_16391,N_14452,N_11244);
or U16392 (N_16392,N_10461,N_11237);
and U16393 (N_16393,N_10475,N_10862);
nor U16394 (N_16394,N_12858,N_14776);
xor U16395 (N_16395,N_12208,N_12753);
or U16396 (N_16396,N_10430,N_10890);
nor U16397 (N_16397,N_11227,N_14056);
xor U16398 (N_16398,N_10454,N_11815);
or U16399 (N_16399,N_11403,N_14566);
or U16400 (N_16400,N_11716,N_12055);
and U16401 (N_16401,N_11872,N_13254);
and U16402 (N_16402,N_12790,N_12239);
nand U16403 (N_16403,N_10084,N_13783);
xor U16404 (N_16404,N_10715,N_12910);
xnor U16405 (N_16405,N_12526,N_10892);
nor U16406 (N_16406,N_11294,N_14209);
and U16407 (N_16407,N_10834,N_10712);
nand U16408 (N_16408,N_12608,N_13797);
xor U16409 (N_16409,N_14152,N_10517);
nand U16410 (N_16410,N_10777,N_13681);
or U16411 (N_16411,N_10271,N_12407);
xnor U16412 (N_16412,N_12662,N_14579);
and U16413 (N_16413,N_12686,N_13138);
nand U16414 (N_16414,N_10722,N_10103);
nand U16415 (N_16415,N_13269,N_13126);
xnor U16416 (N_16416,N_14635,N_12597);
nor U16417 (N_16417,N_12856,N_10319);
nor U16418 (N_16418,N_11335,N_13911);
nand U16419 (N_16419,N_11997,N_12377);
and U16420 (N_16420,N_14479,N_13469);
nand U16421 (N_16421,N_14098,N_13490);
or U16422 (N_16422,N_11497,N_13773);
or U16423 (N_16423,N_10707,N_11595);
or U16424 (N_16424,N_11214,N_14948);
xnor U16425 (N_16425,N_10773,N_13326);
and U16426 (N_16426,N_14308,N_12524);
nor U16427 (N_16427,N_13447,N_12872);
nor U16428 (N_16428,N_14616,N_13370);
xor U16429 (N_16429,N_10848,N_13864);
and U16430 (N_16430,N_10930,N_11042);
xor U16431 (N_16431,N_10913,N_11728);
nor U16432 (N_16432,N_11875,N_10569);
nand U16433 (N_16433,N_12076,N_13562);
xor U16434 (N_16434,N_12447,N_11022);
or U16435 (N_16435,N_13737,N_14560);
xnor U16436 (N_16436,N_10926,N_13173);
xor U16437 (N_16437,N_13660,N_13776);
or U16438 (N_16438,N_13334,N_10357);
xnor U16439 (N_16439,N_11927,N_12803);
nor U16440 (N_16440,N_13085,N_14299);
nor U16441 (N_16441,N_10153,N_11509);
nor U16442 (N_16442,N_12749,N_12813);
xor U16443 (N_16443,N_13575,N_10662);
and U16444 (N_16444,N_13820,N_13113);
nor U16445 (N_16445,N_11923,N_13951);
xnor U16446 (N_16446,N_11680,N_14119);
and U16447 (N_16447,N_13969,N_10670);
xor U16448 (N_16448,N_14668,N_10098);
nor U16449 (N_16449,N_13587,N_12572);
nand U16450 (N_16450,N_11906,N_14577);
nand U16451 (N_16451,N_10545,N_13998);
and U16452 (N_16452,N_12440,N_14669);
nand U16453 (N_16453,N_10904,N_11353);
nand U16454 (N_16454,N_11429,N_12272);
xor U16455 (N_16455,N_13506,N_12751);
or U16456 (N_16456,N_11246,N_11460);
xnor U16457 (N_16457,N_13862,N_12028);
nand U16458 (N_16458,N_11689,N_11690);
xor U16459 (N_16459,N_12927,N_14736);
and U16460 (N_16460,N_12415,N_13002);
and U16461 (N_16461,N_12423,N_12800);
or U16462 (N_16462,N_13056,N_14666);
nor U16463 (N_16463,N_13300,N_14354);
and U16464 (N_16464,N_14349,N_13049);
or U16465 (N_16465,N_13514,N_11084);
and U16466 (N_16466,N_10301,N_10572);
xor U16467 (N_16467,N_13629,N_13947);
and U16468 (N_16468,N_12529,N_14983);
xnor U16469 (N_16469,N_13549,N_14377);
or U16470 (N_16470,N_13434,N_11647);
xnor U16471 (N_16471,N_10291,N_12304);
xor U16472 (N_16472,N_11874,N_14673);
xor U16473 (N_16473,N_11984,N_10668);
and U16474 (N_16474,N_12602,N_13568);
or U16475 (N_16475,N_13599,N_11463);
xor U16476 (N_16476,N_12846,N_11164);
or U16477 (N_16477,N_10821,N_12093);
xor U16478 (N_16478,N_10718,N_10048);
nor U16479 (N_16479,N_11619,N_11541);
xor U16480 (N_16480,N_11348,N_10595);
and U16481 (N_16481,N_11362,N_14366);
nand U16482 (N_16482,N_13982,N_10505);
nor U16483 (N_16483,N_12451,N_11120);
nor U16484 (N_16484,N_12849,N_11956);
xnor U16485 (N_16485,N_10696,N_13676);
nor U16486 (N_16486,N_14217,N_12361);
nor U16487 (N_16487,N_11221,N_14982);
xor U16488 (N_16488,N_14728,N_11425);
nand U16489 (N_16489,N_11064,N_14604);
xnor U16490 (N_16490,N_13912,N_11500);
nor U16491 (N_16491,N_12353,N_13218);
xor U16492 (N_16492,N_10326,N_12179);
xor U16493 (N_16493,N_10938,N_12230);
and U16494 (N_16494,N_10338,N_13130);
xnor U16495 (N_16495,N_14297,N_13972);
or U16496 (N_16496,N_12523,N_10058);
or U16497 (N_16497,N_12129,N_14298);
xnor U16498 (N_16498,N_14327,N_14228);
or U16499 (N_16499,N_11673,N_13647);
nand U16500 (N_16500,N_14628,N_11079);
nand U16501 (N_16501,N_12180,N_14408);
or U16502 (N_16502,N_10294,N_10390);
xnor U16503 (N_16503,N_11917,N_11954);
xor U16504 (N_16504,N_13413,N_10646);
nor U16505 (N_16505,N_12963,N_14025);
xor U16506 (N_16506,N_13499,N_10024);
nand U16507 (N_16507,N_10035,N_12338);
or U16508 (N_16508,N_11201,N_12263);
xor U16509 (N_16509,N_14663,N_10120);
and U16510 (N_16510,N_14816,N_11340);
and U16511 (N_16511,N_11394,N_10854);
nand U16512 (N_16512,N_12921,N_14910);
nand U16513 (N_16513,N_11586,N_12647);
nand U16514 (N_16514,N_14833,N_11694);
xnor U16515 (N_16515,N_10081,N_11115);
nand U16516 (N_16516,N_12289,N_14454);
nor U16517 (N_16517,N_12428,N_11894);
and U16518 (N_16518,N_12705,N_11216);
or U16519 (N_16519,N_13531,N_13763);
nand U16520 (N_16520,N_14853,N_10622);
and U16521 (N_16521,N_11054,N_14337);
nand U16522 (N_16522,N_10659,N_11192);
nor U16523 (N_16523,N_10941,N_12569);
or U16524 (N_16524,N_14720,N_13732);
and U16525 (N_16525,N_13669,N_12902);
nor U16526 (N_16526,N_13476,N_12911);
nor U16527 (N_16527,N_13892,N_13604);
nor U16528 (N_16528,N_13185,N_14743);
xnor U16529 (N_16529,N_14365,N_14353);
xnor U16530 (N_16530,N_12883,N_14334);
nor U16531 (N_16531,N_13858,N_11382);
nand U16532 (N_16532,N_13555,N_14123);
or U16533 (N_16533,N_11764,N_13275);
nor U16534 (N_16534,N_11834,N_14204);
nor U16535 (N_16535,N_13582,N_12771);
nor U16536 (N_16536,N_11877,N_10229);
and U16537 (N_16537,N_12373,N_11878);
and U16538 (N_16538,N_13927,N_10292);
nor U16539 (N_16539,N_14498,N_11240);
or U16540 (N_16540,N_10516,N_13782);
xnor U16541 (N_16541,N_13609,N_12726);
or U16542 (N_16542,N_11261,N_14478);
nand U16543 (N_16543,N_12892,N_11138);
nor U16544 (N_16544,N_14957,N_13793);
nor U16545 (N_16545,N_10614,N_13468);
or U16546 (N_16546,N_12537,N_10523);
and U16547 (N_16547,N_10564,N_14157);
xor U16548 (N_16548,N_11324,N_11342);
and U16549 (N_16549,N_12417,N_13563);
xor U16550 (N_16550,N_14469,N_11349);
nor U16551 (N_16551,N_14868,N_10963);
and U16552 (N_16552,N_13849,N_11387);
nor U16553 (N_16553,N_10681,N_12541);
nor U16554 (N_16554,N_10615,N_11501);
or U16555 (N_16555,N_12772,N_10434);
nor U16556 (N_16556,N_10289,N_12333);
and U16557 (N_16557,N_13422,N_11049);
xor U16558 (N_16558,N_10376,N_14762);
and U16559 (N_16559,N_14996,N_11302);
nor U16560 (N_16560,N_14394,N_13146);
and U16561 (N_16561,N_14439,N_12853);
or U16562 (N_16562,N_14268,N_13353);
nand U16563 (N_16563,N_14778,N_13695);
or U16564 (N_16564,N_11466,N_10194);
and U16565 (N_16565,N_12635,N_10573);
nand U16566 (N_16566,N_10751,N_11591);
nand U16567 (N_16567,N_12561,N_14179);
or U16568 (N_16568,N_12284,N_12880);
nor U16569 (N_16569,N_14746,N_12485);
or U16570 (N_16570,N_12041,N_13608);
nand U16571 (N_16571,N_12368,N_13443);
nor U16572 (N_16572,N_14372,N_11404);
and U16573 (N_16573,N_13023,N_10154);
xnor U16574 (N_16574,N_12216,N_11928);
nand U16575 (N_16575,N_13354,N_11223);
nand U16576 (N_16576,N_12681,N_13281);
nor U16577 (N_16577,N_11590,N_14825);
or U16578 (N_16578,N_13946,N_12989);
nand U16579 (N_16579,N_10360,N_13683);
nand U16580 (N_16580,N_13143,N_12951);
xor U16581 (N_16581,N_10962,N_13325);
xnor U16582 (N_16582,N_13464,N_12925);
nand U16583 (N_16583,N_10169,N_11985);
nor U16584 (N_16584,N_12363,N_10844);
and U16585 (N_16585,N_13203,N_10624);
or U16586 (N_16586,N_14427,N_13635);
and U16587 (N_16587,N_14312,N_11380);
xor U16588 (N_16588,N_12474,N_13750);
and U16589 (N_16589,N_13154,N_10004);
xor U16590 (N_16590,N_13960,N_11021);
xnor U16591 (N_16591,N_12432,N_11010);
nor U16592 (N_16592,N_10244,N_14716);
xnor U16593 (N_16593,N_14742,N_11852);
xnor U16594 (N_16594,N_12568,N_13755);
xor U16595 (N_16595,N_13306,N_13157);
and U16596 (N_16596,N_11829,N_13930);
xnor U16597 (N_16597,N_11083,N_13351);
nand U16598 (N_16598,N_13075,N_14861);
xnor U16599 (N_16599,N_10506,N_14967);
nor U16600 (N_16600,N_14793,N_12630);
nand U16601 (N_16601,N_12830,N_14080);
xnor U16602 (N_16602,N_11736,N_14805);
xnor U16603 (N_16603,N_11552,N_14817);
or U16604 (N_16604,N_13617,N_14586);
or U16605 (N_16605,N_12754,N_12699);
or U16606 (N_16606,N_13140,N_14526);
or U16607 (N_16607,N_12969,N_10460);
nand U16608 (N_16608,N_11175,N_12479);
xor U16609 (N_16609,N_11939,N_10515);
or U16610 (N_16610,N_11507,N_10453);
and U16611 (N_16611,N_12017,N_13386);
and U16612 (N_16612,N_14223,N_11198);
nand U16613 (N_16613,N_12401,N_14419);
nand U16614 (N_16614,N_12508,N_12125);
nor U16615 (N_16615,N_10085,N_13959);
nor U16616 (N_16616,N_12347,N_13378);
or U16617 (N_16617,N_12934,N_14802);
nor U16618 (N_16618,N_10640,N_12192);
and U16619 (N_16619,N_10825,N_13339);
and U16620 (N_16620,N_11165,N_10811);
or U16621 (N_16621,N_10462,N_11656);
nor U16622 (N_16622,N_11204,N_10439);
nand U16623 (N_16623,N_13357,N_14221);
nor U16624 (N_16624,N_10709,N_13907);
nand U16625 (N_16625,N_14774,N_13088);
xor U16626 (N_16626,N_12336,N_14621);
nand U16627 (N_16627,N_12111,N_13610);
nand U16628 (N_16628,N_10970,N_12009);
xnor U16629 (N_16629,N_12799,N_14525);
nor U16630 (N_16630,N_11767,N_14961);
or U16631 (N_16631,N_14769,N_14873);
and U16632 (N_16632,N_11260,N_10579);
nor U16633 (N_16633,N_10014,N_12639);
nor U16634 (N_16634,N_14293,N_13736);
xnor U16635 (N_16635,N_10031,N_12410);
or U16636 (N_16636,N_10620,N_12745);
nand U16637 (N_16637,N_14878,N_12752);
xnor U16638 (N_16638,N_11438,N_12104);
or U16639 (N_16639,N_12720,N_12984);
and U16640 (N_16640,N_14338,N_12704);
or U16641 (N_16641,N_10275,N_11149);
and U16642 (N_16642,N_11034,N_14958);
and U16643 (N_16643,N_11315,N_14220);
xor U16644 (N_16644,N_10594,N_11422);
nand U16645 (N_16645,N_14554,N_14522);
xnor U16646 (N_16646,N_12320,N_14199);
nand U16647 (N_16647,N_12861,N_13317);
and U16648 (N_16648,N_11864,N_10839);
nor U16649 (N_16649,N_12785,N_11459);
nor U16650 (N_16650,N_10996,N_14661);
xnor U16651 (N_16651,N_12792,N_10823);
xor U16652 (N_16652,N_12204,N_13356);
nand U16653 (N_16653,N_11097,N_10205);
nor U16654 (N_16654,N_11453,N_14094);
nand U16655 (N_16655,N_14906,N_14019);
and U16656 (N_16656,N_11778,N_13333);
nor U16657 (N_16657,N_12791,N_14766);
xnor U16658 (N_16658,N_10998,N_12806);
nor U16659 (N_16659,N_13200,N_11849);
or U16660 (N_16660,N_12992,N_10358);
xor U16661 (N_16661,N_12525,N_13058);
or U16662 (N_16662,N_12721,N_11131);
and U16663 (N_16663,N_12469,N_11162);
xor U16664 (N_16664,N_12898,N_11824);
nand U16665 (N_16665,N_13234,N_12161);
xnor U16666 (N_16666,N_13856,N_11464);
and U16667 (N_16667,N_14986,N_10866);
or U16668 (N_16668,N_13800,N_10241);
xor U16669 (N_16669,N_10472,N_13973);
nand U16670 (N_16670,N_13223,N_10168);
nand U16671 (N_16671,N_10802,N_11897);
xnor U16672 (N_16672,N_13163,N_12802);
nand U16673 (N_16673,N_11957,N_14952);
and U16674 (N_16674,N_12824,N_10142);
nand U16675 (N_16675,N_11428,N_10528);
nand U16676 (N_16676,N_12733,N_11999);
and U16677 (N_16677,N_10948,N_13786);
and U16678 (N_16678,N_14517,N_11494);
nand U16679 (N_16679,N_10252,N_10072);
or U16680 (N_16680,N_12303,N_14164);
nor U16681 (N_16681,N_14506,N_13486);
nand U16682 (N_16682,N_11066,N_10140);
and U16683 (N_16683,N_13148,N_12834);
nor U16684 (N_16684,N_14627,N_12805);
or U16685 (N_16685,N_11360,N_12138);
or U16686 (N_16686,N_10403,N_10628);
nor U16687 (N_16687,N_12673,N_13242);
nand U16688 (N_16688,N_14434,N_14850);
xnor U16689 (N_16689,N_12980,N_12243);
and U16690 (N_16690,N_10762,N_11812);
nand U16691 (N_16691,N_10254,N_14964);
and U16692 (N_16692,N_10988,N_10969);
nor U16693 (N_16693,N_11200,N_11427);
xor U16694 (N_16694,N_12215,N_13213);
nand U16695 (N_16695,N_13623,N_12781);
xnor U16696 (N_16696,N_14572,N_10136);
nand U16697 (N_16697,N_11866,N_13756);
xor U16698 (N_16698,N_10625,N_11833);
nand U16699 (N_16699,N_14819,N_12827);
xor U16700 (N_16700,N_12578,N_14789);
and U16701 (N_16701,N_12050,N_12264);
and U16702 (N_16702,N_10703,N_12048);
xor U16703 (N_16703,N_14640,N_11378);
xor U16704 (N_16704,N_13387,N_12619);
xnor U16705 (N_16705,N_13641,N_12300);
xnor U16706 (N_16706,N_14010,N_14401);
nand U16707 (N_16707,N_14283,N_12322);
xnor U16708 (N_16708,N_12102,N_12873);
or U16709 (N_16709,N_11706,N_10500);
nor U16710 (N_16710,N_14788,N_10951);
xor U16711 (N_16711,N_10495,N_11727);
xor U16712 (N_16712,N_10510,N_12134);
nand U16713 (N_16713,N_14907,N_13455);
nor U16714 (N_16714,N_11609,N_10160);
nand U16715 (N_16715,N_14534,N_14014);
or U16716 (N_16716,N_14971,N_14143);
xor U16717 (N_16717,N_13346,N_13497);
and U16718 (N_16718,N_11193,N_14900);
nor U16719 (N_16719,N_13899,N_12655);
and U16720 (N_16720,N_10145,N_10774);
or U16721 (N_16721,N_14931,N_14424);
nor U16722 (N_16722,N_12562,N_13112);
nand U16723 (N_16723,N_12071,N_14351);
and U16724 (N_16724,N_12594,N_11760);
or U16725 (N_16725,N_14131,N_13838);
xnor U16726 (N_16726,N_10206,N_12374);
nand U16727 (N_16727,N_13814,N_12527);
or U16728 (N_16728,N_10725,N_10051);
nand U16729 (N_16729,N_10022,N_10747);
xor U16730 (N_16730,N_14523,N_12614);
nor U16731 (N_16731,N_11759,N_13046);
or U16732 (N_16732,N_10177,N_11352);
or U16733 (N_16733,N_11512,N_11418);
and U16734 (N_16734,N_10509,N_13125);
nand U16735 (N_16735,N_14061,N_12329);
xor U16736 (N_16736,N_14091,N_12727);
or U16737 (N_16737,N_14990,N_10540);
and U16738 (N_16738,N_11317,N_12581);
nand U16739 (N_16739,N_13070,N_14148);
and U16740 (N_16740,N_14665,N_14382);
and U16741 (N_16741,N_13284,N_13449);
nand U16742 (N_16742,N_13159,N_14169);
nor U16743 (N_16743,N_11783,N_11222);
nand U16744 (N_16744,N_10407,N_11395);
nor U16745 (N_16745,N_11791,N_12466);
nand U16746 (N_16746,N_13433,N_12400);
and U16747 (N_16747,N_13060,N_10079);
xnor U16748 (N_16748,N_12199,N_12509);
or U16749 (N_16749,N_14841,N_10054);
and U16750 (N_16750,N_11077,N_13962);
xnor U16751 (N_16751,N_12257,N_10945);
or U16752 (N_16752,N_13680,N_12903);
and U16753 (N_16753,N_10959,N_10456);
or U16754 (N_16754,N_10212,N_14782);
nand U16755 (N_16755,N_10772,N_10409);
xnor U16756 (N_16756,N_10919,N_11524);
and U16757 (N_16757,N_12131,N_13651);
and U16758 (N_16758,N_12646,N_10611);
nand U16759 (N_16759,N_14532,N_11366);
and U16760 (N_16760,N_11684,N_12837);
nor U16761 (N_16761,N_11139,N_14855);
nor U16762 (N_16762,N_12573,N_13726);
nor U16763 (N_16763,N_13771,N_12098);
xnor U16764 (N_16764,N_14800,N_12118);
xor U16765 (N_16765,N_11527,N_10918);
nand U16766 (N_16766,N_10603,N_11122);
or U16767 (N_16767,N_14300,N_10694);
nand U16768 (N_16768,N_13713,N_12040);
nand U16769 (N_16769,N_11605,N_13456);
or U16770 (N_16770,N_13217,N_12382);
nand U16771 (N_16771,N_13174,N_11546);
and U16772 (N_16772,N_12867,N_13051);
xnor U16773 (N_16773,N_12519,N_10581);
xnor U16774 (N_16774,N_12908,N_11958);
xnor U16775 (N_16775,N_12229,N_13106);
or U16776 (N_16776,N_14858,N_13416);
and U16777 (N_16777,N_10087,N_10401);
or U16778 (N_16778,N_10942,N_12430);
nand U16779 (N_16779,N_11014,N_11663);
or U16780 (N_16780,N_13160,N_10069);
nand U16781 (N_16781,N_10245,N_13652);
and U16782 (N_16782,N_12169,N_13248);
xor U16783 (N_16783,N_14278,N_11670);
nor U16784 (N_16784,N_14155,N_11757);
nand U16785 (N_16785,N_13436,N_12923);
and U16786 (N_16786,N_11629,N_10477);
or U16787 (N_16787,N_14403,N_11093);
nand U16788 (N_16788,N_14404,N_10742);
and U16789 (N_16789,N_10558,N_13485);
xnor U16790 (N_16790,N_11071,N_11206);
xnor U16791 (N_16791,N_12110,N_14575);
nand U16792 (N_16792,N_10492,N_10075);
nand U16793 (N_16793,N_12649,N_12495);
xnor U16794 (N_16794,N_12043,N_11484);
nand U16795 (N_16795,N_10385,N_12155);
nand U16796 (N_16796,N_12177,N_10379);
and U16797 (N_16797,N_12281,N_14813);
nor U16798 (N_16798,N_14367,N_10417);
nand U16799 (N_16799,N_12074,N_10304);
nor U16800 (N_16800,N_10026,N_10637);
xor U16801 (N_16801,N_13520,N_13419);
xor U16802 (N_16802,N_12937,N_14060);
nand U16803 (N_16803,N_11207,N_14181);
or U16804 (N_16804,N_10977,N_14136);
nor U16805 (N_16805,N_11212,N_11125);
or U16806 (N_16806,N_13289,N_11959);
xnor U16807 (N_16807,N_14975,N_11406);
and U16808 (N_16808,N_12936,N_12633);
nand U16809 (N_16809,N_14044,N_10097);
and U16810 (N_16810,N_13751,N_11091);
and U16811 (N_16811,N_11994,N_13521);
nand U16812 (N_16812,N_11105,N_12566);
nor U16813 (N_16813,N_13731,N_11150);
or U16814 (N_16814,N_14145,N_13993);
or U16815 (N_16815,N_12042,N_10754);
nor U16816 (N_16816,N_11945,N_12769);
xor U16817 (N_16817,N_14797,N_14928);
xnor U16818 (N_16818,N_10374,N_12045);
nor U16819 (N_16819,N_13278,N_13632);
or U16820 (N_16820,N_12089,N_14754);
or U16821 (N_16821,N_10005,N_12008);
and U16822 (N_16822,N_10577,N_12631);
xnor U16823 (N_16823,N_14105,N_14066);
nand U16824 (N_16824,N_11827,N_10425);
and U16825 (N_16825,N_12839,N_10550);
or U16826 (N_16826,N_12077,N_13948);
xor U16827 (N_16827,N_11517,N_10279);
or U16828 (N_16828,N_12724,N_10032);
xnor U16829 (N_16829,N_11328,N_12385);
or U16830 (N_16830,N_10451,N_10708);
nand U16831 (N_16831,N_13404,N_11465);
or U16832 (N_16832,N_12262,N_14395);
nor U16833 (N_16833,N_12137,N_12404);
xnor U16834 (N_16834,N_12214,N_10513);
nor U16835 (N_16835,N_14709,N_10312);
and U16836 (N_16836,N_11993,N_12617);
xnor U16837 (N_16837,N_12706,N_11610);
xnor U16838 (N_16838,N_12316,N_14749);
nor U16839 (N_16839,N_14074,N_12296);
and U16840 (N_16840,N_11480,N_14068);
nand U16841 (N_16841,N_12436,N_13550);
or U16842 (N_16842,N_12577,N_11525);
xor U16843 (N_16843,N_12246,N_13031);
xnor U16844 (N_16844,N_11354,N_12123);
and U16845 (N_16845,N_13512,N_12907);
and U16846 (N_16846,N_14027,N_13371);
and U16847 (N_16847,N_11743,N_14132);
nor U16848 (N_16848,N_12641,N_11604);
xor U16849 (N_16849,N_10056,N_14536);
and U16850 (N_16850,N_11025,N_10382);
nor U16851 (N_16851,N_11132,N_10973);
xor U16852 (N_16852,N_11190,N_10843);
or U16853 (N_16853,N_11919,N_11177);
or U16854 (N_16854,N_10413,N_11651);
nand U16855 (N_16855,N_12162,N_13441);
or U16856 (N_16856,N_12722,N_12443);
xnor U16857 (N_16857,N_10306,N_13781);
xor U16858 (N_16858,N_13410,N_10479);
or U16859 (N_16859,N_11592,N_13487);
and U16860 (N_16860,N_12375,N_14647);
nor U16861 (N_16861,N_12665,N_14812);
and U16862 (N_16862,N_10514,N_14588);
or U16863 (N_16863,N_11548,N_13452);
nand U16864 (N_16864,N_10925,N_12124);
nor U16865 (N_16865,N_13590,N_13065);
or U16866 (N_16866,N_14023,N_11250);
or U16867 (N_16867,N_12472,N_11901);
or U16868 (N_16868,N_10464,N_11776);
nand U16869 (N_16869,N_14729,N_14991);
nand U16870 (N_16870,N_14885,N_11879);
xnor U16871 (N_16871,N_10130,N_11709);
or U16872 (N_16872,N_11535,N_13738);
xnor U16873 (N_16873,N_10373,N_13270);
nor U16874 (N_16874,N_13179,N_14561);
or U16875 (N_16875,N_12949,N_14016);
and U16876 (N_16876,N_11325,N_13027);
nor U16877 (N_16877,N_12086,N_10394);
xnor U16878 (N_16878,N_11979,N_10687);
xnor U16879 (N_16879,N_10490,N_10397);
and U16880 (N_16880,N_12999,N_12740);
xnor U16881 (N_16881,N_12914,N_12586);
nand U16882 (N_16882,N_10870,N_14093);
or U16883 (N_16883,N_14024,N_10724);
nand U16884 (N_16884,N_13246,N_10129);
nor U16885 (N_16885,N_13900,N_14073);
nor U16886 (N_16886,N_12522,N_14780);
nand U16887 (N_16887,N_10123,N_11400);
or U16888 (N_16888,N_10496,N_11857);
and U16889 (N_16889,N_12616,N_10282);
nor U16890 (N_16890,N_10562,N_13262);
nand U16891 (N_16891,N_14893,N_14648);
nor U16892 (N_16892,N_10463,N_13533);
xnor U16893 (N_16893,N_11589,N_14018);
or U16894 (N_16894,N_10423,N_12061);
and U16895 (N_16895,N_13071,N_11526);
nand U16896 (N_16896,N_14894,N_11296);
xor U16897 (N_16897,N_11777,N_13198);
nand U16898 (N_16898,N_10183,N_14444);
xor U16899 (N_16899,N_14637,N_11796);
and U16900 (N_16900,N_10957,N_14656);
and U16901 (N_16901,N_13192,N_11702);
nand U16902 (N_16902,N_13505,N_12557);
and U16903 (N_16903,N_12940,N_10260);
nor U16904 (N_16904,N_12483,N_12782);
nor U16905 (N_16905,N_13523,N_11419);
and U16906 (N_16906,N_12904,N_14341);
and U16907 (N_16907,N_13238,N_12325);
nor U16908 (N_16908,N_10449,N_14531);
nand U16909 (N_16909,N_13308,N_12801);
and U16910 (N_16910,N_14849,N_11649);
xor U16911 (N_16911,N_14756,N_11104);
and U16912 (N_16912,N_12728,N_12173);
nand U16913 (N_16913,N_11393,N_13005);
nand U16914 (N_16914,N_12915,N_13831);
xnor U16915 (N_16915,N_13094,N_12075);
nand U16916 (N_16916,N_11282,N_10188);
xor U16917 (N_16917,N_11140,N_14876);
or U16918 (N_16918,N_14189,N_11855);
xor U16919 (N_16919,N_13142,N_13739);
and U16920 (N_16920,N_10924,N_14681);
nand U16921 (N_16921,N_13658,N_13903);
xor U16922 (N_16922,N_14178,N_14264);
nor U16923 (N_16923,N_12675,N_12638);
and U16924 (N_16924,N_13804,N_14475);
nor U16925 (N_16925,N_12735,N_11785);
xnor U16926 (N_16926,N_13576,N_14213);
xnor U16927 (N_16927,N_11062,N_12399);
or U16928 (N_16928,N_12698,N_14158);
and U16929 (N_16929,N_14092,N_11390);
and U16930 (N_16930,N_14430,N_14807);
or U16931 (N_16931,N_13175,N_13673);
nand U16932 (N_16932,N_12342,N_14147);
xnor U16933 (N_16933,N_10002,N_10285);
nand U16934 (N_16934,N_14095,N_12267);
nand U16935 (N_16935,N_11823,N_11005);
xor U16936 (N_16936,N_14339,N_13980);
nor U16937 (N_16937,N_11124,N_12546);
nor U16938 (N_16938,N_13313,N_13859);
nor U16939 (N_16939,N_12536,N_10091);
and U16940 (N_16940,N_10636,N_10551);
or U16941 (N_16941,N_11249,N_10955);
and U16942 (N_16942,N_14916,N_12455);
xnor U16943 (N_16943,N_13813,N_11916);
and U16944 (N_16944,N_11117,N_14225);
or U16945 (N_16945,N_14515,N_10235);
and U16946 (N_16946,N_13233,N_14316);
nor U16947 (N_16947,N_10896,N_13502);
nand U16948 (N_16948,N_13435,N_12494);
xnor U16949 (N_16949,N_10406,N_11483);
xor U16950 (N_16950,N_14590,N_10469);
and U16951 (N_16951,N_13730,N_14938);
and U16952 (N_16952,N_12659,N_11924);
and U16953 (N_16953,N_14939,N_10214);
nor U16954 (N_16954,N_14600,N_14449);
nand U16955 (N_16955,N_11606,N_13878);
nor U16956 (N_16956,N_11771,N_12454);
and U16957 (N_16957,N_13987,N_13151);
nor U16958 (N_16958,N_14795,N_14243);
nand U16959 (N_16959,N_14234,N_12166);
nor U16960 (N_16960,N_13181,N_12544);
and U16961 (N_16961,N_12393,N_13103);
or U16962 (N_16962,N_14570,N_10012);
nand U16963 (N_16963,N_13393,N_13290);
or U16964 (N_16964,N_10178,N_12738);
nand U16965 (N_16965,N_14398,N_13942);
nand U16966 (N_16966,N_13789,N_10690);
and U16967 (N_16967,N_10107,N_12593);
nor U16968 (N_16968,N_14623,N_11297);
nand U16969 (N_16969,N_12036,N_11486);
or U16970 (N_16970,N_10225,N_14578);
nand U16971 (N_16971,N_14154,N_10766);
nand U16972 (N_16972,N_12560,N_10237);
nand U16973 (N_16973,N_11868,N_10546);
and U16974 (N_16974,N_12319,N_13235);
nand U16975 (N_16975,N_12332,N_12618);
xor U16976 (N_16976,N_12596,N_13099);
xor U16977 (N_16977,N_11566,N_13400);
and U16978 (N_16978,N_10045,N_14726);
or U16979 (N_16979,N_13164,N_12198);
or U16980 (N_16980,N_10635,N_11451);
and U16981 (N_16981,N_10660,N_13527);
and U16982 (N_16982,N_12819,N_10234);
xor U16983 (N_16983,N_13280,N_14423);
nand U16984 (N_16984,N_13347,N_14935);
xnor U16985 (N_16985,N_10799,N_14005);
or U16986 (N_16986,N_13331,N_12768);
or U16987 (N_16987,N_11533,N_14649);
nand U16988 (N_16988,N_13064,N_11964);
and U16989 (N_16989,N_10278,N_13225);
or U16990 (N_16990,N_14064,N_14999);
nor U16991 (N_16991,N_12863,N_12083);
or U16992 (N_16992,N_11599,N_11379);
xnor U16993 (N_16993,N_11381,N_12674);
or U16994 (N_16994,N_10929,N_14488);
or U16995 (N_16995,N_11892,N_10872);
nor U16996 (N_16996,N_11098,N_14765);
nor U16997 (N_16997,N_12265,N_14989);
xor U16998 (N_16998,N_11032,N_12715);
and U16999 (N_16999,N_10976,N_13355);
or U17000 (N_17000,N_10432,N_13977);
or U17001 (N_17001,N_12444,N_13618);
nor U17002 (N_17002,N_14962,N_11755);
nand U17003 (N_17003,N_13578,N_11818);
xor U17004 (N_17004,N_14804,N_14946);
and U17005 (N_17005,N_12767,N_12463);
or U17006 (N_17006,N_12416,N_13734);
xnor U17007 (N_17007,N_11278,N_12047);
xor U17008 (N_17008,N_12141,N_13318);
nor U17009 (N_17009,N_14932,N_13906);
xor U17010 (N_17010,N_11543,N_11862);
xnor U17011 (N_17011,N_14035,N_13634);
or U17012 (N_17012,N_12225,N_10967);
or U17013 (N_17013,N_13997,N_11813);
nand U17014 (N_17014,N_11594,N_10650);
xnor U17015 (N_17015,N_12426,N_13309);
xor U17016 (N_17016,N_12979,N_14696);
and U17017 (N_17017,N_11768,N_12773);
or U17018 (N_17018,N_13967,N_14317);
and U17019 (N_17019,N_12299,N_13186);
nand U17020 (N_17020,N_10676,N_13598);
and U17021 (N_17021,N_14692,N_10362);
nand U17022 (N_17022,N_13020,N_14657);
nor U17023 (N_17023,N_14441,N_10209);
or U17024 (N_17024,N_13753,N_14257);
nor U17025 (N_17025,N_13470,N_14512);
nor U17026 (N_17026,N_11281,N_10608);
nor U17027 (N_17027,N_10667,N_12421);
nor U17028 (N_17028,N_14301,N_10043);
nand U17029 (N_17029,N_10029,N_10684);
nor U17030 (N_17030,N_13474,N_11986);
nand U17031 (N_17031,N_12766,N_14565);
or U17032 (N_17032,N_12732,N_13132);
nand U17033 (N_17033,N_11057,N_13936);
xor U17034 (N_17034,N_11659,N_11002);
nand U17035 (N_17035,N_11809,N_13069);
nor U17036 (N_17036,N_12532,N_14443);
xnor U17037 (N_17037,N_10547,N_11171);
and U17038 (N_17038,N_14450,N_14730);
or U17039 (N_17039,N_14626,N_10933);
nor U17040 (N_17040,N_14820,N_11899);
xnor U17041 (N_17041,N_12250,N_12734);
nor U17042 (N_17042,N_10182,N_14834);
and U17043 (N_17043,N_14605,N_11633);
nand U17044 (N_17044,N_12518,N_10412);
xnor U17045 (N_17045,N_12488,N_10753);
nand U17046 (N_17046,N_13935,N_12312);
or U17047 (N_17047,N_13388,N_12945);
and U17048 (N_17048,N_10750,N_11218);
nor U17049 (N_17049,N_13168,N_10452);
nand U17050 (N_17050,N_11226,N_10491);
or U17051 (N_17051,N_11128,N_10822);
xor U17052 (N_17052,N_11747,N_13498);
nor U17053 (N_17053,N_14713,N_10732);
and U17054 (N_17054,N_10131,N_10361);
nand U17055 (N_17055,N_10484,N_13121);
nand U17056 (N_17056,N_10619,N_11130);
and U17057 (N_17057,N_12591,N_13411);
nor U17058 (N_17058,N_12542,N_10329);
xor U17059 (N_17059,N_13566,N_11363);
xnor U17060 (N_17060,N_10420,N_14109);
nand U17061 (N_17061,N_11414,N_11653);
nand U17062 (N_17062,N_10960,N_14185);
nand U17063 (N_17063,N_13222,N_14556);
nand U17064 (N_17064,N_14124,N_12441);
nand U17065 (N_17065,N_11367,N_14658);
xor U17066 (N_17066,N_12489,N_14174);
nand U17067 (N_17067,N_14677,N_14603);
and U17068 (N_17068,N_13725,N_14348);
and U17069 (N_17069,N_13701,N_10590);
nand U17070 (N_17070,N_10150,N_13477);
nand U17071 (N_17071,N_12998,N_12187);
xor U17072 (N_17072,N_13824,N_13158);
nand U17073 (N_17073,N_12130,N_14970);
and U17074 (N_17074,N_14326,N_14580);
nor U17075 (N_17075,N_11980,N_10845);
and U17076 (N_17076,N_12707,N_12150);
nor U17077 (N_17077,N_10305,N_12850);
and U17078 (N_17078,N_10486,N_13591);
or U17079 (N_17079,N_11371,N_10331);
or U17080 (N_17080,N_14902,N_10605);
or U17081 (N_17081,N_12027,N_14120);
nand U17082 (N_17082,N_10971,N_12301);
nor U17083 (N_17083,N_13282,N_14500);
and U17084 (N_17084,N_12985,N_12314);
nand U17085 (N_17085,N_14951,N_10502);
or U17086 (N_17086,N_12233,N_11643);
and U17087 (N_17087,N_13025,N_10219);
nand U17088 (N_17088,N_12059,N_11682);
nor U17089 (N_17089,N_11922,N_10840);
and U17090 (N_17090,N_14416,N_10835);
or U17091 (N_17091,N_13979,N_14625);
xnor U17092 (N_17092,N_10369,N_14917);
xor U17093 (N_17093,N_14513,N_11705);
nor U17094 (N_17094,N_13709,N_11744);
nand U17095 (N_17095,N_14573,N_12015);
xor U17096 (N_17096,N_10946,N_11627);
nor U17097 (N_17097,N_10468,N_14102);
and U17098 (N_17098,N_14863,N_13594);
or U17099 (N_17099,N_11470,N_12097);
xnor U17100 (N_17100,N_10171,N_10868);
and U17101 (N_17101,N_14038,N_11489);
xnor U17102 (N_17102,N_13914,N_11799);
and U17103 (N_17103,N_14913,N_10061);
xor U17104 (N_17104,N_14882,N_12412);
xor U17105 (N_17105,N_11202,N_14346);
nand U17106 (N_17106,N_13798,N_10852);
xor U17107 (N_17107,N_13722,N_12826);
nor U17108 (N_17108,N_11805,N_10286);
xor U17109 (N_17109,N_12930,N_13708);
nand U17110 (N_17110,N_10519,N_13014);
nand U17111 (N_17111,N_10906,N_12808);
xor U17112 (N_17112,N_11413,N_12957);
nand U17113 (N_17113,N_13648,N_13415);
or U17114 (N_17114,N_12651,N_13274);
xnor U17115 (N_17115,N_10989,N_13294);
or U17116 (N_17116,N_14979,N_11692);
nor U17117 (N_17117,N_10733,N_12115);
and U17118 (N_17118,N_11087,N_12545);
nand U17119 (N_17119,N_13266,N_12946);
xnor U17120 (N_17120,N_13059,N_14429);
nand U17121 (N_17121,N_11991,N_10232);
nor U17122 (N_17122,N_12938,N_12476);
or U17123 (N_17123,N_10782,N_14595);
or U17124 (N_17124,N_11529,N_13530);
and U17125 (N_17125,N_12140,N_14599);
and U17126 (N_17126,N_14883,N_14218);
xor U17127 (N_17127,N_10699,N_12152);
or U17128 (N_17128,N_13780,N_11700);
nor U17129 (N_17129,N_12484,N_12276);
nand U17130 (N_17130,N_12513,N_13842);
nand U17131 (N_17131,N_14520,N_12231);
nand U17132 (N_17132,N_14822,N_10769);
xor U17133 (N_17133,N_14411,N_13570);
or U17134 (N_17134,N_10600,N_10082);
and U17135 (N_17135,N_13276,N_10114);
and U17136 (N_17136,N_10787,N_14818);
nor U17137 (N_17137,N_13605,N_11802);
nor U17138 (N_17138,N_13794,N_14710);
and U17139 (N_17139,N_10474,N_13265);
and U17140 (N_17140,N_13391,N_11790);
and U17141 (N_17141,N_11155,N_12661);
xor U17142 (N_17142,N_14722,N_14723);
and U17143 (N_17143,N_13840,N_14029);
or U17144 (N_17144,N_12678,N_14889);
nand U17145 (N_17145,N_12978,N_10861);
or U17146 (N_17146,N_12044,N_14949);
or U17147 (N_17147,N_10000,N_10673);
nand U17148 (N_17148,N_10847,N_13214);
or U17149 (N_17149,N_14751,N_11810);
or U17150 (N_17150,N_14057,N_12521);
nor U17151 (N_17151,N_12235,N_11341);
xor U17152 (N_17152,N_11551,N_13272);
nand U17153 (N_17153,N_11967,N_12932);
and U17154 (N_17154,N_11086,N_10654);
and U17155 (N_17155,N_12538,N_13484);
nand U17156 (N_17156,N_13122,N_10195);
and U17157 (N_17157,N_12132,N_13424);
nor U17158 (N_17158,N_12351,N_11047);
and U17159 (N_17159,N_13978,N_12372);
xnor U17160 (N_17160,N_14270,N_11411);
or U17161 (N_17161,N_10207,N_14548);
xnor U17162 (N_17162,N_13923,N_10041);
or U17163 (N_17163,N_11801,N_14034);
nor U17164 (N_17164,N_14407,N_12922);
nand U17165 (N_17165,N_11211,N_11056);
nor U17166 (N_17166,N_11721,N_10148);
or U17167 (N_17167,N_12343,N_11166);
and U17168 (N_17168,N_14879,N_10354);
nor U17169 (N_17169,N_10503,N_13021);
xnor U17170 (N_17170,N_13169,N_13352);
nor U17171 (N_17171,N_10333,N_13588);
xnor U17172 (N_17172,N_12713,N_13397);
xor U17173 (N_17173,N_12405,N_11628);
or U17174 (N_17174,N_10735,N_14077);
and U17175 (N_17175,N_11582,N_12832);
and U17176 (N_17176,N_13255,N_13665);
nor U17177 (N_17177,N_11230,N_13440);
and U17178 (N_17178,N_13981,N_10193);
nand U17179 (N_17179,N_13705,N_13324);
xnor U17180 (N_17180,N_14438,N_14004);
or U17181 (N_17181,N_12278,N_13045);
or U17182 (N_17182,N_14745,N_14552);
nand U17183 (N_17183,N_12600,N_14759);
nand U17184 (N_17184,N_10618,N_11417);
nor U17185 (N_17185,N_10428,N_10534);
or U17186 (N_17186,N_10731,N_12226);
nand U17187 (N_17187,N_12462,N_11836);
nand U17188 (N_17188,N_12514,N_11336);
or U17189 (N_17189,N_10511,N_10748);
nor U17190 (N_17190,N_13846,N_13314);
or U17191 (N_17191,N_14838,N_12869);
and U17192 (N_17192,N_11559,N_10838);
xnor U17193 (N_17193,N_12082,N_14146);
xnor U17194 (N_17194,N_11170,N_10457);
or U17195 (N_17195,N_11433,N_13822);
and U17196 (N_17196,N_10961,N_14968);
or U17197 (N_17197,N_13558,N_11961);
nand U17198 (N_17198,N_11275,N_10038);
nor U17199 (N_17199,N_12168,N_14631);
nand U17200 (N_17200,N_13471,N_10116);
xor U17201 (N_17201,N_14465,N_11455);
or U17202 (N_17202,N_12330,N_12900);
nand U17203 (N_17203,N_11101,N_13104);
xor U17204 (N_17204,N_12916,N_13873);
nor U17205 (N_17205,N_13127,N_12750);
or U17206 (N_17206,N_14428,N_11637);
nor U17207 (N_17207,N_10414,N_10015);
xnor U17208 (N_17208,N_13478,N_11081);
nand U17209 (N_17209,N_13119,N_12860);
nand U17210 (N_17210,N_12176,N_11941);
nor U17211 (N_17211,N_14557,N_11712);
or U17212 (N_17212,N_11276,N_11069);
xnor U17213 (N_17213,N_11051,N_13201);
or U17214 (N_17214,N_12464,N_11557);
nor U17215 (N_17215,N_12933,N_14620);
nand U17216 (N_17216,N_10126,N_11724);
xor U17217 (N_17217,N_12778,N_11830);
nand U17218 (N_17218,N_14373,N_11787);
and U17219 (N_17219,N_13450,N_12411);
nand U17220 (N_17220,N_11332,N_12626);
nand U17221 (N_17221,N_13852,N_12091);
and U17222 (N_17222,N_10830,N_12425);
xnor U17223 (N_17223,N_14363,N_10006);
and U17224 (N_17224,N_14796,N_14127);
nor U17225 (N_17225,N_14667,N_13501);
and U17226 (N_17226,N_10947,N_14076);
and U17227 (N_17227,N_12010,N_14356);
and U17228 (N_17228,N_14277,N_11542);
nor U17229 (N_17229,N_14693,N_11900);
xor U17230 (N_17230,N_10901,N_13319);
nand U17231 (N_17231,N_11504,N_12378);
nand U17232 (N_17232,N_14744,N_14457);
nand U17233 (N_17233,N_11388,N_12595);
or U17234 (N_17234,N_10339,N_10196);
nor U17235 (N_17235,N_13310,N_14871);
nand U17236 (N_17236,N_12551,N_12840);
nand U17237 (N_17237,N_14231,N_12458);
nor U17238 (N_17238,N_13999,N_13931);
or U17239 (N_17239,N_13446,N_12531);
nor U17240 (N_17240,N_13057,N_11842);
nor U17241 (N_17241,N_13577,N_11270);
or U17242 (N_17242,N_10934,N_10088);
xnor U17243 (N_17243,N_11327,N_13572);
xnor U17244 (N_17244,N_11646,N_14453);
nand U17245 (N_17245,N_13868,N_11307);
nand U17246 (N_17246,N_14229,N_11410);
nor U17247 (N_17247,N_10686,N_10980);
or U17248 (N_17248,N_14770,N_14362);
and U17249 (N_17249,N_11881,N_10074);
xnor U17250 (N_17250,N_14017,N_14205);
or U17251 (N_17251,N_14790,N_10121);
xnor U17252 (N_17252,N_11468,N_12456);
or U17253 (N_17253,N_13124,N_13792);
or U17254 (N_17254,N_10663,N_10105);
and U17255 (N_17255,N_13332,N_12088);
xnor U17256 (N_17256,N_14862,N_10810);
or U17257 (N_17257,N_10018,N_13467);
xnor U17258 (N_17258,N_10985,N_14836);
or U17259 (N_17259,N_13638,N_12958);
nand U17260 (N_17260,N_10199,N_10927);
nand U17261 (N_17261,N_12975,N_13296);
or U17262 (N_17262,N_14466,N_13974);
or U17263 (N_17263,N_14121,N_10060);
and U17264 (N_17264,N_11272,N_13541);
and U17265 (N_17265,N_11640,N_10691);
xor U17266 (N_17266,N_11645,N_13559);
nand U17267 (N_17267,N_14082,N_14190);
or U17268 (N_17268,N_12473,N_11740);
or U17269 (N_17269,N_10485,N_10179);
nor U17270 (N_17270,N_13430,N_13423);
and U17271 (N_17271,N_13757,N_10247);
nand U17272 (N_17272,N_10816,N_10797);
and U17273 (N_17273,N_12905,N_13863);
and U17274 (N_17274,N_11846,N_11095);
and U17275 (N_17275,N_12627,N_10701);
nor U17276 (N_17276,N_12038,N_14680);
nand U17277 (N_17277,N_10034,N_10549);
nor U17278 (N_17278,N_14405,N_14563);
and U17279 (N_17279,N_13943,N_12868);
nor U17280 (N_17280,N_13791,N_13368);
nor U17281 (N_17281,N_10327,N_11839);
and U17282 (N_17282,N_11735,N_13747);
or U17283 (N_17283,N_14090,N_12390);
and U17284 (N_17284,N_13348,N_10669);
nand U17285 (N_17285,N_11886,N_13247);
and U17286 (N_17286,N_12409,N_10264);
xor U17287 (N_17287,N_14347,N_11213);
nor U17288 (N_17288,N_11009,N_14456);
nor U17289 (N_17289,N_13884,N_11603);
or U17290 (N_17290,N_13399,N_13957);
or U17291 (N_17291,N_14409,N_12433);
nand U17292 (N_17292,N_11615,N_13086);
or U17293 (N_17293,N_10903,N_10695);
nor U17294 (N_17294,N_13293,N_14002);
nand U17295 (N_17295,N_11972,N_13162);
nor U17296 (N_17296,N_12174,N_10334);
or U17297 (N_17297,N_13645,N_11458);
xor U17298 (N_17298,N_10067,N_10248);
xnor U17299 (N_17299,N_12438,N_10885);
nand U17300 (N_17300,N_10593,N_11884);
and U17301 (N_17301,N_10283,N_14772);
and U17302 (N_17302,N_11208,N_10238);
xor U17303 (N_17303,N_11607,N_14927);
nand U17304 (N_17304,N_10112,N_12847);
xnor U17305 (N_17305,N_12823,N_12643);
nand U17306 (N_17306,N_12656,N_14113);
and U17307 (N_17307,N_12663,N_10086);
or U17308 (N_17308,N_14504,N_14995);
xor U17309 (N_17309,N_11333,N_11268);
and U17310 (N_17310,N_14773,N_11571);
or U17311 (N_17311,N_11650,N_14864);
nand U17312 (N_17312,N_14447,N_10431);
xor U17313 (N_17313,N_13534,N_14758);
and U17314 (N_17314,N_12011,N_14622);
xnor U17315 (N_17315,N_13184,N_12582);
nor U17316 (N_17316,N_11365,N_12210);
nand U17317 (N_17317,N_11337,N_12360);
and U17318 (N_17318,N_14011,N_14485);
nor U17319 (N_17319,N_11068,N_14118);
nand U17320 (N_17320,N_11786,N_12211);
nor U17321 (N_17321,N_10202,N_14307);
nor U17322 (N_17322,N_13659,N_13564);
nand U17323 (N_17323,N_11000,N_11185);
and U17324 (N_17324,N_12335,N_12703);
xnor U17325 (N_17325,N_11291,N_11262);
xnor U17326 (N_17326,N_12549,N_14844);
xor U17327 (N_17327,N_12171,N_11734);
nor U17328 (N_17328,N_13438,N_10610);
nand U17329 (N_17329,N_11499,N_14767);
and U17330 (N_17330,N_13767,N_12835);
or U17331 (N_17331,N_12499,N_10940);
and U17332 (N_17332,N_11046,N_10710);
and U17333 (N_17333,N_10101,N_10849);
or U17334 (N_17334,N_14188,N_14151);
nor U17335 (N_17335,N_10949,N_10520);
xnor U17336 (N_17336,N_14055,N_14388);
or U17337 (N_17337,N_10111,N_12251);
nand U17338 (N_17338,N_13312,N_11142);
or U17339 (N_17339,N_10749,N_14524);
nor U17340 (N_17340,N_10905,N_12054);
and U17341 (N_17341,N_10161,N_12147);
xor U17342 (N_17342,N_12356,N_11995);
or U17343 (N_17343,N_10809,N_13492);
nand U17344 (N_17344,N_11626,N_14445);
or U17345 (N_17345,N_11949,N_11195);
and U17346 (N_17346,N_11639,N_12308);
nand U17347 (N_17347,N_12364,N_13034);
or U17348 (N_17348,N_13087,N_13971);
nand U17349 (N_17349,N_10999,N_12962);
and U17350 (N_17350,N_11007,N_13061);
and U17351 (N_17351,N_10165,N_11089);
or U17352 (N_17352,N_13136,N_14321);
xor U17353 (N_17353,N_11096,N_10530);
xor U17354 (N_17354,N_11391,N_10422);
and U17355 (N_17355,N_12467,N_12402);
and U17356 (N_17356,N_14806,N_13716);
and U17357 (N_17357,N_11119,N_11952);
nor U17358 (N_17358,N_10410,N_10824);
and U17359 (N_17359,N_10284,N_10765);
xor U17360 (N_17360,N_11435,N_11267);
and U17361 (N_17361,N_13827,N_10923);
xnor U17362 (N_17362,N_14084,N_12660);
or U17363 (N_17363,N_12212,N_11828);
or U17364 (N_17364,N_10246,N_11067);
and U17365 (N_17365,N_14319,N_11495);
xnor U17366 (N_17366,N_13679,N_12024);
xnor U17367 (N_17367,N_10826,N_14613);
or U17368 (N_17368,N_10411,N_13620);
nor U17369 (N_17369,N_10675,N_10779);
or U17370 (N_17370,N_11329,N_14330);
xnor U17371 (N_17371,N_14461,N_11519);
xor U17372 (N_17372,N_10198,N_14203);
or U17373 (N_17373,N_14567,N_13196);
or U17374 (N_17374,N_10979,N_13553);
and U17375 (N_17375,N_14381,N_13772);
nand U17376 (N_17376,N_13775,N_13829);
nand U17377 (N_17377,N_11585,N_10739);
nor U17378 (N_17378,N_10553,N_14930);
and U17379 (N_17379,N_10399,N_12680);
xnor U17380 (N_17380,N_12202,N_11808);
or U17381 (N_17381,N_13837,N_11987);
xnor U17382 (N_17382,N_10062,N_10055);
xnor U17383 (N_17383,N_10796,N_13080);
nor U17384 (N_17384,N_14839,N_11950);
or U17385 (N_17385,N_10221,N_11641);
and U17386 (N_17386,N_10288,N_12995);
and U17387 (N_17387,N_12510,N_10236);
nor U17388 (N_17388,N_11797,N_10025);
nand U17389 (N_17389,N_10313,N_11885);
and U17390 (N_17390,N_13696,N_10997);
nand U17391 (N_17391,N_14083,N_11717);
and U17392 (N_17392,N_11547,N_11023);
nand U17393 (N_17393,N_12741,N_12078);
nor U17394 (N_17394,N_10155,N_12968);
nor U17395 (N_17395,N_10364,N_14685);
nor U17396 (N_17396,N_10337,N_12955);
nand U17397 (N_17397,N_11235,N_13503);
xor U17398 (N_17398,N_12060,N_10755);
nor U17399 (N_17399,N_12744,N_13698);
or U17400 (N_17400,N_12057,N_11044);
or U17401 (N_17401,N_10347,N_13062);
xor U17402 (N_17402,N_13996,N_10172);
nor U17403 (N_17403,N_10266,N_12079);
and U17404 (N_17404,N_13195,N_12427);
and U17405 (N_17405,N_10889,N_13596);
nand U17406 (N_17406,N_11518,N_11040);
or U17407 (N_17407,N_12983,N_14959);
and U17408 (N_17408,N_10152,N_12870);
nand U17409 (N_17409,N_13955,N_10679);
nor U17410 (N_17410,N_11351,N_13437);
and U17411 (N_17411,N_10798,N_12762);
and U17412 (N_17412,N_14926,N_12453);
nor U17413 (N_17413,N_12589,N_12158);
xor U17414 (N_17414,N_14614,N_12144);
nor U17415 (N_17415,N_14126,N_11563);
nor U17416 (N_17416,N_11346,N_14391);
nor U17417 (N_17417,N_14378,N_11781);
or U17418 (N_17418,N_12528,N_14974);
nor U17419 (N_17419,N_12774,N_11677);
and U17420 (N_17420,N_10587,N_11920);
and U17421 (N_17421,N_12014,N_13956);
nand U17422 (N_17422,N_10532,N_13337);
nor U17423 (N_17423,N_11156,N_12584);
xnor U17424 (N_17424,N_11847,N_13161);
xnor U17425 (N_17425,N_10104,N_11472);
nor U17426 (N_17426,N_12080,N_11045);
nand U17427 (N_17427,N_11209,N_10808);
and U17428 (N_17428,N_12650,N_12730);
nor U17429 (N_17429,N_11456,N_13024);
nor U17430 (N_17430,N_11729,N_13557);
nor U17431 (N_17431,N_13082,N_12223);
and U17432 (N_17432,N_11436,N_13628);
nor U17433 (N_17433,N_13345,N_14571);
nand U17434 (N_17434,N_13524,N_10180);
and U17435 (N_17435,N_12815,N_10879);
nand U17436 (N_17436,N_10118,N_13493);
or U17437 (N_17437,N_13675,N_10536);
nor U17438 (N_17438,N_12776,N_12228);
xnor U17439 (N_17439,N_12058,N_14420);
nand U17440 (N_17440,N_13407,N_10604);
nand U17441 (N_17441,N_13167,N_11596);
nor U17442 (N_17442,N_12023,N_10688);
and U17443 (N_17443,N_12729,N_12275);
or U17444 (N_17444,N_12974,N_13090);
nor U17445 (N_17445,N_10800,N_13153);
nand U17446 (N_17446,N_11369,N_13026);
xor U17447 (N_17447,N_12711,N_14393);
nor U17448 (N_17448,N_12889,N_10853);
or U17449 (N_17449,N_10956,N_10344);
or U17450 (N_17450,N_11076,N_13778);
xnor U17451 (N_17451,N_13581,N_10680);
and U17452 (N_17452,N_13461,N_13556);
nor U17453 (N_17453,N_14477,N_12282);
or U17454 (N_17454,N_13547,N_13053);
and U17455 (N_17455,N_14687,N_12973);
xor U17456 (N_17456,N_12445,N_10071);
and U17457 (N_17457,N_10855,N_13428);
nor U17458 (N_17458,N_12959,N_10185);
and U17459 (N_17459,N_12709,N_10529);
xnor U17460 (N_17460,N_13078,N_12632);
and U17461 (N_17461,N_14000,N_12095);
or U17462 (N_17462,N_12972,N_12601);
xor U17463 (N_17463,N_13664,N_10591);
or U17464 (N_17464,N_10070,N_14139);
and U17465 (N_17465,N_13908,N_14111);
xor U17466 (N_17466,N_12327,N_12576);
nand U17467 (N_17467,N_11618,N_14684);
or U17468 (N_17468,N_10119,N_12793);
nor U17469 (N_17469,N_14717,N_11467);
and U17470 (N_17470,N_10052,N_14259);
xnor U17471 (N_17471,N_10606,N_12657);
or U17472 (N_17472,N_12954,N_12624);
or U17473 (N_17473,N_11505,N_12986);
nand U17474 (N_17474,N_11766,N_11475);
or U17475 (N_17475,N_10936,N_12334);
or U17476 (N_17476,N_13287,N_13754);
nor U17477 (N_17477,N_14182,N_13925);
xor U17478 (N_17478,N_10044,N_11357);
xor U17479 (N_17479,N_10563,N_12717);
or U17480 (N_17480,N_12067,N_12305);
xor U17481 (N_17481,N_10584,N_12783);
xor U17482 (N_17482,N_14331,N_13742);
nand U17483 (N_17483,N_10613,N_10875);
nand U17484 (N_17484,N_11194,N_12069);
and U17485 (N_17485,N_14258,N_10598);
nor U17486 (N_17486,N_10878,N_13178);
or U17487 (N_17487,N_10276,N_13504);
nor U17488 (N_17488,N_10554,N_11017);
xnor U17489 (N_17489,N_14431,N_13496);
xor U17490 (N_17490,N_11576,N_14489);
and U17491 (N_17491,N_14610,N_10100);
nand U17492 (N_17492,N_13904,N_14026);
nor U17493 (N_17493,N_13047,N_11442);
nand U17494 (N_17494,N_14675,N_12022);
and U17495 (N_17495,N_13990,N_11538);
xnor U17496 (N_17496,N_11715,N_11254);
nor U17497 (N_17497,N_12640,N_10678);
nand U17498 (N_17498,N_10778,N_10398);
nand U17499 (N_17499,N_13602,N_10224);
nand U17500 (N_17500,N_10887,N_14843);
and U17501 (N_17501,N_14330,N_11538);
or U17502 (N_17502,N_11534,N_14593);
and U17503 (N_17503,N_10160,N_11573);
and U17504 (N_17504,N_13788,N_13468);
and U17505 (N_17505,N_13861,N_10835);
xor U17506 (N_17506,N_13855,N_13556);
xnor U17507 (N_17507,N_10149,N_11272);
xor U17508 (N_17508,N_14914,N_11613);
and U17509 (N_17509,N_11637,N_10424);
or U17510 (N_17510,N_12080,N_12758);
or U17511 (N_17511,N_11024,N_14408);
nor U17512 (N_17512,N_12118,N_10869);
nor U17513 (N_17513,N_12004,N_12039);
or U17514 (N_17514,N_11537,N_13145);
or U17515 (N_17515,N_10362,N_12567);
nor U17516 (N_17516,N_13281,N_12427);
and U17517 (N_17517,N_14295,N_12572);
or U17518 (N_17518,N_12266,N_11234);
and U17519 (N_17519,N_13430,N_11233);
or U17520 (N_17520,N_12255,N_11307);
nor U17521 (N_17521,N_10336,N_10421);
or U17522 (N_17522,N_10926,N_13856);
or U17523 (N_17523,N_14980,N_10800);
xnor U17524 (N_17524,N_13762,N_14062);
or U17525 (N_17525,N_12845,N_11821);
xnor U17526 (N_17526,N_13511,N_11469);
or U17527 (N_17527,N_11922,N_10800);
and U17528 (N_17528,N_13197,N_14275);
nor U17529 (N_17529,N_13895,N_12445);
nand U17530 (N_17530,N_11607,N_10608);
nor U17531 (N_17531,N_10139,N_13051);
xnor U17532 (N_17532,N_11218,N_11396);
nor U17533 (N_17533,N_11013,N_13548);
or U17534 (N_17534,N_14739,N_11567);
nand U17535 (N_17535,N_11049,N_13627);
or U17536 (N_17536,N_14030,N_10727);
xnor U17537 (N_17537,N_10889,N_14491);
xor U17538 (N_17538,N_13474,N_10599);
or U17539 (N_17539,N_10214,N_14103);
xnor U17540 (N_17540,N_12549,N_10022);
xor U17541 (N_17541,N_11639,N_13441);
and U17542 (N_17542,N_14462,N_12070);
or U17543 (N_17543,N_14595,N_12336);
or U17544 (N_17544,N_11096,N_10667);
nand U17545 (N_17545,N_12841,N_11537);
or U17546 (N_17546,N_14261,N_11636);
xnor U17547 (N_17547,N_11044,N_10172);
nand U17548 (N_17548,N_14729,N_10113);
xor U17549 (N_17549,N_14229,N_11060);
nand U17550 (N_17550,N_12066,N_13514);
or U17551 (N_17551,N_11976,N_13691);
xnor U17552 (N_17552,N_12896,N_13931);
and U17553 (N_17553,N_10785,N_14858);
xnor U17554 (N_17554,N_12158,N_13192);
or U17555 (N_17555,N_13602,N_10016);
nand U17556 (N_17556,N_10007,N_11889);
nor U17557 (N_17557,N_11768,N_11123);
xor U17558 (N_17558,N_12196,N_10793);
or U17559 (N_17559,N_13991,N_11391);
or U17560 (N_17560,N_13355,N_12447);
or U17561 (N_17561,N_10714,N_14836);
nand U17562 (N_17562,N_13808,N_13613);
xnor U17563 (N_17563,N_10523,N_13188);
and U17564 (N_17564,N_12847,N_11626);
nor U17565 (N_17565,N_14391,N_10746);
or U17566 (N_17566,N_13395,N_14593);
nor U17567 (N_17567,N_10608,N_14808);
xor U17568 (N_17568,N_11253,N_12783);
xor U17569 (N_17569,N_10406,N_14193);
nor U17570 (N_17570,N_13822,N_10858);
nand U17571 (N_17571,N_14433,N_10251);
and U17572 (N_17572,N_14693,N_14355);
nand U17573 (N_17573,N_14045,N_13316);
or U17574 (N_17574,N_13507,N_11815);
and U17575 (N_17575,N_10721,N_10049);
and U17576 (N_17576,N_10982,N_14243);
or U17577 (N_17577,N_10463,N_12892);
and U17578 (N_17578,N_12086,N_14483);
or U17579 (N_17579,N_10870,N_12282);
or U17580 (N_17580,N_12399,N_14872);
nand U17581 (N_17581,N_13482,N_14803);
or U17582 (N_17582,N_14585,N_13693);
nor U17583 (N_17583,N_12053,N_13010);
or U17584 (N_17584,N_11443,N_11059);
and U17585 (N_17585,N_10972,N_11917);
or U17586 (N_17586,N_11951,N_10205);
nor U17587 (N_17587,N_11333,N_11161);
nor U17588 (N_17588,N_10336,N_12913);
xor U17589 (N_17589,N_11173,N_10347);
xnor U17590 (N_17590,N_12938,N_13902);
or U17591 (N_17591,N_10125,N_13259);
nor U17592 (N_17592,N_12286,N_11100);
xor U17593 (N_17593,N_14536,N_14026);
nor U17594 (N_17594,N_14672,N_14243);
xor U17595 (N_17595,N_13412,N_12911);
nor U17596 (N_17596,N_12257,N_11463);
or U17597 (N_17597,N_13384,N_11501);
nor U17598 (N_17598,N_10991,N_13246);
nand U17599 (N_17599,N_11569,N_11114);
xnor U17600 (N_17600,N_13464,N_13458);
and U17601 (N_17601,N_13313,N_12764);
nand U17602 (N_17602,N_11249,N_11379);
or U17603 (N_17603,N_12701,N_14769);
xor U17604 (N_17604,N_11620,N_14246);
nand U17605 (N_17605,N_13327,N_10324);
xor U17606 (N_17606,N_13981,N_12675);
nand U17607 (N_17607,N_12500,N_10055);
xnor U17608 (N_17608,N_14721,N_13475);
xor U17609 (N_17609,N_12526,N_13849);
xor U17610 (N_17610,N_12649,N_11976);
xor U17611 (N_17611,N_11184,N_10717);
and U17612 (N_17612,N_13421,N_11357);
xnor U17613 (N_17613,N_14720,N_12316);
nor U17614 (N_17614,N_11014,N_10485);
or U17615 (N_17615,N_13258,N_10156);
xnor U17616 (N_17616,N_11811,N_12992);
or U17617 (N_17617,N_10900,N_13503);
xor U17618 (N_17618,N_10476,N_13900);
nor U17619 (N_17619,N_11084,N_12627);
nor U17620 (N_17620,N_11781,N_12833);
nand U17621 (N_17621,N_12252,N_14747);
nand U17622 (N_17622,N_12315,N_10047);
nor U17623 (N_17623,N_13985,N_13804);
and U17624 (N_17624,N_11543,N_14879);
nand U17625 (N_17625,N_10340,N_12522);
and U17626 (N_17626,N_14318,N_14162);
nor U17627 (N_17627,N_10170,N_11107);
or U17628 (N_17628,N_10883,N_12177);
xnor U17629 (N_17629,N_11139,N_13371);
nand U17630 (N_17630,N_12559,N_14627);
and U17631 (N_17631,N_12915,N_14522);
nand U17632 (N_17632,N_14082,N_12421);
nand U17633 (N_17633,N_12499,N_10967);
nor U17634 (N_17634,N_10873,N_10890);
nand U17635 (N_17635,N_11224,N_11920);
xor U17636 (N_17636,N_14491,N_11623);
xor U17637 (N_17637,N_13824,N_11110);
and U17638 (N_17638,N_13130,N_13887);
or U17639 (N_17639,N_10907,N_14359);
and U17640 (N_17640,N_10612,N_13916);
or U17641 (N_17641,N_10070,N_11210);
nor U17642 (N_17642,N_13236,N_12684);
xor U17643 (N_17643,N_12581,N_11838);
nand U17644 (N_17644,N_10472,N_10779);
nor U17645 (N_17645,N_11369,N_10151);
xor U17646 (N_17646,N_12162,N_13412);
or U17647 (N_17647,N_14444,N_10988);
or U17648 (N_17648,N_14220,N_10773);
xor U17649 (N_17649,N_10144,N_14568);
xnor U17650 (N_17650,N_11289,N_14978);
nor U17651 (N_17651,N_13127,N_14277);
and U17652 (N_17652,N_10779,N_14206);
and U17653 (N_17653,N_13540,N_11174);
nand U17654 (N_17654,N_13260,N_11960);
or U17655 (N_17655,N_14810,N_14259);
nand U17656 (N_17656,N_11402,N_13137);
or U17657 (N_17657,N_11876,N_10211);
nor U17658 (N_17658,N_11794,N_12881);
or U17659 (N_17659,N_14488,N_14260);
nand U17660 (N_17660,N_11209,N_13056);
xnor U17661 (N_17661,N_13167,N_13534);
and U17662 (N_17662,N_12117,N_10432);
xor U17663 (N_17663,N_13103,N_13857);
nor U17664 (N_17664,N_12279,N_11913);
nor U17665 (N_17665,N_13720,N_13830);
or U17666 (N_17666,N_10879,N_10249);
nand U17667 (N_17667,N_12925,N_11169);
nand U17668 (N_17668,N_12768,N_13811);
or U17669 (N_17669,N_14854,N_10029);
or U17670 (N_17670,N_10936,N_14447);
nor U17671 (N_17671,N_11902,N_12364);
xnor U17672 (N_17672,N_12206,N_13074);
and U17673 (N_17673,N_14728,N_14120);
and U17674 (N_17674,N_12939,N_10709);
nor U17675 (N_17675,N_10371,N_10551);
nor U17676 (N_17676,N_12124,N_14654);
or U17677 (N_17677,N_12475,N_11566);
nand U17678 (N_17678,N_12825,N_12076);
and U17679 (N_17679,N_12696,N_14805);
nor U17680 (N_17680,N_10230,N_11535);
nand U17681 (N_17681,N_14862,N_13662);
or U17682 (N_17682,N_11907,N_10328);
nand U17683 (N_17683,N_12405,N_13502);
or U17684 (N_17684,N_14784,N_13285);
or U17685 (N_17685,N_14799,N_10734);
or U17686 (N_17686,N_12189,N_10989);
and U17687 (N_17687,N_13561,N_10592);
nor U17688 (N_17688,N_10256,N_11484);
xnor U17689 (N_17689,N_12142,N_10027);
xor U17690 (N_17690,N_14081,N_12286);
xnor U17691 (N_17691,N_11074,N_13293);
xor U17692 (N_17692,N_13541,N_14705);
and U17693 (N_17693,N_13755,N_10225);
nand U17694 (N_17694,N_12866,N_12876);
nor U17695 (N_17695,N_13729,N_10120);
and U17696 (N_17696,N_13247,N_14571);
nor U17697 (N_17697,N_11089,N_14302);
xor U17698 (N_17698,N_11204,N_14449);
nand U17699 (N_17699,N_13127,N_13086);
or U17700 (N_17700,N_13329,N_13676);
nor U17701 (N_17701,N_13380,N_13892);
or U17702 (N_17702,N_10057,N_10404);
or U17703 (N_17703,N_12360,N_11583);
or U17704 (N_17704,N_13694,N_12927);
xnor U17705 (N_17705,N_10566,N_14500);
xor U17706 (N_17706,N_11908,N_11846);
xor U17707 (N_17707,N_11190,N_10443);
or U17708 (N_17708,N_10953,N_13219);
and U17709 (N_17709,N_13112,N_10641);
xnor U17710 (N_17710,N_13626,N_14996);
nor U17711 (N_17711,N_10453,N_14161);
nand U17712 (N_17712,N_14543,N_14030);
or U17713 (N_17713,N_12705,N_13876);
and U17714 (N_17714,N_14493,N_13090);
nor U17715 (N_17715,N_13939,N_14526);
nor U17716 (N_17716,N_13799,N_10338);
xor U17717 (N_17717,N_13240,N_12624);
and U17718 (N_17718,N_14747,N_13613);
and U17719 (N_17719,N_12888,N_10327);
and U17720 (N_17720,N_11495,N_11670);
or U17721 (N_17721,N_12455,N_12782);
xnor U17722 (N_17722,N_12195,N_12269);
nor U17723 (N_17723,N_10014,N_11676);
nand U17724 (N_17724,N_10885,N_12884);
nand U17725 (N_17725,N_14254,N_14097);
or U17726 (N_17726,N_14036,N_11220);
or U17727 (N_17727,N_12181,N_11328);
and U17728 (N_17728,N_12177,N_10018);
nand U17729 (N_17729,N_14291,N_13172);
and U17730 (N_17730,N_11437,N_11509);
and U17731 (N_17731,N_11757,N_11106);
and U17732 (N_17732,N_13872,N_14775);
nand U17733 (N_17733,N_11267,N_14006);
xor U17734 (N_17734,N_10461,N_13215);
and U17735 (N_17735,N_10204,N_12474);
or U17736 (N_17736,N_14434,N_10731);
nor U17737 (N_17737,N_10942,N_10427);
xor U17738 (N_17738,N_12615,N_11070);
xnor U17739 (N_17739,N_10009,N_14106);
xnor U17740 (N_17740,N_10370,N_13257);
xor U17741 (N_17741,N_10270,N_14078);
or U17742 (N_17742,N_13747,N_10293);
xor U17743 (N_17743,N_12942,N_10099);
and U17744 (N_17744,N_12838,N_10488);
and U17745 (N_17745,N_10559,N_13725);
and U17746 (N_17746,N_14625,N_10694);
and U17747 (N_17747,N_10131,N_13709);
nor U17748 (N_17748,N_12211,N_11590);
or U17749 (N_17749,N_14797,N_12308);
xnor U17750 (N_17750,N_13382,N_12492);
and U17751 (N_17751,N_12479,N_14221);
or U17752 (N_17752,N_12641,N_11829);
nand U17753 (N_17753,N_12183,N_10460);
and U17754 (N_17754,N_14263,N_12840);
nand U17755 (N_17755,N_12922,N_12974);
xnor U17756 (N_17756,N_14115,N_14259);
nand U17757 (N_17757,N_12411,N_10669);
or U17758 (N_17758,N_14892,N_10848);
xnor U17759 (N_17759,N_10650,N_10983);
nand U17760 (N_17760,N_11740,N_13204);
or U17761 (N_17761,N_13568,N_10552);
nand U17762 (N_17762,N_11610,N_11409);
or U17763 (N_17763,N_10214,N_10286);
nand U17764 (N_17764,N_12324,N_10773);
or U17765 (N_17765,N_12856,N_13199);
nor U17766 (N_17766,N_11113,N_12533);
nand U17767 (N_17767,N_14445,N_10594);
nand U17768 (N_17768,N_13824,N_11491);
nand U17769 (N_17769,N_11496,N_10424);
nand U17770 (N_17770,N_12834,N_10042);
nand U17771 (N_17771,N_14455,N_12536);
nor U17772 (N_17772,N_10816,N_10371);
xor U17773 (N_17773,N_13268,N_13160);
and U17774 (N_17774,N_13348,N_10168);
nor U17775 (N_17775,N_10742,N_13060);
xor U17776 (N_17776,N_11482,N_10976);
xor U17777 (N_17777,N_14996,N_10784);
and U17778 (N_17778,N_14309,N_11252);
and U17779 (N_17779,N_11644,N_10991);
xor U17780 (N_17780,N_10687,N_12717);
nor U17781 (N_17781,N_11872,N_11253);
and U17782 (N_17782,N_13360,N_13364);
or U17783 (N_17783,N_11559,N_13155);
xor U17784 (N_17784,N_14539,N_13812);
and U17785 (N_17785,N_11057,N_12978);
or U17786 (N_17786,N_10286,N_13216);
nand U17787 (N_17787,N_11007,N_12873);
xor U17788 (N_17788,N_13192,N_14529);
or U17789 (N_17789,N_10405,N_13769);
and U17790 (N_17790,N_11162,N_12050);
nand U17791 (N_17791,N_11036,N_14806);
xnor U17792 (N_17792,N_13435,N_12315);
and U17793 (N_17793,N_14926,N_14226);
xnor U17794 (N_17794,N_14392,N_12196);
nor U17795 (N_17795,N_10259,N_14900);
or U17796 (N_17796,N_12785,N_13274);
xnor U17797 (N_17797,N_14764,N_10088);
xor U17798 (N_17798,N_13672,N_10831);
nand U17799 (N_17799,N_12225,N_13720);
nand U17800 (N_17800,N_13919,N_11402);
xor U17801 (N_17801,N_10246,N_12639);
or U17802 (N_17802,N_11910,N_10832);
and U17803 (N_17803,N_13815,N_12415);
nor U17804 (N_17804,N_12195,N_14527);
nand U17805 (N_17805,N_12517,N_11007);
and U17806 (N_17806,N_14321,N_10329);
nor U17807 (N_17807,N_13976,N_14841);
nand U17808 (N_17808,N_10654,N_14623);
nor U17809 (N_17809,N_12361,N_13868);
and U17810 (N_17810,N_10726,N_10354);
nand U17811 (N_17811,N_10546,N_10450);
and U17812 (N_17812,N_10678,N_14926);
or U17813 (N_17813,N_14600,N_11762);
xor U17814 (N_17814,N_10407,N_14950);
nand U17815 (N_17815,N_12926,N_14095);
xor U17816 (N_17816,N_10834,N_13847);
xor U17817 (N_17817,N_14492,N_11339);
and U17818 (N_17818,N_12706,N_14249);
nand U17819 (N_17819,N_13548,N_14839);
and U17820 (N_17820,N_10101,N_14032);
and U17821 (N_17821,N_13726,N_14025);
nand U17822 (N_17822,N_12998,N_12751);
xor U17823 (N_17823,N_10332,N_12206);
nor U17824 (N_17824,N_11319,N_10578);
nor U17825 (N_17825,N_13362,N_12031);
nand U17826 (N_17826,N_13069,N_13065);
or U17827 (N_17827,N_12422,N_12879);
xor U17828 (N_17828,N_12814,N_14875);
or U17829 (N_17829,N_11454,N_12318);
nand U17830 (N_17830,N_14443,N_10050);
nor U17831 (N_17831,N_10842,N_11079);
nand U17832 (N_17832,N_13039,N_10079);
nand U17833 (N_17833,N_14937,N_14730);
nor U17834 (N_17834,N_13692,N_10513);
and U17835 (N_17835,N_14908,N_10637);
or U17836 (N_17836,N_13424,N_10117);
nor U17837 (N_17837,N_14515,N_12900);
and U17838 (N_17838,N_10580,N_14421);
nor U17839 (N_17839,N_12218,N_12393);
xor U17840 (N_17840,N_13897,N_14150);
xor U17841 (N_17841,N_10161,N_13457);
xnor U17842 (N_17842,N_11374,N_14894);
nand U17843 (N_17843,N_11448,N_11867);
nand U17844 (N_17844,N_12481,N_11869);
nand U17845 (N_17845,N_13201,N_12572);
xnor U17846 (N_17846,N_13223,N_14449);
nand U17847 (N_17847,N_12536,N_11682);
nor U17848 (N_17848,N_12981,N_10613);
or U17849 (N_17849,N_10147,N_14944);
xor U17850 (N_17850,N_13628,N_14516);
nor U17851 (N_17851,N_14773,N_13741);
and U17852 (N_17852,N_11080,N_11502);
nor U17853 (N_17853,N_13511,N_12997);
and U17854 (N_17854,N_14457,N_14821);
and U17855 (N_17855,N_14686,N_11053);
nand U17856 (N_17856,N_13983,N_14220);
nor U17857 (N_17857,N_12375,N_13769);
and U17858 (N_17858,N_10050,N_12404);
and U17859 (N_17859,N_13584,N_10247);
nand U17860 (N_17860,N_10756,N_10744);
or U17861 (N_17861,N_12316,N_14738);
nor U17862 (N_17862,N_13572,N_14314);
and U17863 (N_17863,N_14678,N_13689);
and U17864 (N_17864,N_13471,N_12627);
and U17865 (N_17865,N_12959,N_13610);
xnor U17866 (N_17866,N_10713,N_11637);
or U17867 (N_17867,N_11235,N_14305);
nor U17868 (N_17868,N_12290,N_10599);
nand U17869 (N_17869,N_11345,N_10226);
or U17870 (N_17870,N_13444,N_11503);
xor U17871 (N_17871,N_13053,N_11092);
or U17872 (N_17872,N_12390,N_14476);
nor U17873 (N_17873,N_11675,N_10931);
nor U17874 (N_17874,N_10752,N_13694);
xor U17875 (N_17875,N_12985,N_14683);
or U17876 (N_17876,N_10269,N_12846);
and U17877 (N_17877,N_14340,N_14956);
or U17878 (N_17878,N_14879,N_14766);
nor U17879 (N_17879,N_14735,N_11434);
xor U17880 (N_17880,N_11078,N_11596);
nor U17881 (N_17881,N_13818,N_12662);
and U17882 (N_17882,N_11747,N_13551);
nor U17883 (N_17883,N_12260,N_12704);
nand U17884 (N_17884,N_11458,N_14844);
or U17885 (N_17885,N_10928,N_10127);
xnor U17886 (N_17886,N_11648,N_12379);
or U17887 (N_17887,N_11768,N_13687);
or U17888 (N_17888,N_13505,N_10226);
nand U17889 (N_17889,N_14099,N_14731);
or U17890 (N_17890,N_11923,N_10630);
nor U17891 (N_17891,N_12133,N_10742);
and U17892 (N_17892,N_14887,N_12406);
nor U17893 (N_17893,N_13355,N_13108);
xnor U17894 (N_17894,N_14126,N_12529);
and U17895 (N_17895,N_12665,N_12704);
nor U17896 (N_17896,N_10477,N_14438);
nor U17897 (N_17897,N_14111,N_13450);
nor U17898 (N_17898,N_10974,N_13927);
or U17899 (N_17899,N_12137,N_13732);
xnor U17900 (N_17900,N_13321,N_14879);
nand U17901 (N_17901,N_10287,N_10463);
nor U17902 (N_17902,N_13947,N_14877);
and U17903 (N_17903,N_14308,N_14153);
or U17904 (N_17904,N_11807,N_14687);
and U17905 (N_17905,N_14648,N_10160);
or U17906 (N_17906,N_13846,N_10465);
nand U17907 (N_17907,N_12392,N_11927);
and U17908 (N_17908,N_13129,N_12140);
nand U17909 (N_17909,N_10918,N_11283);
nor U17910 (N_17910,N_11051,N_11691);
or U17911 (N_17911,N_12607,N_11946);
and U17912 (N_17912,N_12836,N_14016);
and U17913 (N_17913,N_12555,N_13865);
and U17914 (N_17914,N_14925,N_14309);
xnor U17915 (N_17915,N_12250,N_10102);
nor U17916 (N_17916,N_11265,N_11239);
nand U17917 (N_17917,N_12191,N_13252);
or U17918 (N_17918,N_10439,N_11102);
or U17919 (N_17919,N_14280,N_13786);
nand U17920 (N_17920,N_10244,N_14686);
xor U17921 (N_17921,N_13339,N_12580);
nand U17922 (N_17922,N_10901,N_12438);
and U17923 (N_17923,N_10160,N_11793);
or U17924 (N_17924,N_13182,N_14097);
nand U17925 (N_17925,N_14823,N_11859);
xor U17926 (N_17926,N_12868,N_14126);
nand U17927 (N_17927,N_13094,N_11768);
or U17928 (N_17928,N_11191,N_11158);
or U17929 (N_17929,N_12585,N_10450);
xnor U17930 (N_17930,N_13381,N_13020);
nor U17931 (N_17931,N_14034,N_10973);
nand U17932 (N_17932,N_13474,N_13127);
xor U17933 (N_17933,N_14806,N_11749);
xnor U17934 (N_17934,N_12524,N_14959);
nand U17935 (N_17935,N_13804,N_14956);
nor U17936 (N_17936,N_10755,N_13947);
xnor U17937 (N_17937,N_12104,N_13768);
and U17938 (N_17938,N_13880,N_13539);
xor U17939 (N_17939,N_13591,N_13537);
xnor U17940 (N_17940,N_10952,N_13488);
nand U17941 (N_17941,N_11143,N_11900);
or U17942 (N_17942,N_11895,N_11262);
xnor U17943 (N_17943,N_14933,N_10551);
or U17944 (N_17944,N_14288,N_11582);
nand U17945 (N_17945,N_13256,N_11428);
nor U17946 (N_17946,N_12370,N_13855);
or U17947 (N_17947,N_11624,N_13008);
nor U17948 (N_17948,N_14663,N_14888);
and U17949 (N_17949,N_14970,N_10200);
nor U17950 (N_17950,N_13698,N_10383);
and U17951 (N_17951,N_12664,N_10437);
xor U17952 (N_17952,N_13286,N_10574);
xnor U17953 (N_17953,N_11352,N_12400);
nor U17954 (N_17954,N_14854,N_12604);
nand U17955 (N_17955,N_11933,N_11529);
nand U17956 (N_17956,N_12230,N_11668);
xnor U17957 (N_17957,N_12828,N_13221);
xor U17958 (N_17958,N_13624,N_13818);
and U17959 (N_17959,N_13652,N_14369);
nand U17960 (N_17960,N_12560,N_14497);
nand U17961 (N_17961,N_13387,N_14681);
and U17962 (N_17962,N_10740,N_11375);
nand U17963 (N_17963,N_10193,N_13366);
nor U17964 (N_17964,N_11639,N_10804);
nand U17965 (N_17965,N_12512,N_13750);
nand U17966 (N_17966,N_13581,N_11616);
xnor U17967 (N_17967,N_12014,N_13532);
or U17968 (N_17968,N_12082,N_14647);
or U17969 (N_17969,N_14484,N_14074);
xor U17970 (N_17970,N_10265,N_10778);
nor U17971 (N_17971,N_12053,N_14529);
nand U17972 (N_17972,N_11202,N_14181);
nand U17973 (N_17973,N_10736,N_13831);
and U17974 (N_17974,N_12861,N_12943);
and U17975 (N_17975,N_10905,N_10200);
xor U17976 (N_17976,N_12879,N_14227);
xor U17977 (N_17977,N_10813,N_10189);
nor U17978 (N_17978,N_14318,N_11944);
xor U17979 (N_17979,N_10810,N_14468);
nand U17980 (N_17980,N_13486,N_11835);
nor U17981 (N_17981,N_14307,N_10269);
nor U17982 (N_17982,N_12821,N_14755);
xor U17983 (N_17983,N_12449,N_13949);
and U17984 (N_17984,N_13504,N_11283);
nor U17985 (N_17985,N_11718,N_12235);
nor U17986 (N_17986,N_13908,N_11665);
or U17987 (N_17987,N_14124,N_11123);
xor U17988 (N_17988,N_12566,N_10458);
or U17989 (N_17989,N_12377,N_12744);
or U17990 (N_17990,N_13288,N_13024);
or U17991 (N_17991,N_12547,N_10974);
or U17992 (N_17992,N_13743,N_14943);
nand U17993 (N_17993,N_13529,N_14480);
nor U17994 (N_17994,N_11735,N_10641);
or U17995 (N_17995,N_11052,N_11015);
nor U17996 (N_17996,N_12780,N_14433);
xnor U17997 (N_17997,N_13468,N_14451);
nor U17998 (N_17998,N_14539,N_10172);
or U17999 (N_17999,N_11053,N_13402);
nor U18000 (N_18000,N_11871,N_12965);
and U18001 (N_18001,N_13602,N_10816);
nand U18002 (N_18002,N_13044,N_10525);
xor U18003 (N_18003,N_10031,N_14591);
nand U18004 (N_18004,N_12749,N_10410);
nor U18005 (N_18005,N_12414,N_12111);
xor U18006 (N_18006,N_12353,N_13814);
or U18007 (N_18007,N_10992,N_10835);
nor U18008 (N_18008,N_10997,N_13020);
or U18009 (N_18009,N_12067,N_12478);
and U18010 (N_18010,N_13088,N_14575);
or U18011 (N_18011,N_11126,N_14978);
xor U18012 (N_18012,N_13842,N_11794);
xnor U18013 (N_18013,N_14443,N_10988);
nand U18014 (N_18014,N_13710,N_13929);
nand U18015 (N_18015,N_10041,N_10901);
nor U18016 (N_18016,N_14177,N_13310);
or U18017 (N_18017,N_14045,N_11874);
xnor U18018 (N_18018,N_10364,N_12595);
nor U18019 (N_18019,N_12298,N_12661);
nor U18020 (N_18020,N_10369,N_11301);
or U18021 (N_18021,N_13498,N_12465);
xor U18022 (N_18022,N_11482,N_11313);
and U18023 (N_18023,N_13664,N_14490);
or U18024 (N_18024,N_14551,N_13783);
or U18025 (N_18025,N_14244,N_13486);
and U18026 (N_18026,N_11271,N_11468);
nand U18027 (N_18027,N_11884,N_14680);
nor U18028 (N_18028,N_11593,N_11142);
nor U18029 (N_18029,N_13499,N_12238);
nor U18030 (N_18030,N_10324,N_13791);
nand U18031 (N_18031,N_11844,N_13792);
nor U18032 (N_18032,N_13777,N_12903);
nand U18033 (N_18033,N_11113,N_13548);
nand U18034 (N_18034,N_12516,N_12861);
and U18035 (N_18035,N_13160,N_13663);
nor U18036 (N_18036,N_11845,N_14918);
nor U18037 (N_18037,N_12045,N_12920);
nor U18038 (N_18038,N_10752,N_11432);
nor U18039 (N_18039,N_11018,N_13603);
nand U18040 (N_18040,N_14896,N_12059);
or U18041 (N_18041,N_13004,N_10706);
or U18042 (N_18042,N_10081,N_10390);
nand U18043 (N_18043,N_11981,N_14639);
nor U18044 (N_18044,N_10771,N_11128);
xnor U18045 (N_18045,N_13938,N_11741);
nor U18046 (N_18046,N_14423,N_10195);
nor U18047 (N_18047,N_10331,N_12902);
nand U18048 (N_18048,N_10127,N_10641);
and U18049 (N_18049,N_10089,N_12578);
or U18050 (N_18050,N_11039,N_13456);
nor U18051 (N_18051,N_14236,N_12903);
xor U18052 (N_18052,N_10698,N_10893);
nor U18053 (N_18053,N_13567,N_11831);
and U18054 (N_18054,N_10875,N_13556);
and U18055 (N_18055,N_14188,N_10956);
or U18056 (N_18056,N_13269,N_14877);
and U18057 (N_18057,N_12014,N_10951);
xor U18058 (N_18058,N_12695,N_13367);
and U18059 (N_18059,N_10997,N_12682);
xnor U18060 (N_18060,N_12723,N_12747);
xor U18061 (N_18061,N_14776,N_12334);
xor U18062 (N_18062,N_10168,N_13559);
xnor U18063 (N_18063,N_13601,N_14389);
or U18064 (N_18064,N_11554,N_11985);
and U18065 (N_18065,N_14528,N_11569);
nor U18066 (N_18066,N_11306,N_12247);
and U18067 (N_18067,N_14868,N_11294);
nor U18068 (N_18068,N_13309,N_10506);
and U18069 (N_18069,N_12251,N_11006);
and U18070 (N_18070,N_12123,N_10757);
nand U18071 (N_18071,N_10845,N_12291);
nand U18072 (N_18072,N_12579,N_13598);
and U18073 (N_18073,N_11878,N_13100);
and U18074 (N_18074,N_13892,N_11694);
nand U18075 (N_18075,N_10761,N_10850);
nor U18076 (N_18076,N_10051,N_14685);
nand U18077 (N_18077,N_10374,N_11459);
and U18078 (N_18078,N_13365,N_11816);
or U18079 (N_18079,N_13368,N_11750);
and U18080 (N_18080,N_14211,N_13634);
xnor U18081 (N_18081,N_11926,N_13341);
nor U18082 (N_18082,N_10163,N_11825);
nand U18083 (N_18083,N_13250,N_12011);
nor U18084 (N_18084,N_13102,N_11653);
and U18085 (N_18085,N_11623,N_13653);
nand U18086 (N_18086,N_11698,N_11259);
or U18087 (N_18087,N_13917,N_11588);
or U18088 (N_18088,N_11587,N_14823);
or U18089 (N_18089,N_14845,N_13993);
and U18090 (N_18090,N_11392,N_12763);
xor U18091 (N_18091,N_12441,N_10610);
xnor U18092 (N_18092,N_14543,N_11316);
nor U18093 (N_18093,N_12440,N_14190);
nand U18094 (N_18094,N_14411,N_13207);
nand U18095 (N_18095,N_11822,N_12940);
nor U18096 (N_18096,N_12841,N_11401);
and U18097 (N_18097,N_12899,N_14655);
nor U18098 (N_18098,N_12743,N_11866);
xor U18099 (N_18099,N_12887,N_14819);
or U18100 (N_18100,N_14014,N_12393);
nor U18101 (N_18101,N_11872,N_11194);
nand U18102 (N_18102,N_13717,N_10475);
nor U18103 (N_18103,N_13804,N_14962);
xnor U18104 (N_18104,N_12078,N_11109);
xnor U18105 (N_18105,N_10261,N_11607);
or U18106 (N_18106,N_10618,N_11413);
and U18107 (N_18107,N_11266,N_13525);
nor U18108 (N_18108,N_14992,N_14328);
nor U18109 (N_18109,N_14388,N_13921);
nor U18110 (N_18110,N_10522,N_13360);
xnor U18111 (N_18111,N_13039,N_11282);
xnor U18112 (N_18112,N_11055,N_11297);
or U18113 (N_18113,N_11141,N_11298);
and U18114 (N_18114,N_11088,N_10852);
or U18115 (N_18115,N_11461,N_11694);
nor U18116 (N_18116,N_12818,N_11213);
nor U18117 (N_18117,N_13057,N_14071);
and U18118 (N_18118,N_11948,N_13867);
nand U18119 (N_18119,N_11884,N_11896);
or U18120 (N_18120,N_12817,N_11682);
or U18121 (N_18121,N_10534,N_13819);
nor U18122 (N_18122,N_13198,N_12290);
and U18123 (N_18123,N_12541,N_13818);
nor U18124 (N_18124,N_13937,N_14678);
and U18125 (N_18125,N_14747,N_14915);
nor U18126 (N_18126,N_12864,N_11985);
nand U18127 (N_18127,N_10362,N_13866);
and U18128 (N_18128,N_10099,N_11892);
nor U18129 (N_18129,N_10503,N_10346);
nand U18130 (N_18130,N_13491,N_10130);
nand U18131 (N_18131,N_13470,N_12556);
nand U18132 (N_18132,N_13835,N_11589);
nand U18133 (N_18133,N_11572,N_13267);
nand U18134 (N_18134,N_10286,N_14099);
and U18135 (N_18135,N_11153,N_10852);
nor U18136 (N_18136,N_11917,N_13213);
nor U18137 (N_18137,N_14321,N_13611);
xor U18138 (N_18138,N_10097,N_12897);
nand U18139 (N_18139,N_12985,N_13535);
nand U18140 (N_18140,N_14335,N_11698);
and U18141 (N_18141,N_14208,N_13023);
nand U18142 (N_18142,N_11828,N_10428);
or U18143 (N_18143,N_14042,N_14215);
nand U18144 (N_18144,N_10961,N_13951);
and U18145 (N_18145,N_11860,N_13255);
or U18146 (N_18146,N_11619,N_12064);
nand U18147 (N_18147,N_13868,N_14417);
or U18148 (N_18148,N_12546,N_13123);
xnor U18149 (N_18149,N_12458,N_13288);
nor U18150 (N_18150,N_10622,N_13156);
nand U18151 (N_18151,N_13442,N_11756);
or U18152 (N_18152,N_12283,N_14006);
and U18153 (N_18153,N_13415,N_10947);
nor U18154 (N_18154,N_13953,N_13927);
nor U18155 (N_18155,N_10320,N_13116);
nor U18156 (N_18156,N_10928,N_13329);
and U18157 (N_18157,N_10801,N_11669);
nand U18158 (N_18158,N_12321,N_13420);
or U18159 (N_18159,N_13962,N_12617);
or U18160 (N_18160,N_14580,N_12080);
and U18161 (N_18161,N_12722,N_11855);
xnor U18162 (N_18162,N_10996,N_10204);
nor U18163 (N_18163,N_12296,N_13619);
xnor U18164 (N_18164,N_13177,N_12982);
nand U18165 (N_18165,N_13309,N_12456);
or U18166 (N_18166,N_13261,N_10289);
xnor U18167 (N_18167,N_11562,N_13085);
xor U18168 (N_18168,N_11910,N_11592);
or U18169 (N_18169,N_14376,N_11006);
nor U18170 (N_18170,N_12309,N_10725);
and U18171 (N_18171,N_10956,N_13937);
and U18172 (N_18172,N_11672,N_10376);
nor U18173 (N_18173,N_13604,N_13350);
nand U18174 (N_18174,N_12010,N_11455);
or U18175 (N_18175,N_12936,N_13248);
nor U18176 (N_18176,N_13904,N_13131);
xor U18177 (N_18177,N_13772,N_11076);
nor U18178 (N_18178,N_12050,N_11349);
nand U18179 (N_18179,N_13216,N_14087);
nand U18180 (N_18180,N_11866,N_11962);
xnor U18181 (N_18181,N_13530,N_10839);
xnor U18182 (N_18182,N_12103,N_13167);
nand U18183 (N_18183,N_10803,N_12398);
or U18184 (N_18184,N_11818,N_13974);
xor U18185 (N_18185,N_13342,N_13614);
or U18186 (N_18186,N_12254,N_10226);
nand U18187 (N_18187,N_14008,N_12765);
or U18188 (N_18188,N_14086,N_12048);
nor U18189 (N_18189,N_14311,N_11687);
or U18190 (N_18190,N_14952,N_11054);
and U18191 (N_18191,N_10529,N_11067);
nand U18192 (N_18192,N_11284,N_14061);
nand U18193 (N_18193,N_11827,N_13221);
xnor U18194 (N_18194,N_13517,N_12947);
or U18195 (N_18195,N_10428,N_14157);
nand U18196 (N_18196,N_14360,N_14326);
xor U18197 (N_18197,N_10194,N_10120);
xor U18198 (N_18198,N_13148,N_13192);
or U18199 (N_18199,N_13997,N_14233);
or U18200 (N_18200,N_12846,N_12294);
xnor U18201 (N_18201,N_10880,N_14873);
xor U18202 (N_18202,N_11565,N_10133);
or U18203 (N_18203,N_12310,N_14745);
xnor U18204 (N_18204,N_12792,N_13418);
nand U18205 (N_18205,N_14482,N_14889);
xor U18206 (N_18206,N_13491,N_11561);
nand U18207 (N_18207,N_10691,N_12480);
nand U18208 (N_18208,N_14832,N_14357);
and U18209 (N_18209,N_12311,N_12298);
nor U18210 (N_18210,N_12960,N_14904);
and U18211 (N_18211,N_14002,N_10867);
nor U18212 (N_18212,N_14508,N_12899);
nand U18213 (N_18213,N_13415,N_10003);
nor U18214 (N_18214,N_11451,N_14856);
nor U18215 (N_18215,N_12107,N_12883);
xor U18216 (N_18216,N_11278,N_12635);
nor U18217 (N_18217,N_12080,N_10394);
and U18218 (N_18218,N_11642,N_10301);
nor U18219 (N_18219,N_13958,N_13314);
nand U18220 (N_18220,N_11950,N_13582);
xor U18221 (N_18221,N_11581,N_13959);
or U18222 (N_18222,N_13733,N_10335);
nor U18223 (N_18223,N_12067,N_11276);
xor U18224 (N_18224,N_11515,N_11662);
nor U18225 (N_18225,N_12862,N_12638);
nand U18226 (N_18226,N_12554,N_13864);
nor U18227 (N_18227,N_14290,N_12256);
or U18228 (N_18228,N_13240,N_13348);
nand U18229 (N_18229,N_14878,N_13568);
and U18230 (N_18230,N_13535,N_10388);
xor U18231 (N_18231,N_10021,N_11597);
xor U18232 (N_18232,N_10191,N_13749);
nor U18233 (N_18233,N_13831,N_14168);
or U18234 (N_18234,N_12807,N_11472);
nand U18235 (N_18235,N_13804,N_12581);
or U18236 (N_18236,N_13225,N_10640);
nor U18237 (N_18237,N_14711,N_14662);
xor U18238 (N_18238,N_10959,N_10443);
xor U18239 (N_18239,N_13180,N_11499);
nand U18240 (N_18240,N_10055,N_10121);
xnor U18241 (N_18241,N_14287,N_14650);
nor U18242 (N_18242,N_11087,N_11366);
nor U18243 (N_18243,N_11168,N_10188);
or U18244 (N_18244,N_12129,N_11480);
and U18245 (N_18245,N_14257,N_12598);
and U18246 (N_18246,N_14631,N_13019);
nand U18247 (N_18247,N_13265,N_14458);
xor U18248 (N_18248,N_14892,N_10609);
xor U18249 (N_18249,N_14534,N_12979);
xor U18250 (N_18250,N_13995,N_11484);
xnor U18251 (N_18251,N_14572,N_13240);
and U18252 (N_18252,N_11439,N_11302);
nor U18253 (N_18253,N_10322,N_13645);
xnor U18254 (N_18254,N_12785,N_10383);
and U18255 (N_18255,N_13062,N_12927);
and U18256 (N_18256,N_10081,N_13093);
and U18257 (N_18257,N_12020,N_12290);
xnor U18258 (N_18258,N_11561,N_12630);
xor U18259 (N_18259,N_14406,N_10923);
nor U18260 (N_18260,N_13906,N_13122);
nor U18261 (N_18261,N_13777,N_14263);
nor U18262 (N_18262,N_14306,N_12802);
nand U18263 (N_18263,N_12317,N_13116);
nand U18264 (N_18264,N_13723,N_13344);
nand U18265 (N_18265,N_10968,N_11093);
and U18266 (N_18266,N_11122,N_10905);
or U18267 (N_18267,N_10725,N_10536);
xnor U18268 (N_18268,N_10759,N_14812);
nand U18269 (N_18269,N_10908,N_11427);
xnor U18270 (N_18270,N_11716,N_11524);
and U18271 (N_18271,N_14520,N_11260);
nand U18272 (N_18272,N_11948,N_12970);
or U18273 (N_18273,N_12354,N_10039);
or U18274 (N_18274,N_14346,N_14298);
and U18275 (N_18275,N_11845,N_11040);
nor U18276 (N_18276,N_12740,N_12794);
nor U18277 (N_18277,N_10449,N_10839);
or U18278 (N_18278,N_11499,N_11957);
nor U18279 (N_18279,N_13742,N_13511);
nor U18280 (N_18280,N_13742,N_10859);
and U18281 (N_18281,N_10012,N_14079);
and U18282 (N_18282,N_11734,N_14365);
and U18283 (N_18283,N_11327,N_14955);
or U18284 (N_18284,N_12511,N_14909);
nand U18285 (N_18285,N_11215,N_14873);
nand U18286 (N_18286,N_11562,N_14426);
and U18287 (N_18287,N_14774,N_11778);
and U18288 (N_18288,N_12260,N_12541);
or U18289 (N_18289,N_11083,N_11728);
xnor U18290 (N_18290,N_14512,N_12591);
and U18291 (N_18291,N_11754,N_14135);
nor U18292 (N_18292,N_12131,N_14401);
xnor U18293 (N_18293,N_13172,N_13706);
nand U18294 (N_18294,N_14567,N_11826);
nand U18295 (N_18295,N_11865,N_13196);
and U18296 (N_18296,N_14431,N_12521);
and U18297 (N_18297,N_14510,N_11034);
and U18298 (N_18298,N_11053,N_12472);
xnor U18299 (N_18299,N_12445,N_13083);
or U18300 (N_18300,N_13289,N_10566);
xor U18301 (N_18301,N_13429,N_12767);
xor U18302 (N_18302,N_13718,N_10071);
nand U18303 (N_18303,N_13524,N_14858);
or U18304 (N_18304,N_11947,N_13251);
xnor U18305 (N_18305,N_10808,N_12021);
nor U18306 (N_18306,N_11189,N_14139);
xnor U18307 (N_18307,N_13445,N_12932);
nand U18308 (N_18308,N_13820,N_12984);
and U18309 (N_18309,N_12319,N_11166);
or U18310 (N_18310,N_11684,N_12181);
xor U18311 (N_18311,N_10499,N_13071);
nor U18312 (N_18312,N_11780,N_10535);
or U18313 (N_18313,N_11574,N_13472);
xor U18314 (N_18314,N_11347,N_11520);
or U18315 (N_18315,N_12264,N_10966);
or U18316 (N_18316,N_14647,N_10272);
nor U18317 (N_18317,N_13998,N_12395);
and U18318 (N_18318,N_10092,N_14000);
xor U18319 (N_18319,N_12469,N_14784);
and U18320 (N_18320,N_14252,N_13430);
nor U18321 (N_18321,N_12362,N_14296);
nand U18322 (N_18322,N_11526,N_13671);
and U18323 (N_18323,N_14954,N_10226);
or U18324 (N_18324,N_14868,N_10132);
xor U18325 (N_18325,N_12507,N_12915);
nand U18326 (N_18326,N_12247,N_12321);
xnor U18327 (N_18327,N_11830,N_13178);
or U18328 (N_18328,N_12096,N_11349);
or U18329 (N_18329,N_11299,N_12031);
nor U18330 (N_18330,N_11717,N_10747);
xor U18331 (N_18331,N_10344,N_13982);
nor U18332 (N_18332,N_10397,N_13710);
and U18333 (N_18333,N_14988,N_11682);
xnor U18334 (N_18334,N_13053,N_12135);
and U18335 (N_18335,N_14603,N_10522);
and U18336 (N_18336,N_11317,N_11657);
nor U18337 (N_18337,N_14790,N_13631);
and U18338 (N_18338,N_14360,N_14112);
nor U18339 (N_18339,N_13591,N_14129);
and U18340 (N_18340,N_13886,N_10196);
or U18341 (N_18341,N_12464,N_12924);
or U18342 (N_18342,N_14532,N_14239);
or U18343 (N_18343,N_13951,N_12273);
or U18344 (N_18344,N_11315,N_13681);
xnor U18345 (N_18345,N_14253,N_14181);
nor U18346 (N_18346,N_12591,N_14252);
or U18347 (N_18347,N_13072,N_10978);
nand U18348 (N_18348,N_13307,N_13103);
or U18349 (N_18349,N_12989,N_12351);
nor U18350 (N_18350,N_12980,N_14775);
nand U18351 (N_18351,N_11247,N_12763);
nor U18352 (N_18352,N_11435,N_12191);
nand U18353 (N_18353,N_11394,N_10063);
and U18354 (N_18354,N_10906,N_10390);
xnor U18355 (N_18355,N_11932,N_14511);
nand U18356 (N_18356,N_12942,N_13093);
nor U18357 (N_18357,N_13143,N_10108);
xor U18358 (N_18358,N_12731,N_10062);
nor U18359 (N_18359,N_14476,N_11702);
nand U18360 (N_18360,N_13842,N_12176);
nand U18361 (N_18361,N_14335,N_13590);
xor U18362 (N_18362,N_10931,N_13069);
nand U18363 (N_18363,N_13485,N_11860);
xor U18364 (N_18364,N_11776,N_10438);
nand U18365 (N_18365,N_14841,N_12146);
xor U18366 (N_18366,N_10187,N_13420);
xor U18367 (N_18367,N_12179,N_12504);
xor U18368 (N_18368,N_12826,N_10215);
nand U18369 (N_18369,N_12294,N_14306);
nand U18370 (N_18370,N_10926,N_13285);
and U18371 (N_18371,N_12319,N_10974);
nor U18372 (N_18372,N_12466,N_10965);
nor U18373 (N_18373,N_12756,N_11389);
xnor U18374 (N_18374,N_12628,N_12279);
and U18375 (N_18375,N_13448,N_13082);
xnor U18376 (N_18376,N_14307,N_11479);
nand U18377 (N_18377,N_12830,N_11044);
or U18378 (N_18378,N_14524,N_14970);
and U18379 (N_18379,N_12330,N_14360);
nor U18380 (N_18380,N_14615,N_12161);
and U18381 (N_18381,N_12147,N_13854);
xor U18382 (N_18382,N_11799,N_12102);
nor U18383 (N_18383,N_13085,N_13917);
xor U18384 (N_18384,N_10208,N_10742);
nor U18385 (N_18385,N_14117,N_14382);
xnor U18386 (N_18386,N_11009,N_12339);
or U18387 (N_18387,N_14403,N_12948);
or U18388 (N_18388,N_12836,N_10630);
nand U18389 (N_18389,N_11852,N_12195);
xor U18390 (N_18390,N_14123,N_10736);
nand U18391 (N_18391,N_14867,N_11139);
xor U18392 (N_18392,N_13286,N_10161);
or U18393 (N_18393,N_12751,N_11985);
or U18394 (N_18394,N_11172,N_13455);
or U18395 (N_18395,N_12712,N_11219);
nor U18396 (N_18396,N_10622,N_14522);
nand U18397 (N_18397,N_11810,N_11106);
nand U18398 (N_18398,N_11798,N_10838);
nand U18399 (N_18399,N_13387,N_13231);
xnor U18400 (N_18400,N_12807,N_14980);
nor U18401 (N_18401,N_11838,N_14892);
nor U18402 (N_18402,N_11755,N_11021);
or U18403 (N_18403,N_12384,N_10702);
or U18404 (N_18404,N_14656,N_12188);
nand U18405 (N_18405,N_14580,N_10989);
xor U18406 (N_18406,N_12974,N_11966);
nor U18407 (N_18407,N_10715,N_10757);
and U18408 (N_18408,N_10993,N_10984);
nor U18409 (N_18409,N_11484,N_10053);
or U18410 (N_18410,N_12211,N_14201);
xnor U18411 (N_18411,N_14453,N_14224);
and U18412 (N_18412,N_12601,N_12956);
xor U18413 (N_18413,N_10828,N_14752);
or U18414 (N_18414,N_13318,N_11933);
nand U18415 (N_18415,N_13810,N_12893);
xor U18416 (N_18416,N_14856,N_14142);
or U18417 (N_18417,N_13460,N_12112);
nand U18418 (N_18418,N_11192,N_11325);
nand U18419 (N_18419,N_12107,N_12150);
and U18420 (N_18420,N_10104,N_12422);
nor U18421 (N_18421,N_11496,N_12335);
xnor U18422 (N_18422,N_10378,N_12487);
nor U18423 (N_18423,N_12399,N_10160);
nand U18424 (N_18424,N_12086,N_13252);
and U18425 (N_18425,N_13521,N_14601);
and U18426 (N_18426,N_11636,N_12227);
nand U18427 (N_18427,N_12676,N_11079);
nand U18428 (N_18428,N_14041,N_12012);
xor U18429 (N_18429,N_14773,N_10878);
or U18430 (N_18430,N_10349,N_12961);
and U18431 (N_18431,N_10967,N_10896);
xnor U18432 (N_18432,N_11296,N_11661);
nor U18433 (N_18433,N_13524,N_11182);
nor U18434 (N_18434,N_13817,N_13700);
xnor U18435 (N_18435,N_11463,N_10629);
or U18436 (N_18436,N_14430,N_13932);
nand U18437 (N_18437,N_14683,N_11287);
and U18438 (N_18438,N_12405,N_13314);
xnor U18439 (N_18439,N_10265,N_14978);
and U18440 (N_18440,N_13966,N_12035);
xor U18441 (N_18441,N_13037,N_11918);
xnor U18442 (N_18442,N_13098,N_11789);
xor U18443 (N_18443,N_14086,N_12442);
nand U18444 (N_18444,N_14139,N_14191);
xor U18445 (N_18445,N_10000,N_14481);
nand U18446 (N_18446,N_12317,N_12920);
nor U18447 (N_18447,N_12057,N_13308);
and U18448 (N_18448,N_11706,N_12691);
xor U18449 (N_18449,N_11388,N_11034);
and U18450 (N_18450,N_13734,N_14070);
xor U18451 (N_18451,N_13827,N_11998);
nand U18452 (N_18452,N_10259,N_11621);
nor U18453 (N_18453,N_14658,N_10483);
or U18454 (N_18454,N_11193,N_14145);
and U18455 (N_18455,N_12617,N_14998);
xor U18456 (N_18456,N_11065,N_11530);
and U18457 (N_18457,N_10452,N_10547);
and U18458 (N_18458,N_12607,N_13783);
or U18459 (N_18459,N_14593,N_14609);
xor U18460 (N_18460,N_14882,N_13417);
nor U18461 (N_18461,N_11107,N_13075);
nand U18462 (N_18462,N_11704,N_14641);
xnor U18463 (N_18463,N_12788,N_14536);
nor U18464 (N_18464,N_10428,N_13777);
nor U18465 (N_18465,N_13198,N_11110);
nor U18466 (N_18466,N_13637,N_11107);
nor U18467 (N_18467,N_11613,N_10174);
xnor U18468 (N_18468,N_12478,N_13636);
xnor U18469 (N_18469,N_11548,N_10096);
and U18470 (N_18470,N_14916,N_10939);
nand U18471 (N_18471,N_11539,N_13282);
and U18472 (N_18472,N_14095,N_10032);
nand U18473 (N_18473,N_13838,N_11808);
nor U18474 (N_18474,N_14038,N_10360);
xor U18475 (N_18475,N_12487,N_11175);
or U18476 (N_18476,N_14231,N_13249);
nand U18477 (N_18477,N_13719,N_11040);
nor U18478 (N_18478,N_12454,N_11752);
nor U18479 (N_18479,N_14868,N_12952);
nand U18480 (N_18480,N_11683,N_13810);
and U18481 (N_18481,N_14314,N_12603);
or U18482 (N_18482,N_12166,N_12309);
and U18483 (N_18483,N_14061,N_13797);
xor U18484 (N_18484,N_11707,N_10041);
nor U18485 (N_18485,N_11744,N_12327);
nor U18486 (N_18486,N_14317,N_11468);
or U18487 (N_18487,N_11707,N_10458);
or U18488 (N_18488,N_12932,N_11619);
or U18489 (N_18489,N_14173,N_11682);
or U18490 (N_18490,N_14617,N_13887);
nand U18491 (N_18491,N_11792,N_11518);
nor U18492 (N_18492,N_11553,N_11915);
nor U18493 (N_18493,N_13024,N_11524);
nor U18494 (N_18494,N_13164,N_10999);
or U18495 (N_18495,N_10592,N_14343);
or U18496 (N_18496,N_13098,N_11932);
xor U18497 (N_18497,N_12053,N_11877);
nand U18498 (N_18498,N_12211,N_14378);
xor U18499 (N_18499,N_13890,N_13784);
xnor U18500 (N_18500,N_13372,N_11940);
xor U18501 (N_18501,N_12061,N_14950);
nor U18502 (N_18502,N_12781,N_12491);
xor U18503 (N_18503,N_10349,N_12951);
nand U18504 (N_18504,N_13458,N_11862);
xor U18505 (N_18505,N_14097,N_12331);
and U18506 (N_18506,N_14142,N_13394);
nor U18507 (N_18507,N_14001,N_13650);
or U18508 (N_18508,N_12053,N_13348);
and U18509 (N_18509,N_13015,N_13022);
nand U18510 (N_18510,N_14954,N_12375);
nor U18511 (N_18511,N_14675,N_14128);
and U18512 (N_18512,N_11075,N_10196);
xnor U18513 (N_18513,N_12904,N_11982);
and U18514 (N_18514,N_12312,N_12391);
and U18515 (N_18515,N_11926,N_14372);
xnor U18516 (N_18516,N_11986,N_13778);
nor U18517 (N_18517,N_11868,N_13045);
and U18518 (N_18518,N_14203,N_13868);
and U18519 (N_18519,N_11862,N_12664);
and U18520 (N_18520,N_12050,N_11914);
nor U18521 (N_18521,N_13310,N_12587);
nor U18522 (N_18522,N_10773,N_10257);
nand U18523 (N_18523,N_10590,N_10630);
xnor U18524 (N_18524,N_12465,N_12139);
xnor U18525 (N_18525,N_12630,N_12816);
or U18526 (N_18526,N_14166,N_14761);
or U18527 (N_18527,N_14575,N_13098);
and U18528 (N_18528,N_14902,N_13966);
xor U18529 (N_18529,N_11752,N_14392);
xnor U18530 (N_18530,N_12371,N_10417);
xnor U18531 (N_18531,N_10349,N_14982);
nand U18532 (N_18532,N_11441,N_13164);
nor U18533 (N_18533,N_12324,N_10435);
xor U18534 (N_18534,N_12379,N_11225);
or U18535 (N_18535,N_12289,N_12697);
xor U18536 (N_18536,N_11245,N_11474);
nor U18537 (N_18537,N_10189,N_10329);
nand U18538 (N_18538,N_12114,N_13189);
or U18539 (N_18539,N_12960,N_14506);
nand U18540 (N_18540,N_10590,N_12370);
nand U18541 (N_18541,N_11576,N_11953);
xor U18542 (N_18542,N_11704,N_14217);
or U18543 (N_18543,N_11850,N_10926);
or U18544 (N_18544,N_14940,N_10165);
xor U18545 (N_18545,N_10266,N_12876);
nor U18546 (N_18546,N_12771,N_14272);
nor U18547 (N_18547,N_13366,N_14239);
or U18548 (N_18548,N_14985,N_14895);
or U18549 (N_18549,N_14670,N_12288);
xnor U18550 (N_18550,N_12575,N_13292);
nand U18551 (N_18551,N_13888,N_13433);
xnor U18552 (N_18552,N_13240,N_12342);
nand U18553 (N_18553,N_12750,N_14219);
or U18554 (N_18554,N_10733,N_10952);
and U18555 (N_18555,N_12994,N_10389);
or U18556 (N_18556,N_11482,N_10271);
xor U18557 (N_18557,N_13020,N_11017);
xor U18558 (N_18558,N_14813,N_14133);
and U18559 (N_18559,N_13322,N_12592);
and U18560 (N_18560,N_14065,N_11473);
or U18561 (N_18561,N_11063,N_10285);
or U18562 (N_18562,N_13189,N_14426);
xnor U18563 (N_18563,N_14480,N_12809);
nor U18564 (N_18564,N_12385,N_14740);
xnor U18565 (N_18565,N_12297,N_11955);
nor U18566 (N_18566,N_13584,N_14802);
or U18567 (N_18567,N_14628,N_14559);
or U18568 (N_18568,N_13216,N_13251);
or U18569 (N_18569,N_14822,N_13204);
nand U18570 (N_18570,N_13157,N_14274);
nor U18571 (N_18571,N_12964,N_10923);
nand U18572 (N_18572,N_13512,N_14858);
and U18573 (N_18573,N_14209,N_13058);
nor U18574 (N_18574,N_12271,N_13691);
nand U18575 (N_18575,N_11074,N_14104);
xor U18576 (N_18576,N_10907,N_11672);
nand U18577 (N_18577,N_14074,N_10865);
nor U18578 (N_18578,N_10244,N_10577);
or U18579 (N_18579,N_14088,N_12096);
nand U18580 (N_18580,N_10164,N_13596);
nor U18581 (N_18581,N_12242,N_14053);
xnor U18582 (N_18582,N_13884,N_12337);
xor U18583 (N_18583,N_14241,N_11206);
xnor U18584 (N_18584,N_14890,N_14954);
xor U18585 (N_18585,N_14959,N_11076);
nand U18586 (N_18586,N_10470,N_13486);
nor U18587 (N_18587,N_13517,N_13012);
and U18588 (N_18588,N_12664,N_12357);
xor U18589 (N_18589,N_14009,N_14673);
and U18590 (N_18590,N_14538,N_13225);
nand U18591 (N_18591,N_11778,N_11105);
nor U18592 (N_18592,N_13761,N_10028);
xnor U18593 (N_18593,N_13369,N_10040);
or U18594 (N_18594,N_13594,N_11930);
or U18595 (N_18595,N_10958,N_10566);
and U18596 (N_18596,N_12435,N_13442);
and U18597 (N_18597,N_14803,N_14244);
nor U18598 (N_18598,N_14039,N_13199);
xnor U18599 (N_18599,N_13482,N_13526);
nor U18600 (N_18600,N_11946,N_10836);
and U18601 (N_18601,N_12693,N_14942);
and U18602 (N_18602,N_14310,N_10628);
nor U18603 (N_18603,N_14235,N_12443);
or U18604 (N_18604,N_14539,N_13675);
nor U18605 (N_18605,N_13172,N_14138);
nor U18606 (N_18606,N_13757,N_11575);
nand U18607 (N_18607,N_10589,N_13163);
nor U18608 (N_18608,N_13041,N_12321);
nand U18609 (N_18609,N_10621,N_10740);
and U18610 (N_18610,N_10632,N_13327);
nor U18611 (N_18611,N_10977,N_12427);
and U18612 (N_18612,N_10819,N_14939);
nand U18613 (N_18613,N_11188,N_11791);
and U18614 (N_18614,N_11923,N_14369);
nor U18615 (N_18615,N_12902,N_12157);
nor U18616 (N_18616,N_14486,N_13107);
nor U18617 (N_18617,N_10807,N_14913);
or U18618 (N_18618,N_11456,N_10602);
nor U18619 (N_18619,N_12361,N_11937);
or U18620 (N_18620,N_12805,N_11185);
nor U18621 (N_18621,N_11901,N_11957);
xnor U18622 (N_18622,N_11121,N_14725);
nor U18623 (N_18623,N_10825,N_11114);
nor U18624 (N_18624,N_10601,N_13425);
nand U18625 (N_18625,N_10944,N_14348);
and U18626 (N_18626,N_14937,N_11645);
or U18627 (N_18627,N_12149,N_12720);
and U18628 (N_18628,N_10161,N_10578);
nor U18629 (N_18629,N_13222,N_12176);
xor U18630 (N_18630,N_13481,N_12798);
nor U18631 (N_18631,N_13849,N_12850);
nor U18632 (N_18632,N_13406,N_13279);
nor U18633 (N_18633,N_14416,N_13176);
nand U18634 (N_18634,N_14545,N_13274);
nor U18635 (N_18635,N_10232,N_10519);
nand U18636 (N_18636,N_10112,N_14302);
nor U18637 (N_18637,N_14424,N_11445);
nor U18638 (N_18638,N_14144,N_14659);
and U18639 (N_18639,N_13112,N_13078);
xor U18640 (N_18640,N_13668,N_10031);
and U18641 (N_18641,N_13955,N_10161);
or U18642 (N_18642,N_12230,N_13995);
nand U18643 (N_18643,N_11797,N_10404);
and U18644 (N_18644,N_13031,N_11342);
xnor U18645 (N_18645,N_13119,N_12212);
or U18646 (N_18646,N_11612,N_10097);
and U18647 (N_18647,N_11147,N_12420);
xor U18648 (N_18648,N_11006,N_12854);
and U18649 (N_18649,N_13509,N_12029);
nand U18650 (N_18650,N_10349,N_14789);
nand U18651 (N_18651,N_12718,N_14958);
and U18652 (N_18652,N_11751,N_12423);
and U18653 (N_18653,N_11236,N_10663);
and U18654 (N_18654,N_14669,N_13973);
nor U18655 (N_18655,N_12478,N_13769);
nand U18656 (N_18656,N_13992,N_11265);
nor U18657 (N_18657,N_13685,N_13105);
and U18658 (N_18658,N_11638,N_13788);
nor U18659 (N_18659,N_14300,N_14592);
and U18660 (N_18660,N_11424,N_10135);
xnor U18661 (N_18661,N_11878,N_12758);
xor U18662 (N_18662,N_10492,N_11296);
xnor U18663 (N_18663,N_14941,N_12069);
nand U18664 (N_18664,N_14084,N_11266);
or U18665 (N_18665,N_10162,N_14484);
and U18666 (N_18666,N_12662,N_13670);
xor U18667 (N_18667,N_13363,N_11534);
xor U18668 (N_18668,N_10827,N_11103);
nand U18669 (N_18669,N_14308,N_12429);
or U18670 (N_18670,N_13508,N_13305);
and U18671 (N_18671,N_11548,N_10399);
nand U18672 (N_18672,N_13760,N_13683);
xnor U18673 (N_18673,N_10117,N_10070);
nand U18674 (N_18674,N_12075,N_11486);
and U18675 (N_18675,N_11863,N_10146);
nor U18676 (N_18676,N_12064,N_13580);
and U18677 (N_18677,N_10133,N_12278);
and U18678 (N_18678,N_13946,N_13321);
xor U18679 (N_18679,N_10894,N_12327);
nor U18680 (N_18680,N_10134,N_14365);
and U18681 (N_18681,N_13027,N_10972);
nor U18682 (N_18682,N_14187,N_10639);
xor U18683 (N_18683,N_13184,N_10564);
nand U18684 (N_18684,N_12914,N_13826);
xnor U18685 (N_18685,N_14248,N_13018);
xor U18686 (N_18686,N_14469,N_10769);
nor U18687 (N_18687,N_12484,N_13237);
and U18688 (N_18688,N_12139,N_13387);
and U18689 (N_18689,N_13569,N_14283);
nor U18690 (N_18690,N_12220,N_13369);
and U18691 (N_18691,N_10598,N_13208);
xor U18692 (N_18692,N_14632,N_14391);
and U18693 (N_18693,N_12202,N_13426);
xor U18694 (N_18694,N_11215,N_14214);
or U18695 (N_18695,N_11138,N_10464);
nand U18696 (N_18696,N_13158,N_14575);
xnor U18697 (N_18697,N_14279,N_13809);
nand U18698 (N_18698,N_14744,N_12352);
or U18699 (N_18699,N_13064,N_10765);
nor U18700 (N_18700,N_12457,N_11787);
and U18701 (N_18701,N_12045,N_14154);
nor U18702 (N_18702,N_13861,N_12394);
or U18703 (N_18703,N_13292,N_11567);
and U18704 (N_18704,N_10274,N_10067);
xor U18705 (N_18705,N_12623,N_11803);
xor U18706 (N_18706,N_14860,N_12756);
xnor U18707 (N_18707,N_13559,N_14995);
nor U18708 (N_18708,N_11494,N_14732);
xor U18709 (N_18709,N_11285,N_13447);
nor U18710 (N_18710,N_14747,N_13308);
xor U18711 (N_18711,N_14088,N_12716);
nand U18712 (N_18712,N_12145,N_11205);
and U18713 (N_18713,N_13659,N_10403);
or U18714 (N_18714,N_10424,N_13475);
or U18715 (N_18715,N_12556,N_14272);
nand U18716 (N_18716,N_14011,N_11991);
or U18717 (N_18717,N_14368,N_12033);
nand U18718 (N_18718,N_12191,N_14393);
or U18719 (N_18719,N_10150,N_14895);
and U18720 (N_18720,N_14748,N_12892);
and U18721 (N_18721,N_11688,N_11376);
nand U18722 (N_18722,N_12262,N_14539);
nor U18723 (N_18723,N_12263,N_11957);
xnor U18724 (N_18724,N_10851,N_11959);
nor U18725 (N_18725,N_12768,N_10372);
or U18726 (N_18726,N_12905,N_11232);
and U18727 (N_18727,N_11990,N_13078);
or U18728 (N_18728,N_14652,N_14535);
or U18729 (N_18729,N_12208,N_12792);
nor U18730 (N_18730,N_11203,N_12943);
xor U18731 (N_18731,N_14338,N_12007);
nor U18732 (N_18732,N_11627,N_14669);
nand U18733 (N_18733,N_11892,N_12461);
and U18734 (N_18734,N_10772,N_12516);
or U18735 (N_18735,N_11101,N_14742);
xnor U18736 (N_18736,N_13445,N_10715);
xor U18737 (N_18737,N_12643,N_14885);
xnor U18738 (N_18738,N_11432,N_10094);
nand U18739 (N_18739,N_12635,N_14302);
or U18740 (N_18740,N_11724,N_14309);
nor U18741 (N_18741,N_10475,N_11640);
nand U18742 (N_18742,N_12503,N_11427);
nand U18743 (N_18743,N_12617,N_10990);
nor U18744 (N_18744,N_14844,N_13322);
xor U18745 (N_18745,N_14623,N_11268);
or U18746 (N_18746,N_14186,N_13723);
nor U18747 (N_18747,N_13798,N_10592);
and U18748 (N_18748,N_11003,N_14967);
xnor U18749 (N_18749,N_14976,N_12785);
and U18750 (N_18750,N_11471,N_11043);
and U18751 (N_18751,N_14402,N_13152);
nand U18752 (N_18752,N_13101,N_11163);
or U18753 (N_18753,N_13972,N_11402);
xor U18754 (N_18754,N_14219,N_10197);
and U18755 (N_18755,N_13885,N_11029);
or U18756 (N_18756,N_11125,N_13940);
nand U18757 (N_18757,N_12195,N_10409);
xor U18758 (N_18758,N_10378,N_11812);
and U18759 (N_18759,N_14514,N_10691);
nand U18760 (N_18760,N_10217,N_10312);
or U18761 (N_18761,N_13412,N_14489);
nor U18762 (N_18762,N_12950,N_13032);
xor U18763 (N_18763,N_10252,N_10272);
nor U18764 (N_18764,N_10293,N_12961);
or U18765 (N_18765,N_13262,N_12632);
nand U18766 (N_18766,N_12857,N_11688);
xor U18767 (N_18767,N_11241,N_11974);
nor U18768 (N_18768,N_11642,N_14728);
or U18769 (N_18769,N_13562,N_12763);
nand U18770 (N_18770,N_13240,N_13608);
xnor U18771 (N_18771,N_12235,N_11145);
or U18772 (N_18772,N_13915,N_10413);
and U18773 (N_18773,N_12768,N_14154);
xor U18774 (N_18774,N_14212,N_12823);
or U18775 (N_18775,N_12200,N_11661);
and U18776 (N_18776,N_12391,N_10060);
or U18777 (N_18777,N_11856,N_12886);
nor U18778 (N_18778,N_13944,N_11868);
nor U18779 (N_18779,N_11543,N_13074);
xnor U18780 (N_18780,N_12280,N_14772);
nor U18781 (N_18781,N_10630,N_11496);
and U18782 (N_18782,N_10018,N_13404);
nand U18783 (N_18783,N_14948,N_11731);
and U18784 (N_18784,N_12769,N_11148);
xor U18785 (N_18785,N_10460,N_12486);
xor U18786 (N_18786,N_13257,N_14815);
xnor U18787 (N_18787,N_13145,N_14561);
nor U18788 (N_18788,N_12066,N_14338);
or U18789 (N_18789,N_10191,N_14888);
nand U18790 (N_18790,N_11085,N_14497);
nor U18791 (N_18791,N_10258,N_13239);
nand U18792 (N_18792,N_14530,N_11221);
or U18793 (N_18793,N_11141,N_10493);
nand U18794 (N_18794,N_12741,N_10248);
or U18795 (N_18795,N_14967,N_11565);
or U18796 (N_18796,N_14627,N_10875);
and U18797 (N_18797,N_11398,N_10884);
nand U18798 (N_18798,N_14177,N_14120);
xnor U18799 (N_18799,N_11976,N_12643);
xnor U18800 (N_18800,N_12529,N_13154);
nand U18801 (N_18801,N_10178,N_14419);
xor U18802 (N_18802,N_14441,N_12155);
nand U18803 (N_18803,N_10925,N_13127);
nor U18804 (N_18804,N_10708,N_10003);
and U18805 (N_18805,N_13327,N_11490);
or U18806 (N_18806,N_11399,N_12441);
and U18807 (N_18807,N_14125,N_10970);
and U18808 (N_18808,N_12167,N_14839);
and U18809 (N_18809,N_14319,N_11987);
nor U18810 (N_18810,N_11025,N_11166);
xnor U18811 (N_18811,N_13543,N_10588);
or U18812 (N_18812,N_10212,N_10897);
and U18813 (N_18813,N_10716,N_13362);
nor U18814 (N_18814,N_11323,N_12293);
nand U18815 (N_18815,N_14241,N_12934);
or U18816 (N_18816,N_12433,N_14739);
and U18817 (N_18817,N_14573,N_10049);
nand U18818 (N_18818,N_14333,N_14847);
and U18819 (N_18819,N_12572,N_14858);
nor U18820 (N_18820,N_13824,N_11051);
nand U18821 (N_18821,N_14638,N_11630);
and U18822 (N_18822,N_12162,N_10224);
and U18823 (N_18823,N_13544,N_11205);
nand U18824 (N_18824,N_12016,N_11886);
nand U18825 (N_18825,N_12808,N_10995);
xnor U18826 (N_18826,N_11523,N_10739);
and U18827 (N_18827,N_14512,N_11678);
nand U18828 (N_18828,N_12145,N_14360);
and U18829 (N_18829,N_13023,N_10820);
or U18830 (N_18830,N_13146,N_12563);
nor U18831 (N_18831,N_14852,N_11589);
xor U18832 (N_18832,N_11358,N_14749);
nand U18833 (N_18833,N_10666,N_11924);
xor U18834 (N_18834,N_14725,N_10554);
nand U18835 (N_18835,N_10158,N_11242);
or U18836 (N_18836,N_14024,N_13937);
nand U18837 (N_18837,N_12690,N_10996);
nor U18838 (N_18838,N_14623,N_10097);
and U18839 (N_18839,N_14177,N_10455);
nor U18840 (N_18840,N_11077,N_13290);
nor U18841 (N_18841,N_13866,N_11816);
or U18842 (N_18842,N_12286,N_13906);
xor U18843 (N_18843,N_14742,N_13860);
and U18844 (N_18844,N_13574,N_13947);
nand U18845 (N_18845,N_10854,N_10018);
nor U18846 (N_18846,N_10637,N_11979);
and U18847 (N_18847,N_12380,N_14851);
nand U18848 (N_18848,N_13793,N_13522);
nand U18849 (N_18849,N_13724,N_13638);
and U18850 (N_18850,N_10195,N_12612);
nand U18851 (N_18851,N_11234,N_10794);
nand U18852 (N_18852,N_14724,N_11990);
or U18853 (N_18853,N_10645,N_13138);
and U18854 (N_18854,N_10886,N_13422);
nor U18855 (N_18855,N_13520,N_11460);
nor U18856 (N_18856,N_13937,N_10073);
xor U18857 (N_18857,N_13628,N_10808);
and U18858 (N_18858,N_13017,N_12417);
nor U18859 (N_18859,N_14243,N_11567);
and U18860 (N_18860,N_13014,N_13066);
or U18861 (N_18861,N_11615,N_14458);
nand U18862 (N_18862,N_12944,N_12714);
nand U18863 (N_18863,N_13207,N_10245);
nor U18864 (N_18864,N_12356,N_12360);
nor U18865 (N_18865,N_14018,N_14270);
xor U18866 (N_18866,N_10311,N_10392);
xnor U18867 (N_18867,N_10378,N_10598);
nor U18868 (N_18868,N_14768,N_10291);
and U18869 (N_18869,N_12216,N_12590);
nor U18870 (N_18870,N_11700,N_11663);
and U18871 (N_18871,N_13362,N_11027);
and U18872 (N_18872,N_12750,N_14001);
or U18873 (N_18873,N_13562,N_11537);
nand U18874 (N_18874,N_11785,N_14370);
xnor U18875 (N_18875,N_10296,N_11290);
nor U18876 (N_18876,N_11648,N_12835);
xor U18877 (N_18877,N_12364,N_10243);
or U18878 (N_18878,N_10594,N_10956);
nor U18879 (N_18879,N_13255,N_12474);
nand U18880 (N_18880,N_14672,N_11659);
and U18881 (N_18881,N_10172,N_13912);
nand U18882 (N_18882,N_14900,N_11350);
nor U18883 (N_18883,N_11828,N_11665);
nand U18884 (N_18884,N_14395,N_10286);
nor U18885 (N_18885,N_12373,N_10830);
nand U18886 (N_18886,N_13005,N_13929);
and U18887 (N_18887,N_13005,N_11022);
nand U18888 (N_18888,N_11269,N_14165);
xnor U18889 (N_18889,N_10009,N_14398);
and U18890 (N_18890,N_12640,N_12890);
or U18891 (N_18891,N_13081,N_12188);
or U18892 (N_18892,N_13718,N_14588);
and U18893 (N_18893,N_11645,N_13364);
nor U18894 (N_18894,N_11508,N_14822);
nor U18895 (N_18895,N_12275,N_11609);
or U18896 (N_18896,N_14644,N_11209);
and U18897 (N_18897,N_13486,N_10049);
nand U18898 (N_18898,N_13455,N_13702);
nand U18899 (N_18899,N_11432,N_14133);
or U18900 (N_18900,N_10184,N_10761);
nor U18901 (N_18901,N_14269,N_13919);
and U18902 (N_18902,N_10011,N_12967);
or U18903 (N_18903,N_14065,N_11153);
or U18904 (N_18904,N_11387,N_10156);
xnor U18905 (N_18905,N_10735,N_14618);
nand U18906 (N_18906,N_14845,N_10985);
xnor U18907 (N_18907,N_11284,N_10158);
or U18908 (N_18908,N_10911,N_13406);
nand U18909 (N_18909,N_13198,N_12025);
nor U18910 (N_18910,N_12681,N_12655);
and U18911 (N_18911,N_12465,N_12097);
nand U18912 (N_18912,N_12815,N_13987);
and U18913 (N_18913,N_10538,N_12646);
and U18914 (N_18914,N_14691,N_10105);
and U18915 (N_18915,N_13800,N_12655);
or U18916 (N_18916,N_12972,N_14881);
or U18917 (N_18917,N_12223,N_13090);
xnor U18918 (N_18918,N_11298,N_10112);
nand U18919 (N_18919,N_14384,N_12083);
nor U18920 (N_18920,N_14142,N_11817);
nor U18921 (N_18921,N_14268,N_10275);
or U18922 (N_18922,N_14358,N_12285);
xnor U18923 (N_18923,N_12431,N_10780);
or U18924 (N_18924,N_14296,N_13900);
nor U18925 (N_18925,N_12077,N_11219);
or U18926 (N_18926,N_14814,N_11116);
or U18927 (N_18927,N_11631,N_12192);
and U18928 (N_18928,N_14896,N_12150);
and U18929 (N_18929,N_10574,N_14332);
xnor U18930 (N_18930,N_14702,N_11668);
nand U18931 (N_18931,N_10245,N_13922);
nand U18932 (N_18932,N_11687,N_11467);
nand U18933 (N_18933,N_12804,N_14167);
or U18934 (N_18934,N_10074,N_14342);
and U18935 (N_18935,N_10449,N_14166);
and U18936 (N_18936,N_11569,N_13496);
nor U18937 (N_18937,N_14800,N_12675);
xor U18938 (N_18938,N_13663,N_13348);
nand U18939 (N_18939,N_14125,N_10588);
xor U18940 (N_18940,N_14396,N_14937);
or U18941 (N_18941,N_13498,N_14098);
and U18942 (N_18942,N_14044,N_12260);
and U18943 (N_18943,N_12621,N_14675);
and U18944 (N_18944,N_13518,N_14706);
xnor U18945 (N_18945,N_13306,N_11091);
and U18946 (N_18946,N_13748,N_12633);
xnor U18947 (N_18947,N_10275,N_11310);
or U18948 (N_18948,N_13677,N_12840);
or U18949 (N_18949,N_12927,N_14035);
nor U18950 (N_18950,N_13650,N_11896);
xor U18951 (N_18951,N_13755,N_10974);
nor U18952 (N_18952,N_10429,N_14725);
nor U18953 (N_18953,N_14275,N_10842);
nor U18954 (N_18954,N_11236,N_10324);
xnor U18955 (N_18955,N_10883,N_13233);
nand U18956 (N_18956,N_11586,N_14238);
xor U18957 (N_18957,N_14993,N_12118);
nor U18958 (N_18958,N_10563,N_12417);
and U18959 (N_18959,N_14735,N_10213);
nand U18960 (N_18960,N_11896,N_11323);
and U18961 (N_18961,N_11621,N_13888);
and U18962 (N_18962,N_13676,N_11139);
or U18963 (N_18963,N_10251,N_13481);
nand U18964 (N_18964,N_13270,N_14738);
nand U18965 (N_18965,N_12332,N_14964);
xnor U18966 (N_18966,N_12950,N_13730);
nor U18967 (N_18967,N_14304,N_10980);
nand U18968 (N_18968,N_13912,N_11874);
nand U18969 (N_18969,N_13746,N_14104);
xor U18970 (N_18970,N_13124,N_12051);
nand U18971 (N_18971,N_13892,N_10125);
xor U18972 (N_18972,N_14231,N_13971);
xnor U18973 (N_18973,N_11464,N_14490);
nand U18974 (N_18974,N_13387,N_13853);
or U18975 (N_18975,N_12267,N_10827);
or U18976 (N_18976,N_12324,N_11591);
or U18977 (N_18977,N_13071,N_10539);
or U18978 (N_18978,N_14975,N_10990);
or U18979 (N_18979,N_12703,N_13998);
nand U18980 (N_18980,N_10489,N_13885);
nor U18981 (N_18981,N_13028,N_11876);
and U18982 (N_18982,N_14003,N_14065);
nand U18983 (N_18983,N_13263,N_13738);
nor U18984 (N_18984,N_14591,N_12474);
and U18985 (N_18985,N_14226,N_12172);
nand U18986 (N_18986,N_13031,N_14337);
nand U18987 (N_18987,N_10073,N_12923);
xnor U18988 (N_18988,N_14015,N_10680);
xor U18989 (N_18989,N_14795,N_11234);
xnor U18990 (N_18990,N_12807,N_10848);
and U18991 (N_18991,N_12353,N_11995);
nor U18992 (N_18992,N_11938,N_10935);
or U18993 (N_18993,N_10248,N_12149);
or U18994 (N_18994,N_12515,N_10181);
nor U18995 (N_18995,N_11502,N_11467);
xnor U18996 (N_18996,N_14827,N_14795);
nor U18997 (N_18997,N_10276,N_14526);
or U18998 (N_18998,N_12808,N_13652);
nor U18999 (N_18999,N_10886,N_10187);
and U19000 (N_19000,N_13620,N_11152);
nand U19001 (N_19001,N_14922,N_10777);
nor U19002 (N_19002,N_13849,N_10331);
and U19003 (N_19003,N_14206,N_13896);
and U19004 (N_19004,N_13816,N_11395);
nand U19005 (N_19005,N_13495,N_13138);
or U19006 (N_19006,N_11852,N_14709);
nor U19007 (N_19007,N_10560,N_13988);
or U19008 (N_19008,N_14747,N_14717);
and U19009 (N_19009,N_14537,N_12978);
nand U19010 (N_19010,N_14707,N_11062);
nand U19011 (N_19011,N_13716,N_10551);
and U19012 (N_19012,N_12539,N_13391);
and U19013 (N_19013,N_11229,N_11137);
nand U19014 (N_19014,N_13679,N_13608);
xor U19015 (N_19015,N_11220,N_14738);
or U19016 (N_19016,N_14113,N_13848);
or U19017 (N_19017,N_11688,N_12902);
nand U19018 (N_19018,N_11145,N_10755);
nor U19019 (N_19019,N_12342,N_13276);
nand U19020 (N_19020,N_12740,N_14120);
nor U19021 (N_19021,N_12553,N_13370);
or U19022 (N_19022,N_10346,N_12332);
xnor U19023 (N_19023,N_13311,N_10015);
nand U19024 (N_19024,N_12641,N_11507);
or U19025 (N_19025,N_11812,N_10905);
or U19026 (N_19026,N_10085,N_11549);
and U19027 (N_19027,N_11536,N_14076);
xor U19028 (N_19028,N_13798,N_10178);
nor U19029 (N_19029,N_11534,N_10327);
and U19030 (N_19030,N_11663,N_13840);
or U19031 (N_19031,N_11189,N_11470);
nand U19032 (N_19032,N_12280,N_13699);
and U19033 (N_19033,N_14778,N_14756);
nor U19034 (N_19034,N_12234,N_11952);
nand U19035 (N_19035,N_10220,N_10934);
nor U19036 (N_19036,N_13275,N_13096);
and U19037 (N_19037,N_11836,N_13566);
or U19038 (N_19038,N_14695,N_13235);
xor U19039 (N_19039,N_12442,N_13288);
nor U19040 (N_19040,N_10037,N_11453);
or U19041 (N_19041,N_12267,N_11947);
xor U19042 (N_19042,N_13816,N_10449);
xor U19043 (N_19043,N_13006,N_11815);
nand U19044 (N_19044,N_12747,N_11818);
or U19045 (N_19045,N_13800,N_10138);
or U19046 (N_19046,N_12310,N_11092);
nand U19047 (N_19047,N_12404,N_14159);
nor U19048 (N_19048,N_12326,N_13094);
or U19049 (N_19049,N_11332,N_11383);
xnor U19050 (N_19050,N_11474,N_13152);
and U19051 (N_19051,N_14489,N_12558);
or U19052 (N_19052,N_11875,N_14128);
or U19053 (N_19053,N_10709,N_11891);
nor U19054 (N_19054,N_13878,N_12070);
or U19055 (N_19055,N_14857,N_13942);
and U19056 (N_19056,N_13600,N_13868);
or U19057 (N_19057,N_10539,N_11958);
nor U19058 (N_19058,N_13700,N_12569);
nor U19059 (N_19059,N_11960,N_14068);
and U19060 (N_19060,N_10568,N_11548);
nand U19061 (N_19061,N_11850,N_10869);
nand U19062 (N_19062,N_13744,N_12989);
xor U19063 (N_19063,N_11519,N_13611);
xnor U19064 (N_19064,N_12520,N_10969);
xor U19065 (N_19065,N_14394,N_14974);
xor U19066 (N_19066,N_10712,N_13713);
nor U19067 (N_19067,N_10177,N_11585);
nand U19068 (N_19068,N_14107,N_12244);
and U19069 (N_19069,N_13499,N_13992);
nor U19070 (N_19070,N_11690,N_14550);
xor U19071 (N_19071,N_13748,N_11963);
or U19072 (N_19072,N_11000,N_13410);
xnor U19073 (N_19073,N_14017,N_10731);
and U19074 (N_19074,N_13250,N_13043);
nand U19075 (N_19075,N_11076,N_11407);
or U19076 (N_19076,N_13939,N_10099);
xnor U19077 (N_19077,N_10369,N_12009);
or U19078 (N_19078,N_10971,N_14451);
and U19079 (N_19079,N_10919,N_11850);
nand U19080 (N_19080,N_11544,N_13784);
nor U19081 (N_19081,N_14110,N_12401);
and U19082 (N_19082,N_11756,N_10748);
nand U19083 (N_19083,N_11076,N_13808);
or U19084 (N_19084,N_12838,N_10366);
or U19085 (N_19085,N_13884,N_10712);
nand U19086 (N_19086,N_12939,N_13275);
and U19087 (N_19087,N_10853,N_14324);
nand U19088 (N_19088,N_13865,N_14620);
nor U19089 (N_19089,N_11133,N_12844);
nand U19090 (N_19090,N_11128,N_10357);
and U19091 (N_19091,N_10818,N_14279);
nor U19092 (N_19092,N_12723,N_11152);
xnor U19093 (N_19093,N_10283,N_14940);
nor U19094 (N_19094,N_13526,N_10269);
xnor U19095 (N_19095,N_12710,N_13346);
or U19096 (N_19096,N_11007,N_12928);
nor U19097 (N_19097,N_13028,N_12387);
or U19098 (N_19098,N_10318,N_11517);
and U19099 (N_19099,N_14106,N_11957);
or U19100 (N_19100,N_12534,N_13393);
nand U19101 (N_19101,N_12986,N_12513);
and U19102 (N_19102,N_10609,N_11269);
and U19103 (N_19103,N_14769,N_11267);
nor U19104 (N_19104,N_13271,N_14385);
nand U19105 (N_19105,N_10313,N_14038);
nor U19106 (N_19106,N_14009,N_10490);
or U19107 (N_19107,N_12891,N_14619);
xnor U19108 (N_19108,N_11071,N_11510);
and U19109 (N_19109,N_14036,N_12150);
xnor U19110 (N_19110,N_14261,N_14139);
or U19111 (N_19111,N_14769,N_13779);
and U19112 (N_19112,N_12364,N_10689);
nor U19113 (N_19113,N_10956,N_14873);
or U19114 (N_19114,N_14625,N_13942);
xor U19115 (N_19115,N_11760,N_11329);
xnor U19116 (N_19116,N_11007,N_14079);
or U19117 (N_19117,N_12302,N_10437);
nand U19118 (N_19118,N_10791,N_12299);
and U19119 (N_19119,N_11844,N_11356);
nand U19120 (N_19120,N_12132,N_11968);
and U19121 (N_19121,N_11598,N_11364);
xnor U19122 (N_19122,N_12800,N_14014);
nand U19123 (N_19123,N_10112,N_12598);
or U19124 (N_19124,N_12387,N_13511);
or U19125 (N_19125,N_11798,N_13973);
xnor U19126 (N_19126,N_13215,N_11415);
and U19127 (N_19127,N_12261,N_14815);
nand U19128 (N_19128,N_13290,N_13332);
xor U19129 (N_19129,N_13886,N_13428);
nor U19130 (N_19130,N_11915,N_11750);
xor U19131 (N_19131,N_14665,N_13808);
or U19132 (N_19132,N_12595,N_12692);
nand U19133 (N_19133,N_10964,N_10968);
nand U19134 (N_19134,N_12823,N_10830);
xor U19135 (N_19135,N_11266,N_12088);
and U19136 (N_19136,N_10261,N_10702);
nor U19137 (N_19137,N_14229,N_10716);
nor U19138 (N_19138,N_11466,N_11862);
or U19139 (N_19139,N_13462,N_12287);
nor U19140 (N_19140,N_12314,N_11770);
or U19141 (N_19141,N_12317,N_14708);
nand U19142 (N_19142,N_10180,N_14203);
and U19143 (N_19143,N_10632,N_11613);
and U19144 (N_19144,N_11685,N_11980);
and U19145 (N_19145,N_14651,N_12919);
or U19146 (N_19146,N_14809,N_11130);
nand U19147 (N_19147,N_12359,N_14512);
and U19148 (N_19148,N_11932,N_10157);
or U19149 (N_19149,N_11439,N_10364);
xor U19150 (N_19150,N_11369,N_12213);
nand U19151 (N_19151,N_13583,N_10949);
nor U19152 (N_19152,N_14692,N_13961);
or U19153 (N_19153,N_12066,N_12030);
and U19154 (N_19154,N_10780,N_11963);
nand U19155 (N_19155,N_10195,N_11361);
nand U19156 (N_19156,N_11167,N_14369);
or U19157 (N_19157,N_10032,N_12004);
nor U19158 (N_19158,N_14680,N_14517);
nand U19159 (N_19159,N_13208,N_13513);
and U19160 (N_19160,N_12231,N_12725);
xor U19161 (N_19161,N_10041,N_10343);
and U19162 (N_19162,N_12959,N_13210);
xor U19163 (N_19163,N_14024,N_12112);
nand U19164 (N_19164,N_11686,N_13702);
or U19165 (N_19165,N_10158,N_14411);
or U19166 (N_19166,N_14708,N_12052);
xor U19167 (N_19167,N_14142,N_11031);
nand U19168 (N_19168,N_12460,N_14813);
and U19169 (N_19169,N_14989,N_11909);
nor U19170 (N_19170,N_14900,N_12453);
or U19171 (N_19171,N_13947,N_10102);
and U19172 (N_19172,N_13234,N_12491);
or U19173 (N_19173,N_13322,N_14945);
xnor U19174 (N_19174,N_12591,N_10024);
nand U19175 (N_19175,N_14762,N_10452);
xor U19176 (N_19176,N_14582,N_11458);
nor U19177 (N_19177,N_14172,N_14042);
and U19178 (N_19178,N_12093,N_13645);
nor U19179 (N_19179,N_13229,N_11638);
or U19180 (N_19180,N_14508,N_10361);
nor U19181 (N_19181,N_13781,N_14683);
and U19182 (N_19182,N_13610,N_10666);
or U19183 (N_19183,N_11403,N_14533);
xor U19184 (N_19184,N_10483,N_14890);
nand U19185 (N_19185,N_11813,N_12993);
nand U19186 (N_19186,N_12394,N_10322);
xor U19187 (N_19187,N_10178,N_12881);
nand U19188 (N_19188,N_12261,N_13824);
or U19189 (N_19189,N_11333,N_12317);
and U19190 (N_19190,N_10985,N_11611);
or U19191 (N_19191,N_14083,N_14569);
nand U19192 (N_19192,N_14138,N_11558);
xor U19193 (N_19193,N_14982,N_13680);
or U19194 (N_19194,N_10828,N_10429);
nor U19195 (N_19195,N_12613,N_13572);
and U19196 (N_19196,N_14458,N_10440);
nand U19197 (N_19197,N_14718,N_12724);
nor U19198 (N_19198,N_12854,N_12989);
or U19199 (N_19199,N_13145,N_12304);
nor U19200 (N_19200,N_14740,N_10863);
xnor U19201 (N_19201,N_13571,N_11203);
and U19202 (N_19202,N_12053,N_12695);
xor U19203 (N_19203,N_10661,N_14577);
nand U19204 (N_19204,N_13592,N_12209);
and U19205 (N_19205,N_13957,N_14133);
nand U19206 (N_19206,N_10847,N_12104);
nand U19207 (N_19207,N_10637,N_10324);
xnor U19208 (N_19208,N_13106,N_14207);
or U19209 (N_19209,N_13242,N_11142);
xnor U19210 (N_19210,N_12906,N_14643);
nor U19211 (N_19211,N_10879,N_10217);
and U19212 (N_19212,N_14705,N_14767);
and U19213 (N_19213,N_12156,N_10383);
xor U19214 (N_19214,N_14201,N_13153);
nand U19215 (N_19215,N_11295,N_14734);
xor U19216 (N_19216,N_14114,N_11274);
and U19217 (N_19217,N_11433,N_12829);
nor U19218 (N_19218,N_13444,N_14875);
nand U19219 (N_19219,N_14871,N_10022);
xnor U19220 (N_19220,N_14052,N_11903);
nand U19221 (N_19221,N_12372,N_10594);
or U19222 (N_19222,N_12949,N_13861);
nand U19223 (N_19223,N_13798,N_10868);
and U19224 (N_19224,N_12735,N_12301);
and U19225 (N_19225,N_13732,N_10090);
and U19226 (N_19226,N_10799,N_10218);
or U19227 (N_19227,N_14416,N_13475);
nand U19228 (N_19228,N_12068,N_13606);
and U19229 (N_19229,N_11089,N_14769);
or U19230 (N_19230,N_12222,N_13609);
nand U19231 (N_19231,N_14221,N_14479);
or U19232 (N_19232,N_14467,N_12777);
xnor U19233 (N_19233,N_12143,N_13813);
or U19234 (N_19234,N_13588,N_12154);
xnor U19235 (N_19235,N_11201,N_11017);
or U19236 (N_19236,N_10707,N_12996);
xor U19237 (N_19237,N_11844,N_13164);
and U19238 (N_19238,N_10288,N_10633);
nor U19239 (N_19239,N_10780,N_11767);
nor U19240 (N_19240,N_14957,N_10511);
xor U19241 (N_19241,N_10005,N_13834);
or U19242 (N_19242,N_10677,N_10763);
xor U19243 (N_19243,N_12656,N_10581);
nor U19244 (N_19244,N_13451,N_13752);
nand U19245 (N_19245,N_10724,N_13503);
or U19246 (N_19246,N_13697,N_12418);
nor U19247 (N_19247,N_12326,N_13051);
or U19248 (N_19248,N_11980,N_12052);
xor U19249 (N_19249,N_14703,N_14245);
nand U19250 (N_19250,N_10464,N_14244);
and U19251 (N_19251,N_11149,N_13172);
xnor U19252 (N_19252,N_10896,N_10613);
and U19253 (N_19253,N_10033,N_13450);
and U19254 (N_19254,N_11141,N_11515);
xor U19255 (N_19255,N_12926,N_10890);
xnor U19256 (N_19256,N_13840,N_11271);
nor U19257 (N_19257,N_12307,N_10796);
or U19258 (N_19258,N_13782,N_12926);
nor U19259 (N_19259,N_13408,N_13070);
or U19260 (N_19260,N_14424,N_11979);
and U19261 (N_19261,N_14223,N_14220);
xor U19262 (N_19262,N_12815,N_13093);
nor U19263 (N_19263,N_11567,N_10675);
nor U19264 (N_19264,N_14402,N_13965);
nor U19265 (N_19265,N_12394,N_12886);
xor U19266 (N_19266,N_11577,N_14522);
nand U19267 (N_19267,N_12133,N_10382);
nor U19268 (N_19268,N_10502,N_10000);
nand U19269 (N_19269,N_12435,N_13339);
and U19270 (N_19270,N_14689,N_10523);
or U19271 (N_19271,N_12457,N_12445);
or U19272 (N_19272,N_11232,N_13351);
nor U19273 (N_19273,N_13572,N_13406);
nor U19274 (N_19274,N_10452,N_13261);
nor U19275 (N_19275,N_13579,N_13149);
and U19276 (N_19276,N_13917,N_13352);
nand U19277 (N_19277,N_13329,N_13874);
nor U19278 (N_19278,N_10726,N_11363);
nand U19279 (N_19279,N_13097,N_10922);
or U19280 (N_19280,N_10309,N_10467);
or U19281 (N_19281,N_14314,N_10868);
nand U19282 (N_19282,N_10146,N_10844);
nand U19283 (N_19283,N_11092,N_14694);
xnor U19284 (N_19284,N_13452,N_14865);
xor U19285 (N_19285,N_11280,N_12221);
nor U19286 (N_19286,N_12576,N_14242);
nand U19287 (N_19287,N_10111,N_11532);
nor U19288 (N_19288,N_10621,N_11524);
nor U19289 (N_19289,N_12550,N_12124);
nand U19290 (N_19290,N_14003,N_10813);
xnor U19291 (N_19291,N_13112,N_14049);
nor U19292 (N_19292,N_13076,N_11046);
or U19293 (N_19293,N_13056,N_11052);
or U19294 (N_19294,N_13840,N_12675);
nor U19295 (N_19295,N_13852,N_11019);
nor U19296 (N_19296,N_11144,N_14220);
nand U19297 (N_19297,N_13341,N_14412);
xnor U19298 (N_19298,N_10890,N_13014);
xor U19299 (N_19299,N_12370,N_13189);
or U19300 (N_19300,N_11703,N_11791);
nor U19301 (N_19301,N_11739,N_13515);
and U19302 (N_19302,N_11180,N_11123);
and U19303 (N_19303,N_11876,N_14381);
nand U19304 (N_19304,N_11962,N_10909);
nor U19305 (N_19305,N_10227,N_10558);
nand U19306 (N_19306,N_10320,N_14919);
xor U19307 (N_19307,N_11401,N_12917);
xor U19308 (N_19308,N_10929,N_12528);
or U19309 (N_19309,N_13401,N_11767);
xnor U19310 (N_19310,N_10874,N_11414);
and U19311 (N_19311,N_14491,N_13611);
or U19312 (N_19312,N_14658,N_14966);
and U19313 (N_19313,N_13743,N_11773);
and U19314 (N_19314,N_10284,N_13688);
xor U19315 (N_19315,N_11537,N_10159);
or U19316 (N_19316,N_12030,N_12827);
and U19317 (N_19317,N_11574,N_14986);
nand U19318 (N_19318,N_10163,N_10849);
or U19319 (N_19319,N_14815,N_12556);
nand U19320 (N_19320,N_11081,N_11194);
or U19321 (N_19321,N_14870,N_11066);
or U19322 (N_19322,N_13081,N_10031);
and U19323 (N_19323,N_14879,N_11442);
nand U19324 (N_19324,N_12427,N_14724);
and U19325 (N_19325,N_12340,N_12450);
xnor U19326 (N_19326,N_13918,N_13950);
and U19327 (N_19327,N_13207,N_10645);
and U19328 (N_19328,N_14990,N_13918);
nor U19329 (N_19329,N_13828,N_12676);
xor U19330 (N_19330,N_13701,N_14329);
and U19331 (N_19331,N_12961,N_14156);
or U19332 (N_19332,N_11244,N_14728);
and U19333 (N_19333,N_11822,N_11052);
nor U19334 (N_19334,N_13513,N_11037);
nor U19335 (N_19335,N_13184,N_11227);
and U19336 (N_19336,N_10314,N_14728);
nor U19337 (N_19337,N_12478,N_14010);
nand U19338 (N_19338,N_13956,N_11689);
or U19339 (N_19339,N_13410,N_14579);
nand U19340 (N_19340,N_13720,N_10255);
or U19341 (N_19341,N_13426,N_14774);
or U19342 (N_19342,N_10262,N_10564);
xor U19343 (N_19343,N_14481,N_14380);
nand U19344 (N_19344,N_12441,N_12773);
or U19345 (N_19345,N_10748,N_14204);
nor U19346 (N_19346,N_10016,N_12698);
and U19347 (N_19347,N_10410,N_12496);
or U19348 (N_19348,N_10384,N_11567);
or U19349 (N_19349,N_10416,N_11796);
nand U19350 (N_19350,N_13041,N_11368);
nand U19351 (N_19351,N_11286,N_13364);
nor U19352 (N_19352,N_13404,N_14224);
nor U19353 (N_19353,N_10789,N_14476);
and U19354 (N_19354,N_13387,N_10101);
and U19355 (N_19355,N_10382,N_12943);
nor U19356 (N_19356,N_12000,N_11790);
or U19357 (N_19357,N_11564,N_14681);
nand U19358 (N_19358,N_11779,N_14638);
nor U19359 (N_19359,N_10285,N_13291);
or U19360 (N_19360,N_14146,N_11034);
and U19361 (N_19361,N_13822,N_13760);
nor U19362 (N_19362,N_13328,N_12205);
and U19363 (N_19363,N_11525,N_13530);
nor U19364 (N_19364,N_12419,N_13743);
nor U19365 (N_19365,N_12662,N_11002);
or U19366 (N_19366,N_12135,N_12485);
nor U19367 (N_19367,N_12232,N_11835);
xnor U19368 (N_19368,N_14829,N_11443);
or U19369 (N_19369,N_11726,N_12525);
and U19370 (N_19370,N_11727,N_10385);
and U19371 (N_19371,N_12415,N_14273);
or U19372 (N_19372,N_11307,N_12108);
xnor U19373 (N_19373,N_12956,N_12914);
nor U19374 (N_19374,N_14637,N_11178);
xor U19375 (N_19375,N_12359,N_11900);
nand U19376 (N_19376,N_14540,N_12828);
xnor U19377 (N_19377,N_11856,N_11721);
nand U19378 (N_19378,N_11410,N_14994);
or U19379 (N_19379,N_14153,N_14884);
nor U19380 (N_19380,N_14031,N_13110);
xor U19381 (N_19381,N_14528,N_11289);
nor U19382 (N_19382,N_10050,N_13473);
xnor U19383 (N_19383,N_12465,N_12423);
nand U19384 (N_19384,N_10114,N_13405);
or U19385 (N_19385,N_12461,N_11598);
nand U19386 (N_19386,N_11880,N_10770);
xnor U19387 (N_19387,N_14166,N_10769);
and U19388 (N_19388,N_11745,N_13063);
nand U19389 (N_19389,N_14240,N_13659);
nor U19390 (N_19390,N_13065,N_11339);
or U19391 (N_19391,N_14150,N_13311);
nor U19392 (N_19392,N_11524,N_10994);
and U19393 (N_19393,N_12368,N_10624);
and U19394 (N_19394,N_12354,N_14539);
nor U19395 (N_19395,N_11281,N_13920);
and U19396 (N_19396,N_12027,N_14798);
or U19397 (N_19397,N_12738,N_12787);
and U19398 (N_19398,N_13045,N_10415);
or U19399 (N_19399,N_10723,N_11370);
and U19400 (N_19400,N_10633,N_10688);
or U19401 (N_19401,N_11730,N_11605);
nor U19402 (N_19402,N_13771,N_14092);
and U19403 (N_19403,N_12771,N_12667);
xor U19404 (N_19404,N_10003,N_13649);
or U19405 (N_19405,N_10496,N_12253);
nor U19406 (N_19406,N_12391,N_13675);
xnor U19407 (N_19407,N_14707,N_14405);
and U19408 (N_19408,N_11971,N_11469);
and U19409 (N_19409,N_11370,N_11088);
xnor U19410 (N_19410,N_13208,N_10507);
nand U19411 (N_19411,N_11251,N_14061);
or U19412 (N_19412,N_10648,N_11296);
nor U19413 (N_19413,N_13819,N_12745);
or U19414 (N_19414,N_14609,N_11781);
and U19415 (N_19415,N_13752,N_13642);
nand U19416 (N_19416,N_14954,N_11738);
or U19417 (N_19417,N_12000,N_12882);
nor U19418 (N_19418,N_10662,N_10358);
nor U19419 (N_19419,N_10281,N_14018);
and U19420 (N_19420,N_10555,N_10568);
xnor U19421 (N_19421,N_10289,N_13885);
and U19422 (N_19422,N_11967,N_14412);
or U19423 (N_19423,N_13574,N_11544);
nand U19424 (N_19424,N_10298,N_14623);
nand U19425 (N_19425,N_10539,N_14133);
or U19426 (N_19426,N_11216,N_11256);
or U19427 (N_19427,N_14946,N_12304);
and U19428 (N_19428,N_12462,N_10732);
xnor U19429 (N_19429,N_14459,N_14214);
xor U19430 (N_19430,N_11728,N_14231);
or U19431 (N_19431,N_12075,N_11738);
and U19432 (N_19432,N_10492,N_12547);
nand U19433 (N_19433,N_13035,N_13557);
and U19434 (N_19434,N_10451,N_14426);
nand U19435 (N_19435,N_13376,N_11929);
nor U19436 (N_19436,N_13167,N_14362);
nor U19437 (N_19437,N_13234,N_12248);
nor U19438 (N_19438,N_10679,N_12694);
nor U19439 (N_19439,N_12082,N_13510);
nand U19440 (N_19440,N_11206,N_14373);
xnor U19441 (N_19441,N_14708,N_13732);
nor U19442 (N_19442,N_14945,N_13776);
and U19443 (N_19443,N_14699,N_11778);
or U19444 (N_19444,N_13144,N_14002);
or U19445 (N_19445,N_10497,N_11028);
xnor U19446 (N_19446,N_12290,N_10174);
nand U19447 (N_19447,N_12080,N_14620);
nand U19448 (N_19448,N_11226,N_14793);
nor U19449 (N_19449,N_14818,N_14853);
or U19450 (N_19450,N_13103,N_11289);
or U19451 (N_19451,N_13195,N_12487);
or U19452 (N_19452,N_10017,N_13234);
or U19453 (N_19453,N_10639,N_12393);
and U19454 (N_19454,N_10218,N_13681);
nand U19455 (N_19455,N_10433,N_12900);
nor U19456 (N_19456,N_13172,N_10015);
nor U19457 (N_19457,N_13877,N_13759);
or U19458 (N_19458,N_13630,N_14907);
or U19459 (N_19459,N_14908,N_11907);
nand U19460 (N_19460,N_10084,N_10827);
nor U19461 (N_19461,N_14596,N_13314);
nor U19462 (N_19462,N_11658,N_11466);
nand U19463 (N_19463,N_10289,N_11915);
nor U19464 (N_19464,N_11403,N_14313);
nand U19465 (N_19465,N_14606,N_11595);
nor U19466 (N_19466,N_11165,N_12217);
and U19467 (N_19467,N_13321,N_13773);
xnor U19468 (N_19468,N_13891,N_11251);
and U19469 (N_19469,N_13352,N_10061);
or U19470 (N_19470,N_12675,N_13457);
nand U19471 (N_19471,N_11853,N_12512);
or U19472 (N_19472,N_13505,N_14630);
nor U19473 (N_19473,N_10898,N_11644);
or U19474 (N_19474,N_13392,N_10579);
and U19475 (N_19475,N_13800,N_14408);
and U19476 (N_19476,N_14227,N_14409);
nand U19477 (N_19477,N_14182,N_14647);
and U19478 (N_19478,N_12917,N_13511);
nor U19479 (N_19479,N_10509,N_13328);
and U19480 (N_19480,N_14919,N_14336);
or U19481 (N_19481,N_10320,N_12403);
nor U19482 (N_19482,N_13028,N_13008);
nor U19483 (N_19483,N_11574,N_13727);
nand U19484 (N_19484,N_10944,N_11174);
nor U19485 (N_19485,N_12292,N_12066);
or U19486 (N_19486,N_10603,N_13390);
nor U19487 (N_19487,N_11416,N_14640);
nor U19488 (N_19488,N_12177,N_14211);
nand U19489 (N_19489,N_13065,N_14320);
or U19490 (N_19490,N_11952,N_11453);
or U19491 (N_19491,N_14006,N_10166);
xor U19492 (N_19492,N_14586,N_10888);
or U19493 (N_19493,N_14219,N_12852);
nor U19494 (N_19494,N_12780,N_11955);
nand U19495 (N_19495,N_11395,N_10500);
and U19496 (N_19496,N_10107,N_13816);
or U19497 (N_19497,N_11028,N_10443);
or U19498 (N_19498,N_14498,N_12401);
nor U19499 (N_19499,N_14731,N_13963);
nor U19500 (N_19500,N_11402,N_10389);
or U19501 (N_19501,N_12821,N_13690);
xor U19502 (N_19502,N_14712,N_10182);
xnor U19503 (N_19503,N_10060,N_13700);
xor U19504 (N_19504,N_12651,N_11493);
nand U19505 (N_19505,N_12423,N_10717);
nand U19506 (N_19506,N_11212,N_13613);
nor U19507 (N_19507,N_11364,N_13712);
nor U19508 (N_19508,N_10904,N_12171);
or U19509 (N_19509,N_14143,N_10546);
xor U19510 (N_19510,N_13477,N_10148);
nand U19511 (N_19511,N_11750,N_10902);
xnor U19512 (N_19512,N_10498,N_14415);
nor U19513 (N_19513,N_10700,N_12596);
xnor U19514 (N_19514,N_13476,N_12493);
or U19515 (N_19515,N_14477,N_14735);
nor U19516 (N_19516,N_10358,N_12939);
nand U19517 (N_19517,N_10243,N_14981);
and U19518 (N_19518,N_10055,N_11944);
xor U19519 (N_19519,N_13206,N_11698);
and U19520 (N_19520,N_11251,N_14609);
xnor U19521 (N_19521,N_14186,N_10192);
nand U19522 (N_19522,N_11198,N_13551);
nand U19523 (N_19523,N_14008,N_13558);
or U19524 (N_19524,N_10579,N_12903);
nand U19525 (N_19525,N_12374,N_12856);
and U19526 (N_19526,N_12455,N_10606);
nor U19527 (N_19527,N_14049,N_11707);
nand U19528 (N_19528,N_10831,N_12970);
nor U19529 (N_19529,N_11552,N_13783);
or U19530 (N_19530,N_10025,N_11260);
xor U19531 (N_19531,N_12321,N_11598);
nor U19532 (N_19532,N_11740,N_12637);
nand U19533 (N_19533,N_14240,N_13119);
and U19534 (N_19534,N_11071,N_12580);
or U19535 (N_19535,N_11364,N_12582);
xnor U19536 (N_19536,N_12757,N_10385);
nor U19537 (N_19537,N_12268,N_13515);
nor U19538 (N_19538,N_13462,N_12650);
xor U19539 (N_19539,N_14309,N_10505);
nand U19540 (N_19540,N_10568,N_14437);
and U19541 (N_19541,N_11762,N_13979);
xnor U19542 (N_19542,N_14131,N_12589);
or U19543 (N_19543,N_14536,N_14622);
nor U19544 (N_19544,N_11090,N_13437);
nor U19545 (N_19545,N_13089,N_14145);
nand U19546 (N_19546,N_13313,N_10365);
nand U19547 (N_19547,N_12563,N_11033);
xor U19548 (N_19548,N_13945,N_14649);
nor U19549 (N_19549,N_13344,N_10974);
xnor U19550 (N_19550,N_10646,N_13941);
xnor U19551 (N_19551,N_10442,N_14804);
nor U19552 (N_19552,N_13082,N_10915);
nor U19553 (N_19553,N_12551,N_12445);
xnor U19554 (N_19554,N_13097,N_10903);
nand U19555 (N_19555,N_13477,N_11534);
and U19556 (N_19556,N_11846,N_13265);
and U19557 (N_19557,N_11321,N_12090);
nor U19558 (N_19558,N_10227,N_11913);
nor U19559 (N_19559,N_12605,N_14578);
nand U19560 (N_19560,N_13393,N_10594);
and U19561 (N_19561,N_13279,N_12851);
nand U19562 (N_19562,N_12040,N_12849);
xor U19563 (N_19563,N_10250,N_11951);
or U19564 (N_19564,N_11735,N_14670);
nand U19565 (N_19565,N_13163,N_10933);
nand U19566 (N_19566,N_10692,N_12408);
or U19567 (N_19567,N_10312,N_14205);
nand U19568 (N_19568,N_13243,N_11329);
xnor U19569 (N_19569,N_14393,N_13777);
nand U19570 (N_19570,N_10203,N_13015);
and U19571 (N_19571,N_14351,N_11008);
nor U19572 (N_19572,N_14185,N_10147);
nor U19573 (N_19573,N_10592,N_11988);
and U19574 (N_19574,N_10664,N_10499);
xnor U19575 (N_19575,N_11342,N_11409);
or U19576 (N_19576,N_12521,N_10575);
nor U19577 (N_19577,N_14668,N_10797);
xor U19578 (N_19578,N_12967,N_12535);
xnor U19579 (N_19579,N_14095,N_11776);
xnor U19580 (N_19580,N_10049,N_10632);
or U19581 (N_19581,N_12337,N_12564);
and U19582 (N_19582,N_11017,N_11846);
nor U19583 (N_19583,N_12228,N_11750);
or U19584 (N_19584,N_13859,N_14347);
and U19585 (N_19585,N_11824,N_12971);
nor U19586 (N_19586,N_10601,N_14658);
nor U19587 (N_19587,N_11972,N_12712);
xnor U19588 (N_19588,N_13750,N_11048);
nor U19589 (N_19589,N_10465,N_10684);
nand U19590 (N_19590,N_11687,N_10649);
nor U19591 (N_19591,N_14677,N_13013);
nand U19592 (N_19592,N_14445,N_12802);
and U19593 (N_19593,N_12784,N_11352);
or U19594 (N_19594,N_12571,N_11024);
and U19595 (N_19595,N_11556,N_11053);
and U19596 (N_19596,N_13922,N_14208);
or U19597 (N_19597,N_14949,N_14257);
xor U19598 (N_19598,N_13868,N_12926);
xor U19599 (N_19599,N_14866,N_11370);
nor U19600 (N_19600,N_10804,N_11391);
xnor U19601 (N_19601,N_14511,N_10777);
nor U19602 (N_19602,N_11257,N_13503);
and U19603 (N_19603,N_10835,N_12297);
nor U19604 (N_19604,N_10416,N_11315);
nor U19605 (N_19605,N_13685,N_13112);
nand U19606 (N_19606,N_14855,N_11416);
or U19607 (N_19607,N_10498,N_11516);
and U19608 (N_19608,N_10254,N_14290);
nand U19609 (N_19609,N_11159,N_11930);
and U19610 (N_19610,N_10429,N_12764);
xor U19611 (N_19611,N_12346,N_11907);
nor U19612 (N_19612,N_10375,N_13120);
xor U19613 (N_19613,N_10585,N_12398);
nand U19614 (N_19614,N_14502,N_14566);
nand U19615 (N_19615,N_12315,N_14307);
nand U19616 (N_19616,N_10623,N_11649);
nand U19617 (N_19617,N_14052,N_10513);
nand U19618 (N_19618,N_13347,N_12522);
nor U19619 (N_19619,N_10130,N_11037);
and U19620 (N_19620,N_11418,N_12148);
and U19621 (N_19621,N_11088,N_12707);
nor U19622 (N_19622,N_11419,N_12038);
nor U19623 (N_19623,N_11218,N_11312);
or U19624 (N_19624,N_12382,N_11297);
or U19625 (N_19625,N_13288,N_12737);
or U19626 (N_19626,N_10495,N_14398);
nor U19627 (N_19627,N_11687,N_14418);
or U19628 (N_19628,N_11291,N_10831);
or U19629 (N_19629,N_12641,N_10195);
xor U19630 (N_19630,N_11183,N_11859);
nor U19631 (N_19631,N_14240,N_10965);
nor U19632 (N_19632,N_12335,N_10338);
nor U19633 (N_19633,N_11611,N_13742);
and U19634 (N_19634,N_14775,N_11239);
nor U19635 (N_19635,N_14426,N_13784);
nand U19636 (N_19636,N_11125,N_10440);
and U19637 (N_19637,N_12312,N_12311);
xnor U19638 (N_19638,N_12622,N_10605);
nand U19639 (N_19639,N_11890,N_11090);
nand U19640 (N_19640,N_10226,N_11895);
or U19641 (N_19641,N_13201,N_10121);
nor U19642 (N_19642,N_10568,N_11657);
nand U19643 (N_19643,N_10591,N_14174);
nor U19644 (N_19644,N_11555,N_13101);
and U19645 (N_19645,N_13314,N_13640);
or U19646 (N_19646,N_10646,N_11461);
and U19647 (N_19647,N_14973,N_13815);
nand U19648 (N_19648,N_13025,N_13341);
nand U19649 (N_19649,N_10522,N_10488);
and U19650 (N_19650,N_14351,N_13343);
nand U19651 (N_19651,N_14583,N_11999);
or U19652 (N_19652,N_12739,N_13739);
or U19653 (N_19653,N_14844,N_14916);
nor U19654 (N_19654,N_11680,N_14837);
nor U19655 (N_19655,N_13292,N_11181);
and U19656 (N_19656,N_13963,N_14989);
and U19657 (N_19657,N_11914,N_10330);
nand U19658 (N_19658,N_13489,N_11324);
or U19659 (N_19659,N_11700,N_14472);
nand U19660 (N_19660,N_11056,N_14617);
nor U19661 (N_19661,N_11052,N_10514);
xnor U19662 (N_19662,N_14406,N_11017);
nor U19663 (N_19663,N_12325,N_14216);
nand U19664 (N_19664,N_14571,N_10933);
nor U19665 (N_19665,N_14022,N_10462);
or U19666 (N_19666,N_12872,N_12841);
or U19667 (N_19667,N_11844,N_12458);
and U19668 (N_19668,N_13780,N_10437);
and U19669 (N_19669,N_14495,N_12725);
nand U19670 (N_19670,N_12414,N_11415);
nor U19671 (N_19671,N_10633,N_10906);
xor U19672 (N_19672,N_12175,N_12014);
nand U19673 (N_19673,N_14861,N_11068);
nor U19674 (N_19674,N_12596,N_13012);
nor U19675 (N_19675,N_13364,N_13681);
nor U19676 (N_19676,N_11406,N_13555);
nor U19677 (N_19677,N_14339,N_13246);
and U19678 (N_19678,N_12188,N_14109);
or U19679 (N_19679,N_13864,N_11973);
xnor U19680 (N_19680,N_10930,N_11670);
and U19681 (N_19681,N_11506,N_14204);
nand U19682 (N_19682,N_13323,N_13546);
and U19683 (N_19683,N_13705,N_11837);
xnor U19684 (N_19684,N_14791,N_10493);
or U19685 (N_19685,N_13404,N_11049);
xnor U19686 (N_19686,N_14822,N_11891);
nor U19687 (N_19687,N_12886,N_13590);
or U19688 (N_19688,N_11464,N_14741);
nand U19689 (N_19689,N_14183,N_13566);
xnor U19690 (N_19690,N_14685,N_14210);
xnor U19691 (N_19691,N_10734,N_14076);
xor U19692 (N_19692,N_12884,N_11394);
xnor U19693 (N_19693,N_10867,N_12955);
xor U19694 (N_19694,N_14211,N_12272);
nand U19695 (N_19695,N_12566,N_12476);
nand U19696 (N_19696,N_10971,N_10666);
xor U19697 (N_19697,N_10324,N_12893);
and U19698 (N_19698,N_11254,N_14168);
and U19699 (N_19699,N_13885,N_13813);
and U19700 (N_19700,N_14399,N_14224);
nand U19701 (N_19701,N_11332,N_14243);
or U19702 (N_19702,N_12010,N_12429);
xor U19703 (N_19703,N_14045,N_13966);
nand U19704 (N_19704,N_11594,N_14165);
xor U19705 (N_19705,N_10507,N_14694);
xor U19706 (N_19706,N_13682,N_14323);
and U19707 (N_19707,N_10983,N_11307);
or U19708 (N_19708,N_13802,N_13172);
nor U19709 (N_19709,N_11283,N_10044);
nand U19710 (N_19710,N_14533,N_14596);
and U19711 (N_19711,N_14717,N_14339);
nand U19712 (N_19712,N_14633,N_10013);
nor U19713 (N_19713,N_14556,N_11660);
or U19714 (N_19714,N_10419,N_14284);
and U19715 (N_19715,N_12699,N_11258);
xnor U19716 (N_19716,N_14427,N_13653);
or U19717 (N_19717,N_11254,N_10736);
nor U19718 (N_19718,N_12386,N_11920);
nor U19719 (N_19719,N_10804,N_13888);
nor U19720 (N_19720,N_11677,N_12933);
nor U19721 (N_19721,N_13525,N_12787);
or U19722 (N_19722,N_10774,N_11687);
xor U19723 (N_19723,N_13291,N_12545);
nor U19724 (N_19724,N_12417,N_13434);
nor U19725 (N_19725,N_11617,N_13649);
nor U19726 (N_19726,N_12383,N_10944);
xnor U19727 (N_19727,N_11552,N_11974);
xnor U19728 (N_19728,N_12618,N_11114);
xnor U19729 (N_19729,N_10864,N_10183);
and U19730 (N_19730,N_10753,N_11875);
or U19731 (N_19731,N_12950,N_10632);
nand U19732 (N_19732,N_12765,N_10703);
or U19733 (N_19733,N_14168,N_13409);
nand U19734 (N_19734,N_10008,N_11206);
xnor U19735 (N_19735,N_13003,N_10599);
or U19736 (N_19736,N_12554,N_14979);
nor U19737 (N_19737,N_11628,N_13297);
xor U19738 (N_19738,N_11549,N_11032);
and U19739 (N_19739,N_14228,N_14525);
xor U19740 (N_19740,N_12556,N_10456);
or U19741 (N_19741,N_13461,N_10600);
or U19742 (N_19742,N_13068,N_14603);
and U19743 (N_19743,N_13015,N_12845);
xor U19744 (N_19744,N_12945,N_12616);
xor U19745 (N_19745,N_11305,N_10123);
and U19746 (N_19746,N_11994,N_11436);
or U19747 (N_19747,N_13102,N_12573);
nand U19748 (N_19748,N_10194,N_10286);
xnor U19749 (N_19749,N_11564,N_10721);
nand U19750 (N_19750,N_13027,N_14208);
and U19751 (N_19751,N_11995,N_11052);
and U19752 (N_19752,N_11096,N_14772);
nand U19753 (N_19753,N_14063,N_12109);
or U19754 (N_19754,N_14744,N_13636);
or U19755 (N_19755,N_12437,N_13453);
or U19756 (N_19756,N_13244,N_13355);
nor U19757 (N_19757,N_11848,N_11815);
or U19758 (N_19758,N_10508,N_14193);
or U19759 (N_19759,N_11134,N_11956);
or U19760 (N_19760,N_12638,N_12377);
and U19761 (N_19761,N_12140,N_14418);
and U19762 (N_19762,N_12942,N_14313);
and U19763 (N_19763,N_14874,N_14123);
and U19764 (N_19764,N_12074,N_13595);
and U19765 (N_19765,N_14052,N_14851);
or U19766 (N_19766,N_13430,N_10682);
or U19767 (N_19767,N_14931,N_13684);
nor U19768 (N_19768,N_10960,N_14862);
nor U19769 (N_19769,N_10242,N_11783);
nand U19770 (N_19770,N_10518,N_10377);
or U19771 (N_19771,N_14087,N_11335);
or U19772 (N_19772,N_14285,N_11959);
or U19773 (N_19773,N_13353,N_11118);
nor U19774 (N_19774,N_12063,N_10810);
or U19775 (N_19775,N_10949,N_12144);
nor U19776 (N_19776,N_12250,N_12287);
xor U19777 (N_19777,N_10475,N_10868);
and U19778 (N_19778,N_12492,N_14099);
nor U19779 (N_19779,N_13745,N_10161);
and U19780 (N_19780,N_14137,N_12860);
or U19781 (N_19781,N_11388,N_13764);
nor U19782 (N_19782,N_12247,N_10240);
and U19783 (N_19783,N_11868,N_10530);
or U19784 (N_19784,N_14093,N_11689);
nand U19785 (N_19785,N_13203,N_11347);
or U19786 (N_19786,N_13513,N_11468);
xnor U19787 (N_19787,N_14539,N_13100);
nand U19788 (N_19788,N_11680,N_12080);
nand U19789 (N_19789,N_10935,N_11573);
xnor U19790 (N_19790,N_14603,N_13614);
nand U19791 (N_19791,N_11917,N_12989);
nor U19792 (N_19792,N_10195,N_12807);
xnor U19793 (N_19793,N_13471,N_11726);
nand U19794 (N_19794,N_13086,N_11123);
xnor U19795 (N_19795,N_10676,N_13129);
or U19796 (N_19796,N_12154,N_10507);
nand U19797 (N_19797,N_11328,N_10937);
xor U19798 (N_19798,N_14517,N_14370);
xnor U19799 (N_19799,N_13709,N_11164);
xnor U19800 (N_19800,N_13626,N_12538);
xnor U19801 (N_19801,N_12626,N_14863);
xor U19802 (N_19802,N_10220,N_11541);
nor U19803 (N_19803,N_11862,N_14437);
nor U19804 (N_19804,N_14843,N_14966);
nand U19805 (N_19805,N_11624,N_12292);
xor U19806 (N_19806,N_13531,N_14060);
or U19807 (N_19807,N_13701,N_11373);
xor U19808 (N_19808,N_10264,N_14913);
nand U19809 (N_19809,N_11661,N_10977);
nor U19810 (N_19810,N_10452,N_12092);
xor U19811 (N_19811,N_13965,N_10078);
or U19812 (N_19812,N_12762,N_11964);
nand U19813 (N_19813,N_12194,N_12786);
xnor U19814 (N_19814,N_12498,N_10339);
and U19815 (N_19815,N_10123,N_13191);
nor U19816 (N_19816,N_12734,N_13998);
nand U19817 (N_19817,N_10626,N_10177);
nor U19818 (N_19818,N_13802,N_11992);
xnor U19819 (N_19819,N_10345,N_11844);
nor U19820 (N_19820,N_13871,N_10928);
xor U19821 (N_19821,N_12927,N_10247);
nor U19822 (N_19822,N_13815,N_10195);
and U19823 (N_19823,N_10465,N_12712);
and U19824 (N_19824,N_10808,N_13885);
nor U19825 (N_19825,N_14400,N_10363);
xnor U19826 (N_19826,N_13786,N_12451);
xor U19827 (N_19827,N_12739,N_10059);
xor U19828 (N_19828,N_14689,N_13406);
nand U19829 (N_19829,N_13230,N_14339);
nand U19830 (N_19830,N_14612,N_11227);
and U19831 (N_19831,N_10792,N_13930);
nand U19832 (N_19832,N_14472,N_12089);
nor U19833 (N_19833,N_11365,N_13063);
or U19834 (N_19834,N_14870,N_11716);
xnor U19835 (N_19835,N_10769,N_14490);
nor U19836 (N_19836,N_10699,N_13980);
or U19837 (N_19837,N_10090,N_12627);
or U19838 (N_19838,N_10163,N_11032);
nor U19839 (N_19839,N_10992,N_12910);
xor U19840 (N_19840,N_14776,N_11522);
nor U19841 (N_19841,N_11572,N_14222);
or U19842 (N_19842,N_13639,N_14570);
nand U19843 (N_19843,N_13412,N_10636);
xnor U19844 (N_19844,N_13936,N_12511);
nand U19845 (N_19845,N_11317,N_11448);
and U19846 (N_19846,N_11380,N_14990);
xor U19847 (N_19847,N_13834,N_10367);
xnor U19848 (N_19848,N_11404,N_13896);
nand U19849 (N_19849,N_11898,N_10254);
xor U19850 (N_19850,N_11339,N_11244);
nand U19851 (N_19851,N_12077,N_12099);
nand U19852 (N_19852,N_11991,N_12140);
and U19853 (N_19853,N_14600,N_10501);
xnor U19854 (N_19854,N_14235,N_12039);
and U19855 (N_19855,N_12365,N_10914);
or U19856 (N_19856,N_14138,N_13405);
nor U19857 (N_19857,N_14435,N_13384);
or U19858 (N_19858,N_14495,N_10093);
and U19859 (N_19859,N_14751,N_14356);
xor U19860 (N_19860,N_12591,N_10147);
nor U19861 (N_19861,N_14558,N_10043);
xnor U19862 (N_19862,N_11754,N_11621);
nor U19863 (N_19863,N_10473,N_12686);
xor U19864 (N_19864,N_11820,N_10534);
and U19865 (N_19865,N_11185,N_11782);
nand U19866 (N_19866,N_12800,N_12096);
nand U19867 (N_19867,N_13559,N_12830);
and U19868 (N_19868,N_14793,N_13616);
nor U19869 (N_19869,N_14943,N_10342);
xnor U19870 (N_19870,N_14952,N_14724);
and U19871 (N_19871,N_13879,N_14709);
or U19872 (N_19872,N_14289,N_10260);
nor U19873 (N_19873,N_14899,N_14955);
and U19874 (N_19874,N_13853,N_12927);
and U19875 (N_19875,N_13505,N_11841);
nand U19876 (N_19876,N_10871,N_12504);
and U19877 (N_19877,N_10933,N_13951);
nor U19878 (N_19878,N_14980,N_10191);
and U19879 (N_19879,N_14730,N_13502);
xnor U19880 (N_19880,N_13768,N_10031);
xnor U19881 (N_19881,N_14857,N_12824);
or U19882 (N_19882,N_13167,N_12747);
nor U19883 (N_19883,N_14045,N_14013);
or U19884 (N_19884,N_11745,N_11548);
or U19885 (N_19885,N_10874,N_10954);
nor U19886 (N_19886,N_14205,N_12030);
and U19887 (N_19887,N_13221,N_12480);
or U19888 (N_19888,N_11218,N_11555);
and U19889 (N_19889,N_11439,N_12920);
or U19890 (N_19890,N_11630,N_14548);
or U19891 (N_19891,N_14886,N_10430);
nor U19892 (N_19892,N_10830,N_13326);
or U19893 (N_19893,N_12294,N_11096);
nand U19894 (N_19894,N_12972,N_13193);
nor U19895 (N_19895,N_14654,N_14150);
or U19896 (N_19896,N_12433,N_14284);
nor U19897 (N_19897,N_12866,N_11496);
xnor U19898 (N_19898,N_13519,N_14170);
and U19899 (N_19899,N_11783,N_14964);
nand U19900 (N_19900,N_10078,N_10888);
xnor U19901 (N_19901,N_10064,N_12199);
nor U19902 (N_19902,N_12449,N_10627);
or U19903 (N_19903,N_12399,N_12539);
or U19904 (N_19904,N_10119,N_12106);
xor U19905 (N_19905,N_11285,N_14272);
nor U19906 (N_19906,N_12150,N_14424);
nor U19907 (N_19907,N_10561,N_14560);
nor U19908 (N_19908,N_11517,N_11318);
and U19909 (N_19909,N_11280,N_14458);
nor U19910 (N_19910,N_14206,N_14874);
and U19911 (N_19911,N_10900,N_12951);
nor U19912 (N_19912,N_12872,N_13101);
or U19913 (N_19913,N_10578,N_10122);
xor U19914 (N_19914,N_14562,N_13076);
xor U19915 (N_19915,N_13171,N_11879);
and U19916 (N_19916,N_13104,N_14787);
nor U19917 (N_19917,N_12208,N_12335);
and U19918 (N_19918,N_10923,N_10471);
nor U19919 (N_19919,N_14501,N_10814);
xnor U19920 (N_19920,N_10986,N_11371);
nand U19921 (N_19921,N_11858,N_14312);
xor U19922 (N_19922,N_13152,N_13535);
and U19923 (N_19923,N_12479,N_14192);
nor U19924 (N_19924,N_11210,N_11186);
nand U19925 (N_19925,N_13432,N_11015);
and U19926 (N_19926,N_12114,N_11943);
xnor U19927 (N_19927,N_12293,N_14196);
nand U19928 (N_19928,N_12220,N_10041);
and U19929 (N_19929,N_12975,N_12870);
nand U19930 (N_19930,N_10600,N_11430);
or U19931 (N_19931,N_14858,N_12631);
nand U19932 (N_19932,N_14533,N_10191);
xor U19933 (N_19933,N_13080,N_14737);
and U19934 (N_19934,N_10626,N_12524);
nor U19935 (N_19935,N_13323,N_13496);
and U19936 (N_19936,N_13461,N_13027);
xor U19937 (N_19937,N_12829,N_13803);
nor U19938 (N_19938,N_12687,N_11010);
xor U19939 (N_19939,N_13829,N_12695);
or U19940 (N_19940,N_13997,N_14387);
or U19941 (N_19941,N_11125,N_12199);
or U19942 (N_19942,N_10240,N_10328);
nor U19943 (N_19943,N_14571,N_12483);
or U19944 (N_19944,N_14479,N_12327);
nand U19945 (N_19945,N_14790,N_12542);
xnor U19946 (N_19946,N_12987,N_10857);
nand U19947 (N_19947,N_14727,N_10937);
nand U19948 (N_19948,N_12427,N_14062);
and U19949 (N_19949,N_12653,N_13322);
nand U19950 (N_19950,N_11664,N_10982);
and U19951 (N_19951,N_13251,N_12948);
xnor U19952 (N_19952,N_12579,N_10485);
or U19953 (N_19953,N_12412,N_13485);
nor U19954 (N_19954,N_10425,N_13042);
nor U19955 (N_19955,N_10745,N_11710);
nor U19956 (N_19956,N_13702,N_10434);
or U19957 (N_19957,N_13343,N_12043);
nor U19958 (N_19958,N_13625,N_14541);
xnor U19959 (N_19959,N_14747,N_13984);
xor U19960 (N_19960,N_13350,N_12100);
nor U19961 (N_19961,N_12088,N_11776);
or U19962 (N_19962,N_12277,N_10692);
xnor U19963 (N_19963,N_10075,N_10054);
xnor U19964 (N_19964,N_11881,N_12726);
and U19965 (N_19965,N_10918,N_10505);
and U19966 (N_19966,N_12058,N_13362);
and U19967 (N_19967,N_10796,N_11891);
nand U19968 (N_19968,N_11741,N_14962);
or U19969 (N_19969,N_10980,N_14704);
nor U19970 (N_19970,N_12269,N_13605);
nor U19971 (N_19971,N_11799,N_10116);
nor U19972 (N_19972,N_14073,N_10746);
and U19973 (N_19973,N_12375,N_10577);
xnor U19974 (N_19974,N_13449,N_12806);
and U19975 (N_19975,N_12973,N_11943);
nand U19976 (N_19976,N_10450,N_14803);
and U19977 (N_19977,N_12310,N_10396);
nand U19978 (N_19978,N_11900,N_14533);
nand U19979 (N_19979,N_10567,N_12249);
xor U19980 (N_19980,N_11972,N_10977);
xnor U19981 (N_19981,N_10164,N_12405);
and U19982 (N_19982,N_14643,N_11935);
nand U19983 (N_19983,N_14959,N_10381);
or U19984 (N_19984,N_14319,N_13534);
and U19985 (N_19985,N_11196,N_10123);
nand U19986 (N_19986,N_13667,N_13811);
xor U19987 (N_19987,N_13591,N_13863);
and U19988 (N_19988,N_11436,N_14923);
and U19989 (N_19989,N_13095,N_13461);
nor U19990 (N_19990,N_13683,N_11530);
nand U19991 (N_19991,N_11995,N_13439);
nand U19992 (N_19992,N_10866,N_10897);
or U19993 (N_19993,N_12002,N_13092);
xnor U19994 (N_19994,N_13313,N_12343);
xnor U19995 (N_19995,N_10298,N_11578);
xnor U19996 (N_19996,N_13582,N_12551);
nor U19997 (N_19997,N_14188,N_10276);
xor U19998 (N_19998,N_12547,N_11524);
nand U19999 (N_19999,N_12125,N_13575);
and UO_0 (O_0,N_17439,N_16727);
xor UO_1 (O_1,N_15851,N_15391);
nand UO_2 (O_2,N_16456,N_16592);
nand UO_3 (O_3,N_17579,N_15969);
and UO_4 (O_4,N_18833,N_15560);
nor UO_5 (O_5,N_19348,N_16708);
nor UO_6 (O_6,N_16987,N_15842);
nand UO_7 (O_7,N_15399,N_15197);
xnor UO_8 (O_8,N_17879,N_18609);
xnor UO_9 (O_9,N_19434,N_15323);
nor UO_10 (O_10,N_19750,N_16489);
xor UO_11 (O_11,N_17937,N_19586);
or UO_12 (O_12,N_19024,N_18610);
and UO_13 (O_13,N_18840,N_18666);
nor UO_14 (O_14,N_16659,N_17122);
and UO_15 (O_15,N_16466,N_18208);
xnor UO_16 (O_16,N_15302,N_17338);
or UO_17 (O_17,N_18559,N_18126);
nand UO_18 (O_18,N_15108,N_18916);
xnor UO_19 (O_19,N_16684,N_16296);
and UO_20 (O_20,N_15263,N_18365);
nand UO_21 (O_21,N_15376,N_17656);
nor UO_22 (O_22,N_15480,N_16743);
nor UO_23 (O_23,N_17827,N_19698);
or UO_24 (O_24,N_17914,N_17595);
xnor UO_25 (O_25,N_16681,N_17905);
and UO_26 (O_26,N_16918,N_16971);
or UO_27 (O_27,N_16236,N_17723);
xor UO_28 (O_28,N_17095,N_19834);
xnor UO_29 (O_29,N_18817,N_15992);
nor UO_30 (O_30,N_17391,N_18147);
nor UO_31 (O_31,N_18615,N_15821);
xnor UO_32 (O_32,N_19200,N_18520);
and UO_33 (O_33,N_18130,N_15184);
nand UO_34 (O_34,N_19438,N_18663);
or UO_35 (O_35,N_15023,N_17539);
nand UO_36 (O_36,N_16406,N_16945);
and UO_37 (O_37,N_16598,N_17941);
nand UO_38 (O_38,N_15653,N_15609);
nor UO_39 (O_39,N_16650,N_17846);
nand UO_40 (O_40,N_18456,N_15107);
nand UO_41 (O_41,N_16356,N_16087);
and UO_42 (O_42,N_19784,N_17986);
and UO_43 (O_43,N_18503,N_15695);
nand UO_44 (O_44,N_18254,N_18891);
xor UO_45 (O_45,N_17714,N_15975);
nand UO_46 (O_46,N_17239,N_17818);
nor UO_47 (O_47,N_18472,N_17763);
nor UO_48 (O_48,N_17629,N_17868);
nor UO_49 (O_49,N_17284,N_19042);
nor UO_50 (O_50,N_17070,N_17952);
xor UO_51 (O_51,N_17869,N_19849);
nand UO_52 (O_52,N_15146,N_15577);
and UO_53 (O_53,N_17458,N_18748);
and UO_54 (O_54,N_15087,N_17526);
xnor UO_55 (O_55,N_15699,N_17408);
xnor UO_56 (O_56,N_15491,N_17464);
xnor UO_57 (O_57,N_18272,N_17079);
xnor UO_58 (O_58,N_17100,N_18252);
nand UO_59 (O_59,N_15908,N_15034);
xor UO_60 (O_60,N_18718,N_15164);
or UO_61 (O_61,N_15886,N_16639);
nand UO_62 (O_62,N_18979,N_19796);
or UO_63 (O_63,N_15060,N_19667);
nand UO_64 (O_64,N_16979,N_16013);
or UO_65 (O_65,N_19824,N_16313);
or UO_66 (O_66,N_15503,N_18211);
or UO_67 (O_67,N_16404,N_19265);
or UO_68 (O_68,N_16314,N_15589);
nand UO_69 (O_69,N_15642,N_15050);
and UO_70 (O_70,N_16662,N_16306);
xor UO_71 (O_71,N_15183,N_17590);
and UO_72 (O_72,N_18243,N_18440);
and UO_73 (O_73,N_17253,N_18716);
and UO_74 (O_74,N_16323,N_19004);
nand UO_75 (O_75,N_17883,N_17547);
xnor UO_76 (O_76,N_19106,N_19829);
nand UO_77 (O_77,N_16431,N_19765);
xnor UO_78 (O_78,N_18062,N_16744);
or UO_79 (O_79,N_16029,N_18552);
xnor UO_80 (O_80,N_17000,N_16795);
nand UO_81 (O_81,N_16965,N_19813);
xor UO_82 (O_82,N_15047,N_16112);
nor UO_83 (O_83,N_16993,N_17979);
nor UO_84 (O_84,N_18069,N_16173);
xnor UO_85 (O_85,N_19056,N_17775);
nor UO_86 (O_86,N_17616,N_15586);
and UO_87 (O_87,N_19221,N_18002);
and UO_88 (O_88,N_16104,N_15168);
and UO_89 (O_89,N_17807,N_19192);
xor UO_90 (O_90,N_15896,N_19022);
and UO_91 (O_91,N_19055,N_17360);
xnor UO_92 (O_92,N_19939,N_17323);
or UO_93 (O_93,N_15703,N_15418);
or UO_94 (O_94,N_17867,N_18136);
and UO_95 (O_95,N_17913,N_18360);
nor UO_96 (O_96,N_18774,N_18318);
nand UO_97 (O_97,N_15457,N_19462);
or UO_98 (O_98,N_18868,N_18164);
nand UO_99 (O_99,N_19312,N_18006);
nor UO_100 (O_100,N_16585,N_15248);
or UO_101 (O_101,N_17944,N_17811);
nor UO_102 (O_102,N_17535,N_15421);
xnor UO_103 (O_103,N_18512,N_19903);
or UO_104 (O_104,N_19260,N_19583);
nor UO_105 (O_105,N_16887,N_18315);
nand UO_106 (O_106,N_16819,N_18707);
nand UO_107 (O_107,N_18303,N_18181);
nand UO_108 (O_108,N_17374,N_15917);
nand UO_109 (O_109,N_18495,N_17481);
nor UO_110 (O_110,N_19689,N_15620);
or UO_111 (O_111,N_15537,N_15788);
and UO_112 (O_112,N_17097,N_16068);
nand UO_113 (O_113,N_17383,N_16136);
nand UO_114 (O_114,N_17537,N_16920);
and UO_115 (O_115,N_18016,N_17687);
or UO_116 (O_116,N_16687,N_17437);
nand UO_117 (O_117,N_15453,N_15637);
nand UO_118 (O_118,N_18633,N_17243);
xnor UO_119 (O_119,N_17780,N_17131);
and UO_120 (O_120,N_19984,N_19594);
nand UO_121 (O_121,N_19340,N_17828);
nand UO_122 (O_122,N_17705,N_19660);
and UO_123 (O_123,N_16972,N_17959);
and UO_124 (O_124,N_17193,N_16596);
and UO_125 (O_125,N_15603,N_15394);
and UO_126 (O_126,N_16259,N_15354);
nor UO_127 (O_127,N_18038,N_15211);
nor UO_128 (O_128,N_19785,N_15657);
nor UO_129 (O_129,N_15742,N_15199);
or UO_130 (O_130,N_17845,N_16245);
nor UO_131 (O_131,N_18644,N_15329);
nor UO_132 (O_132,N_15527,N_17291);
nand UO_133 (O_133,N_18641,N_19579);
nand UO_134 (O_134,N_17771,N_15835);
xnor UO_135 (O_135,N_16605,N_15624);
and UO_136 (O_136,N_19815,N_15760);
and UO_137 (O_137,N_18330,N_17171);
and UO_138 (O_138,N_18905,N_18008);
nand UO_139 (O_139,N_17228,N_16936);
nor UO_140 (O_140,N_15782,N_17270);
and UO_141 (O_141,N_17303,N_16193);
xor UO_142 (O_142,N_16811,N_17030);
and UO_143 (O_143,N_16672,N_19988);
nor UO_144 (O_144,N_19792,N_16869);
and UO_145 (O_145,N_15535,N_15841);
nand UO_146 (O_146,N_18203,N_15629);
xnor UO_147 (O_147,N_19492,N_18811);
and UO_148 (O_148,N_19751,N_16165);
xor UO_149 (O_149,N_18753,N_16902);
or UO_150 (O_150,N_19968,N_18441);
and UO_151 (O_151,N_18986,N_17322);
nand UO_152 (O_152,N_16262,N_17394);
xor UO_153 (O_153,N_18083,N_19344);
nand UO_154 (O_154,N_15683,N_18651);
or UO_155 (O_155,N_18776,N_17466);
nor UO_156 (O_156,N_17511,N_15849);
or UO_157 (O_157,N_16118,N_18971);
nor UO_158 (O_158,N_17601,N_15334);
xnor UO_159 (O_159,N_15918,N_19054);
xnor UO_160 (O_160,N_19182,N_19880);
nand UO_161 (O_161,N_16086,N_17700);
nor UO_162 (O_162,N_17915,N_15987);
nand UO_163 (O_163,N_19453,N_15346);
and UO_164 (O_164,N_19623,N_18909);
or UO_165 (O_165,N_19333,N_17278);
and UO_166 (O_166,N_16837,N_15820);
and UO_167 (O_167,N_16721,N_19725);
nor UO_168 (O_168,N_15832,N_19907);
nand UO_169 (O_169,N_18406,N_17636);
nand UO_170 (O_170,N_16571,N_19266);
or UO_171 (O_171,N_17877,N_18127);
xor UO_172 (O_172,N_17974,N_18158);
nand UO_173 (O_173,N_19239,N_16510);
nor UO_174 (O_174,N_17888,N_19954);
and UO_175 (O_175,N_16527,N_18681);
and UO_176 (O_176,N_15651,N_19037);
and UO_177 (O_177,N_17584,N_16617);
or UO_178 (O_178,N_17320,N_17365);
and UO_179 (O_179,N_16186,N_15954);
nand UO_180 (O_180,N_17908,N_16254);
nor UO_181 (O_181,N_15118,N_16564);
or UO_182 (O_182,N_17621,N_19670);
xor UO_183 (O_183,N_16577,N_16771);
or UO_184 (O_184,N_16606,N_16781);
nor UO_185 (O_185,N_17088,N_16647);
xnor UO_186 (O_186,N_16940,N_16707);
or UO_187 (O_187,N_17376,N_17693);
and UO_188 (O_188,N_18457,N_15831);
and UO_189 (O_189,N_17151,N_15481);
nor UO_190 (O_190,N_16853,N_17615);
xor UO_191 (O_191,N_19145,N_16656);
and UO_192 (O_192,N_16303,N_16109);
xnor UO_193 (O_193,N_19040,N_16238);
nor UO_194 (O_194,N_16559,N_16786);
or UO_195 (O_195,N_16504,N_15972);
xor UO_196 (O_196,N_16753,N_16115);
or UO_197 (O_197,N_16586,N_19257);
or UO_198 (O_198,N_19140,N_19914);
nand UO_199 (O_199,N_19994,N_15644);
nand UO_200 (O_200,N_17533,N_17810);
xnor UO_201 (O_201,N_19119,N_16439);
and UO_202 (O_202,N_15521,N_16052);
xnor UO_203 (O_203,N_18572,N_18411);
nand UO_204 (O_204,N_16507,N_15648);
nor UO_205 (O_205,N_16151,N_15003);
and UO_206 (O_206,N_18936,N_17544);
and UO_207 (O_207,N_16692,N_18383);
xnor UO_208 (O_208,N_15966,N_16712);
or UO_209 (O_209,N_19541,N_17377);
and UO_210 (O_210,N_17143,N_15486);
nor UO_211 (O_211,N_16745,N_16310);
or UO_212 (O_212,N_19771,N_19190);
xnor UO_213 (O_213,N_18198,N_18858);
nor UO_214 (O_214,N_18860,N_19697);
nand UO_215 (O_215,N_15568,N_19301);
nand UO_216 (O_216,N_19857,N_19514);
or UO_217 (O_217,N_15317,N_16098);
and UO_218 (O_218,N_19878,N_16409);
nor UO_219 (O_219,N_15132,N_17738);
xor UO_220 (O_220,N_15887,N_18570);
xnor UO_221 (O_221,N_16523,N_16694);
nor UO_222 (O_222,N_19000,N_15476);
and UO_223 (O_223,N_17611,N_18483);
nand UO_224 (O_224,N_17205,N_18799);
nor UO_225 (O_225,N_16216,N_16007);
xor UO_226 (O_226,N_15024,N_18628);
nand UO_227 (O_227,N_15726,N_16642);
and UO_228 (O_228,N_16123,N_16248);
xor UO_229 (O_229,N_16363,N_16604);
and UO_230 (O_230,N_18638,N_15358);
and UO_231 (O_231,N_18820,N_16061);
xnor UO_232 (O_232,N_16355,N_19683);
or UO_233 (O_233,N_16195,N_17178);
xor UO_234 (O_234,N_19261,N_16509);
nor UO_235 (O_235,N_15951,N_16572);
xor UO_236 (O_236,N_19322,N_15335);
or UO_237 (O_237,N_17475,N_16106);
nor UO_238 (O_238,N_17163,N_17002);
nor UO_239 (O_239,N_16437,N_17059);
nor UO_240 (O_240,N_17972,N_15069);
nor UO_241 (O_241,N_17459,N_18058);
nand UO_242 (O_242,N_18773,N_19881);
or UO_243 (O_243,N_18373,N_18851);
or UO_244 (O_244,N_16565,N_15479);
xnor UO_245 (O_245,N_18113,N_19235);
nor UO_246 (O_246,N_17823,N_18410);
or UO_247 (O_247,N_18169,N_16501);
nand UO_248 (O_248,N_19736,N_16562);
and UO_249 (O_249,N_15282,N_18747);
xor UO_250 (O_250,N_16122,N_19155);
and UO_251 (O_251,N_17436,N_17482);
nand UO_252 (O_252,N_16963,N_18005);
nand UO_253 (O_253,N_17499,N_17689);
and UO_254 (O_254,N_17352,N_19110);
xnor UO_255 (O_255,N_17474,N_16796);
xor UO_256 (O_256,N_17919,N_16638);
and UO_257 (O_257,N_17119,N_16344);
nor UO_258 (O_258,N_17203,N_18845);
nand UO_259 (O_259,N_15412,N_16171);
nand UO_260 (O_260,N_19194,N_19211);
nand UO_261 (O_261,N_16986,N_19326);
nand UO_262 (O_262,N_17370,N_16590);
nor UO_263 (O_263,N_19028,N_18217);
xnor UO_264 (O_264,N_16872,N_17757);
nand UO_265 (O_265,N_17060,N_17123);
nor UO_266 (O_266,N_18742,N_19280);
and UO_267 (O_267,N_16257,N_16066);
xor UO_268 (O_268,N_18645,N_15297);
xor UO_269 (O_269,N_16010,N_16557);
and UO_270 (O_270,N_18975,N_19089);
xor UO_271 (O_271,N_15121,N_16839);
and UO_272 (O_272,N_15371,N_15794);
and UO_273 (O_273,N_15370,N_18786);
or UO_274 (O_274,N_17234,N_19294);
nor UO_275 (O_275,N_15165,N_17053);
or UO_276 (O_276,N_17754,N_17036);
xor UO_277 (O_277,N_18515,N_17973);
and UO_278 (O_278,N_17640,N_15551);
and UO_279 (O_279,N_15676,N_18830);
nand UO_280 (O_280,N_15492,N_18731);
and UO_281 (O_281,N_19847,N_18004);
nor UO_282 (O_282,N_16239,N_16922);
and UO_283 (O_283,N_15454,N_17819);
and UO_284 (O_284,N_16612,N_18070);
xnor UO_285 (O_285,N_16824,N_17028);
or UO_286 (O_286,N_16543,N_16567);
nand UO_287 (O_287,N_18746,N_15174);
and UO_288 (O_288,N_15380,N_16256);
xnor UO_289 (O_289,N_15538,N_17166);
and UO_290 (O_290,N_19252,N_16121);
nor UO_291 (O_291,N_15905,N_17411);
or UO_292 (O_292,N_16031,N_16568);
or UO_293 (O_293,N_16822,N_17730);
and UO_294 (O_294,N_16932,N_18403);
nor UO_295 (O_295,N_15331,N_15743);
and UO_296 (O_296,N_16401,N_15257);
and UO_297 (O_297,N_19786,N_19485);
xnor UO_298 (O_298,N_19700,N_18962);
nand UO_299 (O_299,N_18536,N_16646);
nor UO_300 (O_300,N_17460,N_18894);
or UO_301 (O_301,N_16584,N_16937);
xor UO_302 (O_302,N_18598,N_18930);
nor UO_303 (O_303,N_16032,N_17485);
and UO_304 (O_304,N_18863,N_19940);
or UO_305 (O_305,N_16263,N_15242);
xor UO_306 (O_306,N_15460,N_16370);
or UO_307 (O_307,N_17855,N_19398);
nand UO_308 (O_308,N_18445,N_16299);
xor UO_309 (O_309,N_15919,N_18375);
nor UO_310 (O_310,N_15715,N_19549);
nor UO_311 (O_311,N_18513,N_19998);
or UO_312 (O_312,N_19659,N_18701);
or UO_313 (O_313,N_17412,N_19086);
nand UO_314 (O_314,N_16172,N_18745);
xor UO_315 (O_315,N_17951,N_15433);
nand UO_316 (O_316,N_18104,N_15408);
or UO_317 (O_317,N_18730,N_19428);
nor UO_318 (O_318,N_16907,N_15301);
nand UO_319 (O_319,N_16283,N_15103);
xor UO_320 (O_320,N_18761,N_17495);
nor UO_321 (O_321,N_19618,N_18394);
or UO_322 (O_322,N_15296,N_19402);
or UO_323 (O_323,N_15536,N_16196);
nor UO_324 (O_324,N_16761,N_19937);
or UO_325 (O_325,N_17026,N_15946);
xnor UO_326 (O_326,N_16482,N_18199);
xnor UO_327 (O_327,N_18221,N_16494);
or UO_328 (O_328,N_16410,N_15645);
and UO_329 (O_329,N_16374,N_15670);
nor UO_330 (O_330,N_19656,N_16497);
nor UO_331 (O_331,N_17442,N_19757);
nor UO_332 (O_332,N_19682,N_16889);
or UO_333 (O_333,N_19916,N_19507);
nor UO_334 (O_334,N_19922,N_16290);
xnor UO_335 (O_335,N_15030,N_17562);
nand UO_336 (O_336,N_18084,N_19488);
nand UO_337 (O_337,N_15084,N_18150);
nand UO_338 (O_338,N_16422,N_15096);
nor UO_339 (O_339,N_15617,N_16487);
and UO_340 (O_340,N_15855,N_15294);
nand UO_341 (O_341,N_16664,N_16170);
nand UO_342 (O_342,N_15104,N_17204);
nand UO_343 (O_343,N_17786,N_15449);
or UO_344 (O_344,N_16884,N_18956);
or UO_345 (O_345,N_19639,N_16524);
nor UO_346 (O_346,N_17066,N_19853);
xnor UO_347 (O_347,N_18308,N_16957);
and UO_348 (O_348,N_19566,N_17638);
and UO_349 (O_349,N_15866,N_16520);
nor UO_350 (O_350,N_18591,N_18289);
nand UO_351 (O_351,N_18056,N_17334);
or UO_352 (O_352,N_19619,N_16322);
or UO_353 (O_353,N_16483,N_16446);
nand UO_354 (O_354,N_18251,N_18990);
or UO_355 (O_355,N_18093,N_18319);
nor UO_356 (O_356,N_16676,N_19473);
and UO_357 (O_357,N_15100,N_15220);
and UO_358 (O_358,N_18655,N_15076);
or UO_359 (O_359,N_19888,N_17633);
xor UO_360 (O_360,N_15126,N_15193);
nor UO_361 (O_361,N_19482,N_15834);
and UO_362 (O_362,N_17130,N_17190);
nand UO_363 (O_363,N_15732,N_17565);
nand UO_364 (O_364,N_18808,N_17753);
or UO_365 (O_365,N_15665,N_16769);
nor UO_366 (O_366,N_17713,N_19097);
nor UO_367 (O_367,N_15816,N_17658);
xnor UO_368 (O_368,N_16198,N_18565);
or UO_369 (O_369,N_17364,N_17512);
nand UO_370 (O_370,N_15779,N_18311);
xor UO_371 (O_371,N_15347,N_16113);
nand UO_372 (O_372,N_17309,N_17349);
nor UO_373 (O_373,N_18557,N_16677);
nand UO_374 (O_374,N_18895,N_17024);
nand UO_375 (O_375,N_15562,N_16070);
or UO_376 (O_376,N_17453,N_19490);
xnor UO_377 (O_377,N_16127,N_16030);
nor UO_378 (O_378,N_17822,N_15770);
and UO_379 (O_379,N_16009,N_16209);
nor UO_380 (O_380,N_16633,N_19727);
nand UO_381 (O_381,N_17039,N_16375);
xnor UO_382 (O_382,N_19175,N_15110);
nor UO_383 (O_383,N_15028,N_15571);
nor UO_384 (O_384,N_19944,N_18727);
nand UO_385 (O_385,N_17671,N_18577);
and UO_386 (O_386,N_17206,N_17357);
and UO_387 (O_387,N_17379,N_18316);
xor UO_388 (O_388,N_18902,N_19993);
or UO_389 (O_389,N_16108,N_19892);
nor UO_390 (O_390,N_18756,N_17058);
or UO_391 (O_391,N_15662,N_18949);
and UO_392 (O_392,N_18053,N_18549);
xnor UO_393 (O_393,N_17864,N_17675);
nand UO_394 (O_394,N_19752,N_16991);
nor UO_395 (O_395,N_15725,N_16832);
xnor UO_396 (O_396,N_17704,N_15148);
and UO_397 (O_397,N_15952,N_18458);
or UO_398 (O_398,N_18506,N_17113);
and UO_399 (O_399,N_19666,N_19645);
xnor UO_400 (O_400,N_15585,N_19422);
xnor UO_401 (O_401,N_15417,N_19804);
and UO_402 (O_402,N_15077,N_18992);
xnor UO_403 (O_403,N_18751,N_15352);
and UO_404 (O_404,N_19191,N_15434);
nand UO_405 (O_405,N_15928,N_16411);
nor UO_406 (O_406,N_15752,N_16640);
nand UO_407 (O_407,N_17273,N_16843);
xnor UO_408 (O_408,N_17676,N_18976);
nor UO_409 (O_409,N_18369,N_18706);
xor UO_410 (O_410,N_15507,N_19258);
and UO_411 (O_411,N_17701,N_15160);
and UO_412 (O_412,N_17965,N_16615);
xor UO_413 (O_413,N_16159,N_18029);
or UO_414 (O_414,N_15403,N_17970);
xnor UO_415 (O_415,N_16829,N_19608);
nor UO_416 (O_416,N_18602,N_17985);
nand UO_417 (O_417,N_16966,N_16451);
and UO_418 (O_418,N_19284,N_19927);
nand UO_419 (O_419,N_16773,N_16124);
or UO_420 (O_420,N_17497,N_15128);
and UO_421 (O_421,N_18357,N_16386);
or UO_422 (O_422,N_18259,N_15280);
and UO_423 (O_423,N_16474,N_18623);
nor UO_424 (O_424,N_18561,N_19864);
nand UO_425 (O_425,N_16454,N_17553);
nor UO_426 (O_426,N_18744,N_19179);
nor UO_427 (O_427,N_17312,N_18447);
xnor UO_428 (O_428,N_15123,N_19377);
nor UO_429 (O_429,N_16412,N_19909);
nand UO_430 (O_430,N_15031,N_15012);
and UO_431 (O_431,N_15221,N_18166);
xor UO_432 (O_432,N_15252,N_15543);
or UO_433 (O_433,N_16138,N_18195);
and UO_434 (O_434,N_16490,N_16861);
nor UO_435 (O_435,N_15278,N_18214);
nand UO_436 (O_436,N_18819,N_15540);
nand UO_437 (O_437,N_18111,N_19545);
xnor UO_438 (O_438,N_17441,N_16449);
nor UO_439 (O_439,N_16189,N_19099);
xor UO_440 (O_440,N_15680,N_16886);
and UO_441 (O_441,N_17012,N_18980);
xnor UO_442 (O_442,N_17917,N_19693);
or UO_443 (O_443,N_16854,N_18687);
xor UO_444 (O_444,N_19928,N_19195);
nor UO_445 (O_445,N_18178,N_19768);
nand UO_446 (O_446,N_18914,N_18409);
and UO_447 (O_447,N_18276,N_19256);
or UO_448 (O_448,N_16505,N_17225);
nand UO_449 (O_449,N_16663,N_16613);
nor UO_450 (O_450,N_18209,N_16391);
or UO_451 (O_451,N_16426,N_19297);
nand UO_452 (O_452,N_16111,N_15898);
xnor UO_453 (O_453,N_19064,N_19068);
nand UO_454 (O_454,N_15894,N_19758);
and UO_455 (O_455,N_18290,N_19924);
xor UO_456 (O_456,N_18959,N_15903);
xor UO_457 (O_457,N_18759,N_18911);
xor UO_458 (O_458,N_16128,N_19646);
nand UO_459 (O_459,N_18770,N_19003);
or UO_460 (O_460,N_15267,N_17473);
nor UO_461 (O_461,N_15616,N_15411);
and UO_462 (O_462,N_19711,N_17212);
or UO_463 (O_463,N_16095,N_15923);
nor UO_464 (O_464,N_18291,N_17522);
and UO_465 (O_465,N_15934,N_18385);
or UO_466 (O_466,N_19255,N_17957);
xor UO_467 (O_467,N_16390,N_15111);
or UO_468 (O_468,N_15663,N_19742);
or UO_469 (O_469,N_18446,N_19959);
or UO_470 (O_470,N_15061,N_17355);
xnor UO_471 (O_471,N_18678,N_17644);
nor UO_472 (O_472,N_19368,N_18190);
xor UO_473 (O_473,N_19250,N_19637);
or UO_474 (O_474,N_18977,N_15435);
nand UO_475 (O_475,N_18155,N_15180);
xnor UO_476 (O_476,N_18376,N_15879);
and UO_477 (O_477,N_19894,N_17668);
and UO_478 (O_478,N_18064,N_18815);
nor UO_479 (O_479,N_19862,N_19946);
and UO_480 (O_480,N_17594,N_15496);
xor UO_481 (O_481,N_18342,N_19088);
nor UO_482 (O_482,N_18599,N_18923);
nor UO_483 (O_483,N_15432,N_18258);
xor UO_484 (O_484,N_17410,N_15468);
xnor UO_485 (O_485,N_19811,N_19827);
or UO_486 (O_486,N_17162,N_17592);
or UO_487 (O_487,N_19574,N_19216);
nand UO_488 (O_488,N_17837,N_19593);
nand UO_489 (O_489,N_15225,N_19033);
or UO_490 (O_490,N_19609,N_19884);
nand UO_491 (O_491,N_15630,N_18050);
xor UO_492 (O_492,N_16174,N_15428);
nand UO_493 (O_493,N_17093,N_15385);
or UO_494 (O_494,N_15340,N_19925);
nand UO_495 (O_495,N_16213,N_17816);
nor UO_496 (O_496,N_16955,N_16481);
nor UO_497 (O_497,N_16873,N_19472);
xnor UO_498 (O_498,N_16736,N_18380);
and UO_499 (O_499,N_16661,N_18402);
or UO_500 (O_500,N_16142,N_17479);
and UO_501 (O_501,N_16594,N_15765);
nand UO_502 (O_502,N_17477,N_15861);
nand UO_503 (O_503,N_18304,N_18887);
nand UO_504 (O_504,N_17593,N_19197);
and UO_505 (O_505,N_18202,N_18499);
and UO_506 (O_506,N_15163,N_18110);
or UO_507 (O_507,N_15927,N_17413);
nor UO_508 (O_508,N_16673,N_17733);
nor UO_509 (O_509,N_15819,N_19331);
nand UO_510 (O_510,N_18961,N_15759);
or UO_511 (O_511,N_17796,N_19318);
nor UO_512 (O_512,N_19675,N_15693);
nand UO_513 (O_513,N_17496,N_15505);
and UO_514 (O_514,N_16100,N_16740);
xor UO_515 (O_515,N_15569,N_15544);
xnor UO_516 (O_516,N_15388,N_15504);
xor UO_517 (O_517,N_19912,N_19287);
and UO_518 (O_518,N_18118,N_15169);
or UO_519 (O_519,N_15666,N_15349);
xor UO_520 (O_520,N_19278,N_16397);
or UO_521 (O_521,N_15313,N_16133);
nor UO_522 (O_522,N_18073,N_19231);
nor UO_523 (O_523,N_16017,N_15499);
nor UO_524 (O_524,N_18379,N_19530);
xnor UO_525 (O_525,N_19409,N_16710);
or UO_526 (O_526,N_16418,N_17933);
xnor UO_527 (O_527,N_19264,N_19731);
nand UO_528 (O_528,N_19214,N_18032);
and UO_529 (O_529,N_16758,N_16794);
nor UO_530 (O_530,N_17380,N_19797);
nor UO_531 (O_531,N_19807,N_18043);
and UO_532 (O_532,N_18485,N_18099);
nor UO_533 (O_533,N_18484,N_18648);
or UO_534 (O_534,N_18302,N_19662);
and UO_535 (O_535,N_15845,N_16560);
and UO_536 (O_536,N_17926,N_17878);
or UO_537 (O_537,N_18344,N_17385);
nand UO_538 (O_538,N_18794,N_16608);
nor UO_539 (O_539,N_15705,N_19654);
xor UO_540 (O_540,N_18893,N_17343);
xor UO_541 (O_541,N_15643,N_18771);
nand UO_542 (O_542,N_15902,N_18809);
xor UO_543 (O_543,N_18465,N_18569);
and UO_544 (O_544,N_15520,N_15808);
xor UO_545 (O_545,N_16654,N_19652);
nand UO_546 (O_546,N_15885,N_17238);
nand UO_547 (O_547,N_19778,N_15858);
nor UO_548 (O_548,N_18452,N_15395);
nand UO_549 (O_549,N_17259,N_15539);
nor UO_550 (O_550,N_18014,N_15092);
xor UO_551 (O_551,N_19327,N_18048);
nand UO_552 (O_552,N_18408,N_19962);
nand UO_553 (O_553,N_19369,N_15701);
nor UO_554 (O_554,N_16395,N_16836);
and UO_555 (O_555,N_18821,N_17257);
xor UO_556 (O_556,N_15260,N_19595);
or UO_557 (O_557,N_19446,N_16442);
or UO_558 (O_558,N_18711,N_19874);
and UO_559 (O_559,N_15251,N_16950);
nand UO_560 (O_560,N_18985,N_17174);
nand UO_561 (O_561,N_19406,N_19178);
nor UO_562 (O_562,N_15344,N_18066);
nand UO_563 (O_563,N_18493,N_17141);
xor UO_564 (O_564,N_19904,N_19276);
and UO_565 (O_565,N_19354,N_16243);
and UO_566 (O_566,N_17549,N_18030);
and UO_567 (O_567,N_18240,N_19364);
and UO_568 (O_568,N_17798,N_19607);
nor UO_569 (O_569,N_17314,N_16152);
nand UO_570 (O_570,N_17290,N_17604);
xor UO_571 (O_571,N_16156,N_16139);
or UO_572 (O_572,N_18805,N_18886);
and UO_573 (O_573,N_18608,N_18954);
nor UO_574 (O_574,N_17932,N_15157);
nand UO_575 (O_575,N_15541,N_15565);
nand UO_576 (O_576,N_19226,N_18600);
or UO_577 (O_577,N_17199,N_19684);
nand UO_578 (O_578,N_18896,N_16434);
xor UO_579 (O_579,N_16168,N_19127);
nand UO_580 (O_580,N_17463,N_19734);
nand UO_581 (O_581,N_19374,N_19375);
or UO_582 (O_582,N_18517,N_19578);
xor UO_583 (O_583,N_16665,N_19897);
or UO_584 (O_584,N_18582,N_17324);
nand UO_585 (O_585,N_19615,N_17774);
and UO_586 (O_586,N_19941,N_19568);
and UO_587 (O_587,N_19337,N_18673);
nand UO_588 (O_588,N_19102,N_18688);
xnor UO_589 (O_589,N_18947,N_19043);
and UO_590 (O_590,N_15679,N_19410);
xor UO_591 (O_591,N_15716,N_17369);
and UO_592 (O_592,N_15304,N_18141);
xor UO_593 (O_593,N_18089,N_19069);
nand UO_594 (O_594,N_18906,N_15658);
or UO_595 (O_595,N_17582,N_15307);
nor UO_596 (O_596,N_15054,N_17975);
nor UO_597 (O_597,N_15864,N_17898);
or UO_598 (O_598,N_15423,N_19220);
xnor UO_599 (O_599,N_18667,N_17673);
or UO_600 (O_600,N_16982,N_17637);
nor UO_601 (O_601,N_18574,N_16561);
xor UO_602 (O_602,N_15372,N_17814);
nand UO_603 (O_603,N_19091,N_18948);
and UO_604 (O_604,N_17236,N_17386);
nand UO_605 (O_605,N_17462,N_17895);
nor UO_606 (O_606,N_15497,N_17461);
nor UO_607 (O_607,N_18732,N_19933);
nand UO_608 (O_608,N_18596,N_19180);
nor UO_609 (O_609,N_17783,N_16377);
xor UO_610 (O_610,N_19060,N_16246);
xor UO_611 (O_611,N_15079,N_17403);
xor UO_612 (O_612,N_19712,N_17685);
or UO_613 (O_613,N_19748,N_18684);
nand UO_614 (O_614,N_15450,N_19724);
nor UO_615 (O_615,N_18991,N_18873);
nand UO_616 (O_616,N_19219,N_17202);
or UO_617 (O_617,N_17083,N_16748);
and UO_618 (O_618,N_16316,N_18871);
nand UO_619 (O_619,N_17373,N_16117);
or UO_620 (O_620,N_19644,N_18487);
and UO_621 (O_621,N_19431,N_17622);
nand UO_622 (O_622,N_19334,N_15074);
and UO_623 (O_623,N_16408,N_18931);
and UO_624 (O_624,N_15964,N_15707);
nor UO_625 (O_625,N_16103,N_15974);
or UO_626 (O_626,N_16805,N_15200);
xor UO_627 (O_627,N_17504,N_15098);
xnor UO_628 (O_628,N_19961,N_16441);
and UO_629 (O_629,N_15690,N_15033);
nand UO_630 (O_630,N_17682,N_19224);
xor UO_631 (O_631,N_17308,N_18367);
nor UO_632 (O_632,N_15222,N_16833);
xnor UO_633 (O_633,N_18323,N_15189);
and UO_634 (O_634,N_16402,N_16427);
or UO_635 (O_635,N_19115,N_18844);
nand UO_636 (O_636,N_17498,N_19141);
or UO_637 (O_637,N_16366,N_15817);
nor UO_638 (O_638,N_17766,N_15945);
and UO_639 (O_639,N_19715,N_15558);
or UO_640 (O_640,N_16293,N_17177);
or UO_641 (O_641,N_19048,N_18431);
and UO_642 (O_642,N_19339,N_15002);
nand UO_643 (O_643,N_15375,N_17250);
nand UO_644 (O_644,N_18542,N_17581);
nor UO_645 (O_645,N_18420,N_15612);
xnor UO_646 (O_646,N_19934,N_15192);
nand UO_647 (O_647,N_16720,N_18958);
and UO_648 (O_648,N_19906,N_15382);
xor UO_649 (O_649,N_16201,N_15162);
and UO_650 (O_650,N_16167,N_16840);
nor UO_651 (O_651,N_19467,N_18401);
or UO_652 (O_652,N_17849,N_15800);
xor UO_653 (O_653,N_17984,N_16295);
nand UO_654 (O_654,N_18527,N_18419);
xor UO_655 (O_655,N_17189,N_15379);
and UO_656 (O_656,N_17222,N_19974);
or UO_657 (O_657,N_19215,N_17127);
nand UO_658 (O_658,N_16580,N_18109);
nand UO_659 (O_659,N_16129,N_19762);
nor UO_660 (O_660,N_15212,N_15791);
or UO_661 (O_661,N_17605,N_18065);
or UO_662 (O_662,N_18144,N_16860);
nand UO_663 (O_663,N_18965,N_18077);
or UO_664 (O_664,N_15531,N_15733);
and UO_665 (O_665,N_18614,N_18942);
nand UO_666 (O_666,N_17906,N_17226);
and UO_667 (O_667,N_16946,N_16110);
or UO_668 (O_668,N_19782,N_18097);
xor UO_669 (O_669,N_18966,N_17598);
xnor UO_670 (O_670,N_17105,N_16462);
nand UO_671 (O_671,N_19366,N_18611);
and UO_672 (O_672,N_16141,N_19148);
and UO_673 (O_673,N_18031,N_16277);
or UO_674 (O_674,N_15194,N_16655);
and UO_675 (O_675,N_19965,N_15723);
or UO_676 (O_676,N_16043,N_18295);
nor UO_677 (O_677,N_19302,N_18218);
xnor UO_678 (O_678,N_15724,N_15990);
nand UO_679 (O_679,N_18554,N_17054);
and UO_680 (O_680,N_15055,N_17168);
nor UO_681 (O_681,N_18232,N_18970);
nor UO_682 (O_682,N_15692,N_19249);
and UO_683 (O_683,N_19193,N_15328);
nor UO_684 (O_684,N_15881,N_18355);
xor UO_685 (O_685,N_16757,N_15602);
xnor UO_686 (O_686,N_19576,N_17390);
nor UO_687 (O_687,N_19589,N_17620);
nor UO_688 (O_688,N_18359,N_18296);
nor UO_689 (O_689,N_17118,N_15091);
or UO_690 (O_690,N_17697,N_16146);
or UO_691 (O_691,N_17528,N_16900);
or UO_692 (O_692,N_16683,N_15190);
and UO_693 (O_693,N_17833,N_17524);
and UO_694 (O_694,N_15948,N_16048);
or UO_695 (O_695,N_18424,N_18242);
and UO_696 (O_696,N_18106,N_16522);
or UO_697 (O_697,N_18335,N_16949);
xor UO_698 (O_698,N_15681,N_16845);
nand UO_699 (O_699,N_16219,N_19017);
or UO_700 (O_700,N_17111,N_16336);
xnor UO_701 (O_701,N_18249,N_17527);
nand UO_702 (O_702,N_16200,N_18103);
xor UO_703 (O_703,N_17388,N_19365);
xor UO_704 (O_704,N_17790,N_16868);
or UO_705 (O_705,N_18352,N_16157);
and UO_706 (O_706,N_15057,N_17251);
or UO_707 (O_707,N_19995,N_15066);
or UO_708 (O_708,N_17992,N_15806);
nor UO_709 (O_709,N_19531,N_16304);
nand UO_710 (O_710,N_16333,N_18690);
and UO_711 (O_711,N_19803,N_18102);
or UO_712 (O_712,N_15444,N_18767);
or UO_713 (O_713,N_18042,N_16641);
and UO_714 (O_714,N_18219,N_17861);
and UO_715 (O_715,N_17812,N_19898);
xnor UO_716 (O_716,N_17655,N_16610);
nor UO_717 (O_717,N_18326,N_15566);
nor UO_718 (O_718,N_18443,N_17874);
nand UO_719 (O_719,N_18489,N_18883);
or UO_720 (O_720,N_18504,N_17392);
nor UO_721 (O_721,N_18583,N_18281);
xor UO_722 (O_722,N_19963,N_16616);
or UO_723 (O_723,N_19572,N_16082);
nand UO_724 (O_724,N_16635,N_17021);
and UO_725 (O_725,N_18778,N_17313);
xnor UO_726 (O_726,N_19363,N_16653);
nand UO_727 (O_727,N_19653,N_17587);
nor UO_728 (O_728,N_18910,N_18855);
nor UO_729 (O_729,N_15308,N_18525);
nor UO_730 (O_730,N_16153,N_15916);
nor UO_731 (O_731,N_17341,N_18792);
or UO_732 (O_732,N_19164,N_16116);
nand UO_733 (O_733,N_15249,N_16459);
xnor UO_734 (O_734,N_19674,N_17254);
nand UO_735 (O_735,N_16415,N_17019);
nand UO_736 (O_736,N_17302,N_16495);
xnor UO_737 (O_737,N_16755,N_15384);
nand UO_738 (O_738,N_17745,N_19196);
nor UO_739 (O_739,N_19501,N_19606);
or UO_740 (O_740,N_16539,N_15768);
nor UO_741 (O_741,N_17617,N_17519);
nand UO_742 (O_742,N_19987,N_17169);
and UO_743 (O_743,N_15722,N_19439);
nand UO_744 (O_744,N_17078,N_18734);
xor UO_745 (O_745,N_15563,N_17393);
xnor UO_746 (O_746,N_18726,N_15082);
nor UO_747 (O_747,N_17211,N_16380);
nand UO_748 (O_748,N_16498,N_16595);
xor UO_749 (O_749,N_17187,N_17044);
xnor UO_750 (O_750,N_18735,N_18879);
and UO_751 (O_751,N_16515,N_19065);
or UO_752 (O_752,N_16686,N_19990);
xnor UO_753 (O_753,N_19016,N_15477);
and UO_754 (O_754,N_19822,N_16947);
nand UO_755 (O_755,N_17742,N_18140);
nor UO_756 (O_756,N_19112,N_18550);
xor UO_757 (O_757,N_18474,N_15549);
nand UO_758 (O_758,N_15766,N_16798);
xnor UO_759 (O_759,N_17872,N_16667);
or UO_760 (O_760,N_19458,N_15592);
nand UO_761 (O_761,N_18625,N_17440);
nand UO_762 (O_762,N_15512,N_17948);
nand UO_763 (O_763,N_18382,N_16199);
nand UO_764 (O_764,N_16000,N_15745);
nor UO_765 (O_765,N_19858,N_18248);
nor UO_766 (O_766,N_19031,N_17423);
or UO_767 (O_767,N_17842,N_17472);
xor UO_768 (O_768,N_16698,N_17694);
or UO_769 (O_769,N_19479,N_17400);
and UO_770 (O_770,N_18739,N_18500);
or UO_771 (O_771,N_17076,N_19186);
nand UO_772 (O_772,N_17285,N_16701);
nand UO_773 (O_773,N_19053,N_16626);
or UO_774 (O_774,N_19930,N_19980);
and UO_775 (O_775,N_15553,N_15139);
or UO_776 (O_776,N_15440,N_16326);
nor UO_777 (O_777,N_16964,N_18925);
nand UO_778 (O_778,N_18939,N_16651);
or UO_779 (O_779,N_17577,N_18544);
xor UO_780 (O_780,N_19701,N_18356);
nor UO_781 (O_781,N_15939,N_17396);
nor UO_782 (O_782,N_16774,N_19399);
nor UO_783 (O_783,N_18468,N_18236);
nor UO_784 (O_784,N_16999,N_15839);
nand UO_785 (O_785,N_17128,N_17330);
nor UO_786 (O_786,N_19117,N_19832);
nor UO_787 (O_787,N_16044,N_15027);
or UO_788 (O_788,N_16080,N_18719);
nand UO_789 (O_789,N_16147,N_17561);
or UO_790 (O_790,N_15750,N_15207);
or UO_791 (O_791,N_17608,N_19663);
nand UO_792 (O_792,N_17480,N_18865);
nand UO_793 (O_793,N_19177,N_15171);
nand UO_794 (O_794,N_15911,N_19919);
nand UO_795 (O_795,N_17505,N_17667);
or UO_796 (O_796,N_18665,N_19396);
or UO_797 (O_797,N_17891,N_15312);
and UO_798 (O_798,N_17358,N_17074);
xor UO_799 (O_799,N_17103,N_15137);
and UO_800 (O_800,N_19493,N_17557);
and UO_801 (O_801,N_15198,N_19910);
nor UO_802 (O_802,N_19584,N_19132);
or UO_803 (O_803,N_16455,N_18328);
and UO_804 (O_804,N_15986,N_19816);
and UO_805 (O_805,N_19855,N_18675);
nand UO_806 (O_806,N_16852,N_19159);
or UO_807 (O_807,N_15270,N_18505);
nand UO_808 (O_808,N_17699,N_15892);
or UO_809 (O_809,N_16447,N_15049);
or UO_810 (O_810,N_19316,N_18912);
and UO_811 (O_811,N_16929,N_18679);
and UO_812 (O_812,N_18548,N_17316);
xor UO_813 (O_813,N_17692,N_15293);
and UO_814 (O_814,N_18193,N_19310);
or UO_815 (O_815,N_16652,N_15719);
and UO_816 (O_816,N_17126,N_18621);
nor UO_817 (O_817,N_19708,N_16849);
xor UO_818 (O_818,N_16841,N_15610);
and UO_819 (O_819,N_15938,N_19714);
or UO_820 (O_820,N_16614,N_15133);
or UO_821 (O_821,N_18124,N_16994);
nand UO_822 (O_822,N_16581,N_18670);
xor UO_823 (O_823,N_18646,N_17530);
and UO_824 (O_824,N_16844,N_17175);
and UO_825 (O_825,N_15170,N_18892);
or UO_826 (O_826,N_16237,N_18529);
and UO_827 (O_827,N_19678,N_19992);
or UO_828 (O_828,N_15140,N_16908);
or UO_829 (O_829,N_18063,N_18568);
nand UO_830 (O_830,N_19819,N_18277);
xnor UO_831 (O_831,N_15529,N_15796);
nand UO_832 (O_832,N_19958,N_16813);
nand UO_833 (O_833,N_16440,N_16179);
or UO_834 (O_834,N_19007,N_19810);
and UO_835 (O_835,N_15962,N_19496);
and UO_836 (O_836,N_18901,N_18842);
nand UO_837 (O_837,N_17839,N_19917);
nor UO_838 (O_838,N_15337,N_17049);
nor UO_839 (O_839,N_18703,N_18510);
or UO_840 (O_840,N_15465,N_16563);
nand UO_841 (O_841,N_18783,N_17034);
nand UO_842 (O_842,N_15554,N_16019);
xnor UO_843 (O_843,N_16154,N_19041);
and UO_844 (O_844,N_15144,N_15226);
and UO_845 (O_845,N_15223,N_17125);
and UO_846 (O_846,N_19323,N_19845);
nor UO_847 (O_847,N_18601,N_19146);
nor UO_848 (O_848,N_15125,N_19361);
nand UO_849 (O_849,N_15276,N_19926);
nor UO_850 (O_850,N_15994,N_15772);
and UO_851 (O_851,N_15516,N_18967);
nor UO_852 (O_852,N_16697,N_16062);
nand UO_853 (O_853,N_16001,N_16272);
xor UO_854 (O_854,N_15627,N_18603);
nor UO_855 (O_855,N_16658,N_17218);
and UO_856 (O_856,N_17736,N_18227);
nand UO_857 (O_857,N_16948,N_15037);
nand UO_858 (O_858,N_16232,N_17977);
or UO_859 (O_859,N_19213,N_19866);
xnor UO_860 (O_860,N_15736,N_16298);
nand UO_861 (O_861,N_15095,N_19124);
or UO_862 (O_862,N_19135,N_19760);
or UO_863 (O_863,N_16570,N_16679);
and UO_864 (O_864,N_17850,N_17244);
and UO_865 (O_865,N_16496,N_16770);
nor UO_866 (O_866,N_19184,N_18163);
nand UO_867 (O_867,N_16901,N_18306);
or UO_868 (O_868,N_18765,N_16143);
nand UO_869 (O_869,N_19978,N_15924);
or UO_870 (O_870,N_16335,N_19019);
or UO_871 (O_871,N_16126,N_17680);
xor UO_872 (O_872,N_18068,N_16913);
xor UO_873 (O_873,N_19338,N_18371);
nand UO_874 (O_874,N_15883,N_15618);
and UO_875 (O_875,N_16742,N_18334);
nand UO_876 (O_876,N_19315,N_15405);
and UO_877 (O_877,N_19142,N_19872);
or UO_878 (O_878,N_19756,N_16984);
and UO_879 (O_879,N_15570,N_18780);
nor UO_880 (O_880,N_19547,N_16024);
and UO_881 (O_881,N_17890,N_15784);
or UO_882 (O_882,N_18708,N_15639);
nor UO_883 (O_883,N_17672,N_15704);
nand UO_884 (O_884,N_15634,N_15459);
nand UO_885 (O_885,N_18133,N_19274);
xor UO_886 (O_886,N_18286,N_15868);
and UO_887 (O_887,N_16911,N_15774);
nand UO_888 (O_888,N_19347,N_17146);
nor UO_889 (O_889,N_19118,N_18885);
xnor UO_890 (O_890,N_16749,N_17075);
xor UO_891 (O_891,N_19508,N_15735);
and UO_892 (O_892,N_16855,N_18584);
or UO_893 (O_893,N_15749,N_19581);
nand UO_894 (O_894,N_17724,N_19475);
nand UO_895 (O_895,N_17478,N_16210);
nor UO_896 (O_896,N_18275,N_15201);
nand UO_897 (O_897,N_17057,N_17191);
and UO_898 (O_898,N_15320,N_16599);
or UO_899 (O_899,N_16597,N_16718);
xnor UO_900 (O_900,N_18872,N_16284);
nor UO_901 (O_901,N_19058,N_18482);
nand UO_902 (O_902,N_15489,N_19299);
xnor UO_903 (O_903,N_19776,N_19749);
or UO_904 (O_904,N_18471,N_17298);
nand UO_905 (O_905,N_16371,N_15259);
and UO_906 (O_906,N_18037,N_16624);
nor UO_907 (O_907,N_19755,N_19694);
nand UO_908 (O_908,N_15426,N_16834);
nor UO_909 (O_909,N_15576,N_15191);
nand UO_910 (O_910,N_16925,N_17326);
xor UO_911 (O_911,N_15097,N_15094);
nor UO_912 (O_912,N_18336,N_19021);
and UO_913 (O_913,N_16413,N_18120);
nand UO_914 (O_914,N_18952,N_16725);
xnor UO_915 (O_915,N_15673,N_19015);
and UO_916 (O_916,N_19861,N_15262);
or UO_917 (O_917,N_19830,N_16428);
and UO_918 (O_918,N_17716,N_17493);
xor UO_919 (O_919,N_16021,N_19718);
xor UO_920 (O_920,N_16003,N_19309);
nand UO_921 (O_921,N_17678,N_19125);
and UO_922 (O_922,N_17525,N_19745);
xnor UO_923 (O_923,N_16040,N_18161);
nor UO_924 (O_924,N_17688,N_18437);
and UO_925 (O_925,N_15266,N_16340);
nor UO_926 (O_926,N_18374,N_18395);
or UO_927 (O_927,N_18157,N_15915);
or UO_928 (O_928,N_16751,N_19151);
nand UO_929 (O_929,N_17991,N_15447);
and UO_930 (O_930,N_15390,N_16385);
xnor UO_931 (O_931,N_15598,N_15482);
and UO_932 (O_932,N_19672,N_17232);
nor UO_933 (O_933,N_15172,N_18475);
nor UO_934 (O_934,N_15195,N_18880);
nand UO_935 (O_935,N_17372,N_19113);
or UO_936 (O_936,N_17061,N_18652);
and UO_937 (O_937,N_15601,N_19449);
nor UO_938 (O_938,N_16004,N_19918);
or UO_939 (O_939,N_17395,N_18094);
xnor UO_940 (O_940,N_19032,N_18677);
and UO_941 (O_941,N_16703,N_18321);
xor UO_942 (O_942,N_19836,N_15793);
nor UO_943 (O_943,N_19035,N_17209);
nor UO_944 (O_944,N_16724,N_15599);
nand UO_945 (O_945,N_18717,N_15007);
nor UO_946 (O_946,N_19080,N_17843);
or UO_947 (O_947,N_16517,N_15674);
or UO_948 (O_948,N_18189,N_18092);
and UO_949 (O_949,N_15580,N_19335);
or UO_950 (O_950,N_17064,N_15215);
xnor UO_951 (O_951,N_18266,N_16914);
nor UO_952 (O_952,N_16166,N_17283);
nor UO_953 (O_953,N_19066,N_16526);
nand UO_954 (O_954,N_15524,N_19483);
nand UO_955 (O_955,N_18676,N_15114);
and UO_956 (O_956,N_19212,N_16800);
or UO_957 (O_957,N_15763,N_15178);
nand UO_958 (O_958,N_18898,N_17248);
and UO_959 (O_959,N_18035,N_18838);
and UO_960 (O_960,N_19039,N_18686);
xnor UO_961 (O_961,N_18049,N_16988);
xor UO_962 (O_962,N_19920,N_19788);
or UO_963 (O_963,N_18455,N_18831);
and UO_964 (O_964,N_18387,N_17514);
xor UO_965 (O_965,N_15708,N_19900);
nor UO_966 (O_966,N_16513,N_18867);
and UO_967 (O_967,N_17773,N_17296);
and UO_968 (O_968,N_19198,N_19764);
nand UO_969 (O_969,N_16308,N_17732);
xor UO_970 (O_970,N_17426,N_18606);
xor UO_971 (O_971,N_18516,N_15824);
nand UO_972 (O_972,N_16808,N_19295);
xor UO_973 (O_973,N_18829,N_19733);
nor UO_974 (O_974,N_15850,N_15348);
nand UO_975 (O_975,N_15064,N_15778);
nand UO_976 (O_976,N_17467,N_15016);
nor UO_977 (O_977,N_17646,N_19156);
nand UO_978 (O_978,N_18003,N_18810);
and UO_979 (O_979,N_18822,N_17318);
nand UO_980 (O_980,N_18801,N_17600);
or UO_981 (O_981,N_19769,N_17703);
nand UO_982 (O_982,N_16625,N_18337);
or UO_983 (O_983,N_15048,N_19103);
nor UO_984 (O_984,N_15628,N_16857);
nor UO_985 (O_985,N_19498,N_18796);
or UO_986 (O_986,N_18046,N_16799);
or UO_987 (O_987,N_15686,N_17764);
xnor UO_988 (O_988,N_18757,N_16883);
or UO_989 (O_989,N_17051,N_17242);
xnor UO_990 (O_990,N_19465,N_18764);
or UO_991 (O_991,N_17077,N_15255);
and UO_992 (O_992,N_16162,N_19741);
or UO_993 (O_993,N_16018,N_19870);
xor UO_994 (O_994,N_16342,N_16379);
nand UO_995 (O_995,N_15112,N_15289);
xor UO_996 (O_996,N_16812,N_19972);
xor UO_997 (O_997,N_17586,N_17017);
nand UO_998 (O_998,N_17041,N_16183);
or UO_999 (O_999,N_17084,N_15461);
or UO_1000 (O_1000,N_15228,N_15351);
xor UO_1001 (O_1001,N_17328,N_15277);
or UO_1002 (O_1002,N_19999,N_17825);
and UO_1003 (O_1003,N_17431,N_16814);
nand UO_1004 (O_1004,N_15365,N_16942);
xnor UO_1005 (O_1005,N_19229,N_16255);
nor UO_1006 (O_1006,N_15517,N_18055);
nor UO_1007 (O_1007,N_16445,N_19759);
xnor UO_1008 (O_1008,N_18372,N_19506);
nor UO_1009 (O_1009,N_19511,N_15982);
and UO_1010 (O_1010,N_17762,N_17500);
nor UO_1011 (O_1011,N_16373,N_17999);
nor UO_1012 (O_1012,N_15045,N_15149);
nor UO_1013 (O_1013,N_16227,N_16768);
xnor UO_1014 (O_1014,N_16892,N_18287);
or UO_1015 (O_1015,N_19687,N_17517);
and UO_1016 (O_1016,N_19378,N_15285);
or UO_1017 (O_1017,N_16780,N_17857);
xnor UO_1018 (O_1018,N_17245,N_19411);
or UO_1019 (O_1019,N_19451,N_17928);
and UO_1020 (O_1020,N_16140,N_15129);
nand UO_1021 (O_1021,N_19136,N_19357);
nor UO_1022 (O_1022,N_17294,N_17747);
or UO_1023 (O_1023,N_18188,N_19794);
nor UO_1024 (O_1024,N_19350,N_18696);
and UO_1025 (O_1025,N_16438,N_16848);
xnor UO_1026 (O_1026,N_15219,N_18469);
nor UO_1027 (O_1027,N_18131,N_19050);
and UO_1028 (O_1028,N_15456,N_19960);
or UO_1029 (O_1029,N_17776,N_16981);
xor UO_1030 (O_1030,N_15286,N_16582);
or UO_1031 (O_1031,N_17606,N_17056);
xor UO_1032 (O_1032,N_17534,N_17106);
or UO_1033 (O_1033,N_16875,N_16877);
xor UO_1034 (O_1034,N_19371,N_16125);
and UO_1035 (O_1035,N_17208,N_17551);
nand UO_1036 (O_1036,N_18257,N_16215);
and UO_1037 (O_1037,N_15847,N_17112);
nand UO_1038 (O_1038,N_16928,N_15208);
xor UO_1039 (O_1039,N_18593,N_16680);
and UO_1040 (O_1040,N_16643,N_19279);
and UO_1041 (O_1041,N_18467,N_15245);
or UO_1042 (O_1042,N_19717,N_18206);
or UO_1043 (O_1043,N_17737,N_18013);
and UO_1044 (O_1044,N_18168,N_15604);
or UO_1045 (O_1045,N_19172,N_15316);
nand UO_1046 (O_1046,N_17927,N_17721);
nand UO_1047 (O_1047,N_17836,N_15989);
and UO_1048 (O_1048,N_18579,N_15976);
nor UO_1049 (O_1049,N_17761,N_17625);
nor UO_1050 (O_1050,N_19332,N_18694);
nor UO_1051 (O_1051,N_16325,N_17804);
xor UO_1052 (O_1052,N_19168,N_16396);
nor UO_1053 (O_1053,N_18205,N_17157);
and UO_1054 (O_1054,N_18090,N_15605);
and UO_1055 (O_1055,N_19466,N_18396);
xnor UO_1056 (O_1056,N_17241,N_19951);
nand UO_1057 (O_1057,N_17639,N_18866);
and UO_1058 (O_1058,N_16354,N_18802);
nand UO_1059 (O_1059,N_15437,N_16777);
nand UO_1060 (O_1060,N_15290,N_19564);
xnor UO_1061 (O_1061,N_19087,N_18151);
nand UO_1062 (O_1062,N_17354,N_19170);
nand UO_1063 (O_1063,N_17870,N_15640);
xor UO_1064 (O_1064,N_15159,N_19267);
xnor UO_1065 (O_1065,N_19380,N_15997);
nor UO_1066 (O_1066,N_19121,N_18558);
and UO_1067 (O_1067,N_19611,N_18793);
and UO_1068 (O_1068,N_17448,N_17135);
or UO_1069 (O_1069,N_17779,N_15753);
nor UO_1070 (O_1070,N_18226,N_19026);
xor UO_1071 (O_1071,N_16331,N_17887);
nor UO_1072 (O_1072,N_15755,N_15356);
nand UO_1073 (O_1073,N_19728,N_16528);
nand UO_1074 (O_1074,N_17220,N_17445);
nor UO_1075 (O_1075,N_15721,N_15210);
xnor UO_1076 (O_1076,N_15833,N_19726);
and UO_1077 (O_1077,N_15136,N_19552);
nor UO_1078 (O_1078,N_16674,N_16324);
nor UO_1079 (O_1079,N_16959,N_17831);
or UO_1080 (O_1080,N_18114,N_19345);
or UO_1081 (O_1081,N_19840,N_15664);
nor UO_1082 (O_1082,N_18129,N_19059);
nand UO_1083 (O_1083,N_18175,N_18597);
nor UO_1084 (O_1084,N_16992,N_17484);
nor UO_1085 (O_1085,N_17817,N_17235);
and UO_1086 (O_1086,N_19610,N_16164);
nor UO_1087 (O_1087,N_19929,N_19876);
or UO_1088 (O_1088,N_15175,N_19905);
and UO_1089 (O_1089,N_15059,N_17133);
nand UO_1090 (O_1090,N_17359,N_19218);
nor UO_1091 (O_1091,N_18397,N_16457);
nor UO_1092 (O_1092,N_16448,N_18790);
or UO_1093 (O_1093,N_18594,N_16054);
nand UO_1094 (O_1094,N_17844,N_15870);
nor UO_1095 (O_1095,N_18743,N_18843);
and UO_1096 (O_1096,N_18749,N_19956);
nor UO_1097 (O_1097,N_17181,N_17559);
or UO_1098 (O_1098,N_18250,N_18231);
nand UO_1099 (O_1099,N_18246,N_16281);
xor UO_1100 (O_1100,N_15474,N_19851);
or UO_1101 (O_1101,N_19246,N_19460);
or UO_1102 (O_1102,N_16041,N_16706);
xnor UO_1103 (O_1103,N_16292,N_15980);
xor UO_1104 (O_1104,N_16473,N_16978);
or UO_1105 (O_1105,N_17214,N_19869);
nor UO_1106 (O_1106,N_16461,N_18023);
and UO_1107 (O_1107,N_18622,N_16204);
and UO_1108 (O_1108,N_15256,N_16990);
xor UO_1109 (O_1109,N_16416,N_17632);
nor UO_1110 (O_1110,N_17532,N_15656);
nand UO_1111 (O_1111,N_17262,N_18521);
nor UO_1112 (O_1112,N_19385,N_19706);
or UO_1113 (O_1113,N_15515,N_19686);
or UO_1114 (O_1114,N_18172,N_15926);
xor UO_1115 (O_1115,N_16338,N_16827);
nand UO_1116 (O_1116,N_18247,N_17515);
nor UO_1117 (O_1117,N_16726,N_16632);
xnor UO_1118 (O_1118,N_19537,N_18261);
xnor UO_1119 (O_1119,N_15672,N_17069);
xor UO_1120 (O_1120,N_16574,N_19577);
nand UO_1121 (O_1121,N_17014,N_19558);
or UO_1122 (O_1122,N_17936,N_19504);
nor UO_1123 (O_1123,N_15801,N_18222);
nor UO_1124 (O_1124,N_19382,N_16784);
or UO_1125 (O_1125,N_16722,N_19413);
or UO_1126 (O_1126,N_15522,N_15455);
xor UO_1127 (O_1127,N_18803,N_18800);
and UO_1128 (O_1128,N_15273,N_17569);
nand UO_1129 (O_1129,N_17159,N_15143);
xnor UO_1130 (O_1130,N_19444,N_16532);
nor UO_1131 (O_1131,N_16191,N_15999);
or UO_1132 (O_1132,N_16289,N_19076);
or UO_1133 (O_1133,N_17404,N_18398);
nor UO_1134 (O_1134,N_18268,N_16058);
or UO_1135 (O_1135,N_17444,N_18491);
and UO_1136 (O_1136,N_18511,N_15400);
xor UO_1137 (O_1137,N_15684,N_17325);
nand UO_1138 (O_1138,N_15101,N_18278);
nand UO_1139 (O_1139,N_16278,N_19442);
and UO_1140 (O_1140,N_16211,N_19641);
nor UO_1141 (O_1141,N_18377,N_15947);
and UO_1142 (O_1142,N_17073,N_18135);
xnor UO_1143 (O_1143,N_17407,N_16847);
or UO_1144 (O_1144,N_16660,N_16305);
or UO_1145 (O_1145,N_17305,N_16573);
nand UO_1146 (O_1146,N_16280,N_15859);
or UO_1147 (O_1147,N_17813,N_19149);
or UO_1148 (O_1148,N_18498,N_16746);
nor UO_1149 (O_1149,N_16894,N_19349);
nand UO_1150 (O_1150,N_19668,N_18769);
or UO_1151 (O_1151,N_16465,N_18262);
nor UO_1152 (O_1152,N_19358,N_19471);
or UO_1153 (O_1153,N_15525,N_18502);
nor UO_1154 (O_1154,N_17677,N_18573);
nand UO_1155 (O_1155,N_15899,N_16266);
and UO_1156 (O_1156,N_15608,N_16763);
nand UO_1157 (O_1157,N_17748,N_15777);
nor UO_1158 (O_1158,N_16102,N_18179);
nand UO_1159 (O_1159,N_17152,N_18045);
xor UO_1160 (O_1160,N_18766,N_15398);
and UO_1161 (O_1161,N_18526,N_16228);
nand UO_1162 (O_1162,N_19270,N_17981);
or UO_1163 (O_1163,N_19012,N_18224);
or UO_1164 (O_1164,N_15591,N_18392);
and UO_1165 (O_1165,N_17782,N_18305);
and UO_1166 (O_1166,N_17186,N_15550);
nand UO_1167 (O_1167,N_16910,N_17198);
nor UO_1168 (O_1168,N_15258,N_17153);
nand UO_1169 (O_1169,N_18442,N_16435);
xor UO_1170 (O_1170,N_16969,N_16600);
or UO_1171 (O_1171,N_18738,N_15243);
nand UO_1172 (O_1172,N_18964,N_18488);
or UO_1173 (O_1173,N_15594,N_17161);
or UO_1174 (O_1174,N_15153,N_18478);
nand UO_1175 (O_1175,N_17121,N_17660);
xnor UO_1176 (O_1176,N_17654,N_19100);
xnor UO_1177 (O_1177,N_17938,N_16621);
nand UO_1178 (O_1178,N_15921,N_17080);
nand UO_1179 (O_1179,N_17575,N_18807);
and UO_1180 (O_1180,N_18659,N_17696);
xor UO_1181 (O_1181,N_15283,N_17363);
and UO_1182 (O_1182,N_18714,N_18021);
nand UO_1183 (O_1183,N_18173,N_18798);
nor UO_1184 (O_1184,N_19798,N_15611);
nor UO_1185 (O_1185,N_15846,N_15361);
nor UO_1186 (O_1186,N_17311,N_18854);
nor UO_1187 (O_1187,N_15093,N_18538);
nor UO_1188 (O_1188,N_19565,N_15490);
xnor UO_1189 (O_1189,N_18481,N_18870);
nand UO_1190 (O_1190,N_16764,N_16939);
or UO_1191 (O_1191,N_17767,N_19046);
nand UO_1192 (O_1192,N_18950,N_18715);
nor UO_1193 (O_1193,N_17164,N_19174);
or UO_1194 (O_1194,N_19539,N_19502);
or UO_1195 (O_1195,N_17715,N_17968);
and UO_1196 (O_1196,N_17666,N_15404);
nor UO_1197 (O_1197,N_16407,N_15925);
xor UO_1198 (O_1198,N_19970,N_16893);
xor UO_1199 (O_1199,N_19109,N_19293);
or UO_1200 (O_1200,N_15287,N_17231);
and UO_1201 (O_1201,N_15579,N_16161);
nand UO_1202 (O_1202,N_19643,N_19390);
nand UO_1203 (O_1203,N_17487,N_17269);
and UO_1204 (O_1204,N_18722,N_16372);
or UO_1205 (O_1205,N_16601,N_16432);
nand UO_1206 (O_1206,N_15424,N_15315);
xor UO_1207 (O_1207,N_18532,N_15812);
and UO_1208 (O_1208,N_17443,N_16815);
nand UO_1209 (O_1209,N_17247,N_19814);
nor UO_1210 (O_1210,N_17545,N_17183);
nand UO_1211 (O_1211,N_19860,N_17884);
xnor UO_1212 (O_1212,N_18545,N_16821);
and UO_1213 (O_1213,N_15667,N_15913);
nand UO_1214 (O_1214,N_17634,N_19828);
and UO_1215 (O_1215,N_15179,N_18200);
nor UO_1216 (O_1216,N_19325,N_18636);
and UO_1217 (O_1217,N_19454,N_16398);
nor UO_1218 (O_1218,N_17307,N_17346);
nor UO_1219 (O_1219,N_18282,N_16318);
or UO_1220 (O_1220,N_19950,N_15702);
nand UO_1221 (O_1221,N_15241,N_16367);
xor UO_1222 (O_1222,N_15940,N_18378);
or UO_1223 (O_1223,N_18143,N_19098);
or UO_1224 (O_1224,N_15936,N_15216);
xnor UO_1225 (O_1225,N_19468,N_17744);
or UO_1226 (O_1226,N_19747,N_18984);
xnor UO_1227 (O_1227,N_19837,N_15880);
or UO_1228 (O_1228,N_16088,N_19244);
or UO_1229 (O_1229,N_18693,N_19152);
nand UO_1230 (O_1230,N_19036,N_19167);
xnor UO_1231 (O_1231,N_16267,N_19775);
or UO_1232 (O_1232,N_19679,N_16915);
and UO_1233 (O_1233,N_15685,N_17770);
xor UO_1234 (O_1234,N_19856,N_16073);
xor UO_1235 (O_1235,N_16012,N_16093);
xor UO_1236 (O_1236,N_19780,N_16871);
nand UO_1237 (O_1237,N_19376,N_19651);
nor UO_1238 (O_1238,N_15406,N_18728);
xnor UO_1239 (O_1239,N_19848,N_18450);
nand UO_1240 (O_1240,N_16057,N_19598);
nor UO_1241 (O_1241,N_19650,N_17924);
and UO_1242 (O_1242,N_16158,N_18818);
xnor UO_1243 (O_1243,N_15386,N_17134);
xor UO_1244 (O_1244,N_17735,N_17086);
and UO_1245 (O_1245,N_19092,N_19831);
xor UO_1246 (O_1246,N_19001,N_18642);
and UO_1247 (O_1247,N_17789,N_17337);
or UO_1248 (O_1248,N_18613,N_17596);
and UO_1249 (O_1249,N_18338,N_18386);
xor UO_1250 (O_1250,N_17904,N_16807);
xor UO_1251 (O_1251,N_18033,N_17287);
nor UO_1252 (O_1252,N_15268,N_16953);
xnor UO_1253 (O_1253,N_18312,N_15506);
or UO_1254 (O_1254,N_15993,N_19932);
nor UO_1255 (O_1255,N_16525,N_16785);
and UO_1256 (O_1256,N_15338,N_19437);
xnor UO_1257 (O_1257,N_16194,N_16247);
and UO_1258 (O_1258,N_16545,N_18981);
nor UO_1259 (O_1259,N_15897,N_16558);
nor UO_1260 (O_1260,N_19973,N_15904);
and UO_1261 (O_1261,N_17402,N_17255);
xor UO_1262 (O_1262,N_18414,N_16301);
nand UO_1263 (O_1263,N_16589,N_19090);
and UO_1264 (O_1264,N_18361,N_15089);
or UO_1265 (O_1265,N_18271,N_15305);
and UO_1266 (O_1266,N_17132,N_18586);
xnor UO_1267 (O_1267,N_17425,N_15026);
and UO_1268 (O_1268,N_18680,N_18174);
xnor UO_1269 (O_1269,N_16734,N_15151);
and UO_1270 (O_1270,N_15826,N_19009);
nor UO_1271 (O_1271,N_15452,N_17930);
nor UO_1272 (O_1272,N_16806,N_16716);
and UO_1273 (O_1273,N_19550,N_17155);
nor UO_1274 (O_1274,N_16468,N_15150);
xor UO_1275 (O_1275,N_18640,N_15314);
nand UO_1276 (O_1276,N_15407,N_15771);
xor UO_1277 (O_1277,N_15762,N_16028);
and UO_1278 (O_1278,N_18878,N_16623);
and UO_1279 (O_1279,N_18399,N_18839);
and UO_1280 (O_1280,N_16491,N_19063);
xor UO_1281 (O_1281,N_15711,N_19761);
or UO_1282 (O_1282,N_17853,N_18595);
xnor UO_1283 (O_1283,N_17013,N_18292);
and UO_1284 (O_1284,N_19821,N_15900);
nor UO_1285 (O_1285,N_19702,N_19657);
nand UO_1286 (O_1286,N_18619,N_18216);
and UO_1287 (O_1287,N_17229,N_15373);
nor UO_1288 (O_1288,N_17045,N_17969);
and UO_1289 (O_1289,N_16591,N_17196);
nor UO_1290 (O_1290,N_17550,N_16362);
nand UO_1291 (O_1291,N_15345,N_18207);
nand UO_1292 (O_1292,N_17554,N_15712);
or UO_1293 (O_1293,N_19696,N_19705);
xnor UO_1294 (O_1294,N_18567,N_15011);
nand UO_1295 (O_1295,N_19474,N_19563);
or UO_1296 (O_1296,N_19503,N_19625);
nand UO_1297 (O_1297,N_15300,N_17741);
nor UO_1298 (O_1298,N_18159,N_15099);
xor UO_1299 (O_1299,N_19557,N_18514);
and UO_1300 (O_1300,N_18197,N_16628);
or UO_1301 (O_1301,N_19052,N_17446);
xnor UO_1302 (O_1302,N_18994,N_16477);
or UO_1303 (O_1303,N_17099,N_18052);
nand UO_1304 (O_1304,N_16188,N_17297);
nor UO_1305 (O_1305,N_18422,N_15797);
nor UO_1306 (O_1306,N_15081,N_16268);
or UO_1307 (O_1307,N_16221,N_17967);
xor UO_1308 (O_1308,N_18919,N_16691);
and UO_1309 (O_1309,N_17435,N_17792);
or UO_1310 (O_1310,N_16696,N_18012);
and UO_1311 (O_1311,N_15787,N_18297);
and UO_1312 (O_1312,N_15232,N_15021);
nand UO_1313 (O_1313,N_15036,N_18078);
xor UO_1314 (O_1314,N_17588,N_16538);
nand UO_1315 (O_1315,N_17847,N_15973);
nor UO_1316 (O_1316,N_19621,N_18576);
nand UO_1317 (O_1317,N_16912,N_15342);
and UO_1318 (O_1318,N_16312,N_16329);
nor UO_1319 (O_1319,N_16933,N_18946);
nor UO_1320 (O_1320,N_18430,N_16711);
nand UO_1321 (O_1321,N_17455,N_16253);
nand UO_1322 (O_1322,N_19500,N_16360);
nand UO_1323 (O_1323,N_17971,N_15567);
nor UO_1324 (O_1324,N_18859,N_19536);
nand UO_1325 (O_1325,N_17489,N_16802);
nand UO_1326 (O_1326,N_18434,N_17434);
nor UO_1327 (O_1327,N_18627,N_17405);
and UO_1328 (O_1328,N_17027,N_19160);
or UO_1329 (O_1329,N_16144,N_19101);
nor UO_1330 (O_1330,N_15075,N_16903);
or UO_1331 (O_1331,N_18464,N_15006);
xor UO_1332 (O_1332,N_17207,N_17107);
and UO_1333 (O_1333,N_16096,N_18196);
or UO_1334 (O_1334,N_18075,N_19082);
nand UO_1335 (O_1335,N_19389,N_18713);
and UO_1336 (O_1336,N_19202,N_15746);
nor UO_1337 (O_1337,N_15677,N_17145);
nor UO_1338 (O_1338,N_18937,N_18832);
nor UO_1339 (O_1339,N_19002,N_16049);
and UO_1340 (O_1340,N_16717,N_15202);
or UO_1341 (O_1341,N_17315,N_16782);
xor UO_1342 (O_1342,N_19942,N_17182);
and UO_1343 (O_1343,N_16436,N_18758);
or UO_1344 (O_1344,N_18750,N_18340);
or UO_1345 (O_1345,N_18697,N_19355);
or UO_1346 (O_1346,N_17626,N_16645);
nor UO_1347 (O_1347,N_17170,N_18988);
xor UO_1348 (O_1348,N_16556,N_15272);
nand UO_1349 (O_1349,N_18436,N_16251);
xor UO_1350 (O_1350,N_15032,N_15872);
nor UO_1351 (O_1351,N_19269,N_15019);
nand UO_1352 (O_1352,N_15058,N_19311);
nor UO_1353 (O_1353,N_18288,N_17613);
nand UO_1354 (O_1354,N_17158,N_15166);
and UO_1355 (O_1355,N_17720,N_17602);
xor UO_1356 (O_1356,N_19773,N_18341);
nand UO_1357 (O_1357,N_19289,N_19591);
xnor UO_1358 (O_1358,N_15971,N_16476);
and UO_1359 (O_1359,N_19423,N_18459);
and UO_1360 (O_1360,N_19166,N_17114);
and UO_1361 (O_1361,N_16693,N_18091);
or UO_1362 (O_1362,N_17438,N_17743);
and UO_1363 (O_1363,N_19356,N_15748);
nor UO_1364 (O_1364,N_18001,N_18082);
and UO_1365 (O_1365,N_15115,N_18953);
xnor UO_1366 (O_1366,N_16033,N_16038);
xnor UO_1367 (O_1367,N_15761,N_19575);
xor UO_1368 (O_1368,N_15269,N_19225);
and UO_1369 (O_1369,N_16444,N_17510);
xor UO_1370 (O_1370,N_17148,N_17649);
nor UO_1371 (O_1371,N_16467,N_19038);
and UO_1372 (O_1372,N_17546,N_17821);
or UO_1373 (O_1373,N_18874,N_16433);
nand UO_1374 (O_1374,N_19128,N_16265);
xnor UO_1375 (O_1375,N_18142,N_18890);
or UO_1376 (O_1376,N_15134,N_16002);
and UO_1377 (O_1377,N_15430,N_18225);
and UO_1378 (O_1378,N_16607,N_16076);
or UO_1379 (O_1379,N_15528,N_18019);
nor UO_1380 (O_1380,N_19971,N_17982);
and UO_1381 (O_1381,N_16264,N_16212);
nand UO_1382 (O_1382,N_15557,N_15678);
nor UO_1383 (O_1383,N_15803,N_18934);
and UO_1384 (O_1384,N_15534,N_16880);
or UO_1385 (O_1385,N_18553,N_19632);
nand UO_1386 (O_1386,N_17020,N_19833);
or UO_1387 (O_1387,N_19183,N_17052);
or UO_1388 (O_1388,N_17256,N_18327);
or UO_1389 (O_1389,N_18531,N_15321);
nand UO_1390 (O_1390,N_15291,N_19171);
nor UO_1391 (O_1391,N_18368,N_16733);
xor UO_1392 (O_1392,N_17188,N_16750);
or UO_1393 (O_1393,N_15593,N_16023);
nor UO_1394 (O_1394,N_19408,N_15135);
nor UO_1395 (O_1395,N_16503,N_18220);
and UO_1396 (O_1396,N_19777,N_17179);
xor UO_1397 (O_1397,N_18418,N_19983);
or UO_1398 (O_1398,N_17854,N_19272);
nor UO_1399 (O_1399,N_15085,N_17031);
xor UO_1400 (O_1400,N_19664,N_19304);
or UO_1401 (O_1401,N_16053,N_15878);
nand UO_1402 (O_1402,N_19217,N_16897);
or UO_1403 (O_1403,N_16611,N_19061);
nand UO_1404 (O_1404,N_17117,N_17612);
or UO_1405 (O_1405,N_16817,N_17876);
or UO_1406 (O_1406,N_19324,N_19953);
and UO_1407 (O_1407,N_17215,N_17894);
and UO_1408 (O_1408,N_16540,N_19240);
xor UO_1409 (O_1409,N_19616,N_18592);
nor UO_1410 (O_1410,N_18927,N_17572);
and UO_1411 (O_1411,N_17729,N_17279);
or UO_1412 (O_1412,N_16101,N_19863);
or UO_1413 (O_1413,N_17674,N_15090);
or UO_1414 (O_1414,N_18989,N_15799);
and UO_1415 (O_1415,N_17138,N_16458);
nand UO_1416 (O_1416,N_15802,N_16704);
and UO_1417 (O_1417,N_19871,N_17389);
and UO_1418 (O_1418,N_15838,N_19432);
or UO_1419 (O_1419,N_17263,N_15729);
nand UO_1420 (O_1420,N_18929,N_17197);
nor UO_1421 (O_1421,N_18921,N_16353);
and UO_1422 (O_1422,N_15720,N_16394);
xor UO_1423 (O_1423,N_17091,N_16508);
and UO_1424 (O_1424,N_18071,N_17994);
xnor UO_1425 (O_1425,N_17521,N_17939);
xor UO_1426 (O_1426,N_19381,N_17252);
and UO_1427 (O_1427,N_18270,N_17371);
nand UO_1428 (O_1428,N_19071,N_15326);
xor UO_1429 (O_1429,N_15495,N_15963);
and UO_1430 (O_1430,N_18881,N_17233);
xnor UO_1431 (O_1431,N_16328,N_17486);
nand UO_1432 (O_1432,N_19419,N_17946);
and UO_1433 (O_1433,N_19709,N_17277);
nand UO_1434 (O_1434,N_17641,N_19957);
or UO_1435 (O_1435,N_17902,N_19153);
nor UO_1436 (O_1436,N_16131,N_18177);
or UO_1437 (O_1437,N_18470,N_16169);
or UO_1438 (O_1438,N_19336,N_19027);
nor UO_1439 (O_1439,N_17327,N_15595);
nor UO_1440 (O_1440,N_16809,N_17907);
or UO_1441 (O_1441,N_17709,N_15463);
nor UO_1442 (O_1442,N_19277,N_16516);
and UO_1443 (O_1443,N_19542,N_17950);
xnor UO_1444 (O_1444,N_15369,N_17643);
nand UO_1445 (O_1445,N_19818,N_15728);
or UO_1446 (O_1446,N_17711,N_18139);
nand UO_1447 (O_1447,N_16546,N_16879);
and UO_1448 (O_1448,N_15020,N_16421);
nor UO_1449 (O_1449,N_18781,N_15324);
or UO_1450 (O_1450,N_18702,N_18274);
or UO_1451 (O_1451,N_16469,N_17739);
nor UO_1452 (O_1452,N_16286,N_16014);
xor UO_1453 (O_1453,N_19138,N_17698);
and UO_1454 (O_1454,N_15607,N_19893);
nand UO_1455 (O_1455,N_19443,N_18772);
nand UO_1456 (O_1456,N_17881,N_18428);
nor UO_1457 (O_1457,N_17424,N_18733);
nand UO_1458 (O_1458,N_19744,N_17653);
nor UO_1459 (O_1459,N_18407,N_18256);
xor UO_1460 (O_1460,N_17043,N_17282);
xnor UO_1461 (O_1461,N_19976,N_18007);
nor UO_1462 (O_1462,N_18105,N_15756);
xnor UO_1463 (O_1463,N_19049,N_19685);
nand UO_1464 (O_1464,N_17165,N_16544);
or UO_1465 (O_1465,N_15660,N_17089);
or UO_1466 (O_1466,N_16618,N_17348);
xor UO_1467 (O_1467,N_18635,N_18951);
and UO_1468 (O_1468,N_15944,N_19008);
nor UO_1469 (O_1469,N_19436,N_19879);
and UO_1470 (O_1470,N_18737,N_16317);
or UO_1471 (O_1471,N_17645,N_18522);
and UO_1472 (O_1472,N_18922,N_15582);
xnor UO_1473 (O_1473,N_17603,N_17449);
nand UO_1474 (O_1474,N_16114,N_18239);
and UO_1475 (O_1475,N_15977,N_19713);
xor UO_1476 (O_1476,N_18523,N_15483);
or UO_1477 (O_1477,N_17465,N_17683);
and UO_1478 (O_1478,N_18888,N_18000);
and UO_1479 (O_1479,N_17734,N_19407);
or UO_1480 (O_1480,N_18689,N_15862);
and UO_1481 (O_1481,N_19613,N_16288);
and UO_1482 (O_1482,N_15564,N_18480);
or UO_1483 (O_1483,N_19491,N_18543);
nor UO_1484 (O_1484,N_15840,N_15327);
nand UO_1485 (O_1485,N_18907,N_15017);
nor UO_1486 (O_1486,N_19996,N_19313);
xor UO_1487 (O_1487,N_17583,N_17038);
xor UO_1488 (O_1488,N_19081,N_18788);
nor UO_1489 (O_1489,N_18310,N_18875);
or UO_1490 (O_1490,N_16074,N_15830);
and UO_1491 (O_1491,N_15067,N_17249);
and UO_1492 (O_1492,N_17124,N_18760);
nand UO_1493 (O_1493,N_15038,N_17200);
nand UO_1494 (O_1494,N_15116,N_15044);
nor UO_1495 (O_1495,N_17848,N_15341);
nand UO_1496 (O_1496,N_17566,N_19846);
and UO_1497 (O_1497,N_19129,N_17062);
and UO_1498 (O_1498,N_15556,N_18944);
nor UO_1499 (O_1499,N_18709,N_19559);
and UO_1500 (O_1500,N_15206,N_16285);
xnor UO_1501 (O_1501,N_15488,N_18009);
and UO_1502 (O_1502,N_18448,N_18185);
or UO_1503 (O_1503,N_16938,N_18253);
and UO_1504 (O_1504,N_17447,N_17841);
xor UO_1505 (O_1505,N_18669,N_16779);
nor UO_1506 (O_1506,N_17258,N_16506);
or UO_1507 (O_1507,N_19676,N_18462);
or UO_1508 (O_1508,N_16766,N_16242);
or UO_1509 (O_1509,N_16207,N_18265);
xor UO_1510 (O_1510,N_19649,N_18162);
or UO_1511 (O_1511,N_17230,N_18363);
xor UO_1512 (O_1512,N_15109,N_18067);
or UO_1513 (O_1513,N_16675,N_17659);
xnor UO_1514 (O_1514,N_16075,N_15906);
nand UO_1515 (O_1515,N_19018,N_18057);
nor UO_1516 (O_1516,N_18740,N_19688);
nand UO_1517 (O_1517,N_19635,N_16094);
or UO_1518 (O_1518,N_17784,N_18563);
and UO_1519 (O_1519,N_16271,N_17599);
xor UO_1520 (O_1520,N_19122,N_17591);
xor UO_1521 (O_1521,N_17921,N_19699);
nor UO_1522 (O_1522,N_19938,N_15029);
or UO_1523 (O_1523,N_16351,N_17875);
nor UO_1524 (O_1524,N_16931,N_16089);
nand UO_1525 (O_1525,N_17450,N_19062);
xor UO_1526 (O_1526,N_16163,N_18349);
and UO_1527 (O_1527,N_15798,N_17457);
or UO_1528 (O_1528,N_15311,N_19116);
and UO_1529 (O_1529,N_16231,N_18685);
xor UO_1530 (O_1530,N_18364,N_18433);
and UO_1531 (O_1531,N_19587,N_17758);
and UO_1532 (O_1532,N_16224,N_17368);
or UO_1533 (O_1533,N_18096,N_15436);
nand UO_1534 (O_1534,N_19817,N_18631);
and UO_1535 (O_1535,N_19013,N_15584);
xnor UO_1536 (O_1536,N_19147,N_15523);
or UO_1537 (O_1537,N_19275,N_19532);
xor UO_1538 (O_1538,N_19875,N_19131);
nor UO_1539 (O_1539,N_18626,N_15955);
xnor UO_1540 (O_1540,N_15588,N_15209);
nand UO_1541 (O_1541,N_19282,N_16552);
xnor UO_1542 (O_1542,N_15901,N_19808);
or UO_1543 (O_1543,N_16260,N_19158);
and UO_1544 (O_1544,N_18284,N_15227);
nand UO_1545 (O_1545,N_15710,N_16760);
nand UO_1546 (O_1546,N_17886,N_15751);
xor UO_1547 (O_1547,N_17717,N_19868);
nand UO_1548 (O_1548,N_17665,N_19290);
or UO_1549 (O_1549,N_17995,N_16334);
xnor UO_1550 (O_1550,N_19783,N_19570);
nand UO_1551 (O_1551,N_16229,N_18393);
xor UO_1552 (O_1552,N_15687,N_19489);
nor UO_1553 (O_1553,N_18152,N_16132);
and UO_1554 (O_1554,N_17068,N_18587);
or UO_1555 (O_1555,N_16576,N_18412);
nand UO_1556 (O_1556,N_16050,N_16593);
xor UO_1557 (O_1557,N_18346,N_19560);
xnor UO_1558 (O_1558,N_19544,N_15389);
nand UO_1559 (O_1559,N_15416,N_16097);
and UO_1560 (O_1560,N_16828,N_17201);
or UO_1561 (O_1561,N_19424,N_16975);
nor UO_1562 (O_1562,N_18125,N_16250);
xnor UO_1563 (O_1563,N_18461,N_18729);
or UO_1564 (O_1564,N_17852,N_17018);
xnor UO_1565 (O_1565,N_16700,N_15920);
or UO_1566 (O_1566,N_17192,N_15467);
nor UO_1567 (O_1567,N_18366,N_19622);
and UO_1568 (O_1568,N_15597,N_16233);
or UO_1569 (O_1569,N_16609,N_19232);
and UO_1570 (O_1570,N_18137,N_15956);
nor UO_1571 (O_1571,N_18530,N_15041);
xor UO_1572 (O_1572,N_18454,N_17788);
nor UO_1573 (O_1573,N_16064,N_17987);
or UO_1574 (O_1574,N_19512,N_18585);
and UO_1575 (O_1575,N_19306,N_15438);
nor UO_1576 (O_1576,N_18900,N_18186);
xor UO_1577 (O_1577,N_17651,N_15131);
nor UO_1578 (O_1578,N_18575,N_16226);
and UO_1579 (O_1579,N_18269,N_15776);
xor UO_1580 (O_1580,N_16512,N_18339);
and UO_1581 (O_1581,N_15353,N_16917);
nand UO_1582 (O_1582,N_19627,N_19227);
nand UO_1583 (O_1583,N_19964,N_15187);
or UO_1584 (O_1584,N_17727,N_16027);
or UO_1585 (O_1585,N_17851,N_15339);
and UO_1586 (O_1586,N_15025,N_17931);
nor UO_1587 (O_1587,N_19655,N_19823);
xnor UO_1588 (O_1588,N_17820,N_15688);
nor UO_1589 (O_1589,N_16346,N_17710);
or UO_1590 (O_1590,N_15815,N_16034);
xnor UO_1591 (O_1591,N_15413,N_17347);
nand UO_1592 (O_1592,N_15730,N_15173);
xor UO_1593 (O_1593,N_15807,N_17267);
or UO_1594 (O_1594,N_17712,N_19262);
nand UO_1595 (O_1595,N_16548,N_15890);
nand UO_1596 (O_1596,N_18836,N_17023);
xor UO_1597 (O_1597,N_17778,N_18081);
xnor UO_1598 (O_1598,N_17516,N_16858);
nor UO_1599 (O_1599,N_16851,N_16752);
nor UO_1600 (O_1600,N_19450,N_18362);
and UO_1601 (O_1601,N_16787,N_17769);
and UO_1602 (O_1602,N_17943,N_17910);
and UO_1603 (O_1603,N_19596,N_19599);
xor UO_1604 (O_1604,N_15022,N_18847);
nand UO_1605 (O_1605,N_18590,N_17976);
nor UO_1606 (O_1606,N_17336,N_15410);
nor UO_1607 (O_1607,N_16954,N_15893);
nand UO_1608 (O_1608,N_18072,N_19204);
xor UO_1609 (O_1609,N_16554,N_15214);
xnor UO_1610 (O_1610,N_19820,N_18123);
nand UO_1611 (O_1611,N_16637,N_18300);
and UO_1612 (O_1612,N_17858,N_18616);
nor UO_1613 (O_1613,N_19590,N_19735);
xor UO_1614 (O_1614,N_19913,N_18917);
xor UO_1615 (O_1615,N_16629,N_16078);
and UO_1616 (O_1616,N_17642,N_18540);
or UO_1617 (O_1617,N_15953,N_15484);
xor UO_1618 (O_1618,N_18479,N_18148);
nand UO_1619 (O_1619,N_15224,N_16688);
xor UO_1620 (O_1620,N_17670,N_19328);
xnor UO_1621 (O_1621,N_15698,N_19209);
xor UO_1622 (O_1622,N_18400,N_15130);
and UO_1623 (O_1623,N_15010,N_19716);
xor UO_1624 (O_1624,N_15626,N_16974);
and UO_1625 (O_1625,N_16493,N_17409);
nor UO_1626 (O_1626,N_16739,N_18969);
and UO_1627 (O_1627,N_17299,N_19991);
and UO_1628 (O_1628,N_18267,N_15138);
xnor UO_1629 (O_1629,N_16689,N_16339);
xnor UO_1630 (O_1630,N_17271,N_18132);
nor UO_1631 (O_1631,N_19981,N_17630);
or UO_1632 (O_1632,N_16891,N_15669);
nand UO_1633 (O_1633,N_15004,N_15088);
or UO_1634 (O_1634,N_18775,N_19873);
and UO_1635 (O_1635,N_19979,N_16419);
and UO_1636 (O_1636,N_19812,N_18624);
nand UO_1637 (O_1637,N_18938,N_16244);
xnor UO_1638 (O_1638,N_16020,N_18795);
or UO_1639 (O_1639,N_15552,N_19403);
or UO_1640 (O_1640,N_16225,N_19181);
nand UO_1641 (O_1641,N_19839,N_15237);
or UO_1642 (O_1642,N_15829,N_19093);
xor UO_1643 (O_1643,N_16463,N_17090);
nand UO_1644 (O_1644,N_15281,N_18167);
and UO_1645 (O_1645,N_19367,N_16870);
xor UO_1646 (O_1646,N_16685,N_15042);
or UO_1647 (O_1647,N_15053,N_18560);
xor UO_1648 (O_1648,N_18182,N_18566);
xnor UO_1649 (O_1649,N_17815,N_17966);
nand UO_1650 (O_1650,N_15854,N_18307);
and UO_1651 (O_1651,N_17610,N_17022);
and UO_1652 (O_1652,N_15810,N_18662);
nand UO_1653 (O_1653,N_19094,N_16364);
or UO_1654 (O_1654,N_19949,N_18507);
nand UO_1655 (O_1655,N_18605,N_18960);
nor UO_1656 (O_1656,N_19404,N_17494);
nor UO_1657 (O_1657,N_18347,N_18806);
nand UO_1658 (O_1658,N_16943,N_17415);
xnor UO_1659 (O_1659,N_19303,N_15631);
nor UO_1660 (O_1660,N_18791,N_17947);
xnor UO_1661 (O_1661,N_15188,N_19047);
xor UO_1662 (O_1662,N_19233,N_19695);
nand UO_1663 (O_1663,N_15619,N_19527);
nand UO_1664 (O_1664,N_19895,N_18027);
nand UO_1665 (O_1665,N_17047,N_16924);
nor UO_1666 (O_1666,N_15425,N_17531);
nand UO_1667 (O_1667,N_18229,N_17541);
xnor UO_1668 (O_1668,N_17401,N_16669);
nor UO_1669 (O_1669,N_18935,N_15572);
and UO_1670 (O_1670,N_16036,N_15442);
and UO_1671 (O_1671,N_17702,N_18998);
xor UO_1672 (O_1672,N_16657,N_18134);
nand UO_1673 (O_1673,N_18301,N_17571);
nor UO_1674 (O_1674,N_19415,N_18425);
and UO_1675 (O_1675,N_17750,N_18589);
nand UO_1676 (O_1676,N_15935,N_18170);
or UO_1677 (O_1677,N_18755,N_16067);
or UO_1678 (O_1678,N_19401,N_19207);
xnor UO_1679 (O_1679,N_15650,N_16261);
and UO_1680 (O_1680,N_18578,N_15709);
or UO_1681 (O_1681,N_16055,N_19300);
or UO_1682 (O_1682,N_17560,N_15848);
nor UO_1683 (O_1683,N_17268,N_19420);
and UO_1684 (O_1684,N_15615,N_19529);
xnor UO_1685 (O_1685,N_16332,N_18389);
or UO_1686 (O_1686,N_17865,N_18435);
or UO_1687 (O_1687,N_16825,N_16202);
nor UO_1688 (O_1688,N_16934,N_15233);
and UO_1689 (O_1689,N_18381,N_19445);
xnor UO_1690 (O_1690,N_16627,N_19480);
and UO_1691 (O_1691,N_17185,N_17140);
and UO_1692 (O_1692,N_19955,N_19455);
and UO_1693 (O_1693,N_17691,N_17116);
nor UO_1694 (O_1694,N_18660,N_17791);
or UO_1695 (O_1695,N_17989,N_16072);
nor UO_1696 (O_1696,N_18309,N_19067);
xnor UO_1697 (O_1697,N_15487,N_17154);
nand UO_1698 (O_1698,N_19281,N_18022);
nand UO_1699 (O_1699,N_16091,N_19882);
and UO_1700 (O_1700,N_17414,N_19516);
xor UO_1701 (O_1701,N_19911,N_19370);
xor UO_1702 (O_1702,N_18149,N_17949);
nor UO_1703 (O_1703,N_15638,N_17962);
or UO_1704 (O_1704,N_16678,N_19908);
nor UO_1705 (O_1705,N_17071,N_15623);
nor UO_1706 (O_1706,N_15343,N_19176);
nor UO_1707 (O_1707,N_19629,N_16022);
or UO_1708 (O_1708,N_16973,N_19523);
nor UO_1709 (O_1709,N_17237,N_15056);
and UO_1710 (O_1710,N_17037,N_15696);
xnor UO_1711 (O_1711,N_15500,N_19681);
nand UO_1712 (O_1712,N_16838,N_18889);
or UO_1713 (O_1713,N_15717,N_17451);
nor UO_1714 (O_1714,N_19732,N_16985);
nor UO_1715 (O_1715,N_19296,N_19931);
or UO_1716 (O_1716,N_16276,N_18466);
nor UO_1717 (O_1717,N_16348,N_19387);
xnor UO_1718 (O_1718,N_18156,N_15985);
nand UO_1719 (O_1719,N_18494,N_19602);
and UO_1720 (O_1720,N_19085,N_18449);
nand UO_1721 (O_1721,N_19852,N_19273);
nand UO_1722 (O_1722,N_19582,N_18519);
and UO_1723 (O_1723,N_19835,N_19452);
xnor UO_1724 (O_1724,N_17266,N_16731);
nand UO_1725 (O_1725,N_18041,N_15789);
nand UO_1726 (O_1726,N_16905,N_15781);
xor UO_1727 (O_1727,N_17706,N_17552);
nand UO_1728 (O_1728,N_16578,N_16803);
nand UO_1729 (O_1729,N_15080,N_15871);
or UO_1730 (O_1730,N_19329,N_17690);
or UO_1731 (O_1731,N_19435,N_17136);
or UO_1732 (O_1732,N_16358,N_17800);
xnor UO_1733 (O_1733,N_19379,N_17096);
nor UO_1734 (O_1734,N_16182,N_17274);
and UO_1735 (O_1735,N_19111,N_16951);
and UO_1736 (O_1736,N_18782,N_16205);
nor UO_1737 (O_1737,N_15758,N_19351);
nand UO_1738 (O_1738,N_19330,N_16521);
nand UO_1739 (O_1739,N_15714,N_19238);
xnor UO_1740 (O_1740,N_18904,N_15937);
nand UO_1741 (O_1741,N_17213,N_16307);
or UO_1742 (O_1742,N_15590,N_16878);
and UO_1743 (O_1743,N_19883,N_19617);
and UO_1744 (O_1744,N_16217,N_19604);
and UO_1745 (O_1745,N_19241,N_15431);
or UO_1746 (O_1746,N_19597,N_18841);
nand UO_1747 (O_1747,N_18899,N_15697);
nand UO_1748 (O_1748,N_15559,N_18405);
xor UO_1749 (O_1749,N_16729,N_15015);
xnor UO_1750 (O_1750,N_17740,N_15827);
or UO_1751 (O_1751,N_16634,N_15072);
xnor UO_1752 (O_1752,N_17609,N_18100);
nor UO_1753 (O_1753,N_16531,N_18629);
nor UO_1754 (O_1754,N_16349,N_16775);
or UO_1755 (O_1755,N_16555,N_19877);
and UO_1756 (O_1756,N_18496,N_19051);
nor UO_1757 (O_1757,N_18194,N_16823);
and UO_1758 (O_1758,N_19448,N_15511);
nand UO_1759 (O_1759,N_18848,N_15445);
nand UO_1760 (O_1760,N_18255,N_18473);
nor UO_1761 (O_1761,N_15000,N_16423);
or UO_1762 (O_1762,N_18486,N_18647);
or UO_1763 (O_1763,N_19123,N_16499);
nand UO_1764 (O_1764,N_19441,N_15888);
xor UO_1765 (O_1765,N_19513,N_18146);
and UO_1766 (O_1766,N_17221,N_19997);
nor UO_1767 (O_1767,N_16297,N_18837);
nor UO_1768 (O_1768,N_17471,N_15264);
or UO_1769 (O_1769,N_19199,N_17387);
nand UO_1770 (O_1770,N_19543,N_17619);
nor UO_1771 (O_1771,N_15102,N_19477);
nand UO_1772 (O_1772,N_18280,N_19841);
xor UO_1773 (O_1773,N_17960,N_19134);
nor UO_1774 (O_1774,N_19203,N_17055);
or UO_1775 (O_1775,N_17317,N_19072);
and UO_1776 (O_1776,N_16788,N_17834);
xor UO_1777 (O_1777,N_19070,N_16486);
nor UO_1778 (O_1778,N_19291,N_16772);
nand UO_1779 (O_1779,N_15319,N_18823);
and UO_1780 (O_1780,N_19107,N_18509);
xnor UO_1781 (O_1781,N_19522,N_19721);
nand UO_1782 (O_1782,N_16867,N_17015);
or UO_1783 (O_1783,N_16234,N_18982);
or UO_1784 (O_1784,N_16090,N_15230);
nand UO_1785 (O_1785,N_16514,N_16916);
xor UO_1786 (O_1786,N_16479,N_16135);
nor UO_1787 (O_1787,N_15231,N_19631);
nor UO_1788 (O_1788,N_15177,N_15910);
or UO_1789 (O_1789,N_17419,N_17983);
and UO_1790 (O_1790,N_19885,N_15573);
nand UO_1791 (O_1791,N_18453,N_19187);
nand UO_1792 (O_1792,N_17160,N_19665);
xnor UO_1793 (O_1793,N_16842,N_16881);
xnor UO_1794 (O_1794,N_17749,N_17918);
or UO_1795 (O_1795,N_17331,N_16728);
or UO_1796 (O_1796,N_17010,N_18556);
and UO_1797 (O_1797,N_19707,N_16519);
nand UO_1798 (O_1798,N_15783,N_19977);
nor UO_1799 (O_1799,N_17087,N_18184);
or UO_1800 (O_1800,N_19201,N_17942);
xnor UO_1801 (O_1801,N_15958,N_18117);
xor UO_1802 (O_1802,N_15217,N_18720);
xor UO_1803 (O_1803,N_19459,N_16500);
nand UO_1804 (O_1804,N_16208,N_18752);
xor UO_1805 (O_1805,N_19393,N_19044);
and UO_1806 (O_1806,N_17344,N_17627);
xnor UO_1807 (O_1807,N_16583,N_19921);
or UO_1808 (O_1808,N_17873,N_15647);
xor UO_1809 (O_1809,N_16359,N_18541);
nand UO_1810 (O_1810,N_18279,N_16134);
nand UO_1811 (O_1811,N_16602,N_17669);
nand UO_1812 (O_1812,N_15860,N_16995);
or UO_1813 (O_1813,N_16699,N_19899);
and UO_1814 (O_1814,N_15961,N_19271);
and UO_1815 (O_1815,N_18741,N_16762);
or UO_1816 (O_1816,N_18682,N_15671);
nor UO_1817 (O_1817,N_16737,N_16747);
xnor UO_1818 (O_1818,N_19738,N_18692);
nor UO_1819 (O_1819,N_17156,N_19320);
xnor UO_1820 (O_1820,N_19025,N_16071);
nor UO_1821 (O_1821,N_17195,N_19228);
xor UO_1822 (O_1822,N_16890,N_17310);
nor UO_1823 (O_1823,N_15843,N_15865);
nand UO_1824 (O_1824,N_19772,N_16776);
nor UO_1825 (O_1825,N_19150,N_17246);
nor UO_1826 (O_1826,N_16961,N_17509);
and UO_1827 (O_1827,N_18637,N_15397);
nand UO_1828 (O_1828,N_16383,N_19165);
nor UO_1829 (O_1829,N_15814,N_15073);
nand UO_1830 (O_1830,N_16092,N_19989);
xor UO_1831 (O_1831,N_19603,N_19634);
and UO_1832 (O_1832,N_16005,N_15186);
nor UO_1833 (O_1833,N_19461,N_17427);
and UO_1834 (O_1834,N_15856,N_15875);
xor UO_1835 (O_1835,N_18223,N_16015);
or UO_1836 (O_1836,N_19319,N_17998);
or UO_1837 (O_1837,N_17340,N_15867);
or UO_1838 (O_1838,N_15409,N_19640);
nor UO_1839 (O_1839,N_19791,N_17456);
and UO_1840 (O_1840,N_16176,N_16898);
and UO_1841 (O_1841,N_18968,N_19647);
xnor UO_1842 (O_1842,N_15981,N_17469);
xnor UO_1843 (O_1843,N_19573,N_16709);
nand UO_1844 (O_1844,N_18427,N_16714);
and UO_1845 (O_1845,N_19342,N_17329);
nor UO_1846 (O_1846,N_19120,N_18238);
or UO_1847 (O_1847,N_15008,N_19210);
xnor UO_1848 (O_1848,N_16735,N_15383);
xnor UO_1849 (O_1849,N_16414,N_16282);
xnor UO_1850 (O_1850,N_16184,N_18814);
nand UO_1851 (O_1851,N_17618,N_18551);
xnor UO_1852 (O_1852,N_18438,N_15943);
or UO_1853 (O_1853,N_17101,N_18213);
or UO_1854 (O_1854,N_17508,N_16187);
xor UO_1855 (O_1855,N_16756,N_18784);
nor UO_1856 (O_1856,N_18546,N_18391);
or UO_1857 (O_1857,N_17585,N_18618);
and UO_1858 (O_1858,N_16327,N_19497);
nor UO_1859 (O_1859,N_17996,N_18664);
or UO_1860 (O_1860,N_16249,N_18804);
or UO_1861 (O_1861,N_19770,N_16006);
and UO_1862 (O_1862,N_19440,N_15229);
and UO_1863 (O_1863,N_18119,N_18059);
and UO_1864 (O_1864,N_15387,N_15822);
and UO_1865 (O_1865,N_17564,N_18643);
or UO_1866 (O_1866,N_17793,N_19915);
nand UO_1867 (O_1867,N_16453,N_18671);
nand UO_1868 (O_1868,N_18691,N_16291);
nand UO_1869 (O_1869,N_17361,N_19006);
nor UO_1870 (O_1870,N_15600,N_15119);
and UO_1871 (O_1871,N_19754,N_15295);
or UO_1872 (O_1872,N_16107,N_16622);
or UO_1873 (O_1873,N_18128,N_17332);
xnor UO_1874 (O_1874,N_19360,N_17801);
nor UO_1875 (O_1875,N_18332,N_16478);
and UO_1876 (O_1876,N_18650,N_17772);
xnor UO_1877 (O_1877,N_17961,N_16989);
and UO_1878 (O_1878,N_17663,N_15244);
and UO_1879 (O_1879,N_16536,N_16025);
nor UO_1880 (O_1880,N_19859,N_16149);
or UO_1881 (O_1881,N_19551,N_15360);
xnor UO_1882 (O_1882,N_15185,N_16472);
nand UO_1883 (O_1883,N_18215,N_18562);
xor UO_1884 (O_1884,N_18656,N_18112);
and UO_1885 (O_1885,N_17889,N_19887);
nand UO_1886 (O_1886,N_16230,N_15739);
nand UO_1887 (O_1887,N_19642,N_18180);
nor UO_1888 (O_1888,N_15764,N_18439);
nand UO_1889 (O_1889,N_19285,N_19967);
nor UO_1890 (O_1890,N_16392,N_19079);
xor UO_1891 (O_1891,N_19518,N_17005);
xor UO_1892 (O_1892,N_15659,N_17540);
or UO_1893 (O_1893,N_18973,N_18539);
nand UO_1894 (O_1894,N_18116,N_18996);
nor UO_1895 (O_1895,N_16388,N_18828);
nand UO_1896 (O_1896,N_16177,N_15009);
nand UO_1897 (O_1897,N_17576,N_19463);
or UO_1898 (O_1898,N_18345,N_19692);
xor UO_1899 (O_1899,N_19425,N_18079);
or UO_1900 (O_1900,N_19553,N_15247);
or UO_1901 (O_1901,N_19105,N_17301);
and UO_1902 (O_1902,N_15548,N_18154);
xnor UO_1903 (O_1903,N_19723,N_19208);
nor UO_1904 (O_1904,N_18145,N_15909);
and UO_1905 (O_1905,N_18856,N_18654);
nand UO_1906 (O_1906,N_19985,N_18244);
and UO_1907 (O_1907,N_15402,N_15309);
nand UO_1908 (O_1908,N_16035,N_16368);
nor UO_1909 (O_1909,N_15367,N_15889);
or UO_1910 (O_1910,N_16569,N_17893);
and UO_1911 (O_1911,N_16810,N_16079);
xnor UO_1912 (O_1912,N_16046,N_15357);
nand UO_1913 (O_1913,N_15429,N_19889);
xor UO_1914 (O_1914,N_18350,N_19524);
or UO_1915 (O_1915,N_15825,N_17109);
xnor UO_1916 (O_1916,N_16343,N_17502);
or UO_1917 (O_1917,N_16529,N_18025);
nor UO_1918 (O_1918,N_15122,N_17797);
or UO_1919 (O_1919,N_15857,N_19935);
or UO_1920 (O_1920,N_17580,N_19626);
nor UO_1921 (O_1921,N_18564,N_16730);
nor UO_1922 (O_1922,N_15532,N_15804);
nor UO_1923 (O_1923,N_17137,N_17048);
nand UO_1924 (O_1924,N_18331,N_15649);
or UO_1925 (O_1925,N_17288,N_19447);
nor UO_1926 (O_1926,N_18390,N_16549);
and UO_1927 (O_1927,N_17501,N_18160);
xnor UO_1928 (O_1928,N_15991,N_19585);
xnor UO_1929 (O_1929,N_16120,N_18263);
and UO_1930 (O_1930,N_16935,N_17624);
and UO_1931 (O_1931,N_18850,N_17108);
or UO_1932 (O_1932,N_16382,N_16369);
or UO_1933 (O_1933,N_16702,N_15288);
nor UO_1934 (O_1934,N_16876,N_19517);
nand UO_1935 (O_1935,N_17094,N_15501);
and UO_1936 (O_1936,N_16636,N_16502);
xnor UO_1937 (O_1937,N_17375,N_16319);
and UO_1938 (O_1938,N_16603,N_16904);
xor UO_1939 (O_1939,N_17104,N_18813);
nor UO_1940 (O_1940,N_19661,N_15470);
nand UO_1941 (O_1941,N_19966,N_15205);
and UO_1942 (O_1942,N_17980,N_18423);
nor UO_1943 (O_1943,N_16732,N_16666);
xor UO_1944 (O_1944,N_15336,N_15914);
xnor UO_1945 (O_1945,N_15661,N_15441);
nor UO_1946 (O_1946,N_16518,N_16357);
nor UO_1947 (O_1947,N_18779,N_19763);
nand UO_1948 (O_1948,N_18533,N_15396);
and UO_1949 (O_1949,N_19305,N_17513);
nor UO_1950 (O_1950,N_15359,N_17406);
nand UO_1951 (O_1951,N_18085,N_15967);
nor UO_1952 (O_1952,N_18789,N_16997);
nor UO_1953 (O_1953,N_17319,N_19478);
nand UO_1954 (O_1954,N_17430,N_18997);
nand UO_1955 (O_1955,N_17367,N_15613);
xor UO_1956 (O_1956,N_18260,N_15837);
or UO_1957 (O_1957,N_17787,N_15422);
nor UO_1958 (O_1958,N_18607,N_16644);
and UO_1959 (O_1959,N_17420,N_15508);
nor UO_1960 (O_1960,N_17964,N_19143);
nor UO_1961 (O_1961,N_16648,N_19456);
nand UO_1962 (O_1962,N_15561,N_16649);
nor UO_1963 (O_1963,N_15475,N_17885);
nand UO_1964 (O_1964,N_17265,N_18698);
and UO_1965 (O_1965,N_16443,N_18388);
nor UO_1966 (O_1966,N_15078,N_19767);
xor UO_1967 (O_1967,N_15381,N_16488);
xor UO_1968 (O_1968,N_16960,N_17718);
and UO_1969 (O_1969,N_18924,N_15706);
or UO_1970 (O_1970,N_17006,N_19850);
or UO_1971 (O_1971,N_15668,N_18264);
xnor UO_1972 (O_1972,N_18477,N_19372);
xor UO_1973 (O_1973,N_16511,N_16302);
nor UO_1974 (O_1974,N_17832,N_17647);
or UO_1975 (O_1975,N_17491,N_16321);
xor UO_1976 (O_1976,N_15239,N_18501);
nor UO_1977 (O_1977,N_18955,N_17098);
or UO_1978 (O_1978,N_15818,N_16534);
xnor UO_1979 (O_1979,N_18657,N_18920);
xnor UO_1980 (O_1980,N_15127,N_17240);
nand UO_1981 (O_1981,N_16790,N_19283);
xor UO_1982 (O_1982,N_19843,N_18834);
nor UO_1983 (O_1983,N_18534,N_16185);
nor UO_1984 (O_1984,N_19230,N_17922);
nand UO_1985 (O_1985,N_16715,N_19083);
or UO_1986 (O_1986,N_15621,N_18036);
nor UO_1987 (O_1987,N_19011,N_19802);
or UO_1988 (O_1988,N_15823,N_17276);
nor UO_1989 (O_1989,N_19620,N_15274);
and UO_1990 (O_1990,N_18620,N_17454);
xnor UO_1991 (O_1991,N_15310,N_17664);
and UO_1992 (O_1992,N_17210,N_17574);
and UO_1993 (O_1993,N_19405,N_16492);
nand UO_1994 (O_1994,N_19719,N_16996);
or UO_1995 (O_1995,N_19173,N_15284);
or UO_1996 (O_1996,N_15907,N_18926);
nor UO_1997 (O_1997,N_15401,N_17934);
nand UO_1998 (O_1998,N_18993,N_19392);
or UO_1999 (O_1999,N_18047,N_16240);
and UO_2000 (O_2000,N_15884,N_15035);
and UO_2001 (O_2001,N_18235,N_15792);
nor UO_2002 (O_2002,N_15469,N_17954);
nand UO_2003 (O_2003,N_16192,N_18816);
or UO_2004 (O_2004,N_18183,N_15530);
nor UO_2005 (O_2005,N_19509,N_18915);
nand UO_2006 (O_2006,N_18762,N_19779);
nand UO_2007 (O_2007,N_16300,N_15740);
nand UO_2008 (O_2008,N_15578,N_19137);
nor UO_2009 (O_2009,N_18723,N_15451);
and UO_2010 (O_2010,N_19795,N_19074);
xnor UO_2011 (O_2011,N_17726,N_19154);
and UO_2012 (O_2012,N_16341,N_15051);
or UO_2013 (O_2013,N_19189,N_18537);
nor UO_2014 (O_2014,N_16337,N_15546);
nand UO_2015 (O_2015,N_17882,N_19945);
nand UO_2016 (O_2016,N_18705,N_17900);
nor UO_2017 (O_2017,N_17923,N_15852);
nand UO_2018 (O_2018,N_17366,N_19556);
xnor UO_2019 (O_2019,N_19799,N_16275);
nor UO_2020 (O_2020,N_17223,N_17488);
and UO_2021 (O_2021,N_15587,N_19671);
nand UO_2022 (O_2022,N_16069,N_19057);
nand UO_2023 (O_2023,N_17661,N_16345);
nor UO_2024 (O_2024,N_17260,N_15236);
nand UO_2025 (O_2025,N_17803,N_16862);
nor UO_2026 (O_2026,N_16294,N_18876);
xor UO_2027 (O_2027,N_17756,N_19108);
nand UO_2028 (O_2028,N_16197,N_18294);
or UO_2029 (O_2029,N_19383,N_16835);
nor UO_2030 (O_2030,N_18108,N_17421);
and UO_2031 (O_2031,N_17345,N_15718);
nor UO_2032 (O_2032,N_16384,N_15419);
nor UO_2033 (O_2033,N_17988,N_16175);
or UO_2034 (O_2034,N_19538,N_15439);
or UO_2035 (O_2035,N_16826,N_17662);
or UO_2036 (O_2036,N_18107,N_16085);
and UO_2037 (O_2037,N_19464,N_15071);
nor UO_2038 (O_2038,N_18668,N_15415);
nand UO_2039 (O_2039,N_18432,N_16270);
nor UO_2040 (O_2040,N_18413,N_19126);
xnor UO_2041 (O_2041,N_17866,N_17759);
xnor UO_2042 (O_2042,N_16042,N_18630);
xor UO_2043 (O_2043,N_19746,N_17144);
and UO_2044 (O_2044,N_17628,N_19510);
nor UO_2045 (O_2045,N_17490,N_15555);
nor UO_2046 (O_2046,N_18039,N_15633);
xnor UO_2047 (O_2047,N_15322,N_19288);
xor UO_2048 (O_2048,N_18777,N_18812);
or UO_2049 (O_2049,N_15043,N_16387);
and UO_2050 (O_2050,N_15646,N_15965);
or UO_2051 (O_2051,N_15167,N_19612);
or UO_2052 (O_2052,N_16630,N_17275);
nor UO_2053 (O_2053,N_19580,N_19525);
and UO_2054 (O_2054,N_15366,N_16767);
and UO_2055 (O_2055,N_16882,N_19774);
or UO_2056 (O_2056,N_16206,N_19969);
nor UO_2057 (O_2057,N_15754,N_16566);
nor UO_2058 (O_2058,N_18649,N_17452);
or UO_2059 (O_2059,N_16378,N_15161);
or UO_2060 (O_2060,N_15318,N_16060);
nand UO_2061 (O_2061,N_18463,N_17631);
xnor UO_2062 (O_2062,N_16475,N_19605);
xnor UO_2063 (O_2063,N_15443,N_18884);
and UO_2064 (O_2064,N_17016,N_19161);
nor UO_2065 (O_2065,N_19251,N_19114);
xor UO_2066 (O_2066,N_16620,N_16130);
nand UO_2067 (O_2067,N_18978,N_18712);
nor UO_2068 (O_2068,N_15757,N_15046);
and UO_2069 (O_2069,N_16039,N_19045);
and UO_2070 (O_2070,N_16719,N_15065);
or UO_2071 (O_2071,N_16804,N_19737);
nand UO_2072 (O_2072,N_19571,N_18853);
nor UO_2073 (O_2073,N_18877,N_15773);
or UO_2074 (O_2074,N_17826,N_17746);
nor UO_2075 (O_2075,N_19391,N_16180);
nand UO_2076 (O_2076,N_16178,N_16970);
or UO_2077 (O_2077,N_15124,N_15581);
or UO_2078 (O_2078,N_15734,N_17573);
or UO_2079 (O_2079,N_18061,N_15874);
and UO_2080 (O_2080,N_16084,N_15960);
nand UO_2081 (O_2081,N_15298,N_18604);
nor UO_2082 (O_2082,N_15068,N_16361);
nor UO_2083 (O_2083,N_15931,N_18710);
nor UO_2084 (O_2084,N_17556,N_15235);
and UO_2085 (O_2085,N_15805,N_17432);
or UO_2086 (O_2086,N_19986,N_18322);
nand UO_2087 (O_2087,N_19317,N_15731);
xor UO_2088 (O_2088,N_19487,N_15203);
nand UO_2089 (O_2089,N_16921,N_15767);
and UO_2090 (O_2090,N_15622,N_17722);
or UO_2091 (O_2091,N_15001,N_15950);
nor UO_2092 (O_2092,N_15895,N_19546);
nor UO_2093 (O_2093,N_17829,N_16429);
or UO_2094 (O_2094,N_15514,N_18404);
nor UO_2095 (O_2095,N_16190,N_15250);
xnor UO_2096 (O_2096,N_15062,N_16741);
and UO_2097 (O_2097,N_16150,N_17194);
nand UO_2098 (O_2098,N_16056,N_17342);
nand UO_2099 (O_2099,N_15545,N_16801);
and UO_2100 (O_2100,N_17295,N_19789);
and UO_2101 (O_2101,N_16926,N_18054);
and UO_2102 (O_2102,N_18212,N_17142);
nor UO_2103 (O_2103,N_18325,N_19569);
and UO_2104 (O_2104,N_17752,N_18763);
nand UO_2105 (O_2105,N_15790,N_18076);
nand UO_2106 (O_2106,N_16274,N_17824);
and UO_2107 (O_2107,N_16051,N_19005);
or UO_2108 (O_2108,N_19630,N_19658);
xnor UO_2109 (O_2109,N_17382,N_16430);
and UO_2110 (O_2110,N_15196,N_15853);
or UO_2111 (O_2111,N_15694,N_19520);
nor UO_2112 (O_2112,N_15493,N_15979);
and UO_2113 (O_2113,N_17880,N_16541);
nor UO_2114 (O_2114,N_16551,N_17567);
nand UO_2115 (O_2115,N_17897,N_17333);
nor UO_2116 (O_2116,N_15246,N_18508);
and UO_2117 (O_2117,N_17483,N_18018);
nand UO_2118 (O_2118,N_15813,N_19010);
xor UO_2119 (O_2119,N_15113,N_19234);
nand UO_2120 (O_2120,N_15978,N_15542);
nor UO_2121 (O_2121,N_16967,N_17802);
or UO_2122 (O_2122,N_19397,N_18683);
xnor UO_2123 (O_2123,N_17172,N_15117);
nand UO_2124 (O_2124,N_17871,N_15877);
nor UO_2125 (O_2125,N_15727,N_15519);
nor UO_2126 (O_2126,N_17081,N_18086);
or UO_2127 (O_2127,N_18351,N_18634);
xnor UO_2128 (O_2128,N_16155,N_19948);
nor UO_2129 (O_2129,N_17428,N_18897);
xor UO_2130 (O_2130,N_17657,N_19710);
and UO_2131 (O_2131,N_17167,N_16258);
or UO_2132 (O_2132,N_16309,N_17558);
nor UO_2133 (O_2133,N_15182,N_16464);
and UO_2134 (O_2134,N_17920,N_17306);
or UO_2135 (O_2135,N_18995,N_16485);
and UO_2136 (O_2136,N_19412,N_17362);
xnor UO_2137 (O_2137,N_15828,N_17384);
nor UO_2138 (O_2138,N_17589,N_17350);
or UO_2139 (O_2139,N_18121,N_19494);
nand UO_2140 (O_2140,N_16588,N_17916);
or UO_2141 (O_2141,N_16830,N_18490);
and UO_2142 (O_2142,N_15018,N_18241);
and UO_2143 (O_2143,N_19600,N_17542);
or UO_2144 (O_2144,N_16856,N_18768);
nand UO_2145 (O_2145,N_15204,N_19624);
or UO_2146 (O_2146,N_19936,N_18518);
nand UO_2147 (O_2147,N_19691,N_19343);
or UO_2148 (O_2148,N_16816,N_15691);
xor UO_2149 (O_2149,N_15655,N_17397);
nand UO_2150 (O_2150,N_16403,N_18492);
nand UO_2151 (O_2151,N_15689,N_17150);
and UO_2152 (O_2152,N_15039,N_17416);
nand UO_2153 (O_2153,N_18588,N_18547);
nor UO_2154 (O_2154,N_17990,N_19188);
xnor UO_2155 (O_2155,N_17065,N_17679);
nand UO_2156 (O_2156,N_16376,N_15462);
xnor UO_2157 (O_2157,N_18040,N_15641);
and UO_2158 (O_2158,N_18957,N_16723);
or UO_2159 (O_2159,N_19793,N_17506);
xnor UO_2160 (O_2160,N_17289,N_18384);
nand UO_2161 (O_2161,N_18283,N_19806);
nor UO_2162 (O_2162,N_16956,N_17217);
or UO_2163 (O_2163,N_15306,N_15547);
xor UO_2164 (O_2164,N_17993,N_15014);
and UO_2165 (O_2165,N_18299,N_16864);
nor UO_2166 (O_2166,N_19023,N_18017);
nand UO_2167 (O_2167,N_15930,N_17548);
or UO_2168 (O_2168,N_17264,N_15700);
nand UO_2169 (O_2169,N_16690,N_16081);
or UO_2170 (O_2170,N_16906,N_17731);
xor UO_2171 (O_2171,N_15780,N_19499);
xnor UO_2172 (O_2172,N_18908,N_19809);
nor UO_2173 (O_2173,N_19248,N_19548);
and UO_2174 (O_2174,N_17856,N_16980);
nor UO_2175 (O_2175,N_16269,N_19521);
nor UO_2176 (O_2176,N_15785,N_19844);
nor UO_2177 (O_2177,N_16713,N_18725);
or UO_2178 (O_2178,N_16145,N_16405);
xor UO_2179 (O_2179,N_19628,N_16668);
xor UO_2180 (O_2180,N_15941,N_16484);
or UO_2181 (O_2181,N_15299,N_19321);
nand UO_2182 (O_2182,N_17695,N_19720);
or UO_2183 (O_2183,N_16393,N_16670);
xnor UO_2184 (O_2184,N_18060,N_17429);
xnor UO_2185 (O_2185,N_15120,N_19476);
and UO_2186 (O_2186,N_17007,N_17102);
nand UO_2187 (O_2187,N_17835,N_19078);
nor UO_2188 (O_2188,N_19144,N_16783);
xnor UO_2189 (O_2189,N_17351,N_16619);
nor UO_2190 (O_2190,N_16909,N_17476);
or UO_2191 (O_2191,N_19353,N_16287);
nand UO_2192 (O_2192,N_18460,N_19703);
nand UO_2193 (O_2193,N_15713,N_15377);
xor UO_2194 (O_2194,N_19729,N_18721);
nor UO_2195 (O_2195,N_18928,N_15596);
nor UO_2196 (O_2196,N_17909,N_18695);
or UO_2197 (O_2197,N_18476,N_17681);
nand UO_2198 (O_2198,N_15995,N_17180);
or UO_2199 (O_2199,N_18444,N_18204);
or UO_2200 (O_2200,N_18348,N_19245);
or UO_2201 (O_2201,N_18201,N_19540);
xnor UO_2202 (O_2202,N_16998,N_15786);
or UO_2203 (O_2203,N_19923,N_16424);
nand UO_2204 (O_2204,N_19562,N_17860);
nor UO_2205 (O_2205,N_17945,N_18581);
xnor UO_2206 (O_2206,N_17538,N_17353);
xnor UO_2207 (O_2207,N_19418,N_17958);
nand UO_2208 (O_2208,N_19528,N_17760);
nor UO_2209 (O_2209,N_17809,N_18153);
or UO_2210 (O_2210,N_15949,N_17040);
nor UO_2211 (O_2211,N_17956,N_18869);
xor UO_2212 (O_2212,N_19263,N_15738);
or UO_2213 (O_2213,N_15070,N_16471);
nor UO_2214 (O_2214,N_18862,N_16530);
and UO_2215 (O_2215,N_15632,N_17008);
xor UO_2216 (O_2216,N_18864,N_16792);
xnor UO_2217 (O_2217,N_15498,N_18320);
and UO_2218 (O_2218,N_18661,N_15040);
and UO_2219 (O_2219,N_17725,N_18087);
and UO_2220 (O_2220,N_17781,N_16059);
nor UO_2221 (O_2221,N_19787,N_15355);
or UO_2222 (O_2222,N_17652,N_19400);
nand UO_2223 (O_2223,N_15526,N_18987);
xnor UO_2224 (O_2224,N_17422,N_18293);
nor UO_2225 (O_2225,N_15654,N_15996);
xnor UO_2226 (O_2226,N_15254,N_18024);
xnor UO_2227 (O_2227,N_17398,N_16389);
or UO_2228 (O_2228,N_17261,N_15509);
xnor UO_2229 (O_2229,N_17892,N_19614);
and UO_2230 (O_2230,N_15863,N_15471);
and UO_2231 (O_2231,N_16535,N_17607);
or UO_2232 (O_2232,N_19020,N_17570);
nor UO_2233 (O_2233,N_18098,N_19421);
and UO_2234 (O_2234,N_16460,N_19766);
and UO_2235 (O_2235,N_16273,N_16791);
or UO_2236 (O_2236,N_16450,N_17381);
nand UO_2237 (O_2237,N_16350,N_18674);
nand UO_2238 (O_2238,N_17356,N_18074);
xnor UO_2239 (O_2239,N_19801,N_16420);
nor UO_2240 (O_2240,N_15446,N_15238);
xor UO_2241 (O_2241,N_17470,N_15882);
nor UO_2242 (O_2242,N_18317,N_16119);
or UO_2243 (O_2243,N_19554,N_16533);
and UO_2244 (O_2244,N_17840,N_15775);
or UO_2245 (O_2245,N_17139,N_15333);
xor UO_2246 (O_2246,N_15984,N_19414);
nand UO_2247 (O_2247,N_18835,N_18941);
xor UO_2248 (O_2248,N_19388,N_19891);
nor UO_2249 (O_2249,N_15275,N_19901);
nand UO_2250 (O_2250,N_15574,N_17115);
nor UO_2251 (O_2251,N_19386,N_15932);
or UO_2252 (O_2252,N_16065,N_19943);
or UO_2253 (O_2253,N_18451,N_17304);
nor UO_2254 (O_2254,N_17009,N_19075);
or UO_2255 (O_2255,N_16976,N_15420);
nand UO_2256 (O_2256,N_18861,N_18617);
and UO_2257 (O_2257,N_15325,N_16919);
nor UO_2258 (O_2258,N_17001,N_17935);
nor UO_2259 (O_2259,N_16077,N_19268);
nor UO_2260 (O_2260,N_19743,N_15968);
xnor UO_2261 (O_2261,N_16241,N_15145);
xor UO_2262 (O_2262,N_18343,N_18612);
or UO_2263 (O_2263,N_17955,N_17520);
nand UO_2264 (O_2264,N_17468,N_17149);
or UO_2265 (O_2265,N_19163,N_17925);
nand UO_2266 (O_2266,N_17953,N_16026);
nor UO_2267 (O_2267,N_16927,N_18827);
nand UO_2268 (O_2268,N_17648,N_17219);
or UO_2269 (O_2269,N_16952,N_17963);
or UO_2270 (O_2270,N_17929,N_19952);
or UO_2271 (O_2271,N_17216,N_15086);
or UO_2272 (O_2272,N_16759,N_16793);
nor UO_2273 (O_2273,N_16818,N_19314);
nor UO_2274 (O_2274,N_19975,N_17003);
xnor UO_2275 (O_2275,N_15368,N_19292);
or UO_2276 (O_2276,N_17067,N_17300);
nor UO_2277 (O_2277,N_19162,N_15614);
and UO_2278 (O_2278,N_19395,N_19781);
and UO_2279 (O_2279,N_18972,N_17518);
xor UO_2280 (O_2280,N_19286,N_16279);
or UO_2281 (O_2281,N_17072,N_17859);
nand UO_2282 (O_2282,N_18020,N_17536);
or UO_2283 (O_2283,N_15052,N_18826);
or UO_2284 (O_2284,N_19890,N_17025);
nor UO_2285 (O_2285,N_16695,N_16888);
nor UO_2286 (O_2286,N_16330,N_16542);
and UO_2287 (O_2287,N_19633,N_15414);
nor UO_2288 (O_2288,N_18943,N_15013);
nand UO_2289 (O_2289,N_16083,N_16214);
and UO_2290 (O_2290,N_17635,N_19825);
nand UO_2291 (O_2291,N_19084,N_15448);
xor UO_2292 (O_2292,N_19223,N_16587);
nor UO_2293 (O_2293,N_16754,N_19308);
nand UO_2294 (O_2294,N_16859,N_16480);
nor UO_2295 (O_2295,N_17563,N_15625);
or UO_2296 (O_2296,N_19139,N_18080);
nand UO_2297 (O_2297,N_17281,N_15083);
nor UO_2298 (O_2298,N_16315,N_19648);
and UO_2299 (O_2299,N_19298,N_19535);
nand UO_2300 (O_2300,N_19730,N_18639);
xor UO_2301 (O_2301,N_15933,N_19352);
nand UO_2302 (O_2302,N_16347,N_16218);
nand UO_2303 (O_2303,N_15502,N_16352);
nor UO_2304 (O_2304,N_18354,N_17755);
nand UO_2305 (O_2305,N_17862,N_17286);
xor UO_2306 (O_2306,N_17863,N_16865);
nand UO_2307 (O_2307,N_17492,N_18421);
xor UO_2308 (O_2308,N_16452,N_19259);
nand UO_2309 (O_2309,N_16765,N_16223);
nand UO_2310 (O_2310,N_18700,N_16537);
or UO_2311 (O_2311,N_15106,N_17176);
nand UO_2312 (O_2312,N_15330,N_18724);
or UO_2313 (O_2313,N_18672,N_18846);
nand UO_2314 (O_2314,N_15478,N_16220);
nand UO_2315 (O_2315,N_18314,N_19096);
nor UO_2316 (O_2316,N_17339,N_15795);
nand UO_2317 (O_2317,N_19346,N_15261);
or UO_2318 (O_2318,N_17050,N_16968);
nor UO_2319 (O_2319,N_19133,N_15844);
or UO_2320 (O_2320,N_18273,N_17503);
and UO_2321 (O_2321,N_18945,N_16962);
nor UO_2322 (O_2322,N_19740,N_19242);
and UO_2323 (O_2323,N_15957,N_15105);
nand UO_2324 (O_2324,N_19867,N_16850);
xnor UO_2325 (O_2325,N_19307,N_19169);
or UO_2326 (O_2326,N_19384,N_17046);
nand UO_2327 (O_2327,N_17765,N_18415);
or UO_2328 (O_2328,N_15983,N_16977);
and UO_2329 (O_2329,N_15922,N_17768);
nand UO_2330 (O_2330,N_18580,N_15741);
nand UO_2331 (O_2331,N_19394,N_18918);
or UO_2332 (O_2332,N_17707,N_17035);
xnor UO_2333 (O_2333,N_19826,N_17578);
nor UO_2334 (O_2334,N_17417,N_18191);
or UO_2335 (O_2335,N_15809,N_17614);
nand UO_2336 (O_2336,N_18913,N_17728);
or UO_2337 (O_2337,N_18882,N_15393);
or UO_2338 (O_2338,N_17896,N_18358);
and UO_2339 (O_2339,N_19206,N_16941);
xnor UO_2340 (O_2340,N_17777,N_17805);
nor UO_2341 (O_2341,N_15141,N_18571);
xnor UO_2342 (O_2342,N_16148,N_17032);
and UO_2343 (O_2343,N_15876,N_16365);
nand UO_2344 (O_2344,N_16311,N_16575);
nor UO_2345 (O_2345,N_17795,N_15682);
and UO_2346 (O_2346,N_18974,N_17110);
nand UO_2347 (O_2347,N_19486,N_17555);
and UO_2348 (O_2348,N_15510,N_17686);
nor UO_2349 (O_2349,N_18785,N_16896);
or UO_2350 (O_2350,N_17011,N_19427);
xor UO_2351 (O_2351,N_17597,N_19690);
xnor UO_2352 (O_2352,N_19247,N_15533);
nor UO_2353 (O_2353,N_15063,N_19505);
nand UO_2354 (O_2354,N_16222,N_16944);
or UO_2355 (O_2355,N_18429,N_18632);
and UO_2356 (O_2356,N_19073,N_17794);
and UO_2357 (O_2357,N_17830,N_15583);
and UO_2358 (O_2358,N_15427,N_15392);
or UO_2359 (O_2359,N_15988,N_19790);
nand UO_2360 (O_2360,N_17272,N_19433);
nand UO_2361 (O_2361,N_16137,N_17684);
or UO_2362 (O_2362,N_18034,N_18932);
nor UO_2363 (O_2363,N_18849,N_18324);
or UO_2364 (O_2364,N_16797,N_15147);
nand UO_2365 (O_2365,N_17708,N_19359);
nand UO_2366 (O_2366,N_15362,N_19416);
nor UO_2367 (O_2367,N_17378,N_18285);
nor UO_2368 (O_2368,N_17335,N_17650);
or UO_2369 (O_2369,N_18535,N_16705);
xor UO_2370 (O_2370,N_16320,N_15218);
nand UO_2371 (O_2371,N_18528,N_17808);
nand UO_2372 (O_2372,N_19185,N_16874);
or UO_2373 (O_2373,N_19842,N_17042);
and UO_2374 (O_2374,N_16930,N_15279);
and UO_2375 (O_2375,N_15970,N_15869);
nor UO_2376 (O_2376,N_15998,N_16099);
nor UO_2377 (O_2377,N_15176,N_16037);
xor UO_2378 (O_2378,N_18095,N_17184);
xnor UO_2379 (O_2379,N_19469,N_15635);
nor UO_2380 (O_2380,N_18704,N_19481);
xor UO_2381 (O_2381,N_16547,N_19534);
nor UO_2382 (O_2382,N_15292,N_16063);
nand UO_2383 (O_2383,N_18230,N_19722);
nand UO_2384 (O_2384,N_18555,N_19014);
or UO_2385 (O_2385,N_15303,N_19896);
nor UO_2386 (O_2386,N_15747,N_19426);
xor UO_2387 (O_2387,N_16425,N_16016);
or UO_2388 (O_2388,N_18940,N_15652);
xnor UO_2389 (O_2389,N_18797,N_18101);
nor UO_2390 (O_2390,N_16671,N_15240);
xor UO_2391 (O_2391,N_19638,N_16550);
xor UO_2392 (O_2392,N_19130,N_17147);
and UO_2393 (O_2393,N_19470,N_17838);
and UO_2394 (O_2394,N_15464,N_15485);
and UO_2395 (O_2395,N_18245,N_16682);
xor UO_2396 (O_2396,N_16399,N_18333);
nand UO_2397 (O_2397,N_17292,N_15912);
xnor UO_2398 (O_2398,N_15332,N_18233);
or UO_2399 (O_2399,N_17785,N_18138);
nand UO_2400 (O_2400,N_18228,N_18417);
nor UO_2401 (O_2401,N_19680,N_17224);
and UO_2402 (O_2402,N_19373,N_15636);
nor UO_2403 (O_2403,N_15265,N_17418);
nor UO_2404 (O_2404,N_15836,N_19157);
nor UO_2405 (O_2405,N_18015,N_18171);
or UO_2406 (O_2406,N_15271,N_19243);
and UO_2407 (O_2407,N_19800,N_17227);
nand UO_2408 (O_2408,N_19555,N_18653);
nand UO_2409 (O_2409,N_18754,N_15364);
nand UO_2410 (O_2410,N_19669,N_15518);
nor UO_2411 (O_2411,N_16011,N_17063);
xnor UO_2412 (O_2412,N_19095,N_19592);
nor UO_2413 (O_2413,N_18115,N_18088);
xor UO_2414 (O_2414,N_17751,N_15350);
nor UO_2415 (O_2415,N_19636,N_15744);
nor UO_2416 (O_2416,N_18298,N_16160);
and UO_2417 (O_2417,N_18983,N_17997);
xnor UO_2418 (O_2418,N_16252,N_18736);
and UO_2419 (O_2419,N_17799,N_19484);
and UO_2420 (O_2420,N_18353,N_19495);
nand UO_2421 (O_2421,N_16899,N_16553);
xor UO_2422 (O_2422,N_19430,N_18122);
nand UO_2423 (O_2423,N_18857,N_18187);
xor UO_2424 (O_2424,N_19237,N_19205);
nor UO_2425 (O_2425,N_19561,N_15575);
and UO_2426 (O_2426,N_16631,N_15959);
xor UO_2427 (O_2427,N_19533,N_19854);
nand UO_2428 (O_2428,N_18028,N_19677);
and UO_2429 (O_2429,N_18497,N_17568);
and UO_2430 (O_2430,N_19567,N_15873);
nor UO_2431 (O_2431,N_19222,N_17004);
nand UO_2432 (O_2432,N_16863,N_19253);
or UO_2433 (O_2433,N_16047,N_17129);
xnor UO_2434 (O_2434,N_15737,N_17321);
xor UO_2435 (O_2435,N_19902,N_15005);
and UO_2436 (O_2436,N_18824,N_17507);
xor UO_2437 (O_2437,N_15234,N_18176);
and UO_2438 (O_2438,N_16738,N_17911);
or UO_2439 (O_2439,N_16105,N_17978);
and UO_2440 (O_2440,N_19865,N_16789);
xnor UO_2441 (O_2441,N_19601,N_16381);
nor UO_2442 (O_2442,N_18237,N_17092);
nand UO_2443 (O_2443,N_18313,N_16885);
nand UO_2444 (O_2444,N_18026,N_19704);
or UO_2445 (O_2445,N_16983,N_19753);
nor UO_2446 (O_2446,N_19417,N_16778);
nand UO_2447 (O_2447,N_19838,N_15769);
nor UO_2448 (O_2448,N_17623,N_17399);
and UO_2449 (O_2449,N_16831,N_17523);
or UO_2450 (O_2450,N_15181,N_19588);
nand UO_2451 (O_2451,N_15378,N_17085);
nor UO_2452 (O_2452,N_18329,N_18416);
or UO_2453 (O_2453,N_17719,N_17173);
xor UO_2454 (O_2454,N_16181,N_16958);
nor UO_2455 (O_2455,N_19077,N_16235);
nor UO_2456 (O_2456,N_15606,N_17543);
nand UO_2457 (O_2457,N_19341,N_19526);
and UO_2458 (O_2458,N_19947,N_15458);
nand UO_2459 (O_2459,N_17901,N_15811);
nor UO_2460 (O_2460,N_18044,N_16045);
and UO_2461 (O_2461,N_18524,N_18370);
xnor UO_2462 (O_2462,N_19034,N_18210);
xnor UO_2463 (O_2463,N_15942,N_15466);
nand UO_2464 (O_2464,N_19362,N_18903);
nor UO_2465 (O_2465,N_19236,N_18963);
nor UO_2466 (O_2466,N_19886,N_17082);
nand UO_2467 (O_2467,N_15494,N_18051);
and UO_2468 (O_2468,N_15929,N_15374);
or UO_2469 (O_2469,N_15154,N_19029);
nor UO_2470 (O_2470,N_19739,N_18234);
or UO_2471 (O_2471,N_19030,N_19429);
nor UO_2472 (O_2472,N_19515,N_16866);
nor UO_2473 (O_2473,N_15152,N_19104);
nand UO_2474 (O_2474,N_18426,N_17899);
nor UO_2475 (O_2475,N_18999,N_16820);
xnor UO_2476 (O_2476,N_16008,N_16470);
xor UO_2477 (O_2477,N_17806,N_19805);
and UO_2478 (O_2478,N_18192,N_19673);
nor UO_2479 (O_2479,N_18658,N_15155);
xnor UO_2480 (O_2480,N_17529,N_15513);
xnor UO_2481 (O_2481,N_15213,N_17940);
xor UO_2482 (O_2482,N_17033,N_18933);
and UO_2483 (O_2483,N_18852,N_17433);
or UO_2484 (O_2484,N_15891,N_16203);
nand UO_2485 (O_2485,N_15363,N_16895);
nor UO_2486 (O_2486,N_15158,N_16400);
nor UO_2487 (O_2487,N_15253,N_15142);
and UO_2488 (O_2488,N_16923,N_18010);
nor UO_2489 (O_2489,N_17912,N_19254);
nand UO_2490 (O_2490,N_19982,N_15675);
xnor UO_2491 (O_2491,N_17903,N_19519);
and UO_2492 (O_2492,N_17029,N_15473);
xor UO_2493 (O_2493,N_15472,N_18699);
nand UO_2494 (O_2494,N_18165,N_17280);
or UO_2495 (O_2495,N_16846,N_16417);
and UO_2496 (O_2496,N_18787,N_16579);
or UO_2497 (O_2497,N_15156,N_17120);
xor UO_2498 (O_2498,N_18825,N_19457);
nor UO_2499 (O_2499,N_17293,N_18011);
endmodule