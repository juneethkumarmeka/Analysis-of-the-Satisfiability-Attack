module basic_500_3000_500_4_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_154,In_448);
nor U1 (N_1,In_311,In_175);
or U2 (N_2,In_399,In_99);
nand U3 (N_3,In_244,In_475);
and U4 (N_4,In_22,In_21);
nand U5 (N_5,In_77,In_170);
xnor U6 (N_6,In_206,In_379);
xnor U7 (N_7,In_239,In_120);
xnor U8 (N_8,In_419,In_462);
nor U9 (N_9,In_414,In_288);
nand U10 (N_10,In_113,In_488);
and U11 (N_11,In_85,In_376);
nand U12 (N_12,In_400,In_299);
or U13 (N_13,In_439,In_396);
nand U14 (N_14,In_271,In_408);
xor U15 (N_15,In_269,In_200);
nor U16 (N_16,In_88,In_221);
nor U17 (N_17,In_342,In_493);
or U18 (N_18,In_330,In_483);
and U19 (N_19,In_132,In_178);
or U20 (N_20,In_160,In_263);
nand U21 (N_21,In_315,In_297);
or U22 (N_22,In_52,In_56);
or U23 (N_23,In_225,In_235);
nand U24 (N_24,In_286,In_322);
nand U25 (N_25,In_228,In_60);
and U26 (N_26,In_144,In_267);
nor U27 (N_27,In_54,In_82);
and U28 (N_28,In_147,In_385);
nor U29 (N_29,In_309,In_280);
xor U30 (N_30,In_50,In_308);
and U31 (N_31,In_199,In_116);
and U32 (N_32,In_422,In_4);
nor U33 (N_33,In_340,In_354);
and U34 (N_34,In_205,In_404);
and U35 (N_35,In_153,In_146);
nor U36 (N_36,In_166,In_119);
nor U37 (N_37,In_40,In_53);
xor U38 (N_38,In_167,In_69);
or U39 (N_39,In_245,In_435);
or U40 (N_40,In_403,In_91);
xnor U41 (N_41,In_209,In_183);
and U42 (N_42,In_361,In_370);
or U43 (N_43,In_430,In_378);
nand U44 (N_44,In_461,In_23);
xor U45 (N_45,In_432,In_27);
or U46 (N_46,In_14,In_496);
xnor U47 (N_47,In_445,In_94);
nand U48 (N_48,In_44,In_355);
xnor U49 (N_49,In_446,In_103);
and U50 (N_50,In_145,In_443);
or U51 (N_51,In_287,In_498);
nor U52 (N_52,In_464,In_185);
or U53 (N_53,In_331,In_426);
or U54 (N_54,In_352,In_150);
nor U55 (N_55,In_274,In_480);
xnor U56 (N_56,In_424,In_407);
and U57 (N_57,In_316,In_490);
xor U58 (N_58,In_97,In_236);
nand U59 (N_59,In_328,In_148);
nand U60 (N_60,In_394,In_230);
xnor U61 (N_61,In_468,In_36);
nor U62 (N_62,In_420,In_484);
and U63 (N_63,In_250,In_358);
or U64 (N_64,In_261,In_492);
nand U65 (N_65,In_135,In_359);
nor U66 (N_66,In_19,In_243);
xor U67 (N_67,In_26,In_465);
nand U68 (N_68,In_171,In_124);
nor U69 (N_69,In_179,In_393);
and U70 (N_70,In_363,In_278);
and U71 (N_71,In_382,In_471);
nand U72 (N_72,In_248,In_275);
xor U73 (N_73,In_59,In_104);
xnor U74 (N_74,In_126,In_128);
xor U75 (N_75,In_102,In_159);
nand U76 (N_76,In_497,In_454);
xor U77 (N_77,In_11,In_325);
and U78 (N_78,In_115,In_133);
nor U79 (N_79,In_2,In_350);
xnor U80 (N_80,In_70,In_8);
nor U81 (N_81,In_257,In_142);
xor U82 (N_82,In_117,In_143);
and U83 (N_83,In_442,In_74);
and U84 (N_84,In_140,In_392);
nor U85 (N_85,In_93,In_182);
xnor U86 (N_86,In_90,In_195);
xor U87 (N_87,In_216,In_42);
or U88 (N_88,In_138,In_292);
or U89 (N_89,In_34,In_181);
nand U90 (N_90,In_418,In_73);
xnor U91 (N_91,In_335,In_270);
xor U92 (N_92,In_253,In_212);
or U93 (N_93,In_196,In_406);
nor U94 (N_94,In_62,In_158);
xnor U95 (N_95,In_486,In_479);
nor U96 (N_96,In_217,In_177);
xnor U97 (N_97,In_321,In_298);
or U98 (N_98,In_118,In_203);
nor U99 (N_99,In_95,In_37);
xnor U100 (N_100,In_398,In_189);
nand U101 (N_101,In_81,In_106);
and U102 (N_102,In_49,In_86);
xor U103 (N_103,In_223,In_323);
nand U104 (N_104,In_360,In_38);
or U105 (N_105,In_459,In_65);
nand U106 (N_106,In_341,In_425);
xnor U107 (N_107,In_444,In_24);
or U108 (N_108,In_247,In_463);
and U109 (N_109,In_187,In_469);
or U110 (N_110,In_318,In_242);
nor U111 (N_111,In_57,In_482);
xnor U112 (N_112,In_282,In_326);
and U113 (N_113,In_213,In_381);
and U114 (N_114,In_114,In_285);
xnor U115 (N_115,In_43,In_423);
and U116 (N_116,In_35,In_305);
nor U117 (N_117,In_281,In_89);
or U118 (N_118,In_460,In_6);
and U119 (N_119,In_332,In_191);
and U120 (N_120,In_207,In_470);
and U121 (N_121,In_259,In_169);
nand U122 (N_122,In_306,In_333);
and U123 (N_123,In_180,In_174);
xor U124 (N_124,In_33,In_374);
xnor U125 (N_125,In_87,In_47);
or U126 (N_126,In_410,In_457);
xor U127 (N_127,In_96,In_421);
nor U128 (N_128,In_110,In_415);
xor U129 (N_129,In_413,In_238);
and U130 (N_130,In_17,In_487);
xnor U131 (N_131,In_112,In_266);
nand U132 (N_132,In_327,In_351);
xor U133 (N_133,In_208,In_391);
and U134 (N_134,In_339,In_329);
nor U135 (N_135,In_428,In_473);
xor U136 (N_136,In_176,In_64);
nand U137 (N_137,In_80,In_198);
nor U138 (N_138,In_122,In_397);
nand U139 (N_139,In_449,In_338);
nand U140 (N_140,In_313,In_163);
nand U141 (N_141,In_436,In_173);
nor U142 (N_142,In_450,In_485);
or U143 (N_143,In_455,In_277);
and U144 (N_144,In_71,In_211);
nor U145 (N_145,In_232,In_386);
and U146 (N_146,In_109,In_139);
xnor U147 (N_147,In_320,In_452);
and U148 (N_148,In_362,In_268);
xor U149 (N_149,In_226,In_188);
nand U150 (N_150,In_390,In_258);
nand U151 (N_151,In_499,In_151);
xnor U152 (N_152,In_39,In_210);
nor U153 (N_153,In_165,In_383);
or U154 (N_154,In_314,In_201);
nor U155 (N_155,In_18,In_447);
nor U156 (N_156,In_495,In_494);
nor U157 (N_157,In_29,In_79);
or U158 (N_158,In_51,In_251);
nor U159 (N_159,In_416,In_237);
xnor U160 (N_160,In_5,In_260);
xnor U161 (N_161,In_186,In_219);
xor U162 (N_162,In_409,In_367);
xnor U163 (N_163,In_265,In_125);
and U164 (N_164,In_458,In_105);
nor U165 (N_165,In_255,In_429);
nand U166 (N_166,In_231,In_7);
xnor U167 (N_167,In_215,In_155);
xnor U168 (N_168,In_453,In_149);
and U169 (N_169,In_369,In_312);
xnor U170 (N_170,In_344,In_387);
nand U171 (N_171,In_302,In_346);
nor U172 (N_172,In_256,In_375);
and U173 (N_173,In_276,In_131);
nor U174 (N_174,In_440,In_84);
nand U175 (N_175,In_254,In_295);
nand U176 (N_176,In_184,In_78);
or U177 (N_177,In_83,In_476);
nor U178 (N_178,In_30,In_46);
and U179 (N_179,In_290,In_371);
nor U180 (N_180,In_197,In_218);
and U181 (N_181,In_249,In_222);
nor U182 (N_182,In_405,In_161);
nor U183 (N_183,In_273,In_12);
and U184 (N_184,In_129,In_347);
xnor U185 (N_185,In_466,In_101);
or U186 (N_186,In_491,In_152);
xor U187 (N_187,In_1,In_301);
xor U188 (N_188,In_388,In_127);
or U189 (N_189,In_411,In_241);
or U190 (N_190,In_224,In_0);
nor U191 (N_191,In_427,In_204);
xor U192 (N_192,In_55,In_438);
or U193 (N_193,In_368,In_348);
nand U194 (N_194,In_193,In_310);
nand U195 (N_195,In_252,In_172);
or U196 (N_196,In_227,In_412);
nor U197 (N_197,In_296,In_58);
nand U198 (N_198,In_389,In_451);
nor U199 (N_199,In_433,In_220);
xnor U200 (N_200,In_395,In_272);
and U201 (N_201,In_41,In_75);
xnor U202 (N_202,In_123,In_107);
nand U203 (N_203,In_63,In_214);
or U204 (N_204,In_334,In_337);
nand U205 (N_205,In_137,In_264);
nor U206 (N_206,In_304,In_474);
nor U207 (N_207,In_202,In_111);
nand U208 (N_208,In_168,In_353);
nand U209 (N_209,In_467,In_324);
nor U210 (N_210,In_229,In_356);
nand U211 (N_211,In_134,In_293);
xnor U212 (N_212,In_31,In_364);
nand U213 (N_213,In_98,In_291);
and U214 (N_214,In_303,In_9);
xor U215 (N_215,In_141,In_76);
xnor U216 (N_216,In_16,In_164);
nor U217 (N_217,In_130,In_162);
or U218 (N_218,In_431,In_156);
nor U219 (N_219,In_262,In_45);
nand U220 (N_220,In_279,In_349);
xnor U221 (N_221,In_489,In_336);
and U222 (N_222,In_357,In_66);
xor U223 (N_223,In_345,In_481);
xor U224 (N_224,In_233,In_192);
and U225 (N_225,In_108,In_61);
nor U226 (N_226,In_373,In_100);
nor U227 (N_227,In_240,In_15);
and U228 (N_228,In_67,In_3);
and U229 (N_229,In_13,In_401);
and U230 (N_230,In_307,In_402);
xnor U231 (N_231,In_294,In_289);
nand U232 (N_232,In_372,In_477);
and U233 (N_233,In_25,In_434);
xor U234 (N_234,In_283,In_377);
or U235 (N_235,In_48,In_72);
xnor U236 (N_236,In_472,In_441);
nand U237 (N_237,In_380,In_121);
and U238 (N_238,In_478,In_437);
and U239 (N_239,In_343,In_366);
and U240 (N_240,In_246,In_68);
nor U241 (N_241,In_384,In_300);
or U242 (N_242,In_92,In_234);
and U243 (N_243,In_136,In_456);
nand U244 (N_244,In_157,In_190);
nand U245 (N_245,In_284,In_20);
nand U246 (N_246,In_365,In_28);
or U247 (N_247,In_194,In_417);
nand U248 (N_248,In_319,In_10);
or U249 (N_249,In_32,In_317);
nand U250 (N_250,In_124,In_496);
or U251 (N_251,In_332,In_330);
nor U252 (N_252,In_102,In_284);
nand U253 (N_253,In_216,In_164);
nand U254 (N_254,In_239,In_434);
nand U255 (N_255,In_91,In_86);
or U256 (N_256,In_114,In_277);
nand U257 (N_257,In_421,In_103);
xnor U258 (N_258,In_270,In_199);
or U259 (N_259,In_483,In_102);
or U260 (N_260,In_372,In_366);
nor U261 (N_261,In_95,In_261);
or U262 (N_262,In_138,In_403);
or U263 (N_263,In_411,In_416);
xor U264 (N_264,In_295,In_37);
nand U265 (N_265,In_28,In_285);
and U266 (N_266,In_241,In_290);
xor U267 (N_267,In_229,In_313);
and U268 (N_268,In_279,In_218);
nand U269 (N_269,In_339,In_409);
nor U270 (N_270,In_212,In_77);
nor U271 (N_271,In_373,In_54);
nand U272 (N_272,In_1,In_68);
and U273 (N_273,In_224,In_499);
or U274 (N_274,In_74,In_241);
xnor U275 (N_275,In_9,In_63);
nor U276 (N_276,In_63,In_451);
and U277 (N_277,In_401,In_296);
nor U278 (N_278,In_470,In_292);
xnor U279 (N_279,In_481,In_175);
nor U280 (N_280,In_133,In_178);
nor U281 (N_281,In_323,In_301);
and U282 (N_282,In_426,In_278);
nand U283 (N_283,In_408,In_186);
and U284 (N_284,In_89,In_462);
and U285 (N_285,In_289,In_182);
nor U286 (N_286,In_75,In_27);
or U287 (N_287,In_22,In_139);
or U288 (N_288,In_52,In_155);
and U289 (N_289,In_435,In_307);
or U290 (N_290,In_309,In_192);
nor U291 (N_291,In_51,In_270);
or U292 (N_292,In_326,In_175);
xor U293 (N_293,In_412,In_42);
and U294 (N_294,In_90,In_79);
nor U295 (N_295,In_126,In_21);
nand U296 (N_296,In_321,In_188);
nand U297 (N_297,In_35,In_143);
xnor U298 (N_298,In_256,In_32);
or U299 (N_299,In_284,In_185);
nand U300 (N_300,In_265,In_305);
nand U301 (N_301,In_342,In_336);
nor U302 (N_302,In_153,In_8);
xor U303 (N_303,In_409,In_169);
nand U304 (N_304,In_337,In_172);
xor U305 (N_305,In_119,In_424);
nand U306 (N_306,In_76,In_455);
xnor U307 (N_307,In_334,In_227);
or U308 (N_308,In_470,In_332);
nor U309 (N_309,In_421,In_16);
or U310 (N_310,In_275,In_151);
nand U311 (N_311,In_226,In_250);
or U312 (N_312,In_40,In_439);
and U313 (N_313,In_153,In_209);
nand U314 (N_314,In_14,In_162);
nor U315 (N_315,In_377,In_99);
nand U316 (N_316,In_447,In_205);
and U317 (N_317,In_166,In_191);
nor U318 (N_318,In_371,In_352);
or U319 (N_319,In_54,In_156);
xnor U320 (N_320,In_106,In_317);
and U321 (N_321,In_319,In_372);
and U322 (N_322,In_100,In_51);
or U323 (N_323,In_362,In_259);
nor U324 (N_324,In_278,In_207);
and U325 (N_325,In_156,In_69);
nor U326 (N_326,In_277,In_322);
or U327 (N_327,In_446,In_193);
nor U328 (N_328,In_469,In_34);
and U329 (N_329,In_184,In_492);
or U330 (N_330,In_5,In_464);
nor U331 (N_331,In_182,In_164);
nand U332 (N_332,In_301,In_198);
xor U333 (N_333,In_260,In_466);
and U334 (N_334,In_453,In_318);
nor U335 (N_335,In_292,In_283);
nor U336 (N_336,In_235,In_379);
nand U337 (N_337,In_447,In_364);
xnor U338 (N_338,In_32,In_258);
nand U339 (N_339,In_53,In_336);
nand U340 (N_340,In_220,In_113);
xor U341 (N_341,In_279,In_201);
xnor U342 (N_342,In_32,In_474);
or U343 (N_343,In_2,In_438);
or U344 (N_344,In_216,In_320);
and U345 (N_345,In_294,In_384);
nor U346 (N_346,In_264,In_427);
or U347 (N_347,In_137,In_1);
nand U348 (N_348,In_196,In_234);
nand U349 (N_349,In_69,In_449);
nor U350 (N_350,In_338,In_446);
xor U351 (N_351,In_428,In_274);
xnor U352 (N_352,In_57,In_254);
nor U353 (N_353,In_263,In_143);
nand U354 (N_354,In_275,In_381);
nand U355 (N_355,In_66,In_191);
or U356 (N_356,In_283,In_444);
xnor U357 (N_357,In_335,In_278);
or U358 (N_358,In_94,In_276);
nand U359 (N_359,In_344,In_30);
nor U360 (N_360,In_113,In_462);
xnor U361 (N_361,In_435,In_182);
and U362 (N_362,In_474,In_490);
nand U363 (N_363,In_184,In_123);
and U364 (N_364,In_132,In_264);
and U365 (N_365,In_218,In_299);
xor U366 (N_366,In_301,In_364);
nand U367 (N_367,In_202,In_310);
nor U368 (N_368,In_18,In_101);
and U369 (N_369,In_353,In_326);
nor U370 (N_370,In_480,In_183);
nand U371 (N_371,In_60,In_292);
xor U372 (N_372,In_443,In_391);
nor U373 (N_373,In_314,In_277);
and U374 (N_374,In_351,In_115);
nor U375 (N_375,In_271,In_413);
nor U376 (N_376,In_135,In_367);
and U377 (N_377,In_240,In_9);
nand U378 (N_378,In_257,In_210);
and U379 (N_379,In_99,In_176);
nor U380 (N_380,In_147,In_442);
nand U381 (N_381,In_408,In_19);
nor U382 (N_382,In_277,In_172);
nand U383 (N_383,In_463,In_130);
nand U384 (N_384,In_458,In_344);
nand U385 (N_385,In_139,In_222);
and U386 (N_386,In_324,In_475);
nand U387 (N_387,In_340,In_83);
nor U388 (N_388,In_420,In_149);
xnor U389 (N_389,In_111,In_451);
nand U390 (N_390,In_79,In_87);
xor U391 (N_391,In_331,In_242);
nand U392 (N_392,In_408,In_47);
nor U393 (N_393,In_60,In_388);
or U394 (N_394,In_105,In_8);
and U395 (N_395,In_191,In_322);
nor U396 (N_396,In_177,In_387);
nand U397 (N_397,In_58,In_36);
and U398 (N_398,In_232,In_362);
and U399 (N_399,In_492,In_470);
or U400 (N_400,In_39,In_390);
and U401 (N_401,In_140,In_43);
nand U402 (N_402,In_230,In_302);
nor U403 (N_403,In_359,In_344);
nand U404 (N_404,In_16,In_375);
nor U405 (N_405,In_102,In_168);
xnor U406 (N_406,In_288,In_55);
and U407 (N_407,In_298,In_6);
nand U408 (N_408,In_187,In_352);
and U409 (N_409,In_445,In_267);
nor U410 (N_410,In_225,In_264);
or U411 (N_411,In_414,In_58);
nor U412 (N_412,In_280,In_84);
or U413 (N_413,In_230,In_94);
nand U414 (N_414,In_54,In_295);
nor U415 (N_415,In_53,In_203);
xnor U416 (N_416,In_224,In_30);
xnor U417 (N_417,In_231,In_456);
nor U418 (N_418,In_7,In_291);
and U419 (N_419,In_4,In_89);
and U420 (N_420,In_352,In_356);
nor U421 (N_421,In_217,In_487);
and U422 (N_422,In_196,In_117);
or U423 (N_423,In_67,In_225);
or U424 (N_424,In_416,In_242);
xor U425 (N_425,In_15,In_254);
or U426 (N_426,In_380,In_46);
xnor U427 (N_427,In_479,In_81);
or U428 (N_428,In_319,In_49);
and U429 (N_429,In_421,In_373);
nand U430 (N_430,In_172,In_58);
and U431 (N_431,In_460,In_111);
xor U432 (N_432,In_403,In_226);
or U433 (N_433,In_70,In_187);
nor U434 (N_434,In_234,In_471);
and U435 (N_435,In_206,In_75);
nor U436 (N_436,In_397,In_425);
and U437 (N_437,In_468,In_262);
nor U438 (N_438,In_351,In_349);
nand U439 (N_439,In_109,In_320);
nand U440 (N_440,In_57,In_5);
and U441 (N_441,In_75,In_238);
nor U442 (N_442,In_49,In_150);
xor U443 (N_443,In_140,In_176);
xnor U444 (N_444,In_72,In_390);
nor U445 (N_445,In_327,In_205);
and U446 (N_446,In_479,In_393);
nand U447 (N_447,In_25,In_422);
xnor U448 (N_448,In_496,In_236);
nor U449 (N_449,In_37,In_274);
xnor U450 (N_450,In_165,In_82);
and U451 (N_451,In_333,In_195);
or U452 (N_452,In_325,In_16);
or U453 (N_453,In_360,In_420);
nor U454 (N_454,In_156,In_366);
nor U455 (N_455,In_179,In_242);
nand U456 (N_456,In_450,In_16);
nor U457 (N_457,In_202,In_81);
nor U458 (N_458,In_388,In_357);
or U459 (N_459,In_1,In_142);
or U460 (N_460,In_168,In_388);
nor U461 (N_461,In_188,In_206);
or U462 (N_462,In_108,In_235);
nand U463 (N_463,In_446,In_218);
nand U464 (N_464,In_382,In_196);
and U465 (N_465,In_160,In_152);
and U466 (N_466,In_365,In_114);
nand U467 (N_467,In_434,In_381);
nor U468 (N_468,In_213,In_303);
or U469 (N_469,In_192,In_414);
and U470 (N_470,In_46,In_302);
or U471 (N_471,In_294,In_160);
nor U472 (N_472,In_117,In_97);
xor U473 (N_473,In_375,In_380);
and U474 (N_474,In_36,In_417);
nor U475 (N_475,In_96,In_147);
xnor U476 (N_476,In_248,In_340);
nand U477 (N_477,In_473,In_467);
nand U478 (N_478,In_106,In_470);
nor U479 (N_479,In_3,In_126);
nor U480 (N_480,In_55,In_198);
nor U481 (N_481,In_472,In_47);
xnor U482 (N_482,In_73,In_179);
and U483 (N_483,In_348,In_461);
or U484 (N_484,In_496,In_208);
or U485 (N_485,In_130,In_429);
xor U486 (N_486,In_484,In_404);
nor U487 (N_487,In_375,In_140);
or U488 (N_488,In_291,In_402);
nand U489 (N_489,In_232,In_169);
nor U490 (N_490,In_92,In_498);
nand U491 (N_491,In_395,In_295);
nor U492 (N_492,In_81,In_75);
nor U493 (N_493,In_424,In_187);
nand U494 (N_494,In_134,In_76);
nor U495 (N_495,In_166,In_253);
nand U496 (N_496,In_356,In_306);
and U497 (N_497,In_140,In_187);
nand U498 (N_498,In_279,In_244);
nor U499 (N_499,In_139,In_424);
nand U500 (N_500,In_476,In_65);
xor U501 (N_501,In_382,In_96);
nand U502 (N_502,In_381,In_178);
or U503 (N_503,In_355,In_155);
xor U504 (N_504,In_449,In_3);
nand U505 (N_505,In_45,In_204);
or U506 (N_506,In_379,In_221);
or U507 (N_507,In_96,In_412);
nand U508 (N_508,In_425,In_6);
xnor U509 (N_509,In_402,In_175);
nor U510 (N_510,In_262,In_76);
or U511 (N_511,In_409,In_133);
and U512 (N_512,In_152,In_259);
and U513 (N_513,In_48,In_391);
and U514 (N_514,In_2,In_146);
xnor U515 (N_515,In_96,In_146);
nor U516 (N_516,In_117,In_113);
nor U517 (N_517,In_303,In_41);
nor U518 (N_518,In_336,In_430);
xnor U519 (N_519,In_148,In_252);
nor U520 (N_520,In_99,In_322);
nor U521 (N_521,In_342,In_120);
xor U522 (N_522,In_378,In_495);
and U523 (N_523,In_63,In_286);
nand U524 (N_524,In_200,In_474);
xor U525 (N_525,In_359,In_236);
and U526 (N_526,In_309,In_355);
nand U527 (N_527,In_358,In_164);
xnor U528 (N_528,In_252,In_233);
xnor U529 (N_529,In_32,In_273);
or U530 (N_530,In_351,In_398);
nor U531 (N_531,In_396,In_194);
xor U532 (N_532,In_114,In_352);
xnor U533 (N_533,In_110,In_371);
nor U534 (N_534,In_496,In_159);
nor U535 (N_535,In_64,In_236);
or U536 (N_536,In_164,In_135);
and U537 (N_537,In_167,In_214);
nor U538 (N_538,In_416,In_466);
and U539 (N_539,In_332,In_264);
nand U540 (N_540,In_434,In_52);
nor U541 (N_541,In_265,In_456);
or U542 (N_542,In_383,In_231);
xnor U543 (N_543,In_20,In_350);
nand U544 (N_544,In_361,In_486);
xor U545 (N_545,In_459,In_244);
xnor U546 (N_546,In_335,In_112);
xnor U547 (N_547,In_461,In_410);
nand U548 (N_548,In_466,In_393);
and U549 (N_549,In_163,In_46);
or U550 (N_550,In_16,In_163);
nor U551 (N_551,In_362,In_334);
xnor U552 (N_552,In_255,In_411);
nor U553 (N_553,In_394,In_76);
nand U554 (N_554,In_374,In_212);
or U555 (N_555,In_496,In_381);
nor U556 (N_556,In_161,In_400);
nor U557 (N_557,In_180,In_246);
nand U558 (N_558,In_405,In_402);
xor U559 (N_559,In_26,In_409);
nor U560 (N_560,In_219,In_94);
and U561 (N_561,In_249,In_51);
xnor U562 (N_562,In_481,In_277);
and U563 (N_563,In_141,In_449);
xor U564 (N_564,In_41,In_406);
nand U565 (N_565,In_261,In_61);
nor U566 (N_566,In_6,In_208);
and U567 (N_567,In_452,In_225);
and U568 (N_568,In_327,In_386);
nand U569 (N_569,In_172,In_431);
or U570 (N_570,In_366,In_395);
nand U571 (N_571,In_336,In_241);
or U572 (N_572,In_354,In_246);
or U573 (N_573,In_394,In_157);
xnor U574 (N_574,In_324,In_224);
nor U575 (N_575,In_207,In_312);
and U576 (N_576,In_475,In_161);
nand U577 (N_577,In_209,In_147);
nor U578 (N_578,In_156,In_367);
or U579 (N_579,In_421,In_190);
xnor U580 (N_580,In_354,In_351);
nor U581 (N_581,In_259,In_47);
nor U582 (N_582,In_384,In_145);
and U583 (N_583,In_461,In_440);
and U584 (N_584,In_302,In_490);
and U585 (N_585,In_51,In_153);
xnor U586 (N_586,In_74,In_267);
nand U587 (N_587,In_471,In_384);
or U588 (N_588,In_121,In_333);
xor U589 (N_589,In_456,In_371);
or U590 (N_590,In_161,In_42);
and U591 (N_591,In_399,In_69);
nor U592 (N_592,In_87,In_5);
xnor U593 (N_593,In_215,In_163);
and U594 (N_594,In_209,In_244);
and U595 (N_595,In_449,In_176);
or U596 (N_596,In_493,In_142);
xor U597 (N_597,In_128,In_231);
and U598 (N_598,In_6,In_260);
and U599 (N_599,In_109,In_79);
or U600 (N_600,In_118,In_177);
nor U601 (N_601,In_5,In_218);
xor U602 (N_602,In_343,In_184);
xor U603 (N_603,In_211,In_24);
nor U604 (N_604,In_344,In_377);
xor U605 (N_605,In_72,In_373);
and U606 (N_606,In_45,In_474);
or U607 (N_607,In_243,In_144);
and U608 (N_608,In_373,In_45);
nor U609 (N_609,In_29,In_467);
xnor U610 (N_610,In_252,In_285);
or U611 (N_611,In_27,In_244);
and U612 (N_612,In_265,In_405);
nand U613 (N_613,In_318,In_460);
and U614 (N_614,In_53,In_382);
or U615 (N_615,In_169,In_350);
and U616 (N_616,In_87,In_6);
nand U617 (N_617,In_423,In_155);
nand U618 (N_618,In_469,In_311);
or U619 (N_619,In_381,In_339);
nand U620 (N_620,In_152,In_126);
nor U621 (N_621,In_272,In_131);
nand U622 (N_622,In_321,In_194);
and U623 (N_623,In_308,In_327);
nor U624 (N_624,In_130,In_232);
or U625 (N_625,In_390,In_358);
nor U626 (N_626,In_190,In_177);
nor U627 (N_627,In_463,In_99);
nand U628 (N_628,In_456,In_454);
xor U629 (N_629,In_294,In_273);
nand U630 (N_630,In_193,In_271);
nor U631 (N_631,In_388,In_106);
xor U632 (N_632,In_424,In_127);
nand U633 (N_633,In_107,In_358);
nor U634 (N_634,In_369,In_343);
and U635 (N_635,In_37,In_187);
xor U636 (N_636,In_74,In_474);
xor U637 (N_637,In_156,In_106);
and U638 (N_638,In_413,In_469);
xnor U639 (N_639,In_41,In_297);
nand U640 (N_640,In_428,In_455);
and U641 (N_641,In_103,In_338);
nor U642 (N_642,In_186,In_444);
nand U643 (N_643,In_37,In_363);
nand U644 (N_644,In_368,In_160);
xnor U645 (N_645,In_238,In_449);
nor U646 (N_646,In_375,In_247);
nand U647 (N_647,In_124,In_265);
and U648 (N_648,In_477,In_375);
nor U649 (N_649,In_316,In_232);
or U650 (N_650,In_405,In_267);
or U651 (N_651,In_21,In_135);
xnor U652 (N_652,In_13,In_33);
nor U653 (N_653,In_428,In_137);
or U654 (N_654,In_84,In_313);
xnor U655 (N_655,In_291,In_404);
and U656 (N_656,In_81,In_107);
and U657 (N_657,In_301,In_148);
xnor U658 (N_658,In_184,In_357);
or U659 (N_659,In_299,In_194);
and U660 (N_660,In_279,In_422);
or U661 (N_661,In_123,In_96);
nor U662 (N_662,In_223,In_495);
and U663 (N_663,In_129,In_96);
nand U664 (N_664,In_274,In_102);
or U665 (N_665,In_389,In_234);
nor U666 (N_666,In_239,In_329);
nand U667 (N_667,In_457,In_426);
nand U668 (N_668,In_64,In_359);
and U669 (N_669,In_380,In_272);
nand U670 (N_670,In_277,In_136);
and U671 (N_671,In_427,In_297);
nand U672 (N_672,In_419,In_193);
nand U673 (N_673,In_84,In_65);
nor U674 (N_674,In_173,In_460);
nor U675 (N_675,In_423,In_4);
xnor U676 (N_676,In_163,In_21);
nor U677 (N_677,In_363,In_120);
or U678 (N_678,In_317,In_91);
or U679 (N_679,In_388,In_320);
nor U680 (N_680,In_452,In_439);
nand U681 (N_681,In_13,In_70);
xor U682 (N_682,In_234,In_302);
nor U683 (N_683,In_494,In_95);
xnor U684 (N_684,In_216,In_455);
or U685 (N_685,In_231,In_118);
nor U686 (N_686,In_209,In_110);
and U687 (N_687,In_302,In_39);
and U688 (N_688,In_88,In_245);
or U689 (N_689,In_373,In_433);
xnor U690 (N_690,In_368,In_367);
or U691 (N_691,In_342,In_152);
and U692 (N_692,In_309,In_223);
or U693 (N_693,In_364,In_231);
nor U694 (N_694,In_214,In_291);
xnor U695 (N_695,In_272,In_480);
nand U696 (N_696,In_377,In_216);
nor U697 (N_697,In_133,In_336);
and U698 (N_698,In_297,In_498);
and U699 (N_699,In_281,In_31);
nand U700 (N_700,In_131,In_49);
or U701 (N_701,In_486,In_330);
nand U702 (N_702,In_127,In_183);
or U703 (N_703,In_62,In_0);
nor U704 (N_704,In_345,In_251);
xor U705 (N_705,In_337,In_441);
or U706 (N_706,In_375,In_431);
nor U707 (N_707,In_119,In_17);
and U708 (N_708,In_107,In_101);
nand U709 (N_709,In_96,In_437);
and U710 (N_710,In_169,In_42);
and U711 (N_711,In_34,In_410);
nor U712 (N_712,In_488,In_4);
nor U713 (N_713,In_50,In_163);
xor U714 (N_714,In_438,In_124);
nor U715 (N_715,In_262,In_200);
nor U716 (N_716,In_275,In_231);
or U717 (N_717,In_43,In_367);
and U718 (N_718,In_100,In_41);
or U719 (N_719,In_12,In_255);
and U720 (N_720,In_400,In_167);
or U721 (N_721,In_46,In_68);
xnor U722 (N_722,In_470,In_270);
nand U723 (N_723,In_22,In_499);
xnor U724 (N_724,In_287,In_496);
and U725 (N_725,In_461,In_130);
nor U726 (N_726,In_279,In_54);
nand U727 (N_727,In_225,In_475);
or U728 (N_728,In_70,In_154);
nor U729 (N_729,In_199,In_234);
nand U730 (N_730,In_399,In_474);
and U731 (N_731,In_192,In_440);
or U732 (N_732,In_30,In_24);
nor U733 (N_733,In_116,In_328);
and U734 (N_734,In_419,In_488);
and U735 (N_735,In_154,In_484);
and U736 (N_736,In_120,In_402);
or U737 (N_737,In_474,In_480);
or U738 (N_738,In_124,In_94);
or U739 (N_739,In_355,In_32);
xor U740 (N_740,In_413,In_258);
nor U741 (N_741,In_251,In_38);
or U742 (N_742,In_496,In_215);
or U743 (N_743,In_74,In_371);
xnor U744 (N_744,In_155,In_47);
nor U745 (N_745,In_251,In_260);
or U746 (N_746,In_246,In_190);
nand U747 (N_747,In_175,In_299);
nand U748 (N_748,In_399,In_254);
xnor U749 (N_749,In_427,In_179);
nand U750 (N_750,N_262,N_203);
nor U751 (N_751,N_217,N_403);
xnor U752 (N_752,N_272,N_127);
nand U753 (N_753,N_42,N_341);
and U754 (N_754,N_125,N_484);
or U755 (N_755,N_181,N_316);
nand U756 (N_756,N_64,N_200);
and U757 (N_757,N_558,N_307);
nand U758 (N_758,N_164,N_730);
nor U759 (N_759,N_71,N_556);
and U760 (N_760,N_617,N_221);
nor U761 (N_761,N_573,N_627);
nor U762 (N_762,N_734,N_199);
xnor U763 (N_763,N_479,N_186);
nand U764 (N_764,N_655,N_140);
xnor U765 (N_765,N_615,N_303);
xor U766 (N_766,N_438,N_69);
xor U767 (N_767,N_687,N_511);
or U768 (N_768,N_674,N_582);
nor U769 (N_769,N_253,N_277);
xor U770 (N_770,N_78,N_294);
or U771 (N_771,N_683,N_95);
nand U772 (N_772,N_52,N_173);
or U773 (N_773,N_535,N_255);
nand U774 (N_774,N_317,N_352);
or U775 (N_775,N_565,N_232);
xnor U776 (N_776,N_624,N_409);
nand U777 (N_777,N_494,N_439);
nor U778 (N_778,N_265,N_292);
xor U779 (N_779,N_254,N_637);
nor U780 (N_780,N_109,N_612);
xor U781 (N_781,N_376,N_447);
nand U782 (N_782,N_51,N_118);
and U783 (N_783,N_562,N_508);
nor U784 (N_784,N_260,N_408);
nand U785 (N_785,N_611,N_521);
and U786 (N_786,N_168,N_205);
nor U787 (N_787,N_259,N_311);
nand U788 (N_788,N_87,N_645);
nor U789 (N_789,N_679,N_153);
nand U790 (N_790,N_339,N_407);
xnor U791 (N_791,N_183,N_257);
and U792 (N_792,N_510,N_418);
or U793 (N_793,N_746,N_157);
or U794 (N_794,N_24,N_583);
nand U795 (N_795,N_400,N_274);
nor U796 (N_796,N_246,N_513);
nor U797 (N_797,N_98,N_401);
xnor U798 (N_798,N_685,N_365);
or U799 (N_799,N_549,N_336);
and U800 (N_800,N_697,N_735);
nor U801 (N_801,N_239,N_606);
nand U802 (N_802,N_374,N_481);
or U803 (N_803,N_666,N_60);
xnor U804 (N_804,N_444,N_67);
or U805 (N_805,N_487,N_233);
nand U806 (N_806,N_563,N_660);
or U807 (N_807,N_198,N_538);
or U808 (N_808,N_680,N_11);
or U809 (N_809,N_218,N_58);
nor U810 (N_810,N_229,N_711);
nor U811 (N_811,N_120,N_35);
nand U812 (N_812,N_602,N_544);
and U813 (N_813,N_267,N_626);
xor U814 (N_814,N_672,N_344);
nor U815 (N_815,N_422,N_603);
nand U816 (N_816,N_471,N_426);
nand U817 (N_817,N_31,N_117);
nand U818 (N_818,N_144,N_428);
or U819 (N_819,N_543,N_643);
or U820 (N_820,N_727,N_696);
or U821 (N_821,N_13,N_248);
and U822 (N_822,N_701,N_12);
and U823 (N_823,N_387,N_45);
xnor U824 (N_824,N_247,N_595);
or U825 (N_825,N_113,N_326);
nand U826 (N_826,N_367,N_364);
xor U827 (N_827,N_665,N_673);
or U828 (N_828,N_80,N_642);
nand U829 (N_829,N_178,N_128);
or U830 (N_830,N_56,N_103);
xnor U831 (N_831,N_420,N_472);
nand U832 (N_832,N_397,N_518);
xnor U833 (N_833,N_502,N_542);
nor U834 (N_834,N_179,N_288);
and U835 (N_835,N_749,N_162);
nor U836 (N_836,N_550,N_41);
and U837 (N_837,N_499,N_610);
or U838 (N_838,N_335,N_351);
nand U839 (N_839,N_245,N_419);
nand U840 (N_840,N_314,N_713);
xnor U841 (N_841,N_105,N_366);
nand U842 (N_842,N_313,N_92);
and U843 (N_843,N_664,N_532);
nor U844 (N_844,N_442,N_86);
and U845 (N_845,N_273,N_141);
nor U846 (N_846,N_85,N_358);
xor U847 (N_847,N_89,N_96);
xnor U848 (N_848,N_15,N_70);
and U849 (N_849,N_159,N_656);
nand U850 (N_850,N_619,N_715);
or U851 (N_851,N_119,N_379);
nor U852 (N_852,N_576,N_68);
or U853 (N_853,N_709,N_516);
and U854 (N_854,N_413,N_286);
nor U855 (N_855,N_73,N_594);
or U856 (N_856,N_309,N_658);
nor U857 (N_857,N_54,N_353);
nand U858 (N_858,N_618,N_240);
xnor U859 (N_859,N_414,N_28);
xor U860 (N_860,N_670,N_567);
nand U861 (N_861,N_402,N_553);
nor U862 (N_862,N_75,N_150);
nand U863 (N_863,N_281,N_388);
nand U864 (N_864,N_210,N_321);
and U865 (N_865,N_546,N_710);
and U866 (N_866,N_725,N_410);
xor U867 (N_867,N_584,N_427);
nand U868 (N_868,N_686,N_505);
xor U869 (N_869,N_135,N_706);
and U870 (N_870,N_600,N_234);
or U871 (N_871,N_574,N_596);
or U872 (N_872,N_434,N_74);
or U873 (N_873,N_498,N_26);
nand U874 (N_874,N_623,N_393);
and U875 (N_875,N_129,N_88);
or U876 (N_876,N_305,N_340);
or U877 (N_877,N_417,N_638);
and U878 (N_878,N_431,N_346);
nand U879 (N_879,N_738,N_650);
nand U880 (N_880,N_302,N_279);
nor U881 (N_881,N_32,N_312);
and U882 (N_882,N_327,N_284);
nand U883 (N_883,N_328,N_158);
or U884 (N_884,N_289,N_228);
and U885 (N_885,N_264,N_545);
xor U886 (N_886,N_256,N_509);
or U887 (N_887,N_112,N_446);
or U888 (N_888,N_720,N_390);
nor U889 (N_889,N_458,N_18);
nor U890 (N_890,N_130,N_160);
nor U891 (N_891,N_65,N_383);
nor U892 (N_892,N_139,N_122);
nor U893 (N_893,N_172,N_121);
nand U894 (N_894,N_244,N_593);
nand U895 (N_895,N_251,N_377);
xnor U896 (N_896,N_592,N_478);
nor U897 (N_897,N_632,N_304);
nand U898 (N_898,N_136,N_382);
and U899 (N_899,N_504,N_693);
and U900 (N_900,N_375,N_4);
and U901 (N_901,N_450,N_741);
nand U902 (N_902,N_519,N_620);
nand U903 (N_903,N_213,N_241);
nand U904 (N_904,N_182,N_733);
or U905 (N_905,N_412,N_537);
and U906 (N_906,N_275,N_722);
and U907 (N_907,N_476,N_634);
nor U908 (N_908,N_671,N_224);
nand U909 (N_909,N_528,N_644);
nor U910 (N_910,N_635,N_718);
nor U911 (N_911,N_588,N_466);
nand U912 (N_912,N_622,N_628);
xor U913 (N_913,N_467,N_712);
or U914 (N_914,N_290,N_116);
nand U915 (N_915,N_9,N_453);
xnor U916 (N_916,N_395,N_525);
xnor U917 (N_917,N_227,N_47);
nor U918 (N_918,N_278,N_470);
nand U919 (N_919,N_455,N_193);
xnor U920 (N_920,N_743,N_194);
nand U921 (N_921,N_99,N_111);
or U922 (N_922,N_580,N_394);
nand U923 (N_923,N_315,N_299);
nor U924 (N_924,N_226,N_266);
nand U925 (N_925,N_404,N_250);
and U926 (N_926,N_359,N_94);
nor U927 (N_927,N_212,N_222);
and U928 (N_928,N_649,N_391);
or U929 (N_929,N_448,N_678);
and U930 (N_930,N_347,N_561);
or U931 (N_931,N_399,N_30);
nor U932 (N_932,N_406,N_451);
xor U933 (N_933,N_700,N_114);
nand U934 (N_934,N_325,N_270);
nor U935 (N_935,N_308,N_177);
nor U936 (N_936,N_386,N_654);
nor U937 (N_937,N_682,N_318);
nor U938 (N_938,N_601,N_380);
or U939 (N_939,N_430,N_0);
and U940 (N_940,N_296,N_134);
xnor U941 (N_941,N_560,N_243);
and U942 (N_942,N_287,N_398);
xnor U943 (N_943,N_322,N_231);
xnor U944 (N_944,N_40,N_357);
and U945 (N_945,N_263,N_491);
and U946 (N_946,N_577,N_372);
nand U947 (N_947,N_348,N_371);
and U948 (N_948,N_384,N_677);
and U949 (N_949,N_719,N_21);
nand U950 (N_950,N_483,N_166);
nor U951 (N_951,N_667,N_310);
nand U952 (N_952,N_539,N_625);
xor U953 (N_953,N_554,N_27);
nand U954 (N_954,N_66,N_517);
xor U955 (N_955,N_732,N_728);
nor U956 (N_956,N_614,N_605);
or U957 (N_957,N_101,N_43);
and U958 (N_958,N_690,N_640);
nor U959 (N_959,N_526,N_176);
or U960 (N_960,N_167,N_488);
xnor U961 (N_961,N_530,N_587);
nor U962 (N_962,N_146,N_49);
or U963 (N_963,N_571,N_416);
xor U964 (N_964,N_586,N_653);
nor U965 (N_965,N_559,N_342);
or U966 (N_966,N_154,N_2);
or U967 (N_967,N_124,N_661);
or U968 (N_968,N_541,N_22);
or U969 (N_969,N_138,N_350);
nand U970 (N_970,N_575,N_590);
or U971 (N_971,N_283,N_214);
or U972 (N_972,N_57,N_648);
or U973 (N_973,N_295,N_515);
and U974 (N_974,N_202,N_108);
or U975 (N_975,N_362,N_411);
and U976 (N_976,N_378,N_684);
or U977 (N_977,N_440,N_23);
xor U978 (N_978,N_717,N_578);
xnor U979 (N_979,N_482,N_306);
nor U980 (N_980,N_83,N_707);
or U981 (N_981,N_512,N_659);
nand U982 (N_982,N_454,N_529);
and U983 (N_983,N_17,N_195);
or U984 (N_984,N_676,N_360);
and U985 (N_985,N_230,N_189);
and U986 (N_986,N_506,N_465);
and U987 (N_987,N_631,N_564);
nand U988 (N_988,N_156,N_503);
and U989 (N_989,N_609,N_170);
nand U990 (N_990,N_81,N_389);
and U991 (N_991,N_581,N_201);
xor U992 (N_992,N_681,N_36);
or U993 (N_993,N_55,N_460);
and U994 (N_994,N_107,N_492);
nand U995 (N_995,N_25,N_16);
or U996 (N_996,N_531,N_84);
or U997 (N_997,N_744,N_46);
xnor U998 (N_998,N_459,N_361);
nor U999 (N_999,N_197,N_208);
nor U1000 (N_1000,N_363,N_337);
nor U1001 (N_1001,N_90,N_557);
and U1002 (N_1002,N_249,N_333);
xnor U1003 (N_1003,N_82,N_276);
xor U1004 (N_1004,N_745,N_219);
and U1005 (N_1005,N_19,N_106);
nand U1006 (N_1006,N_669,N_485);
and U1007 (N_1007,N_691,N_271);
and U1008 (N_1008,N_207,N_432);
nand U1009 (N_1009,N_143,N_385);
nand U1010 (N_1010,N_3,N_211);
nand U1011 (N_1011,N_613,N_527);
nor U1012 (N_1012,N_196,N_433);
and U1013 (N_1013,N_258,N_209);
or U1014 (N_1014,N_486,N_100);
or U1015 (N_1015,N_437,N_716);
nand U1016 (N_1016,N_332,N_345);
nand U1017 (N_1017,N_185,N_282);
nor U1018 (N_1018,N_126,N_552);
and U1019 (N_1019,N_591,N_423);
nor U1020 (N_1020,N_147,N_748);
xor U1021 (N_1021,N_191,N_238);
nand U1022 (N_1022,N_721,N_269);
nor U1023 (N_1023,N_174,N_373);
nand U1024 (N_1024,N_489,N_97);
nand U1025 (N_1025,N_441,N_39);
nand U1026 (N_1026,N_14,N_705);
nor U1027 (N_1027,N_425,N_547);
nor U1028 (N_1028,N_598,N_343);
xnor U1029 (N_1029,N_731,N_44);
nor U1030 (N_1030,N_616,N_142);
or U1031 (N_1031,N_657,N_534);
nand U1032 (N_1032,N_452,N_497);
xnor U1033 (N_1033,N_38,N_698);
and U1034 (N_1034,N_520,N_464);
or U1035 (N_1035,N_72,N_102);
or U1036 (N_1036,N_688,N_8);
nor U1037 (N_1037,N_714,N_297);
and U1038 (N_1038,N_93,N_742);
or U1039 (N_1039,N_572,N_220);
nor U1040 (N_1040,N_692,N_242);
and U1041 (N_1041,N_501,N_568);
nand U1042 (N_1042,N_76,N_729);
nor U1043 (N_1043,N_639,N_349);
nand U1044 (N_1044,N_20,N_694);
or U1045 (N_1045,N_1,N_5);
nor U1046 (N_1046,N_215,N_368);
nor U1047 (N_1047,N_555,N_169);
and U1048 (N_1048,N_702,N_689);
or U1049 (N_1049,N_708,N_291);
and U1050 (N_1050,N_443,N_338);
nor U1051 (N_1051,N_500,N_331);
and U1052 (N_1052,N_225,N_330);
and U1053 (N_1053,N_236,N_187);
or U1054 (N_1054,N_695,N_115);
and U1055 (N_1055,N_490,N_123);
nor U1056 (N_1056,N_171,N_533);
nand U1057 (N_1057,N_536,N_474);
nor U1058 (N_1058,N_405,N_175);
or U1059 (N_1059,N_137,N_651);
xnor U1060 (N_1060,N_355,N_323);
and U1061 (N_1061,N_110,N_381);
or U1062 (N_1062,N_462,N_704);
nor U1063 (N_1063,N_320,N_29);
and U1064 (N_1064,N_737,N_468);
nor U1065 (N_1065,N_151,N_324);
xor U1066 (N_1066,N_608,N_6);
and U1067 (N_1067,N_62,N_190);
nand U1068 (N_1068,N_566,N_133);
xor U1069 (N_1069,N_740,N_652);
and U1070 (N_1070,N_597,N_463);
nand U1071 (N_1071,N_223,N_461);
nor U1072 (N_1072,N_10,N_50);
nor U1073 (N_1073,N_421,N_569);
or U1074 (N_1074,N_445,N_496);
xor U1075 (N_1075,N_34,N_514);
and U1076 (N_1076,N_59,N_132);
xor U1077 (N_1077,N_285,N_429);
nor U1078 (N_1078,N_216,N_724);
nand U1079 (N_1079,N_235,N_579);
nor U1080 (N_1080,N_630,N_449);
xnor U1081 (N_1081,N_280,N_300);
nand U1082 (N_1082,N_61,N_206);
nand U1083 (N_1083,N_599,N_334);
or U1084 (N_1084,N_524,N_723);
and U1085 (N_1085,N_252,N_354);
xnor U1086 (N_1086,N_237,N_152);
nand U1087 (N_1087,N_415,N_646);
and U1088 (N_1088,N_165,N_53);
nand U1089 (N_1089,N_104,N_493);
and U1090 (N_1090,N_63,N_155);
xnor U1091 (N_1091,N_356,N_149);
nor U1092 (N_1092,N_739,N_621);
nor U1093 (N_1093,N_7,N_161);
or U1094 (N_1094,N_663,N_522);
xnor U1095 (N_1095,N_37,N_469);
xor U1096 (N_1096,N_629,N_329);
and U1097 (N_1097,N_145,N_475);
or U1098 (N_1098,N_424,N_77);
nand U1099 (N_1099,N_633,N_523);
and U1100 (N_1100,N_293,N_726);
xor U1101 (N_1101,N_319,N_507);
and U1102 (N_1102,N_551,N_435);
xnor U1103 (N_1103,N_192,N_456);
nand U1104 (N_1104,N_585,N_392);
or U1105 (N_1105,N_261,N_268);
and U1106 (N_1106,N_647,N_369);
or U1107 (N_1107,N_747,N_736);
and U1108 (N_1108,N_641,N_636);
xor U1109 (N_1109,N_188,N_184);
nor U1110 (N_1110,N_675,N_589);
nor U1111 (N_1111,N_604,N_607);
and U1112 (N_1112,N_703,N_301);
and U1113 (N_1113,N_131,N_436);
nor U1114 (N_1114,N_548,N_163);
xnor U1115 (N_1115,N_662,N_495);
or U1116 (N_1116,N_480,N_79);
nand U1117 (N_1117,N_396,N_668);
nand U1118 (N_1118,N_204,N_477);
nor U1119 (N_1119,N_699,N_48);
and U1120 (N_1120,N_457,N_33);
or U1121 (N_1121,N_540,N_473);
nor U1122 (N_1122,N_570,N_91);
nand U1123 (N_1123,N_370,N_298);
nor U1124 (N_1124,N_148,N_180);
xnor U1125 (N_1125,N_100,N_170);
nor U1126 (N_1126,N_121,N_35);
nand U1127 (N_1127,N_39,N_426);
xnor U1128 (N_1128,N_346,N_157);
nor U1129 (N_1129,N_614,N_135);
xnor U1130 (N_1130,N_72,N_168);
and U1131 (N_1131,N_155,N_450);
or U1132 (N_1132,N_205,N_272);
and U1133 (N_1133,N_79,N_145);
or U1134 (N_1134,N_665,N_205);
xnor U1135 (N_1135,N_492,N_210);
xor U1136 (N_1136,N_740,N_452);
nand U1137 (N_1137,N_144,N_157);
xor U1138 (N_1138,N_664,N_7);
xor U1139 (N_1139,N_515,N_284);
or U1140 (N_1140,N_68,N_496);
and U1141 (N_1141,N_463,N_605);
nand U1142 (N_1142,N_722,N_324);
or U1143 (N_1143,N_30,N_444);
and U1144 (N_1144,N_614,N_421);
or U1145 (N_1145,N_684,N_550);
and U1146 (N_1146,N_615,N_53);
nor U1147 (N_1147,N_412,N_151);
and U1148 (N_1148,N_723,N_384);
or U1149 (N_1149,N_288,N_538);
and U1150 (N_1150,N_707,N_704);
nand U1151 (N_1151,N_727,N_75);
xnor U1152 (N_1152,N_712,N_8);
or U1153 (N_1153,N_195,N_554);
or U1154 (N_1154,N_519,N_418);
or U1155 (N_1155,N_606,N_351);
xnor U1156 (N_1156,N_330,N_243);
xnor U1157 (N_1157,N_218,N_724);
nand U1158 (N_1158,N_643,N_101);
xor U1159 (N_1159,N_547,N_186);
xor U1160 (N_1160,N_650,N_544);
nor U1161 (N_1161,N_604,N_193);
xor U1162 (N_1162,N_31,N_269);
nand U1163 (N_1163,N_361,N_395);
or U1164 (N_1164,N_384,N_75);
nand U1165 (N_1165,N_32,N_116);
xnor U1166 (N_1166,N_379,N_558);
nor U1167 (N_1167,N_353,N_37);
or U1168 (N_1168,N_302,N_222);
nor U1169 (N_1169,N_136,N_172);
nand U1170 (N_1170,N_38,N_462);
xnor U1171 (N_1171,N_410,N_696);
and U1172 (N_1172,N_72,N_600);
or U1173 (N_1173,N_368,N_321);
nor U1174 (N_1174,N_524,N_163);
xnor U1175 (N_1175,N_550,N_209);
nand U1176 (N_1176,N_679,N_213);
nand U1177 (N_1177,N_740,N_473);
xnor U1178 (N_1178,N_41,N_530);
nor U1179 (N_1179,N_394,N_589);
nand U1180 (N_1180,N_344,N_535);
xor U1181 (N_1181,N_185,N_747);
nor U1182 (N_1182,N_325,N_17);
or U1183 (N_1183,N_345,N_178);
nor U1184 (N_1184,N_739,N_610);
xor U1185 (N_1185,N_607,N_143);
xnor U1186 (N_1186,N_281,N_644);
or U1187 (N_1187,N_653,N_158);
and U1188 (N_1188,N_579,N_605);
xnor U1189 (N_1189,N_647,N_152);
nor U1190 (N_1190,N_145,N_547);
or U1191 (N_1191,N_716,N_514);
and U1192 (N_1192,N_158,N_485);
or U1193 (N_1193,N_94,N_614);
or U1194 (N_1194,N_118,N_286);
nand U1195 (N_1195,N_654,N_544);
and U1196 (N_1196,N_570,N_566);
xnor U1197 (N_1197,N_273,N_735);
or U1198 (N_1198,N_585,N_80);
or U1199 (N_1199,N_355,N_62);
nor U1200 (N_1200,N_463,N_386);
nor U1201 (N_1201,N_54,N_717);
xnor U1202 (N_1202,N_336,N_183);
or U1203 (N_1203,N_40,N_483);
and U1204 (N_1204,N_697,N_378);
xnor U1205 (N_1205,N_481,N_575);
nor U1206 (N_1206,N_26,N_482);
xor U1207 (N_1207,N_593,N_196);
xor U1208 (N_1208,N_236,N_109);
xor U1209 (N_1209,N_258,N_629);
nand U1210 (N_1210,N_343,N_449);
nand U1211 (N_1211,N_280,N_380);
or U1212 (N_1212,N_317,N_636);
nand U1213 (N_1213,N_313,N_242);
and U1214 (N_1214,N_720,N_236);
nor U1215 (N_1215,N_224,N_483);
xor U1216 (N_1216,N_238,N_567);
and U1217 (N_1217,N_307,N_468);
xnor U1218 (N_1218,N_197,N_103);
xor U1219 (N_1219,N_670,N_116);
nor U1220 (N_1220,N_314,N_397);
nor U1221 (N_1221,N_709,N_62);
or U1222 (N_1222,N_55,N_336);
nor U1223 (N_1223,N_454,N_138);
or U1224 (N_1224,N_212,N_105);
nand U1225 (N_1225,N_18,N_639);
nor U1226 (N_1226,N_385,N_371);
and U1227 (N_1227,N_473,N_719);
or U1228 (N_1228,N_442,N_121);
nand U1229 (N_1229,N_259,N_291);
nor U1230 (N_1230,N_308,N_95);
nor U1231 (N_1231,N_557,N_280);
xnor U1232 (N_1232,N_197,N_611);
xnor U1233 (N_1233,N_478,N_579);
or U1234 (N_1234,N_678,N_218);
nor U1235 (N_1235,N_611,N_517);
or U1236 (N_1236,N_393,N_433);
or U1237 (N_1237,N_319,N_238);
xnor U1238 (N_1238,N_189,N_332);
nand U1239 (N_1239,N_569,N_294);
nand U1240 (N_1240,N_732,N_354);
or U1241 (N_1241,N_390,N_124);
nor U1242 (N_1242,N_35,N_575);
xnor U1243 (N_1243,N_8,N_678);
xor U1244 (N_1244,N_317,N_355);
nand U1245 (N_1245,N_363,N_335);
nor U1246 (N_1246,N_613,N_3);
and U1247 (N_1247,N_500,N_393);
and U1248 (N_1248,N_551,N_550);
nand U1249 (N_1249,N_181,N_170);
or U1250 (N_1250,N_420,N_598);
and U1251 (N_1251,N_34,N_210);
xor U1252 (N_1252,N_742,N_154);
xor U1253 (N_1253,N_449,N_292);
or U1254 (N_1254,N_361,N_327);
or U1255 (N_1255,N_168,N_49);
and U1256 (N_1256,N_582,N_3);
xnor U1257 (N_1257,N_732,N_341);
nor U1258 (N_1258,N_409,N_496);
or U1259 (N_1259,N_218,N_328);
and U1260 (N_1260,N_625,N_156);
nand U1261 (N_1261,N_427,N_432);
or U1262 (N_1262,N_501,N_627);
and U1263 (N_1263,N_193,N_247);
xnor U1264 (N_1264,N_410,N_130);
xor U1265 (N_1265,N_546,N_207);
or U1266 (N_1266,N_61,N_611);
nor U1267 (N_1267,N_421,N_617);
nor U1268 (N_1268,N_216,N_79);
and U1269 (N_1269,N_279,N_262);
or U1270 (N_1270,N_391,N_333);
nor U1271 (N_1271,N_55,N_726);
xnor U1272 (N_1272,N_304,N_567);
or U1273 (N_1273,N_598,N_730);
or U1274 (N_1274,N_338,N_283);
nand U1275 (N_1275,N_573,N_302);
nor U1276 (N_1276,N_621,N_3);
nor U1277 (N_1277,N_643,N_36);
or U1278 (N_1278,N_338,N_394);
nand U1279 (N_1279,N_739,N_325);
xnor U1280 (N_1280,N_732,N_748);
and U1281 (N_1281,N_564,N_42);
or U1282 (N_1282,N_493,N_601);
nand U1283 (N_1283,N_665,N_301);
and U1284 (N_1284,N_493,N_606);
nand U1285 (N_1285,N_617,N_741);
nand U1286 (N_1286,N_468,N_359);
and U1287 (N_1287,N_663,N_158);
xnor U1288 (N_1288,N_329,N_288);
or U1289 (N_1289,N_510,N_523);
xnor U1290 (N_1290,N_164,N_426);
nor U1291 (N_1291,N_299,N_46);
nand U1292 (N_1292,N_742,N_291);
nand U1293 (N_1293,N_70,N_693);
xnor U1294 (N_1294,N_234,N_651);
nor U1295 (N_1295,N_189,N_411);
nor U1296 (N_1296,N_144,N_746);
or U1297 (N_1297,N_345,N_55);
xnor U1298 (N_1298,N_255,N_558);
and U1299 (N_1299,N_146,N_54);
and U1300 (N_1300,N_476,N_155);
or U1301 (N_1301,N_392,N_569);
nor U1302 (N_1302,N_71,N_410);
nor U1303 (N_1303,N_719,N_11);
and U1304 (N_1304,N_587,N_20);
xor U1305 (N_1305,N_431,N_453);
xor U1306 (N_1306,N_713,N_589);
and U1307 (N_1307,N_220,N_336);
or U1308 (N_1308,N_322,N_395);
nand U1309 (N_1309,N_350,N_487);
xor U1310 (N_1310,N_22,N_211);
or U1311 (N_1311,N_225,N_494);
and U1312 (N_1312,N_335,N_99);
and U1313 (N_1313,N_281,N_597);
or U1314 (N_1314,N_575,N_22);
xor U1315 (N_1315,N_210,N_274);
nor U1316 (N_1316,N_396,N_51);
xor U1317 (N_1317,N_158,N_622);
nor U1318 (N_1318,N_454,N_307);
nor U1319 (N_1319,N_315,N_233);
and U1320 (N_1320,N_728,N_736);
nor U1321 (N_1321,N_559,N_395);
nor U1322 (N_1322,N_548,N_202);
nand U1323 (N_1323,N_172,N_342);
nand U1324 (N_1324,N_332,N_701);
nand U1325 (N_1325,N_345,N_310);
or U1326 (N_1326,N_203,N_563);
xor U1327 (N_1327,N_94,N_232);
and U1328 (N_1328,N_577,N_85);
xor U1329 (N_1329,N_23,N_88);
and U1330 (N_1330,N_593,N_710);
and U1331 (N_1331,N_551,N_218);
and U1332 (N_1332,N_639,N_571);
xnor U1333 (N_1333,N_32,N_499);
nor U1334 (N_1334,N_355,N_679);
xnor U1335 (N_1335,N_698,N_605);
nor U1336 (N_1336,N_287,N_365);
or U1337 (N_1337,N_17,N_278);
and U1338 (N_1338,N_499,N_612);
xnor U1339 (N_1339,N_99,N_578);
or U1340 (N_1340,N_328,N_648);
xnor U1341 (N_1341,N_745,N_118);
nor U1342 (N_1342,N_140,N_469);
nand U1343 (N_1343,N_133,N_465);
and U1344 (N_1344,N_438,N_16);
nand U1345 (N_1345,N_9,N_302);
nor U1346 (N_1346,N_64,N_1);
xnor U1347 (N_1347,N_23,N_124);
xor U1348 (N_1348,N_367,N_465);
xnor U1349 (N_1349,N_136,N_378);
or U1350 (N_1350,N_364,N_434);
and U1351 (N_1351,N_469,N_507);
and U1352 (N_1352,N_560,N_186);
nand U1353 (N_1353,N_222,N_619);
xnor U1354 (N_1354,N_438,N_35);
nand U1355 (N_1355,N_445,N_580);
and U1356 (N_1356,N_439,N_398);
and U1357 (N_1357,N_39,N_157);
nor U1358 (N_1358,N_710,N_626);
nor U1359 (N_1359,N_238,N_334);
xnor U1360 (N_1360,N_613,N_412);
and U1361 (N_1361,N_84,N_426);
nor U1362 (N_1362,N_255,N_23);
or U1363 (N_1363,N_203,N_161);
or U1364 (N_1364,N_119,N_19);
nand U1365 (N_1365,N_699,N_141);
nor U1366 (N_1366,N_533,N_236);
xor U1367 (N_1367,N_643,N_683);
nand U1368 (N_1368,N_289,N_450);
xnor U1369 (N_1369,N_71,N_649);
and U1370 (N_1370,N_361,N_488);
or U1371 (N_1371,N_563,N_736);
nor U1372 (N_1372,N_508,N_242);
nor U1373 (N_1373,N_266,N_44);
or U1374 (N_1374,N_90,N_548);
and U1375 (N_1375,N_306,N_391);
nand U1376 (N_1376,N_151,N_184);
nor U1377 (N_1377,N_633,N_666);
xnor U1378 (N_1378,N_65,N_52);
nor U1379 (N_1379,N_152,N_421);
nor U1380 (N_1380,N_509,N_312);
nand U1381 (N_1381,N_509,N_385);
and U1382 (N_1382,N_304,N_67);
xnor U1383 (N_1383,N_144,N_358);
nor U1384 (N_1384,N_345,N_622);
xnor U1385 (N_1385,N_130,N_221);
and U1386 (N_1386,N_723,N_551);
nand U1387 (N_1387,N_67,N_432);
nor U1388 (N_1388,N_324,N_247);
xor U1389 (N_1389,N_366,N_30);
and U1390 (N_1390,N_568,N_199);
or U1391 (N_1391,N_508,N_311);
xnor U1392 (N_1392,N_396,N_681);
nand U1393 (N_1393,N_76,N_509);
nand U1394 (N_1394,N_562,N_379);
xor U1395 (N_1395,N_428,N_557);
or U1396 (N_1396,N_409,N_230);
and U1397 (N_1397,N_582,N_337);
nor U1398 (N_1398,N_261,N_418);
and U1399 (N_1399,N_260,N_37);
nor U1400 (N_1400,N_617,N_467);
or U1401 (N_1401,N_394,N_397);
and U1402 (N_1402,N_719,N_660);
and U1403 (N_1403,N_292,N_104);
nand U1404 (N_1404,N_629,N_673);
and U1405 (N_1405,N_3,N_366);
nand U1406 (N_1406,N_552,N_67);
nor U1407 (N_1407,N_250,N_635);
nand U1408 (N_1408,N_207,N_253);
or U1409 (N_1409,N_365,N_76);
and U1410 (N_1410,N_274,N_688);
or U1411 (N_1411,N_206,N_113);
nor U1412 (N_1412,N_298,N_227);
nor U1413 (N_1413,N_457,N_37);
and U1414 (N_1414,N_310,N_405);
xnor U1415 (N_1415,N_637,N_178);
nand U1416 (N_1416,N_143,N_676);
and U1417 (N_1417,N_144,N_457);
nand U1418 (N_1418,N_162,N_600);
nor U1419 (N_1419,N_748,N_268);
nand U1420 (N_1420,N_463,N_213);
and U1421 (N_1421,N_55,N_636);
nor U1422 (N_1422,N_10,N_581);
or U1423 (N_1423,N_379,N_381);
nor U1424 (N_1424,N_219,N_236);
and U1425 (N_1425,N_516,N_41);
and U1426 (N_1426,N_243,N_112);
nand U1427 (N_1427,N_185,N_281);
and U1428 (N_1428,N_313,N_219);
and U1429 (N_1429,N_377,N_176);
nand U1430 (N_1430,N_565,N_408);
nor U1431 (N_1431,N_69,N_539);
nor U1432 (N_1432,N_163,N_390);
xor U1433 (N_1433,N_231,N_281);
nor U1434 (N_1434,N_505,N_597);
xnor U1435 (N_1435,N_76,N_221);
nor U1436 (N_1436,N_170,N_183);
xor U1437 (N_1437,N_66,N_395);
or U1438 (N_1438,N_580,N_601);
nor U1439 (N_1439,N_289,N_29);
nand U1440 (N_1440,N_412,N_377);
xor U1441 (N_1441,N_667,N_177);
or U1442 (N_1442,N_334,N_515);
nand U1443 (N_1443,N_14,N_726);
nor U1444 (N_1444,N_255,N_47);
xor U1445 (N_1445,N_64,N_184);
nand U1446 (N_1446,N_394,N_204);
nand U1447 (N_1447,N_472,N_13);
or U1448 (N_1448,N_348,N_582);
or U1449 (N_1449,N_176,N_89);
nand U1450 (N_1450,N_668,N_207);
or U1451 (N_1451,N_407,N_302);
xnor U1452 (N_1452,N_302,N_216);
xor U1453 (N_1453,N_213,N_537);
xnor U1454 (N_1454,N_1,N_588);
or U1455 (N_1455,N_649,N_431);
and U1456 (N_1456,N_254,N_715);
nor U1457 (N_1457,N_126,N_652);
xor U1458 (N_1458,N_443,N_400);
nor U1459 (N_1459,N_310,N_194);
xor U1460 (N_1460,N_662,N_474);
nand U1461 (N_1461,N_149,N_642);
nand U1462 (N_1462,N_157,N_632);
and U1463 (N_1463,N_126,N_261);
and U1464 (N_1464,N_459,N_194);
xor U1465 (N_1465,N_220,N_543);
or U1466 (N_1466,N_251,N_109);
xnor U1467 (N_1467,N_364,N_210);
or U1468 (N_1468,N_402,N_451);
nor U1469 (N_1469,N_331,N_632);
and U1470 (N_1470,N_226,N_290);
and U1471 (N_1471,N_207,N_560);
or U1472 (N_1472,N_326,N_506);
or U1473 (N_1473,N_469,N_493);
xor U1474 (N_1474,N_212,N_591);
or U1475 (N_1475,N_420,N_71);
nand U1476 (N_1476,N_608,N_138);
nand U1477 (N_1477,N_58,N_93);
and U1478 (N_1478,N_395,N_214);
nand U1479 (N_1479,N_164,N_742);
nand U1480 (N_1480,N_743,N_351);
and U1481 (N_1481,N_61,N_493);
and U1482 (N_1482,N_438,N_653);
xor U1483 (N_1483,N_160,N_83);
and U1484 (N_1484,N_454,N_333);
and U1485 (N_1485,N_426,N_102);
and U1486 (N_1486,N_397,N_642);
xnor U1487 (N_1487,N_485,N_532);
or U1488 (N_1488,N_151,N_417);
xor U1489 (N_1489,N_365,N_0);
nor U1490 (N_1490,N_110,N_384);
and U1491 (N_1491,N_586,N_193);
or U1492 (N_1492,N_278,N_144);
nand U1493 (N_1493,N_374,N_369);
nand U1494 (N_1494,N_615,N_82);
nor U1495 (N_1495,N_204,N_590);
and U1496 (N_1496,N_220,N_3);
nand U1497 (N_1497,N_678,N_433);
nand U1498 (N_1498,N_373,N_426);
nand U1499 (N_1499,N_317,N_106);
nor U1500 (N_1500,N_783,N_998);
or U1501 (N_1501,N_1386,N_971);
xnor U1502 (N_1502,N_1367,N_1389);
or U1503 (N_1503,N_1262,N_1366);
and U1504 (N_1504,N_1381,N_1083);
and U1505 (N_1505,N_757,N_1337);
and U1506 (N_1506,N_1498,N_1138);
or U1507 (N_1507,N_1313,N_1466);
or U1508 (N_1508,N_1006,N_1155);
and U1509 (N_1509,N_1148,N_1424);
nor U1510 (N_1510,N_803,N_1426);
and U1511 (N_1511,N_965,N_821);
and U1512 (N_1512,N_1432,N_952);
xnor U1513 (N_1513,N_1210,N_860);
or U1514 (N_1514,N_903,N_1286);
or U1515 (N_1515,N_832,N_1361);
and U1516 (N_1516,N_1315,N_923);
nor U1517 (N_1517,N_1117,N_1174);
and U1518 (N_1518,N_1312,N_1160);
xor U1519 (N_1519,N_1238,N_817);
xnor U1520 (N_1520,N_1398,N_1070);
nor U1521 (N_1521,N_984,N_1063);
or U1522 (N_1522,N_1412,N_1157);
nand U1523 (N_1523,N_892,N_1438);
or U1524 (N_1524,N_1360,N_1047);
or U1525 (N_1525,N_888,N_874);
and U1526 (N_1526,N_1031,N_766);
nand U1527 (N_1527,N_954,N_1411);
or U1528 (N_1528,N_1491,N_1374);
nor U1529 (N_1529,N_829,N_936);
xor U1530 (N_1530,N_964,N_879);
xor U1531 (N_1531,N_1284,N_949);
nor U1532 (N_1532,N_809,N_1053);
or U1533 (N_1533,N_867,N_988);
and U1534 (N_1534,N_1205,N_950);
xnor U1535 (N_1535,N_801,N_1280);
and U1536 (N_1536,N_768,N_1255);
nand U1537 (N_1537,N_1292,N_1257);
and U1538 (N_1538,N_1377,N_1087);
and U1539 (N_1539,N_939,N_953);
or U1540 (N_1540,N_1145,N_828);
or U1541 (N_1541,N_1215,N_1153);
xor U1542 (N_1542,N_762,N_1239);
and U1543 (N_1543,N_1154,N_1346);
nand U1544 (N_1544,N_922,N_1476);
xnor U1545 (N_1545,N_802,N_1102);
xor U1546 (N_1546,N_1372,N_1109);
nand U1547 (N_1547,N_1427,N_1396);
and U1548 (N_1548,N_855,N_905);
nand U1549 (N_1549,N_1460,N_919);
nand U1550 (N_1550,N_987,N_916);
nand U1551 (N_1551,N_1314,N_1442);
xnor U1552 (N_1552,N_1190,N_1142);
or U1553 (N_1553,N_1482,N_1402);
nand U1554 (N_1554,N_1444,N_887);
and U1555 (N_1555,N_1196,N_1410);
nand U1556 (N_1556,N_1058,N_1199);
xor U1557 (N_1557,N_920,N_1098);
nor U1558 (N_1558,N_1128,N_1005);
nand U1559 (N_1559,N_1177,N_1025);
nand U1560 (N_1560,N_1124,N_1114);
or U1561 (N_1561,N_1089,N_1221);
xor U1562 (N_1562,N_1146,N_1198);
nor U1563 (N_1563,N_1173,N_1450);
nand U1564 (N_1564,N_1038,N_773);
xnor U1565 (N_1565,N_1363,N_1375);
or U1566 (N_1566,N_1197,N_1028);
or U1567 (N_1567,N_1263,N_847);
or U1568 (N_1568,N_1297,N_846);
and U1569 (N_1569,N_883,N_1066);
nor U1570 (N_1570,N_1429,N_932);
nand U1571 (N_1571,N_1464,N_991);
nor U1572 (N_1572,N_1171,N_1493);
or U1573 (N_1573,N_1225,N_951);
nor U1574 (N_1574,N_851,N_1468);
or U1575 (N_1575,N_1104,N_1116);
xor U1576 (N_1576,N_935,N_1399);
nand U1577 (N_1577,N_1243,N_861);
nand U1578 (N_1578,N_1009,N_1191);
nor U1579 (N_1579,N_1162,N_862);
and U1580 (N_1580,N_1144,N_1400);
nor U1581 (N_1581,N_1483,N_1169);
nor U1582 (N_1582,N_1044,N_1336);
xor U1583 (N_1583,N_1338,N_1194);
nor U1584 (N_1584,N_1395,N_871);
nand U1585 (N_1585,N_958,N_1134);
nand U1586 (N_1586,N_1289,N_1248);
and U1587 (N_1587,N_1451,N_799);
nor U1588 (N_1588,N_979,N_1441);
nor U1589 (N_1589,N_878,N_782);
nor U1590 (N_1590,N_1165,N_1081);
nor U1591 (N_1591,N_1164,N_1040);
nor U1592 (N_1592,N_752,N_1206);
or U1593 (N_1593,N_1224,N_1309);
nand U1594 (N_1594,N_1329,N_1497);
or U1595 (N_1595,N_1492,N_1016);
xor U1596 (N_1596,N_1094,N_1187);
nor U1597 (N_1597,N_841,N_859);
xnor U1598 (N_1598,N_800,N_1203);
nand U1599 (N_1599,N_1136,N_1282);
and U1600 (N_1600,N_1074,N_764);
or U1601 (N_1601,N_1151,N_1027);
and U1602 (N_1602,N_1419,N_1328);
xor U1603 (N_1603,N_941,N_1310);
nand U1604 (N_1604,N_1179,N_1068);
nand U1605 (N_1605,N_854,N_823);
or U1606 (N_1606,N_1277,N_822);
and U1607 (N_1607,N_1307,N_995);
and U1608 (N_1608,N_1489,N_1091);
or U1609 (N_1609,N_1260,N_1007);
and U1610 (N_1610,N_1067,N_1075);
nand U1611 (N_1611,N_1368,N_960);
xnor U1612 (N_1612,N_818,N_787);
xor U1613 (N_1613,N_1456,N_1204);
xnor U1614 (N_1614,N_1088,N_918);
nor U1615 (N_1615,N_842,N_1234);
and U1616 (N_1616,N_1457,N_908);
or U1617 (N_1617,N_772,N_804);
nor U1618 (N_1618,N_1084,N_1235);
or U1619 (N_1619,N_982,N_778);
xnor U1620 (N_1620,N_1101,N_1388);
nand U1621 (N_1621,N_912,N_869);
or U1622 (N_1622,N_1061,N_843);
nand U1623 (N_1623,N_1259,N_776);
and U1624 (N_1624,N_1471,N_1200);
and U1625 (N_1625,N_1474,N_1334);
nor U1626 (N_1626,N_980,N_1010);
and U1627 (N_1627,N_1317,N_1214);
xor U1628 (N_1628,N_994,N_754);
and U1629 (N_1629,N_1452,N_1106);
nor U1630 (N_1630,N_1454,N_1046);
nand U1631 (N_1631,N_1390,N_1343);
or U1632 (N_1632,N_1271,N_1041);
or U1633 (N_1633,N_1150,N_884);
nand U1634 (N_1634,N_1030,N_1032);
xor U1635 (N_1635,N_1062,N_877);
xnor U1636 (N_1636,N_1222,N_895);
xnor U1637 (N_1637,N_1125,N_1287);
and U1638 (N_1638,N_1416,N_989);
and U1639 (N_1639,N_788,N_1405);
nor U1640 (N_1640,N_1281,N_1472);
nand U1641 (N_1641,N_898,N_845);
nand U1642 (N_1642,N_1135,N_956);
xor U1643 (N_1643,N_1488,N_1440);
nand U1644 (N_1644,N_1261,N_835);
and U1645 (N_1645,N_881,N_1325);
nand U1646 (N_1646,N_1278,N_1433);
and U1647 (N_1647,N_986,N_1035);
xnor U1648 (N_1648,N_1288,N_990);
and U1649 (N_1649,N_1496,N_962);
nor U1650 (N_1650,N_1176,N_1274);
and U1651 (N_1651,N_1100,N_819);
and U1652 (N_1652,N_1244,N_1409);
nand U1653 (N_1653,N_1423,N_1342);
xnor U1654 (N_1654,N_1002,N_1455);
nand U1655 (N_1655,N_1226,N_793);
nor U1656 (N_1656,N_807,N_1026);
or U1657 (N_1657,N_947,N_1355);
nand U1658 (N_1658,N_1024,N_1495);
or U1659 (N_1659,N_1401,N_1439);
xor U1660 (N_1660,N_1323,N_1283);
or U1661 (N_1661,N_1479,N_902);
nand U1662 (N_1662,N_1186,N_1121);
and U1663 (N_1663,N_1163,N_955);
xor U1664 (N_1664,N_929,N_1189);
nor U1665 (N_1665,N_1275,N_1347);
xor U1666 (N_1666,N_1242,N_1348);
nand U1667 (N_1667,N_978,N_996);
xor U1668 (N_1668,N_1233,N_780);
and U1669 (N_1669,N_1172,N_1216);
xor U1670 (N_1670,N_1111,N_1126);
nor U1671 (N_1671,N_1227,N_767);
and U1672 (N_1672,N_993,N_1185);
nand U1673 (N_1673,N_1080,N_901);
or U1674 (N_1674,N_1267,N_1324);
or U1675 (N_1675,N_1004,N_1385);
and U1676 (N_1676,N_1059,N_1078);
and U1677 (N_1677,N_1076,N_1108);
nand U1678 (N_1678,N_792,N_981);
nand U1679 (N_1679,N_1060,N_1137);
xnor U1680 (N_1680,N_1015,N_1300);
or U1681 (N_1681,N_1000,N_1331);
and U1682 (N_1682,N_1332,N_1453);
nand U1683 (N_1683,N_1487,N_1321);
nor U1684 (N_1684,N_863,N_1037);
xor U1685 (N_1685,N_1384,N_870);
or U1686 (N_1686,N_824,N_839);
and U1687 (N_1687,N_1178,N_1301);
and U1688 (N_1688,N_1379,N_774);
and U1689 (N_1689,N_1320,N_1333);
nor U1690 (N_1690,N_858,N_928);
nand U1691 (N_1691,N_1480,N_1490);
nand U1692 (N_1692,N_910,N_868);
and U1693 (N_1693,N_1129,N_825);
and U1694 (N_1694,N_1090,N_938);
and U1695 (N_1695,N_1220,N_1478);
xnor U1696 (N_1696,N_1017,N_1443);
and U1697 (N_1697,N_1430,N_1449);
nor U1698 (N_1698,N_1036,N_794);
xor U1699 (N_1699,N_1152,N_970);
or U1700 (N_1700,N_1296,N_1014);
xnor U1701 (N_1701,N_1254,N_1435);
or U1702 (N_1702,N_945,N_805);
and U1703 (N_1703,N_1358,N_827);
xnor U1704 (N_1704,N_1229,N_853);
and U1705 (N_1705,N_913,N_810);
xor U1706 (N_1706,N_992,N_1417);
and U1707 (N_1707,N_831,N_1459);
xor U1708 (N_1708,N_1158,N_1258);
and U1709 (N_1709,N_1484,N_999);
and U1710 (N_1710,N_1276,N_760);
xor U1711 (N_1711,N_1170,N_1079);
nor U1712 (N_1712,N_930,N_915);
nand U1713 (N_1713,N_1241,N_937);
nor U1714 (N_1714,N_833,N_789);
or U1715 (N_1715,N_972,N_1291);
nand U1716 (N_1716,N_1404,N_1130);
xnor U1717 (N_1717,N_1359,N_1064);
or U1718 (N_1718,N_961,N_1056);
nand U1719 (N_1719,N_806,N_1393);
or U1720 (N_1720,N_1118,N_756);
xnor U1721 (N_1721,N_872,N_1308);
nand U1722 (N_1722,N_1351,N_1103);
or U1723 (N_1723,N_779,N_897);
xnor U1724 (N_1724,N_1223,N_1295);
nand U1725 (N_1725,N_816,N_834);
and U1726 (N_1726,N_1008,N_1467);
nand U1727 (N_1727,N_891,N_1085);
nor U1728 (N_1728,N_943,N_1202);
and U1729 (N_1729,N_1183,N_933);
xnor U1730 (N_1730,N_866,N_797);
nand U1731 (N_1731,N_808,N_1231);
and U1732 (N_1732,N_894,N_1113);
and U1733 (N_1733,N_944,N_1373);
xor U1734 (N_1734,N_1132,N_1119);
and U1735 (N_1735,N_1049,N_1378);
and U1736 (N_1736,N_777,N_1264);
xnor U1737 (N_1737,N_1473,N_1311);
and U1738 (N_1738,N_1156,N_957);
xor U1739 (N_1739,N_909,N_1122);
or U1740 (N_1740,N_1391,N_759);
xor U1741 (N_1741,N_857,N_1318);
xnor U1742 (N_1742,N_1270,N_1376);
and U1743 (N_1743,N_885,N_1462);
or U1744 (N_1744,N_927,N_1256);
nor U1745 (N_1745,N_1445,N_1465);
nor U1746 (N_1746,N_865,N_790);
or U1747 (N_1747,N_1394,N_849);
xnor U1748 (N_1748,N_983,N_1237);
nor U1749 (N_1749,N_1072,N_1349);
nor U1750 (N_1750,N_1131,N_1249);
xor U1751 (N_1751,N_966,N_1065);
xnor U1752 (N_1752,N_1340,N_1236);
and U1753 (N_1753,N_769,N_848);
or U1754 (N_1754,N_914,N_1356);
nor U1755 (N_1755,N_934,N_820);
nand U1756 (N_1756,N_1413,N_1246);
and U1757 (N_1757,N_1011,N_1149);
and U1758 (N_1758,N_1043,N_977);
and U1759 (N_1759,N_921,N_1357);
nand U1760 (N_1760,N_1212,N_1327);
nand U1761 (N_1761,N_924,N_1364);
xnor U1762 (N_1762,N_967,N_1322);
or U1763 (N_1763,N_1201,N_765);
nor U1764 (N_1764,N_1230,N_1175);
nor U1765 (N_1765,N_1167,N_1217);
or U1766 (N_1766,N_1304,N_1252);
nor U1767 (N_1767,N_1208,N_813);
nor U1768 (N_1768,N_1339,N_836);
xnor U1769 (N_1769,N_890,N_1069);
and U1770 (N_1770,N_837,N_1034);
and U1771 (N_1771,N_864,N_1184);
nor U1772 (N_1772,N_1019,N_911);
nand U1773 (N_1773,N_1245,N_1469);
and U1774 (N_1774,N_1481,N_770);
xor U1775 (N_1775,N_1168,N_791);
nand U1776 (N_1776,N_1071,N_1120);
nand U1777 (N_1777,N_876,N_1253);
nor U1778 (N_1778,N_1494,N_751);
nor U1779 (N_1779,N_785,N_1437);
xor U1780 (N_1780,N_1166,N_907);
nor U1781 (N_1781,N_1247,N_1485);
nand U1782 (N_1782,N_1422,N_1029);
xor U1783 (N_1783,N_1048,N_1285);
nand U1784 (N_1784,N_761,N_1268);
xnor U1785 (N_1785,N_1326,N_844);
nand U1786 (N_1786,N_758,N_1054);
or U1787 (N_1787,N_1362,N_889);
nor U1788 (N_1788,N_1209,N_931);
nand U1789 (N_1789,N_880,N_1023);
nor U1790 (N_1790,N_1018,N_1182);
xor U1791 (N_1791,N_1434,N_753);
and U1792 (N_1792,N_1097,N_899);
or U1793 (N_1793,N_1380,N_1415);
nor U1794 (N_1794,N_1279,N_1093);
nor U1795 (N_1795,N_1387,N_850);
xnor U1796 (N_1796,N_1448,N_1050);
and U1797 (N_1797,N_1051,N_1045);
or U1798 (N_1798,N_1350,N_1306);
or U1799 (N_1799,N_750,N_997);
or U1800 (N_1800,N_1003,N_975);
xor U1801 (N_1801,N_1188,N_873);
or U1802 (N_1802,N_904,N_1436);
and U1803 (N_1803,N_1302,N_796);
and U1804 (N_1804,N_968,N_1013);
nand U1805 (N_1805,N_1266,N_1218);
and U1806 (N_1806,N_893,N_1341);
nand U1807 (N_1807,N_1139,N_1055);
nor U1808 (N_1808,N_1293,N_830);
or U1809 (N_1809,N_1073,N_1316);
and U1810 (N_1810,N_815,N_1475);
or U1811 (N_1811,N_1133,N_1499);
and U1812 (N_1812,N_1159,N_1039);
nand U1813 (N_1813,N_1353,N_1446);
nand U1814 (N_1814,N_917,N_1141);
xnor U1815 (N_1815,N_1033,N_1107);
xnor U1816 (N_1816,N_1207,N_925);
or U1817 (N_1817,N_826,N_1265);
nand U1818 (N_1818,N_1408,N_1352);
nand U1819 (N_1819,N_976,N_1250);
nand U1820 (N_1820,N_1290,N_1335);
or U1821 (N_1821,N_1228,N_798);
nand U1822 (N_1822,N_1319,N_1305);
nand U1823 (N_1823,N_1365,N_1077);
xor U1824 (N_1824,N_1458,N_1299);
or U1825 (N_1825,N_856,N_1330);
nor U1826 (N_1826,N_1181,N_882);
or U1827 (N_1827,N_1345,N_1082);
xor U1828 (N_1828,N_1382,N_1269);
nand U1829 (N_1829,N_814,N_1123);
or U1830 (N_1830,N_1294,N_1470);
nor U1831 (N_1831,N_1042,N_812);
nand U1832 (N_1832,N_1192,N_1406);
nor U1833 (N_1833,N_1105,N_1195);
nor U1834 (N_1834,N_1112,N_1147);
or U1835 (N_1835,N_1407,N_1232);
xor U1836 (N_1836,N_781,N_1052);
or U1837 (N_1837,N_926,N_1421);
or U1838 (N_1838,N_784,N_1303);
or U1839 (N_1839,N_755,N_1211);
and U1840 (N_1840,N_838,N_1012);
nand U1841 (N_1841,N_886,N_1096);
xor U1842 (N_1842,N_1397,N_1369);
nand U1843 (N_1843,N_1022,N_1001);
and U1844 (N_1844,N_1180,N_1092);
or U1845 (N_1845,N_1463,N_786);
xor U1846 (N_1846,N_985,N_1477);
nor U1847 (N_1847,N_1193,N_940);
xnor U1848 (N_1848,N_1431,N_1354);
nand U1849 (N_1849,N_1461,N_1115);
and U1850 (N_1850,N_1420,N_1213);
or U1851 (N_1851,N_1344,N_1020);
nor U1852 (N_1852,N_852,N_1251);
and U1853 (N_1853,N_775,N_795);
xor U1854 (N_1854,N_948,N_1086);
nand U1855 (N_1855,N_1418,N_1414);
nand U1856 (N_1856,N_896,N_973);
or U1857 (N_1857,N_1240,N_1273);
or U1858 (N_1858,N_1298,N_1272);
nand U1859 (N_1859,N_763,N_1161);
nor U1860 (N_1860,N_906,N_959);
xor U1861 (N_1861,N_946,N_963);
nand U1862 (N_1862,N_811,N_1057);
nor U1863 (N_1863,N_1127,N_1371);
nor U1864 (N_1864,N_1392,N_1099);
and U1865 (N_1865,N_900,N_1447);
or U1866 (N_1866,N_1425,N_1110);
nand U1867 (N_1867,N_1140,N_1486);
nor U1868 (N_1868,N_1370,N_875);
nand U1869 (N_1869,N_1219,N_1403);
or U1870 (N_1870,N_974,N_771);
nand U1871 (N_1871,N_1143,N_1095);
nor U1872 (N_1872,N_969,N_1021);
xor U1873 (N_1873,N_1428,N_1383);
nor U1874 (N_1874,N_840,N_942);
or U1875 (N_1875,N_843,N_912);
nand U1876 (N_1876,N_1006,N_1022);
nor U1877 (N_1877,N_1226,N_1033);
xnor U1878 (N_1878,N_1013,N_852);
nand U1879 (N_1879,N_941,N_1399);
nor U1880 (N_1880,N_1013,N_1399);
and U1881 (N_1881,N_848,N_1107);
nand U1882 (N_1882,N_1285,N_1185);
xor U1883 (N_1883,N_1156,N_1058);
nor U1884 (N_1884,N_1376,N_1399);
or U1885 (N_1885,N_1067,N_1307);
nand U1886 (N_1886,N_1415,N_950);
nand U1887 (N_1887,N_1268,N_1167);
xor U1888 (N_1888,N_1289,N_1447);
xnor U1889 (N_1889,N_1189,N_1339);
or U1890 (N_1890,N_1019,N_995);
nor U1891 (N_1891,N_1334,N_848);
and U1892 (N_1892,N_1062,N_1465);
xnor U1893 (N_1893,N_1135,N_1490);
nor U1894 (N_1894,N_1406,N_1041);
xor U1895 (N_1895,N_1144,N_890);
nor U1896 (N_1896,N_865,N_1060);
xnor U1897 (N_1897,N_1139,N_1220);
or U1898 (N_1898,N_846,N_1174);
xnor U1899 (N_1899,N_1298,N_966);
and U1900 (N_1900,N_1066,N_996);
or U1901 (N_1901,N_785,N_1084);
nor U1902 (N_1902,N_1277,N_1186);
xor U1903 (N_1903,N_1050,N_1033);
xnor U1904 (N_1904,N_1201,N_1431);
nor U1905 (N_1905,N_1104,N_1175);
or U1906 (N_1906,N_1029,N_1103);
xnor U1907 (N_1907,N_1493,N_1366);
nand U1908 (N_1908,N_1449,N_1490);
or U1909 (N_1909,N_962,N_1169);
or U1910 (N_1910,N_871,N_786);
nor U1911 (N_1911,N_835,N_1440);
or U1912 (N_1912,N_1406,N_1214);
nand U1913 (N_1913,N_1181,N_985);
nand U1914 (N_1914,N_1223,N_754);
or U1915 (N_1915,N_1237,N_1236);
and U1916 (N_1916,N_1377,N_1120);
or U1917 (N_1917,N_802,N_1026);
and U1918 (N_1918,N_875,N_833);
and U1919 (N_1919,N_1156,N_1307);
or U1920 (N_1920,N_1219,N_1033);
and U1921 (N_1921,N_1019,N_1347);
and U1922 (N_1922,N_1154,N_937);
nor U1923 (N_1923,N_922,N_1345);
nand U1924 (N_1924,N_769,N_912);
nor U1925 (N_1925,N_869,N_1328);
nand U1926 (N_1926,N_863,N_1009);
or U1927 (N_1927,N_1489,N_1328);
xnor U1928 (N_1928,N_1231,N_1420);
or U1929 (N_1929,N_821,N_1493);
xnor U1930 (N_1930,N_1339,N_1248);
nand U1931 (N_1931,N_1270,N_1489);
and U1932 (N_1932,N_931,N_1382);
and U1933 (N_1933,N_1146,N_922);
nor U1934 (N_1934,N_1292,N_1076);
nand U1935 (N_1935,N_1281,N_1280);
and U1936 (N_1936,N_1056,N_1452);
xnor U1937 (N_1937,N_1471,N_955);
xnor U1938 (N_1938,N_1014,N_1127);
nand U1939 (N_1939,N_1110,N_938);
or U1940 (N_1940,N_1080,N_868);
nand U1941 (N_1941,N_754,N_1310);
nor U1942 (N_1942,N_1094,N_773);
or U1943 (N_1943,N_882,N_820);
nor U1944 (N_1944,N_792,N_1448);
or U1945 (N_1945,N_1118,N_1009);
nand U1946 (N_1946,N_852,N_1020);
xnor U1947 (N_1947,N_1441,N_1410);
and U1948 (N_1948,N_1082,N_1068);
nor U1949 (N_1949,N_1224,N_1411);
nor U1950 (N_1950,N_976,N_968);
xor U1951 (N_1951,N_893,N_1485);
nor U1952 (N_1952,N_1061,N_952);
xor U1953 (N_1953,N_929,N_1360);
nor U1954 (N_1954,N_839,N_942);
nor U1955 (N_1955,N_1499,N_1147);
and U1956 (N_1956,N_1110,N_816);
nand U1957 (N_1957,N_834,N_783);
nor U1958 (N_1958,N_907,N_862);
nand U1959 (N_1959,N_1496,N_1320);
nor U1960 (N_1960,N_764,N_828);
xor U1961 (N_1961,N_918,N_1366);
xnor U1962 (N_1962,N_1067,N_936);
xnor U1963 (N_1963,N_1115,N_1359);
nand U1964 (N_1964,N_1134,N_1072);
and U1965 (N_1965,N_1308,N_1054);
and U1966 (N_1966,N_1437,N_1467);
or U1967 (N_1967,N_1136,N_760);
nand U1968 (N_1968,N_1058,N_1197);
and U1969 (N_1969,N_1061,N_1067);
xnor U1970 (N_1970,N_1270,N_1190);
xnor U1971 (N_1971,N_1436,N_1240);
nor U1972 (N_1972,N_1459,N_1014);
and U1973 (N_1973,N_1061,N_1000);
nand U1974 (N_1974,N_1176,N_1245);
xnor U1975 (N_1975,N_1296,N_1141);
nor U1976 (N_1976,N_1352,N_1288);
xor U1977 (N_1977,N_1294,N_785);
or U1978 (N_1978,N_1304,N_784);
nor U1979 (N_1979,N_1178,N_967);
nor U1980 (N_1980,N_1045,N_1031);
and U1981 (N_1981,N_1171,N_1254);
or U1982 (N_1982,N_1357,N_897);
nor U1983 (N_1983,N_1440,N_1258);
nand U1984 (N_1984,N_1071,N_847);
nor U1985 (N_1985,N_1138,N_999);
and U1986 (N_1986,N_933,N_963);
nor U1987 (N_1987,N_759,N_1219);
nor U1988 (N_1988,N_1414,N_1365);
and U1989 (N_1989,N_924,N_1201);
and U1990 (N_1990,N_1477,N_1146);
nor U1991 (N_1991,N_910,N_799);
xor U1992 (N_1992,N_797,N_1352);
nand U1993 (N_1993,N_1158,N_1054);
nand U1994 (N_1994,N_1034,N_1471);
and U1995 (N_1995,N_1342,N_1106);
and U1996 (N_1996,N_809,N_1441);
and U1997 (N_1997,N_1141,N_1217);
xnor U1998 (N_1998,N_750,N_1026);
nand U1999 (N_1999,N_1040,N_760);
xor U2000 (N_2000,N_1448,N_1463);
nand U2001 (N_2001,N_1076,N_1214);
or U2002 (N_2002,N_1152,N_965);
nor U2003 (N_2003,N_1038,N_1304);
nor U2004 (N_2004,N_1105,N_1284);
and U2005 (N_2005,N_1387,N_1014);
or U2006 (N_2006,N_1392,N_1057);
nor U2007 (N_2007,N_904,N_885);
nor U2008 (N_2008,N_1167,N_814);
and U2009 (N_2009,N_1325,N_1134);
xor U2010 (N_2010,N_818,N_959);
or U2011 (N_2011,N_996,N_761);
or U2012 (N_2012,N_911,N_1392);
and U2013 (N_2013,N_1154,N_1445);
xor U2014 (N_2014,N_872,N_1340);
xnor U2015 (N_2015,N_897,N_902);
nor U2016 (N_2016,N_765,N_1123);
nand U2017 (N_2017,N_1051,N_1375);
xor U2018 (N_2018,N_1163,N_852);
nor U2019 (N_2019,N_1322,N_754);
or U2020 (N_2020,N_852,N_897);
xor U2021 (N_2021,N_1398,N_1474);
and U2022 (N_2022,N_1134,N_912);
nor U2023 (N_2023,N_1208,N_1414);
xor U2024 (N_2024,N_1243,N_1247);
nand U2025 (N_2025,N_1286,N_1385);
or U2026 (N_2026,N_818,N_1321);
nand U2027 (N_2027,N_1425,N_1346);
nor U2028 (N_2028,N_1012,N_1228);
or U2029 (N_2029,N_861,N_1450);
nand U2030 (N_2030,N_772,N_1093);
xor U2031 (N_2031,N_1289,N_1292);
nor U2032 (N_2032,N_1211,N_769);
xnor U2033 (N_2033,N_1453,N_1477);
nor U2034 (N_2034,N_1307,N_911);
and U2035 (N_2035,N_1262,N_1348);
or U2036 (N_2036,N_1264,N_1155);
or U2037 (N_2037,N_1350,N_1172);
nor U2038 (N_2038,N_907,N_1482);
nand U2039 (N_2039,N_807,N_1406);
nor U2040 (N_2040,N_1429,N_787);
or U2041 (N_2041,N_1484,N_1079);
xnor U2042 (N_2042,N_1338,N_1400);
nor U2043 (N_2043,N_994,N_1459);
and U2044 (N_2044,N_997,N_1367);
nor U2045 (N_2045,N_977,N_1187);
and U2046 (N_2046,N_961,N_1353);
or U2047 (N_2047,N_922,N_1090);
or U2048 (N_2048,N_1435,N_1006);
and U2049 (N_2049,N_1249,N_1455);
or U2050 (N_2050,N_955,N_1107);
or U2051 (N_2051,N_932,N_1335);
or U2052 (N_2052,N_1123,N_1233);
and U2053 (N_2053,N_886,N_1454);
or U2054 (N_2054,N_874,N_1131);
nand U2055 (N_2055,N_802,N_800);
nand U2056 (N_2056,N_1375,N_1010);
xor U2057 (N_2057,N_751,N_905);
xor U2058 (N_2058,N_1044,N_1316);
and U2059 (N_2059,N_1288,N_1234);
and U2060 (N_2060,N_823,N_1063);
nor U2061 (N_2061,N_1205,N_786);
or U2062 (N_2062,N_1347,N_1285);
xnor U2063 (N_2063,N_1138,N_1210);
nor U2064 (N_2064,N_1271,N_1069);
nor U2065 (N_2065,N_1447,N_1305);
nand U2066 (N_2066,N_1352,N_1028);
and U2067 (N_2067,N_1439,N_1138);
nor U2068 (N_2068,N_1391,N_1481);
xnor U2069 (N_2069,N_986,N_1447);
nand U2070 (N_2070,N_1134,N_897);
and U2071 (N_2071,N_1429,N_866);
or U2072 (N_2072,N_1289,N_842);
nand U2073 (N_2073,N_1237,N_1386);
nand U2074 (N_2074,N_1213,N_1293);
nand U2075 (N_2075,N_1324,N_1257);
and U2076 (N_2076,N_1255,N_1287);
and U2077 (N_2077,N_1380,N_1366);
or U2078 (N_2078,N_1234,N_1438);
and U2079 (N_2079,N_1055,N_1456);
nand U2080 (N_2080,N_1108,N_1179);
and U2081 (N_2081,N_844,N_1265);
nor U2082 (N_2082,N_1280,N_1248);
xnor U2083 (N_2083,N_1335,N_1136);
or U2084 (N_2084,N_1067,N_895);
and U2085 (N_2085,N_990,N_1041);
or U2086 (N_2086,N_1102,N_1068);
nor U2087 (N_2087,N_900,N_1147);
or U2088 (N_2088,N_1175,N_945);
or U2089 (N_2089,N_1416,N_1492);
and U2090 (N_2090,N_1032,N_1443);
and U2091 (N_2091,N_790,N_1220);
xnor U2092 (N_2092,N_1305,N_1056);
nand U2093 (N_2093,N_1433,N_1392);
nand U2094 (N_2094,N_1464,N_952);
xor U2095 (N_2095,N_1073,N_1026);
or U2096 (N_2096,N_1241,N_1220);
and U2097 (N_2097,N_1405,N_1482);
and U2098 (N_2098,N_1128,N_1373);
nor U2099 (N_2099,N_1285,N_966);
or U2100 (N_2100,N_1173,N_1177);
nor U2101 (N_2101,N_1488,N_1218);
xor U2102 (N_2102,N_896,N_1289);
nand U2103 (N_2103,N_756,N_844);
nor U2104 (N_2104,N_873,N_1164);
xnor U2105 (N_2105,N_1059,N_1125);
or U2106 (N_2106,N_1425,N_843);
nand U2107 (N_2107,N_1159,N_1300);
nand U2108 (N_2108,N_976,N_875);
or U2109 (N_2109,N_807,N_860);
xor U2110 (N_2110,N_936,N_1375);
or U2111 (N_2111,N_1417,N_1411);
nand U2112 (N_2112,N_1076,N_1478);
nand U2113 (N_2113,N_1050,N_1091);
xnor U2114 (N_2114,N_991,N_1383);
xnor U2115 (N_2115,N_856,N_1154);
nand U2116 (N_2116,N_1002,N_904);
or U2117 (N_2117,N_1395,N_953);
nor U2118 (N_2118,N_830,N_1173);
xnor U2119 (N_2119,N_755,N_1344);
or U2120 (N_2120,N_1180,N_1134);
xnor U2121 (N_2121,N_1490,N_898);
nand U2122 (N_2122,N_1184,N_1165);
xor U2123 (N_2123,N_1137,N_1401);
nor U2124 (N_2124,N_1040,N_820);
nand U2125 (N_2125,N_1413,N_900);
or U2126 (N_2126,N_1498,N_1491);
and U2127 (N_2127,N_1201,N_1370);
xor U2128 (N_2128,N_861,N_1490);
and U2129 (N_2129,N_1100,N_1125);
and U2130 (N_2130,N_938,N_1466);
or U2131 (N_2131,N_1066,N_1379);
nand U2132 (N_2132,N_1185,N_938);
nand U2133 (N_2133,N_776,N_1073);
nor U2134 (N_2134,N_927,N_1103);
and U2135 (N_2135,N_836,N_960);
or U2136 (N_2136,N_854,N_1364);
xor U2137 (N_2137,N_1347,N_1382);
nand U2138 (N_2138,N_1470,N_1141);
and U2139 (N_2139,N_977,N_1095);
or U2140 (N_2140,N_1037,N_940);
or U2141 (N_2141,N_1053,N_1252);
and U2142 (N_2142,N_944,N_1424);
or U2143 (N_2143,N_1031,N_1370);
xor U2144 (N_2144,N_1271,N_1157);
or U2145 (N_2145,N_1076,N_1470);
xnor U2146 (N_2146,N_759,N_1071);
xor U2147 (N_2147,N_1059,N_998);
nand U2148 (N_2148,N_952,N_1467);
nor U2149 (N_2149,N_873,N_1081);
xnor U2150 (N_2150,N_1373,N_817);
xor U2151 (N_2151,N_997,N_776);
or U2152 (N_2152,N_772,N_868);
nand U2153 (N_2153,N_1343,N_1267);
and U2154 (N_2154,N_860,N_859);
and U2155 (N_2155,N_819,N_970);
nand U2156 (N_2156,N_921,N_1179);
or U2157 (N_2157,N_1165,N_1384);
xor U2158 (N_2158,N_979,N_981);
or U2159 (N_2159,N_1451,N_1393);
xnor U2160 (N_2160,N_755,N_1047);
xnor U2161 (N_2161,N_1190,N_1188);
or U2162 (N_2162,N_933,N_1361);
nor U2163 (N_2163,N_1343,N_1309);
xnor U2164 (N_2164,N_1143,N_1179);
and U2165 (N_2165,N_780,N_1337);
nor U2166 (N_2166,N_822,N_1092);
nor U2167 (N_2167,N_756,N_1350);
nand U2168 (N_2168,N_788,N_1384);
xor U2169 (N_2169,N_1195,N_1322);
nand U2170 (N_2170,N_1038,N_988);
nand U2171 (N_2171,N_1345,N_1201);
or U2172 (N_2172,N_1060,N_1340);
and U2173 (N_2173,N_1140,N_753);
or U2174 (N_2174,N_989,N_1213);
nand U2175 (N_2175,N_961,N_787);
xnor U2176 (N_2176,N_1280,N_847);
xnor U2177 (N_2177,N_884,N_980);
and U2178 (N_2178,N_1090,N_1359);
nor U2179 (N_2179,N_801,N_1214);
or U2180 (N_2180,N_1485,N_782);
xor U2181 (N_2181,N_1265,N_1406);
or U2182 (N_2182,N_1374,N_772);
xnor U2183 (N_2183,N_834,N_1422);
and U2184 (N_2184,N_998,N_797);
nor U2185 (N_2185,N_847,N_771);
or U2186 (N_2186,N_1399,N_1416);
nor U2187 (N_2187,N_960,N_1197);
xnor U2188 (N_2188,N_1227,N_866);
and U2189 (N_2189,N_1319,N_931);
xnor U2190 (N_2190,N_1333,N_1150);
nor U2191 (N_2191,N_828,N_1309);
or U2192 (N_2192,N_1171,N_784);
xnor U2193 (N_2193,N_1440,N_998);
nor U2194 (N_2194,N_1344,N_888);
xnor U2195 (N_2195,N_1280,N_1407);
nor U2196 (N_2196,N_1286,N_1238);
and U2197 (N_2197,N_1128,N_1085);
nor U2198 (N_2198,N_1123,N_776);
nor U2199 (N_2199,N_921,N_1225);
or U2200 (N_2200,N_1455,N_1400);
xnor U2201 (N_2201,N_1410,N_1250);
nor U2202 (N_2202,N_979,N_1099);
nor U2203 (N_2203,N_1010,N_1271);
or U2204 (N_2204,N_830,N_1322);
nand U2205 (N_2205,N_1399,N_778);
or U2206 (N_2206,N_1039,N_1080);
or U2207 (N_2207,N_782,N_758);
xnor U2208 (N_2208,N_1057,N_779);
nand U2209 (N_2209,N_945,N_860);
nor U2210 (N_2210,N_1175,N_1033);
nor U2211 (N_2211,N_946,N_1356);
xnor U2212 (N_2212,N_833,N_1155);
or U2213 (N_2213,N_843,N_785);
or U2214 (N_2214,N_1457,N_1113);
nor U2215 (N_2215,N_820,N_1260);
and U2216 (N_2216,N_1323,N_843);
and U2217 (N_2217,N_809,N_1178);
nand U2218 (N_2218,N_922,N_1424);
and U2219 (N_2219,N_1301,N_1243);
xor U2220 (N_2220,N_1207,N_1370);
or U2221 (N_2221,N_853,N_1365);
xnor U2222 (N_2222,N_1188,N_1052);
and U2223 (N_2223,N_1227,N_791);
xor U2224 (N_2224,N_1097,N_965);
xor U2225 (N_2225,N_1069,N_1467);
and U2226 (N_2226,N_1143,N_772);
or U2227 (N_2227,N_975,N_846);
or U2228 (N_2228,N_1015,N_1271);
nor U2229 (N_2229,N_985,N_765);
or U2230 (N_2230,N_1136,N_1141);
xnor U2231 (N_2231,N_1354,N_1276);
or U2232 (N_2232,N_1319,N_1083);
nand U2233 (N_2233,N_1069,N_1134);
xnor U2234 (N_2234,N_1171,N_786);
or U2235 (N_2235,N_955,N_1329);
xnor U2236 (N_2236,N_1458,N_833);
nor U2237 (N_2237,N_1020,N_776);
nand U2238 (N_2238,N_1419,N_1044);
and U2239 (N_2239,N_1040,N_1496);
nand U2240 (N_2240,N_800,N_1487);
nand U2241 (N_2241,N_1437,N_1473);
xnor U2242 (N_2242,N_1033,N_1312);
xor U2243 (N_2243,N_772,N_1249);
and U2244 (N_2244,N_1492,N_1342);
xor U2245 (N_2245,N_1189,N_842);
and U2246 (N_2246,N_1474,N_877);
and U2247 (N_2247,N_766,N_802);
and U2248 (N_2248,N_1270,N_880);
or U2249 (N_2249,N_829,N_1005);
nand U2250 (N_2250,N_1646,N_2080);
and U2251 (N_2251,N_2098,N_1848);
nor U2252 (N_2252,N_1862,N_1523);
nor U2253 (N_2253,N_2018,N_1503);
xnor U2254 (N_2254,N_1795,N_2115);
nand U2255 (N_2255,N_1650,N_1853);
and U2256 (N_2256,N_1543,N_2203);
nor U2257 (N_2257,N_1665,N_1689);
or U2258 (N_2258,N_1778,N_1831);
xor U2259 (N_2259,N_1903,N_1547);
and U2260 (N_2260,N_1579,N_2228);
or U2261 (N_2261,N_1866,N_1777);
or U2262 (N_2262,N_1633,N_2200);
nand U2263 (N_2263,N_2027,N_1983);
nand U2264 (N_2264,N_2186,N_1590);
nor U2265 (N_2265,N_2248,N_1695);
nand U2266 (N_2266,N_2044,N_2064);
nand U2267 (N_2267,N_2007,N_1905);
xnor U2268 (N_2268,N_1554,N_1673);
nor U2269 (N_2269,N_1643,N_2135);
and U2270 (N_2270,N_2198,N_2218);
or U2271 (N_2271,N_2170,N_2013);
nor U2272 (N_2272,N_1892,N_1515);
and U2273 (N_2273,N_2028,N_1992);
xor U2274 (N_2274,N_1644,N_1782);
nor U2275 (N_2275,N_1698,N_1833);
or U2276 (N_2276,N_1636,N_2168);
and U2277 (N_2277,N_2059,N_1685);
or U2278 (N_2278,N_1790,N_1712);
nor U2279 (N_2279,N_1530,N_1655);
nor U2280 (N_2280,N_1700,N_1789);
or U2281 (N_2281,N_1787,N_2081);
and U2282 (N_2282,N_1599,N_1568);
or U2283 (N_2283,N_1508,N_1522);
nand U2284 (N_2284,N_1708,N_1783);
or U2285 (N_2285,N_1950,N_1731);
nor U2286 (N_2286,N_1813,N_2237);
or U2287 (N_2287,N_2026,N_2214);
or U2288 (N_2288,N_1607,N_1762);
xnor U2289 (N_2289,N_2210,N_1760);
xnor U2290 (N_2290,N_1586,N_1948);
nor U2291 (N_2291,N_1742,N_1781);
nand U2292 (N_2292,N_1583,N_1682);
xor U2293 (N_2293,N_2223,N_1964);
and U2294 (N_2294,N_1951,N_1668);
nand U2295 (N_2295,N_1516,N_1737);
xnor U2296 (N_2296,N_1580,N_1811);
or U2297 (N_2297,N_2088,N_1563);
nand U2298 (N_2298,N_1854,N_1672);
or U2299 (N_2299,N_1872,N_1574);
nor U2300 (N_2300,N_2151,N_2085);
and U2301 (N_2301,N_1880,N_2144);
xnor U2302 (N_2302,N_1691,N_2153);
nand U2303 (N_2303,N_2131,N_1722);
and U2304 (N_2304,N_2076,N_2101);
or U2305 (N_2305,N_1955,N_1770);
xor U2306 (N_2306,N_2053,N_1775);
nor U2307 (N_2307,N_2208,N_1727);
nor U2308 (N_2308,N_2147,N_1603);
xor U2309 (N_2309,N_2244,N_1578);
xnor U2310 (N_2310,N_1832,N_1640);
or U2311 (N_2311,N_2219,N_1944);
xor U2312 (N_2312,N_1763,N_1843);
or U2313 (N_2313,N_2104,N_2241);
nand U2314 (N_2314,N_1864,N_1834);
nor U2315 (N_2315,N_1662,N_1622);
xor U2316 (N_2316,N_2204,N_1765);
and U2317 (N_2317,N_2021,N_1559);
and U2318 (N_2318,N_2196,N_2079);
xor U2319 (N_2319,N_1767,N_2012);
and U2320 (N_2320,N_1774,N_2145);
or U2321 (N_2321,N_2169,N_1873);
or U2322 (N_2322,N_1819,N_1533);
xnor U2323 (N_2323,N_1616,N_2141);
xor U2324 (N_2324,N_1661,N_1581);
and U2325 (N_2325,N_1684,N_1965);
xor U2326 (N_2326,N_2162,N_1696);
nand U2327 (N_2327,N_1815,N_1575);
and U2328 (N_2328,N_1754,N_2226);
or U2329 (N_2329,N_1658,N_1663);
nand U2330 (N_2330,N_2060,N_1694);
xnor U2331 (N_2331,N_1692,N_2035);
and U2332 (N_2332,N_1923,N_2122);
and U2333 (N_2333,N_1536,N_1541);
and U2334 (N_2334,N_1999,N_2054);
and U2335 (N_2335,N_1676,N_2042);
xor U2336 (N_2336,N_2087,N_1558);
nand U2337 (N_2337,N_1764,N_1576);
nand U2338 (N_2338,N_1513,N_1693);
xnor U2339 (N_2339,N_1988,N_1981);
and U2340 (N_2340,N_2225,N_1863);
or U2341 (N_2341,N_1728,N_1982);
or U2342 (N_2342,N_2047,N_1934);
and U2343 (N_2343,N_1657,N_1935);
and U2344 (N_2344,N_2154,N_1920);
nor U2345 (N_2345,N_1562,N_1875);
or U2346 (N_2346,N_1734,N_1915);
nor U2347 (N_2347,N_1500,N_1931);
xnor U2348 (N_2348,N_1674,N_1651);
xnor U2349 (N_2349,N_1861,N_2230);
nor U2350 (N_2350,N_1652,N_1921);
nor U2351 (N_2351,N_2234,N_1720);
nand U2352 (N_2352,N_2068,N_2002);
nand U2353 (N_2353,N_1614,N_2213);
nand U2354 (N_2354,N_2177,N_1512);
and U2355 (N_2355,N_2051,N_1970);
nand U2356 (N_2356,N_1838,N_2197);
nand U2357 (N_2357,N_2201,N_1667);
and U2358 (N_2358,N_1740,N_1532);
nor U2359 (N_2359,N_2073,N_1572);
nor U2360 (N_2360,N_1625,N_1598);
xnor U2361 (N_2361,N_1874,N_2065);
nand U2362 (N_2362,N_2030,N_1749);
nand U2363 (N_2363,N_1876,N_1971);
xor U2364 (N_2364,N_2119,N_1912);
nand U2365 (N_2365,N_1933,N_1882);
nand U2366 (N_2366,N_1542,N_2231);
nand U2367 (N_2367,N_1546,N_2138);
and U2368 (N_2368,N_2167,N_1814);
xor U2369 (N_2369,N_1859,N_1552);
nand U2370 (N_2370,N_1701,N_1937);
or U2371 (N_2371,N_2149,N_1842);
xor U2372 (N_2372,N_1871,N_2001);
or U2373 (N_2373,N_2015,N_1753);
and U2374 (N_2374,N_1733,N_1884);
and U2375 (N_2375,N_2023,N_1630);
or U2376 (N_2376,N_2247,N_2074);
xor U2377 (N_2377,N_1836,N_2194);
xor U2378 (N_2378,N_1639,N_2233);
and U2379 (N_2379,N_1945,N_1706);
or U2380 (N_2380,N_1628,N_1823);
and U2381 (N_2381,N_2077,N_2063);
and U2382 (N_2382,N_2032,N_2150);
or U2383 (N_2383,N_2031,N_1953);
xnor U2384 (N_2384,N_2140,N_2100);
xnor U2385 (N_2385,N_1642,N_1804);
nand U2386 (N_2386,N_1669,N_1867);
xor U2387 (N_2387,N_1901,N_2185);
and U2388 (N_2388,N_2020,N_1670);
nor U2389 (N_2389,N_1688,N_1545);
nor U2390 (N_2390,N_1961,N_2157);
nand U2391 (N_2391,N_1845,N_1844);
nand U2392 (N_2392,N_1514,N_2224);
nor U2393 (N_2393,N_1621,N_2121);
or U2394 (N_2394,N_1947,N_1835);
and U2395 (N_2395,N_1664,N_1817);
or U2396 (N_2396,N_1610,N_1697);
nand U2397 (N_2397,N_1878,N_1713);
or U2398 (N_2398,N_2103,N_2179);
or U2399 (N_2399,N_1679,N_1724);
nand U2400 (N_2400,N_2058,N_2025);
nand U2401 (N_2401,N_2057,N_1703);
nor U2402 (N_2402,N_1641,N_1769);
nand U2403 (N_2403,N_1656,N_1645);
xor U2404 (N_2404,N_1710,N_1678);
or U2405 (N_2405,N_1735,N_2084);
nand U2406 (N_2406,N_1840,N_1881);
nand U2407 (N_2407,N_1918,N_1932);
nor U2408 (N_2408,N_2046,N_1699);
or U2409 (N_2409,N_1868,N_1551);
and U2410 (N_2410,N_1914,N_2055);
or U2411 (N_2411,N_1807,N_1537);
xnor U2412 (N_2412,N_1925,N_1707);
xnor U2413 (N_2413,N_1821,N_2212);
and U2414 (N_2414,N_1974,N_1509);
and U2415 (N_2415,N_1759,N_1946);
nand U2416 (N_2416,N_2215,N_2182);
nor U2417 (N_2417,N_1850,N_2134);
and U2418 (N_2418,N_2217,N_1776);
xor U2419 (N_2419,N_1890,N_1896);
or U2420 (N_2420,N_2242,N_1612);
xnor U2421 (N_2421,N_1567,N_1561);
xnor U2422 (N_2422,N_2156,N_1966);
nor U2423 (N_2423,N_2071,N_1675);
nor U2424 (N_2424,N_2236,N_1739);
xnor U2425 (N_2425,N_1573,N_2038);
xnor U2426 (N_2426,N_1565,N_2128);
or U2427 (N_2427,N_1886,N_2041);
xor U2428 (N_2428,N_2091,N_1623);
nand U2429 (N_2429,N_1705,N_1761);
nand U2430 (N_2430,N_2113,N_1564);
xnor U2431 (N_2431,N_2174,N_1847);
nand U2432 (N_2432,N_2034,N_1994);
and U2433 (N_2433,N_1906,N_2029);
and U2434 (N_2434,N_1987,N_2190);
nor U2435 (N_2435,N_1587,N_2019);
xnor U2436 (N_2436,N_2067,N_1887);
or U2437 (N_2437,N_1680,N_1802);
nor U2438 (N_2438,N_1540,N_1852);
nor U2439 (N_2439,N_1608,N_2235);
nor U2440 (N_2440,N_1595,N_2093);
nor U2441 (N_2441,N_1785,N_1780);
xor U2442 (N_2442,N_2152,N_2243);
or U2443 (N_2443,N_2092,N_2052);
nand U2444 (N_2444,N_1986,N_2178);
xor U2445 (N_2445,N_2061,N_1592);
or U2446 (N_2446,N_2075,N_2078);
or U2447 (N_2447,N_1810,N_1615);
nor U2448 (N_2448,N_2024,N_1827);
and U2449 (N_2449,N_2143,N_2183);
nand U2450 (N_2450,N_2089,N_1746);
nor U2451 (N_2451,N_1726,N_1985);
nor U2452 (N_2452,N_1527,N_2094);
and U2453 (N_2453,N_1959,N_1526);
nand U2454 (N_2454,N_1855,N_1858);
or U2455 (N_2455,N_2008,N_2112);
xor U2456 (N_2456,N_1911,N_2114);
or U2457 (N_2457,N_1738,N_2207);
nand U2458 (N_2458,N_2069,N_1752);
nor U2459 (N_2459,N_2107,N_1539);
or U2460 (N_2460,N_2221,N_1809);
nand U2461 (N_2461,N_2003,N_1963);
nor U2462 (N_2462,N_2083,N_1569);
xnor U2463 (N_2463,N_2123,N_2011);
or U2464 (N_2464,N_1960,N_2146);
nor U2465 (N_2465,N_2161,N_1857);
xnor U2466 (N_2466,N_1617,N_2232);
and U2467 (N_2467,N_1619,N_2192);
nand U2468 (N_2468,N_2133,N_2111);
or U2469 (N_2469,N_2189,N_1624);
xor U2470 (N_2470,N_1635,N_1609);
and U2471 (N_2471,N_1709,N_1799);
nor U2472 (N_2472,N_1812,N_1956);
nor U2473 (N_2473,N_2191,N_2159);
nor U2474 (N_2474,N_2049,N_1751);
and U2475 (N_2475,N_1520,N_1747);
nor U2476 (N_2476,N_1756,N_1877);
nor U2477 (N_2477,N_2195,N_2238);
xor U2478 (N_2478,N_1566,N_1632);
xnor U2479 (N_2479,N_1553,N_1556);
xor U2480 (N_2480,N_2142,N_1681);
and U2481 (N_2481,N_1797,N_1805);
xor U2482 (N_2482,N_2014,N_1683);
nor U2483 (N_2483,N_2096,N_1557);
nor U2484 (N_2484,N_1743,N_2095);
nor U2485 (N_2485,N_1927,N_1779);
or U2486 (N_2486,N_1943,N_1659);
and U2487 (N_2487,N_1570,N_2164);
and U2488 (N_2488,N_1941,N_1972);
or U2489 (N_2489,N_1647,N_1800);
xor U2490 (N_2490,N_1788,N_1507);
nor U2491 (N_2491,N_1597,N_1648);
or U2492 (N_2492,N_1588,N_1730);
and U2493 (N_2493,N_2005,N_1571);
nand U2494 (N_2494,N_1957,N_1690);
nand U2495 (N_2495,N_2016,N_1980);
nor U2496 (N_2496,N_1550,N_1631);
or U2497 (N_2497,N_2160,N_2181);
nand U2498 (N_2498,N_2099,N_2163);
and U2499 (N_2499,N_2036,N_1816);
and U2500 (N_2500,N_1968,N_1806);
and U2501 (N_2501,N_2043,N_2216);
xnor U2502 (N_2502,N_1771,N_1702);
xnor U2503 (N_2503,N_2176,N_1525);
nand U2504 (N_2504,N_2037,N_2105);
nand U2505 (N_2505,N_1582,N_1794);
xnor U2506 (N_2506,N_1518,N_1841);
nand U2507 (N_2507,N_2129,N_1506);
and U2508 (N_2508,N_1792,N_2211);
xor U2509 (N_2509,N_1786,N_1677);
xnor U2510 (N_2510,N_2109,N_1666);
or U2511 (N_2511,N_1904,N_2116);
nand U2512 (N_2512,N_1654,N_1627);
nor U2513 (N_2513,N_1711,N_1936);
xor U2514 (N_2514,N_1725,N_1894);
xor U2515 (N_2515,N_1538,N_2006);
nor U2516 (N_2516,N_1535,N_1846);
xor U2517 (N_2517,N_1851,N_1791);
nand U2518 (N_2518,N_2120,N_1993);
or U2519 (N_2519,N_1618,N_1721);
nand U2520 (N_2520,N_2097,N_1919);
and U2521 (N_2521,N_1849,N_1501);
and U2522 (N_2522,N_1548,N_1891);
xor U2523 (N_2523,N_1917,N_1924);
xor U2524 (N_2524,N_2039,N_1908);
nand U2525 (N_2525,N_1758,N_1606);
xnor U2526 (N_2526,N_2062,N_1995);
nand U2527 (N_2527,N_1913,N_2188);
and U2528 (N_2528,N_1589,N_2206);
nor U2529 (N_2529,N_1653,N_2048);
xor U2530 (N_2530,N_2000,N_2066);
or U2531 (N_2531,N_1549,N_1715);
xor U2532 (N_2532,N_1818,N_1748);
nand U2533 (N_2533,N_1649,N_2193);
or U2534 (N_2534,N_1502,N_1870);
nand U2535 (N_2535,N_1704,N_2086);
or U2536 (N_2536,N_1784,N_1605);
or U2537 (N_2537,N_1601,N_1744);
and U2538 (N_2538,N_1865,N_1973);
nor U2539 (N_2539,N_1928,N_2229);
nor U2540 (N_2540,N_1954,N_1510);
xor U2541 (N_2541,N_1902,N_2117);
xnor U2542 (N_2542,N_2102,N_1634);
nand U2543 (N_2543,N_2240,N_1793);
nand U2544 (N_2544,N_1732,N_1638);
nor U2545 (N_2545,N_1895,N_1958);
nand U2546 (N_2546,N_1837,N_1907);
and U2547 (N_2547,N_1729,N_1736);
xnor U2548 (N_2548,N_1996,N_2246);
and U2549 (N_2549,N_1517,N_2173);
nor U2550 (N_2550,N_1591,N_1997);
xor U2551 (N_2551,N_1584,N_2239);
xor U2552 (N_2552,N_1808,N_1629);
nand U2553 (N_2553,N_1885,N_1967);
and U2554 (N_2554,N_2072,N_2199);
nor U2555 (N_2555,N_1828,N_2130);
xor U2556 (N_2556,N_1757,N_1637);
xor U2557 (N_2557,N_1975,N_1671);
nand U2558 (N_2558,N_2127,N_2137);
nor U2559 (N_2559,N_2040,N_2209);
nand U2560 (N_2560,N_1560,N_2165);
or U2561 (N_2561,N_1686,N_1626);
and U2562 (N_2562,N_1990,N_2249);
nor U2563 (N_2563,N_1984,N_1521);
nand U2564 (N_2564,N_1529,N_1938);
nor U2565 (N_2565,N_1929,N_1949);
xnor U2566 (N_2566,N_1883,N_1897);
nand U2567 (N_2567,N_1796,N_2155);
nor U2568 (N_2568,N_2180,N_1723);
or U2569 (N_2569,N_1745,N_2045);
or U2570 (N_2570,N_1604,N_1528);
and U2571 (N_2571,N_1860,N_2050);
nand U2572 (N_2572,N_1976,N_2010);
nor U2573 (N_2573,N_2022,N_2172);
nor U2574 (N_2574,N_1824,N_1544);
nand U2575 (N_2575,N_1600,N_2132);
or U2576 (N_2576,N_2220,N_1534);
nor U2577 (N_2577,N_1620,N_1926);
nand U2578 (N_2578,N_2202,N_1755);
nor U2579 (N_2579,N_2175,N_1798);
nor U2580 (N_2580,N_1922,N_1801);
nor U2581 (N_2581,N_2082,N_1899);
and U2582 (N_2582,N_2148,N_1717);
xnor U2583 (N_2583,N_1820,N_2126);
or U2584 (N_2584,N_1803,N_1504);
and U2585 (N_2585,N_2125,N_1660);
and U2586 (N_2586,N_1531,N_1519);
and U2587 (N_2587,N_1830,N_2136);
nor U2588 (N_2588,N_1869,N_1714);
and U2589 (N_2589,N_2033,N_1594);
xor U2590 (N_2590,N_1719,N_1825);
nor U2591 (N_2591,N_1888,N_1613);
and U2592 (N_2592,N_1750,N_1593);
nor U2593 (N_2593,N_1977,N_1505);
xor U2594 (N_2594,N_1979,N_2009);
and U2595 (N_2595,N_2124,N_2070);
or U2596 (N_2596,N_1773,N_1829);
xor U2597 (N_2597,N_2090,N_1991);
xor U2598 (N_2598,N_1524,N_1596);
nor U2599 (N_2599,N_1768,N_2245);
or U2600 (N_2600,N_1930,N_2004);
xor U2601 (N_2601,N_1910,N_1962);
xnor U2602 (N_2602,N_1585,N_2110);
xor U2603 (N_2603,N_2184,N_2056);
or U2604 (N_2604,N_2205,N_2106);
nand U2605 (N_2605,N_1939,N_1577);
or U2606 (N_2606,N_2187,N_2166);
xor U2607 (N_2607,N_1940,N_1952);
or U2608 (N_2608,N_1826,N_1898);
and U2609 (N_2609,N_2158,N_2118);
or U2610 (N_2610,N_1839,N_1856);
and U2611 (N_2611,N_1741,N_1716);
or U2612 (N_2612,N_1942,N_1602);
and U2613 (N_2613,N_1909,N_1989);
nand U2614 (N_2614,N_1889,N_1766);
nand U2615 (N_2615,N_1969,N_1900);
nand U2616 (N_2616,N_1822,N_1611);
or U2617 (N_2617,N_1879,N_2171);
nand U2618 (N_2618,N_2017,N_1555);
xnor U2619 (N_2619,N_2108,N_1718);
nor U2620 (N_2620,N_1772,N_1916);
nor U2621 (N_2621,N_1978,N_1998);
nor U2622 (N_2622,N_1511,N_2222);
and U2623 (N_2623,N_1893,N_1687);
nor U2624 (N_2624,N_2227,N_2139);
and U2625 (N_2625,N_2109,N_1786);
nand U2626 (N_2626,N_1510,N_1913);
nor U2627 (N_2627,N_2009,N_1928);
nand U2628 (N_2628,N_2052,N_2114);
nor U2629 (N_2629,N_1553,N_2227);
nand U2630 (N_2630,N_1968,N_1840);
and U2631 (N_2631,N_1513,N_1559);
nor U2632 (N_2632,N_1661,N_1569);
and U2633 (N_2633,N_1857,N_1711);
nor U2634 (N_2634,N_1625,N_1934);
nand U2635 (N_2635,N_1904,N_2126);
xnor U2636 (N_2636,N_1680,N_2139);
xnor U2637 (N_2637,N_2096,N_2109);
and U2638 (N_2638,N_1616,N_1923);
nor U2639 (N_2639,N_1607,N_1980);
nor U2640 (N_2640,N_1652,N_2241);
xnor U2641 (N_2641,N_1795,N_1705);
nand U2642 (N_2642,N_2142,N_2051);
or U2643 (N_2643,N_2231,N_2164);
nand U2644 (N_2644,N_1810,N_2145);
and U2645 (N_2645,N_1524,N_2099);
and U2646 (N_2646,N_1548,N_1689);
and U2647 (N_2647,N_1660,N_1893);
or U2648 (N_2648,N_1525,N_1959);
and U2649 (N_2649,N_2077,N_2182);
or U2650 (N_2650,N_1577,N_2192);
and U2651 (N_2651,N_2187,N_2066);
xor U2652 (N_2652,N_2010,N_2029);
nand U2653 (N_2653,N_1660,N_2182);
and U2654 (N_2654,N_1928,N_2220);
nor U2655 (N_2655,N_2165,N_1860);
nor U2656 (N_2656,N_2178,N_1677);
and U2657 (N_2657,N_1865,N_1600);
nand U2658 (N_2658,N_2196,N_2167);
and U2659 (N_2659,N_2098,N_1719);
and U2660 (N_2660,N_1760,N_2190);
xor U2661 (N_2661,N_2072,N_2037);
xnor U2662 (N_2662,N_2239,N_1514);
and U2663 (N_2663,N_2090,N_2218);
xor U2664 (N_2664,N_2117,N_1852);
xor U2665 (N_2665,N_1733,N_2163);
xor U2666 (N_2666,N_1842,N_1725);
and U2667 (N_2667,N_1517,N_2163);
xor U2668 (N_2668,N_2129,N_1791);
or U2669 (N_2669,N_1950,N_1580);
xnor U2670 (N_2670,N_1556,N_2084);
or U2671 (N_2671,N_2222,N_2230);
or U2672 (N_2672,N_1798,N_2081);
or U2673 (N_2673,N_1842,N_2120);
nand U2674 (N_2674,N_1864,N_1778);
nor U2675 (N_2675,N_1661,N_1975);
xnor U2676 (N_2676,N_1786,N_1938);
xnor U2677 (N_2677,N_2045,N_1963);
nor U2678 (N_2678,N_1585,N_1747);
xnor U2679 (N_2679,N_1659,N_2069);
nor U2680 (N_2680,N_2019,N_1829);
nand U2681 (N_2681,N_2018,N_2121);
xnor U2682 (N_2682,N_2060,N_2073);
nand U2683 (N_2683,N_1943,N_2080);
nor U2684 (N_2684,N_1808,N_1920);
and U2685 (N_2685,N_1996,N_1834);
and U2686 (N_2686,N_1613,N_1760);
and U2687 (N_2687,N_1601,N_2010);
nor U2688 (N_2688,N_2184,N_1879);
nand U2689 (N_2689,N_1552,N_1554);
or U2690 (N_2690,N_2175,N_1737);
nor U2691 (N_2691,N_1970,N_1694);
or U2692 (N_2692,N_1651,N_1859);
and U2693 (N_2693,N_2140,N_1996);
or U2694 (N_2694,N_1556,N_1937);
and U2695 (N_2695,N_1536,N_1769);
xor U2696 (N_2696,N_1894,N_1604);
xor U2697 (N_2697,N_1695,N_1703);
nor U2698 (N_2698,N_2086,N_2010);
xor U2699 (N_2699,N_1770,N_2161);
xor U2700 (N_2700,N_2050,N_2119);
or U2701 (N_2701,N_1775,N_2059);
or U2702 (N_2702,N_2062,N_1915);
nor U2703 (N_2703,N_1827,N_1622);
or U2704 (N_2704,N_1722,N_1845);
and U2705 (N_2705,N_1931,N_1941);
or U2706 (N_2706,N_1711,N_1741);
xnor U2707 (N_2707,N_2037,N_1993);
xnor U2708 (N_2708,N_1936,N_1737);
and U2709 (N_2709,N_1818,N_2171);
xor U2710 (N_2710,N_1527,N_1636);
nor U2711 (N_2711,N_2207,N_1606);
or U2712 (N_2712,N_1660,N_1906);
or U2713 (N_2713,N_1610,N_1646);
nor U2714 (N_2714,N_1621,N_1649);
nand U2715 (N_2715,N_1558,N_1992);
xor U2716 (N_2716,N_1715,N_2210);
xnor U2717 (N_2717,N_2101,N_2182);
and U2718 (N_2718,N_2144,N_1978);
xnor U2719 (N_2719,N_2119,N_1528);
nor U2720 (N_2720,N_1664,N_1701);
and U2721 (N_2721,N_1606,N_1510);
nor U2722 (N_2722,N_2071,N_2193);
or U2723 (N_2723,N_1686,N_1553);
nand U2724 (N_2724,N_2222,N_1558);
and U2725 (N_2725,N_2141,N_1952);
or U2726 (N_2726,N_1874,N_2199);
or U2727 (N_2727,N_1603,N_1573);
nor U2728 (N_2728,N_2144,N_1518);
xnor U2729 (N_2729,N_1591,N_2115);
nand U2730 (N_2730,N_1716,N_1979);
or U2731 (N_2731,N_2226,N_1731);
nor U2732 (N_2732,N_1609,N_1766);
or U2733 (N_2733,N_1873,N_2234);
and U2734 (N_2734,N_1811,N_2146);
nand U2735 (N_2735,N_1550,N_1828);
xnor U2736 (N_2736,N_2015,N_2054);
nor U2737 (N_2737,N_1811,N_2170);
nand U2738 (N_2738,N_1881,N_2163);
nand U2739 (N_2739,N_1858,N_1638);
xor U2740 (N_2740,N_1665,N_2012);
and U2741 (N_2741,N_2090,N_1619);
or U2742 (N_2742,N_1523,N_1723);
xor U2743 (N_2743,N_1946,N_2245);
and U2744 (N_2744,N_1906,N_2156);
xor U2745 (N_2745,N_2245,N_1939);
or U2746 (N_2746,N_1567,N_1903);
or U2747 (N_2747,N_1567,N_1944);
nor U2748 (N_2748,N_2187,N_2113);
nand U2749 (N_2749,N_1510,N_1941);
xor U2750 (N_2750,N_1804,N_2199);
nor U2751 (N_2751,N_2127,N_1937);
nor U2752 (N_2752,N_1778,N_1795);
nor U2753 (N_2753,N_2230,N_1604);
nand U2754 (N_2754,N_1867,N_1861);
nor U2755 (N_2755,N_2015,N_1999);
xor U2756 (N_2756,N_1830,N_1639);
nor U2757 (N_2757,N_1786,N_1980);
or U2758 (N_2758,N_2026,N_1515);
or U2759 (N_2759,N_1820,N_1975);
and U2760 (N_2760,N_1521,N_2071);
xnor U2761 (N_2761,N_2083,N_2169);
nand U2762 (N_2762,N_1899,N_1693);
nor U2763 (N_2763,N_2212,N_1948);
nor U2764 (N_2764,N_1611,N_2200);
xnor U2765 (N_2765,N_2041,N_2132);
and U2766 (N_2766,N_1795,N_2135);
nor U2767 (N_2767,N_1543,N_1575);
nand U2768 (N_2768,N_1940,N_2095);
and U2769 (N_2769,N_2216,N_1995);
nor U2770 (N_2770,N_1854,N_1974);
xor U2771 (N_2771,N_2082,N_2153);
and U2772 (N_2772,N_2179,N_1782);
and U2773 (N_2773,N_1856,N_2030);
and U2774 (N_2774,N_2220,N_2081);
xnor U2775 (N_2775,N_2093,N_2224);
and U2776 (N_2776,N_2208,N_2021);
nand U2777 (N_2777,N_1769,N_2090);
and U2778 (N_2778,N_1561,N_2061);
nand U2779 (N_2779,N_1559,N_1617);
xor U2780 (N_2780,N_1553,N_1831);
and U2781 (N_2781,N_1668,N_1832);
and U2782 (N_2782,N_2132,N_2233);
or U2783 (N_2783,N_1580,N_2138);
xor U2784 (N_2784,N_1768,N_2175);
nand U2785 (N_2785,N_1621,N_2212);
or U2786 (N_2786,N_1817,N_1804);
nor U2787 (N_2787,N_1784,N_1816);
xor U2788 (N_2788,N_1875,N_1937);
xor U2789 (N_2789,N_1728,N_1623);
xor U2790 (N_2790,N_1638,N_1665);
nor U2791 (N_2791,N_1719,N_1879);
and U2792 (N_2792,N_1814,N_1770);
nand U2793 (N_2793,N_2058,N_2087);
nand U2794 (N_2794,N_1549,N_2213);
and U2795 (N_2795,N_1835,N_1648);
or U2796 (N_2796,N_2101,N_2097);
or U2797 (N_2797,N_1816,N_1663);
nor U2798 (N_2798,N_1727,N_2048);
and U2799 (N_2799,N_2111,N_1516);
xnor U2800 (N_2800,N_1644,N_2112);
nand U2801 (N_2801,N_1739,N_1945);
or U2802 (N_2802,N_1556,N_1539);
or U2803 (N_2803,N_2065,N_1629);
and U2804 (N_2804,N_1716,N_2205);
and U2805 (N_2805,N_1566,N_2222);
xnor U2806 (N_2806,N_1971,N_2176);
xnor U2807 (N_2807,N_1831,N_1532);
nand U2808 (N_2808,N_1906,N_2249);
nor U2809 (N_2809,N_1726,N_2114);
xnor U2810 (N_2810,N_2122,N_2020);
nor U2811 (N_2811,N_1804,N_2212);
nor U2812 (N_2812,N_2203,N_1520);
and U2813 (N_2813,N_2157,N_2075);
nor U2814 (N_2814,N_1572,N_1968);
nor U2815 (N_2815,N_2185,N_1820);
or U2816 (N_2816,N_2151,N_2246);
nand U2817 (N_2817,N_2078,N_1697);
nand U2818 (N_2818,N_1539,N_2167);
or U2819 (N_2819,N_1580,N_2189);
or U2820 (N_2820,N_2145,N_1633);
nand U2821 (N_2821,N_1625,N_1777);
xnor U2822 (N_2822,N_2062,N_2164);
xnor U2823 (N_2823,N_1525,N_2002);
xnor U2824 (N_2824,N_1909,N_1904);
or U2825 (N_2825,N_1805,N_1812);
nand U2826 (N_2826,N_2177,N_2067);
or U2827 (N_2827,N_1565,N_2162);
xor U2828 (N_2828,N_1717,N_2236);
and U2829 (N_2829,N_1857,N_1587);
xor U2830 (N_2830,N_1851,N_1682);
nor U2831 (N_2831,N_1964,N_1578);
xor U2832 (N_2832,N_2149,N_1822);
and U2833 (N_2833,N_1729,N_1516);
nor U2834 (N_2834,N_1593,N_1733);
nand U2835 (N_2835,N_2193,N_1586);
xnor U2836 (N_2836,N_2128,N_1553);
or U2837 (N_2837,N_1883,N_1508);
nand U2838 (N_2838,N_1693,N_1830);
nor U2839 (N_2839,N_2151,N_1860);
or U2840 (N_2840,N_2196,N_1555);
or U2841 (N_2841,N_1961,N_1944);
xnor U2842 (N_2842,N_1852,N_1792);
nor U2843 (N_2843,N_1923,N_1641);
nand U2844 (N_2844,N_1648,N_1637);
or U2845 (N_2845,N_1918,N_2243);
xor U2846 (N_2846,N_2163,N_1736);
xnor U2847 (N_2847,N_1760,N_1716);
nand U2848 (N_2848,N_1669,N_1739);
nand U2849 (N_2849,N_1798,N_1508);
or U2850 (N_2850,N_1505,N_1998);
xnor U2851 (N_2851,N_1825,N_1915);
nor U2852 (N_2852,N_1866,N_1911);
xor U2853 (N_2853,N_1932,N_1650);
nor U2854 (N_2854,N_1615,N_2029);
nand U2855 (N_2855,N_2231,N_1677);
nor U2856 (N_2856,N_1804,N_1840);
xor U2857 (N_2857,N_1669,N_1637);
nand U2858 (N_2858,N_1941,N_2071);
xor U2859 (N_2859,N_2048,N_1882);
or U2860 (N_2860,N_2114,N_2107);
xor U2861 (N_2861,N_2196,N_1553);
or U2862 (N_2862,N_2239,N_1854);
or U2863 (N_2863,N_2182,N_1796);
and U2864 (N_2864,N_1962,N_2037);
nor U2865 (N_2865,N_1994,N_2087);
xor U2866 (N_2866,N_2058,N_1792);
and U2867 (N_2867,N_1806,N_1999);
xnor U2868 (N_2868,N_1571,N_1995);
and U2869 (N_2869,N_1863,N_2028);
nand U2870 (N_2870,N_2082,N_2197);
or U2871 (N_2871,N_2220,N_1527);
or U2872 (N_2872,N_1507,N_1845);
nor U2873 (N_2873,N_1542,N_1556);
nor U2874 (N_2874,N_1802,N_1857);
or U2875 (N_2875,N_1739,N_1909);
or U2876 (N_2876,N_1925,N_2078);
xnor U2877 (N_2877,N_1887,N_1844);
and U2878 (N_2878,N_1688,N_2201);
or U2879 (N_2879,N_2165,N_1975);
or U2880 (N_2880,N_1780,N_1620);
or U2881 (N_2881,N_2077,N_1770);
and U2882 (N_2882,N_2232,N_2101);
nand U2883 (N_2883,N_2069,N_2136);
and U2884 (N_2884,N_1684,N_2246);
nand U2885 (N_2885,N_1960,N_1956);
nand U2886 (N_2886,N_2066,N_2154);
nor U2887 (N_2887,N_2152,N_1929);
and U2888 (N_2888,N_1624,N_2066);
nor U2889 (N_2889,N_1587,N_2003);
xnor U2890 (N_2890,N_1947,N_2134);
nand U2891 (N_2891,N_1956,N_1577);
xnor U2892 (N_2892,N_1915,N_2110);
xnor U2893 (N_2893,N_1937,N_2034);
nand U2894 (N_2894,N_2089,N_1692);
nor U2895 (N_2895,N_1831,N_2042);
xor U2896 (N_2896,N_1854,N_1614);
xnor U2897 (N_2897,N_2051,N_2222);
nand U2898 (N_2898,N_1796,N_1529);
or U2899 (N_2899,N_1844,N_2145);
or U2900 (N_2900,N_1841,N_1543);
nand U2901 (N_2901,N_2036,N_1888);
nand U2902 (N_2902,N_1519,N_1870);
nand U2903 (N_2903,N_1734,N_2051);
xor U2904 (N_2904,N_1506,N_2125);
and U2905 (N_2905,N_2122,N_2236);
nor U2906 (N_2906,N_1704,N_1572);
xnor U2907 (N_2907,N_2241,N_1752);
and U2908 (N_2908,N_1582,N_2018);
or U2909 (N_2909,N_2025,N_1539);
nand U2910 (N_2910,N_1714,N_1599);
nor U2911 (N_2911,N_1829,N_2180);
nor U2912 (N_2912,N_1886,N_1569);
and U2913 (N_2913,N_1705,N_1988);
and U2914 (N_2914,N_2024,N_2093);
nand U2915 (N_2915,N_2201,N_1947);
or U2916 (N_2916,N_2196,N_1950);
nor U2917 (N_2917,N_1940,N_2152);
nand U2918 (N_2918,N_1544,N_1521);
nor U2919 (N_2919,N_1996,N_2149);
and U2920 (N_2920,N_2106,N_1825);
and U2921 (N_2921,N_1945,N_1851);
nand U2922 (N_2922,N_1768,N_2237);
nand U2923 (N_2923,N_1971,N_1976);
xnor U2924 (N_2924,N_1742,N_1804);
and U2925 (N_2925,N_2138,N_1538);
xor U2926 (N_2926,N_2064,N_1727);
nor U2927 (N_2927,N_2113,N_1538);
nand U2928 (N_2928,N_2175,N_1752);
and U2929 (N_2929,N_1954,N_1645);
or U2930 (N_2930,N_2115,N_2166);
xor U2931 (N_2931,N_1840,N_1627);
or U2932 (N_2932,N_2226,N_1628);
or U2933 (N_2933,N_2057,N_2197);
xnor U2934 (N_2934,N_1970,N_1967);
nor U2935 (N_2935,N_1667,N_1727);
or U2936 (N_2936,N_2169,N_2140);
nor U2937 (N_2937,N_1534,N_2024);
and U2938 (N_2938,N_1512,N_1531);
xor U2939 (N_2939,N_1511,N_1629);
nor U2940 (N_2940,N_2133,N_2208);
or U2941 (N_2941,N_1892,N_1548);
xnor U2942 (N_2942,N_1879,N_1794);
and U2943 (N_2943,N_1853,N_2026);
nand U2944 (N_2944,N_1780,N_2000);
nor U2945 (N_2945,N_1647,N_1870);
xnor U2946 (N_2946,N_1625,N_2215);
or U2947 (N_2947,N_1715,N_1710);
nand U2948 (N_2948,N_1950,N_2013);
nand U2949 (N_2949,N_1554,N_2196);
or U2950 (N_2950,N_2080,N_1526);
xor U2951 (N_2951,N_1661,N_2159);
nor U2952 (N_2952,N_2068,N_2018);
nor U2953 (N_2953,N_1669,N_1890);
or U2954 (N_2954,N_2089,N_2209);
xor U2955 (N_2955,N_2096,N_2066);
nand U2956 (N_2956,N_2236,N_2204);
nand U2957 (N_2957,N_2010,N_1633);
or U2958 (N_2958,N_1919,N_1543);
nor U2959 (N_2959,N_2164,N_1501);
nand U2960 (N_2960,N_2013,N_1861);
nand U2961 (N_2961,N_1628,N_1691);
nand U2962 (N_2962,N_2162,N_1694);
or U2963 (N_2963,N_1757,N_1641);
nand U2964 (N_2964,N_2116,N_2083);
or U2965 (N_2965,N_1591,N_1872);
or U2966 (N_2966,N_1585,N_1993);
or U2967 (N_2967,N_2099,N_2230);
xnor U2968 (N_2968,N_1754,N_1631);
nor U2969 (N_2969,N_2121,N_2083);
xor U2970 (N_2970,N_2083,N_2096);
and U2971 (N_2971,N_1549,N_2223);
xor U2972 (N_2972,N_2149,N_1853);
nor U2973 (N_2973,N_1577,N_2193);
nor U2974 (N_2974,N_1890,N_1534);
or U2975 (N_2975,N_1616,N_1738);
and U2976 (N_2976,N_1882,N_2198);
xor U2977 (N_2977,N_1515,N_2089);
nor U2978 (N_2978,N_2237,N_1504);
and U2979 (N_2979,N_1536,N_2134);
nor U2980 (N_2980,N_2151,N_1665);
and U2981 (N_2981,N_1535,N_1590);
or U2982 (N_2982,N_1791,N_2236);
nand U2983 (N_2983,N_2072,N_2158);
and U2984 (N_2984,N_1569,N_1575);
nor U2985 (N_2985,N_1681,N_1721);
and U2986 (N_2986,N_1620,N_1719);
nand U2987 (N_2987,N_2184,N_1753);
xnor U2988 (N_2988,N_2191,N_2149);
and U2989 (N_2989,N_1951,N_2232);
and U2990 (N_2990,N_1735,N_1572);
nor U2991 (N_2991,N_1580,N_1775);
nand U2992 (N_2992,N_1546,N_2071);
or U2993 (N_2993,N_1960,N_1714);
and U2994 (N_2994,N_1954,N_1518);
nor U2995 (N_2995,N_1583,N_1689);
nand U2996 (N_2996,N_1749,N_1673);
xor U2997 (N_2997,N_1568,N_1647);
and U2998 (N_2998,N_2033,N_1899);
or U2999 (N_2999,N_1940,N_1814);
nor UO_0 (O_0,N_2854,N_2407);
and UO_1 (O_1,N_2431,N_2288);
nand UO_2 (O_2,N_2957,N_2852);
nor UO_3 (O_3,N_2322,N_2881);
xor UO_4 (O_4,N_2297,N_2324);
xnor UO_5 (O_5,N_2755,N_2848);
xnor UO_6 (O_6,N_2263,N_2303);
xnor UO_7 (O_7,N_2445,N_2552);
xor UO_8 (O_8,N_2292,N_2284);
xnor UO_9 (O_9,N_2337,N_2627);
xor UO_10 (O_10,N_2912,N_2658);
nand UO_11 (O_11,N_2513,N_2287);
or UO_12 (O_12,N_2868,N_2795);
xor UO_13 (O_13,N_2908,N_2611);
xnor UO_14 (O_14,N_2849,N_2365);
nor UO_15 (O_15,N_2969,N_2580);
xnor UO_16 (O_16,N_2869,N_2539);
and UO_17 (O_17,N_2613,N_2759);
or UO_18 (O_18,N_2491,N_2743);
xor UO_19 (O_19,N_2979,N_2838);
or UO_20 (O_20,N_2452,N_2326);
or UO_21 (O_21,N_2254,N_2440);
or UO_22 (O_22,N_2680,N_2345);
nand UO_23 (O_23,N_2449,N_2919);
and UO_24 (O_24,N_2739,N_2765);
nand UO_25 (O_25,N_2764,N_2258);
or UO_26 (O_26,N_2545,N_2994);
xnor UO_27 (O_27,N_2520,N_2479);
nand UO_28 (O_28,N_2895,N_2836);
and UO_29 (O_29,N_2887,N_2295);
or UO_30 (O_30,N_2846,N_2753);
and UO_31 (O_31,N_2812,N_2703);
nand UO_32 (O_32,N_2830,N_2293);
xor UO_33 (O_33,N_2712,N_2896);
nor UO_34 (O_34,N_2581,N_2530);
xnor UO_35 (O_35,N_2467,N_2571);
and UO_36 (O_36,N_2387,N_2644);
and UO_37 (O_37,N_2570,N_2374);
nor UO_38 (O_38,N_2600,N_2772);
or UO_39 (O_39,N_2857,N_2873);
nand UO_40 (O_40,N_2515,N_2397);
or UO_41 (O_41,N_2259,N_2261);
xor UO_42 (O_42,N_2933,N_2867);
or UO_43 (O_43,N_2891,N_2777);
and UO_44 (O_44,N_2949,N_2503);
xnor UO_45 (O_45,N_2874,N_2648);
nand UO_46 (O_46,N_2475,N_2304);
and UO_47 (O_47,N_2332,N_2606);
nand UO_48 (O_48,N_2321,N_2549);
nand UO_49 (O_49,N_2670,N_2690);
xnor UO_50 (O_50,N_2628,N_2853);
nor UO_51 (O_51,N_2529,N_2694);
nand UO_52 (O_52,N_2499,N_2952);
xnor UO_53 (O_53,N_2740,N_2507);
or UO_54 (O_54,N_2927,N_2910);
nor UO_55 (O_55,N_2706,N_2920);
and UO_56 (O_56,N_2342,N_2855);
nor UO_57 (O_57,N_2481,N_2464);
or UO_58 (O_58,N_2566,N_2421);
and UO_59 (O_59,N_2885,N_2892);
nand UO_60 (O_60,N_2900,N_2972);
xor UO_61 (O_61,N_2934,N_2935);
or UO_62 (O_62,N_2422,N_2450);
or UO_63 (O_63,N_2792,N_2403);
nor UO_64 (O_64,N_2405,N_2542);
and UO_65 (O_65,N_2540,N_2872);
nand UO_66 (O_66,N_2357,N_2681);
nor UO_67 (O_67,N_2575,N_2831);
nor UO_68 (O_68,N_2859,N_2889);
nor UO_69 (O_69,N_2594,N_2569);
nor UO_70 (O_70,N_2909,N_2842);
nor UO_71 (O_71,N_2386,N_2769);
or UO_72 (O_72,N_2604,N_2428);
or UO_73 (O_73,N_2301,N_2265);
xor UO_74 (O_74,N_2799,N_2330);
nor UO_75 (O_75,N_2578,N_2696);
or UO_76 (O_76,N_2748,N_2442);
nor UO_77 (O_77,N_2937,N_2646);
nor UO_78 (O_78,N_2635,N_2730);
nor UO_79 (O_79,N_2702,N_2745);
xnor UO_80 (O_80,N_2388,N_2583);
nor UO_81 (O_81,N_2724,N_2923);
nand UO_82 (O_82,N_2984,N_2424);
xor UO_83 (O_83,N_2557,N_2733);
nor UO_84 (O_84,N_2416,N_2823);
and UO_85 (O_85,N_2822,N_2797);
or UO_86 (O_86,N_2310,N_2472);
xor UO_87 (O_87,N_2942,N_2713);
and UO_88 (O_88,N_2672,N_2573);
and UO_89 (O_89,N_2269,N_2533);
or UO_90 (O_90,N_2944,N_2932);
or UO_91 (O_91,N_2951,N_2804);
and UO_92 (O_92,N_2928,N_2538);
or UO_93 (O_93,N_2541,N_2897);
nor UO_94 (O_94,N_2615,N_2390);
nor UO_95 (O_95,N_2877,N_2563);
nand UO_96 (O_96,N_2856,N_2929);
and UO_97 (O_97,N_2470,N_2858);
xor UO_98 (O_98,N_2903,N_2788);
nand UO_99 (O_99,N_2722,N_2662);
xnor UO_100 (O_100,N_2808,N_2385);
xnor UO_101 (O_101,N_2921,N_2446);
or UO_102 (O_102,N_2953,N_2947);
xnor UO_103 (O_103,N_2294,N_2590);
and UO_104 (O_104,N_2360,N_2786);
xnor UO_105 (O_105,N_2531,N_2266);
and UO_106 (O_106,N_2970,N_2805);
nand UO_107 (O_107,N_2302,N_2410);
and UO_108 (O_108,N_2819,N_2567);
nor UO_109 (O_109,N_2977,N_2863);
xor UO_110 (O_110,N_2262,N_2882);
and UO_111 (O_111,N_2279,N_2883);
and UO_112 (O_112,N_2653,N_2377);
xnor UO_113 (O_113,N_2641,N_2906);
nor UO_114 (O_114,N_2603,N_2950);
and UO_115 (O_115,N_2311,N_2492);
xnor UO_116 (O_116,N_2483,N_2943);
or UO_117 (O_117,N_2916,N_2589);
or UO_118 (O_118,N_2577,N_2700);
and UO_119 (O_119,N_2298,N_2666);
nand UO_120 (O_120,N_2392,N_2664);
and UO_121 (O_121,N_2760,N_2427);
xor UO_122 (O_122,N_2956,N_2462);
xnor UO_123 (O_123,N_2723,N_2276);
and UO_124 (O_124,N_2809,N_2794);
or UO_125 (O_125,N_2353,N_2349);
xnor UO_126 (O_126,N_2985,N_2558);
nor UO_127 (O_127,N_2582,N_2551);
nand UO_128 (O_128,N_2899,N_2290);
or UO_129 (O_129,N_2766,N_2546);
xnor UO_130 (O_130,N_2514,N_2574);
and UO_131 (O_131,N_2963,N_2731);
nor UO_132 (O_132,N_2843,N_2964);
xnor UO_133 (O_133,N_2693,N_2645);
nand UO_134 (O_134,N_2775,N_2750);
nor UO_135 (O_135,N_2742,N_2612);
nor UO_136 (O_136,N_2343,N_2496);
xnor UO_137 (O_137,N_2468,N_2461);
nand UO_138 (O_138,N_2938,N_2255);
xor UO_139 (O_139,N_2598,N_2665);
nor UO_140 (O_140,N_2966,N_2423);
or UO_141 (O_141,N_2380,N_2835);
xor UO_142 (O_142,N_2283,N_2682);
nand UO_143 (O_143,N_2289,N_2880);
and UO_144 (O_144,N_2413,N_2820);
nor UO_145 (O_145,N_2597,N_2331);
nand UO_146 (O_146,N_2443,N_2691);
nand UO_147 (O_147,N_2465,N_2476);
nor UO_148 (O_148,N_2918,N_2780);
and UO_149 (O_149,N_2497,N_2992);
xor UO_150 (O_150,N_2528,N_2318);
nand UO_151 (O_151,N_2996,N_2975);
or UO_152 (O_152,N_2523,N_2274);
and UO_153 (O_153,N_2751,N_2411);
and UO_154 (O_154,N_2605,N_2381);
xor UO_155 (O_155,N_2654,N_2791);
xor UO_156 (O_156,N_2404,N_2257);
xor UO_157 (O_157,N_2814,N_2320);
nor UO_158 (O_158,N_2516,N_2323);
nor UO_159 (O_159,N_2584,N_2555);
or UO_160 (O_160,N_2596,N_2562);
nand UO_161 (O_161,N_2264,N_2968);
nand UO_162 (O_162,N_2587,N_2911);
nand UO_163 (O_163,N_2828,N_2990);
or UO_164 (O_164,N_2463,N_2399);
nor UO_165 (O_165,N_2409,N_2798);
nand UO_166 (O_166,N_2510,N_2998);
or UO_167 (O_167,N_2622,N_2632);
or UO_168 (O_168,N_2778,N_2761);
or UO_169 (O_169,N_2369,N_2710);
nor UO_170 (O_170,N_2457,N_2640);
and UO_171 (O_171,N_2466,N_2459);
or UO_172 (O_172,N_2291,N_2732);
nand UO_173 (O_173,N_2401,N_2862);
and UO_174 (O_174,N_2608,N_2363);
xor UO_175 (O_175,N_2671,N_2384);
or UO_176 (O_176,N_2768,N_2618);
nor UO_177 (O_177,N_2741,N_2500);
xor UO_178 (O_178,N_2636,N_2537);
and UO_179 (O_179,N_2486,N_2746);
or UO_180 (O_180,N_2824,N_2678);
nor UO_181 (O_181,N_2432,N_2915);
and UO_182 (O_182,N_2735,N_2926);
nor UO_183 (O_183,N_2800,N_2829);
or UO_184 (O_184,N_2425,N_2660);
nor UO_185 (O_185,N_2999,N_2316);
xnor UO_186 (O_186,N_2752,N_2488);
or UO_187 (O_187,N_2941,N_2727);
or UO_188 (O_188,N_2275,N_2817);
or UO_189 (O_189,N_2988,N_2347);
nor UO_190 (O_190,N_2356,N_2861);
nor UO_191 (O_191,N_2663,N_2803);
or UO_192 (O_192,N_2339,N_2965);
or UO_193 (O_193,N_2429,N_2398);
xnor UO_194 (O_194,N_2754,N_2256);
nand UO_195 (O_195,N_2736,N_2451);
and UO_196 (O_196,N_2319,N_2879);
xor UO_197 (O_197,N_2726,N_2689);
or UO_198 (O_198,N_2890,N_2839);
and UO_199 (O_199,N_2783,N_2917);
or UO_200 (O_200,N_2441,N_2980);
and UO_201 (O_201,N_2286,N_2400);
or UO_202 (O_202,N_2453,N_2484);
or UO_203 (O_203,N_2375,N_2565);
nor UO_204 (O_204,N_2904,N_2834);
and UO_205 (O_205,N_2536,N_2674);
xnor UO_206 (O_206,N_2981,N_2866);
nor UO_207 (O_207,N_2554,N_2273);
nand UO_208 (O_208,N_2699,N_2436);
or UO_209 (O_209,N_2454,N_2773);
xnor UO_210 (O_210,N_2989,N_2329);
or UO_211 (O_211,N_2278,N_2480);
or UO_212 (O_212,N_2687,N_2361);
or UO_213 (O_213,N_2876,N_2406);
nor UO_214 (O_214,N_2717,N_2816);
xnor UO_215 (O_215,N_2414,N_2490);
and UO_216 (O_216,N_2901,N_2827);
or UO_217 (O_217,N_2352,N_2758);
and UO_218 (O_218,N_2512,N_2821);
nor UO_219 (O_219,N_2522,N_2493);
xnor UO_220 (O_220,N_2744,N_2971);
nor UO_221 (O_221,N_2708,N_2373);
nand UO_222 (O_222,N_2308,N_2253);
xor UO_223 (O_223,N_2378,N_2907);
nand UO_224 (O_224,N_2793,N_2556);
xnor UO_225 (O_225,N_2576,N_2844);
nand UO_226 (O_226,N_2864,N_2435);
nand UO_227 (O_227,N_2677,N_2517);
xor UO_228 (O_228,N_2946,N_2905);
or UO_229 (O_229,N_2315,N_2757);
and UO_230 (O_230,N_2502,N_2350);
and UO_231 (O_231,N_2945,N_2930);
and UO_232 (O_232,N_2782,N_2300);
nor UO_233 (O_233,N_2894,N_2679);
nand UO_234 (O_234,N_2607,N_2371);
xor UO_235 (O_235,N_2806,N_2630);
or UO_236 (O_236,N_2417,N_2433);
nor UO_237 (O_237,N_2995,N_2643);
nor UO_238 (O_238,N_2925,N_2747);
or UO_239 (O_239,N_2495,N_2367);
nand UO_240 (O_240,N_2477,N_2282);
xor UO_241 (O_241,N_2620,N_2796);
nor UO_242 (O_242,N_2610,N_2922);
or UO_243 (O_243,N_2973,N_2368);
nor UO_244 (O_244,N_2351,N_2647);
nand UO_245 (O_245,N_2826,N_2978);
nor UO_246 (O_246,N_2599,N_2684);
nor UO_247 (O_247,N_2588,N_2637);
xor UO_248 (O_248,N_2616,N_2355);
nor UO_249 (O_249,N_2277,N_2376);
or UO_250 (O_250,N_2591,N_2306);
or UO_251 (O_251,N_2914,N_2455);
or UO_252 (O_252,N_2312,N_2787);
xor UO_253 (O_253,N_2408,N_2667);
and UO_254 (O_254,N_2313,N_2870);
or UO_255 (O_255,N_2617,N_2333);
nand UO_256 (O_256,N_2701,N_2811);
and UO_257 (O_257,N_2372,N_2737);
nand UO_258 (O_258,N_2958,N_2832);
nor UO_259 (O_259,N_2714,N_2716);
nand UO_260 (O_260,N_2886,N_2358);
and UO_261 (O_261,N_2725,N_2650);
or UO_262 (O_262,N_2801,N_2639);
xor UO_263 (O_263,N_2448,N_2344);
and UO_264 (O_264,N_2550,N_2469);
or UO_265 (O_265,N_2655,N_2781);
xor UO_266 (O_266,N_2592,N_2354);
nand UO_267 (O_267,N_2718,N_2729);
and UO_268 (O_268,N_2784,N_2893);
and UO_269 (O_269,N_2370,N_2532);
nor UO_270 (O_270,N_2389,N_2456);
nand UO_271 (O_271,N_2847,N_2524);
and UO_272 (O_272,N_2692,N_2704);
xnor UO_273 (O_273,N_2705,N_2837);
and UO_274 (O_274,N_2790,N_2394);
or UO_275 (O_275,N_2268,N_2865);
nand UO_276 (O_276,N_2991,N_2335);
or UO_277 (O_277,N_2993,N_2767);
nand UO_278 (O_278,N_2651,N_2683);
xnor UO_279 (O_279,N_2395,N_2260);
or UO_280 (O_280,N_2625,N_2974);
nand UO_281 (O_281,N_2948,N_2738);
or UO_282 (O_282,N_2711,N_2676);
xnor UO_283 (O_283,N_2494,N_2875);
and UO_284 (O_284,N_2506,N_2478);
and UO_285 (O_285,N_2888,N_2884);
nand UO_286 (O_286,N_2504,N_2967);
nand UO_287 (O_287,N_2771,N_2314);
nand UO_288 (O_288,N_2547,N_2366);
xor UO_289 (O_289,N_2444,N_2698);
or UO_290 (O_290,N_2825,N_2633);
or UO_291 (O_291,N_2460,N_2818);
xor UO_292 (O_292,N_2346,N_2521);
xor UO_293 (O_293,N_2252,N_2983);
and UO_294 (O_294,N_2585,N_2661);
or UO_295 (O_295,N_2810,N_2695);
and UO_296 (O_296,N_2638,N_2334);
nor UO_297 (O_297,N_2997,N_2634);
xor UO_298 (O_298,N_2609,N_2774);
and UO_299 (O_299,N_2447,N_2626);
nand UO_300 (O_300,N_2489,N_2940);
nor UO_301 (O_301,N_2415,N_2841);
nand UO_302 (O_302,N_2393,N_2527);
xor UO_303 (O_303,N_2707,N_2721);
xnor UO_304 (O_304,N_2325,N_2382);
xnor UO_305 (O_305,N_2341,N_2813);
and UO_306 (O_306,N_2749,N_2487);
or UO_307 (O_307,N_2762,N_2601);
nand UO_308 (O_308,N_2986,N_2623);
or UO_309 (O_309,N_2756,N_2685);
xnor UO_310 (O_310,N_2624,N_2535);
or UO_311 (O_311,N_2675,N_2338);
xnor UO_312 (O_312,N_2564,N_2299);
xnor UO_313 (O_313,N_2579,N_2391);
or UO_314 (O_314,N_2340,N_2720);
nand UO_315 (O_315,N_2437,N_2418);
and UO_316 (O_316,N_2619,N_2402);
or UO_317 (O_317,N_2709,N_2482);
and UO_318 (O_318,N_2327,N_2763);
or UO_319 (O_319,N_2438,N_2544);
xnor UO_320 (O_320,N_2924,N_2396);
xnor UO_321 (O_321,N_2419,N_2548);
nand UO_322 (O_322,N_2614,N_2250);
nor UO_323 (O_323,N_2595,N_2328);
nand UO_324 (O_324,N_2802,N_2296);
nand UO_325 (O_325,N_2383,N_2776);
nand UO_326 (O_326,N_2458,N_2270);
xnor UO_327 (O_327,N_2697,N_2789);
or UO_328 (O_328,N_2734,N_2631);
xor UO_329 (O_329,N_2359,N_2267);
or UO_330 (O_330,N_2560,N_2526);
nand UO_331 (O_331,N_2348,N_2379);
nor UO_332 (O_332,N_2426,N_2474);
or UO_333 (O_333,N_2987,N_2961);
nand UO_334 (O_334,N_2307,N_2572);
xnor UO_335 (O_335,N_2534,N_2362);
nor UO_336 (O_336,N_2364,N_2939);
nor UO_337 (O_337,N_2982,N_2656);
nor UO_338 (O_338,N_2833,N_2669);
nand UO_339 (O_339,N_2686,N_2518);
nand UO_340 (O_340,N_2807,N_2509);
and UO_341 (O_341,N_2501,N_2629);
xnor UO_342 (O_342,N_2593,N_2336);
xor UO_343 (O_343,N_2430,N_2902);
or UO_344 (O_344,N_2959,N_2851);
nor UO_345 (O_345,N_2955,N_2719);
nor UO_346 (O_346,N_2715,N_2543);
xnor UO_347 (O_347,N_2898,N_2770);
and UO_348 (O_348,N_2850,N_2960);
nand UO_349 (O_349,N_2659,N_2471);
and UO_350 (O_350,N_2954,N_2485);
nand UO_351 (O_351,N_2439,N_2434);
or UO_352 (O_352,N_2586,N_2649);
or UO_353 (O_353,N_2642,N_2561);
nand UO_354 (O_354,N_2525,N_2317);
or UO_355 (O_355,N_2309,N_2913);
xor UO_356 (O_356,N_2281,N_2845);
nor UO_357 (O_357,N_2511,N_2420);
or UO_358 (O_358,N_2305,N_2519);
or UO_359 (O_359,N_2285,N_2553);
xnor UO_360 (O_360,N_2251,N_2931);
nand UO_361 (O_361,N_2602,N_2568);
and UO_362 (O_362,N_2673,N_2668);
nor UO_363 (O_363,N_2840,N_2779);
nand UO_364 (O_364,N_2559,N_2878);
and UO_365 (O_365,N_2688,N_2652);
nor UO_366 (O_366,N_2412,N_2505);
nand UO_367 (O_367,N_2272,N_2860);
and UO_368 (O_368,N_2728,N_2271);
nand UO_369 (O_369,N_2976,N_2962);
and UO_370 (O_370,N_2815,N_2621);
xor UO_371 (O_371,N_2936,N_2498);
nor UO_372 (O_372,N_2508,N_2473);
nor UO_373 (O_373,N_2657,N_2871);
or UO_374 (O_374,N_2280,N_2785);
nand UO_375 (O_375,N_2570,N_2562);
or UO_376 (O_376,N_2620,N_2662);
nor UO_377 (O_377,N_2388,N_2773);
or UO_378 (O_378,N_2309,N_2336);
and UO_379 (O_379,N_2805,N_2884);
nor UO_380 (O_380,N_2738,N_2571);
and UO_381 (O_381,N_2924,N_2936);
nand UO_382 (O_382,N_2779,N_2379);
nand UO_383 (O_383,N_2327,N_2916);
or UO_384 (O_384,N_2822,N_2785);
nor UO_385 (O_385,N_2435,N_2932);
nand UO_386 (O_386,N_2501,N_2785);
xor UO_387 (O_387,N_2574,N_2896);
nand UO_388 (O_388,N_2747,N_2810);
xnor UO_389 (O_389,N_2524,N_2353);
and UO_390 (O_390,N_2905,N_2443);
and UO_391 (O_391,N_2251,N_2827);
or UO_392 (O_392,N_2626,N_2700);
nand UO_393 (O_393,N_2476,N_2304);
nor UO_394 (O_394,N_2649,N_2267);
nand UO_395 (O_395,N_2906,N_2743);
nor UO_396 (O_396,N_2760,N_2353);
xnor UO_397 (O_397,N_2864,N_2872);
xnor UO_398 (O_398,N_2496,N_2726);
nor UO_399 (O_399,N_2418,N_2508);
and UO_400 (O_400,N_2843,N_2765);
nor UO_401 (O_401,N_2385,N_2994);
nand UO_402 (O_402,N_2981,N_2606);
nand UO_403 (O_403,N_2490,N_2930);
xor UO_404 (O_404,N_2301,N_2801);
and UO_405 (O_405,N_2948,N_2850);
nor UO_406 (O_406,N_2905,N_2496);
and UO_407 (O_407,N_2369,N_2803);
xor UO_408 (O_408,N_2473,N_2932);
xor UO_409 (O_409,N_2821,N_2588);
and UO_410 (O_410,N_2924,N_2770);
xnor UO_411 (O_411,N_2924,N_2854);
and UO_412 (O_412,N_2482,N_2457);
nor UO_413 (O_413,N_2395,N_2467);
nand UO_414 (O_414,N_2977,N_2941);
nand UO_415 (O_415,N_2634,N_2866);
xor UO_416 (O_416,N_2779,N_2901);
or UO_417 (O_417,N_2759,N_2554);
or UO_418 (O_418,N_2356,N_2543);
nand UO_419 (O_419,N_2918,N_2357);
or UO_420 (O_420,N_2975,N_2643);
nand UO_421 (O_421,N_2309,N_2761);
and UO_422 (O_422,N_2692,N_2254);
and UO_423 (O_423,N_2985,N_2929);
or UO_424 (O_424,N_2722,N_2601);
and UO_425 (O_425,N_2682,N_2567);
or UO_426 (O_426,N_2537,N_2975);
or UO_427 (O_427,N_2924,N_2645);
nand UO_428 (O_428,N_2525,N_2856);
xor UO_429 (O_429,N_2901,N_2431);
nand UO_430 (O_430,N_2928,N_2649);
or UO_431 (O_431,N_2764,N_2862);
and UO_432 (O_432,N_2736,N_2354);
xnor UO_433 (O_433,N_2746,N_2360);
nor UO_434 (O_434,N_2735,N_2547);
or UO_435 (O_435,N_2590,N_2801);
nor UO_436 (O_436,N_2441,N_2673);
or UO_437 (O_437,N_2762,N_2946);
or UO_438 (O_438,N_2939,N_2859);
or UO_439 (O_439,N_2301,N_2972);
and UO_440 (O_440,N_2388,N_2958);
nand UO_441 (O_441,N_2889,N_2853);
nor UO_442 (O_442,N_2883,N_2427);
and UO_443 (O_443,N_2733,N_2504);
xor UO_444 (O_444,N_2305,N_2301);
and UO_445 (O_445,N_2692,N_2532);
or UO_446 (O_446,N_2417,N_2648);
nor UO_447 (O_447,N_2396,N_2649);
xor UO_448 (O_448,N_2319,N_2784);
nand UO_449 (O_449,N_2591,N_2338);
or UO_450 (O_450,N_2882,N_2863);
xnor UO_451 (O_451,N_2866,N_2712);
nor UO_452 (O_452,N_2394,N_2831);
or UO_453 (O_453,N_2697,N_2746);
and UO_454 (O_454,N_2324,N_2812);
and UO_455 (O_455,N_2738,N_2813);
nor UO_456 (O_456,N_2500,N_2865);
or UO_457 (O_457,N_2610,N_2486);
and UO_458 (O_458,N_2259,N_2787);
xor UO_459 (O_459,N_2286,N_2319);
nand UO_460 (O_460,N_2310,N_2594);
nor UO_461 (O_461,N_2305,N_2971);
xor UO_462 (O_462,N_2428,N_2633);
nor UO_463 (O_463,N_2256,N_2532);
or UO_464 (O_464,N_2916,N_2500);
nor UO_465 (O_465,N_2283,N_2814);
or UO_466 (O_466,N_2762,N_2602);
xnor UO_467 (O_467,N_2308,N_2471);
nand UO_468 (O_468,N_2905,N_2997);
or UO_469 (O_469,N_2557,N_2831);
xor UO_470 (O_470,N_2639,N_2642);
nand UO_471 (O_471,N_2284,N_2995);
and UO_472 (O_472,N_2360,N_2315);
or UO_473 (O_473,N_2701,N_2438);
or UO_474 (O_474,N_2613,N_2619);
nor UO_475 (O_475,N_2619,N_2638);
nor UO_476 (O_476,N_2838,N_2590);
xnor UO_477 (O_477,N_2583,N_2600);
and UO_478 (O_478,N_2707,N_2611);
nor UO_479 (O_479,N_2287,N_2959);
xor UO_480 (O_480,N_2535,N_2270);
or UO_481 (O_481,N_2672,N_2335);
and UO_482 (O_482,N_2393,N_2452);
xnor UO_483 (O_483,N_2859,N_2999);
nand UO_484 (O_484,N_2590,N_2647);
xor UO_485 (O_485,N_2489,N_2532);
nor UO_486 (O_486,N_2940,N_2628);
nand UO_487 (O_487,N_2324,N_2765);
nand UO_488 (O_488,N_2535,N_2854);
nand UO_489 (O_489,N_2575,N_2448);
or UO_490 (O_490,N_2493,N_2638);
and UO_491 (O_491,N_2305,N_2734);
or UO_492 (O_492,N_2906,N_2839);
or UO_493 (O_493,N_2912,N_2583);
nor UO_494 (O_494,N_2318,N_2586);
nor UO_495 (O_495,N_2641,N_2955);
xnor UO_496 (O_496,N_2655,N_2795);
nand UO_497 (O_497,N_2751,N_2583);
nor UO_498 (O_498,N_2959,N_2530);
nand UO_499 (O_499,N_2326,N_2774);
endmodule