module basic_500_3000_500_6_levels_1xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_298,In_343);
and U1 (N_1,In_412,In_476);
and U2 (N_2,In_431,In_114);
and U3 (N_3,In_103,In_232);
and U4 (N_4,In_36,In_300);
and U5 (N_5,In_393,In_189);
nand U6 (N_6,In_165,In_29);
and U7 (N_7,In_489,In_54);
and U8 (N_8,In_321,In_310);
nand U9 (N_9,In_279,In_374);
nand U10 (N_10,In_311,In_244);
nand U11 (N_11,In_32,In_175);
and U12 (N_12,In_127,In_337);
nor U13 (N_13,In_149,In_87);
nor U14 (N_14,In_433,In_107);
nand U15 (N_15,In_1,In_88);
nor U16 (N_16,In_340,In_69);
and U17 (N_17,In_402,In_193);
nand U18 (N_18,In_330,In_483);
and U19 (N_19,In_62,In_58);
nor U20 (N_20,In_257,In_109);
or U21 (N_21,In_215,In_465);
or U22 (N_22,In_98,In_264);
and U23 (N_23,In_43,In_451);
nand U24 (N_24,In_450,In_275);
nor U25 (N_25,In_247,In_91);
nand U26 (N_26,In_185,In_28);
nand U27 (N_27,In_409,In_125);
nor U28 (N_28,In_205,In_394);
nor U29 (N_29,In_137,In_434);
or U30 (N_30,In_403,In_414);
or U31 (N_31,In_26,In_346);
and U32 (N_32,In_324,In_130);
or U33 (N_33,In_280,In_80);
and U34 (N_34,In_316,In_436);
nor U35 (N_35,In_372,In_376);
and U36 (N_36,In_268,In_25);
and U37 (N_37,In_482,In_435);
or U38 (N_38,In_235,In_77);
nand U39 (N_39,In_404,In_115);
nand U40 (N_40,In_56,In_371);
nor U41 (N_41,In_428,In_464);
nand U42 (N_42,In_240,In_475);
nor U43 (N_43,In_20,In_196);
nand U44 (N_44,In_288,In_242);
nand U45 (N_45,In_64,In_430);
nor U46 (N_46,In_407,In_363);
or U47 (N_47,In_417,In_128);
and U48 (N_48,In_273,In_454);
nand U49 (N_49,In_229,In_463);
or U50 (N_50,In_492,In_460);
xnor U51 (N_51,In_429,In_24);
and U52 (N_52,In_85,In_367);
xnor U53 (N_53,In_78,In_203);
nand U54 (N_54,In_283,In_361);
or U55 (N_55,In_124,In_270);
nor U56 (N_56,In_183,In_437);
nor U57 (N_57,In_16,In_142);
nand U58 (N_58,In_152,In_167);
nor U59 (N_59,In_491,In_369);
or U60 (N_60,In_269,In_466);
nor U61 (N_61,In_206,In_154);
nand U62 (N_62,In_220,In_89);
nor U63 (N_63,In_312,In_14);
and U64 (N_64,In_291,In_186);
nand U65 (N_65,In_117,In_397);
nor U66 (N_66,In_155,In_405);
nor U67 (N_67,In_19,In_234);
nor U68 (N_68,In_79,In_82);
nand U69 (N_69,In_216,In_471);
and U70 (N_70,In_163,In_325);
nand U71 (N_71,In_387,In_188);
and U72 (N_72,In_357,In_101);
nor U73 (N_73,In_76,In_131);
or U74 (N_74,In_256,In_329);
or U75 (N_75,In_105,In_418);
or U76 (N_76,In_45,In_389);
and U77 (N_77,In_478,In_219);
nor U78 (N_78,In_455,In_265);
or U79 (N_79,In_156,In_81);
nand U80 (N_80,In_453,In_495);
nand U81 (N_81,In_446,In_60);
nor U82 (N_82,In_97,In_364);
and U83 (N_83,In_208,In_135);
and U84 (N_84,In_116,In_170);
nand U85 (N_85,In_384,In_487);
nand U86 (N_86,In_222,In_334);
nand U87 (N_87,In_74,In_299);
or U88 (N_88,In_493,In_323);
and U89 (N_89,In_419,In_315);
xnor U90 (N_90,In_248,In_342);
and U91 (N_91,In_438,In_326);
nand U92 (N_92,In_192,In_339);
or U93 (N_93,In_285,In_11);
nor U94 (N_94,In_366,In_352);
nand U95 (N_95,In_319,In_295);
nor U96 (N_96,In_468,In_469);
and U97 (N_97,In_245,In_282);
nand U98 (N_98,In_249,In_160);
nand U99 (N_99,In_9,In_401);
or U100 (N_100,In_47,In_171);
nor U101 (N_101,In_210,In_44);
or U102 (N_102,In_217,In_182);
or U103 (N_103,In_383,In_306);
nor U104 (N_104,In_49,In_48);
or U105 (N_105,In_209,In_34);
nor U106 (N_106,In_61,In_95);
nand U107 (N_107,In_121,In_345);
nand U108 (N_108,In_94,In_174);
nor U109 (N_109,In_169,In_146);
nand U110 (N_110,In_370,In_253);
nor U111 (N_111,In_133,In_496);
and U112 (N_112,In_153,In_227);
nor U113 (N_113,In_486,In_309);
and U114 (N_114,In_301,In_31);
or U115 (N_115,In_379,In_444);
or U116 (N_116,In_138,In_373);
or U117 (N_117,In_66,In_349);
nand U118 (N_118,In_336,In_120);
or U119 (N_119,In_385,In_72);
or U120 (N_120,In_250,In_30);
nor U121 (N_121,In_427,In_314);
nor U122 (N_122,In_202,In_70);
and U123 (N_123,In_347,In_335);
nand U124 (N_124,In_259,In_195);
and U125 (N_125,In_37,In_328);
nor U126 (N_126,In_260,In_425);
xnor U127 (N_127,In_254,In_441);
nor U128 (N_128,In_447,In_246);
and U129 (N_129,In_477,In_302);
or U130 (N_130,In_375,In_168);
and U131 (N_131,In_184,In_327);
nand U132 (N_132,In_461,In_392);
nor U133 (N_133,In_129,In_2);
and U134 (N_134,In_12,In_83);
or U135 (N_135,In_65,In_17);
nor U136 (N_136,In_173,In_297);
nand U137 (N_137,In_6,In_200);
nor U138 (N_138,In_204,In_422);
or U139 (N_139,In_41,In_408);
nand U140 (N_140,In_225,In_7);
and U141 (N_141,In_424,In_307);
nor U142 (N_142,In_157,In_214);
nand U143 (N_143,In_462,In_172);
nor U144 (N_144,In_218,In_287);
nor U145 (N_145,In_176,In_318);
or U146 (N_146,In_488,In_150);
nand U147 (N_147,In_286,In_110);
and U148 (N_148,In_144,In_358);
xor U149 (N_149,In_399,In_191);
nand U150 (N_150,In_223,In_386);
and U151 (N_151,In_360,In_67);
nand U152 (N_152,In_320,In_395);
nand U153 (N_153,In_236,In_39);
nand U154 (N_154,In_481,In_166);
nand U155 (N_155,In_296,In_57);
or U156 (N_156,In_344,In_305);
nand U157 (N_157,In_415,In_426);
nand U158 (N_158,In_113,In_457);
nor U159 (N_159,In_178,In_106);
or U160 (N_160,In_239,In_377);
and U161 (N_161,In_0,In_151);
or U162 (N_162,In_52,In_499);
or U163 (N_163,In_22,In_241);
or U164 (N_164,In_33,In_304);
and U165 (N_165,In_388,In_252);
nor U166 (N_166,In_272,In_449);
nor U167 (N_167,In_255,In_490);
or U168 (N_168,In_3,In_458);
and U169 (N_169,In_293,In_46);
nor U170 (N_170,In_303,In_382);
and U171 (N_171,In_289,In_8);
or U172 (N_172,In_390,In_143);
or U173 (N_173,In_398,In_15);
and U174 (N_174,In_396,In_443);
or U175 (N_175,In_356,In_221);
nand U176 (N_176,In_145,In_442);
or U177 (N_177,In_132,In_140);
nor U178 (N_178,In_456,In_480);
and U179 (N_179,In_276,In_55);
nand U180 (N_180,In_262,In_452);
nand U181 (N_181,In_237,In_484);
nor U182 (N_182,In_84,In_365);
nor U183 (N_183,In_23,In_50);
nand U184 (N_184,In_277,In_148);
nor U185 (N_185,In_164,In_432);
nor U186 (N_186,In_292,In_212);
nand U187 (N_187,In_119,In_448);
nand U188 (N_188,In_359,In_35);
nand U189 (N_189,In_99,In_473);
nand U190 (N_190,In_134,In_93);
or U191 (N_191,In_368,In_263);
or U192 (N_192,In_421,In_51);
or U193 (N_193,In_181,In_420);
nand U194 (N_194,In_381,In_479);
or U195 (N_195,In_281,In_136);
nor U196 (N_196,In_472,In_224);
or U197 (N_197,In_238,In_86);
nor U198 (N_198,In_21,In_122);
or U199 (N_199,In_199,In_271);
or U200 (N_200,In_126,In_187);
and U201 (N_201,In_40,In_211);
or U202 (N_202,In_53,In_294);
nor U203 (N_203,In_179,In_118);
or U204 (N_204,In_42,In_104);
and U205 (N_205,In_362,In_333);
or U206 (N_206,In_96,In_351);
nand U207 (N_207,In_180,In_102);
nand U208 (N_208,In_213,In_338);
nor U209 (N_209,In_75,In_201);
nor U210 (N_210,In_13,In_228);
and U211 (N_211,In_158,In_38);
and U212 (N_212,In_226,In_284);
nand U213 (N_213,In_231,In_162);
and U214 (N_214,In_498,In_207);
or U215 (N_215,In_59,In_68);
nand U216 (N_216,In_378,In_413);
or U217 (N_217,In_341,In_177);
or U218 (N_218,In_348,In_350);
or U219 (N_219,In_410,In_190);
nor U220 (N_220,In_470,In_290);
nor U221 (N_221,In_90,In_258);
or U222 (N_222,In_251,In_355);
xor U223 (N_223,In_423,In_416);
nor U224 (N_224,In_406,In_439);
or U225 (N_225,In_5,In_100);
or U226 (N_226,In_63,In_497);
or U227 (N_227,In_467,In_274);
xor U228 (N_228,In_391,In_380);
nor U229 (N_229,In_159,In_10);
or U230 (N_230,In_243,In_18);
and U231 (N_231,In_108,In_332);
nor U232 (N_232,In_71,In_194);
nor U233 (N_233,In_123,In_278);
nand U234 (N_234,In_73,In_233);
or U235 (N_235,In_445,In_141);
nand U236 (N_236,In_112,In_331);
and U237 (N_237,In_261,In_147);
nor U238 (N_238,In_230,In_197);
nor U239 (N_239,In_411,In_494);
nor U240 (N_240,In_485,In_267);
nor U241 (N_241,In_474,In_313);
nor U242 (N_242,In_266,In_139);
nand U243 (N_243,In_322,In_111);
nor U244 (N_244,In_161,In_198);
xnor U245 (N_245,In_4,In_459);
and U246 (N_246,In_440,In_354);
nand U247 (N_247,In_308,In_92);
and U248 (N_248,In_353,In_400);
nand U249 (N_249,In_27,In_317);
nor U250 (N_250,In_176,In_316);
and U251 (N_251,In_89,In_86);
nor U252 (N_252,In_444,In_117);
nor U253 (N_253,In_470,In_498);
and U254 (N_254,In_239,In_182);
nor U255 (N_255,In_402,In_202);
nor U256 (N_256,In_378,In_331);
or U257 (N_257,In_112,In_113);
nand U258 (N_258,In_97,In_128);
and U259 (N_259,In_130,In_90);
and U260 (N_260,In_305,In_334);
nand U261 (N_261,In_429,In_108);
nor U262 (N_262,In_335,In_222);
and U263 (N_263,In_360,In_12);
and U264 (N_264,In_97,In_83);
nand U265 (N_265,In_429,In_325);
nand U266 (N_266,In_461,In_150);
nand U267 (N_267,In_428,In_353);
and U268 (N_268,In_181,In_414);
nor U269 (N_269,In_377,In_68);
nor U270 (N_270,In_19,In_299);
or U271 (N_271,In_356,In_214);
nor U272 (N_272,In_253,In_38);
nand U273 (N_273,In_61,In_232);
nor U274 (N_274,In_461,In_111);
nand U275 (N_275,In_37,In_458);
or U276 (N_276,In_36,In_49);
nand U277 (N_277,In_282,In_116);
or U278 (N_278,In_215,In_84);
or U279 (N_279,In_439,In_380);
nand U280 (N_280,In_59,In_274);
nand U281 (N_281,In_60,In_11);
nor U282 (N_282,In_141,In_216);
or U283 (N_283,In_32,In_124);
and U284 (N_284,In_112,In_2);
and U285 (N_285,In_331,In_276);
or U286 (N_286,In_109,In_387);
nand U287 (N_287,In_265,In_401);
or U288 (N_288,In_75,In_294);
and U289 (N_289,In_382,In_14);
and U290 (N_290,In_453,In_445);
or U291 (N_291,In_166,In_253);
nand U292 (N_292,In_486,In_110);
nor U293 (N_293,In_492,In_438);
or U294 (N_294,In_443,In_499);
and U295 (N_295,In_52,In_67);
and U296 (N_296,In_214,In_173);
nor U297 (N_297,In_361,In_262);
and U298 (N_298,In_137,In_485);
nand U299 (N_299,In_229,In_218);
nand U300 (N_300,In_453,In_231);
and U301 (N_301,In_446,In_96);
or U302 (N_302,In_424,In_35);
or U303 (N_303,In_406,In_282);
or U304 (N_304,In_7,In_405);
nor U305 (N_305,In_106,In_445);
or U306 (N_306,In_243,In_103);
or U307 (N_307,In_492,In_175);
nand U308 (N_308,In_12,In_109);
or U309 (N_309,In_489,In_260);
and U310 (N_310,In_57,In_83);
nand U311 (N_311,In_396,In_475);
nand U312 (N_312,In_319,In_90);
nand U313 (N_313,In_167,In_44);
nor U314 (N_314,In_4,In_256);
nor U315 (N_315,In_397,In_262);
and U316 (N_316,In_311,In_456);
nand U317 (N_317,In_428,In_387);
and U318 (N_318,In_218,In_152);
and U319 (N_319,In_356,In_432);
and U320 (N_320,In_184,In_366);
nor U321 (N_321,In_207,In_486);
nor U322 (N_322,In_163,In_247);
and U323 (N_323,In_176,In_136);
nand U324 (N_324,In_231,In_383);
nand U325 (N_325,In_332,In_264);
nand U326 (N_326,In_180,In_124);
nor U327 (N_327,In_66,In_98);
or U328 (N_328,In_494,In_299);
or U329 (N_329,In_25,In_336);
and U330 (N_330,In_151,In_384);
and U331 (N_331,In_77,In_368);
and U332 (N_332,In_104,In_337);
and U333 (N_333,In_7,In_324);
nand U334 (N_334,In_409,In_86);
nand U335 (N_335,In_20,In_293);
or U336 (N_336,In_263,In_264);
and U337 (N_337,In_37,In_99);
and U338 (N_338,In_60,In_185);
or U339 (N_339,In_131,In_377);
and U340 (N_340,In_217,In_220);
nor U341 (N_341,In_402,In_257);
or U342 (N_342,In_224,In_109);
nand U343 (N_343,In_328,In_279);
nor U344 (N_344,In_155,In_346);
or U345 (N_345,In_344,In_156);
nor U346 (N_346,In_81,In_482);
or U347 (N_347,In_372,In_262);
nor U348 (N_348,In_6,In_307);
and U349 (N_349,In_268,In_415);
xor U350 (N_350,In_44,In_304);
nand U351 (N_351,In_32,In_322);
nor U352 (N_352,In_430,In_213);
and U353 (N_353,In_16,In_307);
nand U354 (N_354,In_144,In_88);
nor U355 (N_355,In_141,In_276);
nand U356 (N_356,In_479,In_180);
or U357 (N_357,In_321,In_248);
or U358 (N_358,In_117,In_336);
or U359 (N_359,In_245,In_50);
or U360 (N_360,In_133,In_10);
and U361 (N_361,In_433,In_445);
and U362 (N_362,In_356,In_120);
nand U363 (N_363,In_402,In_120);
and U364 (N_364,In_470,In_443);
nor U365 (N_365,In_341,In_325);
or U366 (N_366,In_165,In_312);
nand U367 (N_367,In_24,In_277);
nand U368 (N_368,In_208,In_161);
and U369 (N_369,In_230,In_0);
and U370 (N_370,In_157,In_354);
and U371 (N_371,In_370,In_73);
nor U372 (N_372,In_194,In_358);
nand U373 (N_373,In_153,In_253);
or U374 (N_374,In_37,In_447);
or U375 (N_375,In_494,In_364);
and U376 (N_376,In_61,In_177);
nor U377 (N_377,In_442,In_300);
or U378 (N_378,In_93,In_153);
nand U379 (N_379,In_337,In_369);
nand U380 (N_380,In_278,In_263);
and U381 (N_381,In_305,In_488);
nor U382 (N_382,In_397,In_437);
nor U383 (N_383,In_210,In_224);
and U384 (N_384,In_199,In_295);
nand U385 (N_385,In_451,In_118);
nor U386 (N_386,In_351,In_68);
and U387 (N_387,In_299,In_396);
nor U388 (N_388,In_55,In_287);
nor U389 (N_389,In_354,In_302);
nand U390 (N_390,In_262,In_194);
nand U391 (N_391,In_378,In_274);
or U392 (N_392,In_266,In_367);
or U393 (N_393,In_91,In_4);
and U394 (N_394,In_311,In_400);
nand U395 (N_395,In_377,In_440);
nand U396 (N_396,In_101,In_324);
nor U397 (N_397,In_261,In_191);
or U398 (N_398,In_439,In_256);
nor U399 (N_399,In_132,In_460);
and U400 (N_400,In_13,In_8);
and U401 (N_401,In_220,In_495);
and U402 (N_402,In_106,In_383);
nand U403 (N_403,In_227,In_134);
and U404 (N_404,In_181,In_310);
or U405 (N_405,In_177,In_357);
and U406 (N_406,In_245,In_133);
and U407 (N_407,In_225,In_75);
nor U408 (N_408,In_139,In_166);
or U409 (N_409,In_360,In_242);
and U410 (N_410,In_32,In_128);
nor U411 (N_411,In_31,In_97);
or U412 (N_412,In_475,In_334);
and U413 (N_413,In_364,In_221);
nor U414 (N_414,In_254,In_128);
and U415 (N_415,In_322,In_479);
or U416 (N_416,In_183,In_34);
or U417 (N_417,In_316,In_386);
and U418 (N_418,In_49,In_198);
or U419 (N_419,In_436,In_54);
or U420 (N_420,In_16,In_264);
nand U421 (N_421,In_133,In_450);
and U422 (N_422,In_243,In_229);
and U423 (N_423,In_215,In_154);
and U424 (N_424,In_73,In_48);
nor U425 (N_425,In_116,In_399);
nand U426 (N_426,In_276,In_81);
or U427 (N_427,In_122,In_431);
nand U428 (N_428,In_225,In_409);
nand U429 (N_429,In_303,In_89);
nand U430 (N_430,In_34,In_496);
or U431 (N_431,In_257,In_337);
nand U432 (N_432,In_395,In_182);
nor U433 (N_433,In_263,In_66);
and U434 (N_434,In_26,In_239);
nor U435 (N_435,In_217,In_50);
nor U436 (N_436,In_337,In_362);
nor U437 (N_437,In_239,In_234);
nand U438 (N_438,In_460,In_102);
or U439 (N_439,In_43,In_91);
nand U440 (N_440,In_179,In_455);
nand U441 (N_441,In_292,In_81);
xnor U442 (N_442,In_54,In_203);
nand U443 (N_443,In_80,In_407);
nand U444 (N_444,In_26,In_159);
and U445 (N_445,In_181,In_485);
nand U446 (N_446,In_137,In_297);
nand U447 (N_447,In_315,In_395);
and U448 (N_448,In_264,In_386);
nor U449 (N_449,In_13,In_349);
nand U450 (N_450,In_215,In_26);
nor U451 (N_451,In_346,In_413);
nand U452 (N_452,In_215,In_64);
nand U453 (N_453,In_66,In_449);
or U454 (N_454,In_285,In_152);
and U455 (N_455,In_163,In_157);
nor U456 (N_456,In_133,In_384);
or U457 (N_457,In_482,In_366);
nand U458 (N_458,In_59,In_326);
nand U459 (N_459,In_333,In_217);
and U460 (N_460,In_151,In_298);
nand U461 (N_461,In_476,In_283);
nor U462 (N_462,In_206,In_95);
nand U463 (N_463,In_212,In_91);
and U464 (N_464,In_462,In_306);
or U465 (N_465,In_71,In_5);
nor U466 (N_466,In_266,In_99);
nand U467 (N_467,In_209,In_421);
nand U468 (N_468,In_295,In_267);
nand U469 (N_469,In_104,In_351);
nand U470 (N_470,In_335,In_285);
nand U471 (N_471,In_410,In_202);
nor U472 (N_472,In_245,In_167);
and U473 (N_473,In_18,In_141);
and U474 (N_474,In_454,In_328);
or U475 (N_475,In_241,In_340);
and U476 (N_476,In_438,In_74);
nor U477 (N_477,In_163,In_40);
nand U478 (N_478,In_413,In_106);
and U479 (N_479,In_101,In_105);
nor U480 (N_480,In_294,In_300);
nand U481 (N_481,In_45,In_133);
or U482 (N_482,In_173,In_27);
or U483 (N_483,In_154,In_392);
and U484 (N_484,In_308,In_341);
and U485 (N_485,In_177,In_191);
nor U486 (N_486,In_318,In_488);
and U487 (N_487,In_452,In_325);
and U488 (N_488,In_454,In_129);
nor U489 (N_489,In_45,In_324);
nand U490 (N_490,In_329,In_214);
or U491 (N_491,In_470,In_196);
nand U492 (N_492,In_450,In_118);
nand U493 (N_493,In_244,In_222);
and U494 (N_494,In_396,In_74);
and U495 (N_495,In_454,In_427);
or U496 (N_496,In_369,In_40);
nand U497 (N_497,In_414,In_465);
and U498 (N_498,In_54,In_76);
and U499 (N_499,In_440,In_459);
and U500 (N_500,N_108,N_345);
nor U501 (N_501,N_82,N_368);
xor U502 (N_502,N_208,N_68);
nand U503 (N_503,N_412,N_118);
nand U504 (N_504,N_361,N_121);
or U505 (N_505,N_396,N_229);
or U506 (N_506,N_239,N_308);
or U507 (N_507,N_314,N_426);
or U508 (N_508,N_437,N_191);
and U509 (N_509,N_321,N_451);
nand U510 (N_510,N_42,N_417);
xor U511 (N_511,N_182,N_416);
nand U512 (N_512,N_401,N_240);
and U513 (N_513,N_178,N_414);
nor U514 (N_514,N_370,N_445);
or U515 (N_515,N_277,N_187);
nand U516 (N_516,N_70,N_129);
nand U517 (N_517,N_474,N_325);
and U518 (N_518,N_464,N_226);
nand U519 (N_519,N_433,N_48);
and U520 (N_520,N_334,N_337);
or U521 (N_521,N_80,N_267);
or U522 (N_522,N_181,N_293);
nand U523 (N_523,N_307,N_406);
and U524 (N_524,N_348,N_237);
nor U525 (N_525,N_31,N_106);
nor U526 (N_526,N_104,N_372);
and U527 (N_527,N_304,N_490);
nor U528 (N_528,N_351,N_193);
nor U529 (N_529,N_312,N_477);
nor U530 (N_530,N_492,N_17);
or U531 (N_531,N_319,N_327);
nand U532 (N_532,N_256,N_263);
nand U533 (N_533,N_50,N_26);
nand U534 (N_534,N_405,N_364);
nand U535 (N_535,N_461,N_134);
nor U536 (N_536,N_192,N_303);
and U537 (N_537,N_421,N_484);
nor U538 (N_538,N_436,N_206);
nand U539 (N_539,N_39,N_144);
or U540 (N_540,N_167,N_175);
or U541 (N_541,N_79,N_404);
nand U542 (N_542,N_491,N_169);
nor U543 (N_543,N_360,N_328);
nand U544 (N_544,N_36,N_194);
or U545 (N_545,N_148,N_349);
or U546 (N_546,N_411,N_95);
nor U547 (N_547,N_60,N_232);
nor U548 (N_548,N_216,N_305);
nand U549 (N_549,N_205,N_18);
or U550 (N_550,N_282,N_90);
nor U551 (N_551,N_183,N_51);
or U552 (N_552,N_107,N_330);
and U553 (N_553,N_355,N_210);
and U554 (N_554,N_21,N_71);
nor U555 (N_555,N_362,N_499);
nor U556 (N_556,N_440,N_266);
and U557 (N_557,N_352,N_343);
and U558 (N_558,N_94,N_16);
and U559 (N_559,N_62,N_127);
or U560 (N_560,N_165,N_201);
nor U561 (N_561,N_139,N_469);
or U562 (N_562,N_120,N_222);
nand U563 (N_563,N_151,N_119);
nor U564 (N_564,N_10,N_297);
nand U565 (N_565,N_3,N_238);
nand U566 (N_566,N_84,N_443);
nor U567 (N_567,N_137,N_203);
nand U568 (N_568,N_11,N_311);
and U569 (N_569,N_444,N_13);
nand U570 (N_570,N_369,N_125);
nand U571 (N_571,N_313,N_158);
xor U572 (N_572,N_176,N_301);
nand U573 (N_573,N_248,N_14);
and U574 (N_574,N_448,N_264);
and U575 (N_575,N_109,N_468);
or U576 (N_576,N_381,N_149);
or U577 (N_577,N_154,N_56);
nand U578 (N_578,N_278,N_57);
nor U579 (N_579,N_259,N_171);
or U580 (N_580,N_66,N_427);
nor U581 (N_581,N_389,N_476);
nor U582 (N_582,N_449,N_124);
nand U583 (N_583,N_460,N_415);
or U584 (N_584,N_288,N_2);
nor U585 (N_585,N_397,N_77);
or U586 (N_586,N_27,N_43);
nor U587 (N_587,N_49,N_418);
nand U588 (N_588,N_356,N_115);
and U589 (N_589,N_399,N_447);
nor U590 (N_590,N_174,N_338);
nand U591 (N_591,N_329,N_22);
and U592 (N_592,N_41,N_357);
nand U593 (N_593,N_392,N_315);
and U594 (N_594,N_497,N_473);
nand U595 (N_595,N_466,N_92);
or U596 (N_596,N_353,N_153);
or U597 (N_597,N_280,N_195);
nor U598 (N_598,N_4,N_310);
nor U599 (N_599,N_88,N_215);
and U600 (N_600,N_33,N_61);
xnor U601 (N_601,N_130,N_471);
nand U602 (N_602,N_20,N_424);
nand U603 (N_603,N_391,N_454);
or U604 (N_604,N_28,N_196);
nor U605 (N_605,N_385,N_204);
nand U606 (N_606,N_260,N_365);
and U607 (N_607,N_270,N_12);
nor U608 (N_608,N_489,N_177);
or U609 (N_609,N_441,N_331);
nor U610 (N_610,N_133,N_91);
and U611 (N_611,N_367,N_220);
nor U612 (N_612,N_488,N_89);
nand U613 (N_613,N_253,N_413);
and U614 (N_614,N_258,N_480);
nand U615 (N_615,N_463,N_1);
nand U616 (N_616,N_211,N_379);
and U617 (N_617,N_387,N_35);
or U618 (N_618,N_294,N_218);
and U619 (N_619,N_147,N_230);
and U620 (N_620,N_431,N_111);
or U621 (N_621,N_390,N_105);
and U622 (N_622,N_213,N_261);
xor U623 (N_623,N_332,N_67);
nor U624 (N_624,N_287,N_428);
nor U625 (N_625,N_117,N_197);
nor U626 (N_626,N_141,N_281);
nor U627 (N_627,N_96,N_470);
or U628 (N_628,N_407,N_429);
nand U629 (N_629,N_273,N_52);
nor U630 (N_630,N_296,N_241);
and U631 (N_631,N_457,N_340);
nand U632 (N_632,N_190,N_402);
and U633 (N_633,N_252,N_157);
and U634 (N_634,N_112,N_378);
nand U635 (N_635,N_170,N_45);
nand U636 (N_636,N_212,N_6);
or U637 (N_637,N_185,N_8);
nor U638 (N_638,N_317,N_452);
nor U639 (N_639,N_269,N_344);
nor U640 (N_640,N_64,N_453);
nor U641 (N_641,N_300,N_347);
or U642 (N_642,N_209,N_236);
nor U643 (N_643,N_65,N_54);
or U644 (N_644,N_290,N_366);
nand U645 (N_645,N_496,N_446);
or U646 (N_646,N_335,N_7);
nand U647 (N_647,N_246,N_122);
nand U648 (N_648,N_359,N_113);
or U649 (N_649,N_32,N_225);
and U650 (N_650,N_101,N_69);
nand U651 (N_651,N_63,N_333);
nor U652 (N_652,N_25,N_168);
or U653 (N_653,N_254,N_99);
nand U654 (N_654,N_495,N_382);
or U655 (N_655,N_493,N_155);
and U656 (N_656,N_373,N_383);
nand U657 (N_657,N_494,N_386);
or U658 (N_658,N_318,N_156);
nor U659 (N_659,N_326,N_47);
and U660 (N_660,N_180,N_339);
nand U661 (N_661,N_255,N_73);
and U662 (N_662,N_419,N_336);
or U663 (N_663,N_250,N_143);
and U664 (N_664,N_102,N_245);
and U665 (N_665,N_83,N_423);
nor U666 (N_666,N_87,N_276);
or U667 (N_667,N_324,N_5);
nand U668 (N_668,N_75,N_78);
nand U669 (N_669,N_15,N_59);
nand U670 (N_670,N_159,N_482);
or U671 (N_671,N_161,N_409);
and U672 (N_672,N_408,N_29);
or U673 (N_673,N_403,N_410);
and U674 (N_674,N_286,N_189);
and U675 (N_675,N_374,N_114);
nor U676 (N_676,N_234,N_478);
and U677 (N_677,N_486,N_291);
nor U678 (N_678,N_432,N_376);
or U679 (N_679,N_465,N_430);
and U680 (N_680,N_289,N_214);
nor U681 (N_681,N_46,N_103);
and U682 (N_682,N_298,N_462);
nand U683 (N_683,N_173,N_322);
nand U684 (N_684,N_199,N_132);
xor U685 (N_685,N_74,N_450);
nand U686 (N_686,N_126,N_400);
nand U687 (N_687,N_274,N_320);
nand U688 (N_688,N_323,N_19);
nor U689 (N_689,N_242,N_24);
nor U690 (N_690,N_309,N_140);
nor U691 (N_691,N_467,N_98);
and U692 (N_692,N_93,N_9);
nor U693 (N_693,N_420,N_72);
nor U694 (N_694,N_142,N_86);
nor U695 (N_695,N_354,N_145);
or U696 (N_696,N_123,N_439);
and U697 (N_697,N_58,N_275);
xnor U698 (N_698,N_76,N_316);
and U699 (N_699,N_341,N_283);
or U700 (N_700,N_247,N_38);
nor U701 (N_701,N_395,N_223);
nand U702 (N_702,N_380,N_188);
or U703 (N_703,N_377,N_224);
nand U704 (N_704,N_302,N_162);
or U705 (N_705,N_388,N_136);
nand U706 (N_706,N_217,N_186);
nor U707 (N_707,N_375,N_172);
nand U708 (N_708,N_479,N_342);
nor U709 (N_709,N_55,N_160);
nor U710 (N_710,N_44,N_422);
nand U711 (N_711,N_306,N_53);
nor U712 (N_712,N_146,N_292);
and U713 (N_713,N_37,N_251);
or U714 (N_714,N_350,N_163);
or U715 (N_715,N_244,N_358);
nor U716 (N_716,N_200,N_425);
and U717 (N_717,N_262,N_23);
nand U718 (N_718,N_498,N_166);
nor U719 (N_719,N_472,N_243);
nor U720 (N_720,N_268,N_202);
nand U721 (N_721,N_458,N_257);
and U722 (N_722,N_299,N_475);
nor U723 (N_723,N_34,N_295);
and U724 (N_724,N_221,N_81);
nor U725 (N_725,N_456,N_442);
nor U726 (N_726,N_231,N_198);
nor U727 (N_727,N_135,N_279);
or U728 (N_728,N_435,N_271);
and U729 (N_729,N_438,N_393);
nand U730 (N_730,N_265,N_284);
or U731 (N_731,N_272,N_434);
nor U732 (N_732,N_138,N_235);
nor U733 (N_733,N_485,N_179);
nor U734 (N_734,N_100,N_131);
and U735 (N_735,N_285,N_249);
nor U736 (N_736,N_227,N_398);
nand U737 (N_737,N_371,N_85);
and U738 (N_738,N_164,N_128);
nand U739 (N_739,N_116,N_455);
and U740 (N_740,N_363,N_346);
and U741 (N_741,N_233,N_30);
nand U742 (N_742,N_483,N_97);
and U743 (N_743,N_394,N_110);
nand U744 (N_744,N_184,N_219);
and U745 (N_745,N_0,N_152);
or U746 (N_746,N_150,N_384);
or U747 (N_747,N_459,N_207);
and U748 (N_748,N_487,N_228);
or U749 (N_749,N_481,N_40);
and U750 (N_750,N_374,N_212);
and U751 (N_751,N_76,N_498);
nor U752 (N_752,N_447,N_389);
or U753 (N_753,N_226,N_222);
and U754 (N_754,N_385,N_268);
nand U755 (N_755,N_242,N_32);
and U756 (N_756,N_453,N_394);
and U757 (N_757,N_306,N_488);
and U758 (N_758,N_391,N_481);
or U759 (N_759,N_344,N_412);
and U760 (N_760,N_159,N_223);
nand U761 (N_761,N_301,N_118);
nor U762 (N_762,N_307,N_250);
and U763 (N_763,N_332,N_498);
and U764 (N_764,N_95,N_421);
nor U765 (N_765,N_451,N_32);
nand U766 (N_766,N_487,N_372);
or U767 (N_767,N_47,N_479);
nand U768 (N_768,N_254,N_330);
nor U769 (N_769,N_219,N_416);
nor U770 (N_770,N_184,N_227);
nor U771 (N_771,N_19,N_231);
nand U772 (N_772,N_23,N_461);
or U773 (N_773,N_4,N_358);
and U774 (N_774,N_379,N_157);
nand U775 (N_775,N_56,N_187);
nand U776 (N_776,N_119,N_83);
nand U777 (N_777,N_286,N_91);
nand U778 (N_778,N_459,N_227);
nand U779 (N_779,N_76,N_117);
nor U780 (N_780,N_35,N_349);
or U781 (N_781,N_287,N_433);
nor U782 (N_782,N_434,N_393);
nor U783 (N_783,N_276,N_209);
and U784 (N_784,N_286,N_127);
nand U785 (N_785,N_78,N_273);
nor U786 (N_786,N_481,N_281);
or U787 (N_787,N_194,N_384);
and U788 (N_788,N_128,N_470);
nor U789 (N_789,N_267,N_13);
and U790 (N_790,N_55,N_233);
nand U791 (N_791,N_364,N_246);
nand U792 (N_792,N_46,N_414);
nor U793 (N_793,N_297,N_418);
nor U794 (N_794,N_170,N_119);
or U795 (N_795,N_376,N_362);
nand U796 (N_796,N_158,N_288);
and U797 (N_797,N_241,N_394);
nand U798 (N_798,N_22,N_78);
nor U799 (N_799,N_440,N_222);
nor U800 (N_800,N_134,N_197);
nand U801 (N_801,N_254,N_421);
nand U802 (N_802,N_128,N_472);
nor U803 (N_803,N_303,N_36);
and U804 (N_804,N_290,N_461);
xnor U805 (N_805,N_28,N_431);
and U806 (N_806,N_206,N_189);
nor U807 (N_807,N_151,N_366);
nor U808 (N_808,N_306,N_425);
nand U809 (N_809,N_355,N_174);
nor U810 (N_810,N_54,N_213);
nand U811 (N_811,N_236,N_41);
and U812 (N_812,N_2,N_185);
nand U813 (N_813,N_167,N_222);
or U814 (N_814,N_262,N_498);
nand U815 (N_815,N_408,N_165);
nand U816 (N_816,N_147,N_212);
and U817 (N_817,N_399,N_183);
or U818 (N_818,N_68,N_152);
nand U819 (N_819,N_381,N_223);
and U820 (N_820,N_44,N_161);
nor U821 (N_821,N_391,N_73);
nor U822 (N_822,N_389,N_465);
nor U823 (N_823,N_218,N_196);
nand U824 (N_824,N_449,N_305);
nor U825 (N_825,N_78,N_51);
or U826 (N_826,N_400,N_47);
and U827 (N_827,N_386,N_208);
and U828 (N_828,N_320,N_362);
nor U829 (N_829,N_493,N_366);
nand U830 (N_830,N_301,N_108);
nor U831 (N_831,N_160,N_14);
or U832 (N_832,N_262,N_382);
nor U833 (N_833,N_495,N_302);
nor U834 (N_834,N_245,N_3);
nor U835 (N_835,N_314,N_439);
nand U836 (N_836,N_241,N_307);
nor U837 (N_837,N_65,N_166);
or U838 (N_838,N_285,N_146);
or U839 (N_839,N_186,N_224);
nor U840 (N_840,N_338,N_298);
xor U841 (N_841,N_72,N_113);
or U842 (N_842,N_6,N_236);
or U843 (N_843,N_259,N_187);
xor U844 (N_844,N_26,N_81);
and U845 (N_845,N_362,N_0);
nor U846 (N_846,N_466,N_462);
and U847 (N_847,N_387,N_252);
nor U848 (N_848,N_415,N_142);
nor U849 (N_849,N_242,N_403);
or U850 (N_850,N_190,N_148);
nor U851 (N_851,N_108,N_61);
nand U852 (N_852,N_300,N_123);
nor U853 (N_853,N_160,N_124);
and U854 (N_854,N_425,N_253);
nand U855 (N_855,N_467,N_269);
nor U856 (N_856,N_243,N_234);
nand U857 (N_857,N_386,N_394);
nand U858 (N_858,N_131,N_345);
and U859 (N_859,N_307,N_224);
or U860 (N_860,N_455,N_280);
nor U861 (N_861,N_166,N_215);
nand U862 (N_862,N_308,N_393);
nand U863 (N_863,N_151,N_195);
and U864 (N_864,N_257,N_155);
nand U865 (N_865,N_48,N_329);
nor U866 (N_866,N_97,N_211);
and U867 (N_867,N_106,N_304);
nor U868 (N_868,N_163,N_278);
or U869 (N_869,N_309,N_298);
and U870 (N_870,N_389,N_49);
and U871 (N_871,N_489,N_365);
and U872 (N_872,N_294,N_131);
nor U873 (N_873,N_403,N_238);
nor U874 (N_874,N_407,N_5);
nor U875 (N_875,N_431,N_153);
or U876 (N_876,N_459,N_252);
nor U877 (N_877,N_120,N_2);
or U878 (N_878,N_231,N_157);
nor U879 (N_879,N_425,N_340);
nor U880 (N_880,N_486,N_207);
nor U881 (N_881,N_282,N_5);
and U882 (N_882,N_483,N_480);
and U883 (N_883,N_196,N_392);
or U884 (N_884,N_499,N_163);
or U885 (N_885,N_483,N_393);
and U886 (N_886,N_132,N_315);
nand U887 (N_887,N_151,N_240);
and U888 (N_888,N_418,N_308);
or U889 (N_889,N_276,N_13);
or U890 (N_890,N_401,N_296);
nand U891 (N_891,N_458,N_3);
nand U892 (N_892,N_272,N_447);
or U893 (N_893,N_73,N_473);
and U894 (N_894,N_296,N_7);
nand U895 (N_895,N_192,N_497);
nor U896 (N_896,N_306,N_28);
xnor U897 (N_897,N_78,N_323);
and U898 (N_898,N_311,N_434);
nand U899 (N_899,N_115,N_21);
or U900 (N_900,N_212,N_19);
nand U901 (N_901,N_319,N_471);
nor U902 (N_902,N_201,N_332);
nor U903 (N_903,N_423,N_19);
nor U904 (N_904,N_355,N_279);
or U905 (N_905,N_269,N_114);
and U906 (N_906,N_472,N_140);
nor U907 (N_907,N_117,N_271);
nand U908 (N_908,N_298,N_79);
or U909 (N_909,N_61,N_447);
or U910 (N_910,N_241,N_32);
and U911 (N_911,N_123,N_11);
and U912 (N_912,N_13,N_401);
or U913 (N_913,N_21,N_429);
and U914 (N_914,N_143,N_331);
nor U915 (N_915,N_419,N_182);
and U916 (N_916,N_102,N_27);
and U917 (N_917,N_257,N_427);
or U918 (N_918,N_446,N_19);
and U919 (N_919,N_462,N_451);
and U920 (N_920,N_105,N_448);
or U921 (N_921,N_167,N_148);
and U922 (N_922,N_341,N_223);
and U923 (N_923,N_191,N_232);
or U924 (N_924,N_101,N_62);
nor U925 (N_925,N_178,N_465);
nand U926 (N_926,N_495,N_439);
or U927 (N_927,N_94,N_431);
nor U928 (N_928,N_282,N_188);
nor U929 (N_929,N_388,N_69);
and U930 (N_930,N_282,N_326);
or U931 (N_931,N_58,N_248);
or U932 (N_932,N_52,N_221);
nor U933 (N_933,N_121,N_365);
and U934 (N_934,N_100,N_476);
and U935 (N_935,N_317,N_371);
nor U936 (N_936,N_139,N_122);
nand U937 (N_937,N_385,N_193);
nor U938 (N_938,N_320,N_86);
or U939 (N_939,N_276,N_428);
nor U940 (N_940,N_168,N_398);
and U941 (N_941,N_300,N_137);
or U942 (N_942,N_218,N_110);
or U943 (N_943,N_427,N_399);
nand U944 (N_944,N_41,N_285);
or U945 (N_945,N_92,N_439);
nand U946 (N_946,N_94,N_341);
or U947 (N_947,N_497,N_459);
nand U948 (N_948,N_196,N_437);
xor U949 (N_949,N_316,N_291);
or U950 (N_950,N_253,N_324);
nand U951 (N_951,N_158,N_360);
nor U952 (N_952,N_214,N_394);
nand U953 (N_953,N_288,N_194);
nor U954 (N_954,N_312,N_292);
and U955 (N_955,N_417,N_370);
or U956 (N_956,N_17,N_444);
nor U957 (N_957,N_166,N_130);
or U958 (N_958,N_8,N_124);
nand U959 (N_959,N_156,N_228);
nand U960 (N_960,N_167,N_404);
nor U961 (N_961,N_281,N_8);
nand U962 (N_962,N_487,N_473);
and U963 (N_963,N_372,N_260);
or U964 (N_964,N_423,N_322);
nor U965 (N_965,N_64,N_374);
or U966 (N_966,N_165,N_197);
nand U967 (N_967,N_320,N_246);
xor U968 (N_968,N_448,N_345);
or U969 (N_969,N_226,N_67);
nand U970 (N_970,N_86,N_127);
nand U971 (N_971,N_35,N_494);
or U972 (N_972,N_419,N_324);
or U973 (N_973,N_380,N_219);
or U974 (N_974,N_465,N_151);
nor U975 (N_975,N_89,N_476);
nand U976 (N_976,N_437,N_406);
and U977 (N_977,N_317,N_168);
or U978 (N_978,N_483,N_173);
nor U979 (N_979,N_350,N_286);
nor U980 (N_980,N_115,N_86);
and U981 (N_981,N_163,N_463);
nand U982 (N_982,N_167,N_336);
and U983 (N_983,N_415,N_289);
or U984 (N_984,N_499,N_409);
and U985 (N_985,N_267,N_387);
or U986 (N_986,N_23,N_398);
or U987 (N_987,N_466,N_249);
and U988 (N_988,N_352,N_203);
and U989 (N_989,N_140,N_203);
and U990 (N_990,N_185,N_206);
nor U991 (N_991,N_217,N_151);
nand U992 (N_992,N_388,N_173);
nand U993 (N_993,N_112,N_440);
nor U994 (N_994,N_194,N_175);
nor U995 (N_995,N_76,N_273);
nor U996 (N_996,N_270,N_486);
or U997 (N_997,N_396,N_92);
nor U998 (N_998,N_361,N_451);
nor U999 (N_999,N_134,N_487);
and U1000 (N_1000,N_895,N_679);
or U1001 (N_1001,N_920,N_863);
nand U1002 (N_1002,N_781,N_577);
nor U1003 (N_1003,N_988,N_632);
nand U1004 (N_1004,N_866,N_598);
or U1005 (N_1005,N_543,N_756);
nor U1006 (N_1006,N_586,N_809);
or U1007 (N_1007,N_892,N_626);
nor U1008 (N_1008,N_842,N_827);
or U1009 (N_1009,N_891,N_942);
and U1010 (N_1010,N_867,N_785);
nand U1011 (N_1011,N_629,N_656);
or U1012 (N_1012,N_545,N_881);
nand U1013 (N_1013,N_735,N_528);
nor U1014 (N_1014,N_934,N_654);
nor U1015 (N_1015,N_771,N_912);
and U1016 (N_1016,N_535,N_683);
and U1017 (N_1017,N_906,N_864);
and U1018 (N_1018,N_713,N_753);
nor U1019 (N_1019,N_612,N_831);
nand U1020 (N_1020,N_986,N_611);
xnor U1021 (N_1021,N_798,N_633);
and U1022 (N_1022,N_599,N_525);
or U1023 (N_1023,N_605,N_813);
and U1024 (N_1024,N_759,N_662);
nand U1025 (N_1025,N_570,N_590);
and U1026 (N_1026,N_919,N_510);
nor U1027 (N_1027,N_954,N_976);
and U1028 (N_1028,N_932,N_925);
and U1029 (N_1029,N_663,N_806);
nor U1030 (N_1030,N_544,N_603);
nor U1031 (N_1031,N_928,N_747);
and U1032 (N_1032,N_989,N_826);
nand U1033 (N_1033,N_847,N_762);
and U1034 (N_1034,N_944,N_960);
nand U1035 (N_1035,N_969,N_768);
and U1036 (N_1036,N_873,N_896);
nor U1037 (N_1037,N_997,N_567);
nor U1038 (N_1038,N_961,N_608);
or U1039 (N_1039,N_914,N_744);
nand U1040 (N_1040,N_795,N_773);
and U1041 (N_1041,N_856,N_887);
nor U1042 (N_1042,N_623,N_999);
nand U1043 (N_1043,N_810,N_751);
and U1044 (N_1044,N_874,N_538);
and U1045 (N_1045,N_956,N_576);
or U1046 (N_1046,N_503,N_916);
nand U1047 (N_1047,N_651,N_898);
nor U1048 (N_1048,N_572,N_852);
nor U1049 (N_1049,N_804,N_776);
and U1050 (N_1050,N_950,N_647);
and U1051 (N_1051,N_834,N_921);
nand U1052 (N_1052,N_723,N_929);
nor U1053 (N_1053,N_573,N_500);
and U1054 (N_1054,N_837,N_615);
nand U1055 (N_1055,N_995,N_708);
nand U1056 (N_1056,N_861,N_696);
or U1057 (N_1057,N_924,N_522);
and U1058 (N_1058,N_902,N_689);
and U1059 (N_1059,N_560,N_981);
nor U1060 (N_1060,N_817,N_802);
xor U1061 (N_1061,N_565,N_564);
nor U1062 (N_1062,N_843,N_816);
and U1063 (N_1063,N_517,N_886);
nand U1064 (N_1064,N_641,N_774);
nor U1065 (N_1065,N_945,N_964);
or U1066 (N_1066,N_582,N_606);
or U1067 (N_1067,N_628,N_955);
or U1068 (N_1068,N_868,N_691);
nor U1069 (N_1069,N_501,N_716);
or U1070 (N_1070,N_515,N_855);
and U1071 (N_1071,N_659,N_669);
nor U1072 (N_1072,N_518,N_943);
and U1073 (N_1073,N_637,N_903);
and U1074 (N_1074,N_550,N_636);
or U1075 (N_1075,N_514,N_740);
nor U1076 (N_1076,N_521,N_765);
or U1077 (N_1077,N_504,N_549);
nor U1078 (N_1078,N_604,N_882);
or U1079 (N_1079,N_602,N_695);
or U1080 (N_1080,N_799,N_711);
or U1081 (N_1081,N_739,N_980);
nor U1082 (N_1082,N_678,N_959);
nor U1083 (N_1083,N_918,N_870);
nand U1084 (N_1084,N_542,N_951);
nand U1085 (N_1085,N_655,N_991);
and U1086 (N_1086,N_613,N_973);
or U1087 (N_1087,N_534,N_814);
nand U1088 (N_1088,N_748,N_650);
and U1089 (N_1089,N_539,N_645);
nor U1090 (N_1090,N_985,N_705);
nor U1091 (N_1091,N_783,N_936);
nand U1092 (N_1092,N_559,N_687);
nor U1093 (N_1093,N_766,N_984);
and U1094 (N_1094,N_622,N_899);
or U1095 (N_1095,N_832,N_931);
nand U1096 (N_1096,N_859,N_681);
or U1097 (N_1097,N_581,N_548);
nor U1098 (N_1098,N_523,N_509);
or U1099 (N_1099,N_725,N_835);
nand U1100 (N_1100,N_644,N_901);
or U1101 (N_1101,N_853,N_782);
or U1102 (N_1102,N_587,N_977);
nand U1103 (N_1103,N_600,N_734);
or U1104 (N_1104,N_619,N_697);
and U1105 (N_1105,N_682,N_851);
or U1106 (N_1106,N_524,N_718);
and U1107 (N_1107,N_822,N_738);
nor U1108 (N_1108,N_532,N_933);
or U1109 (N_1109,N_704,N_631);
or U1110 (N_1110,N_990,N_743);
and U1111 (N_1111,N_648,N_724);
nor U1112 (N_1112,N_583,N_967);
nor U1113 (N_1113,N_818,N_639);
nand U1114 (N_1114,N_888,N_878);
nor U1115 (N_1115,N_609,N_516);
and U1116 (N_1116,N_983,N_700);
nand U1117 (N_1117,N_607,N_601);
and U1118 (N_1118,N_927,N_812);
or U1119 (N_1119,N_975,N_833);
nor U1120 (N_1120,N_617,N_685);
or U1121 (N_1121,N_911,N_506);
xor U1122 (N_1122,N_800,N_953);
or U1123 (N_1123,N_665,N_701);
or U1124 (N_1124,N_915,N_917);
nand U1125 (N_1125,N_937,N_974);
or U1126 (N_1126,N_998,N_884);
and U1127 (N_1127,N_760,N_946);
and U1128 (N_1128,N_555,N_568);
and U1129 (N_1129,N_698,N_889);
nor U1130 (N_1130,N_963,N_792);
nor U1131 (N_1131,N_657,N_805);
nand U1132 (N_1132,N_846,N_947);
and U1133 (N_1133,N_820,N_894);
nand U1134 (N_1134,N_670,N_726);
and U1135 (N_1135,N_597,N_996);
nor U1136 (N_1136,N_923,N_883);
nand U1137 (N_1137,N_745,N_594);
nor U1138 (N_1138,N_869,N_746);
or U1139 (N_1139,N_571,N_758);
and U1140 (N_1140,N_703,N_780);
or U1141 (N_1141,N_970,N_618);
and U1142 (N_1142,N_763,N_652);
nand U1143 (N_1143,N_966,N_699);
or U1144 (N_1144,N_530,N_845);
and U1145 (N_1145,N_502,N_674);
or U1146 (N_1146,N_803,N_791);
or U1147 (N_1147,N_821,N_860);
nand U1148 (N_1148,N_558,N_592);
nor U1149 (N_1149,N_677,N_707);
and U1150 (N_1150,N_635,N_987);
or U1151 (N_1151,N_526,N_926);
nand U1152 (N_1152,N_513,N_625);
nand U1153 (N_1153,N_972,N_693);
and U1154 (N_1154,N_643,N_680);
nand U1155 (N_1155,N_938,N_624);
or U1156 (N_1156,N_710,N_880);
nor U1157 (N_1157,N_585,N_978);
or U1158 (N_1158,N_653,N_709);
nor U1159 (N_1159,N_640,N_939);
nor U1160 (N_1160,N_930,N_666);
nand U1161 (N_1161,N_540,N_507);
xor U1162 (N_1162,N_714,N_630);
or U1163 (N_1163,N_825,N_563);
nor U1164 (N_1164,N_819,N_958);
nor U1165 (N_1165,N_579,N_910);
nor U1166 (N_1166,N_547,N_553);
nand U1167 (N_1167,N_661,N_994);
nand U1168 (N_1168,N_672,N_569);
or U1169 (N_1169,N_556,N_638);
nor U1170 (N_1170,N_566,N_634);
or U1171 (N_1171,N_909,N_667);
nor U1172 (N_1172,N_658,N_589);
nor U1173 (N_1173,N_962,N_575);
or U1174 (N_1174,N_770,N_948);
nand U1175 (N_1175,N_764,N_900);
and U1176 (N_1176,N_720,N_775);
nor U1177 (N_1177,N_620,N_839);
or U1178 (N_1178,N_591,N_732);
nand U1179 (N_1179,N_536,N_907);
and U1180 (N_1180,N_777,N_527);
or U1181 (N_1181,N_574,N_684);
or U1182 (N_1182,N_801,N_757);
or U1183 (N_1183,N_840,N_529);
nor U1184 (N_1184,N_706,N_811);
and U1185 (N_1185,N_668,N_646);
nor U1186 (N_1186,N_541,N_596);
nand U1187 (N_1187,N_676,N_979);
and U1188 (N_1188,N_836,N_621);
nand U1189 (N_1189,N_971,N_787);
or U1190 (N_1190,N_686,N_779);
xnor U1191 (N_1191,N_824,N_849);
nand U1192 (N_1192,N_841,N_721);
and U1193 (N_1193,N_719,N_935);
xnor U1194 (N_1194,N_742,N_790);
or U1195 (N_1195,N_511,N_554);
nand U1196 (N_1196,N_561,N_858);
and U1197 (N_1197,N_844,N_904);
nand U1198 (N_1198,N_627,N_546);
and U1199 (N_1199,N_664,N_968);
or U1200 (N_1200,N_578,N_551);
or U1201 (N_1201,N_614,N_741);
or U1202 (N_1202,N_784,N_797);
or U1203 (N_1203,N_660,N_865);
and U1204 (N_1204,N_610,N_692);
nand U1205 (N_1205,N_728,N_702);
nand U1206 (N_1206,N_897,N_690);
nor U1207 (N_1207,N_727,N_673);
or U1208 (N_1208,N_731,N_830);
nand U1209 (N_1209,N_722,N_675);
or U1210 (N_1210,N_940,N_649);
and U1211 (N_1211,N_786,N_793);
nand U1212 (N_1212,N_890,N_941);
nor U1213 (N_1213,N_828,N_580);
nand U1214 (N_1214,N_694,N_755);
or U1215 (N_1215,N_922,N_557);
nand U1216 (N_1216,N_688,N_761);
and U1217 (N_1217,N_769,N_715);
or U1218 (N_1218,N_562,N_992);
nor U1219 (N_1219,N_584,N_750);
and U1220 (N_1220,N_616,N_519);
nand U1221 (N_1221,N_512,N_794);
xor U1222 (N_1222,N_877,N_885);
nor U1223 (N_1223,N_533,N_908);
or U1224 (N_1224,N_796,N_850);
nand U1225 (N_1225,N_862,N_807);
or U1226 (N_1226,N_593,N_730);
and U1227 (N_1227,N_808,N_712);
nand U1228 (N_1228,N_982,N_893);
nand U1229 (N_1229,N_729,N_505);
and U1230 (N_1230,N_531,N_736);
or U1231 (N_1231,N_752,N_552);
nor U1232 (N_1232,N_854,N_789);
nand U1233 (N_1233,N_879,N_949);
and U1234 (N_1234,N_717,N_588);
nand U1235 (N_1235,N_733,N_508);
or U1236 (N_1236,N_913,N_871);
or U1237 (N_1237,N_778,N_815);
or U1238 (N_1238,N_848,N_829);
nand U1239 (N_1239,N_788,N_952);
nand U1240 (N_1240,N_876,N_857);
nor U1241 (N_1241,N_737,N_993);
nor U1242 (N_1242,N_767,N_965);
nand U1243 (N_1243,N_671,N_772);
or U1244 (N_1244,N_872,N_905);
nand U1245 (N_1245,N_537,N_823);
and U1246 (N_1246,N_875,N_957);
nor U1247 (N_1247,N_595,N_749);
nor U1248 (N_1248,N_838,N_520);
nor U1249 (N_1249,N_642,N_754);
nand U1250 (N_1250,N_907,N_792);
or U1251 (N_1251,N_840,N_753);
and U1252 (N_1252,N_727,N_528);
or U1253 (N_1253,N_784,N_811);
and U1254 (N_1254,N_817,N_656);
nand U1255 (N_1255,N_666,N_777);
nor U1256 (N_1256,N_614,N_935);
or U1257 (N_1257,N_758,N_682);
nor U1258 (N_1258,N_512,N_624);
or U1259 (N_1259,N_646,N_985);
nand U1260 (N_1260,N_695,N_667);
nor U1261 (N_1261,N_978,N_676);
nor U1262 (N_1262,N_832,N_684);
nand U1263 (N_1263,N_891,N_810);
nand U1264 (N_1264,N_935,N_579);
and U1265 (N_1265,N_955,N_562);
or U1266 (N_1266,N_609,N_904);
or U1267 (N_1267,N_956,N_950);
nor U1268 (N_1268,N_671,N_515);
nor U1269 (N_1269,N_555,N_526);
or U1270 (N_1270,N_971,N_735);
nor U1271 (N_1271,N_708,N_556);
or U1272 (N_1272,N_585,N_756);
nor U1273 (N_1273,N_937,N_518);
nand U1274 (N_1274,N_540,N_838);
or U1275 (N_1275,N_837,N_960);
nor U1276 (N_1276,N_513,N_881);
nor U1277 (N_1277,N_993,N_527);
nand U1278 (N_1278,N_932,N_913);
nor U1279 (N_1279,N_617,N_926);
or U1280 (N_1280,N_904,N_695);
or U1281 (N_1281,N_692,N_657);
nor U1282 (N_1282,N_664,N_953);
nor U1283 (N_1283,N_661,N_838);
or U1284 (N_1284,N_974,N_990);
nand U1285 (N_1285,N_526,N_891);
and U1286 (N_1286,N_634,N_928);
and U1287 (N_1287,N_930,N_994);
and U1288 (N_1288,N_776,N_650);
or U1289 (N_1289,N_573,N_809);
and U1290 (N_1290,N_805,N_541);
and U1291 (N_1291,N_824,N_970);
or U1292 (N_1292,N_772,N_638);
nor U1293 (N_1293,N_553,N_590);
nand U1294 (N_1294,N_894,N_792);
nand U1295 (N_1295,N_573,N_585);
nand U1296 (N_1296,N_852,N_768);
nand U1297 (N_1297,N_953,N_819);
nand U1298 (N_1298,N_914,N_505);
nand U1299 (N_1299,N_573,N_745);
nor U1300 (N_1300,N_770,N_535);
and U1301 (N_1301,N_799,N_569);
or U1302 (N_1302,N_835,N_941);
nand U1303 (N_1303,N_595,N_999);
nand U1304 (N_1304,N_981,N_692);
nor U1305 (N_1305,N_549,N_671);
nor U1306 (N_1306,N_864,N_855);
and U1307 (N_1307,N_667,N_520);
nand U1308 (N_1308,N_511,N_872);
and U1309 (N_1309,N_683,N_667);
or U1310 (N_1310,N_570,N_971);
nor U1311 (N_1311,N_854,N_713);
nand U1312 (N_1312,N_794,N_971);
nand U1313 (N_1313,N_938,N_529);
or U1314 (N_1314,N_596,N_943);
or U1315 (N_1315,N_712,N_666);
or U1316 (N_1316,N_711,N_551);
or U1317 (N_1317,N_972,N_727);
or U1318 (N_1318,N_782,N_984);
nand U1319 (N_1319,N_535,N_698);
nor U1320 (N_1320,N_720,N_908);
nand U1321 (N_1321,N_874,N_714);
or U1322 (N_1322,N_600,N_725);
nand U1323 (N_1323,N_601,N_851);
nand U1324 (N_1324,N_532,N_979);
or U1325 (N_1325,N_739,N_535);
or U1326 (N_1326,N_829,N_999);
nor U1327 (N_1327,N_677,N_838);
or U1328 (N_1328,N_661,N_537);
or U1329 (N_1329,N_698,N_525);
and U1330 (N_1330,N_758,N_924);
and U1331 (N_1331,N_838,N_599);
or U1332 (N_1332,N_601,N_713);
and U1333 (N_1333,N_736,N_807);
or U1334 (N_1334,N_506,N_746);
nor U1335 (N_1335,N_648,N_769);
nor U1336 (N_1336,N_718,N_855);
nand U1337 (N_1337,N_729,N_724);
nor U1338 (N_1338,N_969,N_867);
nor U1339 (N_1339,N_871,N_652);
and U1340 (N_1340,N_704,N_964);
and U1341 (N_1341,N_755,N_936);
and U1342 (N_1342,N_953,N_679);
nand U1343 (N_1343,N_741,N_900);
and U1344 (N_1344,N_572,N_799);
nor U1345 (N_1345,N_734,N_799);
nand U1346 (N_1346,N_599,N_617);
xor U1347 (N_1347,N_893,N_874);
and U1348 (N_1348,N_585,N_653);
xnor U1349 (N_1349,N_642,N_948);
or U1350 (N_1350,N_844,N_709);
or U1351 (N_1351,N_707,N_634);
and U1352 (N_1352,N_777,N_900);
or U1353 (N_1353,N_503,N_919);
or U1354 (N_1354,N_898,N_668);
nor U1355 (N_1355,N_827,N_961);
or U1356 (N_1356,N_808,N_605);
nor U1357 (N_1357,N_525,N_578);
nand U1358 (N_1358,N_803,N_802);
or U1359 (N_1359,N_658,N_616);
or U1360 (N_1360,N_824,N_695);
nand U1361 (N_1361,N_713,N_732);
nor U1362 (N_1362,N_717,N_932);
or U1363 (N_1363,N_675,N_955);
nor U1364 (N_1364,N_972,N_793);
nand U1365 (N_1365,N_909,N_685);
nor U1366 (N_1366,N_976,N_590);
nand U1367 (N_1367,N_969,N_584);
nand U1368 (N_1368,N_507,N_898);
nand U1369 (N_1369,N_849,N_872);
and U1370 (N_1370,N_897,N_923);
or U1371 (N_1371,N_874,N_534);
nor U1372 (N_1372,N_739,N_743);
nor U1373 (N_1373,N_612,N_609);
and U1374 (N_1374,N_770,N_866);
nor U1375 (N_1375,N_812,N_679);
and U1376 (N_1376,N_566,N_564);
nor U1377 (N_1377,N_923,N_871);
nor U1378 (N_1378,N_939,N_866);
nand U1379 (N_1379,N_782,N_642);
nor U1380 (N_1380,N_549,N_834);
nand U1381 (N_1381,N_649,N_872);
nor U1382 (N_1382,N_862,N_625);
nand U1383 (N_1383,N_846,N_708);
nor U1384 (N_1384,N_759,N_534);
nand U1385 (N_1385,N_597,N_886);
and U1386 (N_1386,N_954,N_646);
nand U1387 (N_1387,N_548,N_992);
nand U1388 (N_1388,N_984,N_900);
nand U1389 (N_1389,N_570,N_886);
or U1390 (N_1390,N_574,N_519);
nor U1391 (N_1391,N_937,N_663);
nand U1392 (N_1392,N_741,N_976);
and U1393 (N_1393,N_506,N_740);
nand U1394 (N_1394,N_553,N_778);
xnor U1395 (N_1395,N_636,N_795);
nor U1396 (N_1396,N_800,N_585);
or U1397 (N_1397,N_538,N_718);
and U1398 (N_1398,N_820,N_884);
nor U1399 (N_1399,N_722,N_664);
and U1400 (N_1400,N_647,N_519);
nor U1401 (N_1401,N_509,N_706);
nand U1402 (N_1402,N_692,N_843);
and U1403 (N_1403,N_861,N_597);
and U1404 (N_1404,N_825,N_770);
or U1405 (N_1405,N_676,N_535);
or U1406 (N_1406,N_845,N_858);
or U1407 (N_1407,N_517,N_625);
nor U1408 (N_1408,N_538,N_692);
nor U1409 (N_1409,N_848,N_660);
and U1410 (N_1410,N_995,N_693);
and U1411 (N_1411,N_513,N_571);
nand U1412 (N_1412,N_707,N_776);
nor U1413 (N_1413,N_541,N_976);
or U1414 (N_1414,N_647,N_774);
and U1415 (N_1415,N_661,N_691);
nand U1416 (N_1416,N_773,N_827);
nor U1417 (N_1417,N_593,N_976);
nor U1418 (N_1418,N_938,N_976);
nand U1419 (N_1419,N_741,N_571);
nand U1420 (N_1420,N_507,N_888);
nor U1421 (N_1421,N_798,N_781);
and U1422 (N_1422,N_860,N_778);
and U1423 (N_1423,N_711,N_504);
nand U1424 (N_1424,N_559,N_858);
and U1425 (N_1425,N_730,N_771);
nor U1426 (N_1426,N_512,N_921);
and U1427 (N_1427,N_997,N_673);
nand U1428 (N_1428,N_716,N_824);
or U1429 (N_1429,N_952,N_967);
nand U1430 (N_1430,N_988,N_684);
nand U1431 (N_1431,N_948,N_769);
and U1432 (N_1432,N_906,N_538);
nand U1433 (N_1433,N_935,N_722);
nand U1434 (N_1434,N_568,N_639);
xnor U1435 (N_1435,N_962,N_804);
or U1436 (N_1436,N_877,N_732);
and U1437 (N_1437,N_977,N_952);
nor U1438 (N_1438,N_924,N_742);
nor U1439 (N_1439,N_984,N_873);
nor U1440 (N_1440,N_508,N_959);
nand U1441 (N_1441,N_731,N_553);
or U1442 (N_1442,N_687,N_960);
and U1443 (N_1443,N_826,N_651);
nor U1444 (N_1444,N_748,N_763);
nand U1445 (N_1445,N_512,N_563);
nand U1446 (N_1446,N_592,N_596);
nand U1447 (N_1447,N_662,N_622);
or U1448 (N_1448,N_926,N_787);
and U1449 (N_1449,N_620,N_989);
nor U1450 (N_1450,N_589,N_945);
or U1451 (N_1451,N_840,N_895);
and U1452 (N_1452,N_775,N_737);
nor U1453 (N_1453,N_654,N_562);
nand U1454 (N_1454,N_692,N_812);
or U1455 (N_1455,N_779,N_529);
nand U1456 (N_1456,N_920,N_914);
nor U1457 (N_1457,N_773,N_791);
xnor U1458 (N_1458,N_735,N_595);
nand U1459 (N_1459,N_656,N_594);
nor U1460 (N_1460,N_912,N_809);
nand U1461 (N_1461,N_781,N_594);
and U1462 (N_1462,N_584,N_930);
or U1463 (N_1463,N_735,N_935);
and U1464 (N_1464,N_739,N_580);
nor U1465 (N_1465,N_535,N_704);
nor U1466 (N_1466,N_909,N_569);
nand U1467 (N_1467,N_919,N_901);
and U1468 (N_1468,N_998,N_591);
nand U1469 (N_1469,N_718,N_744);
nand U1470 (N_1470,N_927,N_673);
and U1471 (N_1471,N_675,N_747);
or U1472 (N_1472,N_654,N_917);
nor U1473 (N_1473,N_978,N_699);
nor U1474 (N_1474,N_968,N_516);
nand U1475 (N_1475,N_666,N_900);
or U1476 (N_1476,N_823,N_587);
and U1477 (N_1477,N_697,N_654);
or U1478 (N_1478,N_773,N_986);
or U1479 (N_1479,N_825,N_930);
and U1480 (N_1480,N_735,N_868);
xnor U1481 (N_1481,N_556,N_845);
or U1482 (N_1482,N_619,N_526);
and U1483 (N_1483,N_767,N_543);
and U1484 (N_1484,N_682,N_905);
and U1485 (N_1485,N_648,N_758);
nor U1486 (N_1486,N_811,N_694);
nor U1487 (N_1487,N_931,N_864);
and U1488 (N_1488,N_525,N_985);
nor U1489 (N_1489,N_781,N_573);
or U1490 (N_1490,N_754,N_703);
and U1491 (N_1491,N_734,N_893);
nand U1492 (N_1492,N_599,N_880);
nand U1493 (N_1493,N_892,N_583);
or U1494 (N_1494,N_551,N_875);
or U1495 (N_1495,N_503,N_866);
nand U1496 (N_1496,N_925,N_797);
and U1497 (N_1497,N_772,N_694);
and U1498 (N_1498,N_659,N_608);
nor U1499 (N_1499,N_814,N_965);
or U1500 (N_1500,N_1130,N_1330);
nor U1501 (N_1501,N_1292,N_1029);
nor U1502 (N_1502,N_1228,N_1472);
nor U1503 (N_1503,N_1202,N_1038);
nand U1504 (N_1504,N_1063,N_1105);
and U1505 (N_1505,N_1271,N_1093);
nand U1506 (N_1506,N_1272,N_1416);
and U1507 (N_1507,N_1434,N_1327);
or U1508 (N_1508,N_1408,N_1142);
nand U1509 (N_1509,N_1139,N_1156);
and U1510 (N_1510,N_1109,N_1265);
or U1511 (N_1511,N_1147,N_1134);
nor U1512 (N_1512,N_1457,N_1005);
nand U1513 (N_1513,N_1468,N_1192);
nand U1514 (N_1514,N_1369,N_1480);
nand U1515 (N_1515,N_1396,N_1390);
and U1516 (N_1516,N_1388,N_1169);
or U1517 (N_1517,N_1240,N_1184);
nand U1518 (N_1518,N_1489,N_1064);
and U1519 (N_1519,N_1232,N_1027);
or U1520 (N_1520,N_1441,N_1471);
nor U1521 (N_1521,N_1190,N_1333);
or U1522 (N_1522,N_1309,N_1291);
and U1523 (N_1523,N_1280,N_1487);
or U1524 (N_1524,N_1306,N_1371);
nor U1525 (N_1525,N_1338,N_1188);
or U1526 (N_1526,N_1001,N_1322);
nand U1527 (N_1527,N_1117,N_1294);
nand U1528 (N_1528,N_1079,N_1279);
and U1529 (N_1529,N_1124,N_1080);
nand U1530 (N_1530,N_1435,N_1128);
or U1531 (N_1531,N_1082,N_1494);
or U1532 (N_1532,N_1380,N_1421);
nor U1533 (N_1533,N_1177,N_1493);
and U1534 (N_1534,N_1496,N_1159);
nand U1535 (N_1535,N_1165,N_1164);
or U1536 (N_1536,N_1437,N_1400);
or U1537 (N_1537,N_1049,N_1497);
nor U1538 (N_1538,N_1384,N_1483);
and U1539 (N_1539,N_1211,N_1004);
and U1540 (N_1540,N_1344,N_1321);
nand U1541 (N_1541,N_1474,N_1368);
nand U1542 (N_1542,N_1436,N_1178);
and U1543 (N_1543,N_1351,N_1432);
and U1544 (N_1544,N_1254,N_1046);
nand U1545 (N_1545,N_1060,N_1170);
or U1546 (N_1546,N_1357,N_1106);
nand U1547 (N_1547,N_1449,N_1256);
or U1548 (N_1548,N_1405,N_1462);
nor U1549 (N_1549,N_1212,N_1348);
and U1550 (N_1550,N_1205,N_1023);
nor U1551 (N_1551,N_1347,N_1477);
nor U1552 (N_1552,N_1073,N_1255);
nor U1553 (N_1553,N_1055,N_1131);
and U1554 (N_1554,N_1331,N_1197);
and U1555 (N_1555,N_1041,N_1445);
nand U1556 (N_1556,N_1375,N_1206);
and U1557 (N_1557,N_1218,N_1207);
nor U1558 (N_1558,N_1334,N_1310);
or U1559 (N_1559,N_1411,N_1492);
or U1560 (N_1560,N_1168,N_1026);
nand U1561 (N_1561,N_1266,N_1373);
or U1562 (N_1562,N_1267,N_1329);
nor U1563 (N_1563,N_1446,N_1141);
and U1564 (N_1564,N_1340,N_1094);
nor U1565 (N_1565,N_1158,N_1448);
and U1566 (N_1566,N_1070,N_1013);
and U1567 (N_1567,N_1398,N_1113);
or U1568 (N_1568,N_1420,N_1459);
and U1569 (N_1569,N_1418,N_1257);
nand U1570 (N_1570,N_1378,N_1428);
and U1571 (N_1571,N_1059,N_1018);
or U1572 (N_1572,N_1006,N_1406);
and U1573 (N_1573,N_1253,N_1458);
and U1574 (N_1574,N_1083,N_1008);
nor U1575 (N_1575,N_1074,N_1163);
and U1576 (N_1576,N_1157,N_1189);
nor U1577 (N_1577,N_1431,N_1403);
and U1578 (N_1578,N_1311,N_1374);
nor U1579 (N_1579,N_1176,N_1488);
and U1580 (N_1580,N_1098,N_1215);
nand U1581 (N_1581,N_1221,N_1414);
or U1582 (N_1582,N_1456,N_1412);
nor U1583 (N_1583,N_1317,N_1498);
nand U1584 (N_1584,N_1103,N_1440);
and U1585 (N_1585,N_1076,N_1243);
and U1586 (N_1586,N_1182,N_1315);
nand U1587 (N_1587,N_1484,N_1187);
nor U1588 (N_1588,N_1146,N_1316);
and U1589 (N_1589,N_1166,N_1479);
nand U1590 (N_1590,N_1324,N_1282);
nor U1591 (N_1591,N_1033,N_1068);
or U1592 (N_1592,N_1464,N_1425);
or U1593 (N_1593,N_1423,N_1236);
and U1594 (N_1594,N_1478,N_1352);
nand U1595 (N_1595,N_1220,N_1495);
and U1596 (N_1596,N_1290,N_1143);
and U1597 (N_1597,N_1328,N_1057);
and U1598 (N_1598,N_1210,N_1318);
or U1599 (N_1599,N_1119,N_1360);
or U1600 (N_1600,N_1248,N_1410);
and U1601 (N_1601,N_1230,N_1090);
or U1602 (N_1602,N_1470,N_1066);
and U1603 (N_1603,N_1081,N_1469);
and U1604 (N_1604,N_1299,N_1237);
or U1605 (N_1605,N_1071,N_1454);
or U1606 (N_1606,N_1407,N_1426);
nand U1607 (N_1607,N_1002,N_1343);
and U1608 (N_1608,N_1288,N_1439);
nand U1609 (N_1609,N_1012,N_1115);
nor U1610 (N_1610,N_1376,N_1224);
and U1611 (N_1611,N_1377,N_1427);
nand U1612 (N_1612,N_1155,N_1121);
nand U1613 (N_1613,N_1302,N_1089);
nand U1614 (N_1614,N_1028,N_1137);
nor U1615 (N_1615,N_1171,N_1020);
or U1616 (N_1616,N_1335,N_1465);
or U1617 (N_1617,N_1138,N_1091);
nor U1618 (N_1618,N_1096,N_1017);
nand U1619 (N_1619,N_1153,N_1185);
and U1620 (N_1620,N_1261,N_1429);
and U1621 (N_1621,N_1350,N_1251);
nor U1622 (N_1622,N_1056,N_1490);
xor U1623 (N_1623,N_1363,N_1362);
nor U1624 (N_1624,N_1194,N_1172);
or U1625 (N_1625,N_1175,N_1241);
nor U1626 (N_1626,N_1140,N_1305);
nor U1627 (N_1627,N_1387,N_1499);
and U1628 (N_1628,N_1450,N_1107);
and U1629 (N_1629,N_1354,N_1397);
nand U1630 (N_1630,N_1133,N_1278);
and U1631 (N_1631,N_1009,N_1413);
nand U1632 (N_1632,N_1295,N_1225);
or U1633 (N_1633,N_1162,N_1148);
nor U1634 (N_1634,N_1067,N_1249);
nand U1635 (N_1635,N_1246,N_1264);
and U1636 (N_1636,N_1000,N_1303);
or U1637 (N_1637,N_1036,N_1275);
nor U1638 (N_1638,N_1242,N_1053);
or U1639 (N_1639,N_1003,N_1262);
nor U1640 (N_1640,N_1084,N_1342);
and U1641 (N_1641,N_1011,N_1268);
nand U1642 (N_1642,N_1095,N_1393);
nor U1643 (N_1643,N_1485,N_1438);
nand U1644 (N_1644,N_1208,N_1379);
and U1645 (N_1645,N_1307,N_1269);
nor U1646 (N_1646,N_1409,N_1135);
or U1647 (N_1647,N_1301,N_1419);
or U1648 (N_1648,N_1092,N_1451);
nand U1649 (N_1649,N_1108,N_1223);
and U1650 (N_1650,N_1200,N_1024);
and U1651 (N_1651,N_1238,N_1402);
nand U1652 (N_1652,N_1136,N_1010);
or U1653 (N_1653,N_1149,N_1424);
nand U1654 (N_1654,N_1195,N_1120);
and U1655 (N_1655,N_1281,N_1179);
or U1656 (N_1656,N_1222,N_1078);
or U1657 (N_1657,N_1442,N_1300);
nor U1658 (N_1658,N_1312,N_1346);
or U1659 (N_1659,N_1122,N_1355);
nand U1660 (N_1660,N_1100,N_1482);
nor U1661 (N_1661,N_1048,N_1326);
and U1662 (N_1662,N_1198,N_1389);
or U1663 (N_1663,N_1069,N_1339);
nor U1664 (N_1664,N_1430,N_1394);
or U1665 (N_1665,N_1042,N_1235);
nor U1666 (N_1666,N_1160,N_1250);
nor U1667 (N_1667,N_1452,N_1144);
nor U1668 (N_1668,N_1461,N_1399);
nand U1669 (N_1669,N_1116,N_1463);
or U1670 (N_1670,N_1286,N_1319);
nor U1671 (N_1671,N_1353,N_1088);
nand U1672 (N_1672,N_1021,N_1025);
and U1673 (N_1673,N_1051,N_1385);
nor U1674 (N_1674,N_1132,N_1356);
nor U1675 (N_1675,N_1129,N_1361);
nand U1676 (N_1676,N_1433,N_1320);
nor U1677 (N_1677,N_1337,N_1030);
and U1678 (N_1678,N_1382,N_1112);
and U1679 (N_1679,N_1453,N_1386);
nor U1680 (N_1680,N_1359,N_1101);
nand U1681 (N_1681,N_1031,N_1467);
and U1682 (N_1682,N_1022,N_1481);
and U1683 (N_1683,N_1044,N_1443);
and U1684 (N_1684,N_1364,N_1150);
or U1685 (N_1685,N_1277,N_1476);
nor U1686 (N_1686,N_1199,N_1161);
xor U1687 (N_1687,N_1231,N_1422);
nor U1688 (N_1688,N_1263,N_1077);
or U1689 (N_1689,N_1314,N_1110);
or U1690 (N_1690,N_1007,N_1270);
nand U1691 (N_1691,N_1287,N_1118);
nor U1692 (N_1692,N_1173,N_1383);
nand U1693 (N_1693,N_1114,N_1234);
nor U1694 (N_1694,N_1391,N_1058);
and U1695 (N_1695,N_1219,N_1447);
or U1696 (N_1696,N_1372,N_1154);
or U1697 (N_1697,N_1336,N_1039);
and U1698 (N_1698,N_1325,N_1313);
nand U1699 (N_1699,N_1019,N_1181);
or U1700 (N_1700,N_1061,N_1045);
or U1701 (N_1701,N_1104,N_1349);
nor U1702 (N_1702,N_1304,N_1050);
nand U1703 (N_1703,N_1111,N_1216);
nand U1704 (N_1704,N_1460,N_1415);
nor U1705 (N_1705,N_1259,N_1284);
nand U1706 (N_1706,N_1308,N_1473);
and U1707 (N_1707,N_1099,N_1125);
or U1708 (N_1708,N_1035,N_1401);
and U1709 (N_1709,N_1167,N_1047);
and U1710 (N_1710,N_1323,N_1475);
or U1711 (N_1711,N_1126,N_1367);
nand U1712 (N_1712,N_1404,N_1151);
nand U1713 (N_1713,N_1332,N_1054);
and U1714 (N_1714,N_1486,N_1040);
or U1715 (N_1715,N_1193,N_1203);
or U1716 (N_1716,N_1014,N_1183);
nand U1717 (N_1717,N_1097,N_1227);
or U1718 (N_1718,N_1201,N_1085);
nand U1719 (N_1719,N_1252,N_1075);
nor U1720 (N_1720,N_1417,N_1209);
nand U1721 (N_1721,N_1226,N_1296);
nor U1722 (N_1722,N_1358,N_1062);
and U1723 (N_1723,N_1217,N_1273);
and U1724 (N_1724,N_1127,N_1087);
and U1725 (N_1725,N_1444,N_1298);
and U1726 (N_1726,N_1214,N_1072);
and U1727 (N_1727,N_1260,N_1086);
nor U1728 (N_1728,N_1037,N_1244);
or U1729 (N_1729,N_1289,N_1345);
nand U1730 (N_1730,N_1065,N_1196);
or U1731 (N_1731,N_1395,N_1258);
nor U1732 (N_1732,N_1123,N_1245);
nand U1733 (N_1733,N_1043,N_1293);
nand U1734 (N_1734,N_1145,N_1466);
nand U1735 (N_1735,N_1276,N_1186);
or U1736 (N_1736,N_1034,N_1285);
or U1737 (N_1737,N_1274,N_1102);
or U1738 (N_1738,N_1191,N_1052);
or U1739 (N_1739,N_1370,N_1341);
nor U1740 (N_1740,N_1365,N_1015);
nand U1741 (N_1741,N_1032,N_1366);
xnor U1742 (N_1742,N_1381,N_1239);
and U1743 (N_1743,N_1204,N_1174);
nand U1744 (N_1744,N_1016,N_1297);
nand U1745 (N_1745,N_1229,N_1247);
and U1746 (N_1746,N_1213,N_1455);
nor U1747 (N_1747,N_1180,N_1392);
or U1748 (N_1748,N_1283,N_1152);
and U1749 (N_1749,N_1491,N_1233);
and U1750 (N_1750,N_1255,N_1289);
nor U1751 (N_1751,N_1456,N_1403);
nand U1752 (N_1752,N_1458,N_1313);
nand U1753 (N_1753,N_1180,N_1204);
nand U1754 (N_1754,N_1016,N_1304);
and U1755 (N_1755,N_1359,N_1157);
and U1756 (N_1756,N_1260,N_1211);
or U1757 (N_1757,N_1180,N_1279);
nand U1758 (N_1758,N_1414,N_1494);
and U1759 (N_1759,N_1175,N_1046);
nand U1760 (N_1760,N_1231,N_1337);
nand U1761 (N_1761,N_1161,N_1313);
nor U1762 (N_1762,N_1255,N_1208);
or U1763 (N_1763,N_1408,N_1212);
and U1764 (N_1764,N_1064,N_1386);
xor U1765 (N_1765,N_1416,N_1068);
nor U1766 (N_1766,N_1239,N_1272);
or U1767 (N_1767,N_1253,N_1105);
nor U1768 (N_1768,N_1419,N_1244);
nand U1769 (N_1769,N_1130,N_1013);
nand U1770 (N_1770,N_1181,N_1309);
nand U1771 (N_1771,N_1280,N_1418);
or U1772 (N_1772,N_1365,N_1400);
nor U1773 (N_1773,N_1223,N_1467);
and U1774 (N_1774,N_1132,N_1237);
and U1775 (N_1775,N_1022,N_1092);
nor U1776 (N_1776,N_1448,N_1256);
and U1777 (N_1777,N_1412,N_1028);
nand U1778 (N_1778,N_1319,N_1361);
or U1779 (N_1779,N_1282,N_1067);
nand U1780 (N_1780,N_1244,N_1267);
and U1781 (N_1781,N_1490,N_1019);
or U1782 (N_1782,N_1499,N_1257);
nor U1783 (N_1783,N_1000,N_1022);
and U1784 (N_1784,N_1020,N_1141);
or U1785 (N_1785,N_1145,N_1025);
nor U1786 (N_1786,N_1468,N_1295);
nand U1787 (N_1787,N_1388,N_1244);
nand U1788 (N_1788,N_1119,N_1497);
or U1789 (N_1789,N_1055,N_1339);
or U1790 (N_1790,N_1499,N_1254);
nor U1791 (N_1791,N_1089,N_1491);
nand U1792 (N_1792,N_1174,N_1056);
or U1793 (N_1793,N_1159,N_1314);
and U1794 (N_1794,N_1200,N_1381);
nand U1795 (N_1795,N_1104,N_1294);
or U1796 (N_1796,N_1238,N_1147);
nor U1797 (N_1797,N_1338,N_1128);
and U1798 (N_1798,N_1279,N_1453);
xnor U1799 (N_1799,N_1006,N_1264);
or U1800 (N_1800,N_1141,N_1094);
xor U1801 (N_1801,N_1004,N_1104);
and U1802 (N_1802,N_1222,N_1133);
nor U1803 (N_1803,N_1158,N_1473);
nor U1804 (N_1804,N_1426,N_1236);
nand U1805 (N_1805,N_1212,N_1170);
nand U1806 (N_1806,N_1335,N_1007);
and U1807 (N_1807,N_1013,N_1488);
and U1808 (N_1808,N_1043,N_1246);
and U1809 (N_1809,N_1436,N_1104);
and U1810 (N_1810,N_1410,N_1495);
nor U1811 (N_1811,N_1451,N_1456);
nand U1812 (N_1812,N_1383,N_1412);
nand U1813 (N_1813,N_1392,N_1327);
nor U1814 (N_1814,N_1014,N_1471);
or U1815 (N_1815,N_1116,N_1083);
nor U1816 (N_1816,N_1257,N_1046);
or U1817 (N_1817,N_1392,N_1137);
nor U1818 (N_1818,N_1095,N_1154);
nor U1819 (N_1819,N_1071,N_1120);
and U1820 (N_1820,N_1055,N_1340);
nor U1821 (N_1821,N_1141,N_1413);
or U1822 (N_1822,N_1248,N_1252);
nor U1823 (N_1823,N_1232,N_1152);
or U1824 (N_1824,N_1259,N_1096);
nand U1825 (N_1825,N_1108,N_1034);
nor U1826 (N_1826,N_1451,N_1168);
and U1827 (N_1827,N_1114,N_1057);
and U1828 (N_1828,N_1005,N_1269);
or U1829 (N_1829,N_1231,N_1002);
and U1830 (N_1830,N_1229,N_1144);
nor U1831 (N_1831,N_1492,N_1045);
nor U1832 (N_1832,N_1211,N_1119);
and U1833 (N_1833,N_1249,N_1170);
and U1834 (N_1834,N_1420,N_1317);
xor U1835 (N_1835,N_1361,N_1002);
and U1836 (N_1836,N_1277,N_1140);
or U1837 (N_1837,N_1093,N_1115);
or U1838 (N_1838,N_1095,N_1255);
nor U1839 (N_1839,N_1444,N_1484);
or U1840 (N_1840,N_1086,N_1408);
and U1841 (N_1841,N_1492,N_1184);
and U1842 (N_1842,N_1490,N_1043);
nor U1843 (N_1843,N_1417,N_1418);
or U1844 (N_1844,N_1171,N_1088);
or U1845 (N_1845,N_1199,N_1454);
or U1846 (N_1846,N_1457,N_1418);
nand U1847 (N_1847,N_1181,N_1412);
and U1848 (N_1848,N_1255,N_1225);
or U1849 (N_1849,N_1272,N_1025);
nand U1850 (N_1850,N_1195,N_1125);
nor U1851 (N_1851,N_1364,N_1304);
nand U1852 (N_1852,N_1090,N_1298);
or U1853 (N_1853,N_1337,N_1227);
nor U1854 (N_1854,N_1436,N_1105);
nor U1855 (N_1855,N_1080,N_1232);
nor U1856 (N_1856,N_1268,N_1365);
nor U1857 (N_1857,N_1078,N_1372);
and U1858 (N_1858,N_1058,N_1277);
nor U1859 (N_1859,N_1396,N_1000);
nor U1860 (N_1860,N_1457,N_1355);
and U1861 (N_1861,N_1399,N_1221);
nor U1862 (N_1862,N_1415,N_1457);
xnor U1863 (N_1863,N_1169,N_1277);
nand U1864 (N_1864,N_1007,N_1108);
nor U1865 (N_1865,N_1276,N_1470);
and U1866 (N_1866,N_1143,N_1153);
and U1867 (N_1867,N_1443,N_1078);
nand U1868 (N_1868,N_1155,N_1449);
nand U1869 (N_1869,N_1257,N_1461);
or U1870 (N_1870,N_1079,N_1071);
xnor U1871 (N_1871,N_1497,N_1271);
nand U1872 (N_1872,N_1209,N_1239);
and U1873 (N_1873,N_1204,N_1112);
nor U1874 (N_1874,N_1159,N_1458);
and U1875 (N_1875,N_1012,N_1290);
and U1876 (N_1876,N_1404,N_1442);
nor U1877 (N_1877,N_1324,N_1292);
and U1878 (N_1878,N_1149,N_1228);
or U1879 (N_1879,N_1113,N_1014);
nand U1880 (N_1880,N_1243,N_1294);
or U1881 (N_1881,N_1243,N_1335);
or U1882 (N_1882,N_1207,N_1132);
nand U1883 (N_1883,N_1324,N_1274);
or U1884 (N_1884,N_1338,N_1324);
nor U1885 (N_1885,N_1172,N_1240);
nand U1886 (N_1886,N_1101,N_1371);
or U1887 (N_1887,N_1195,N_1112);
or U1888 (N_1888,N_1421,N_1189);
and U1889 (N_1889,N_1496,N_1095);
nor U1890 (N_1890,N_1236,N_1463);
and U1891 (N_1891,N_1288,N_1386);
nor U1892 (N_1892,N_1171,N_1499);
or U1893 (N_1893,N_1496,N_1489);
nand U1894 (N_1894,N_1200,N_1032);
nand U1895 (N_1895,N_1094,N_1201);
and U1896 (N_1896,N_1424,N_1402);
nand U1897 (N_1897,N_1136,N_1256);
nor U1898 (N_1898,N_1357,N_1132);
or U1899 (N_1899,N_1487,N_1093);
or U1900 (N_1900,N_1481,N_1384);
nor U1901 (N_1901,N_1001,N_1009);
nand U1902 (N_1902,N_1115,N_1045);
and U1903 (N_1903,N_1172,N_1187);
and U1904 (N_1904,N_1324,N_1199);
and U1905 (N_1905,N_1093,N_1415);
or U1906 (N_1906,N_1330,N_1234);
nand U1907 (N_1907,N_1496,N_1230);
nand U1908 (N_1908,N_1250,N_1499);
nor U1909 (N_1909,N_1085,N_1253);
and U1910 (N_1910,N_1300,N_1074);
nand U1911 (N_1911,N_1134,N_1359);
or U1912 (N_1912,N_1071,N_1292);
and U1913 (N_1913,N_1332,N_1187);
nand U1914 (N_1914,N_1000,N_1340);
nand U1915 (N_1915,N_1179,N_1341);
nor U1916 (N_1916,N_1318,N_1440);
nand U1917 (N_1917,N_1445,N_1087);
nand U1918 (N_1918,N_1081,N_1368);
nand U1919 (N_1919,N_1132,N_1341);
or U1920 (N_1920,N_1259,N_1008);
nand U1921 (N_1921,N_1359,N_1108);
and U1922 (N_1922,N_1227,N_1020);
or U1923 (N_1923,N_1467,N_1370);
xnor U1924 (N_1924,N_1116,N_1020);
nor U1925 (N_1925,N_1215,N_1345);
nor U1926 (N_1926,N_1277,N_1111);
nor U1927 (N_1927,N_1053,N_1027);
nor U1928 (N_1928,N_1351,N_1327);
nor U1929 (N_1929,N_1023,N_1394);
and U1930 (N_1930,N_1054,N_1246);
or U1931 (N_1931,N_1214,N_1105);
and U1932 (N_1932,N_1366,N_1395);
and U1933 (N_1933,N_1335,N_1403);
or U1934 (N_1934,N_1313,N_1071);
nand U1935 (N_1935,N_1067,N_1109);
nor U1936 (N_1936,N_1382,N_1040);
nand U1937 (N_1937,N_1383,N_1177);
and U1938 (N_1938,N_1409,N_1177);
nor U1939 (N_1939,N_1103,N_1400);
and U1940 (N_1940,N_1424,N_1306);
or U1941 (N_1941,N_1434,N_1275);
and U1942 (N_1942,N_1270,N_1420);
nand U1943 (N_1943,N_1474,N_1216);
and U1944 (N_1944,N_1284,N_1129);
or U1945 (N_1945,N_1145,N_1381);
or U1946 (N_1946,N_1066,N_1025);
and U1947 (N_1947,N_1449,N_1402);
and U1948 (N_1948,N_1004,N_1412);
or U1949 (N_1949,N_1190,N_1025);
and U1950 (N_1950,N_1052,N_1314);
nand U1951 (N_1951,N_1419,N_1136);
nand U1952 (N_1952,N_1115,N_1440);
or U1953 (N_1953,N_1495,N_1000);
or U1954 (N_1954,N_1024,N_1377);
and U1955 (N_1955,N_1014,N_1451);
nand U1956 (N_1956,N_1228,N_1275);
nor U1957 (N_1957,N_1487,N_1045);
nor U1958 (N_1958,N_1407,N_1478);
nand U1959 (N_1959,N_1158,N_1316);
nor U1960 (N_1960,N_1161,N_1328);
xor U1961 (N_1961,N_1092,N_1079);
and U1962 (N_1962,N_1154,N_1146);
nand U1963 (N_1963,N_1444,N_1031);
nor U1964 (N_1964,N_1318,N_1084);
or U1965 (N_1965,N_1074,N_1155);
nor U1966 (N_1966,N_1164,N_1314);
or U1967 (N_1967,N_1387,N_1047);
and U1968 (N_1968,N_1447,N_1380);
and U1969 (N_1969,N_1235,N_1010);
nand U1970 (N_1970,N_1031,N_1377);
and U1971 (N_1971,N_1013,N_1198);
nand U1972 (N_1972,N_1268,N_1290);
and U1973 (N_1973,N_1273,N_1001);
nand U1974 (N_1974,N_1291,N_1053);
nor U1975 (N_1975,N_1216,N_1247);
and U1976 (N_1976,N_1463,N_1454);
nor U1977 (N_1977,N_1160,N_1325);
or U1978 (N_1978,N_1294,N_1066);
nor U1979 (N_1979,N_1317,N_1209);
and U1980 (N_1980,N_1058,N_1359);
and U1981 (N_1981,N_1010,N_1122);
and U1982 (N_1982,N_1162,N_1384);
nand U1983 (N_1983,N_1184,N_1093);
and U1984 (N_1984,N_1410,N_1144);
nor U1985 (N_1985,N_1134,N_1210);
nor U1986 (N_1986,N_1372,N_1461);
nor U1987 (N_1987,N_1006,N_1176);
and U1988 (N_1988,N_1045,N_1129);
nand U1989 (N_1989,N_1170,N_1121);
or U1990 (N_1990,N_1267,N_1399);
and U1991 (N_1991,N_1116,N_1374);
or U1992 (N_1992,N_1121,N_1400);
nor U1993 (N_1993,N_1471,N_1001);
or U1994 (N_1994,N_1030,N_1478);
or U1995 (N_1995,N_1117,N_1166);
or U1996 (N_1996,N_1417,N_1119);
nand U1997 (N_1997,N_1484,N_1015);
nand U1998 (N_1998,N_1037,N_1469);
nor U1999 (N_1999,N_1489,N_1269);
and U2000 (N_2000,N_1879,N_1817);
nor U2001 (N_2001,N_1683,N_1996);
nand U2002 (N_2002,N_1506,N_1829);
nand U2003 (N_2003,N_1516,N_1505);
or U2004 (N_2004,N_1566,N_1905);
or U2005 (N_2005,N_1990,N_1724);
or U2006 (N_2006,N_1735,N_1973);
and U2007 (N_2007,N_1748,N_1596);
nor U2008 (N_2008,N_1877,N_1605);
or U2009 (N_2009,N_1593,N_1772);
or U2010 (N_2010,N_1625,N_1921);
nor U2011 (N_2011,N_1843,N_1549);
or U2012 (N_2012,N_1894,N_1550);
nor U2013 (N_2013,N_1527,N_1552);
xnor U2014 (N_2014,N_1760,N_1776);
and U2015 (N_2015,N_1948,N_1531);
nand U2016 (N_2016,N_1989,N_1560);
nor U2017 (N_2017,N_1887,N_1547);
nand U2018 (N_2018,N_1753,N_1961);
or U2019 (N_2019,N_1876,N_1752);
nor U2020 (N_2020,N_1568,N_1640);
nand U2021 (N_2021,N_1974,N_1788);
nor U2022 (N_2022,N_1922,N_1624);
and U2023 (N_2023,N_1586,N_1738);
and U2024 (N_2024,N_1874,N_1626);
or U2025 (N_2025,N_1576,N_1662);
or U2026 (N_2026,N_1551,N_1591);
nand U2027 (N_2027,N_1813,N_1639);
and U2028 (N_2028,N_1627,N_1908);
nand U2029 (N_2029,N_1558,N_1595);
nand U2030 (N_2030,N_1691,N_1616);
xnor U2031 (N_2031,N_1925,N_1823);
nor U2032 (N_2032,N_1521,N_1722);
and U2033 (N_2033,N_1802,N_1953);
and U2034 (N_2034,N_1963,N_1962);
and U2035 (N_2035,N_1744,N_1597);
nand U2036 (N_2036,N_1617,N_1969);
nand U2037 (N_2037,N_1548,N_1573);
xor U2038 (N_2038,N_1808,N_1795);
nand U2039 (N_2039,N_1608,N_1806);
nand U2040 (N_2040,N_1858,N_1889);
and U2041 (N_2041,N_1733,N_1821);
nor U2042 (N_2042,N_1666,N_1682);
nor U2043 (N_2043,N_1863,N_1714);
and U2044 (N_2044,N_1717,N_1998);
or U2045 (N_2045,N_1827,N_1575);
and U2046 (N_2046,N_1931,N_1571);
or U2047 (N_2047,N_1898,N_1539);
or U2048 (N_2048,N_1705,N_1530);
and U2049 (N_2049,N_1517,N_1967);
nor U2050 (N_2050,N_1654,N_1728);
nor U2051 (N_2051,N_1762,N_1611);
or U2052 (N_2052,N_1901,N_1696);
nor U2053 (N_2053,N_1606,N_1871);
nand U2054 (N_2054,N_1747,N_1939);
nor U2055 (N_2055,N_1952,N_1833);
and U2056 (N_2056,N_1830,N_1656);
nor U2057 (N_2057,N_1870,N_1542);
nor U2058 (N_2058,N_1679,N_1950);
and U2059 (N_2059,N_1763,N_1859);
nor U2060 (N_2060,N_1756,N_1565);
nand U2061 (N_2061,N_1668,N_1839);
and U2062 (N_2062,N_1881,N_1731);
nand U2063 (N_2063,N_1522,N_1848);
and U2064 (N_2064,N_1884,N_1726);
or U2065 (N_2065,N_1604,N_1840);
and U2066 (N_2066,N_1955,N_1533);
nor U2067 (N_2067,N_1780,N_1792);
and U2068 (N_2068,N_1805,N_1867);
and U2069 (N_2069,N_1811,N_1592);
or U2070 (N_2070,N_1688,N_1966);
and U2071 (N_2071,N_1982,N_1510);
and U2072 (N_2072,N_1759,N_1750);
xor U2073 (N_2073,N_1997,N_1983);
nand U2074 (N_2074,N_1689,N_1652);
nand U2075 (N_2075,N_1826,N_1841);
nand U2076 (N_2076,N_1746,N_1959);
or U2077 (N_2077,N_1937,N_1873);
nor U2078 (N_2078,N_1562,N_1951);
nand U2079 (N_2079,N_1653,N_1799);
nor U2080 (N_2080,N_1754,N_1947);
and U2081 (N_2081,N_1540,N_1941);
nand U2082 (N_2082,N_1999,N_1984);
nor U2083 (N_2083,N_1703,N_1587);
or U2084 (N_2084,N_1701,N_1633);
nor U2085 (N_2085,N_1686,N_1559);
nand U2086 (N_2086,N_1651,N_1767);
nand U2087 (N_2087,N_1782,N_1872);
or U2088 (N_2088,N_1807,N_1720);
nor U2089 (N_2089,N_1786,N_1938);
or U2090 (N_2090,N_1890,N_1737);
nor U2091 (N_2091,N_1702,N_1642);
nor U2092 (N_2092,N_1958,N_1825);
nand U2093 (N_2093,N_1924,N_1553);
or U2094 (N_2094,N_1758,N_1866);
and U2095 (N_2095,N_1743,N_1646);
and U2096 (N_2096,N_1675,N_1897);
or U2097 (N_2097,N_1868,N_1920);
nor U2098 (N_2098,N_1790,N_1844);
nor U2099 (N_2099,N_1725,N_1512);
or U2100 (N_2100,N_1745,N_1561);
nor U2101 (N_2101,N_1658,N_1878);
nand U2102 (N_2102,N_1945,N_1892);
or U2103 (N_2103,N_1610,N_1800);
nand U2104 (N_2104,N_1797,N_1665);
or U2105 (N_2105,N_1578,N_1854);
or U2106 (N_2106,N_1770,N_1783);
nor U2107 (N_2107,N_1520,N_1956);
or U2108 (N_2108,N_1850,N_1710);
and U2109 (N_2109,N_1853,N_1957);
nand U2110 (N_2110,N_1534,N_1970);
nor U2111 (N_2111,N_1977,N_1557);
and U2112 (N_2112,N_1695,N_1532);
nor U2113 (N_2113,N_1971,N_1669);
nor U2114 (N_2114,N_1769,N_1768);
and U2115 (N_2115,N_1819,N_1960);
and U2116 (N_2116,N_1933,N_1875);
and U2117 (N_2117,N_1538,N_1932);
and U2118 (N_2118,N_1810,N_1609);
or U2119 (N_2119,N_1899,N_1739);
and U2120 (N_2120,N_1765,N_1985);
and U2121 (N_2121,N_1677,N_1755);
nand U2122 (N_2122,N_1991,N_1836);
nor U2123 (N_2123,N_1507,N_1647);
xor U2124 (N_2124,N_1523,N_1828);
or U2125 (N_2125,N_1599,N_1504);
nor U2126 (N_2126,N_1598,N_1700);
or U2127 (N_2127,N_1751,N_1981);
nand U2128 (N_2128,N_1775,N_1995);
and U2129 (N_2129,N_1911,N_1930);
or U2130 (N_2130,N_1661,N_1893);
nor U2131 (N_2131,N_1685,N_1513);
nor U2132 (N_2132,N_1741,N_1896);
and U2133 (N_2133,N_1988,N_1919);
nor U2134 (N_2134,N_1546,N_1706);
nor U2135 (N_2135,N_1734,N_1529);
or U2136 (N_2136,N_1729,N_1883);
nor U2137 (N_2137,N_1888,N_1926);
nand U2138 (N_2138,N_1508,N_1994);
nand U2139 (N_2139,N_1637,N_1614);
nor U2140 (N_2140,N_1612,N_1629);
nand U2141 (N_2141,N_1912,N_1917);
and U2142 (N_2142,N_1712,N_1992);
and U2143 (N_2143,N_1774,N_1655);
nor U2144 (N_2144,N_1902,N_1856);
and U2145 (N_2145,N_1946,N_1766);
or U2146 (N_2146,N_1906,N_1684);
and U2147 (N_2147,N_1928,N_1721);
nor U2148 (N_2148,N_1518,N_1537);
nor U2149 (N_2149,N_1690,N_1667);
and U2150 (N_2150,N_1944,N_1978);
and U2151 (N_2151,N_1727,N_1882);
or U2152 (N_2152,N_1972,N_1847);
or U2153 (N_2153,N_1601,N_1736);
nand U2154 (N_2154,N_1861,N_1880);
nand U2155 (N_2155,N_1923,N_1891);
and U2156 (N_2156,N_1832,N_1980);
nor U2157 (N_2157,N_1918,N_1670);
xor U2158 (N_2158,N_1694,N_1975);
nand U2159 (N_2159,N_1659,N_1818);
and U2160 (N_2160,N_1903,N_1812);
nand U2161 (N_2161,N_1641,N_1781);
nor U2162 (N_2162,N_1676,N_1968);
nand U2163 (N_2163,N_1509,N_1657);
and U2164 (N_2164,N_1784,N_1886);
nand U2165 (N_2165,N_1789,N_1663);
and U2166 (N_2166,N_1764,N_1628);
or U2167 (N_2167,N_1577,N_1773);
or U2168 (N_2168,N_1809,N_1620);
nor U2169 (N_2169,N_1622,N_1794);
or U2170 (N_2170,N_1778,N_1541);
nand U2171 (N_2171,N_1572,N_1555);
and U2172 (N_2172,N_1942,N_1916);
or U2173 (N_2173,N_1602,N_1680);
or U2174 (N_2174,N_1503,N_1954);
nand U2175 (N_2175,N_1849,N_1934);
and U2176 (N_2176,N_1525,N_1846);
and U2177 (N_2177,N_1927,N_1915);
nor U2178 (N_2178,N_1643,N_1619);
nor U2179 (N_2179,N_1708,N_1636);
and U2180 (N_2180,N_1793,N_1623);
nor U2181 (N_2181,N_1615,N_1771);
and U2182 (N_2182,N_1574,N_1822);
nor U2183 (N_2183,N_1835,N_1749);
and U2184 (N_2184,N_1965,N_1842);
or U2185 (N_2185,N_1579,N_1787);
nor U2186 (N_2186,N_1582,N_1979);
or U2187 (N_2187,N_1814,N_1885);
or U2188 (N_2188,N_1777,N_1940);
and U2189 (N_2189,N_1929,N_1943);
and U2190 (N_2190,N_1704,N_1693);
and U2191 (N_2191,N_1660,N_1649);
or U2192 (N_2192,N_1935,N_1528);
or U2193 (N_2193,N_1831,N_1820);
nor U2194 (N_2194,N_1590,N_1976);
nand U2195 (N_2195,N_1845,N_1564);
nor U2196 (N_2196,N_1709,N_1600);
and U2197 (N_2197,N_1570,N_1804);
nand U2198 (N_2198,N_1865,N_1993);
or U2199 (N_2199,N_1543,N_1904);
or U2200 (N_2200,N_1581,N_1502);
nor U2201 (N_2201,N_1650,N_1837);
nand U2202 (N_2202,N_1671,N_1757);
or U2203 (N_2203,N_1589,N_1986);
nor U2204 (N_2204,N_1511,N_1535);
nand U2205 (N_2205,N_1583,N_1664);
nand U2206 (N_2206,N_1618,N_1585);
and U2207 (N_2207,N_1588,N_1855);
nand U2208 (N_2208,N_1524,N_1803);
or U2209 (N_2209,N_1711,N_1514);
or U2210 (N_2210,N_1580,N_1678);
or U2211 (N_2211,N_1816,N_1613);
nand U2212 (N_2212,N_1909,N_1697);
nand U2213 (N_2213,N_1556,N_1723);
nor U2214 (N_2214,N_1900,N_1569);
or U2215 (N_2215,N_1544,N_1785);
nor U2216 (N_2216,N_1869,N_1718);
nor U2217 (N_2217,N_1914,N_1862);
nor U2218 (N_2218,N_1567,N_1895);
nor U2219 (N_2219,N_1698,N_1742);
or U2220 (N_2220,N_1607,N_1732);
and U2221 (N_2221,N_1964,N_1791);
nor U2222 (N_2222,N_1621,N_1913);
or U2223 (N_2223,N_1907,N_1936);
nor U2224 (N_2224,N_1864,N_1644);
or U2225 (N_2225,N_1536,N_1632);
and U2226 (N_2226,N_1987,N_1707);
nand U2227 (N_2227,N_1631,N_1672);
nand U2228 (N_2228,N_1515,N_1851);
nand U2229 (N_2229,N_1852,N_1519);
nor U2230 (N_2230,N_1815,N_1545);
or U2231 (N_2231,N_1687,N_1630);
nand U2232 (N_2232,N_1603,N_1634);
nor U2233 (N_2233,N_1681,N_1673);
and U2234 (N_2234,N_1584,N_1801);
nand U2235 (N_2235,N_1838,N_1500);
nor U2236 (N_2236,N_1857,N_1713);
nand U2237 (N_2237,N_1699,N_1779);
nor U2238 (N_2238,N_1740,N_1910);
or U2239 (N_2239,N_1716,N_1648);
nand U2240 (N_2240,N_1645,N_1834);
nor U2241 (N_2241,N_1554,N_1730);
nor U2242 (N_2242,N_1860,N_1824);
nand U2243 (N_2243,N_1674,N_1719);
nand U2244 (N_2244,N_1563,N_1761);
and U2245 (N_2245,N_1501,N_1715);
or U2246 (N_2246,N_1594,N_1692);
and U2247 (N_2247,N_1638,N_1798);
nand U2248 (N_2248,N_1949,N_1635);
nor U2249 (N_2249,N_1526,N_1796);
nand U2250 (N_2250,N_1833,N_1520);
or U2251 (N_2251,N_1979,N_1722);
or U2252 (N_2252,N_1717,N_1891);
nand U2253 (N_2253,N_1542,N_1983);
nand U2254 (N_2254,N_1596,N_1872);
and U2255 (N_2255,N_1576,N_1515);
nand U2256 (N_2256,N_1830,N_1838);
nor U2257 (N_2257,N_1591,N_1715);
and U2258 (N_2258,N_1983,N_1903);
or U2259 (N_2259,N_1529,N_1878);
nand U2260 (N_2260,N_1513,N_1792);
or U2261 (N_2261,N_1789,N_1862);
or U2262 (N_2262,N_1947,N_1976);
nand U2263 (N_2263,N_1956,N_1551);
nand U2264 (N_2264,N_1863,N_1907);
nand U2265 (N_2265,N_1547,N_1991);
xnor U2266 (N_2266,N_1684,N_1719);
or U2267 (N_2267,N_1685,N_1679);
and U2268 (N_2268,N_1856,N_1506);
nand U2269 (N_2269,N_1796,N_1979);
nand U2270 (N_2270,N_1526,N_1985);
or U2271 (N_2271,N_1514,N_1639);
and U2272 (N_2272,N_1735,N_1939);
and U2273 (N_2273,N_1611,N_1933);
nand U2274 (N_2274,N_1855,N_1570);
nor U2275 (N_2275,N_1535,N_1523);
nand U2276 (N_2276,N_1578,N_1803);
or U2277 (N_2277,N_1635,N_1730);
and U2278 (N_2278,N_1739,N_1814);
or U2279 (N_2279,N_1607,N_1835);
nand U2280 (N_2280,N_1793,N_1847);
and U2281 (N_2281,N_1531,N_1767);
and U2282 (N_2282,N_1869,N_1613);
nand U2283 (N_2283,N_1825,N_1688);
or U2284 (N_2284,N_1993,N_1620);
and U2285 (N_2285,N_1578,N_1934);
nor U2286 (N_2286,N_1941,N_1971);
nand U2287 (N_2287,N_1869,N_1745);
nand U2288 (N_2288,N_1529,N_1909);
or U2289 (N_2289,N_1664,N_1557);
and U2290 (N_2290,N_1791,N_1696);
and U2291 (N_2291,N_1587,N_1822);
nand U2292 (N_2292,N_1506,N_1972);
and U2293 (N_2293,N_1536,N_1666);
and U2294 (N_2294,N_1774,N_1536);
and U2295 (N_2295,N_1688,N_1550);
nand U2296 (N_2296,N_1670,N_1869);
or U2297 (N_2297,N_1835,N_1895);
or U2298 (N_2298,N_1900,N_1550);
or U2299 (N_2299,N_1672,N_1962);
and U2300 (N_2300,N_1866,N_1779);
and U2301 (N_2301,N_1530,N_1564);
nor U2302 (N_2302,N_1999,N_1801);
nand U2303 (N_2303,N_1828,N_1682);
nand U2304 (N_2304,N_1881,N_1993);
nor U2305 (N_2305,N_1955,N_1815);
or U2306 (N_2306,N_1569,N_1859);
and U2307 (N_2307,N_1714,N_1842);
nor U2308 (N_2308,N_1961,N_1871);
and U2309 (N_2309,N_1789,N_1636);
nand U2310 (N_2310,N_1580,N_1749);
nand U2311 (N_2311,N_1773,N_1789);
or U2312 (N_2312,N_1796,N_1759);
or U2313 (N_2313,N_1551,N_1760);
nor U2314 (N_2314,N_1786,N_1785);
nand U2315 (N_2315,N_1860,N_1935);
and U2316 (N_2316,N_1550,N_1957);
nand U2317 (N_2317,N_1886,N_1868);
nor U2318 (N_2318,N_1787,N_1805);
nand U2319 (N_2319,N_1553,N_1949);
or U2320 (N_2320,N_1708,N_1577);
nor U2321 (N_2321,N_1950,N_1965);
nand U2322 (N_2322,N_1902,N_1623);
or U2323 (N_2323,N_1963,N_1920);
or U2324 (N_2324,N_1794,N_1786);
nor U2325 (N_2325,N_1773,N_1978);
or U2326 (N_2326,N_1789,N_1586);
and U2327 (N_2327,N_1643,N_1575);
nor U2328 (N_2328,N_1605,N_1902);
and U2329 (N_2329,N_1575,N_1813);
or U2330 (N_2330,N_1523,N_1949);
or U2331 (N_2331,N_1932,N_1754);
nand U2332 (N_2332,N_1559,N_1804);
nor U2333 (N_2333,N_1515,N_1769);
and U2334 (N_2334,N_1777,N_1773);
or U2335 (N_2335,N_1701,N_1670);
nand U2336 (N_2336,N_1531,N_1997);
nor U2337 (N_2337,N_1688,N_1559);
or U2338 (N_2338,N_1825,N_1891);
and U2339 (N_2339,N_1954,N_1766);
and U2340 (N_2340,N_1527,N_1822);
and U2341 (N_2341,N_1587,N_1923);
nor U2342 (N_2342,N_1915,N_1896);
nor U2343 (N_2343,N_1865,N_1803);
and U2344 (N_2344,N_1512,N_1788);
or U2345 (N_2345,N_1644,N_1929);
nor U2346 (N_2346,N_1941,N_1522);
nor U2347 (N_2347,N_1794,N_1760);
nor U2348 (N_2348,N_1503,N_1874);
nor U2349 (N_2349,N_1982,N_1887);
nor U2350 (N_2350,N_1601,N_1646);
and U2351 (N_2351,N_1823,N_1592);
or U2352 (N_2352,N_1669,N_1783);
nor U2353 (N_2353,N_1567,N_1808);
nand U2354 (N_2354,N_1989,N_1860);
or U2355 (N_2355,N_1744,N_1604);
nor U2356 (N_2356,N_1905,N_1706);
and U2357 (N_2357,N_1895,N_1723);
and U2358 (N_2358,N_1692,N_1863);
nor U2359 (N_2359,N_1725,N_1939);
nor U2360 (N_2360,N_1656,N_1956);
or U2361 (N_2361,N_1971,N_1740);
and U2362 (N_2362,N_1603,N_1847);
or U2363 (N_2363,N_1768,N_1884);
nand U2364 (N_2364,N_1625,N_1615);
and U2365 (N_2365,N_1686,N_1825);
nand U2366 (N_2366,N_1836,N_1502);
nor U2367 (N_2367,N_1809,N_1910);
or U2368 (N_2368,N_1602,N_1676);
or U2369 (N_2369,N_1747,N_1999);
nor U2370 (N_2370,N_1863,N_1949);
nor U2371 (N_2371,N_1787,N_1756);
or U2372 (N_2372,N_1514,N_1620);
nand U2373 (N_2373,N_1873,N_1844);
nor U2374 (N_2374,N_1544,N_1944);
nor U2375 (N_2375,N_1651,N_1736);
or U2376 (N_2376,N_1740,N_1643);
nor U2377 (N_2377,N_1818,N_1918);
nand U2378 (N_2378,N_1991,N_1691);
and U2379 (N_2379,N_1649,N_1624);
nor U2380 (N_2380,N_1896,N_1935);
or U2381 (N_2381,N_1787,N_1895);
nor U2382 (N_2382,N_1705,N_1890);
nand U2383 (N_2383,N_1908,N_1754);
or U2384 (N_2384,N_1947,N_1647);
or U2385 (N_2385,N_1862,N_1601);
and U2386 (N_2386,N_1736,N_1535);
nand U2387 (N_2387,N_1743,N_1746);
and U2388 (N_2388,N_1808,N_1862);
nand U2389 (N_2389,N_1817,N_1693);
or U2390 (N_2390,N_1907,N_1965);
nand U2391 (N_2391,N_1965,N_1821);
nand U2392 (N_2392,N_1573,N_1863);
or U2393 (N_2393,N_1529,N_1585);
or U2394 (N_2394,N_1997,N_1999);
nand U2395 (N_2395,N_1687,N_1644);
nor U2396 (N_2396,N_1656,N_1978);
nand U2397 (N_2397,N_1565,N_1976);
nor U2398 (N_2398,N_1859,N_1983);
and U2399 (N_2399,N_1676,N_1954);
nor U2400 (N_2400,N_1650,N_1598);
or U2401 (N_2401,N_1719,N_1985);
or U2402 (N_2402,N_1915,N_1912);
and U2403 (N_2403,N_1925,N_1820);
nand U2404 (N_2404,N_1634,N_1811);
and U2405 (N_2405,N_1734,N_1770);
nand U2406 (N_2406,N_1770,N_1527);
or U2407 (N_2407,N_1761,N_1516);
and U2408 (N_2408,N_1813,N_1746);
nor U2409 (N_2409,N_1812,N_1613);
or U2410 (N_2410,N_1557,N_1975);
and U2411 (N_2411,N_1817,N_1742);
or U2412 (N_2412,N_1617,N_1549);
and U2413 (N_2413,N_1582,N_1605);
and U2414 (N_2414,N_1828,N_1535);
and U2415 (N_2415,N_1974,N_1963);
nor U2416 (N_2416,N_1567,N_1837);
and U2417 (N_2417,N_1762,N_1873);
nor U2418 (N_2418,N_1663,N_1892);
nand U2419 (N_2419,N_1995,N_1646);
and U2420 (N_2420,N_1787,N_1552);
or U2421 (N_2421,N_1797,N_1577);
or U2422 (N_2422,N_1753,N_1924);
nor U2423 (N_2423,N_1858,N_1942);
or U2424 (N_2424,N_1707,N_1500);
nand U2425 (N_2425,N_1636,N_1721);
nor U2426 (N_2426,N_1737,N_1806);
and U2427 (N_2427,N_1856,N_1619);
nor U2428 (N_2428,N_1727,N_1594);
nand U2429 (N_2429,N_1749,N_1942);
nand U2430 (N_2430,N_1546,N_1802);
nor U2431 (N_2431,N_1999,N_1637);
nand U2432 (N_2432,N_1928,N_1896);
and U2433 (N_2433,N_1798,N_1898);
nand U2434 (N_2434,N_1875,N_1522);
or U2435 (N_2435,N_1929,N_1893);
and U2436 (N_2436,N_1675,N_1805);
nor U2437 (N_2437,N_1762,N_1601);
nor U2438 (N_2438,N_1542,N_1650);
and U2439 (N_2439,N_1810,N_1858);
nor U2440 (N_2440,N_1561,N_1625);
nand U2441 (N_2441,N_1677,N_1807);
and U2442 (N_2442,N_1615,N_1857);
or U2443 (N_2443,N_1642,N_1867);
and U2444 (N_2444,N_1888,N_1661);
and U2445 (N_2445,N_1995,N_1702);
or U2446 (N_2446,N_1823,N_1928);
and U2447 (N_2447,N_1723,N_1762);
or U2448 (N_2448,N_1598,N_1543);
or U2449 (N_2449,N_1644,N_1871);
or U2450 (N_2450,N_1756,N_1965);
nor U2451 (N_2451,N_1916,N_1820);
and U2452 (N_2452,N_1941,N_1864);
or U2453 (N_2453,N_1783,N_1884);
nor U2454 (N_2454,N_1739,N_1606);
or U2455 (N_2455,N_1623,N_1651);
or U2456 (N_2456,N_1503,N_1963);
nand U2457 (N_2457,N_1827,N_1758);
nor U2458 (N_2458,N_1503,N_1622);
nand U2459 (N_2459,N_1898,N_1549);
and U2460 (N_2460,N_1725,N_1728);
nand U2461 (N_2461,N_1778,N_1604);
or U2462 (N_2462,N_1666,N_1774);
nor U2463 (N_2463,N_1823,N_1584);
or U2464 (N_2464,N_1725,N_1677);
and U2465 (N_2465,N_1743,N_1817);
nor U2466 (N_2466,N_1822,N_1714);
and U2467 (N_2467,N_1819,N_1907);
and U2468 (N_2468,N_1853,N_1790);
or U2469 (N_2469,N_1779,N_1531);
or U2470 (N_2470,N_1911,N_1778);
nand U2471 (N_2471,N_1529,N_1776);
nand U2472 (N_2472,N_1556,N_1940);
or U2473 (N_2473,N_1861,N_1851);
nor U2474 (N_2474,N_1577,N_1897);
nand U2475 (N_2475,N_1518,N_1790);
or U2476 (N_2476,N_1524,N_1663);
nand U2477 (N_2477,N_1609,N_1793);
nor U2478 (N_2478,N_1551,N_1712);
or U2479 (N_2479,N_1597,N_1698);
and U2480 (N_2480,N_1747,N_1992);
nor U2481 (N_2481,N_1989,N_1975);
nand U2482 (N_2482,N_1604,N_1531);
and U2483 (N_2483,N_1797,N_1887);
nand U2484 (N_2484,N_1986,N_1706);
or U2485 (N_2485,N_1522,N_1917);
and U2486 (N_2486,N_1555,N_1751);
nand U2487 (N_2487,N_1573,N_1521);
and U2488 (N_2488,N_1989,N_1955);
nand U2489 (N_2489,N_1737,N_1835);
nand U2490 (N_2490,N_1504,N_1525);
or U2491 (N_2491,N_1821,N_1673);
nand U2492 (N_2492,N_1627,N_1739);
nand U2493 (N_2493,N_1552,N_1992);
nand U2494 (N_2494,N_1675,N_1613);
nand U2495 (N_2495,N_1533,N_1765);
or U2496 (N_2496,N_1558,N_1638);
or U2497 (N_2497,N_1994,N_1516);
nand U2498 (N_2498,N_1660,N_1798);
and U2499 (N_2499,N_1574,N_1721);
nor U2500 (N_2500,N_2002,N_2388);
nor U2501 (N_2501,N_2258,N_2036);
or U2502 (N_2502,N_2354,N_2172);
or U2503 (N_2503,N_2407,N_2262);
nand U2504 (N_2504,N_2241,N_2086);
nand U2505 (N_2505,N_2192,N_2440);
nor U2506 (N_2506,N_2486,N_2113);
and U2507 (N_2507,N_2482,N_2214);
or U2508 (N_2508,N_2017,N_2398);
nand U2509 (N_2509,N_2225,N_2394);
nor U2510 (N_2510,N_2497,N_2463);
nand U2511 (N_2511,N_2223,N_2282);
nand U2512 (N_2512,N_2469,N_2236);
and U2513 (N_2513,N_2293,N_2273);
and U2514 (N_2514,N_2211,N_2392);
or U2515 (N_2515,N_2404,N_2494);
nor U2516 (N_2516,N_2400,N_2382);
nand U2517 (N_2517,N_2053,N_2033);
nand U2518 (N_2518,N_2366,N_2143);
or U2519 (N_2519,N_2155,N_2302);
nor U2520 (N_2520,N_2003,N_2128);
or U2521 (N_2521,N_2168,N_2091);
nand U2522 (N_2522,N_2240,N_2120);
nor U2523 (N_2523,N_2103,N_2314);
nor U2524 (N_2524,N_2378,N_2106);
or U2525 (N_2525,N_2489,N_2044);
nand U2526 (N_2526,N_2342,N_2186);
and U2527 (N_2527,N_2275,N_2030);
or U2528 (N_2528,N_2268,N_2357);
or U2529 (N_2529,N_2177,N_2391);
nor U2530 (N_2530,N_2100,N_2287);
or U2531 (N_2531,N_2080,N_2251);
and U2532 (N_2532,N_2054,N_2064);
nor U2533 (N_2533,N_2333,N_2456);
nor U2534 (N_2534,N_2291,N_2071);
nor U2535 (N_2535,N_2141,N_2216);
nor U2536 (N_2536,N_2343,N_2008);
nor U2537 (N_2537,N_2427,N_2462);
or U2538 (N_2538,N_2235,N_2477);
and U2539 (N_2539,N_2323,N_2083);
or U2540 (N_2540,N_2358,N_2485);
nand U2541 (N_2541,N_2047,N_2110);
nand U2542 (N_2542,N_2220,N_2156);
or U2543 (N_2543,N_2340,N_2416);
and U2544 (N_2544,N_2350,N_2271);
nor U2545 (N_2545,N_2090,N_2239);
nor U2546 (N_2546,N_2248,N_2237);
or U2547 (N_2547,N_2222,N_2279);
or U2548 (N_2548,N_2260,N_2134);
nand U2549 (N_2549,N_2459,N_2413);
and U2550 (N_2550,N_2067,N_2329);
nor U2551 (N_2551,N_2495,N_2115);
or U2552 (N_2552,N_2180,N_2073);
and U2553 (N_2553,N_2283,N_2153);
nor U2554 (N_2554,N_2377,N_2432);
nand U2555 (N_2555,N_2174,N_2041);
and U2556 (N_2556,N_2060,N_2396);
and U2557 (N_2557,N_2311,N_2453);
and U2558 (N_2558,N_2347,N_2245);
nand U2559 (N_2559,N_2124,N_2082);
and U2560 (N_2560,N_2049,N_2146);
nand U2561 (N_2561,N_2447,N_2270);
and U2562 (N_2562,N_2484,N_2165);
and U2563 (N_2563,N_2249,N_2009);
nor U2564 (N_2564,N_2107,N_2012);
nand U2565 (N_2565,N_2039,N_2175);
or U2566 (N_2566,N_2133,N_2405);
and U2567 (N_2567,N_2170,N_2452);
or U2568 (N_2568,N_2018,N_2108);
and U2569 (N_2569,N_2118,N_2034);
or U2570 (N_2570,N_2490,N_2429);
or U2571 (N_2571,N_2423,N_2042);
nor U2572 (N_2572,N_2367,N_2428);
nor U2573 (N_2573,N_2199,N_2478);
and U2574 (N_2574,N_2243,N_2126);
and U2575 (N_2575,N_2465,N_2070);
nand U2576 (N_2576,N_2238,N_2431);
nand U2577 (N_2577,N_2252,N_2492);
or U2578 (N_2578,N_2443,N_2253);
nand U2579 (N_2579,N_2219,N_2176);
nor U2580 (N_2580,N_2132,N_2406);
nand U2581 (N_2581,N_2137,N_2196);
or U2582 (N_2582,N_2266,N_2163);
nand U2583 (N_2583,N_2210,N_2050);
nand U2584 (N_2584,N_2322,N_2450);
and U2585 (N_2585,N_2373,N_2230);
nand U2586 (N_2586,N_2286,N_2289);
and U2587 (N_2587,N_2109,N_2037);
nand U2588 (N_2588,N_2043,N_2010);
nand U2589 (N_2589,N_2409,N_2221);
nand U2590 (N_2590,N_2346,N_2401);
nand U2591 (N_2591,N_2085,N_2470);
nor U2592 (N_2592,N_2076,N_2062);
nand U2593 (N_2593,N_2442,N_2435);
and U2594 (N_2594,N_2295,N_2006);
or U2595 (N_2595,N_2095,N_2144);
and U2596 (N_2596,N_2345,N_2375);
xnor U2597 (N_2597,N_2261,N_2181);
and U2598 (N_2598,N_2077,N_2119);
nor U2599 (N_2599,N_2046,N_2310);
nor U2600 (N_2600,N_2499,N_2166);
xnor U2601 (N_2601,N_2298,N_2228);
nand U2602 (N_2602,N_2102,N_2264);
and U2603 (N_2603,N_2209,N_2142);
and U2604 (N_2604,N_2386,N_2152);
nand U2605 (N_2605,N_2496,N_2403);
nand U2606 (N_2606,N_2419,N_2059);
nand U2607 (N_2607,N_2438,N_2048);
and U2608 (N_2608,N_2320,N_2184);
and U2609 (N_2609,N_2290,N_2171);
and U2610 (N_2610,N_2362,N_2341);
nand U2611 (N_2611,N_2472,N_2325);
and U2612 (N_2612,N_2361,N_2079);
and U2613 (N_2613,N_2455,N_2246);
nand U2614 (N_2614,N_2127,N_2300);
nand U2615 (N_2615,N_2149,N_2173);
nor U2616 (N_2616,N_2430,N_2093);
nand U2617 (N_2617,N_2097,N_2198);
or U2618 (N_2618,N_2330,N_2277);
nor U2619 (N_2619,N_2092,N_2384);
nand U2620 (N_2620,N_2069,N_2063);
nand U2621 (N_2621,N_2372,N_2191);
or U2622 (N_2622,N_2061,N_2234);
nand U2623 (N_2623,N_2299,N_2139);
and U2624 (N_2624,N_2111,N_2393);
nor U2625 (N_2625,N_2027,N_2474);
nor U2626 (N_2626,N_2158,N_2437);
nand U2627 (N_2627,N_2130,N_2415);
nand U2628 (N_2628,N_2159,N_2278);
nor U2629 (N_2629,N_2331,N_2318);
and U2630 (N_2630,N_2464,N_2259);
or U2631 (N_2631,N_2308,N_2206);
or U2632 (N_2632,N_2138,N_2454);
and U2633 (N_2633,N_2162,N_2292);
or U2634 (N_2634,N_2369,N_2204);
nor U2635 (N_2635,N_2466,N_2116);
and U2636 (N_2636,N_2125,N_2122);
nor U2637 (N_2637,N_2229,N_2352);
nand U2638 (N_2638,N_2312,N_2444);
nand U2639 (N_2639,N_2029,N_2169);
and U2640 (N_2640,N_2038,N_2231);
nor U2641 (N_2641,N_2324,N_2381);
and U2642 (N_2642,N_2194,N_2136);
nand U2643 (N_2643,N_2334,N_2131);
and U2644 (N_2644,N_2021,N_2267);
and U2645 (N_2645,N_2099,N_2483);
and U2646 (N_2646,N_2359,N_2226);
nand U2647 (N_2647,N_2178,N_2274);
nor U2648 (N_2648,N_2232,N_2190);
and U2649 (N_2649,N_2212,N_2439);
nand U2650 (N_2650,N_2461,N_2321);
and U2651 (N_2651,N_2072,N_2183);
nand U2652 (N_2652,N_2436,N_2179);
nor U2653 (N_2653,N_2348,N_2215);
nand U2654 (N_2654,N_2326,N_2397);
and U2655 (N_2655,N_2151,N_2066);
nor U2656 (N_2656,N_2385,N_2414);
nand U2657 (N_2657,N_2389,N_2255);
or U2658 (N_2658,N_2319,N_2150);
nor U2659 (N_2659,N_2123,N_2356);
or U2660 (N_2660,N_2145,N_2412);
nor U2661 (N_2661,N_2218,N_2250);
nand U2662 (N_2662,N_2434,N_2104);
and U2663 (N_2663,N_2317,N_2088);
nor U2664 (N_2664,N_2032,N_2446);
or U2665 (N_2665,N_2313,N_2448);
and U2666 (N_2666,N_2285,N_2476);
xnor U2667 (N_2667,N_2098,N_2185);
nand U2668 (N_2668,N_2084,N_2307);
and U2669 (N_2669,N_2488,N_2004);
and U2670 (N_2670,N_2201,N_2498);
nor U2671 (N_2671,N_2468,N_2114);
and U2672 (N_2672,N_2272,N_2189);
and U2673 (N_2673,N_2424,N_2254);
or U2674 (N_2674,N_2402,N_2303);
nand U2675 (N_2675,N_2227,N_2420);
or U2676 (N_2676,N_2217,N_2441);
or U2677 (N_2677,N_2154,N_2418);
nand U2678 (N_2678,N_2451,N_2460);
nor U2679 (N_2679,N_2368,N_2387);
nor U2680 (N_2680,N_2473,N_2493);
and U2681 (N_2681,N_2074,N_2193);
and U2682 (N_2682,N_2294,N_2425);
nor U2683 (N_2683,N_2339,N_2031);
or U2684 (N_2684,N_2376,N_2297);
nand U2685 (N_2685,N_2395,N_2265);
and U2686 (N_2686,N_2207,N_2015);
and U2687 (N_2687,N_2316,N_2058);
nand U2688 (N_2688,N_2257,N_2305);
and U2689 (N_2689,N_2337,N_2148);
nor U2690 (N_2690,N_2365,N_2019);
nand U2691 (N_2691,N_2491,N_2349);
and U2692 (N_2692,N_2089,N_2160);
nor U2693 (N_2693,N_2399,N_2057);
and U2694 (N_2694,N_2028,N_2315);
and U2695 (N_2695,N_2247,N_2445);
nand U2696 (N_2696,N_2360,N_2203);
xnor U2697 (N_2697,N_2481,N_2263);
nand U2698 (N_2698,N_2288,N_2129);
or U2699 (N_2699,N_2480,N_2202);
nand U2700 (N_2700,N_2055,N_2068);
nor U2701 (N_2701,N_2075,N_2379);
nor U2702 (N_2702,N_2022,N_2001);
nand U2703 (N_2703,N_2433,N_2351);
or U2704 (N_2704,N_2304,N_2421);
nor U2705 (N_2705,N_2167,N_2363);
or U2706 (N_2706,N_2101,N_2205);
or U2707 (N_2707,N_2087,N_2096);
and U2708 (N_2708,N_2200,N_2182);
nand U2709 (N_2709,N_2025,N_2187);
nand U2710 (N_2710,N_2188,N_2479);
nor U2711 (N_2711,N_2208,N_2016);
nand U2712 (N_2712,N_2051,N_2244);
nand U2713 (N_2713,N_2197,N_2422);
nor U2714 (N_2714,N_2335,N_2371);
and U2715 (N_2715,N_2242,N_2309);
nor U2716 (N_2716,N_2471,N_2475);
nor U2717 (N_2717,N_2327,N_2353);
nor U2718 (N_2718,N_2052,N_2449);
nand U2719 (N_2719,N_2284,N_2078);
and U2720 (N_2720,N_2157,N_2195);
nand U2721 (N_2721,N_2344,N_2011);
nand U2722 (N_2722,N_2338,N_2213);
nand U2723 (N_2723,N_2233,N_2105);
or U2724 (N_2724,N_2000,N_2081);
nor U2725 (N_2725,N_2380,N_2020);
nor U2726 (N_2726,N_2121,N_2013);
or U2727 (N_2727,N_2040,N_2417);
or U2728 (N_2728,N_2336,N_2411);
and U2729 (N_2729,N_2094,N_2370);
and U2730 (N_2730,N_2332,N_2390);
nor U2731 (N_2731,N_2487,N_2164);
nand U2732 (N_2732,N_2457,N_2296);
and U2733 (N_2733,N_2135,N_2005);
nand U2734 (N_2734,N_2147,N_2467);
nor U2735 (N_2735,N_2140,N_2117);
nor U2736 (N_2736,N_2023,N_2007);
nor U2737 (N_2737,N_2269,N_2161);
or U2738 (N_2738,N_2301,N_2014);
xnor U2739 (N_2739,N_2374,N_2256);
nor U2740 (N_2740,N_2026,N_2276);
nor U2741 (N_2741,N_2045,N_2056);
and U2742 (N_2742,N_2065,N_2408);
nand U2743 (N_2743,N_2024,N_2280);
nor U2744 (N_2744,N_2112,N_2328);
and U2745 (N_2745,N_2281,N_2306);
or U2746 (N_2746,N_2364,N_2383);
or U2747 (N_2747,N_2426,N_2458);
or U2748 (N_2748,N_2035,N_2410);
nor U2749 (N_2749,N_2224,N_2355);
nor U2750 (N_2750,N_2447,N_2214);
nor U2751 (N_2751,N_2149,N_2472);
nand U2752 (N_2752,N_2070,N_2448);
nand U2753 (N_2753,N_2487,N_2281);
or U2754 (N_2754,N_2099,N_2479);
or U2755 (N_2755,N_2189,N_2016);
or U2756 (N_2756,N_2114,N_2165);
or U2757 (N_2757,N_2450,N_2396);
and U2758 (N_2758,N_2248,N_2342);
or U2759 (N_2759,N_2497,N_2131);
nand U2760 (N_2760,N_2107,N_2182);
nand U2761 (N_2761,N_2415,N_2446);
and U2762 (N_2762,N_2282,N_2458);
nand U2763 (N_2763,N_2482,N_2405);
xor U2764 (N_2764,N_2206,N_2467);
nand U2765 (N_2765,N_2368,N_2494);
nand U2766 (N_2766,N_2484,N_2424);
and U2767 (N_2767,N_2030,N_2318);
and U2768 (N_2768,N_2374,N_2244);
and U2769 (N_2769,N_2389,N_2452);
nand U2770 (N_2770,N_2033,N_2263);
nor U2771 (N_2771,N_2236,N_2424);
and U2772 (N_2772,N_2273,N_2353);
and U2773 (N_2773,N_2182,N_2428);
nor U2774 (N_2774,N_2132,N_2368);
or U2775 (N_2775,N_2288,N_2094);
nor U2776 (N_2776,N_2144,N_2340);
nand U2777 (N_2777,N_2181,N_2196);
or U2778 (N_2778,N_2221,N_2487);
or U2779 (N_2779,N_2127,N_2464);
nand U2780 (N_2780,N_2133,N_2257);
nor U2781 (N_2781,N_2178,N_2267);
or U2782 (N_2782,N_2094,N_2218);
nor U2783 (N_2783,N_2179,N_2210);
xnor U2784 (N_2784,N_2421,N_2259);
nor U2785 (N_2785,N_2344,N_2465);
nor U2786 (N_2786,N_2196,N_2073);
and U2787 (N_2787,N_2169,N_2421);
and U2788 (N_2788,N_2087,N_2161);
nand U2789 (N_2789,N_2412,N_2105);
nand U2790 (N_2790,N_2134,N_2412);
or U2791 (N_2791,N_2117,N_2131);
and U2792 (N_2792,N_2147,N_2087);
and U2793 (N_2793,N_2438,N_2244);
nor U2794 (N_2794,N_2212,N_2028);
nor U2795 (N_2795,N_2320,N_2272);
nand U2796 (N_2796,N_2305,N_2195);
nor U2797 (N_2797,N_2348,N_2055);
and U2798 (N_2798,N_2005,N_2230);
nor U2799 (N_2799,N_2469,N_2033);
xor U2800 (N_2800,N_2385,N_2425);
nand U2801 (N_2801,N_2296,N_2468);
and U2802 (N_2802,N_2100,N_2064);
nand U2803 (N_2803,N_2305,N_2039);
or U2804 (N_2804,N_2299,N_2235);
and U2805 (N_2805,N_2087,N_2083);
and U2806 (N_2806,N_2045,N_2327);
nor U2807 (N_2807,N_2464,N_2185);
nand U2808 (N_2808,N_2189,N_2366);
nor U2809 (N_2809,N_2344,N_2278);
nand U2810 (N_2810,N_2335,N_2492);
or U2811 (N_2811,N_2008,N_2328);
or U2812 (N_2812,N_2078,N_2467);
nand U2813 (N_2813,N_2442,N_2144);
nor U2814 (N_2814,N_2380,N_2249);
nor U2815 (N_2815,N_2163,N_2142);
or U2816 (N_2816,N_2310,N_2464);
and U2817 (N_2817,N_2075,N_2034);
nand U2818 (N_2818,N_2225,N_2177);
nand U2819 (N_2819,N_2310,N_2001);
nand U2820 (N_2820,N_2471,N_2079);
or U2821 (N_2821,N_2411,N_2309);
or U2822 (N_2822,N_2043,N_2419);
nand U2823 (N_2823,N_2243,N_2172);
or U2824 (N_2824,N_2135,N_2259);
and U2825 (N_2825,N_2169,N_2404);
or U2826 (N_2826,N_2117,N_2236);
or U2827 (N_2827,N_2494,N_2471);
nand U2828 (N_2828,N_2247,N_2292);
nand U2829 (N_2829,N_2097,N_2102);
and U2830 (N_2830,N_2153,N_2469);
or U2831 (N_2831,N_2143,N_2417);
and U2832 (N_2832,N_2098,N_2244);
nor U2833 (N_2833,N_2254,N_2468);
and U2834 (N_2834,N_2456,N_2165);
and U2835 (N_2835,N_2082,N_2350);
nor U2836 (N_2836,N_2267,N_2153);
and U2837 (N_2837,N_2127,N_2216);
or U2838 (N_2838,N_2264,N_2236);
nor U2839 (N_2839,N_2384,N_2136);
nor U2840 (N_2840,N_2112,N_2347);
nor U2841 (N_2841,N_2143,N_2060);
nor U2842 (N_2842,N_2197,N_2236);
nor U2843 (N_2843,N_2075,N_2174);
nand U2844 (N_2844,N_2189,N_2345);
or U2845 (N_2845,N_2439,N_2358);
nor U2846 (N_2846,N_2105,N_2446);
nand U2847 (N_2847,N_2197,N_2344);
nand U2848 (N_2848,N_2156,N_2303);
nor U2849 (N_2849,N_2032,N_2010);
nor U2850 (N_2850,N_2092,N_2497);
and U2851 (N_2851,N_2058,N_2237);
nand U2852 (N_2852,N_2029,N_2390);
nand U2853 (N_2853,N_2324,N_2436);
nor U2854 (N_2854,N_2212,N_2260);
nand U2855 (N_2855,N_2277,N_2423);
nor U2856 (N_2856,N_2274,N_2217);
nor U2857 (N_2857,N_2489,N_2412);
and U2858 (N_2858,N_2231,N_2329);
and U2859 (N_2859,N_2277,N_2469);
nor U2860 (N_2860,N_2126,N_2095);
or U2861 (N_2861,N_2194,N_2026);
nand U2862 (N_2862,N_2079,N_2008);
or U2863 (N_2863,N_2499,N_2490);
nand U2864 (N_2864,N_2330,N_2066);
nand U2865 (N_2865,N_2440,N_2090);
or U2866 (N_2866,N_2465,N_2059);
nand U2867 (N_2867,N_2027,N_2239);
and U2868 (N_2868,N_2338,N_2499);
nand U2869 (N_2869,N_2261,N_2380);
and U2870 (N_2870,N_2091,N_2099);
nand U2871 (N_2871,N_2052,N_2443);
nand U2872 (N_2872,N_2230,N_2380);
and U2873 (N_2873,N_2178,N_2151);
nor U2874 (N_2874,N_2107,N_2055);
or U2875 (N_2875,N_2416,N_2376);
nor U2876 (N_2876,N_2357,N_2129);
nand U2877 (N_2877,N_2310,N_2334);
nand U2878 (N_2878,N_2141,N_2093);
nand U2879 (N_2879,N_2446,N_2017);
or U2880 (N_2880,N_2001,N_2134);
nor U2881 (N_2881,N_2340,N_2472);
nand U2882 (N_2882,N_2299,N_2428);
or U2883 (N_2883,N_2150,N_2081);
and U2884 (N_2884,N_2484,N_2062);
nor U2885 (N_2885,N_2304,N_2235);
nand U2886 (N_2886,N_2141,N_2383);
and U2887 (N_2887,N_2179,N_2127);
or U2888 (N_2888,N_2083,N_2160);
nand U2889 (N_2889,N_2383,N_2156);
nor U2890 (N_2890,N_2336,N_2021);
nand U2891 (N_2891,N_2478,N_2497);
or U2892 (N_2892,N_2025,N_2446);
nor U2893 (N_2893,N_2081,N_2178);
nor U2894 (N_2894,N_2358,N_2368);
nand U2895 (N_2895,N_2481,N_2300);
or U2896 (N_2896,N_2182,N_2404);
nand U2897 (N_2897,N_2132,N_2403);
nand U2898 (N_2898,N_2422,N_2125);
and U2899 (N_2899,N_2261,N_2455);
nor U2900 (N_2900,N_2358,N_2429);
or U2901 (N_2901,N_2491,N_2119);
or U2902 (N_2902,N_2157,N_2248);
nor U2903 (N_2903,N_2048,N_2234);
and U2904 (N_2904,N_2349,N_2171);
nand U2905 (N_2905,N_2113,N_2105);
nor U2906 (N_2906,N_2248,N_2194);
or U2907 (N_2907,N_2379,N_2047);
or U2908 (N_2908,N_2314,N_2488);
nand U2909 (N_2909,N_2196,N_2222);
or U2910 (N_2910,N_2278,N_2092);
nand U2911 (N_2911,N_2306,N_2061);
or U2912 (N_2912,N_2030,N_2233);
nor U2913 (N_2913,N_2367,N_2291);
and U2914 (N_2914,N_2191,N_2236);
nor U2915 (N_2915,N_2015,N_2004);
nor U2916 (N_2916,N_2327,N_2185);
nand U2917 (N_2917,N_2243,N_2230);
nor U2918 (N_2918,N_2497,N_2378);
nand U2919 (N_2919,N_2367,N_2385);
nand U2920 (N_2920,N_2321,N_2368);
nand U2921 (N_2921,N_2037,N_2023);
or U2922 (N_2922,N_2357,N_2437);
or U2923 (N_2923,N_2122,N_2481);
nand U2924 (N_2924,N_2093,N_2301);
nor U2925 (N_2925,N_2360,N_2442);
nor U2926 (N_2926,N_2141,N_2392);
and U2927 (N_2927,N_2406,N_2257);
and U2928 (N_2928,N_2070,N_2202);
and U2929 (N_2929,N_2007,N_2380);
or U2930 (N_2930,N_2161,N_2150);
nor U2931 (N_2931,N_2132,N_2486);
or U2932 (N_2932,N_2275,N_2096);
or U2933 (N_2933,N_2377,N_2357);
nand U2934 (N_2934,N_2264,N_2477);
or U2935 (N_2935,N_2220,N_2408);
or U2936 (N_2936,N_2291,N_2265);
nor U2937 (N_2937,N_2295,N_2351);
nand U2938 (N_2938,N_2483,N_2346);
and U2939 (N_2939,N_2215,N_2019);
nand U2940 (N_2940,N_2434,N_2161);
nor U2941 (N_2941,N_2073,N_2145);
nand U2942 (N_2942,N_2340,N_2296);
and U2943 (N_2943,N_2371,N_2441);
nor U2944 (N_2944,N_2349,N_2315);
nand U2945 (N_2945,N_2427,N_2255);
and U2946 (N_2946,N_2069,N_2460);
nor U2947 (N_2947,N_2198,N_2025);
or U2948 (N_2948,N_2052,N_2253);
nor U2949 (N_2949,N_2062,N_2217);
and U2950 (N_2950,N_2028,N_2156);
or U2951 (N_2951,N_2479,N_2394);
or U2952 (N_2952,N_2137,N_2492);
or U2953 (N_2953,N_2143,N_2117);
nor U2954 (N_2954,N_2189,N_2346);
or U2955 (N_2955,N_2188,N_2168);
nand U2956 (N_2956,N_2107,N_2111);
nor U2957 (N_2957,N_2236,N_2432);
nor U2958 (N_2958,N_2176,N_2387);
or U2959 (N_2959,N_2327,N_2031);
nor U2960 (N_2960,N_2395,N_2131);
or U2961 (N_2961,N_2277,N_2054);
and U2962 (N_2962,N_2368,N_2468);
nand U2963 (N_2963,N_2056,N_2488);
nand U2964 (N_2964,N_2041,N_2001);
or U2965 (N_2965,N_2322,N_2221);
or U2966 (N_2966,N_2232,N_2032);
nand U2967 (N_2967,N_2339,N_2226);
and U2968 (N_2968,N_2400,N_2168);
nand U2969 (N_2969,N_2462,N_2279);
nor U2970 (N_2970,N_2365,N_2406);
and U2971 (N_2971,N_2062,N_2052);
or U2972 (N_2972,N_2489,N_2369);
nor U2973 (N_2973,N_2075,N_2268);
nand U2974 (N_2974,N_2321,N_2418);
and U2975 (N_2975,N_2033,N_2088);
xnor U2976 (N_2976,N_2496,N_2359);
nor U2977 (N_2977,N_2287,N_2482);
or U2978 (N_2978,N_2056,N_2264);
nor U2979 (N_2979,N_2499,N_2070);
nand U2980 (N_2980,N_2106,N_2101);
nand U2981 (N_2981,N_2210,N_2101);
nand U2982 (N_2982,N_2004,N_2468);
nor U2983 (N_2983,N_2249,N_2467);
and U2984 (N_2984,N_2115,N_2271);
nor U2985 (N_2985,N_2318,N_2323);
or U2986 (N_2986,N_2345,N_2321);
nor U2987 (N_2987,N_2203,N_2192);
nand U2988 (N_2988,N_2336,N_2236);
nor U2989 (N_2989,N_2089,N_2437);
nand U2990 (N_2990,N_2466,N_2075);
nor U2991 (N_2991,N_2075,N_2318);
or U2992 (N_2992,N_2378,N_2252);
nand U2993 (N_2993,N_2318,N_2145);
or U2994 (N_2994,N_2103,N_2207);
and U2995 (N_2995,N_2227,N_2333);
xnor U2996 (N_2996,N_2085,N_2417);
nand U2997 (N_2997,N_2140,N_2158);
nor U2998 (N_2998,N_2466,N_2048);
nand U2999 (N_2999,N_2208,N_2220);
nor UO_0 (O_0,N_2961,N_2832);
or UO_1 (O_1,N_2552,N_2850);
nor UO_2 (O_2,N_2935,N_2980);
nand UO_3 (O_3,N_2659,N_2804);
or UO_4 (O_4,N_2638,N_2545);
nor UO_5 (O_5,N_2815,N_2555);
and UO_6 (O_6,N_2701,N_2929);
nor UO_7 (O_7,N_2535,N_2778);
nor UO_8 (O_8,N_2729,N_2588);
and UO_9 (O_9,N_2840,N_2847);
nand UO_10 (O_10,N_2707,N_2689);
nor UO_11 (O_11,N_2661,N_2616);
nor UO_12 (O_12,N_2993,N_2735);
nand UO_13 (O_13,N_2767,N_2795);
and UO_14 (O_14,N_2514,N_2699);
or UO_15 (O_15,N_2538,N_2543);
nor UO_16 (O_16,N_2972,N_2754);
nor UO_17 (O_17,N_2906,N_2569);
nand UO_18 (O_18,N_2768,N_2720);
or UO_19 (O_19,N_2919,N_2668);
nor UO_20 (O_20,N_2824,N_2835);
nor UO_21 (O_21,N_2724,N_2725);
and UO_22 (O_22,N_2976,N_2985);
nand UO_23 (O_23,N_2737,N_2758);
nand UO_24 (O_24,N_2665,N_2992);
nor UO_25 (O_25,N_2837,N_2708);
nor UO_26 (O_26,N_2944,N_2710);
nand UO_27 (O_27,N_2994,N_2879);
and UO_28 (O_28,N_2849,N_2641);
or UO_29 (O_29,N_2524,N_2618);
or UO_30 (O_30,N_2749,N_2878);
xor UO_31 (O_31,N_2893,N_2677);
or UO_32 (O_32,N_2572,N_2669);
and UO_33 (O_33,N_2612,N_2958);
and UO_34 (O_34,N_2602,N_2846);
nand UO_35 (O_35,N_2521,N_2627);
or UO_36 (O_36,N_2955,N_2968);
nor UO_37 (O_37,N_2712,N_2862);
nor UO_38 (O_38,N_2554,N_2848);
and UO_39 (O_39,N_2809,N_2694);
and UO_40 (O_40,N_2772,N_2649);
or UO_41 (O_41,N_2765,N_2932);
or UO_42 (O_42,N_2875,N_2648);
nor UO_43 (O_43,N_2800,N_2637);
nor UO_44 (O_44,N_2760,N_2500);
and UO_45 (O_45,N_2723,N_2933);
or UO_46 (O_46,N_2518,N_2506);
nand UO_47 (O_47,N_2951,N_2954);
nand UO_48 (O_48,N_2923,N_2881);
and UO_49 (O_49,N_2709,N_2746);
or UO_50 (O_50,N_2797,N_2647);
nand UO_51 (O_51,N_2692,N_2744);
and UO_52 (O_52,N_2722,N_2567);
and UO_53 (O_53,N_2704,N_2609);
nand UO_54 (O_54,N_2696,N_2546);
xor UO_55 (O_55,N_2788,N_2947);
and UO_56 (O_56,N_2585,N_2789);
nand UO_57 (O_57,N_2711,N_2949);
or UO_58 (O_58,N_2752,N_2913);
nand UO_59 (O_59,N_2808,N_2801);
nand UO_60 (O_60,N_2779,N_2888);
or UO_61 (O_61,N_2916,N_2628);
nand UO_62 (O_62,N_2613,N_2584);
nand UO_63 (O_63,N_2805,N_2956);
or UO_64 (O_64,N_2587,N_2902);
nor UO_65 (O_65,N_2676,N_2642);
nand UO_66 (O_66,N_2666,N_2945);
nor UO_67 (O_67,N_2792,N_2682);
nor UO_68 (O_68,N_2905,N_2730);
and UO_69 (O_69,N_2855,N_2528);
and UO_70 (O_70,N_2581,N_2589);
nor UO_71 (O_71,N_2926,N_2684);
and UO_72 (O_72,N_2565,N_2776);
or UO_73 (O_73,N_2610,N_2925);
and UO_74 (O_74,N_2716,N_2774);
or UO_75 (O_75,N_2871,N_2734);
and UO_76 (O_76,N_2997,N_2928);
nor UO_77 (O_77,N_2784,N_2970);
and UO_78 (O_78,N_2551,N_2502);
nand UO_79 (O_79,N_2510,N_2915);
and UO_80 (O_80,N_2576,N_2889);
or UO_81 (O_81,N_2903,N_2987);
or UO_82 (O_82,N_2831,N_2736);
or UO_83 (O_83,N_2516,N_2683);
and UO_84 (O_84,N_2963,N_2596);
or UO_85 (O_85,N_2592,N_2799);
or UO_86 (O_86,N_2673,N_2501);
and UO_87 (O_87,N_2728,N_2690);
and UO_88 (O_88,N_2941,N_2939);
nand UO_89 (O_89,N_2814,N_2549);
and UO_90 (O_90,N_2988,N_2914);
and UO_91 (O_91,N_2670,N_2912);
nor UO_92 (O_92,N_2845,N_2973);
nand UO_93 (O_93,N_2548,N_2738);
nand UO_94 (O_94,N_2917,N_2898);
nor UO_95 (O_95,N_2859,N_2547);
and UO_96 (O_96,N_2953,N_2529);
and UO_97 (O_97,N_2922,N_2745);
nor UO_98 (O_98,N_2751,N_2851);
and UO_99 (O_99,N_2530,N_2887);
nand UO_100 (O_100,N_2531,N_2975);
nor UO_101 (O_101,N_2757,N_2620);
or UO_102 (O_102,N_2748,N_2523);
nand UO_103 (O_103,N_2532,N_2693);
or UO_104 (O_104,N_2911,N_2622);
and UO_105 (O_105,N_2743,N_2894);
or UO_106 (O_106,N_2901,N_2816);
or UO_107 (O_107,N_2731,N_2654);
nand UO_108 (O_108,N_2962,N_2562);
nand UO_109 (O_109,N_2841,N_2515);
nand UO_110 (O_110,N_2632,N_2866);
or UO_111 (O_111,N_2623,N_2899);
and UO_112 (O_112,N_2578,N_2786);
nor UO_113 (O_113,N_2787,N_2702);
nor UO_114 (O_114,N_2839,N_2721);
or UO_115 (O_115,N_2877,N_2686);
nand UO_116 (O_116,N_2527,N_2582);
and UO_117 (O_117,N_2507,N_2864);
nor UO_118 (O_118,N_2780,N_2769);
nand UO_119 (O_119,N_2553,N_2820);
nand UO_120 (O_120,N_2759,N_2568);
nand UO_121 (O_121,N_2909,N_2950);
and UO_122 (O_122,N_2560,N_2785);
or UO_123 (O_123,N_2873,N_2571);
nand UO_124 (O_124,N_2503,N_2557);
or UO_125 (O_125,N_2936,N_2794);
or UO_126 (O_126,N_2777,N_2671);
nor UO_127 (O_127,N_2965,N_2519);
nand UO_128 (O_128,N_2559,N_2969);
nor UO_129 (O_129,N_2634,N_2825);
nor UO_130 (O_130,N_2924,N_2977);
nor UO_131 (O_131,N_2667,N_2747);
or UO_132 (O_132,N_2896,N_2534);
nand UO_133 (O_133,N_2796,N_2583);
and UO_134 (O_134,N_2750,N_2678);
nor UO_135 (O_135,N_2595,N_2586);
or UO_136 (O_136,N_2826,N_2823);
or UO_137 (O_137,N_2967,N_2940);
nand UO_138 (O_138,N_2869,N_2617);
nor UO_139 (O_139,N_2960,N_2505);
nand UO_140 (O_140,N_2842,N_2513);
xnor UO_141 (O_141,N_2775,N_2580);
nand UO_142 (O_142,N_2998,N_2883);
and UO_143 (O_143,N_2830,N_2811);
or UO_144 (O_144,N_2921,N_2727);
nor UO_145 (O_145,N_2593,N_2604);
or UO_146 (O_146,N_2964,N_2761);
or UO_147 (O_147,N_2890,N_2904);
and UO_148 (O_148,N_2742,N_2542);
xnor UO_149 (O_149,N_2856,N_2626);
xor UO_150 (O_150,N_2817,N_2611);
and UO_151 (O_151,N_2983,N_2573);
and UO_152 (O_152,N_2597,N_2558);
and UO_153 (O_153,N_2766,N_2865);
xor UO_154 (O_154,N_2959,N_2833);
nor UO_155 (O_155,N_2655,N_2601);
nor UO_156 (O_156,N_2931,N_2782);
and UO_157 (O_157,N_2999,N_2783);
or UO_158 (O_158,N_2544,N_2605);
or UO_159 (O_159,N_2679,N_2629);
nor UO_160 (O_160,N_2537,N_2615);
nand UO_161 (O_161,N_2645,N_2812);
nand UO_162 (O_162,N_2658,N_2539);
nand UO_163 (O_163,N_2630,N_2844);
and UO_164 (O_164,N_2753,N_2918);
nor UO_165 (O_165,N_2876,N_2600);
nand UO_166 (O_166,N_2946,N_2662);
nand UO_167 (O_167,N_2719,N_2706);
or UO_168 (O_168,N_2533,N_2663);
nor UO_169 (O_169,N_2900,N_2884);
or UO_170 (O_170,N_2536,N_2764);
nor UO_171 (O_171,N_2691,N_2700);
and UO_172 (O_172,N_2687,N_2836);
nor UO_173 (O_173,N_2781,N_2908);
and UO_174 (O_174,N_2807,N_2829);
and UO_175 (O_175,N_2813,N_2504);
nand UO_176 (O_176,N_2803,N_2644);
or UO_177 (O_177,N_2574,N_2920);
nor UO_178 (O_178,N_2798,N_2793);
or UO_179 (O_179,N_2741,N_2874);
or UO_180 (O_180,N_2755,N_2631);
nand UO_181 (O_181,N_2656,N_2520);
nor UO_182 (O_182,N_2681,N_2575);
nor UO_183 (O_183,N_2640,N_2633);
and UO_184 (O_184,N_2643,N_2621);
nor UO_185 (O_185,N_2927,N_2541);
nand UO_186 (O_186,N_2857,N_2982);
nand UO_187 (O_187,N_2508,N_2948);
and UO_188 (O_188,N_2646,N_2625);
and UO_189 (O_189,N_2608,N_2624);
and UO_190 (O_190,N_2819,N_2550);
nand UO_191 (O_191,N_2981,N_2897);
and UO_192 (O_192,N_2938,N_2930);
and UO_193 (O_193,N_2861,N_2674);
or UO_194 (O_194,N_2957,N_2880);
or UO_195 (O_195,N_2995,N_2853);
xor UO_196 (O_196,N_2996,N_2740);
nor UO_197 (O_197,N_2762,N_2717);
and UO_198 (O_198,N_2713,N_2863);
nor UO_199 (O_199,N_2942,N_2763);
nor UO_200 (O_200,N_2838,N_2697);
nand UO_201 (O_201,N_2886,N_2885);
nand UO_202 (O_202,N_2525,N_2512);
nor UO_203 (O_203,N_2810,N_2652);
or UO_204 (O_204,N_2986,N_2979);
or UO_205 (O_205,N_2688,N_2952);
nor UO_206 (O_206,N_2821,N_2564);
and UO_207 (O_207,N_2556,N_2526);
nand UO_208 (O_208,N_2974,N_2715);
and UO_209 (O_209,N_2718,N_2858);
or UO_210 (O_210,N_2966,N_2790);
nor UO_211 (O_211,N_2714,N_2991);
or UO_212 (O_212,N_2603,N_2685);
nand UO_213 (O_213,N_2854,N_2990);
or UO_214 (O_214,N_2680,N_2522);
and UO_215 (O_215,N_2563,N_2868);
nor UO_216 (O_216,N_2698,N_2822);
or UO_217 (O_217,N_2978,N_2971);
nor UO_218 (O_218,N_2791,N_2771);
or UO_219 (O_219,N_2606,N_2517);
nor UO_220 (O_220,N_2636,N_2540);
nor UO_221 (O_221,N_2834,N_2726);
nand UO_222 (O_222,N_2895,N_2657);
nor UO_223 (O_223,N_2806,N_2860);
nand UO_224 (O_224,N_2577,N_2511);
and UO_225 (O_225,N_2907,N_2570);
nor UO_226 (O_226,N_2695,N_2660);
and UO_227 (O_227,N_2852,N_2590);
and UO_228 (O_228,N_2653,N_2566);
or UO_229 (O_229,N_2705,N_2599);
nand UO_230 (O_230,N_2639,N_2934);
nor UO_231 (O_231,N_2891,N_2989);
nor UO_232 (O_232,N_2827,N_2598);
or UO_233 (O_233,N_2867,N_2770);
nand UO_234 (O_234,N_2910,N_2943);
and UO_235 (O_235,N_2607,N_2703);
and UO_236 (O_236,N_2651,N_2675);
nor UO_237 (O_237,N_2843,N_2591);
and UO_238 (O_238,N_2892,N_2733);
or UO_239 (O_239,N_2937,N_2882);
nor UO_240 (O_240,N_2984,N_2664);
and UO_241 (O_241,N_2872,N_2828);
nand UO_242 (O_242,N_2614,N_2802);
or UO_243 (O_243,N_2739,N_2732);
nor UO_244 (O_244,N_2579,N_2509);
nor UO_245 (O_245,N_2870,N_2773);
nor UO_246 (O_246,N_2818,N_2561);
nand UO_247 (O_247,N_2635,N_2672);
and UO_248 (O_248,N_2650,N_2594);
nand UO_249 (O_249,N_2756,N_2619);
nor UO_250 (O_250,N_2700,N_2936);
nand UO_251 (O_251,N_2744,N_2765);
nand UO_252 (O_252,N_2766,N_2734);
nor UO_253 (O_253,N_2887,N_2514);
nor UO_254 (O_254,N_2578,N_2849);
nor UO_255 (O_255,N_2691,N_2982);
nand UO_256 (O_256,N_2963,N_2833);
nand UO_257 (O_257,N_2953,N_2501);
and UO_258 (O_258,N_2889,N_2742);
or UO_259 (O_259,N_2730,N_2994);
nor UO_260 (O_260,N_2640,N_2713);
nand UO_261 (O_261,N_2606,N_2860);
or UO_262 (O_262,N_2536,N_2701);
nor UO_263 (O_263,N_2950,N_2581);
nor UO_264 (O_264,N_2564,N_2612);
and UO_265 (O_265,N_2867,N_2935);
nor UO_266 (O_266,N_2508,N_2911);
and UO_267 (O_267,N_2693,N_2976);
nor UO_268 (O_268,N_2839,N_2936);
and UO_269 (O_269,N_2588,N_2695);
nor UO_270 (O_270,N_2753,N_2979);
nor UO_271 (O_271,N_2698,N_2881);
nand UO_272 (O_272,N_2887,N_2718);
or UO_273 (O_273,N_2520,N_2987);
nand UO_274 (O_274,N_2842,N_2845);
and UO_275 (O_275,N_2992,N_2996);
and UO_276 (O_276,N_2879,N_2689);
and UO_277 (O_277,N_2861,N_2945);
or UO_278 (O_278,N_2710,N_2889);
nor UO_279 (O_279,N_2693,N_2941);
nor UO_280 (O_280,N_2614,N_2763);
nand UO_281 (O_281,N_2500,N_2980);
nor UO_282 (O_282,N_2669,N_2631);
and UO_283 (O_283,N_2724,N_2965);
nand UO_284 (O_284,N_2752,N_2798);
nand UO_285 (O_285,N_2869,N_2689);
or UO_286 (O_286,N_2851,N_2657);
nand UO_287 (O_287,N_2924,N_2773);
or UO_288 (O_288,N_2704,N_2980);
nand UO_289 (O_289,N_2589,N_2630);
nand UO_290 (O_290,N_2506,N_2725);
nor UO_291 (O_291,N_2688,N_2515);
or UO_292 (O_292,N_2907,N_2526);
nand UO_293 (O_293,N_2552,N_2993);
nor UO_294 (O_294,N_2735,N_2942);
or UO_295 (O_295,N_2669,N_2698);
or UO_296 (O_296,N_2503,N_2548);
nand UO_297 (O_297,N_2635,N_2607);
and UO_298 (O_298,N_2835,N_2983);
or UO_299 (O_299,N_2811,N_2796);
or UO_300 (O_300,N_2988,N_2677);
nand UO_301 (O_301,N_2756,N_2844);
or UO_302 (O_302,N_2536,N_2651);
nor UO_303 (O_303,N_2771,N_2678);
and UO_304 (O_304,N_2898,N_2505);
or UO_305 (O_305,N_2676,N_2610);
nand UO_306 (O_306,N_2914,N_2957);
or UO_307 (O_307,N_2967,N_2552);
nor UO_308 (O_308,N_2969,N_2756);
and UO_309 (O_309,N_2939,N_2901);
nor UO_310 (O_310,N_2890,N_2993);
nand UO_311 (O_311,N_2843,N_2831);
or UO_312 (O_312,N_2705,N_2813);
nor UO_313 (O_313,N_2922,N_2627);
nand UO_314 (O_314,N_2656,N_2740);
nor UO_315 (O_315,N_2791,N_2940);
or UO_316 (O_316,N_2618,N_2858);
nand UO_317 (O_317,N_2825,N_2627);
or UO_318 (O_318,N_2545,N_2507);
and UO_319 (O_319,N_2829,N_2725);
nand UO_320 (O_320,N_2605,N_2919);
or UO_321 (O_321,N_2693,N_2541);
and UO_322 (O_322,N_2781,N_2607);
or UO_323 (O_323,N_2627,N_2636);
nand UO_324 (O_324,N_2565,N_2598);
and UO_325 (O_325,N_2911,N_2563);
or UO_326 (O_326,N_2808,N_2579);
nand UO_327 (O_327,N_2872,N_2506);
or UO_328 (O_328,N_2597,N_2895);
nor UO_329 (O_329,N_2668,N_2581);
or UO_330 (O_330,N_2791,N_2932);
or UO_331 (O_331,N_2581,N_2783);
nand UO_332 (O_332,N_2701,N_2843);
or UO_333 (O_333,N_2868,N_2731);
and UO_334 (O_334,N_2715,N_2650);
nand UO_335 (O_335,N_2996,N_2693);
nand UO_336 (O_336,N_2953,N_2560);
nand UO_337 (O_337,N_2908,N_2775);
nor UO_338 (O_338,N_2591,N_2713);
and UO_339 (O_339,N_2747,N_2623);
and UO_340 (O_340,N_2780,N_2995);
nor UO_341 (O_341,N_2693,N_2910);
and UO_342 (O_342,N_2936,N_2932);
and UO_343 (O_343,N_2815,N_2679);
or UO_344 (O_344,N_2773,N_2966);
or UO_345 (O_345,N_2540,N_2571);
or UO_346 (O_346,N_2700,N_2612);
and UO_347 (O_347,N_2824,N_2724);
and UO_348 (O_348,N_2723,N_2599);
and UO_349 (O_349,N_2682,N_2830);
and UO_350 (O_350,N_2858,N_2750);
or UO_351 (O_351,N_2598,N_2616);
nor UO_352 (O_352,N_2843,N_2710);
and UO_353 (O_353,N_2645,N_2962);
and UO_354 (O_354,N_2843,N_2943);
nor UO_355 (O_355,N_2695,N_2675);
or UO_356 (O_356,N_2522,N_2906);
and UO_357 (O_357,N_2661,N_2952);
nor UO_358 (O_358,N_2862,N_2554);
nor UO_359 (O_359,N_2974,N_2711);
and UO_360 (O_360,N_2932,N_2876);
or UO_361 (O_361,N_2588,N_2626);
or UO_362 (O_362,N_2559,N_2864);
or UO_363 (O_363,N_2670,N_2525);
or UO_364 (O_364,N_2998,N_2857);
nand UO_365 (O_365,N_2531,N_2739);
nor UO_366 (O_366,N_2755,N_2826);
nor UO_367 (O_367,N_2520,N_2816);
nand UO_368 (O_368,N_2783,N_2946);
nor UO_369 (O_369,N_2812,N_2805);
nand UO_370 (O_370,N_2997,N_2783);
and UO_371 (O_371,N_2965,N_2818);
and UO_372 (O_372,N_2689,N_2768);
and UO_373 (O_373,N_2969,N_2988);
and UO_374 (O_374,N_2950,N_2773);
nand UO_375 (O_375,N_2834,N_2688);
nand UO_376 (O_376,N_2631,N_2941);
and UO_377 (O_377,N_2624,N_2944);
nor UO_378 (O_378,N_2562,N_2970);
and UO_379 (O_379,N_2811,N_2978);
and UO_380 (O_380,N_2646,N_2922);
or UO_381 (O_381,N_2676,N_2516);
nand UO_382 (O_382,N_2871,N_2677);
or UO_383 (O_383,N_2903,N_2550);
nor UO_384 (O_384,N_2875,N_2767);
nor UO_385 (O_385,N_2958,N_2969);
and UO_386 (O_386,N_2915,N_2978);
and UO_387 (O_387,N_2547,N_2532);
and UO_388 (O_388,N_2619,N_2579);
nand UO_389 (O_389,N_2737,N_2808);
nand UO_390 (O_390,N_2811,N_2802);
nand UO_391 (O_391,N_2754,N_2942);
and UO_392 (O_392,N_2596,N_2518);
and UO_393 (O_393,N_2624,N_2997);
or UO_394 (O_394,N_2709,N_2680);
nor UO_395 (O_395,N_2849,N_2635);
or UO_396 (O_396,N_2506,N_2957);
or UO_397 (O_397,N_2773,N_2813);
and UO_398 (O_398,N_2966,N_2744);
and UO_399 (O_399,N_2672,N_2549);
and UO_400 (O_400,N_2704,N_2889);
or UO_401 (O_401,N_2579,N_2629);
nor UO_402 (O_402,N_2712,N_2664);
nor UO_403 (O_403,N_2800,N_2550);
or UO_404 (O_404,N_2932,N_2567);
and UO_405 (O_405,N_2809,N_2968);
or UO_406 (O_406,N_2597,N_2608);
or UO_407 (O_407,N_2500,N_2713);
and UO_408 (O_408,N_2895,N_2799);
and UO_409 (O_409,N_2764,N_2926);
and UO_410 (O_410,N_2687,N_2789);
nand UO_411 (O_411,N_2770,N_2620);
nor UO_412 (O_412,N_2634,N_2987);
or UO_413 (O_413,N_2556,N_2878);
nand UO_414 (O_414,N_2897,N_2910);
or UO_415 (O_415,N_2870,N_2586);
and UO_416 (O_416,N_2836,N_2856);
and UO_417 (O_417,N_2667,N_2961);
or UO_418 (O_418,N_2950,N_2809);
nor UO_419 (O_419,N_2608,N_2748);
and UO_420 (O_420,N_2728,N_2909);
nand UO_421 (O_421,N_2608,N_2641);
or UO_422 (O_422,N_2671,N_2549);
nand UO_423 (O_423,N_2937,N_2567);
nor UO_424 (O_424,N_2582,N_2906);
and UO_425 (O_425,N_2732,N_2921);
or UO_426 (O_426,N_2658,N_2716);
xor UO_427 (O_427,N_2800,N_2797);
nor UO_428 (O_428,N_2678,N_2507);
nor UO_429 (O_429,N_2610,N_2844);
nand UO_430 (O_430,N_2983,N_2527);
nand UO_431 (O_431,N_2872,N_2757);
nor UO_432 (O_432,N_2908,N_2844);
and UO_433 (O_433,N_2757,N_2770);
nand UO_434 (O_434,N_2777,N_2857);
nor UO_435 (O_435,N_2715,N_2869);
or UO_436 (O_436,N_2635,N_2868);
nand UO_437 (O_437,N_2780,N_2614);
nand UO_438 (O_438,N_2952,N_2639);
or UO_439 (O_439,N_2516,N_2579);
nor UO_440 (O_440,N_2962,N_2654);
or UO_441 (O_441,N_2884,N_2681);
and UO_442 (O_442,N_2652,N_2820);
or UO_443 (O_443,N_2944,N_2529);
nand UO_444 (O_444,N_2696,N_2901);
nand UO_445 (O_445,N_2752,N_2761);
nand UO_446 (O_446,N_2930,N_2529);
and UO_447 (O_447,N_2847,N_2640);
or UO_448 (O_448,N_2558,N_2798);
nand UO_449 (O_449,N_2699,N_2573);
and UO_450 (O_450,N_2978,N_2535);
and UO_451 (O_451,N_2689,N_2910);
nand UO_452 (O_452,N_2562,N_2641);
and UO_453 (O_453,N_2863,N_2768);
and UO_454 (O_454,N_2845,N_2787);
and UO_455 (O_455,N_2844,N_2975);
or UO_456 (O_456,N_2874,N_2852);
nor UO_457 (O_457,N_2966,N_2834);
nand UO_458 (O_458,N_2870,N_2904);
and UO_459 (O_459,N_2518,N_2945);
nand UO_460 (O_460,N_2508,N_2891);
nor UO_461 (O_461,N_2549,N_2841);
or UO_462 (O_462,N_2711,N_2661);
nand UO_463 (O_463,N_2862,N_2751);
nand UO_464 (O_464,N_2759,N_2735);
nor UO_465 (O_465,N_2809,N_2858);
or UO_466 (O_466,N_2521,N_2758);
or UO_467 (O_467,N_2859,N_2777);
nand UO_468 (O_468,N_2900,N_2707);
or UO_469 (O_469,N_2620,N_2706);
and UO_470 (O_470,N_2815,N_2963);
nor UO_471 (O_471,N_2702,N_2742);
nand UO_472 (O_472,N_2599,N_2867);
and UO_473 (O_473,N_2742,N_2632);
and UO_474 (O_474,N_2637,N_2964);
nand UO_475 (O_475,N_2530,N_2694);
or UO_476 (O_476,N_2813,N_2981);
nor UO_477 (O_477,N_2632,N_2806);
and UO_478 (O_478,N_2612,N_2985);
nand UO_479 (O_479,N_2567,N_2754);
and UO_480 (O_480,N_2913,N_2834);
nand UO_481 (O_481,N_2501,N_2669);
nand UO_482 (O_482,N_2958,N_2920);
nand UO_483 (O_483,N_2713,N_2651);
nor UO_484 (O_484,N_2843,N_2975);
or UO_485 (O_485,N_2973,N_2583);
nor UO_486 (O_486,N_2979,N_2786);
nor UO_487 (O_487,N_2924,N_2562);
nor UO_488 (O_488,N_2612,N_2539);
nor UO_489 (O_489,N_2988,N_2562);
nand UO_490 (O_490,N_2557,N_2775);
nor UO_491 (O_491,N_2992,N_2928);
nor UO_492 (O_492,N_2817,N_2634);
or UO_493 (O_493,N_2503,N_2786);
nor UO_494 (O_494,N_2940,N_2759);
nor UO_495 (O_495,N_2663,N_2862);
or UO_496 (O_496,N_2906,N_2932);
and UO_497 (O_497,N_2769,N_2852);
nor UO_498 (O_498,N_2762,N_2703);
nand UO_499 (O_499,N_2893,N_2765);
endmodule