module basic_500_3000_500_4_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_438,In_320);
xor U1 (N_1,In_295,In_323);
xor U2 (N_2,In_262,In_21);
xnor U3 (N_3,In_368,In_42);
or U4 (N_4,In_7,In_240);
or U5 (N_5,In_330,In_374);
and U6 (N_6,In_12,In_165);
and U7 (N_7,In_243,In_68);
or U8 (N_8,In_465,In_134);
nor U9 (N_9,In_453,In_107);
and U10 (N_10,In_256,In_106);
and U11 (N_11,In_28,In_43);
xor U12 (N_12,In_285,In_226);
nand U13 (N_13,In_124,In_306);
nand U14 (N_14,In_213,In_141);
and U15 (N_15,In_187,In_400);
and U16 (N_16,In_377,In_392);
or U17 (N_17,In_476,In_376);
or U18 (N_18,In_364,In_190);
or U19 (N_19,In_215,In_2);
nor U20 (N_20,In_52,In_89);
xor U21 (N_21,In_200,In_229);
xor U22 (N_22,In_22,In_314);
xor U23 (N_23,In_432,In_211);
nor U24 (N_24,In_34,In_327);
and U25 (N_25,In_383,In_17);
and U26 (N_26,In_279,In_96);
and U27 (N_27,In_55,In_206);
or U28 (N_28,In_110,In_302);
xnor U29 (N_29,In_49,In_430);
nor U30 (N_30,In_56,In_102);
nor U31 (N_31,In_389,In_345);
xnor U32 (N_32,In_337,In_287);
nor U33 (N_33,In_201,In_118);
xor U34 (N_34,In_263,In_91);
and U35 (N_35,In_5,In_177);
nand U36 (N_36,In_322,In_149);
or U37 (N_37,In_253,In_444);
nand U38 (N_38,In_494,In_216);
xnor U39 (N_39,In_203,In_379);
or U40 (N_40,In_181,In_172);
xor U41 (N_41,In_144,In_58);
and U42 (N_42,In_169,In_62);
xnor U43 (N_43,In_398,In_120);
nor U44 (N_44,In_69,In_360);
nor U45 (N_45,In_268,In_157);
xnor U46 (N_46,In_164,In_93);
and U47 (N_47,In_353,In_418);
nand U48 (N_48,In_33,In_159);
nand U49 (N_49,In_207,In_98);
and U50 (N_50,In_171,In_309);
xor U51 (N_51,In_126,In_473);
nand U52 (N_52,In_297,In_127);
nand U53 (N_53,In_275,In_236);
xnor U54 (N_54,In_286,In_303);
or U55 (N_55,In_481,In_245);
or U56 (N_56,In_152,In_411);
nand U57 (N_57,In_45,In_371);
nand U58 (N_58,In_455,In_155);
nand U59 (N_59,In_188,In_274);
nor U60 (N_60,In_202,In_66);
and U61 (N_61,In_409,In_334);
xor U62 (N_62,In_51,In_86);
or U63 (N_63,In_162,In_385);
or U64 (N_64,In_233,In_46);
or U65 (N_65,In_339,In_183);
and U66 (N_66,In_490,In_460);
or U67 (N_67,In_457,In_63);
or U68 (N_68,In_145,In_242);
nor U69 (N_69,In_31,In_394);
or U70 (N_70,In_382,In_496);
and U71 (N_71,In_458,In_269);
and U72 (N_72,In_223,In_402);
nor U73 (N_73,In_447,In_255);
nand U74 (N_74,In_193,In_158);
xnor U75 (N_75,In_259,In_276);
nor U76 (N_76,In_357,In_270);
and U77 (N_77,In_308,In_37);
nor U78 (N_78,In_484,In_387);
and U79 (N_79,In_410,In_341);
nor U80 (N_80,In_142,In_271);
or U81 (N_81,In_60,In_186);
and U82 (N_82,In_273,In_300);
or U83 (N_83,In_347,In_29);
or U84 (N_84,In_264,In_289);
xor U85 (N_85,In_104,In_252);
xnor U86 (N_86,In_122,In_199);
xor U87 (N_87,In_317,In_426);
nor U88 (N_88,In_362,In_113);
nor U89 (N_89,In_340,In_282);
xnor U90 (N_90,In_161,In_332);
nand U91 (N_91,In_227,In_6);
nor U92 (N_92,In_491,In_50);
xnor U93 (N_93,In_54,In_479);
and U94 (N_94,In_160,In_280);
or U95 (N_95,In_417,In_100);
and U96 (N_96,In_76,In_436);
or U97 (N_97,In_194,In_214);
nand U98 (N_98,In_367,In_475);
nand U99 (N_99,In_355,In_131);
xor U100 (N_100,In_407,In_478);
and U101 (N_101,In_18,In_375);
nor U102 (N_102,In_492,In_220);
xnor U103 (N_103,In_112,In_146);
xnor U104 (N_104,In_20,In_210);
or U105 (N_105,In_11,In_442);
xor U106 (N_106,In_167,In_293);
or U107 (N_107,In_349,In_384);
nand U108 (N_108,In_153,In_221);
xor U109 (N_109,In_38,In_468);
xnor U110 (N_110,In_372,In_388);
or U111 (N_111,In_14,In_395);
xor U112 (N_112,In_333,In_1);
nor U113 (N_113,In_284,In_184);
nand U114 (N_114,In_36,In_361);
xnor U115 (N_115,In_448,In_331);
nor U116 (N_116,In_24,In_277);
nor U117 (N_117,In_425,In_163);
xnor U118 (N_118,In_325,In_235);
and U119 (N_119,In_72,In_498);
and U120 (N_120,In_486,In_440);
nor U121 (N_121,In_246,In_378);
nand U122 (N_122,In_4,In_396);
nor U123 (N_123,In_321,In_137);
and U124 (N_124,In_488,In_196);
nor U125 (N_125,In_154,In_487);
nor U126 (N_126,In_182,In_239);
or U127 (N_127,In_125,In_464);
nor U128 (N_128,In_472,In_23);
nand U129 (N_129,In_173,In_354);
nand U130 (N_130,In_316,In_180);
nor U131 (N_131,In_466,In_224);
and U132 (N_132,In_299,In_434);
or U133 (N_133,In_397,In_204);
and U134 (N_134,In_237,In_185);
nor U135 (N_135,In_70,In_129);
nor U136 (N_136,In_150,In_119);
nand U137 (N_137,In_446,In_209);
and U138 (N_138,In_261,In_307);
xnor U139 (N_139,In_168,In_231);
and U140 (N_140,In_393,In_421);
nand U141 (N_141,In_3,In_73);
xor U142 (N_142,In_75,In_195);
or U143 (N_143,In_249,In_391);
nor U144 (N_144,In_318,In_212);
nand U145 (N_145,In_495,In_380);
and U146 (N_146,In_310,In_413);
or U147 (N_147,In_250,In_156);
or U148 (N_148,In_420,In_480);
or U149 (N_149,In_443,In_390);
and U150 (N_150,In_117,In_40);
nand U151 (N_151,In_25,In_412);
nor U152 (N_152,In_433,In_175);
nand U153 (N_153,In_469,In_406);
nor U154 (N_154,In_77,In_366);
nand U155 (N_155,In_272,In_328);
nor U156 (N_156,In_359,In_350);
nand U157 (N_157,In_19,In_8);
nor U158 (N_158,In_133,In_419);
xnor U159 (N_159,In_352,In_462);
nand U160 (N_160,In_44,In_267);
nor U161 (N_161,In_192,In_461);
or U162 (N_162,In_166,In_311);
xor U163 (N_163,In_258,In_228);
or U164 (N_164,In_121,In_454);
or U165 (N_165,In_471,In_401);
or U166 (N_166,In_15,In_427);
or U167 (N_167,In_365,In_288);
nor U168 (N_168,In_429,In_290);
nand U169 (N_169,In_10,In_130);
nor U170 (N_170,In_151,In_416);
nand U171 (N_171,In_94,In_477);
nand U172 (N_172,In_219,In_452);
and U173 (N_173,In_474,In_281);
or U174 (N_174,In_422,In_48);
and U175 (N_175,In_399,In_301);
and U176 (N_176,In_16,In_67);
nor U177 (N_177,In_342,In_428);
nor U178 (N_178,In_450,In_65);
and U179 (N_179,In_27,In_81);
xnor U180 (N_180,In_9,In_338);
and U181 (N_181,In_304,In_74);
xor U182 (N_182,In_441,In_174);
xnor U183 (N_183,In_139,In_176);
nor U184 (N_184,In_248,In_305);
and U185 (N_185,In_489,In_241);
nand U186 (N_186,In_257,In_403);
nor U187 (N_187,In_415,In_108);
nor U188 (N_188,In_265,In_278);
and U189 (N_189,In_266,In_324);
nor U190 (N_190,In_348,In_115);
and U191 (N_191,In_283,In_53);
nand U192 (N_192,In_64,In_197);
nand U193 (N_193,In_111,In_191);
xnor U194 (N_194,In_346,In_456);
nand U195 (N_195,In_232,In_208);
or U196 (N_196,In_205,In_26);
and U197 (N_197,In_449,In_189);
or U198 (N_198,In_71,In_463);
xor U199 (N_199,In_373,In_147);
xnor U200 (N_200,In_140,In_136);
and U201 (N_201,In_312,In_87);
or U202 (N_202,In_381,In_408);
nor U203 (N_203,In_424,In_132);
or U204 (N_204,In_437,In_105);
and U205 (N_205,In_41,In_82);
xor U206 (N_206,In_336,In_222);
nor U207 (N_207,In_0,In_143);
nand U208 (N_208,In_90,In_445);
xor U209 (N_209,In_61,In_30);
nand U210 (N_210,In_198,In_326);
nor U211 (N_211,In_85,In_344);
xor U212 (N_212,In_356,In_88);
xor U213 (N_213,In_386,In_13);
or U214 (N_214,In_116,In_251);
xnor U215 (N_215,In_78,In_319);
or U216 (N_216,In_497,In_493);
and U217 (N_217,In_218,In_178);
xor U218 (N_218,In_260,In_39);
and U219 (N_219,In_298,In_217);
nand U220 (N_220,In_291,In_254);
nor U221 (N_221,In_138,In_95);
or U222 (N_222,In_329,In_369);
nor U223 (N_223,In_114,In_238);
xnor U224 (N_224,In_179,In_313);
and U225 (N_225,In_431,In_483);
xor U226 (N_226,In_225,In_123);
and U227 (N_227,In_99,In_92);
xor U228 (N_228,In_404,In_423);
and U229 (N_229,In_343,In_351);
nand U230 (N_230,In_244,In_57);
and U231 (N_231,In_59,In_79);
nand U232 (N_232,In_370,In_451);
nand U233 (N_233,In_128,In_47);
nor U234 (N_234,In_499,In_459);
or U235 (N_235,In_84,In_234);
or U236 (N_236,In_335,In_35);
and U237 (N_237,In_315,In_439);
nor U238 (N_238,In_470,In_101);
xnor U239 (N_239,In_83,In_363);
and U240 (N_240,In_296,In_358);
and U241 (N_241,In_247,In_292);
or U242 (N_242,In_485,In_109);
nand U243 (N_243,In_148,In_103);
xor U244 (N_244,In_467,In_80);
and U245 (N_245,In_405,In_97);
or U246 (N_246,In_482,In_32);
nor U247 (N_247,In_435,In_230);
and U248 (N_248,In_414,In_135);
nor U249 (N_249,In_170,In_294);
and U250 (N_250,In_373,In_27);
nand U251 (N_251,In_111,In_426);
nand U252 (N_252,In_349,In_51);
and U253 (N_253,In_91,In_232);
or U254 (N_254,In_498,In_499);
xnor U255 (N_255,In_287,In_479);
xor U256 (N_256,In_43,In_211);
nor U257 (N_257,In_74,In_441);
or U258 (N_258,In_223,In_387);
or U259 (N_259,In_111,In_97);
and U260 (N_260,In_178,In_246);
and U261 (N_261,In_344,In_155);
nor U262 (N_262,In_378,In_173);
xnor U263 (N_263,In_354,In_149);
or U264 (N_264,In_119,In_123);
or U265 (N_265,In_471,In_186);
or U266 (N_266,In_340,In_69);
nor U267 (N_267,In_276,In_327);
nor U268 (N_268,In_341,In_438);
xnor U269 (N_269,In_317,In_316);
or U270 (N_270,In_497,In_359);
nand U271 (N_271,In_177,In_327);
or U272 (N_272,In_212,In_388);
xor U273 (N_273,In_445,In_261);
nand U274 (N_274,In_253,In_252);
or U275 (N_275,In_384,In_458);
nor U276 (N_276,In_320,In_483);
xor U277 (N_277,In_191,In_14);
nor U278 (N_278,In_343,In_133);
or U279 (N_279,In_163,In_157);
and U280 (N_280,In_165,In_25);
nand U281 (N_281,In_367,In_321);
nor U282 (N_282,In_100,In_101);
xnor U283 (N_283,In_423,In_356);
nand U284 (N_284,In_257,In_248);
or U285 (N_285,In_361,In_329);
nor U286 (N_286,In_423,In_110);
nand U287 (N_287,In_216,In_143);
and U288 (N_288,In_180,In_446);
and U289 (N_289,In_381,In_293);
xnor U290 (N_290,In_113,In_346);
nor U291 (N_291,In_164,In_261);
and U292 (N_292,In_173,In_40);
nand U293 (N_293,In_207,In_428);
nand U294 (N_294,In_158,In_87);
or U295 (N_295,In_62,In_52);
xor U296 (N_296,In_442,In_87);
nand U297 (N_297,In_49,In_375);
nor U298 (N_298,In_26,In_406);
nand U299 (N_299,In_63,In_96);
or U300 (N_300,In_456,In_350);
nor U301 (N_301,In_114,In_316);
nor U302 (N_302,In_321,In_192);
nor U303 (N_303,In_181,In_274);
nor U304 (N_304,In_165,In_157);
or U305 (N_305,In_248,In_438);
and U306 (N_306,In_54,In_126);
nor U307 (N_307,In_199,In_443);
or U308 (N_308,In_203,In_286);
nand U309 (N_309,In_376,In_252);
and U310 (N_310,In_486,In_144);
nand U311 (N_311,In_116,In_321);
and U312 (N_312,In_109,In_390);
xnor U313 (N_313,In_424,In_43);
nor U314 (N_314,In_287,In_106);
nor U315 (N_315,In_3,In_285);
nor U316 (N_316,In_456,In_53);
xnor U317 (N_317,In_252,In_313);
xnor U318 (N_318,In_66,In_173);
or U319 (N_319,In_431,In_322);
xnor U320 (N_320,In_149,In_151);
nand U321 (N_321,In_15,In_3);
nor U322 (N_322,In_110,In_343);
nand U323 (N_323,In_476,In_281);
nor U324 (N_324,In_487,In_476);
nand U325 (N_325,In_436,In_467);
xor U326 (N_326,In_271,In_164);
and U327 (N_327,In_433,In_299);
nand U328 (N_328,In_289,In_251);
or U329 (N_329,In_82,In_15);
or U330 (N_330,In_170,In_424);
and U331 (N_331,In_328,In_191);
and U332 (N_332,In_260,In_75);
nand U333 (N_333,In_283,In_125);
xnor U334 (N_334,In_475,In_317);
and U335 (N_335,In_236,In_166);
nor U336 (N_336,In_405,In_400);
xor U337 (N_337,In_245,In_292);
or U338 (N_338,In_477,In_309);
nor U339 (N_339,In_49,In_359);
nand U340 (N_340,In_166,In_147);
and U341 (N_341,In_436,In_9);
nand U342 (N_342,In_166,In_160);
nand U343 (N_343,In_5,In_271);
and U344 (N_344,In_395,In_83);
nand U345 (N_345,In_492,In_37);
nor U346 (N_346,In_444,In_449);
nand U347 (N_347,In_402,In_127);
and U348 (N_348,In_330,In_285);
xnor U349 (N_349,In_92,In_24);
xnor U350 (N_350,In_82,In_381);
nor U351 (N_351,In_363,In_364);
nand U352 (N_352,In_134,In_120);
xnor U353 (N_353,In_367,In_132);
nand U354 (N_354,In_198,In_106);
and U355 (N_355,In_348,In_28);
or U356 (N_356,In_419,In_477);
nor U357 (N_357,In_454,In_169);
nor U358 (N_358,In_72,In_444);
or U359 (N_359,In_7,In_297);
nand U360 (N_360,In_424,In_362);
nor U361 (N_361,In_294,In_370);
and U362 (N_362,In_388,In_167);
nand U363 (N_363,In_228,In_15);
and U364 (N_364,In_439,In_475);
or U365 (N_365,In_451,In_147);
and U366 (N_366,In_415,In_461);
or U367 (N_367,In_76,In_182);
or U368 (N_368,In_130,In_488);
and U369 (N_369,In_73,In_0);
nor U370 (N_370,In_247,In_419);
and U371 (N_371,In_122,In_432);
nand U372 (N_372,In_423,In_257);
nor U373 (N_373,In_32,In_340);
nor U374 (N_374,In_1,In_399);
nor U375 (N_375,In_145,In_419);
and U376 (N_376,In_210,In_320);
or U377 (N_377,In_17,In_121);
nand U378 (N_378,In_469,In_190);
and U379 (N_379,In_284,In_441);
or U380 (N_380,In_334,In_48);
nand U381 (N_381,In_459,In_32);
or U382 (N_382,In_174,In_68);
and U383 (N_383,In_251,In_202);
or U384 (N_384,In_328,In_34);
xnor U385 (N_385,In_3,In_152);
xor U386 (N_386,In_447,In_404);
nand U387 (N_387,In_258,In_450);
and U388 (N_388,In_91,In_326);
xnor U389 (N_389,In_14,In_332);
nor U390 (N_390,In_129,In_125);
nor U391 (N_391,In_242,In_258);
nor U392 (N_392,In_207,In_233);
nand U393 (N_393,In_447,In_28);
nor U394 (N_394,In_356,In_478);
xor U395 (N_395,In_195,In_261);
and U396 (N_396,In_405,In_203);
or U397 (N_397,In_167,In_119);
and U398 (N_398,In_216,In_350);
nand U399 (N_399,In_470,In_414);
nand U400 (N_400,In_471,In_116);
and U401 (N_401,In_423,In_442);
or U402 (N_402,In_11,In_407);
nand U403 (N_403,In_120,In_122);
or U404 (N_404,In_122,In_157);
or U405 (N_405,In_394,In_66);
nand U406 (N_406,In_433,In_126);
nor U407 (N_407,In_409,In_362);
nand U408 (N_408,In_193,In_77);
or U409 (N_409,In_194,In_326);
nand U410 (N_410,In_63,In_435);
or U411 (N_411,In_457,In_234);
nand U412 (N_412,In_345,In_221);
and U413 (N_413,In_172,In_297);
nand U414 (N_414,In_42,In_476);
or U415 (N_415,In_335,In_126);
or U416 (N_416,In_260,In_138);
or U417 (N_417,In_242,In_401);
nor U418 (N_418,In_491,In_405);
and U419 (N_419,In_474,In_454);
or U420 (N_420,In_61,In_424);
xor U421 (N_421,In_371,In_407);
or U422 (N_422,In_128,In_49);
and U423 (N_423,In_492,In_135);
xor U424 (N_424,In_374,In_41);
xor U425 (N_425,In_253,In_198);
or U426 (N_426,In_423,In_20);
nor U427 (N_427,In_22,In_175);
and U428 (N_428,In_102,In_477);
or U429 (N_429,In_31,In_406);
nand U430 (N_430,In_115,In_445);
and U431 (N_431,In_290,In_472);
and U432 (N_432,In_477,In_480);
nor U433 (N_433,In_142,In_326);
or U434 (N_434,In_353,In_415);
or U435 (N_435,In_196,In_110);
xor U436 (N_436,In_376,In_318);
and U437 (N_437,In_10,In_152);
xnor U438 (N_438,In_324,In_240);
or U439 (N_439,In_432,In_386);
or U440 (N_440,In_493,In_238);
nor U441 (N_441,In_374,In_458);
or U442 (N_442,In_306,In_78);
or U443 (N_443,In_455,In_94);
nor U444 (N_444,In_275,In_366);
and U445 (N_445,In_438,In_483);
nand U446 (N_446,In_301,In_400);
and U447 (N_447,In_374,In_34);
or U448 (N_448,In_297,In_493);
nand U449 (N_449,In_400,In_214);
and U450 (N_450,In_43,In_318);
and U451 (N_451,In_221,In_44);
xnor U452 (N_452,In_310,In_196);
nand U453 (N_453,In_191,In_274);
nor U454 (N_454,In_237,In_14);
xor U455 (N_455,In_127,In_485);
nor U456 (N_456,In_258,In_26);
nand U457 (N_457,In_402,In_114);
and U458 (N_458,In_18,In_1);
nand U459 (N_459,In_148,In_138);
or U460 (N_460,In_107,In_269);
xor U461 (N_461,In_160,In_483);
or U462 (N_462,In_99,In_457);
nor U463 (N_463,In_318,In_340);
xnor U464 (N_464,In_412,In_463);
xnor U465 (N_465,In_243,In_141);
nand U466 (N_466,In_422,In_19);
and U467 (N_467,In_91,In_386);
nand U468 (N_468,In_384,In_57);
xnor U469 (N_469,In_282,In_440);
or U470 (N_470,In_151,In_287);
and U471 (N_471,In_75,In_381);
and U472 (N_472,In_357,In_146);
nand U473 (N_473,In_480,In_364);
or U474 (N_474,In_30,In_313);
or U475 (N_475,In_422,In_171);
and U476 (N_476,In_208,In_246);
xnor U477 (N_477,In_102,In_62);
or U478 (N_478,In_293,In_319);
nand U479 (N_479,In_54,In_218);
or U480 (N_480,In_422,In_346);
and U481 (N_481,In_170,In_44);
xnor U482 (N_482,In_139,In_340);
or U483 (N_483,In_368,In_96);
xnor U484 (N_484,In_261,In_74);
xor U485 (N_485,In_375,In_397);
or U486 (N_486,In_283,In_51);
nand U487 (N_487,In_123,In_207);
or U488 (N_488,In_479,In_423);
nand U489 (N_489,In_12,In_267);
xor U490 (N_490,In_3,In_335);
nand U491 (N_491,In_147,In_198);
and U492 (N_492,In_44,In_451);
nor U493 (N_493,In_130,In_359);
and U494 (N_494,In_139,In_478);
xnor U495 (N_495,In_282,In_179);
nor U496 (N_496,In_103,In_24);
or U497 (N_497,In_6,In_479);
or U498 (N_498,In_163,In_434);
xor U499 (N_499,In_11,In_340);
and U500 (N_500,In_212,In_45);
and U501 (N_501,In_244,In_309);
or U502 (N_502,In_349,In_210);
and U503 (N_503,In_237,In_474);
xor U504 (N_504,In_403,In_289);
xnor U505 (N_505,In_168,In_100);
xnor U506 (N_506,In_399,In_124);
nor U507 (N_507,In_355,In_362);
and U508 (N_508,In_235,In_26);
nand U509 (N_509,In_98,In_157);
and U510 (N_510,In_58,In_59);
or U511 (N_511,In_38,In_239);
and U512 (N_512,In_238,In_396);
or U513 (N_513,In_261,In_255);
and U514 (N_514,In_206,In_477);
nand U515 (N_515,In_168,In_10);
and U516 (N_516,In_90,In_73);
nor U517 (N_517,In_167,In_260);
and U518 (N_518,In_416,In_439);
nand U519 (N_519,In_423,In_86);
xnor U520 (N_520,In_16,In_152);
and U521 (N_521,In_347,In_395);
nor U522 (N_522,In_197,In_269);
nor U523 (N_523,In_405,In_299);
or U524 (N_524,In_286,In_116);
and U525 (N_525,In_458,In_340);
or U526 (N_526,In_320,In_489);
xor U527 (N_527,In_426,In_316);
xor U528 (N_528,In_226,In_458);
xnor U529 (N_529,In_226,In_455);
nand U530 (N_530,In_350,In_212);
and U531 (N_531,In_454,In_151);
or U532 (N_532,In_294,In_227);
xnor U533 (N_533,In_277,In_430);
and U534 (N_534,In_442,In_30);
nor U535 (N_535,In_388,In_194);
xnor U536 (N_536,In_285,In_275);
nand U537 (N_537,In_303,In_148);
nand U538 (N_538,In_333,In_357);
xor U539 (N_539,In_397,In_94);
xor U540 (N_540,In_322,In_462);
xnor U541 (N_541,In_226,In_144);
or U542 (N_542,In_132,In_20);
nand U543 (N_543,In_280,In_58);
xor U544 (N_544,In_322,In_32);
xor U545 (N_545,In_257,In_61);
xor U546 (N_546,In_190,In_317);
nor U547 (N_547,In_111,In_307);
and U548 (N_548,In_230,In_57);
nand U549 (N_549,In_230,In_372);
xnor U550 (N_550,In_90,In_228);
nor U551 (N_551,In_60,In_20);
or U552 (N_552,In_191,In_317);
or U553 (N_553,In_199,In_448);
xnor U554 (N_554,In_225,In_363);
nor U555 (N_555,In_99,In_84);
nand U556 (N_556,In_316,In_497);
xnor U557 (N_557,In_47,In_171);
nor U558 (N_558,In_330,In_184);
nor U559 (N_559,In_202,In_433);
or U560 (N_560,In_203,In_57);
xor U561 (N_561,In_326,In_325);
or U562 (N_562,In_380,In_425);
nand U563 (N_563,In_336,In_303);
nor U564 (N_564,In_102,In_20);
or U565 (N_565,In_431,In_376);
nand U566 (N_566,In_159,In_329);
and U567 (N_567,In_163,In_412);
and U568 (N_568,In_321,In_462);
or U569 (N_569,In_248,In_206);
nand U570 (N_570,In_252,In_397);
or U571 (N_571,In_38,In_406);
nor U572 (N_572,In_225,In_401);
nor U573 (N_573,In_9,In_206);
or U574 (N_574,In_143,In_106);
and U575 (N_575,In_79,In_20);
nand U576 (N_576,In_117,In_219);
nor U577 (N_577,In_50,In_440);
and U578 (N_578,In_233,In_484);
nor U579 (N_579,In_205,In_119);
nand U580 (N_580,In_193,In_80);
nor U581 (N_581,In_144,In_477);
and U582 (N_582,In_486,In_235);
or U583 (N_583,In_30,In_460);
nand U584 (N_584,In_74,In_318);
or U585 (N_585,In_152,In_323);
nand U586 (N_586,In_34,In_11);
xor U587 (N_587,In_9,In_113);
and U588 (N_588,In_481,In_239);
nor U589 (N_589,In_117,In_87);
nor U590 (N_590,In_126,In_1);
and U591 (N_591,In_138,In_310);
nand U592 (N_592,In_435,In_157);
nand U593 (N_593,In_66,In_56);
nand U594 (N_594,In_221,In_16);
nor U595 (N_595,In_225,In_10);
or U596 (N_596,In_94,In_331);
nand U597 (N_597,In_474,In_40);
nor U598 (N_598,In_338,In_273);
nor U599 (N_599,In_224,In_447);
nor U600 (N_600,In_171,In_119);
and U601 (N_601,In_417,In_251);
nand U602 (N_602,In_1,In_257);
xnor U603 (N_603,In_385,In_157);
and U604 (N_604,In_139,In_238);
nand U605 (N_605,In_414,In_437);
or U606 (N_606,In_266,In_67);
xnor U607 (N_607,In_132,In_142);
nand U608 (N_608,In_56,In_279);
xnor U609 (N_609,In_375,In_293);
nand U610 (N_610,In_225,In_388);
nand U611 (N_611,In_252,In_475);
nor U612 (N_612,In_106,In_118);
nor U613 (N_613,In_85,In_494);
xnor U614 (N_614,In_431,In_217);
nor U615 (N_615,In_189,In_93);
or U616 (N_616,In_5,In_456);
nand U617 (N_617,In_87,In_379);
xor U618 (N_618,In_242,In_448);
and U619 (N_619,In_476,In_221);
and U620 (N_620,In_440,In_149);
nand U621 (N_621,In_231,In_256);
or U622 (N_622,In_74,In_437);
or U623 (N_623,In_337,In_487);
nor U624 (N_624,In_0,In_464);
xnor U625 (N_625,In_53,In_307);
nand U626 (N_626,In_310,In_81);
or U627 (N_627,In_161,In_131);
xnor U628 (N_628,In_155,In_138);
nand U629 (N_629,In_149,In_430);
or U630 (N_630,In_293,In_356);
and U631 (N_631,In_74,In_397);
xor U632 (N_632,In_326,In_463);
nand U633 (N_633,In_223,In_417);
nand U634 (N_634,In_251,In_315);
xor U635 (N_635,In_375,In_391);
nand U636 (N_636,In_180,In_122);
or U637 (N_637,In_159,In_480);
nor U638 (N_638,In_92,In_388);
nor U639 (N_639,In_149,In_141);
or U640 (N_640,In_196,In_61);
nor U641 (N_641,In_413,In_174);
nor U642 (N_642,In_219,In_114);
or U643 (N_643,In_376,In_423);
nand U644 (N_644,In_312,In_24);
or U645 (N_645,In_236,In_389);
nor U646 (N_646,In_3,In_385);
and U647 (N_647,In_190,In_208);
nand U648 (N_648,In_139,In_158);
or U649 (N_649,In_92,In_214);
or U650 (N_650,In_129,In_160);
and U651 (N_651,In_370,In_405);
and U652 (N_652,In_48,In_138);
nor U653 (N_653,In_233,In_200);
and U654 (N_654,In_121,In_478);
or U655 (N_655,In_486,In_78);
nand U656 (N_656,In_373,In_94);
and U657 (N_657,In_323,In_404);
and U658 (N_658,In_235,In_170);
nand U659 (N_659,In_127,In_358);
or U660 (N_660,In_107,In_174);
nand U661 (N_661,In_147,In_211);
or U662 (N_662,In_373,In_346);
and U663 (N_663,In_246,In_473);
nand U664 (N_664,In_403,In_200);
nand U665 (N_665,In_427,In_205);
nor U666 (N_666,In_251,In_99);
xnor U667 (N_667,In_435,In_423);
nand U668 (N_668,In_160,In_297);
and U669 (N_669,In_90,In_128);
nor U670 (N_670,In_58,In_406);
and U671 (N_671,In_408,In_316);
nor U672 (N_672,In_45,In_200);
or U673 (N_673,In_106,In_221);
or U674 (N_674,In_197,In_170);
nor U675 (N_675,In_98,In_417);
and U676 (N_676,In_209,In_124);
xor U677 (N_677,In_208,In_33);
and U678 (N_678,In_278,In_346);
xnor U679 (N_679,In_327,In_95);
or U680 (N_680,In_434,In_353);
and U681 (N_681,In_279,In_156);
nor U682 (N_682,In_12,In_22);
nor U683 (N_683,In_187,In_433);
xnor U684 (N_684,In_247,In_457);
or U685 (N_685,In_473,In_498);
or U686 (N_686,In_350,In_353);
nand U687 (N_687,In_422,In_103);
and U688 (N_688,In_315,In_336);
or U689 (N_689,In_438,In_255);
or U690 (N_690,In_286,In_289);
nor U691 (N_691,In_46,In_327);
or U692 (N_692,In_479,In_265);
and U693 (N_693,In_19,In_492);
or U694 (N_694,In_191,In_467);
or U695 (N_695,In_325,In_341);
nand U696 (N_696,In_264,In_360);
nand U697 (N_697,In_285,In_103);
and U698 (N_698,In_56,In_400);
xor U699 (N_699,In_19,In_88);
or U700 (N_700,In_52,In_332);
nand U701 (N_701,In_371,In_444);
xnor U702 (N_702,In_304,In_41);
nor U703 (N_703,In_226,In_275);
xor U704 (N_704,In_33,In_390);
or U705 (N_705,In_477,In_145);
nor U706 (N_706,In_466,In_145);
and U707 (N_707,In_39,In_165);
nor U708 (N_708,In_410,In_66);
or U709 (N_709,In_10,In_260);
and U710 (N_710,In_405,In_225);
or U711 (N_711,In_252,In_297);
nor U712 (N_712,In_56,In_244);
or U713 (N_713,In_362,In_102);
and U714 (N_714,In_117,In_448);
nor U715 (N_715,In_302,In_49);
nand U716 (N_716,In_455,In_485);
nor U717 (N_717,In_234,In_87);
or U718 (N_718,In_329,In_487);
nand U719 (N_719,In_317,In_117);
xnor U720 (N_720,In_490,In_314);
or U721 (N_721,In_333,In_48);
nand U722 (N_722,In_226,In_495);
nor U723 (N_723,In_72,In_476);
xor U724 (N_724,In_95,In_463);
nor U725 (N_725,In_360,In_167);
xnor U726 (N_726,In_460,In_104);
nand U727 (N_727,In_301,In_66);
nor U728 (N_728,In_217,In_275);
nand U729 (N_729,In_49,In_478);
xnor U730 (N_730,In_470,In_185);
xnor U731 (N_731,In_43,In_279);
xor U732 (N_732,In_56,In_75);
nor U733 (N_733,In_384,In_102);
xor U734 (N_734,In_464,In_346);
nor U735 (N_735,In_25,In_430);
and U736 (N_736,In_200,In_148);
and U737 (N_737,In_426,In_337);
nand U738 (N_738,In_194,In_366);
nand U739 (N_739,In_323,In_169);
xnor U740 (N_740,In_92,In_456);
or U741 (N_741,In_126,In_437);
nand U742 (N_742,In_159,In_405);
and U743 (N_743,In_125,In_318);
or U744 (N_744,In_347,In_216);
or U745 (N_745,In_351,In_378);
nand U746 (N_746,In_124,In_87);
nor U747 (N_747,In_21,In_347);
xor U748 (N_748,In_66,In_352);
nand U749 (N_749,In_301,In_243);
and U750 (N_750,N_688,N_262);
and U751 (N_751,N_62,N_206);
and U752 (N_752,N_265,N_375);
nor U753 (N_753,N_521,N_92);
or U754 (N_754,N_115,N_294);
nand U755 (N_755,N_233,N_647);
nand U756 (N_756,N_378,N_247);
xnor U757 (N_757,N_131,N_31);
or U758 (N_758,N_186,N_185);
nor U759 (N_759,N_473,N_248);
xor U760 (N_760,N_741,N_229);
or U761 (N_761,N_5,N_582);
nand U762 (N_762,N_59,N_729);
and U763 (N_763,N_161,N_138);
nor U764 (N_764,N_197,N_282);
nor U765 (N_765,N_566,N_419);
xor U766 (N_766,N_699,N_142);
or U767 (N_767,N_668,N_71);
nor U768 (N_768,N_103,N_245);
nor U769 (N_769,N_237,N_691);
xnor U770 (N_770,N_682,N_448);
and U771 (N_771,N_725,N_231);
nand U772 (N_772,N_158,N_662);
nor U773 (N_773,N_24,N_174);
xnor U774 (N_774,N_354,N_634);
nor U775 (N_775,N_350,N_433);
xor U776 (N_776,N_496,N_11);
xnor U777 (N_777,N_405,N_361);
and U778 (N_778,N_303,N_539);
nor U779 (N_779,N_167,N_671);
nand U780 (N_780,N_641,N_373);
or U781 (N_781,N_123,N_213);
nand U782 (N_782,N_608,N_722);
nor U783 (N_783,N_430,N_181);
and U784 (N_784,N_68,N_645);
nor U785 (N_785,N_491,N_385);
xnor U786 (N_786,N_441,N_408);
or U787 (N_787,N_575,N_505);
and U788 (N_788,N_162,N_402);
nor U789 (N_789,N_65,N_76);
nand U790 (N_790,N_281,N_222);
and U791 (N_791,N_145,N_79);
or U792 (N_792,N_458,N_555);
and U793 (N_793,N_611,N_207);
nand U794 (N_794,N_4,N_696);
and U795 (N_795,N_352,N_88);
nand U796 (N_796,N_669,N_134);
nor U797 (N_797,N_442,N_193);
xor U798 (N_798,N_58,N_178);
and U799 (N_799,N_531,N_588);
and U800 (N_800,N_326,N_345);
xnor U801 (N_801,N_549,N_100);
nand U802 (N_802,N_93,N_733);
nand U803 (N_803,N_331,N_340);
nand U804 (N_804,N_509,N_417);
or U805 (N_805,N_495,N_409);
xnor U806 (N_806,N_276,N_238);
nand U807 (N_807,N_347,N_426);
nor U808 (N_808,N_613,N_561);
nor U809 (N_809,N_150,N_57);
nor U810 (N_810,N_239,N_199);
or U811 (N_811,N_371,N_601);
nor U812 (N_812,N_342,N_703);
nor U813 (N_813,N_676,N_438);
and U814 (N_814,N_410,N_586);
or U815 (N_815,N_114,N_536);
nor U816 (N_816,N_470,N_716);
or U817 (N_817,N_657,N_344);
or U818 (N_818,N_674,N_396);
nor U819 (N_819,N_453,N_21);
or U820 (N_820,N_631,N_3);
nand U821 (N_821,N_523,N_590);
nand U822 (N_822,N_528,N_388);
xor U823 (N_823,N_450,N_680);
and U824 (N_824,N_60,N_745);
xor U825 (N_825,N_216,N_368);
nand U826 (N_826,N_36,N_715);
nand U827 (N_827,N_72,N_567);
xor U828 (N_828,N_83,N_609);
nor U829 (N_829,N_704,N_32);
nand U830 (N_830,N_126,N_494);
xnor U831 (N_831,N_358,N_220);
or U832 (N_832,N_116,N_295);
nand U833 (N_833,N_292,N_343);
or U834 (N_834,N_141,N_477);
xor U835 (N_835,N_273,N_687);
nor U836 (N_836,N_339,N_66);
or U837 (N_837,N_573,N_70);
xnor U838 (N_838,N_746,N_196);
nor U839 (N_839,N_359,N_501);
and U840 (N_840,N_443,N_532);
or U841 (N_841,N_267,N_259);
xor U842 (N_842,N_12,N_290);
and U843 (N_843,N_382,N_82);
and U844 (N_844,N_425,N_614);
or U845 (N_845,N_377,N_683);
xor U846 (N_846,N_8,N_380);
xor U847 (N_847,N_125,N_133);
xor U848 (N_848,N_61,N_740);
nand U849 (N_849,N_702,N_654);
nor U850 (N_850,N_283,N_297);
xor U851 (N_851,N_249,N_154);
xnor U852 (N_852,N_665,N_395);
and U853 (N_853,N_527,N_323);
xor U854 (N_854,N_315,N_617);
and U855 (N_855,N_192,N_170);
nor U856 (N_856,N_436,N_466);
and U857 (N_857,N_399,N_285);
or U858 (N_858,N_338,N_296);
xor U859 (N_859,N_626,N_204);
or U860 (N_860,N_306,N_101);
xor U861 (N_861,N_498,N_602);
and U862 (N_862,N_45,N_153);
or U863 (N_863,N_490,N_41);
and U864 (N_864,N_708,N_74);
or U865 (N_865,N_263,N_73);
xor U866 (N_866,N_270,N_210);
nor U867 (N_867,N_455,N_554);
xor U868 (N_868,N_493,N_563);
or U869 (N_869,N_42,N_445);
nor U870 (N_870,N_714,N_726);
xor U871 (N_871,N_415,N_387);
and U872 (N_872,N_530,N_413);
or U873 (N_873,N_578,N_581);
xnor U874 (N_874,N_564,N_320);
nand U875 (N_875,N_0,N_289);
nand U876 (N_876,N_19,N_749);
and U877 (N_877,N_401,N_97);
and U878 (N_878,N_463,N_544);
nor U879 (N_879,N_589,N_209);
or U880 (N_880,N_743,N_191);
nand U881 (N_881,N_363,N_705);
and U882 (N_882,N_13,N_164);
and U883 (N_883,N_333,N_362);
or U884 (N_884,N_595,N_597);
and U885 (N_885,N_302,N_291);
or U886 (N_886,N_400,N_475);
or U887 (N_887,N_454,N_310);
xnor U888 (N_888,N_639,N_610);
or U889 (N_889,N_176,N_328);
nor U890 (N_890,N_713,N_85);
nor U891 (N_891,N_353,N_659);
or U892 (N_892,N_271,N_137);
nand U893 (N_893,N_51,N_132);
xor U894 (N_894,N_511,N_288);
nor U895 (N_895,N_481,N_689);
nand U896 (N_896,N_707,N_542);
or U897 (N_897,N_633,N_616);
or U898 (N_898,N_718,N_661);
nand U899 (N_899,N_488,N_421);
nor U900 (N_900,N_44,N_151);
and U901 (N_901,N_166,N_640);
nand U902 (N_902,N_155,N_356);
nor U903 (N_903,N_200,N_658);
nand U904 (N_904,N_479,N_651);
nor U905 (N_905,N_225,N_27);
xnor U906 (N_906,N_428,N_143);
nor U907 (N_907,N_317,N_129);
nand U908 (N_908,N_457,N_656);
nor U909 (N_909,N_46,N_636);
or U910 (N_910,N_619,N_747);
nor U911 (N_911,N_33,N_627);
and U912 (N_912,N_175,N_630);
xnor U913 (N_913,N_223,N_10);
nor U914 (N_914,N_111,N_25);
nand U915 (N_915,N_731,N_712);
xor U916 (N_916,N_230,N_513);
nand U917 (N_917,N_605,N_565);
nor U918 (N_918,N_140,N_414);
or U919 (N_919,N_412,N_355);
nor U920 (N_920,N_337,N_144);
or U921 (N_921,N_105,N_742);
xnor U922 (N_922,N_548,N_615);
xor U923 (N_923,N_20,N_468);
or U924 (N_924,N_330,N_594);
nor U925 (N_925,N_357,N_508);
and U926 (N_926,N_472,N_709);
nand U927 (N_927,N_251,N_35);
xor U928 (N_928,N_246,N_182);
and U929 (N_929,N_275,N_557);
or U930 (N_930,N_489,N_205);
and U931 (N_931,N_525,N_723);
nand U932 (N_932,N_341,N_690);
nor U933 (N_933,N_404,N_467);
nand U934 (N_934,N_679,N_692);
xor U935 (N_935,N_541,N_706);
and U936 (N_936,N_17,N_540);
or U937 (N_937,N_9,N_701);
nand U938 (N_938,N_424,N_560);
xor U939 (N_939,N_451,N_287);
xor U940 (N_940,N_434,N_644);
or U941 (N_941,N_519,N_598);
xnor U942 (N_942,N_304,N_695);
or U943 (N_943,N_201,N_214);
nand U944 (N_944,N_406,N_465);
or U945 (N_945,N_348,N_313);
and U946 (N_946,N_571,N_681);
and U947 (N_947,N_524,N_28);
or U948 (N_948,N_177,N_484);
nor U949 (N_949,N_322,N_556);
and U950 (N_950,N_146,N_535);
nand U951 (N_951,N_600,N_183);
or U952 (N_952,N_96,N_346);
and U953 (N_953,N_208,N_432);
or U954 (N_954,N_537,N_579);
or U955 (N_955,N_711,N_300);
xor U956 (N_956,N_34,N_364);
nand U957 (N_957,N_612,N_266);
xor U958 (N_958,N_121,N_585);
or U959 (N_959,N_40,N_685);
xnor U960 (N_960,N_316,N_215);
and U961 (N_961,N_95,N_301);
nor U962 (N_962,N_739,N_667);
nor U963 (N_963,N_622,N_211);
or U964 (N_964,N_234,N_108);
nand U965 (N_965,N_437,N_336);
xor U966 (N_966,N_515,N_469);
xor U967 (N_967,N_516,N_94);
nor U968 (N_968,N_91,N_666);
or U969 (N_969,N_117,N_135);
xnor U970 (N_970,N_738,N_492);
and U971 (N_971,N_254,N_390);
nand U972 (N_972,N_386,N_156);
and U973 (N_973,N_422,N_360);
nand U974 (N_974,N_243,N_190);
nand U975 (N_975,N_717,N_570);
nor U976 (N_976,N_99,N_648);
xnor U977 (N_977,N_700,N_744);
or U978 (N_978,N_47,N_652);
or U979 (N_979,N_486,N_384);
xnor U980 (N_980,N_50,N_748);
nand U981 (N_981,N_67,N_39);
nor U982 (N_982,N_52,N_698);
nand U983 (N_983,N_366,N_502);
nand U984 (N_984,N_507,N_423);
or U985 (N_985,N_258,N_420);
or U986 (N_986,N_471,N_580);
nand U987 (N_987,N_697,N_591);
nand U988 (N_988,N_512,N_499);
nor U989 (N_989,N_221,N_621);
nand U990 (N_990,N_478,N_553);
nor U991 (N_991,N_212,N_514);
and U992 (N_992,N_632,N_277);
or U993 (N_993,N_311,N_643);
nand U994 (N_994,N_449,N_558);
or U995 (N_995,N_672,N_256);
nor U996 (N_996,N_351,N_280);
and U997 (N_997,N_260,N_124);
or U998 (N_998,N_278,N_224);
nor U999 (N_999,N_187,N_547);
and U1000 (N_1000,N_482,N_653);
nand U1001 (N_1001,N_416,N_628);
and U1002 (N_1002,N_165,N_106);
xor U1003 (N_1003,N_431,N_86);
or U1004 (N_1004,N_568,N_128);
or U1005 (N_1005,N_383,N_506);
and U1006 (N_1006,N_429,N_664);
and U1007 (N_1007,N_533,N_252);
and U1008 (N_1008,N_319,N_389);
nand U1009 (N_1009,N_381,N_15);
nand U1010 (N_1010,N_577,N_370);
nand U1011 (N_1011,N_649,N_329);
xnor U1012 (N_1012,N_241,N_309);
nand U1013 (N_1013,N_675,N_180);
xor U1014 (N_1014,N_157,N_104);
xor U1015 (N_1015,N_195,N_550);
xnor U1016 (N_1016,N_737,N_149);
nor U1017 (N_1017,N_299,N_198);
and U1018 (N_1018,N_179,N_474);
xor U1019 (N_1019,N_526,N_418);
or U1020 (N_1020,N_684,N_269);
nand U1021 (N_1021,N_148,N_456);
xor U1022 (N_1022,N_112,N_462);
and U1023 (N_1023,N_604,N_122);
nand U1024 (N_1024,N_440,N_37);
and U1025 (N_1025,N_736,N_551);
nand U1026 (N_1026,N_485,N_110);
and U1027 (N_1027,N_264,N_274);
and U1028 (N_1028,N_487,N_584);
nor U1029 (N_1029,N_646,N_54);
or U1030 (N_1030,N_253,N_2);
xor U1031 (N_1031,N_1,N_14);
nand U1032 (N_1032,N_724,N_242);
and U1033 (N_1033,N_228,N_332);
xor U1034 (N_1034,N_314,N_435);
xor U1035 (N_1035,N_219,N_75);
xnor U1036 (N_1036,N_147,N_497);
xor U1037 (N_1037,N_618,N_369);
nor U1038 (N_1038,N_624,N_444);
or U1039 (N_1039,N_48,N_98);
nand U1040 (N_1040,N_307,N_394);
nor U1041 (N_1041,N_308,N_673);
or U1042 (N_1042,N_587,N_255);
or U1043 (N_1043,N_43,N_305);
xnor U1044 (N_1044,N_372,N_26);
or U1045 (N_1045,N_407,N_572);
and U1046 (N_1046,N_504,N_293);
or U1047 (N_1047,N_272,N_203);
and U1048 (N_1048,N_78,N_545);
or U1049 (N_1049,N_152,N_226);
nand U1050 (N_1050,N_286,N_374);
xnor U1051 (N_1051,N_284,N_503);
and U1052 (N_1052,N_327,N_120);
nor U1053 (N_1053,N_727,N_459);
and U1054 (N_1054,N_694,N_655);
or U1055 (N_1055,N_599,N_240);
nand U1056 (N_1056,N_49,N_534);
xor U1057 (N_1057,N_7,N_38);
nor U1058 (N_1058,N_660,N_119);
nand U1059 (N_1059,N_173,N_89);
nand U1060 (N_1060,N_257,N_202);
xor U1061 (N_1061,N_169,N_593);
or U1062 (N_1062,N_298,N_734);
xnor U1063 (N_1063,N_427,N_63);
and U1064 (N_1064,N_642,N_510);
xnor U1065 (N_1065,N_393,N_476);
nand U1066 (N_1066,N_693,N_629);
or U1067 (N_1067,N_268,N_194);
xnor U1068 (N_1068,N_102,N_188);
and U1069 (N_1069,N_719,N_29);
and U1070 (N_1070,N_367,N_81);
xor U1071 (N_1071,N_6,N_677);
nor U1072 (N_1072,N_480,N_379);
xor U1073 (N_1073,N_325,N_335);
or U1074 (N_1074,N_500,N_235);
or U1075 (N_1075,N_244,N_638);
or U1076 (N_1076,N_318,N_227);
nand U1077 (N_1077,N_184,N_569);
nor U1078 (N_1078,N_607,N_452);
xor U1079 (N_1079,N_447,N_168);
xnor U1080 (N_1080,N_517,N_543);
or U1081 (N_1081,N_55,N_637);
nor U1082 (N_1082,N_461,N_365);
or U1083 (N_1083,N_650,N_625);
nand U1084 (N_1084,N_136,N_232);
nand U1085 (N_1085,N_218,N_163);
or U1086 (N_1086,N_411,N_446);
nand U1087 (N_1087,N_90,N_576);
xor U1088 (N_1088,N_127,N_189);
xnor U1089 (N_1089,N_16,N_520);
xnor U1090 (N_1090,N_23,N_710);
nand U1091 (N_1091,N_171,N_22);
or U1092 (N_1092,N_518,N_312);
and U1093 (N_1093,N_130,N_139);
or U1094 (N_1094,N_56,N_728);
or U1095 (N_1095,N_522,N_30);
and U1096 (N_1096,N_321,N_670);
and U1097 (N_1097,N_686,N_606);
or U1098 (N_1098,N_107,N_583);
and U1099 (N_1099,N_87,N_663);
xor U1100 (N_1100,N_250,N_217);
xor U1101 (N_1101,N_392,N_460);
or U1102 (N_1102,N_160,N_559);
nor U1103 (N_1103,N_720,N_118);
or U1104 (N_1104,N_620,N_721);
nor U1105 (N_1105,N_349,N_172);
or U1106 (N_1106,N_483,N_529);
xor U1107 (N_1107,N_562,N_398);
or U1108 (N_1108,N_64,N_574);
xnor U1109 (N_1109,N_732,N_69);
nand U1110 (N_1110,N_538,N_439);
nor U1111 (N_1111,N_376,N_635);
nand U1112 (N_1112,N_113,N_403);
or U1113 (N_1113,N_84,N_109);
and U1114 (N_1114,N_334,N_236);
or U1115 (N_1115,N_53,N_391);
nor U1116 (N_1116,N_735,N_80);
nand U1117 (N_1117,N_603,N_552);
or U1118 (N_1118,N_261,N_77);
nand U1119 (N_1119,N_730,N_592);
nand U1120 (N_1120,N_279,N_623);
nor U1121 (N_1121,N_324,N_546);
nand U1122 (N_1122,N_678,N_397);
and U1123 (N_1123,N_596,N_159);
nand U1124 (N_1124,N_464,N_18);
or U1125 (N_1125,N_272,N_31);
and U1126 (N_1126,N_481,N_178);
nor U1127 (N_1127,N_92,N_547);
xnor U1128 (N_1128,N_640,N_388);
or U1129 (N_1129,N_490,N_294);
and U1130 (N_1130,N_344,N_281);
nand U1131 (N_1131,N_346,N_354);
xor U1132 (N_1132,N_206,N_712);
nand U1133 (N_1133,N_132,N_598);
nor U1134 (N_1134,N_520,N_261);
and U1135 (N_1135,N_32,N_320);
nand U1136 (N_1136,N_544,N_278);
xor U1137 (N_1137,N_285,N_450);
nand U1138 (N_1138,N_629,N_142);
nand U1139 (N_1139,N_16,N_598);
and U1140 (N_1140,N_428,N_730);
nor U1141 (N_1141,N_494,N_208);
xor U1142 (N_1142,N_509,N_472);
xor U1143 (N_1143,N_330,N_224);
nor U1144 (N_1144,N_374,N_316);
nor U1145 (N_1145,N_92,N_115);
nand U1146 (N_1146,N_543,N_706);
nand U1147 (N_1147,N_135,N_149);
xor U1148 (N_1148,N_360,N_347);
xor U1149 (N_1149,N_562,N_503);
nand U1150 (N_1150,N_735,N_550);
or U1151 (N_1151,N_460,N_355);
or U1152 (N_1152,N_516,N_513);
nand U1153 (N_1153,N_263,N_362);
or U1154 (N_1154,N_739,N_202);
or U1155 (N_1155,N_141,N_372);
xnor U1156 (N_1156,N_734,N_409);
nor U1157 (N_1157,N_13,N_100);
nor U1158 (N_1158,N_503,N_45);
or U1159 (N_1159,N_345,N_334);
and U1160 (N_1160,N_127,N_436);
or U1161 (N_1161,N_273,N_322);
or U1162 (N_1162,N_657,N_598);
nor U1163 (N_1163,N_60,N_333);
nand U1164 (N_1164,N_357,N_230);
nor U1165 (N_1165,N_207,N_219);
or U1166 (N_1166,N_296,N_74);
xnor U1167 (N_1167,N_423,N_11);
nor U1168 (N_1168,N_418,N_33);
nand U1169 (N_1169,N_312,N_564);
or U1170 (N_1170,N_314,N_671);
and U1171 (N_1171,N_629,N_39);
nand U1172 (N_1172,N_266,N_530);
nor U1173 (N_1173,N_60,N_335);
xor U1174 (N_1174,N_448,N_599);
xnor U1175 (N_1175,N_581,N_389);
nand U1176 (N_1176,N_331,N_397);
nand U1177 (N_1177,N_326,N_557);
or U1178 (N_1178,N_50,N_306);
or U1179 (N_1179,N_403,N_650);
nor U1180 (N_1180,N_110,N_740);
and U1181 (N_1181,N_197,N_120);
nor U1182 (N_1182,N_235,N_635);
nor U1183 (N_1183,N_138,N_544);
xnor U1184 (N_1184,N_79,N_243);
and U1185 (N_1185,N_169,N_622);
nand U1186 (N_1186,N_128,N_361);
xnor U1187 (N_1187,N_544,N_478);
nor U1188 (N_1188,N_195,N_711);
or U1189 (N_1189,N_129,N_47);
xor U1190 (N_1190,N_400,N_687);
or U1191 (N_1191,N_149,N_323);
or U1192 (N_1192,N_199,N_735);
or U1193 (N_1193,N_712,N_671);
nand U1194 (N_1194,N_681,N_526);
xor U1195 (N_1195,N_552,N_696);
xnor U1196 (N_1196,N_138,N_693);
or U1197 (N_1197,N_570,N_610);
and U1198 (N_1198,N_190,N_35);
nand U1199 (N_1199,N_44,N_590);
xor U1200 (N_1200,N_42,N_292);
nand U1201 (N_1201,N_715,N_658);
xor U1202 (N_1202,N_626,N_571);
xor U1203 (N_1203,N_238,N_370);
and U1204 (N_1204,N_120,N_184);
or U1205 (N_1205,N_481,N_558);
and U1206 (N_1206,N_271,N_358);
nor U1207 (N_1207,N_737,N_417);
xnor U1208 (N_1208,N_90,N_34);
or U1209 (N_1209,N_42,N_228);
or U1210 (N_1210,N_715,N_468);
nor U1211 (N_1211,N_261,N_130);
xor U1212 (N_1212,N_33,N_283);
nor U1213 (N_1213,N_411,N_315);
xor U1214 (N_1214,N_27,N_111);
or U1215 (N_1215,N_137,N_492);
xor U1216 (N_1216,N_356,N_532);
xor U1217 (N_1217,N_179,N_220);
or U1218 (N_1218,N_13,N_467);
or U1219 (N_1219,N_362,N_232);
xor U1220 (N_1220,N_416,N_668);
nand U1221 (N_1221,N_264,N_709);
nor U1222 (N_1222,N_550,N_4);
nand U1223 (N_1223,N_303,N_313);
or U1224 (N_1224,N_683,N_111);
xor U1225 (N_1225,N_169,N_240);
xnor U1226 (N_1226,N_559,N_93);
or U1227 (N_1227,N_23,N_403);
and U1228 (N_1228,N_117,N_506);
and U1229 (N_1229,N_587,N_352);
nor U1230 (N_1230,N_167,N_101);
and U1231 (N_1231,N_61,N_321);
nand U1232 (N_1232,N_271,N_554);
nand U1233 (N_1233,N_616,N_186);
and U1234 (N_1234,N_697,N_301);
and U1235 (N_1235,N_443,N_100);
nor U1236 (N_1236,N_708,N_474);
xor U1237 (N_1237,N_382,N_674);
nor U1238 (N_1238,N_372,N_507);
nand U1239 (N_1239,N_211,N_689);
and U1240 (N_1240,N_584,N_21);
xor U1241 (N_1241,N_264,N_419);
nand U1242 (N_1242,N_516,N_481);
nand U1243 (N_1243,N_53,N_699);
or U1244 (N_1244,N_249,N_55);
and U1245 (N_1245,N_236,N_155);
or U1246 (N_1246,N_285,N_178);
and U1247 (N_1247,N_720,N_276);
and U1248 (N_1248,N_110,N_663);
nor U1249 (N_1249,N_214,N_326);
xnor U1250 (N_1250,N_598,N_520);
nor U1251 (N_1251,N_660,N_676);
xnor U1252 (N_1252,N_684,N_673);
and U1253 (N_1253,N_415,N_558);
and U1254 (N_1254,N_0,N_129);
nand U1255 (N_1255,N_187,N_667);
and U1256 (N_1256,N_285,N_460);
nand U1257 (N_1257,N_700,N_192);
nor U1258 (N_1258,N_404,N_45);
or U1259 (N_1259,N_199,N_637);
or U1260 (N_1260,N_14,N_413);
xnor U1261 (N_1261,N_165,N_336);
or U1262 (N_1262,N_256,N_162);
or U1263 (N_1263,N_42,N_582);
nor U1264 (N_1264,N_354,N_223);
and U1265 (N_1265,N_423,N_653);
and U1266 (N_1266,N_2,N_306);
nor U1267 (N_1267,N_98,N_466);
xor U1268 (N_1268,N_692,N_46);
and U1269 (N_1269,N_574,N_326);
and U1270 (N_1270,N_18,N_353);
or U1271 (N_1271,N_552,N_205);
nand U1272 (N_1272,N_128,N_317);
or U1273 (N_1273,N_554,N_16);
xnor U1274 (N_1274,N_722,N_352);
nor U1275 (N_1275,N_267,N_262);
nor U1276 (N_1276,N_614,N_168);
xor U1277 (N_1277,N_14,N_701);
nor U1278 (N_1278,N_116,N_686);
nor U1279 (N_1279,N_173,N_260);
nor U1280 (N_1280,N_173,N_662);
and U1281 (N_1281,N_264,N_676);
and U1282 (N_1282,N_331,N_684);
or U1283 (N_1283,N_341,N_196);
nor U1284 (N_1284,N_617,N_707);
and U1285 (N_1285,N_478,N_572);
and U1286 (N_1286,N_517,N_568);
and U1287 (N_1287,N_363,N_748);
xnor U1288 (N_1288,N_613,N_27);
and U1289 (N_1289,N_490,N_746);
xnor U1290 (N_1290,N_153,N_337);
and U1291 (N_1291,N_684,N_259);
nand U1292 (N_1292,N_261,N_413);
or U1293 (N_1293,N_29,N_595);
nand U1294 (N_1294,N_85,N_710);
and U1295 (N_1295,N_288,N_654);
nand U1296 (N_1296,N_558,N_731);
nand U1297 (N_1297,N_454,N_624);
nand U1298 (N_1298,N_611,N_8);
or U1299 (N_1299,N_68,N_722);
xor U1300 (N_1300,N_423,N_161);
and U1301 (N_1301,N_305,N_201);
xor U1302 (N_1302,N_482,N_419);
and U1303 (N_1303,N_170,N_27);
xor U1304 (N_1304,N_502,N_497);
xor U1305 (N_1305,N_617,N_310);
and U1306 (N_1306,N_0,N_400);
or U1307 (N_1307,N_163,N_277);
or U1308 (N_1308,N_687,N_311);
or U1309 (N_1309,N_258,N_374);
and U1310 (N_1310,N_271,N_627);
nor U1311 (N_1311,N_348,N_266);
and U1312 (N_1312,N_520,N_116);
and U1313 (N_1313,N_48,N_62);
nor U1314 (N_1314,N_245,N_469);
xnor U1315 (N_1315,N_635,N_618);
xor U1316 (N_1316,N_123,N_372);
nand U1317 (N_1317,N_333,N_129);
nor U1318 (N_1318,N_662,N_54);
nor U1319 (N_1319,N_201,N_262);
nand U1320 (N_1320,N_639,N_451);
nor U1321 (N_1321,N_195,N_5);
nor U1322 (N_1322,N_452,N_499);
and U1323 (N_1323,N_148,N_649);
xnor U1324 (N_1324,N_168,N_480);
and U1325 (N_1325,N_65,N_362);
xor U1326 (N_1326,N_356,N_362);
and U1327 (N_1327,N_357,N_61);
nor U1328 (N_1328,N_612,N_242);
or U1329 (N_1329,N_640,N_673);
or U1330 (N_1330,N_661,N_572);
nand U1331 (N_1331,N_35,N_352);
nor U1332 (N_1332,N_495,N_324);
xor U1333 (N_1333,N_474,N_498);
nand U1334 (N_1334,N_118,N_702);
or U1335 (N_1335,N_564,N_18);
nand U1336 (N_1336,N_706,N_537);
or U1337 (N_1337,N_492,N_684);
or U1338 (N_1338,N_72,N_590);
nand U1339 (N_1339,N_126,N_499);
nand U1340 (N_1340,N_78,N_480);
xnor U1341 (N_1341,N_28,N_41);
or U1342 (N_1342,N_369,N_75);
nor U1343 (N_1343,N_243,N_214);
xnor U1344 (N_1344,N_302,N_636);
nor U1345 (N_1345,N_192,N_379);
and U1346 (N_1346,N_238,N_619);
nand U1347 (N_1347,N_75,N_204);
xnor U1348 (N_1348,N_647,N_731);
nor U1349 (N_1349,N_137,N_372);
nor U1350 (N_1350,N_511,N_700);
nand U1351 (N_1351,N_516,N_219);
or U1352 (N_1352,N_175,N_555);
and U1353 (N_1353,N_313,N_575);
xnor U1354 (N_1354,N_695,N_226);
nand U1355 (N_1355,N_594,N_229);
nor U1356 (N_1356,N_665,N_13);
and U1357 (N_1357,N_126,N_721);
and U1358 (N_1358,N_216,N_705);
nor U1359 (N_1359,N_614,N_451);
nand U1360 (N_1360,N_369,N_42);
and U1361 (N_1361,N_636,N_255);
nand U1362 (N_1362,N_310,N_367);
and U1363 (N_1363,N_274,N_605);
and U1364 (N_1364,N_667,N_497);
or U1365 (N_1365,N_31,N_638);
xor U1366 (N_1366,N_652,N_103);
or U1367 (N_1367,N_155,N_352);
or U1368 (N_1368,N_215,N_485);
or U1369 (N_1369,N_438,N_88);
nor U1370 (N_1370,N_212,N_463);
nor U1371 (N_1371,N_583,N_169);
or U1372 (N_1372,N_416,N_148);
and U1373 (N_1373,N_152,N_519);
and U1374 (N_1374,N_353,N_540);
nor U1375 (N_1375,N_359,N_319);
and U1376 (N_1376,N_464,N_192);
or U1377 (N_1377,N_463,N_355);
or U1378 (N_1378,N_665,N_205);
and U1379 (N_1379,N_283,N_7);
and U1380 (N_1380,N_375,N_206);
nand U1381 (N_1381,N_475,N_313);
and U1382 (N_1382,N_367,N_320);
or U1383 (N_1383,N_596,N_27);
nor U1384 (N_1384,N_414,N_287);
and U1385 (N_1385,N_207,N_741);
xor U1386 (N_1386,N_415,N_583);
nor U1387 (N_1387,N_187,N_639);
nand U1388 (N_1388,N_696,N_632);
xnor U1389 (N_1389,N_649,N_743);
nor U1390 (N_1390,N_410,N_537);
xnor U1391 (N_1391,N_547,N_325);
and U1392 (N_1392,N_632,N_594);
or U1393 (N_1393,N_545,N_152);
nor U1394 (N_1394,N_14,N_488);
xor U1395 (N_1395,N_403,N_277);
nor U1396 (N_1396,N_209,N_621);
nor U1397 (N_1397,N_168,N_529);
nand U1398 (N_1398,N_666,N_93);
nor U1399 (N_1399,N_442,N_151);
nor U1400 (N_1400,N_544,N_296);
nor U1401 (N_1401,N_457,N_325);
and U1402 (N_1402,N_360,N_680);
and U1403 (N_1403,N_22,N_716);
and U1404 (N_1404,N_96,N_402);
xor U1405 (N_1405,N_544,N_379);
and U1406 (N_1406,N_632,N_441);
nand U1407 (N_1407,N_368,N_287);
and U1408 (N_1408,N_25,N_579);
nand U1409 (N_1409,N_332,N_746);
and U1410 (N_1410,N_25,N_269);
and U1411 (N_1411,N_13,N_253);
or U1412 (N_1412,N_87,N_646);
nand U1413 (N_1413,N_695,N_227);
and U1414 (N_1414,N_306,N_685);
nor U1415 (N_1415,N_309,N_407);
nand U1416 (N_1416,N_571,N_113);
and U1417 (N_1417,N_548,N_699);
nor U1418 (N_1418,N_128,N_699);
and U1419 (N_1419,N_352,N_744);
nor U1420 (N_1420,N_188,N_623);
and U1421 (N_1421,N_716,N_610);
xor U1422 (N_1422,N_9,N_56);
nand U1423 (N_1423,N_262,N_97);
or U1424 (N_1424,N_163,N_186);
or U1425 (N_1425,N_367,N_471);
nand U1426 (N_1426,N_398,N_128);
and U1427 (N_1427,N_655,N_540);
nand U1428 (N_1428,N_608,N_134);
xnor U1429 (N_1429,N_197,N_290);
or U1430 (N_1430,N_325,N_535);
or U1431 (N_1431,N_568,N_573);
nand U1432 (N_1432,N_42,N_44);
or U1433 (N_1433,N_743,N_577);
nor U1434 (N_1434,N_521,N_702);
or U1435 (N_1435,N_533,N_476);
and U1436 (N_1436,N_650,N_188);
or U1437 (N_1437,N_460,N_528);
and U1438 (N_1438,N_148,N_413);
and U1439 (N_1439,N_70,N_24);
xnor U1440 (N_1440,N_221,N_196);
nand U1441 (N_1441,N_503,N_328);
nand U1442 (N_1442,N_209,N_368);
and U1443 (N_1443,N_679,N_91);
nor U1444 (N_1444,N_169,N_519);
or U1445 (N_1445,N_414,N_320);
nand U1446 (N_1446,N_251,N_192);
or U1447 (N_1447,N_223,N_106);
nand U1448 (N_1448,N_706,N_387);
and U1449 (N_1449,N_368,N_162);
xor U1450 (N_1450,N_742,N_517);
or U1451 (N_1451,N_389,N_223);
nor U1452 (N_1452,N_86,N_221);
nor U1453 (N_1453,N_40,N_520);
nand U1454 (N_1454,N_391,N_360);
or U1455 (N_1455,N_192,N_518);
nand U1456 (N_1456,N_636,N_699);
or U1457 (N_1457,N_639,N_293);
and U1458 (N_1458,N_741,N_38);
xnor U1459 (N_1459,N_567,N_308);
and U1460 (N_1460,N_656,N_268);
nor U1461 (N_1461,N_339,N_631);
xor U1462 (N_1462,N_566,N_719);
nand U1463 (N_1463,N_165,N_514);
and U1464 (N_1464,N_613,N_179);
or U1465 (N_1465,N_138,N_348);
nor U1466 (N_1466,N_456,N_682);
nor U1467 (N_1467,N_156,N_227);
or U1468 (N_1468,N_274,N_360);
nor U1469 (N_1469,N_580,N_398);
nor U1470 (N_1470,N_238,N_695);
and U1471 (N_1471,N_447,N_659);
nand U1472 (N_1472,N_421,N_249);
nor U1473 (N_1473,N_50,N_387);
xor U1474 (N_1474,N_111,N_505);
or U1475 (N_1475,N_188,N_470);
or U1476 (N_1476,N_436,N_275);
nand U1477 (N_1477,N_77,N_495);
xnor U1478 (N_1478,N_315,N_682);
and U1479 (N_1479,N_174,N_581);
nand U1480 (N_1480,N_472,N_2);
and U1481 (N_1481,N_704,N_251);
nand U1482 (N_1482,N_549,N_689);
xnor U1483 (N_1483,N_299,N_119);
and U1484 (N_1484,N_86,N_382);
xor U1485 (N_1485,N_552,N_2);
and U1486 (N_1486,N_578,N_566);
and U1487 (N_1487,N_628,N_86);
nand U1488 (N_1488,N_528,N_733);
nand U1489 (N_1489,N_396,N_14);
or U1490 (N_1490,N_131,N_75);
nand U1491 (N_1491,N_212,N_51);
nor U1492 (N_1492,N_328,N_618);
and U1493 (N_1493,N_493,N_626);
xor U1494 (N_1494,N_308,N_396);
nand U1495 (N_1495,N_277,N_179);
or U1496 (N_1496,N_472,N_156);
nor U1497 (N_1497,N_555,N_290);
and U1498 (N_1498,N_533,N_25);
and U1499 (N_1499,N_616,N_461);
nand U1500 (N_1500,N_1306,N_949);
or U1501 (N_1501,N_794,N_878);
xor U1502 (N_1502,N_1038,N_1226);
xnor U1503 (N_1503,N_1157,N_1060);
nand U1504 (N_1504,N_1327,N_1082);
nand U1505 (N_1505,N_1328,N_1249);
nand U1506 (N_1506,N_1359,N_779);
and U1507 (N_1507,N_1282,N_1325);
and U1508 (N_1508,N_1171,N_1378);
or U1509 (N_1509,N_1417,N_824);
xor U1510 (N_1510,N_813,N_1336);
xnor U1511 (N_1511,N_861,N_1224);
xor U1512 (N_1512,N_1341,N_1002);
or U1513 (N_1513,N_1207,N_1443);
or U1514 (N_1514,N_1009,N_1393);
nor U1515 (N_1515,N_1178,N_767);
nand U1516 (N_1516,N_800,N_1269);
and U1517 (N_1517,N_1143,N_935);
or U1518 (N_1518,N_914,N_1187);
nor U1519 (N_1519,N_1069,N_1026);
xnor U1520 (N_1520,N_835,N_934);
nand U1521 (N_1521,N_869,N_939);
and U1522 (N_1522,N_986,N_1040);
xor U1523 (N_1523,N_1240,N_1189);
nand U1524 (N_1524,N_1130,N_1270);
xnor U1525 (N_1525,N_816,N_1097);
or U1526 (N_1526,N_758,N_918);
or U1527 (N_1527,N_896,N_1441);
nor U1528 (N_1528,N_970,N_1313);
xnor U1529 (N_1529,N_1324,N_1430);
xor U1530 (N_1530,N_1016,N_1035);
nand U1531 (N_1531,N_1278,N_1440);
or U1532 (N_1532,N_1225,N_1010);
and U1533 (N_1533,N_1186,N_1155);
nor U1534 (N_1534,N_757,N_1455);
and U1535 (N_1535,N_1432,N_1316);
nand U1536 (N_1536,N_1364,N_1319);
or U1537 (N_1537,N_1006,N_1193);
nand U1538 (N_1538,N_762,N_852);
xor U1539 (N_1539,N_1073,N_985);
nor U1540 (N_1540,N_778,N_810);
and U1541 (N_1541,N_1416,N_1357);
and U1542 (N_1542,N_1499,N_1438);
xnor U1543 (N_1543,N_797,N_1236);
nand U1544 (N_1544,N_806,N_975);
and U1545 (N_1545,N_981,N_1492);
nor U1546 (N_1546,N_1351,N_1179);
xor U1547 (N_1547,N_1264,N_1201);
and U1548 (N_1548,N_876,N_781);
xnor U1549 (N_1549,N_1283,N_1445);
nand U1550 (N_1550,N_846,N_875);
or U1551 (N_1551,N_965,N_1217);
nand U1552 (N_1552,N_925,N_963);
nand U1553 (N_1553,N_972,N_1109);
and U1554 (N_1554,N_1389,N_1210);
nor U1555 (N_1555,N_1095,N_1106);
and U1556 (N_1556,N_1090,N_941);
nand U1557 (N_1557,N_1120,N_1052);
or U1558 (N_1558,N_1211,N_1202);
and U1559 (N_1559,N_1220,N_1277);
nand U1560 (N_1560,N_857,N_1025);
nand U1561 (N_1561,N_1453,N_1235);
xor U1562 (N_1562,N_1285,N_859);
nand U1563 (N_1563,N_1387,N_1358);
or U1564 (N_1564,N_1005,N_1159);
or U1565 (N_1565,N_988,N_793);
nand U1566 (N_1566,N_1122,N_1491);
and U1567 (N_1567,N_1253,N_1498);
and U1568 (N_1568,N_1185,N_1353);
and U1569 (N_1569,N_1294,N_1295);
and U1570 (N_1570,N_1071,N_1065);
nand U1571 (N_1571,N_1384,N_1369);
nand U1572 (N_1572,N_1054,N_979);
and U1573 (N_1573,N_1388,N_853);
or U1574 (N_1574,N_1134,N_1044);
nor U1575 (N_1575,N_1433,N_948);
nand U1576 (N_1576,N_1028,N_1053);
nor U1577 (N_1577,N_836,N_908);
or U1578 (N_1578,N_1032,N_1067);
xnor U1579 (N_1579,N_976,N_1156);
nand U1580 (N_1580,N_881,N_958);
nor U1581 (N_1581,N_1227,N_1470);
xor U1582 (N_1582,N_821,N_1251);
nand U1583 (N_1583,N_1007,N_1111);
and U1584 (N_1584,N_1472,N_913);
xnor U1585 (N_1585,N_791,N_769);
xnor U1586 (N_1586,N_1373,N_1399);
xor U1587 (N_1587,N_974,N_1160);
nand U1588 (N_1588,N_1061,N_1018);
nor U1589 (N_1589,N_1287,N_1165);
nor U1590 (N_1590,N_843,N_1129);
xnor U1591 (N_1591,N_1188,N_1466);
nor U1592 (N_1592,N_1123,N_885);
nand U1593 (N_1593,N_888,N_795);
and U1594 (N_1594,N_1383,N_1375);
or U1595 (N_1595,N_1233,N_1355);
or U1596 (N_1596,N_1459,N_1495);
and U1597 (N_1597,N_1460,N_1252);
nor U1598 (N_1598,N_1079,N_858);
nor U1599 (N_1599,N_1222,N_1480);
nor U1600 (N_1600,N_1213,N_1320);
nand U1601 (N_1601,N_840,N_865);
xnor U1602 (N_1602,N_833,N_1150);
and U1603 (N_1603,N_1381,N_774);
or U1604 (N_1604,N_1050,N_952);
xor U1605 (N_1605,N_1289,N_919);
nor U1606 (N_1606,N_1442,N_1288);
or U1607 (N_1607,N_1184,N_1036);
nand U1608 (N_1608,N_768,N_1333);
and U1609 (N_1609,N_1274,N_1405);
xor U1610 (N_1610,N_1011,N_1170);
and U1611 (N_1611,N_1221,N_1163);
nand U1612 (N_1612,N_780,N_1337);
xnor U1613 (N_1613,N_790,N_900);
or U1614 (N_1614,N_911,N_1477);
and U1615 (N_1615,N_1033,N_803);
nand U1616 (N_1616,N_1377,N_938);
nor U1617 (N_1617,N_1076,N_1382);
or U1618 (N_1618,N_937,N_867);
xnor U1619 (N_1619,N_1138,N_961);
xnor U1620 (N_1620,N_1250,N_964);
and U1621 (N_1621,N_871,N_1410);
and U1622 (N_1622,N_1142,N_812);
or U1623 (N_1623,N_856,N_1021);
nand U1624 (N_1624,N_1023,N_1194);
nand U1625 (N_1625,N_1401,N_1080);
or U1626 (N_1626,N_1198,N_1141);
and U1627 (N_1627,N_1027,N_923);
xnor U1628 (N_1628,N_1085,N_917);
nand U1629 (N_1629,N_870,N_826);
nor U1630 (N_1630,N_1116,N_1128);
nand U1631 (N_1631,N_1175,N_1368);
and U1632 (N_1632,N_834,N_1094);
or U1633 (N_1633,N_1427,N_788);
and U1634 (N_1634,N_825,N_1012);
or U1635 (N_1635,N_1411,N_924);
nand U1636 (N_1636,N_1110,N_851);
and U1637 (N_1637,N_1068,N_1041);
and U1638 (N_1638,N_1348,N_1371);
nand U1639 (N_1639,N_1243,N_1473);
xor U1640 (N_1640,N_1331,N_1279);
nand U1641 (N_1641,N_932,N_1314);
nand U1642 (N_1642,N_1101,N_1181);
and U1643 (N_1643,N_944,N_1494);
nand U1644 (N_1644,N_933,N_764);
or U1645 (N_1645,N_1267,N_1307);
nor U1646 (N_1646,N_987,N_1431);
or U1647 (N_1647,N_1055,N_1261);
nor U1648 (N_1648,N_804,N_860);
and U1649 (N_1649,N_882,N_844);
or U1650 (N_1650,N_1484,N_1029);
and U1651 (N_1651,N_761,N_922);
xor U1652 (N_1652,N_1063,N_902);
nand U1653 (N_1653,N_808,N_1424);
xor U1654 (N_1654,N_989,N_1390);
nor U1655 (N_1655,N_823,N_1303);
or U1656 (N_1656,N_980,N_1199);
nor U1657 (N_1657,N_893,N_1102);
and U1658 (N_1658,N_837,N_1272);
nor U1659 (N_1659,N_1468,N_905);
xnor U1660 (N_1660,N_1203,N_1229);
nor U1661 (N_1661,N_1449,N_1493);
xor U1662 (N_1662,N_760,N_832);
xor U1663 (N_1663,N_1144,N_880);
or U1664 (N_1664,N_771,N_1245);
or U1665 (N_1665,N_1342,N_1059);
or U1666 (N_1666,N_1121,N_1457);
or U1667 (N_1667,N_894,N_969);
xnor U1668 (N_1668,N_839,N_1452);
and U1669 (N_1669,N_1464,N_1174);
xor U1670 (N_1670,N_920,N_1276);
or U1671 (N_1671,N_959,N_877);
nor U1672 (N_1672,N_1093,N_954);
and U1673 (N_1673,N_814,N_1140);
and U1674 (N_1674,N_890,N_1088);
and U1675 (N_1675,N_968,N_910);
nand U1676 (N_1676,N_1496,N_1352);
xnor U1677 (N_1677,N_1164,N_1479);
nand U1678 (N_1678,N_929,N_1191);
nor U1679 (N_1679,N_1346,N_785);
or U1680 (N_1680,N_1022,N_786);
and U1681 (N_1681,N_830,N_864);
nor U1682 (N_1682,N_775,N_1379);
and U1683 (N_1683,N_966,N_1293);
or U1684 (N_1684,N_1074,N_1192);
nor U1685 (N_1685,N_1487,N_1467);
xor U1686 (N_1686,N_1273,N_784);
nor U1687 (N_1687,N_1209,N_1034);
or U1688 (N_1688,N_1374,N_1343);
nor U1689 (N_1689,N_1112,N_1152);
nor U1690 (N_1690,N_1125,N_909);
nand U1691 (N_1691,N_1380,N_1418);
nand U1692 (N_1692,N_1266,N_1402);
xor U1693 (N_1693,N_1363,N_841);
nor U1694 (N_1694,N_1081,N_1284);
or U1695 (N_1695,N_1204,N_1315);
and U1696 (N_1696,N_993,N_842);
and U1697 (N_1697,N_805,N_1301);
nor U1698 (N_1698,N_1451,N_1195);
or U1699 (N_1699,N_889,N_1231);
nand U1700 (N_1700,N_1237,N_1397);
and U1701 (N_1701,N_1429,N_1238);
or U1702 (N_1702,N_1183,N_1345);
and U1703 (N_1703,N_1197,N_1409);
nand U1704 (N_1704,N_1322,N_1326);
nand U1705 (N_1705,N_942,N_1344);
nor U1706 (N_1706,N_1066,N_1092);
and U1707 (N_1707,N_906,N_796);
or U1708 (N_1708,N_1078,N_1447);
xor U1709 (N_1709,N_754,N_1030);
xor U1710 (N_1710,N_1317,N_872);
nand U1711 (N_1711,N_1394,N_1395);
xnor U1712 (N_1712,N_1434,N_1304);
nor U1713 (N_1713,N_763,N_1362);
xnor U1714 (N_1714,N_1132,N_1015);
or U1715 (N_1715,N_1228,N_811);
xnor U1716 (N_1716,N_977,N_1001);
or U1717 (N_1717,N_829,N_1182);
xor U1718 (N_1718,N_1149,N_994);
and U1719 (N_1719,N_950,N_1070);
nor U1720 (N_1720,N_1039,N_1291);
nor U1721 (N_1721,N_1248,N_792);
and U1722 (N_1722,N_1077,N_854);
and U1723 (N_1723,N_1215,N_1139);
and U1724 (N_1724,N_1017,N_1321);
and U1725 (N_1725,N_1086,N_1113);
and U1726 (N_1726,N_1020,N_995);
or U1727 (N_1727,N_883,N_1478);
or U1728 (N_1728,N_1415,N_898);
xor U1729 (N_1729,N_1161,N_770);
nand U1730 (N_1730,N_789,N_1104);
or U1731 (N_1731,N_1296,N_849);
and U1732 (N_1732,N_1486,N_903);
and U1733 (N_1733,N_798,N_1465);
nand U1734 (N_1734,N_926,N_1099);
xnor U1735 (N_1735,N_931,N_1218);
or U1736 (N_1736,N_1075,N_1045);
nand U1737 (N_1737,N_1311,N_1490);
nand U1738 (N_1738,N_884,N_845);
xnor U1739 (N_1739,N_1043,N_1244);
and U1740 (N_1740,N_1419,N_1297);
nand U1741 (N_1741,N_1376,N_773);
nand U1742 (N_1742,N_1391,N_1392);
and U1743 (N_1743,N_1096,N_1425);
or U1744 (N_1744,N_822,N_992);
or U1745 (N_1745,N_1126,N_1356);
nor U1746 (N_1746,N_1281,N_1058);
nand U1747 (N_1747,N_1107,N_1089);
xnor U1748 (N_1748,N_755,N_1308);
nand U1749 (N_1749,N_887,N_886);
nand U1750 (N_1750,N_1151,N_1414);
xor U1751 (N_1751,N_1103,N_953);
nor U1752 (N_1752,N_1219,N_862);
nor U1753 (N_1753,N_1153,N_1214);
and U1754 (N_1754,N_1361,N_1051);
and U1755 (N_1755,N_1254,N_1312);
nand U1756 (N_1756,N_1256,N_936);
or U1757 (N_1757,N_1292,N_815);
nand U1758 (N_1758,N_1323,N_930);
nor U1759 (N_1759,N_751,N_1056);
or U1760 (N_1760,N_1257,N_1412);
xnor U1761 (N_1761,N_1408,N_1042);
and U1762 (N_1762,N_866,N_1386);
nor U1763 (N_1763,N_772,N_1259);
nand U1764 (N_1764,N_1108,N_973);
nand U1765 (N_1765,N_1309,N_1047);
xor U1766 (N_1766,N_907,N_1435);
nand U1767 (N_1767,N_1439,N_946);
xor U1768 (N_1768,N_783,N_1298);
nand U1769 (N_1769,N_1057,N_1019);
and U1770 (N_1770,N_1485,N_1008);
and U1771 (N_1771,N_895,N_1347);
and U1772 (N_1772,N_978,N_1114);
and U1773 (N_1773,N_1180,N_1048);
or U1774 (N_1774,N_1475,N_782);
and U1775 (N_1775,N_1354,N_904);
nor U1776 (N_1776,N_1413,N_1124);
nand U1777 (N_1777,N_1366,N_1131);
nand U1778 (N_1778,N_1426,N_1037);
nor U1779 (N_1779,N_892,N_756);
nand U1780 (N_1780,N_1208,N_1145);
xor U1781 (N_1781,N_991,N_801);
nand U1782 (N_1782,N_940,N_752);
nand U1783 (N_1783,N_1403,N_1474);
nor U1784 (N_1784,N_1133,N_1423);
nor U1785 (N_1785,N_1137,N_1158);
or U1786 (N_1786,N_1154,N_1476);
or U1787 (N_1787,N_809,N_818);
nor U1788 (N_1788,N_1406,N_1339);
xor U1789 (N_1789,N_1305,N_947);
and U1790 (N_1790,N_1360,N_990);
xor U1791 (N_1791,N_1446,N_1232);
xor U1792 (N_1792,N_1275,N_1448);
and U1793 (N_1793,N_957,N_971);
nand U1794 (N_1794,N_1462,N_1265);
nor U1795 (N_1795,N_999,N_1136);
xor U1796 (N_1796,N_1115,N_1013);
nand U1797 (N_1797,N_1335,N_868);
nand U1798 (N_1798,N_915,N_1200);
or U1799 (N_1799,N_945,N_750);
nor U1800 (N_1800,N_1168,N_777);
xor U1801 (N_1801,N_1064,N_1072);
or U1802 (N_1802,N_828,N_1330);
nand U1803 (N_1803,N_1444,N_807);
or U1804 (N_1804,N_916,N_799);
nor U1805 (N_1805,N_951,N_1046);
and U1806 (N_1806,N_1084,N_1385);
xor U1807 (N_1807,N_996,N_891);
xor U1808 (N_1808,N_1481,N_921);
and U1809 (N_1809,N_759,N_1091);
nor U1810 (N_1810,N_1169,N_899);
nor U1811 (N_1811,N_1290,N_1062);
and U1812 (N_1812,N_1083,N_827);
and U1813 (N_1813,N_765,N_1302);
nand U1814 (N_1814,N_1400,N_850);
nor U1815 (N_1815,N_847,N_956);
xor U1816 (N_1816,N_1398,N_962);
nand U1817 (N_1817,N_1280,N_1310);
nor U1818 (N_1818,N_879,N_831);
nor U1819 (N_1819,N_873,N_1334);
xnor U1820 (N_1820,N_1260,N_1230);
nand U1821 (N_1821,N_802,N_1404);
and U1822 (N_1822,N_1489,N_997);
or U1823 (N_1823,N_1100,N_1087);
xor U1824 (N_1824,N_1014,N_1190);
nor U1825 (N_1825,N_1271,N_1212);
xor U1826 (N_1826,N_1105,N_1483);
and U1827 (N_1827,N_1247,N_820);
and U1828 (N_1828,N_1118,N_1147);
and U1829 (N_1829,N_984,N_1205);
xor U1830 (N_1830,N_817,N_1003);
nand U1831 (N_1831,N_927,N_1223);
or U1832 (N_1832,N_1396,N_1318);
nor U1833 (N_1833,N_1482,N_1268);
nand U1834 (N_1834,N_776,N_1262);
or U1835 (N_1835,N_1436,N_863);
xnor U1836 (N_1836,N_955,N_912);
or U1837 (N_1837,N_1461,N_1299);
nand U1838 (N_1838,N_1177,N_874);
nand U1839 (N_1839,N_1255,N_1167);
or U1840 (N_1840,N_1216,N_1241);
or U1841 (N_1841,N_1365,N_897);
xnor U1842 (N_1842,N_1463,N_1497);
nor U1843 (N_1843,N_1367,N_982);
and U1844 (N_1844,N_819,N_1422);
and U1845 (N_1845,N_1458,N_1146);
and U1846 (N_1846,N_1372,N_1117);
or U1847 (N_1847,N_960,N_1234);
nor U1848 (N_1848,N_1421,N_1471);
or U1849 (N_1849,N_1332,N_1456);
xor U1850 (N_1850,N_1196,N_1428);
or U1851 (N_1851,N_1148,N_1246);
or U1852 (N_1852,N_848,N_1420);
or U1853 (N_1853,N_1206,N_1004);
or U1854 (N_1854,N_766,N_1127);
nor U1855 (N_1855,N_1242,N_1098);
xnor U1856 (N_1856,N_1407,N_1300);
xor U1857 (N_1857,N_1049,N_1258);
or U1858 (N_1858,N_1173,N_1469);
xnor U1859 (N_1859,N_1166,N_1286);
xor U1860 (N_1860,N_753,N_1370);
or U1861 (N_1861,N_1329,N_1000);
nor U1862 (N_1862,N_1350,N_1340);
xnor U1863 (N_1863,N_1263,N_943);
xor U1864 (N_1864,N_1239,N_1437);
and U1865 (N_1865,N_1454,N_1135);
and U1866 (N_1866,N_998,N_1172);
and U1867 (N_1867,N_1031,N_787);
nor U1868 (N_1868,N_1119,N_838);
xnor U1869 (N_1869,N_901,N_983);
and U1870 (N_1870,N_1338,N_1349);
xnor U1871 (N_1871,N_1488,N_855);
nand U1872 (N_1872,N_1024,N_1176);
and U1873 (N_1873,N_967,N_928);
nor U1874 (N_1874,N_1162,N_1450);
xor U1875 (N_1875,N_1231,N_931);
and U1876 (N_1876,N_881,N_1294);
or U1877 (N_1877,N_754,N_833);
or U1878 (N_1878,N_1226,N_1214);
or U1879 (N_1879,N_975,N_1284);
nor U1880 (N_1880,N_1316,N_1110);
nand U1881 (N_1881,N_928,N_1257);
and U1882 (N_1882,N_932,N_1261);
nor U1883 (N_1883,N_853,N_945);
or U1884 (N_1884,N_1176,N_1095);
xor U1885 (N_1885,N_975,N_768);
and U1886 (N_1886,N_842,N_1077);
and U1887 (N_1887,N_1111,N_1256);
and U1888 (N_1888,N_1102,N_1022);
nand U1889 (N_1889,N_856,N_1431);
and U1890 (N_1890,N_913,N_1297);
or U1891 (N_1891,N_775,N_855);
or U1892 (N_1892,N_1440,N_869);
and U1893 (N_1893,N_1077,N_986);
nor U1894 (N_1894,N_910,N_1338);
or U1895 (N_1895,N_1203,N_1039);
nand U1896 (N_1896,N_1156,N_896);
nand U1897 (N_1897,N_1119,N_965);
xor U1898 (N_1898,N_1280,N_822);
xor U1899 (N_1899,N_916,N_1070);
nand U1900 (N_1900,N_1026,N_1230);
xnor U1901 (N_1901,N_1481,N_1278);
or U1902 (N_1902,N_1377,N_1219);
and U1903 (N_1903,N_867,N_1071);
nand U1904 (N_1904,N_1025,N_1321);
or U1905 (N_1905,N_1057,N_1450);
and U1906 (N_1906,N_1343,N_1449);
xnor U1907 (N_1907,N_1469,N_1058);
xnor U1908 (N_1908,N_911,N_1110);
or U1909 (N_1909,N_943,N_1373);
and U1910 (N_1910,N_1031,N_1350);
and U1911 (N_1911,N_1030,N_1354);
and U1912 (N_1912,N_993,N_1203);
nor U1913 (N_1913,N_1260,N_999);
or U1914 (N_1914,N_775,N_875);
and U1915 (N_1915,N_867,N_1084);
xor U1916 (N_1916,N_1498,N_765);
nand U1917 (N_1917,N_1317,N_1188);
and U1918 (N_1918,N_1138,N_1291);
nor U1919 (N_1919,N_1430,N_784);
nor U1920 (N_1920,N_1222,N_1427);
and U1921 (N_1921,N_1170,N_1250);
and U1922 (N_1922,N_1400,N_817);
nor U1923 (N_1923,N_1493,N_758);
nand U1924 (N_1924,N_946,N_1101);
nor U1925 (N_1925,N_970,N_920);
and U1926 (N_1926,N_865,N_1198);
xnor U1927 (N_1927,N_1139,N_1055);
or U1928 (N_1928,N_1175,N_963);
nor U1929 (N_1929,N_845,N_1056);
nor U1930 (N_1930,N_1020,N_1106);
nor U1931 (N_1931,N_995,N_1474);
xor U1932 (N_1932,N_1222,N_1167);
xnor U1933 (N_1933,N_1347,N_1377);
xnor U1934 (N_1934,N_1185,N_1081);
nand U1935 (N_1935,N_918,N_1361);
nand U1936 (N_1936,N_1394,N_1213);
xnor U1937 (N_1937,N_1031,N_1223);
xnor U1938 (N_1938,N_983,N_1160);
or U1939 (N_1939,N_772,N_788);
xor U1940 (N_1940,N_753,N_817);
nand U1941 (N_1941,N_886,N_770);
xor U1942 (N_1942,N_1485,N_1123);
nor U1943 (N_1943,N_809,N_1409);
nand U1944 (N_1944,N_1394,N_1434);
nand U1945 (N_1945,N_1437,N_753);
or U1946 (N_1946,N_1127,N_1184);
xor U1947 (N_1947,N_1300,N_1101);
nand U1948 (N_1948,N_1377,N_857);
nand U1949 (N_1949,N_963,N_1442);
or U1950 (N_1950,N_1389,N_942);
xnor U1951 (N_1951,N_1027,N_753);
xor U1952 (N_1952,N_990,N_1135);
xnor U1953 (N_1953,N_1428,N_885);
nor U1954 (N_1954,N_1323,N_824);
and U1955 (N_1955,N_1308,N_750);
xor U1956 (N_1956,N_966,N_1481);
xor U1957 (N_1957,N_1318,N_1428);
nand U1958 (N_1958,N_1400,N_1196);
or U1959 (N_1959,N_905,N_876);
and U1960 (N_1960,N_1331,N_1016);
xor U1961 (N_1961,N_1421,N_1375);
xnor U1962 (N_1962,N_1133,N_925);
nor U1963 (N_1963,N_1428,N_1063);
nand U1964 (N_1964,N_1459,N_1370);
nand U1965 (N_1965,N_1096,N_1297);
and U1966 (N_1966,N_1101,N_1421);
or U1967 (N_1967,N_902,N_1200);
or U1968 (N_1968,N_1379,N_908);
xnor U1969 (N_1969,N_793,N_1337);
and U1970 (N_1970,N_1242,N_1195);
nor U1971 (N_1971,N_1221,N_802);
nor U1972 (N_1972,N_1288,N_1460);
nor U1973 (N_1973,N_1487,N_972);
and U1974 (N_1974,N_1472,N_1104);
and U1975 (N_1975,N_1168,N_828);
nand U1976 (N_1976,N_1091,N_905);
and U1977 (N_1977,N_1142,N_1167);
nand U1978 (N_1978,N_1217,N_819);
xnor U1979 (N_1979,N_960,N_1457);
and U1980 (N_1980,N_1407,N_779);
or U1981 (N_1981,N_1364,N_1471);
nand U1982 (N_1982,N_1413,N_860);
nand U1983 (N_1983,N_1341,N_1489);
nand U1984 (N_1984,N_922,N_1303);
xor U1985 (N_1985,N_1282,N_841);
xnor U1986 (N_1986,N_936,N_1349);
nor U1987 (N_1987,N_1314,N_1359);
nor U1988 (N_1988,N_882,N_1439);
nor U1989 (N_1989,N_1167,N_1088);
nor U1990 (N_1990,N_1072,N_758);
or U1991 (N_1991,N_764,N_942);
xnor U1992 (N_1992,N_1419,N_1457);
nor U1993 (N_1993,N_851,N_983);
nor U1994 (N_1994,N_1012,N_918);
or U1995 (N_1995,N_1254,N_815);
xnor U1996 (N_1996,N_1186,N_1101);
or U1997 (N_1997,N_1331,N_853);
nand U1998 (N_1998,N_873,N_823);
xor U1999 (N_1999,N_1435,N_1270);
nand U2000 (N_2000,N_1102,N_1337);
xnor U2001 (N_2001,N_1330,N_872);
nor U2002 (N_2002,N_1095,N_987);
xnor U2003 (N_2003,N_1308,N_1246);
nor U2004 (N_2004,N_1417,N_1467);
or U2005 (N_2005,N_999,N_1451);
and U2006 (N_2006,N_793,N_779);
xor U2007 (N_2007,N_1492,N_838);
nand U2008 (N_2008,N_1249,N_1446);
nand U2009 (N_2009,N_1298,N_1140);
and U2010 (N_2010,N_959,N_1074);
or U2011 (N_2011,N_1343,N_835);
nor U2012 (N_2012,N_1145,N_1487);
nor U2013 (N_2013,N_916,N_809);
or U2014 (N_2014,N_1172,N_1215);
nor U2015 (N_2015,N_913,N_1349);
and U2016 (N_2016,N_868,N_1300);
or U2017 (N_2017,N_1463,N_855);
and U2018 (N_2018,N_881,N_866);
and U2019 (N_2019,N_977,N_1495);
nand U2020 (N_2020,N_1316,N_840);
or U2021 (N_2021,N_1119,N_760);
or U2022 (N_2022,N_1172,N_1437);
xor U2023 (N_2023,N_1038,N_938);
or U2024 (N_2024,N_1343,N_760);
or U2025 (N_2025,N_771,N_1420);
or U2026 (N_2026,N_1192,N_838);
xnor U2027 (N_2027,N_956,N_1480);
nand U2028 (N_2028,N_848,N_1388);
xnor U2029 (N_2029,N_1062,N_1289);
or U2030 (N_2030,N_1410,N_1374);
nor U2031 (N_2031,N_766,N_1494);
and U2032 (N_2032,N_1158,N_1380);
nand U2033 (N_2033,N_781,N_1377);
nand U2034 (N_2034,N_1046,N_1405);
nand U2035 (N_2035,N_1074,N_913);
xnor U2036 (N_2036,N_781,N_1090);
and U2037 (N_2037,N_826,N_806);
nor U2038 (N_2038,N_1329,N_1006);
xnor U2039 (N_2039,N_935,N_1428);
nand U2040 (N_2040,N_1325,N_1341);
or U2041 (N_2041,N_1492,N_1225);
nand U2042 (N_2042,N_1227,N_1384);
or U2043 (N_2043,N_1449,N_1336);
and U2044 (N_2044,N_1437,N_1181);
or U2045 (N_2045,N_1205,N_1460);
or U2046 (N_2046,N_851,N_1033);
nor U2047 (N_2047,N_975,N_918);
or U2048 (N_2048,N_940,N_949);
and U2049 (N_2049,N_1405,N_1177);
xnor U2050 (N_2050,N_1200,N_1109);
nor U2051 (N_2051,N_857,N_1395);
nand U2052 (N_2052,N_1168,N_1485);
xnor U2053 (N_2053,N_784,N_1018);
and U2054 (N_2054,N_910,N_1235);
and U2055 (N_2055,N_1008,N_1171);
or U2056 (N_2056,N_976,N_1311);
and U2057 (N_2057,N_888,N_1375);
or U2058 (N_2058,N_1267,N_999);
and U2059 (N_2059,N_1086,N_1253);
and U2060 (N_2060,N_1377,N_924);
or U2061 (N_2061,N_1046,N_1053);
nand U2062 (N_2062,N_1485,N_1027);
nor U2063 (N_2063,N_905,N_1422);
and U2064 (N_2064,N_832,N_1210);
or U2065 (N_2065,N_1376,N_1250);
nand U2066 (N_2066,N_1201,N_1378);
or U2067 (N_2067,N_835,N_798);
nand U2068 (N_2068,N_967,N_1331);
nand U2069 (N_2069,N_915,N_1444);
and U2070 (N_2070,N_987,N_843);
or U2071 (N_2071,N_1304,N_1351);
and U2072 (N_2072,N_1379,N_1304);
nor U2073 (N_2073,N_1234,N_1431);
nand U2074 (N_2074,N_1395,N_1171);
or U2075 (N_2075,N_1118,N_1341);
xnor U2076 (N_2076,N_944,N_1234);
and U2077 (N_2077,N_1148,N_1168);
xor U2078 (N_2078,N_844,N_1173);
xor U2079 (N_2079,N_908,N_802);
or U2080 (N_2080,N_773,N_986);
nor U2081 (N_2081,N_1338,N_1204);
or U2082 (N_2082,N_1037,N_1110);
nand U2083 (N_2083,N_1211,N_778);
nand U2084 (N_2084,N_1026,N_1013);
xor U2085 (N_2085,N_805,N_925);
or U2086 (N_2086,N_1488,N_888);
and U2087 (N_2087,N_965,N_1403);
xnor U2088 (N_2088,N_1136,N_1412);
nand U2089 (N_2089,N_817,N_834);
nor U2090 (N_2090,N_1074,N_968);
nand U2091 (N_2091,N_774,N_1482);
nor U2092 (N_2092,N_1147,N_1013);
nor U2093 (N_2093,N_1033,N_1378);
nor U2094 (N_2094,N_1228,N_1472);
xnor U2095 (N_2095,N_1182,N_774);
and U2096 (N_2096,N_839,N_1171);
nor U2097 (N_2097,N_1002,N_1390);
nand U2098 (N_2098,N_1209,N_831);
xor U2099 (N_2099,N_1391,N_1336);
xnor U2100 (N_2100,N_1009,N_978);
nand U2101 (N_2101,N_772,N_1189);
nand U2102 (N_2102,N_772,N_1013);
xnor U2103 (N_2103,N_1166,N_1056);
or U2104 (N_2104,N_1055,N_966);
nor U2105 (N_2105,N_1367,N_1081);
nand U2106 (N_2106,N_1462,N_811);
xnor U2107 (N_2107,N_1345,N_870);
and U2108 (N_2108,N_1105,N_833);
or U2109 (N_2109,N_1216,N_1452);
or U2110 (N_2110,N_1437,N_1462);
or U2111 (N_2111,N_1345,N_1154);
nor U2112 (N_2112,N_1427,N_1430);
nand U2113 (N_2113,N_1110,N_1123);
or U2114 (N_2114,N_915,N_1220);
xnor U2115 (N_2115,N_1378,N_981);
xor U2116 (N_2116,N_929,N_764);
or U2117 (N_2117,N_1311,N_1472);
xor U2118 (N_2118,N_770,N_1284);
and U2119 (N_2119,N_1399,N_1204);
and U2120 (N_2120,N_904,N_1084);
or U2121 (N_2121,N_1475,N_836);
xor U2122 (N_2122,N_793,N_1341);
or U2123 (N_2123,N_1070,N_886);
nor U2124 (N_2124,N_1186,N_1260);
nand U2125 (N_2125,N_1362,N_1384);
nand U2126 (N_2126,N_1130,N_793);
nand U2127 (N_2127,N_815,N_1026);
and U2128 (N_2128,N_1415,N_942);
xor U2129 (N_2129,N_1055,N_1110);
and U2130 (N_2130,N_960,N_914);
xor U2131 (N_2131,N_1254,N_1034);
or U2132 (N_2132,N_1239,N_829);
xor U2133 (N_2133,N_1109,N_752);
and U2134 (N_2134,N_1483,N_951);
nor U2135 (N_2135,N_1305,N_1271);
and U2136 (N_2136,N_1360,N_1388);
xor U2137 (N_2137,N_1139,N_1448);
nand U2138 (N_2138,N_840,N_1359);
nor U2139 (N_2139,N_1096,N_1400);
nor U2140 (N_2140,N_878,N_1060);
nor U2141 (N_2141,N_824,N_1073);
nand U2142 (N_2142,N_832,N_1035);
xnor U2143 (N_2143,N_1462,N_1301);
nor U2144 (N_2144,N_789,N_1486);
or U2145 (N_2145,N_887,N_1284);
nor U2146 (N_2146,N_1413,N_1136);
nor U2147 (N_2147,N_1135,N_1223);
xor U2148 (N_2148,N_1411,N_950);
or U2149 (N_2149,N_1217,N_1246);
nand U2150 (N_2150,N_1303,N_1446);
xnor U2151 (N_2151,N_1029,N_985);
nor U2152 (N_2152,N_970,N_1410);
or U2153 (N_2153,N_1287,N_993);
or U2154 (N_2154,N_994,N_1477);
xnor U2155 (N_2155,N_1456,N_1047);
or U2156 (N_2156,N_929,N_834);
and U2157 (N_2157,N_1182,N_896);
xnor U2158 (N_2158,N_1070,N_1040);
or U2159 (N_2159,N_1058,N_952);
nor U2160 (N_2160,N_1441,N_1434);
or U2161 (N_2161,N_1170,N_1473);
xor U2162 (N_2162,N_1019,N_764);
nand U2163 (N_2163,N_966,N_954);
nor U2164 (N_2164,N_930,N_909);
xnor U2165 (N_2165,N_1444,N_1326);
nand U2166 (N_2166,N_872,N_1499);
nor U2167 (N_2167,N_1030,N_1280);
or U2168 (N_2168,N_1413,N_1197);
xnor U2169 (N_2169,N_1220,N_1311);
nand U2170 (N_2170,N_1044,N_1132);
xnor U2171 (N_2171,N_1206,N_1292);
xnor U2172 (N_2172,N_1293,N_1402);
nand U2173 (N_2173,N_1254,N_1259);
and U2174 (N_2174,N_1448,N_929);
or U2175 (N_2175,N_1092,N_1374);
and U2176 (N_2176,N_1324,N_852);
xnor U2177 (N_2177,N_956,N_1066);
xnor U2178 (N_2178,N_932,N_1093);
or U2179 (N_2179,N_1009,N_1451);
nor U2180 (N_2180,N_1320,N_1171);
and U2181 (N_2181,N_1270,N_894);
xnor U2182 (N_2182,N_956,N_991);
nor U2183 (N_2183,N_916,N_982);
nor U2184 (N_2184,N_887,N_926);
or U2185 (N_2185,N_1492,N_1489);
nand U2186 (N_2186,N_971,N_856);
or U2187 (N_2187,N_1258,N_873);
xor U2188 (N_2188,N_945,N_1111);
xor U2189 (N_2189,N_1374,N_855);
nand U2190 (N_2190,N_1320,N_966);
or U2191 (N_2191,N_1324,N_1486);
xnor U2192 (N_2192,N_752,N_1241);
nor U2193 (N_2193,N_1293,N_776);
or U2194 (N_2194,N_900,N_1085);
or U2195 (N_2195,N_1137,N_1291);
xor U2196 (N_2196,N_1475,N_1173);
and U2197 (N_2197,N_1011,N_876);
nor U2198 (N_2198,N_1459,N_948);
or U2199 (N_2199,N_1253,N_1337);
xnor U2200 (N_2200,N_811,N_878);
xor U2201 (N_2201,N_1049,N_1415);
and U2202 (N_2202,N_780,N_1278);
xor U2203 (N_2203,N_835,N_780);
and U2204 (N_2204,N_1308,N_1354);
xnor U2205 (N_2205,N_815,N_1311);
nand U2206 (N_2206,N_807,N_942);
xnor U2207 (N_2207,N_1486,N_1460);
and U2208 (N_2208,N_1422,N_830);
nand U2209 (N_2209,N_1067,N_1465);
or U2210 (N_2210,N_1237,N_994);
nor U2211 (N_2211,N_1497,N_1473);
xnor U2212 (N_2212,N_1195,N_1166);
and U2213 (N_2213,N_1300,N_821);
nand U2214 (N_2214,N_1375,N_1376);
xnor U2215 (N_2215,N_1380,N_1088);
xnor U2216 (N_2216,N_874,N_1466);
nand U2217 (N_2217,N_1065,N_1444);
and U2218 (N_2218,N_1453,N_765);
and U2219 (N_2219,N_842,N_1216);
and U2220 (N_2220,N_1031,N_1224);
xor U2221 (N_2221,N_917,N_1099);
and U2222 (N_2222,N_1437,N_1496);
xnor U2223 (N_2223,N_1437,N_1488);
nor U2224 (N_2224,N_1494,N_848);
nor U2225 (N_2225,N_1346,N_927);
xor U2226 (N_2226,N_973,N_1154);
nand U2227 (N_2227,N_1034,N_1372);
or U2228 (N_2228,N_803,N_1391);
and U2229 (N_2229,N_753,N_1234);
or U2230 (N_2230,N_1194,N_844);
and U2231 (N_2231,N_972,N_827);
xor U2232 (N_2232,N_760,N_1007);
nor U2233 (N_2233,N_1058,N_1149);
and U2234 (N_2234,N_1233,N_1010);
and U2235 (N_2235,N_868,N_1140);
xnor U2236 (N_2236,N_1122,N_1105);
xnor U2237 (N_2237,N_1289,N_1034);
and U2238 (N_2238,N_900,N_810);
and U2239 (N_2239,N_1483,N_1007);
xnor U2240 (N_2240,N_1401,N_1222);
or U2241 (N_2241,N_1208,N_910);
and U2242 (N_2242,N_851,N_751);
and U2243 (N_2243,N_1054,N_1036);
xor U2244 (N_2244,N_957,N_852);
or U2245 (N_2245,N_907,N_1084);
xnor U2246 (N_2246,N_832,N_1119);
xor U2247 (N_2247,N_909,N_1497);
nor U2248 (N_2248,N_940,N_936);
nand U2249 (N_2249,N_1052,N_885);
xor U2250 (N_2250,N_2003,N_1502);
or U2251 (N_2251,N_1570,N_1959);
nor U2252 (N_2252,N_1557,N_2036);
nor U2253 (N_2253,N_1800,N_2122);
nor U2254 (N_2254,N_2111,N_1897);
or U2255 (N_2255,N_1874,N_1504);
nor U2256 (N_2256,N_1979,N_1653);
nor U2257 (N_2257,N_2053,N_2045);
or U2258 (N_2258,N_1957,N_2178);
nand U2259 (N_2259,N_1531,N_1796);
nor U2260 (N_2260,N_1672,N_2205);
nand U2261 (N_2261,N_1581,N_1890);
or U2262 (N_2262,N_1788,N_1543);
xnor U2263 (N_2263,N_1555,N_2177);
xnor U2264 (N_2264,N_1759,N_1750);
xnor U2265 (N_2265,N_2030,N_2162);
nor U2266 (N_2266,N_1941,N_1930);
nor U2267 (N_2267,N_1921,N_1873);
xnor U2268 (N_2268,N_1772,N_1815);
and U2269 (N_2269,N_1970,N_2040);
xnor U2270 (N_2270,N_2147,N_1647);
nor U2271 (N_2271,N_2039,N_1735);
or U2272 (N_2272,N_2057,N_1836);
or U2273 (N_2273,N_1592,N_1822);
nor U2274 (N_2274,N_2038,N_1567);
or U2275 (N_2275,N_1881,N_1980);
nor U2276 (N_2276,N_1547,N_1820);
or U2277 (N_2277,N_1965,N_1660);
nand U2278 (N_2278,N_1550,N_1834);
nor U2279 (N_2279,N_2224,N_1829);
and U2280 (N_2280,N_2145,N_1875);
or U2281 (N_2281,N_2107,N_2082);
nand U2282 (N_2282,N_2026,N_2071);
nor U2283 (N_2283,N_1774,N_1801);
xor U2284 (N_2284,N_1743,N_2059);
xnor U2285 (N_2285,N_1642,N_2133);
nand U2286 (N_2286,N_1527,N_2020);
and U2287 (N_2287,N_1992,N_2117);
nand U2288 (N_2288,N_2091,N_1898);
and U2289 (N_2289,N_1655,N_1731);
xnor U2290 (N_2290,N_1817,N_2019);
nand U2291 (N_2291,N_2226,N_2033);
and U2292 (N_2292,N_1943,N_2000);
nor U2293 (N_2293,N_1797,N_1638);
or U2294 (N_2294,N_1689,N_1804);
and U2295 (N_2295,N_2044,N_1784);
or U2296 (N_2296,N_2096,N_1937);
xnor U2297 (N_2297,N_1508,N_2175);
xnor U2298 (N_2298,N_2217,N_1831);
nor U2299 (N_2299,N_1597,N_2208);
and U2300 (N_2300,N_2001,N_2151);
or U2301 (N_2301,N_1764,N_2153);
and U2302 (N_2302,N_1969,N_1859);
xor U2303 (N_2303,N_1795,N_1863);
or U2304 (N_2304,N_2154,N_2123);
xnor U2305 (N_2305,N_1556,N_1753);
nand U2306 (N_2306,N_1621,N_1549);
nor U2307 (N_2307,N_1974,N_1725);
nor U2308 (N_2308,N_1560,N_1553);
xor U2309 (N_2309,N_1563,N_2021);
or U2310 (N_2310,N_2027,N_1682);
xor U2311 (N_2311,N_2167,N_1646);
and U2312 (N_2312,N_2090,N_2109);
nand U2313 (N_2313,N_2120,N_1628);
and U2314 (N_2314,N_2190,N_1610);
or U2315 (N_2315,N_1926,N_1516);
or U2316 (N_2316,N_1712,N_2223);
nand U2317 (N_2317,N_2163,N_1929);
and U2318 (N_2318,N_1634,N_2118);
or U2319 (N_2319,N_2068,N_1709);
and U2320 (N_2320,N_2236,N_1860);
nor U2321 (N_2321,N_1645,N_1765);
or U2322 (N_2322,N_2203,N_2046);
nand U2323 (N_2323,N_1896,N_2127);
and U2324 (N_2324,N_2067,N_1838);
or U2325 (N_2325,N_2006,N_2070);
nand U2326 (N_2326,N_2084,N_1568);
xnor U2327 (N_2327,N_2164,N_1825);
and U2328 (N_2328,N_1826,N_2211);
and U2329 (N_2329,N_1640,N_1604);
nor U2330 (N_2330,N_1912,N_1678);
and U2331 (N_2331,N_1942,N_1850);
and U2332 (N_2332,N_1691,N_1887);
xnor U2333 (N_2333,N_1751,N_2138);
nand U2334 (N_2334,N_1903,N_2139);
and U2335 (N_2335,N_1602,N_1952);
nor U2336 (N_2336,N_1947,N_2061);
xor U2337 (N_2337,N_1893,N_1662);
nor U2338 (N_2338,N_1687,N_1683);
nand U2339 (N_2339,N_1579,N_1586);
nor U2340 (N_2340,N_1847,N_1832);
nand U2341 (N_2341,N_1548,N_1532);
and U2342 (N_2342,N_2014,N_1744);
xor U2343 (N_2343,N_1705,N_1999);
xnor U2344 (N_2344,N_2102,N_2028);
and U2345 (N_2345,N_2227,N_1669);
nor U2346 (N_2346,N_1981,N_1629);
or U2347 (N_2347,N_1790,N_1639);
xor U2348 (N_2348,N_2064,N_1830);
nand U2349 (N_2349,N_1697,N_1685);
xnor U2350 (N_2350,N_1644,N_2148);
xor U2351 (N_2351,N_1840,N_1781);
xor U2352 (N_2352,N_2069,N_2160);
or U2353 (N_2353,N_1916,N_1564);
nand U2354 (N_2354,N_1986,N_1914);
xnor U2355 (N_2355,N_1762,N_2170);
or U2356 (N_2356,N_1983,N_1613);
xor U2357 (N_2357,N_1728,N_2169);
xor U2358 (N_2358,N_1814,N_1741);
nand U2359 (N_2359,N_1919,N_2158);
xnor U2360 (N_2360,N_1805,N_1583);
and U2361 (N_2361,N_1913,N_2018);
nor U2362 (N_2362,N_1944,N_2043);
and U2363 (N_2363,N_2140,N_1618);
xor U2364 (N_2364,N_1552,N_2193);
or U2365 (N_2365,N_2008,N_1542);
nor U2366 (N_2366,N_1673,N_1908);
and U2367 (N_2367,N_1745,N_2197);
nor U2368 (N_2368,N_1871,N_1701);
nand U2369 (N_2369,N_1739,N_1747);
nand U2370 (N_2370,N_1839,N_1848);
nand U2371 (N_2371,N_1761,N_1779);
xor U2372 (N_2372,N_2136,N_1513);
or U2373 (N_2373,N_1541,N_2143);
or U2374 (N_2374,N_2029,N_1982);
and U2375 (N_2375,N_1575,N_1708);
or U2376 (N_2376,N_1948,N_1870);
nand U2377 (N_2377,N_1902,N_1730);
xor U2378 (N_2378,N_2023,N_2228);
xor U2379 (N_2379,N_1540,N_1650);
or U2380 (N_2380,N_2050,N_1923);
nand U2381 (N_2381,N_2249,N_1591);
nor U2382 (N_2382,N_1828,N_1522);
or U2383 (N_2383,N_2168,N_1842);
xor U2384 (N_2384,N_1869,N_1978);
and U2385 (N_2385,N_1837,N_1659);
xnor U2386 (N_2386,N_2213,N_1595);
and U2387 (N_2387,N_1934,N_2076);
xnor U2388 (N_2388,N_1975,N_1577);
nor U2389 (N_2389,N_2088,N_1671);
nand U2390 (N_2390,N_1713,N_2222);
xor U2391 (N_2391,N_1811,N_1688);
nand U2392 (N_2392,N_1964,N_1818);
and U2393 (N_2393,N_1856,N_2199);
nor U2394 (N_2394,N_2002,N_1611);
xor U2395 (N_2395,N_1539,N_1971);
or U2396 (N_2396,N_1715,N_2083);
nor U2397 (N_2397,N_2013,N_1958);
and U2398 (N_2398,N_1833,N_1885);
nand U2399 (N_2399,N_1989,N_1773);
xnor U2400 (N_2400,N_1698,N_2207);
or U2401 (N_2401,N_2142,N_1661);
nor U2402 (N_2402,N_1538,N_1729);
or U2403 (N_2403,N_1905,N_2244);
and U2404 (N_2404,N_1864,N_2051);
nor U2405 (N_2405,N_1955,N_1872);
xnor U2406 (N_2406,N_1658,N_1968);
nand U2407 (N_2407,N_2238,N_1505);
and U2408 (N_2408,N_2128,N_2218);
xnor U2409 (N_2409,N_1737,N_2233);
or U2410 (N_2410,N_1529,N_1588);
or U2411 (N_2411,N_2055,N_1571);
nor U2412 (N_2412,N_2230,N_1598);
xnor U2413 (N_2413,N_1802,N_1614);
or U2414 (N_2414,N_2184,N_1748);
xnor U2415 (N_2415,N_2105,N_1714);
and U2416 (N_2416,N_1584,N_2056);
nor U2417 (N_2417,N_2119,N_1631);
xnor U2418 (N_2418,N_2048,N_1736);
or U2419 (N_2419,N_2210,N_1996);
nor U2420 (N_2420,N_1951,N_1738);
and U2421 (N_2421,N_2146,N_2195);
nand U2422 (N_2422,N_1726,N_1991);
nor U2423 (N_2423,N_2156,N_1782);
xor U2424 (N_2424,N_1630,N_2200);
nand U2425 (N_2425,N_2165,N_1694);
or U2426 (N_2426,N_1813,N_1945);
and U2427 (N_2427,N_1703,N_1977);
nor U2428 (N_2428,N_2075,N_1665);
and U2429 (N_2429,N_2103,N_1973);
nor U2430 (N_2430,N_1733,N_1793);
or U2431 (N_2431,N_2094,N_1904);
and U2432 (N_2432,N_2074,N_1976);
and U2433 (N_2433,N_1767,N_1998);
and U2434 (N_2434,N_1648,N_2034);
nand U2435 (N_2435,N_1972,N_1500);
nor U2436 (N_2436,N_1928,N_2234);
xor U2437 (N_2437,N_1954,N_1769);
xor U2438 (N_2438,N_1511,N_1878);
and U2439 (N_2439,N_1789,N_1867);
or U2440 (N_2440,N_2248,N_2087);
nand U2441 (N_2441,N_2089,N_1809);
and U2442 (N_2442,N_1894,N_1615);
xor U2443 (N_2443,N_1530,N_1651);
and U2444 (N_2444,N_1684,N_1843);
and U2445 (N_2445,N_1721,N_1918);
xnor U2446 (N_2446,N_1900,N_2012);
nor U2447 (N_2447,N_2035,N_1754);
nand U2448 (N_2448,N_2085,N_2204);
or U2449 (N_2449,N_1559,N_1760);
nand U2450 (N_2450,N_1879,N_2010);
and U2451 (N_2451,N_2132,N_1590);
xnor U2452 (N_2452,N_1578,N_2202);
xor U2453 (N_2453,N_1718,N_2191);
nand U2454 (N_2454,N_1625,N_1676);
xnor U2455 (N_2455,N_2209,N_2183);
nand U2456 (N_2456,N_1938,N_1852);
or U2457 (N_2457,N_1605,N_2106);
nand U2458 (N_2458,N_1990,N_2081);
or U2459 (N_2459,N_2116,N_2135);
and U2460 (N_2460,N_2172,N_1536);
nand U2461 (N_2461,N_1775,N_2242);
nor U2462 (N_2462,N_2189,N_1886);
and U2463 (N_2463,N_1791,N_1911);
and U2464 (N_2464,N_1824,N_1596);
and U2465 (N_2465,N_1798,N_2031);
xor U2466 (N_2466,N_1554,N_1656);
nor U2467 (N_2467,N_2159,N_2221);
xnor U2468 (N_2468,N_1692,N_1637);
nor U2469 (N_2469,N_1925,N_2131);
or U2470 (N_2470,N_1643,N_1704);
or U2471 (N_2471,N_1868,N_2141);
nand U2472 (N_2472,N_2115,N_2231);
or U2473 (N_2473,N_1915,N_1967);
and U2474 (N_2474,N_1717,N_1517);
nor U2475 (N_2475,N_1888,N_2182);
or U2476 (N_2476,N_2171,N_2144);
xor U2477 (N_2477,N_1742,N_1846);
nor U2478 (N_2478,N_2093,N_2016);
or U2479 (N_2479,N_1757,N_1649);
xnor U2480 (N_2480,N_2110,N_1624);
xnor U2481 (N_2481,N_1922,N_2086);
and U2482 (N_2482,N_2179,N_1880);
nand U2483 (N_2483,N_2157,N_1652);
nand U2484 (N_2484,N_2247,N_2196);
and U2485 (N_2485,N_1949,N_1528);
and U2486 (N_2486,N_2240,N_2077);
and U2487 (N_2487,N_1695,N_1960);
or U2488 (N_2488,N_1786,N_1901);
xor U2489 (N_2489,N_2166,N_1675);
or U2490 (N_2490,N_2011,N_1699);
or U2491 (N_2491,N_1994,N_1654);
or U2492 (N_2492,N_2101,N_1783);
or U2493 (N_2493,N_1616,N_1962);
xor U2494 (N_2494,N_2235,N_1768);
and U2495 (N_2495,N_1844,N_1876);
or U2496 (N_2496,N_2125,N_2097);
and U2497 (N_2497,N_1756,N_1865);
xnor U2498 (N_2498,N_1627,N_1924);
nor U2499 (N_2499,N_1580,N_1907);
or U2500 (N_2500,N_2073,N_1633);
nand U2501 (N_2501,N_2150,N_2079);
nand U2502 (N_2502,N_1622,N_1574);
and U2503 (N_2503,N_2032,N_2134);
xor U2504 (N_2504,N_2206,N_1988);
and U2505 (N_2505,N_1877,N_1807);
and U2506 (N_2506,N_1518,N_1816);
or U2507 (N_2507,N_2216,N_1895);
and U2508 (N_2508,N_1808,N_1677);
and U2509 (N_2509,N_2220,N_2042);
or U2510 (N_2510,N_1544,N_1749);
nand U2511 (N_2511,N_1724,N_1953);
and U2512 (N_2512,N_1667,N_1700);
nor U2513 (N_2513,N_1693,N_1939);
nor U2514 (N_2514,N_2066,N_1931);
and U2515 (N_2515,N_2058,N_1537);
or U2516 (N_2516,N_1950,N_1589);
nand U2517 (N_2517,N_1770,N_2054);
nand U2518 (N_2518,N_1503,N_1632);
and U2519 (N_2519,N_2173,N_1509);
and U2520 (N_2520,N_1932,N_1906);
xnor U2521 (N_2521,N_2181,N_1849);
or U2522 (N_2522,N_2152,N_1501);
and U2523 (N_2523,N_1702,N_1626);
xor U2524 (N_2524,N_2060,N_1889);
and U2525 (N_2525,N_1812,N_1766);
nand U2526 (N_2526,N_1803,N_1609);
and U2527 (N_2527,N_1546,N_1777);
nand U2528 (N_2528,N_1707,N_1593);
nor U2529 (N_2529,N_2095,N_1956);
nor U2530 (N_2530,N_1594,N_2041);
nor U2531 (N_2531,N_1533,N_2004);
nand U2532 (N_2532,N_1819,N_1523);
nand U2533 (N_2533,N_1883,N_2108);
nor U2534 (N_2534,N_2237,N_1927);
xnor U2535 (N_2535,N_2114,N_2007);
and U2536 (N_2536,N_2187,N_1997);
nand U2537 (N_2537,N_1720,N_1620);
nand U2538 (N_2538,N_2037,N_1619);
nor U2539 (N_2539,N_1861,N_2155);
nor U2540 (N_2540,N_1535,N_1910);
nor U2541 (N_2541,N_1558,N_1519);
xnor U2542 (N_2542,N_2112,N_2015);
or U2543 (N_2543,N_2149,N_1727);
xor U2544 (N_2544,N_1732,N_1681);
and U2545 (N_2545,N_1524,N_2192);
and U2546 (N_2546,N_1966,N_2130);
nor U2547 (N_2547,N_2100,N_1674);
nand U2548 (N_2548,N_1545,N_1785);
nor U2549 (N_2549,N_1940,N_1899);
or U2550 (N_2550,N_1892,N_2113);
or U2551 (N_2551,N_1799,N_2174);
nor U2552 (N_2552,N_2099,N_1551);
and U2553 (N_2553,N_2126,N_2080);
or U2554 (N_2554,N_1569,N_1680);
nand U2555 (N_2555,N_1507,N_2185);
nor U2556 (N_2556,N_2246,N_1821);
or U2557 (N_2557,N_1794,N_2098);
xnor U2558 (N_2558,N_1679,N_2243);
and U2559 (N_2559,N_1623,N_1758);
and U2560 (N_2560,N_1723,N_1585);
and U2561 (N_2561,N_2062,N_2022);
or U2562 (N_2562,N_1582,N_1525);
nand U2563 (N_2563,N_1776,N_1719);
and U2564 (N_2564,N_2047,N_1606);
xnor U2565 (N_2565,N_1686,N_1841);
and U2566 (N_2566,N_1806,N_1506);
nor U2567 (N_2567,N_1909,N_1534);
nand U2568 (N_2568,N_1835,N_2124);
nor U2569 (N_2569,N_1696,N_2201);
nand U2570 (N_2570,N_2232,N_1510);
and U2571 (N_2571,N_1755,N_1882);
nor U2572 (N_2572,N_2176,N_2180);
xor U2573 (N_2573,N_2212,N_2229);
nand U2574 (N_2574,N_1853,N_2049);
xor U2575 (N_2575,N_2137,N_1746);
or U2576 (N_2576,N_2072,N_1607);
nand U2577 (N_2577,N_1993,N_1573);
and U2578 (N_2578,N_1917,N_1792);
or U2579 (N_2579,N_1600,N_2241);
and U2580 (N_2580,N_1933,N_2215);
nor U2581 (N_2581,N_2219,N_1866);
and U2582 (N_2582,N_1780,N_2025);
xor U2583 (N_2583,N_1734,N_1663);
xor U2584 (N_2584,N_2214,N_2194);
or U2585 (N_2585,N_1771,N_1936);
nor U2586 (N_2586,N_1858,N_1587);
and U2587 (N_2587,N_1576,N_1520);
and U2588 (N_2588,N_2104,N_1961);
nand U2589 (N_2589,N_1995,N_1636);
nor U2590 (N_2590,N_2198,N_1763);
nand U2591 (N_2591,N_1710,N_1752);
and U2592 (N_2592,N_1827,N_2009);
nand U2593 (N_2593,N_1635,N_1515);
xnor U2594 (N_2594,N_1884,N_1668);
xor U2595 (N_2595,N_2245,N_1985);
xnor U2596 (N_2596,N_1854,N_1740);
xnor U2597 (N_2597,N_1857,N_1617);
nand U2598 (N_2598,N_1603,N_1845);
nand U2599 (N_2599,N_1561,N_1706);
or U2600 (N_2600,N_1984,N_2063);
or U2601 (N_2601,N_1657,N_2161);
and U2602 (N_2602,N_1608,N_1891);
nand U2603 (N_2603,N_1810,N_2017);
or U2604 (N_2604,N_1572,N_1722);
nor U2605 (N_2605,N_1514,N_1862);
nor U2606 (N_2606,N_1612,N_1935);
xnor U2607 (N_2607,N_1963,N_1946);
nand U2608 (N_2608,N_1778,N_1920);
and U2609 (N_2609,N_1562,N_2239);
and U2610 (N_2610,N_2078,N_1690);
nand U2611 (N_2611,N_2052,N_1664);
xnor U2612 (N_2612,N_1711,N_1565);
xnor U2613 (N_2613,N_2129,N_1787);
xor U2614 (N_2614,N_1599,N_1851);
nand U2615 (N_2615,N_2225,N_1641);
or U2616 (N_2616,N_2188,N_1526);
and U2617 (N_2617,N_1521,N_1666);
xor U2618 (N_2618,N_2005,N_1566);
nor U2619 (N_2619,N_1716,N_1855);
nor U2620 (N_2620,N_2092,N_1987);
or U2621 (N_2621,N_2024,N_1823);
nor U2622 (N_2622,N_2065,N_2121);
and U2623 (N_2623,N_1601,N_2186);
xor U2624 (N_2624,N_1512,N_1670);
nand U2625 (N_2625,N_2065,N_1591);
and U2626 (N_2626,N_1758,N_1536);
nand U2627 (N_2627,N_1668,N_2043);
and U2628 (N_2628,N_1783,N_1701);
nor U2629 (N_2629,N_1841,N_1654);
and U2630 (N_2630,N_1916,N_1691);
or U2631 (N_2631,N_2231,N_2142);
nor U2632 (N_2632,N_1704,N_1646);
xnor U2633 (N_2633,N_1790,N_2232);
nand U2634 (N_2634,N_1538,N_2127);
xnor U2635 (N_2635,N_2040,N_2012);
or U2636 (N_2636,N_1762,N_1882);
nor U2637 (N_2637,N_2120,N_1784);
xnor U2638 (N_2638,N_2205,N_1573);
nor U2639 (N_2639,N_2191,N_1873);
or U2640 (N_2640,N_1542,N_1877);
and U2641 (N_2641,N_1693,N_1702);
or U2642 (N_2642,N_1678,N_1660);
nand U2643 (N_2643,N_1793,N_1831);
and U2644 (N_2644,N_1716,N_1570);
xnor U2645 (N_2645,N_1545,N_2023);
or U2646 (N_2646,N_1537,N_1706);
xor U2647 (N_2647,N_1549,N_1573);
xnor U2648 (N_2648,N_1624,N_1847);
or U2649 (N_2649,N_2239,N_1995);
or U2650 (N_2650,N_2076,N_1868);
nor U2651 (N_2651,N_1736,N_2084);
or U2652 (N_2652,N_1733,N_1592);
nor U2653 (N_2653,N_1519,N_1653);
nand U2654 (N_2654,N_2135,N_1820);
xor U2655 (N_2655,N_1905,N_2025);
or U2656 (N_2656,N_1861,N_1881);
nor U2657 (N_2657,N_1851,N_1598);
and U2658 (N_2658,N_2215,N_1642);
xor U2659 (N_2659,N_2005,N_2042);
and U2660 (N_2660,N_2079,N_1931);
nand U2661 (N_2661,N_1974,N_2170);
and U2662 (N_2662,N_2230,N_1934);
or U2663 (N_2663,N_1760,N_1664);
nand U2664 (N_2664,N_1651,N_2070);
and U2665 (N_2665,N_1970,N_1720);
nand U2666 (N_2666,N_1984,N_2098);
nor U2667 (N_2667,N_1736,N_1792);
nand U2668 (N_2668,N_2105,N_2063);
or U2669 (N_2669,N_1504,N_2089);
nor U2670 (N_2670,N_1615,N_2130);
or U2671 (N_2671,N_1568,N_1854);
and U2672 (N_2672,N_2106,N_2128);
xnor U2673 (N_2673,N_2102,N_2198);
xor U2674 (N_2674,N_1520,N_2182);
xnor U2675 (N_2675,N_1520,N_1699);
or U2676 (N_2676,N_1756,N_2114);
nor U2677 (N_2677,N_1971,N_2126);
nand U2678 (N_2678,N_1834,N_1590);
xnor U2679 (N_2679,N_2245,N_1527);
nand U2680 (N_2680,N_1916,N_1505);
and U2681 (N_2681,N_1525,N_1504);
nor U2682 (N_2682,N_2014,N_2177);
nand U2683 (N_2683,N_1942,N_1741);
and U2684 (N_2684,N_2114,N_1640);
nor U2685 (N_2685,N_1948,N_1862);
or U2686 (N_2686,N_1867,N_1979);
nor U2687 (N_2687,N_1780,N_2150);
nand U2688 (N_2688,N_1890,N_1719);
nor U2689 (N_2689,N_1670,N_1983);
or U2690 (N_2690,N_1868,N_2127);
or U2691 (N_2691,N_2131,N_2177);
and U2692 (N_2692,N_2047,N_2150);
and U2693 (N_2693,N_2084,N_1697);
and U2694 (N_2694,N_1807,N_1858);
nor U2695 (N_2695,N_1623,N_1773);
nand U2696 (N_2696,N_1783,N_1575);
xnor U2697 (N_2697,N_2242,N_1548);
or U2698 (N_2698,N_1944,N_1695);
and U2699 (N_2699,N_2002,N_2182);
or U2700 (N_2700,N_1527,N_2140);
nand U2701 (N_2701,N_1763,N_1515);
or U2702 (N_2702,N_1583,N_2073);
xor U2703 (N_2703,N_1605,N_1511);
and U2704 (N_2704,N_1745,N_1942);
nand U2705 (N_2705,N_1779,N_1843);
nor U2706 (N_2706,N_2176,N_1575);
nand U2707 (N_2707,N_2099,N_1672);
and U2708 (N_2708,N_1971,N_1621);
nand U2709 (N_2709,N_1887,N_2077);
and U2710 (N_2710,N_2249,N_1608);
and U2711 (N_2711,N_1598,N_1732);
or U2712 (N_2712,N_1651,N_2249);
nor U2713 (N_2713,N_1910,N_1719);
nor U2714 (N_2714,N_1548,N_1921);
or U2715 (N_2715,N_1588,N_2069);
and U2716 (N_2716,N_1738,N_2159);
xor U2717 (N_2717,N_1802,N_1864);
nor U2718 (N_2718,N_1789,N_2178);
nand U2719 (N_2719,N_2179,N_1827);
nand U2720 (N_2720,N_1777,N_1897);
xnor U2721 (N_2721,N_2231,N_2179);
or U2722 (N_2722,N_1784,N_2225);
nand U2723 (N_2723,N_2102,N_1561);
xnor U2724 (N_2724,N_1537,N_1555);
xnor U2725 (N_2725,N_1925,N_2143);
xnor U2726 (N_2726,N_2054,N_1855);
or U2727 (N_2727,N_1894,N_1553);
nor U2728 (N_2728,N_2131,N_1652);
xnor U2729 (N_2729,N_2218,N_2039);
nand U2730 (N_2730,N_1713,N_1520);
xnor U2731 (N_2731,N_2214,N_1778);
nand U2732 (N_2732,N_1684,N_1607);
or U2733 (N_2733,N_2166,N_1540);
xor U2734 (N_2734,N_2160,N_1855);
nor U2735 (N_2735,N_1866,N_1838);
and U2736 (N_2736,N_1613,N_1989);
or U2737 (N_2737,N_1831,N_1532);
nand U2738 (N_2738,N_1788,N_2044);
and U2739 (N_2739,N_2003,N_1605);
xor U2740 (N_2740,N_1821,N_2055);
nand U2741 (N_2741,N_1811,N_1575);
or U2742 (N_2742,N_1949,N_1664);
and U2743 (N_2743,N_2144,N_1715);
xor U2744 (N_2744,N_2064,N_1596);
nand U2745 (N_2745,N_2173,N_1648);
and U2746 (N_2746,N_1715,N_2156);
xnor U2747 (N_2747,N_2051,N_1776);
or U2748 (N_2748,N_1605,N_1808);
nand U2749 (N_2749,N_1621,N_1710);
xor U2750 (N_2750,N_2125,N_1797);
and U2751 (N_2751,N_1510,N_2111);
and U2752 (N_2752,N_1686,N_2108);
or U2753 (N_2753,N_1624,N_1740);
or U2754 (N_2754,N_1728,N_2168);
nor U2755 (N_2755,N_1798,N_1738);
nand U2756 (N_2756,N_1522,N_1904);
or U2757 (N_2757,N_1625,N_2231);
nor U2758 (N_2758,N_1670,N_2136);
or U2759 (N_2759,N_1970,N_2037);
and U2760 (N_2760,N_1799,N_1738);
nand U2761 (N_2761,N_1861,N_1520);
and U2762 (N_2762,N_1925,N_1756);
nor U2763 (N_2763,N_2171,N_1720);
and U2764 (N_2764,N_1775,N_1784);
nand U2765 (N_2765,N_1723,N_2175);
xnor U2766 (N_2766,N_2202,N_2222);
nand U2767 (N_2767,N_1595,N_1854);
nand U2768 (N_2768,N_1963,N_1678);
or U2769 (N_2769,N_2102,N_1596);
nand U2770 (N_2770,N_2057,N_1641);
nand U2771 (N_2771,N_1839,N_1552);
or U2772 (N_2772,N_1551,N_2069);
and U2773 (N_2773,N_1565,N_2017);
and U2774 (N_2774,N_1527,N_1823);
nor U2775 (N_2775,N_1840,N_1866);
and U2776 (N_2776,N_1624,N_1964);
nand U2777 (N_2777,N_2037,N_2036);
or U2778 (N_2778,N_2093,N_1845);
nor U2779 (N_2779,N_1781,N_2038);
and U2780 (N_2780,N_1870,N_1953);
and U2781 (N_2781,N_1569,N_2077);
and U2782 (N_2782,N_2067,N_1788);
and U2783 (N_2783,N_1892,N_1943);
nand U2784 (N_2784,N_2000,N_2176);
and U2785 (N_2785,N_2137,N_1681);
nor U2786 (N_2786,N_2013,N_1547);
and U2787 (N_2787,N_1779,N_1627);
nor U2788 (N_2788,N_2006,N_1540);
and U2789 (N_2789,N_1843,N_1670);
xor U2790 (N_2790,N_1665,N_1539);
nor U2791 (N_2791,N_2225,N_1632);
or U2792 (N_2792,N_1884,N_1544);
and U2793 (N_2793,N_2235,N_1752);
or U2794 (N_2794,N_2103,N_1760);
nor U2795 (N_2795,N_1755,N_1920);
xor U2796 (N_2796,N_1762,N_1520);
xnor U2797 (N_2797,N_1602,N_2076);
nor U2798 (N_2798,N_1733,N_1918);
or U2799 (N_2799,N_2081,N_1561);
and U2800 (N_2800,N_2062,N_1994);
nor U2801 (N_2801,N_1999,N_1731);
or U2802 (N_2802,N_1989,N_2069);
nor U2803 (N_2803,N_2028,N_1969);
nand U2804 (N_2804,N_1796,N_1624);
and U2805 (N_2805,N_1537,N_1603);
nand U2806 (N_2806,N_1679,N_1763);
nor U2807 (N_2807,N_2185,N_1849);
and U2808 (N_2808,N_2034,N_1716);
and U2809 (N_2809,N_2100,N_2046);
nand U2810 (N_2810,N_2059,N_1500);
xor U2811 (N_2811,N_1924,N_1904);
and U2812 (N_2812,N_2101,N_1654);
and U2813 (N_2813,N_2237,N_1681);
nand U2814 (N_2814,N_2183,N_2014);
nand U2815 (N_2815,N_1563,N_1613);
nor U2816 (N_2816,N_1667,N_1772);
xor U2817 (N_2817,N_1987,N_2022);
nand U2818 (N_2818,N_1967,N_1714);
xnor U2819 (N_2819,N_1867,N_1648);
and U2820 (N_2820,N_1651,N_2089);
nor U2821 (N_2821,N_1714,N_1792);
or U2822 (N_2822,N_1843,N_1744);
and U2823 (N_2823,N_1922,N_1612);
or U2824 (N_2824,N_1917,N_1645);
or U2825 (N_2825,N_1631,N_2034);
nor U2826 (N_2826,N_2043,N_2146);
nand U2827 (N_2827,N_1614,N_2204);
or U2828 (N_2828,N_1813,N_1636);
nor U2829 (N_2829,N_2108,N_1999);
nor U2830 (N_2830,N_1584,N_2028);
nor U2831 (N_2831,N_1754,N_1612);
nand U2832 (N_2832,N_1901,N_1918);
or U2833 (N_2833,N_1606,N_1614);
and U2834 (N_2834,N_1618,N_2088);
xor U2835 (N_2835,N_1969,N_2228);
nor U2836 (N_2836,N_1509,N_2134);
nand U2837 (N_2837,N_2186,N_2084);
or U2838 (N_2838,N_1835,N_1581);
nor U2839 (N_2839,N_1606,N_1578);
nand U2840 (N_2840,N_1806,N_2249);
xnor U2841 (N_2841,N_2243,N_1586);
or U2842 (N_2842,N_1791,N_1557);
xor U2843 (N_2843,N_1630,N_2069);
nand U2844 (N_2844,N_2036,N_2111);
and U2845 (N_2845,N_1759,N_2026);
nor U2846 (N_2846,N_2214,N_1831);
nand U2847 (N_2847,N_1532,N_2037);
nand U2848 (N_2848,N_1976,N_1666);
or U2849 (N_2849,N_2114,N_1910);
nand U2850 (N_2850,N_1799,N_1529);
nand U2851 (N_2851,N_1767,N_1926);
nand U2852 (N_2852,N_2144,N_1959);
and U2853 (N_2853,N_1544,N_1852);
nor U2854 (N_2854,N_2242,N_1515);
or U2855 (N_2855,N_2241,N_1667);
nor U2856 (N_2856,N_1585,N_1693);
and U2857 (N_2857,N_2241,N_2198);
nand U2858 (N_2858,N_1852,N_2103);
and U2859 (N_2859,N_1650,N_1831);
nand U2860 (N_2860,N_1841,N_2152);
and U2861 (N_2861,N_1977,N_2214);
nor U2862 (N_2862,N_2163,N_1949);
xor U2863 (N_2863,N_1973,N_1565);
and U2864 (N_2864,N_1626,N_2165);
xnor U2865 (N_2865,N_1599,N_2094);
and U2866 (N_2866,N_1918,N_2001);
nand U2867 (N_2867,N_1560,N_2237);
or U2868 (N_2868,N_1862,N_1610);
and U2869 (N_2869,N_2013,N_1816);
xor U2870 (N_2870,N_1627,N_1800);
or U2871 (N_2871,N_2102,N_2206);
or U2872 (N_2872,N_1646,N_1897);
nand U2873 (N_2873,N_2141,N_2170);
nor U2874 (N_2874,N_1828,N_2028);
and U2875 (N_2875,N_1547,N_1515);
nor U2876 (N_2876,N_2249,N_1989);
nor U2877 (N_2877,N_2043,N_1949);
xor U2878 (N_2878,N_1789,N_2139);
or U2879 (N_2879,N_1580,N_2024);
nor U2880 (N_2880,N_1698,N_2227);
nand U2881 (N_2881,N_1697,N_2027);
or U2882 (N_2882,N_1873,N_1652);
xnor U2883 (N_2883,N_2197,N_2164);
xnor U2884 (N_2884,N_2177,N_2112);
nand U2885 (N_2885,N_2077,N_1677);
nand U2886 (N_2886,N_2005,N_2148);
nand U2887 (N_2887,N_2117,N_1606);
and U2888 (N_2888,N_1855,N_1607);
or U2889 (N_2889,N_1595,N_2240);
and U2890 (N_2890,N_2036,N_2201);
xor U2891 (N_2891,N_1702,N_1821);
and U2892 (N_2892,N_1860,N_1659);
or U2893 (N_2893,N_1883,N_1725);
nand U2894 (N_2894,N_1565,N_1851);
xor U2895 (N_2895,N_1827,N_1768);
or U2896 (N_2896,N_1962,N_2038);
or U2897 (N_2897,N_1994,N_1739);
or U2898 (N_2898,N_1690,N_1871);
nor U2899 (N_2899,N_1909,N_1843);
nor U2900 (N_2900,N_2177,N_2012);
or U2901 (N_2901,N_2010,N_2053);
xnor U2902 (N_2902,N_2205,N_1946);
and U2903 (N_2903,N_1675,N_1612);
or U2904 (N_2904,N_2037,N_2245);
xor U2905 (N_2905,N_1719,N_1505);
xnor U2906 (N_2906,N_1518,N_1586);
xor U2907 (N_2907,N_1710,N_1936);
nand U2908 (N_2908,N_2056,N_1570);
nor U2909 (N_2909,N_1884,N_2172);
and U2910 (N_2910,N_1506,N_1919);
nand U2911 (N_2911,N_2229,N_1510);
nand U2912 (N_2912,N_1899,N_1711);
nor U2913 (N_2913,N_2034,N_1579);
nand U2914 (N_2914,N_2138,N_1750);
or U2915 (N_2915,N_1562,N_2106);
or U2916 (N_2916,N_2145,N_1721);
xor U2917 (N_2917,N_2193,N_2180);
nand U2918 (N_2918,N_2017,N_2076);
xor U2919 (N_2919,N_2111,N_1600);
nand U2920 (N_2920,N_1857,N_1793);
or U2921 (N_2921,N_1990,N_2028);
and U2922 (N_2922,N_1833,N_2080);
nand U2923 (N_2923,N_2131,N_1808);
nand U2924 (N_2924,N_1869,N_1984);
nand U2925 (N_2925,N_1557,N_1869);
nor U2926 (N_2926,N_1901,N_1764);
or U2927 (N_2927,N_2112,N_1770);
nand U2928 (N_2928,N_1942,N_1994);
nor U2929 (N_2929,N_2162,N_1505);
nor U2930 (N_2930,N_2046,N_1533);
or U2931 (N_2931,N_2159,N_2073);
nand U2932 (N_2932,N_2140,N_1838);
and U2933 (N_2933,N_2156,N_1690);
or U2934 (N_2934,N_1968,N_2114);
nand U2935 (N_2935,N_2119,N_2136);
or U2936 (N_2936,N_1671,N_2101);
nand U2937 (N_2937,N_2154,N_1523);
and U2938 (N_2938,N_1602,N_1611);
xnor U2939 (N_2939,N_2227,N_1608);
nor U2940 (N_2940,N_2007,N_1636);
or U2941 (N_2941,N_1524,N_1501);
nand U2942 (N_2942,N_1640,N_2002);
xor U2943 (N_2943,N_1501,N_1666);
xor U2944 (N_2944,N_2240,N_1534);
and U2945 (N_2945,N_2211,N_2000);
or U2946 (N_2946,N_2136,N_1978);
nand U2947 (N_2947,N_1978,N_2155);
nand U2948 (N_2948,N_1746,N_1988);
nor U2949 (N_2949,N_1551,N_2093);
xnor U2950 (N_2950,N_1615,N_1511);
nand U2951 (N_2951,N_1775,N_2100);
and U2952 (N_2952,N_1923,N_2094);
nand U2953 (N_2953,N_1731,N_1914);
or U2954 (N_2954,N_1784,N_1551);
xnor U2955 (N_2955,N_1993,N_1761);
xnor U2956 (N_2956,N_1894,N_1660);
nor U2957 (N_2957,N_1992,N_2177);
xor U2958 (N_2958,N_2023,N_1533);
nor U2959 (N_2959,N_1702,N_1866);
nand U2960 (N_2960,N_1682,N_1746);
xnor U2961 (N_2961,N_1990,N_1944);
xnor U2962 (N_2962,N_1865,N_2024);
xor U2963 (N_2963,N_1661,N_1814);
xor U2964 (N_2964,N_1742,N_2131);
or U2965 (N_2965,N_2014,N_2078);
nand U2966 (N_2966,N_2162,N_2048);
or U2967 (N_2967,N_2017,N_2025);
nor U2968 (N_2968,N_2157,N_1723);
or U2969 (N_2969,N_1696,N_1805);
and U2970 (N_2970,N_2016,N_1964);
or U2971 (N_2971,N_2246,N_1522);
or U2972 (N_2972,N_1780,N_1676);
or U2973 (N_2973,N_2125,N_1732);
and U2974 (N_2974,N_1614,N_1967);
xor U2975 (N_2975,N_1548,N_2078);
and U2976 (N_2976,N_1838,N_1698);
nand U2977 (N_2977,N_1833,N_1657);
xnor U2978 (N_2978,N_1809,N_2188);
xnor U2979 (N_2979,N_1518,N_1627);
and U2980 (N_2980,N_2120,N_1575);
nand U2981 (N_2981,N_2162,N_1626);
or U2982 (N_2982,N_1925,N_1759);
and U2983 (N_2983,N_1815,N_1779);
and U2984 (N_2984,N_1796,N_1999);
xor U2985 (N_2985,N_1875,N_1989);
nor U2986 (N_2986,N_1622,N_2184);
or U2987 (N_2987,N_2130,N_1599);
nand U2988 (N_2988,N_1866,N_1568);
and U2989 (N_2989,N_2191,N_2237);
or U2990 (N_2990,N_2063,N_1654);
and U2991 (N_2991,N_1782,N_1978);
and U2992 (N_2992,N_1933,N_2046);
or U2993 (N_2993,N_2234,N_1875);
or U2994 (N_2994,N_1697,N_1961);
or U2995 (N_2995,N_2159,N_1630);
xor U2996 (N_2996,N_1542,N_2193);
or U2997 (N_2997,N_1846,N_1514);
xor U2998 (N_2998,N_2000,N_1923);
and U2999 (N_2999,N_1957,N_1733);
nor UO_0 (O_0,N_2440,N_2592);
nor UO_1 (O_1,N_2741,N_2344);
or UO_2 (O_2,N_2901,N_2300);
nand UO_3 (O_3,N_2808,N_2327);
and UO_4 (O_4,N_2670,N_2257);
and UO_5 (O_5,N_2416,N_2929);
nor UO_6 (O_6,N_2683,N_2462);
nor UO_7 (O_7,N_2654,N_2404);
xnor UO_8 (O_8,N_2943,N_2413);
and UO_9 (O_9,N_2524,N_2915);
or UO_10 (O_10,N_2349,N_2981);
xor UO_11 (O_11,N_2628,N_2730);
and UO_12 (O_12,N_2742,N_2375);
nor UO_13 (O_13,N_2348,N_2704);
and UO_14 (O_14,N_2615,N_2582);
and UO_15 (O_15,N_2378,N_2284);
xor UO_16 (O_16,N_2955,N_2698);
xnor UO_17 (O_17,N_2969,N_2547);
and UO_18 (O_18,N_2429,N_2775);
xor UO_19 (O_19,N_2471,N_2590);
and UO_20 (O_20,N_2398,N_2361);
nor UO_21 (O_21,N_2574,N_2371);
or UO_22 (O_22,N_2987,N_2820);
nor UO_23 (O_23,N_2304,N_2265);
and UO_24 (O_24,N_2934,N_2766);
nor UO_25 (O_25,N_2566,N_2609);
or UO_26 (O_26,N_2713,N_2695);
or UO_27 (O_27,N_2840,N_2897);
and UO_28 (O_28,N_2390,N_2671);
and UO_29 (O_29,N_2858,N_2294);
and UO_30 (O_30,N_2424,N_2627);
xor UO_31 (O_31,N_2639,N_2703);
nand UO_32 (O_32,N_2924,N_2912);
and UO_33 (O_33,N_2707,N_2495);
xnor UO_34 (O_34,N_2382,N_2586);
nor UO_35 (O_35,N_2258,N_2759);
nand UO_36 (O_36,N_2391,N_2965);
nor UO_37 (O_37,N_2485,N_2826);
and UO_38 (O_38,N_2320,N_2283);
and UO_39 (O_39,N_2802,N_2997);
nand UO_40 (O_40,N_2807,N_2461);
xor UO_41 (O_41,N_2958,N_2352);
nand UO_42 (O_42,N_2403,N_2800);
xor UO_43 (O_43,N_2816,N_2844);
or UO_44 (O_44,N_2530,N_2596);
nand UO_45 (O_45,N_2752,N_2922);
nand UO_46 (O_46,N_2666,N_2968);
or UO_47 (O_47,N_2857,N_2303);
and UO_48 (O_48,N_2837,N_2657);
xor UO_49 (O_49,N_2674,N_2815);
or UO_50 (O_50,N_2556,N_2748);
xnor UO_51 (O_51,N_2939,N_2519);
and UO_52 (O_52,N_2921,N_2267);
xor UO_53 (O_53,N_2710,N_2677);
or UO_54 (O_54,N_2942,N_2812);
or UO_55 (O_55,N_2388,N_2863);
nor UO_56 (O_56,N_2291,N_2555);
or UO_57 (O_57,N_2892,N_2493);
and UO_58 (O_58,N_2790,N_2540);
and UO_59 (O_59,N_2268,N_2908);
and UO_60 (O_60,N_2644,N_2684);
and UO_61 (O_61,N_2309,N_2410);
nor UO_62 (O_62,N_2434,N_2467);
and UO_63 (O_63,N_2266,N_2868);
or UO_64 (O_64,N_2894,N_2399);
nor UO_65 (O_65,N_2274,N_2792);
nor UO_66 (O_66,N_2598,N_2720);
nor UO_67 (O_67,N_2708,N_2822);
nor UO_68 (O_68,N_2646,N_2597);
nand UO_69 (O_69,N_2405,N_2636);
nor UO_70 (O_70,N_2805,N_2281);
nor UO_71 (O_71,N_2712,N_2865);
nand UO_72 (O_72,N_2801,N_2269);
xnor UO_73 (O_73,N_2705,N_2570);
or UO_74 (O_74,N_2451,N_2262);
or UO_75 (O_75,N_2867,N_2484);
xor UO_76 (O_76,N_2308,N_2389);
xor UO_77 (O_77,N_2438,N_2446);
or UO_78 (O_78,N_2675,N_2862);
or UO_79 (O_79,N_2907,N_2575);
and UO_80 (O_80,N_2848,N_2458);
and UO_81 (O_81,N_2831,N_2771);
or UO_82 (O_82,N_2412,N_2854);
or UO_83 (O_83,N_2601,N_2548);
or UO_84 (O_84,N_2311,N_2884);
nor UO_85 (O_85,N_2585,N_2750);
and UO_86 (O_86,N_2285,N_2515);
nand UO_87 (O_87,N_2254,N_2895);
nand UO_88 (O_88,N_2838,N_2879);
and UO_89 (O_89,N_2472,N_2558);
xnor UO_90 (O_90,N_2487,N_2717);
and UO_91 (O_91,N_2605,N_2918);
or UO_92 (O_92,N_2692,N_2761);
or UO_93 (O_93,N_2847,N_2439);
xnor UO_94 (O_94,N_2287,N_2364);
nand UO_95 (O_95,N_2803,N_2612);
xnor UO_96 (O_96,N_2629,N_2679);
or UO_97 (O_97,N_2905,N_2441);
nand UO_98 (O_98,N_2278,N_2874);
and UO_99 (O_99,N_2443,N_2937);
nand UO_100 (O_100,N_2641,N_2643);
nor UO_101 (O_101,N_2568,N_2420);
and UO_102 (O_102,N_2367,N_2850);
or UO_103 (O_103,N_2474,N_2406);
and UO_104 (O_104,N_2353,N_2966);
nand UO_105 (O_105,N_2326,N_2632);
nand UO_106 (O_106,N_2588,N_2302);
nand UO_107 (O_107,N_2913,N_2542);
nand UO_108 (O_108,N_2277,N_2749);
nand UO_109 (O_109,N_2743,N_2333);
xor UO_110 (O_110,N_2944,N_2919);
xnor UO_111 (O_111,N_2655,N_2301);
or UO_112 (O_112,N_2562,N_2473);
nand UO_113 (O_113,N_2290,N_2976);
nand UO_114 (O_114,N_2337,N_2888);
xor UO_115 (O_115,N_2984,N_2516);
or UO_116 (O_116,N_2680,N_2572);
or UO_117 (O_117,N_2450,N_2383);
nor UO_118 (O_118,N_2700,N_2756);
or UO_119 (O_119,N_2264,N_2841);
or UO_120 (O_120,N_2673,N_2885);
or UO_121 (O_121,N_2699,N_2975);
and UO_122 (O_122,N_2448,N_2925);
nor UO_123 (O_123,N_2297,N_2830);
nor UO_124 (O_124,N_2397,N_2422);
nor UO_125 (O_125,N_2469,N_2559);
or UO_126 (O_126,N_2456,N_2339);
and UO_127 (O_127,N_2370,N_2251);
nor UO_128 (O_128,N_2619,N_2343);
nand UO_129 (O_129,N_2535,N_2881);
xnor UO_130 (O_130,N_2649,N_2324);
nor UO_131 (O_131,N_2583,N_2538);
and UO_132 (O_132,N_2764,N_2411);
nand UO_133 (O_133,N_2864,N_2634);
nand UO_134 (O_134,N_2444,N_2853);
nor UO_135 (O_135,N_2701,N_2736);
xnor UO_136 (O_136,N_2724,N_2738);
xnor UO_137 (O_137,N_2505,N_2490);
or UO_138 (O_138,N_2319,N_2433);
nor UO_139 (O_139,N_2476,N_2691);
xnor UO_140 (O_140,N_2956,N_2616);
or UO_141 (O_141,N_2543,N_2718);
nor UO_142 (O_142,N_2503,N_2263);
nor UO_143 (O_143,N_2466,N_2656);
nor UO_144 (O_144,N_2739,N_2255);
xnor UO_145 (O_145,N_2332,N_2408);
or UO_146 (O_146,N_2638,N_2521);
xor UO_147 (O_147,N_2647,N_2936);
and UO_148 (O_148,N_2839,N_2386);
and UO_149 (O_149,N_2380,N_2791);
or UO_150 (O_150,N_2475,N_2729);
nor UO_151 (O_151,N_2565,N_2525);
nand UO_152 (O_152,N_2777,N_2664);
and UO_153 (O_153,N_2306,N_2415);
and UO_154 (O_154,N_2366,N_2998);
nor UO_155 (O_155,N_2726,N_2902);
and UO_156 (O_156,N_2381,N_2722);
xor UO_157 (O_157,N_2686,N_2904);
nand UO_158 (O_158,N_2569,N_2401);
xor UO_159 (O_159,N_2793,N_2661);
and UO_160 (O_160,N_2479,N_2829);
nand UO_161 (O_161,N_2614,N_2983);
nor UO_162 (O_162,N_2810,N_2532);
or UO_163 (O_163,N_2781,N_2866);
nor UO_164 (O_164,N_2501,N_2445);
nor UO_165 (O_165,N_2407,N_2906);
nand UO_166 (O_166,N_2607,N_2253);
nand UO_167 (O_167,N_2681,N_2876);
xor UO_168 (O_168,N_2527,N_2914);
xor UO_169 (O_169,N_2788,N_2869);
and UO_170 (O_170,N_2512,N_2312);
or UO_171 (O_171,N_2536,N_2940);
or UO_172 (O_172,N_2359,N_2789);
nor UO_173 (O_173,N_2427,N_2967);
or UO_174 (O_174,N_2676,N_2957);
and UO_175 (O_175,N_2355,N_2552);
and UO_176 (O_176,N_2986,N_2506);
and UO_177 (O_177,N_2325,N_2447);
and UO_178 (O_178,N_2950,N_2425);
nand UO_179 (O_179,N_2604,N_2488);
xnor UO_180 (O_180,N_2694,N_2658);
and UO_181 (O_181,N_2755,N_2814);
and UO_182 (O_182,N_2414,N_2991);
nand UO_183 (O_183,N_2859,N_2457);
nand UO_184 (O_184,N_2331,N_2637);
or UO_185 (O_185,N_2497,N_2533);
nor UO_186 (O_186,N_2977,N_2836);
xnor UO_187 (O_187,N_2642,N_2546);
or UO_188 (O_188,N_2577,N_2785);
xor UO_189 (O_189,N_2368,N_2786);
nand UO_190 (O_190,N_2953,N_2298);
and UO_191 (O_191,N_2843,N_2514);
nand UO_192 (O_192,N_2606,N_2502);
nand UO_193 (O_193,N_2685,N_2280);
and UO_194 (O_194,N_2554,N_2758);
nand UO_195 (O_195,N_2307,N_2377);
and UO_196 (O_196,N_2618,N_2455);
nand UO_197 (O_197,N_2318,N_2809);
and UO_198 (O_198,N_2599,N_2982);
or UO_199 (O_199,N_2464,N_2948);
xor UO_200 (O_200,N_2932,N_2891);
nand UO_201 (O_201,N_2477,N_2608);
nor UO_202 (O_202,N_2295,N_2715);
xnor UO_203 (O_203,N_2567,N_2824);
nor UO_204 (O_204,N_2323,N_2600);
xnor UO_205 (O_205,N_2587,N_2520);
and UO_206 (O_206,N_2350,N_2579);
xnor UO_207 (O_207,N_2633,N_2770);
nand UO_208 (O_208,N_2855,N_2883);
nor UO_209 (O_209,N_2351,N_2498);
and UO_210 (O_210,N_2470,N_2659);
nor UO_211 (O_211,N_2360,N_2395);
nand UO_212 (O_212,N_2910,N_2959);
and UO_213 (O_213,N_2293,N_2418);
xor UO_214 (O_214,N_2688,N_2563);
xnor UO_215 (O_215,N_2819,N_2979);
or UO_216 (O_216,N_2534,N_2875);
or UO_217 (O_217,N_2494,N_2751);
xnor UO_218 (O_218,N_2678,N_2328);
nand UO_219 (O_219,N_2964,N_2768);
nand UO_220 (O_220,N_2553,N_2421);
or UO_221 (O_221,N_2279,N_2354);
and UO_222 (O_222,N_2917,N_2362);
nor UO_223 (O_223,N_2949,N_2622);
and UO_224 (O_224,N_2663,N_2356);
nand UO_225 (O_225,N_2690,N_2322);
nand UO_226 (O_226,N_2341,N_2890);
xor UO_227 (O_227,N_2828,N_2845);
or UO_228 (O_228,N_2988,N_2709);
and UO_229 (O_229,N_2702,N_2511);
nor UO_230 (O_230,N_2896,N_2811);
or UO_231 (O_231,N_2276,N_2817);
and UO_232 (O_232,N_2365,N_2746);
nand UO_233 (O_233,N_2813,N_2760);
nand UO_234 (O_234,N_2486,N_2635);
xor UO_235 (O_235,N_2550,N_2591);
xor UO_236 (O_236,N_2797,N_2316);
xor UO_237 (O_237,N_2626,N_2693);
xor UO_238 (O_238,N_2728,N_2903);
nand UO_239 (O_239,N_2551,N_2711);
and UO_240 (O_240,N_2799,N_2541);
xor UO_241 (O_241,N_2423,N_2772);
nor UO_242 (O_242,N_2483,N_2992);
or UO_243 (O_243,N_2650,N_2767);
nor UO_244 (O_244,N_2878,N_2576);
or UO_245 (O_245,N_2299,N_2744);
xnor UO_246 (O_246,N_2522,N_2780);
nand UO_247 (O_247,N_2500,N_2782);
or UO_248 (O_248,N_2996,N_2727);
nor UO_249 (O_249,N_2453,N_2480);
and UO_250 (O_250,N_2787,N_2539);
or UO_251 (O_251,N_2273,N_2972);
and UO_252 (O_252,N_2594,N_2510);
and UO_253 (O_253,N_2652,N_2970);
or UO_254 (O_254,N_2832,N_2994);
and UO_255 (O_255,N_2459,N_2999);
nor UO_256 (O_256,N_2329,N_2396);
nand UO_257 (O_257,N_2610,N_2776);
and UO_258 (O_258,N_2887,N_2923);
or UO_259 (O_259,N_2426,N_2640);
nand UO_260 (O_260,N_2288,N_2737);
and UO_261 (O_261,N_2667,N_2321);
xnor UO_262 (O_262,N_2893,N_2305);
and UO_263 (O_263,N_2625,N_2825);
or UO_264 (O_264,N_2938,N_2962);
nor UO_265 (O_265,N_2252,N_2669);
nand UO_266 (O_266,N_2507,N_2732);
or UO_267 (O_267,N_2379,N_2261);
nand UO_268 (O_268,N_2765,N_2392);
xnor UO_269 (O_269,N_2376,N_2603);
nand UO_270 (O_270,N_2593,N_2260);
and UO_271 (O_271,N_2804,N_2660);
nand UO_272 (O_272,N_2282,N_2589);
nand UO_273 (O_273,N_2898,N_2584);
and UO_274 (O_274,N_2545,N_2400);
nor UO_275 (O_275,N_2409,N_2911);
and UO_276 (O_276,N_2794,N_2369);
nand UO_277 (O_277,N_2821,N_2842);
or UO_278 (O_278,N_2342,N_2774);
nor UO_279 (O_279,N_2928,N_2849);
and UO_280 (O_280,N_2989,N_2393);
nand UO_281 (O_281,N_2358,N_2385);
xor UO_282 (O_282,N_2315,N_2706);
nand UO_283 (O_283,N_2783,N_2916);
xor UO_284 (O_284,N_2581,N_2463);
and UO_285 (O_285,N_2452,N_2773);
nand UO_286 (O_286,N_2946,N_2431);
and UO_287 (O_287,N_2747,N_2973);
nor UO_288 (O_288,N_2531,N_2990);
or UO_289 (O_289,N_2481,N_2313);
and UO_290 (O_290,N_2733,N_2974);
xnor UO_291 (O_291,N_2544,N_2557);
nor UO_292 (O_292,N_2951,N_2734);
and UO_293 (O_293,N_2716,N_2564);
xor UO_294 (O_294,N_2560,N_2496);
or UO_295 (O_295,N_2769,N_2340);
and UO_296 (O_296,N_2721,N_2631);
and UO_297 (O_297,N_2900,N_2595);
nand UO_298 (O_298,N_2779,N_2714);
xor UO_299 (O_299,N_2334,N_2292);
nor UO_300 (O_300,N_2947,N_2995);
or UO_301 (O_301,N_2933,N_2835);
nor UO_302 (O_302,N_2330,N_2250);
nand UO_303 (O_303,N_2909,N_2602);
nand UO_304 (O_304,N_2952,N_2419);
or UO_305 (O_305,N_2920,N_2578);
or UO_306 (O_306,N_2927,N_2275);
nor UO_307 (O_307,N_2436,N_2296);
or UO_308 (O_308,N_2963,N_2509);
or UO_309 (O_309,N_2662,N_2549);
nor UO_310 (O_310,N_2806,N_2345);
xnor UO_311 (O_311,N_2373,N_2270);
and UO_312 (O_312,N_2271,N_2763);
or UO_313 (O_313,N_2719,N_2363);
nand UO_314 (O_314,N_2272,N_2796);
nor UO_315 (O_315,N_2945,N_2617);
and UO_316 (O_316,N_2665,N_2387);
nor UO_317 (O_317,N_2834,N_2468);
and UO_318 (O_318,N_2518,N_2613);
nand UO_319 (O_319,N_2314,N_2528);
nor UO_320 (O_320,N_2860,N_2336);
xor UO_321 (O_321,N_2523,N_2561);
nand UO_322 (O_322,N_2762,N_2877);
xnor UO_323 (O_323,N_2402,N_2504);
xnor UO_324 (O_324,N_2985,N_2645);
and UO_325 (O_325,N_2757,N_2798);
or UO_326 (O_326,N_2580,N_2571);
nor UO_327 (O_327,N_2889,N_2372);
and UO_328 (O_328,N_2478,N_2795);
and UO_329 (O_329,N_2745,N_2347);
xor UO_330 (O_330,N_2491,N_2449);
nand UO_331 (O_331,N_2697,N_2827);
xor UO_332 (O_332,N_2623,N_2573);
nand UO_333 (O_333,N_2852,N_2653);
nand UO_334 (O_334,N_2286,N_2735);
nand UO_335 (O_335,N_2668,N_2346);
or UO_336 (O_336,N_2621,N_2482);
xor UO_337 (O_337,N_2993,N_2335);
xor UO_338 (O_338,N_2931,N_2870);
xnor UO_339 (O_339,N_2435,N_2256);
nand UO_340 (O_340,N_2417,N_2687);
nand UO_341 (O_341,N_2537,N_2432);
xor UO_342 (O_342,N_2529,N_2851);
nand UO_343 (O_343,N_2846,N_2651);
nand UO_344 (O_344,N_2861,N_2394);
and UO_345 (O_345,N_2428,N_2833);
or UO_346 (O_346,N_2465,N_2784);
nor UO_347 (O_347,N_2454,N_2960);
nand UO_348 (O_348,N_2437,N_2338);
and UO_349 (O_349,N_2880,N_2961);
nor UO_350 (O_350,N_2954,N_2460);
or UO_351 (O_351,N_2725,N_2499);
nand UO_352 (O_352,N_2648,N_2740);
or UO_353 (O_353,N_2508,N_2941);
nand UO_354 (O_354,N_2723,N_2310);
nor UO_355 (O_355,N_2517,N_2442);
and UO_356 (O_356,N_2630,N_2672);
or UO_357 (O_357,N_2935,N_2899);
xnor UO_358 (O_358,N_2357,N_2886);
nor UO_359 (O_359,N_2317,N_2513);
and UO_360 (O_360,N_2696,N_2873);
nand UO_361 (O_361,N_2682,N_2754);
and UO_362 (O_362,N_2980,N_2818);
xor UO_363 (O_363,N_2430,N_2882);
or UO_364 (O_364,N_2753,N_2926);
nor UO_365 (O_365,N_2871,N_2856);
and UO_366 (O_366,N_2872,N_2611);
nand UO_367 (O_367,N_2823,N_2259);
nand UO_368 (O_368,N_2526,N_2289);
and UO_369 (O_369,N_2978,N_2384);
nor UO_370 (O_370,N_2492,N_2374);
nand UO_371 (O_371,N_2620,N_2489);
and UO_372 (O_372,N_2689,N_2731);
or UO_373 (O_373,N_2971,N_2930);
and UO_374 (O_374,N_2778,N_2624);
and UO_375 (O_375,N_2516,N_2419);
and UO_376 (O_376,N_2654,N_2720);
nand UO_377 (O_377,N_2583,N_2817);
nand UO_378 (O_378,N_2946,N_2883);
and UO_379 (O_379,N_2971,N_2449);
and UO_380 (O_380,N_2814,N_2340);
nand UO_381 (O_381,N_2483,N_2881);
or UO_382 (O_382,N_2840,N_2602);
and UO_383 (O_383,N_2319,N_2384);
nor UO_384 (O_384,N_2977,N_2494);
and UO_385 (O_385,N_2551,N_2488);
nor UO_386 (O_386,N_2477,N_2890);
or UO_387 (O_387,N_2310,N_2494);
and UO_388 (O_388,N_2327,N_2344);
nor UO_389 (O_389,N_2364,N_2759);
xnor UO_390 (O_390,N_2790,N_2553);
and UO_391 (O_391,N_2833,N_2871);
nor UO_392 (O_392,N_2618,N_2467);
or UO_393 (O_393,N_2287,N_2578);
or UO_394 (O_394,N_2817,N_2910);
or UO_395 (O_395,N_2675,N_2542);
and UO_396 (O_396,N_2588,N_2699);
nor UO_397 (O_397,N_2452,N_2660);
nand UO_398 (O_398,N_2529,N_2517);
nand UO_399 (O_399,N_2431,N_2741);
and UO_400 (O_400,N_2841,N_2787);
xor UO_401 (O_401,N_2673,N_2258);
and UO_402 (O_402,N_2295,N_2625);
or UO_403 (O_403,N_2402,N_2703);
xnor UO_404 (O_404,N_2934,N_2877);
nand UO_405 (O_405,N_2383,N_2335);
and UO_406 (O_406,N_2648,N_2793);
nand UO_407 (O_407,N_2757,N_2389);
nor UO_408 (O_408,N_2439,N_2725);
xnor UO_409 (O_409,N_2870,N_2839);
xor UO_410 (O_410,N_2961,N_2995);
xnor UO_411 (O_411,N_2359,N_2590);
and UO_412 (O_412,N_2511,N_2447);
nand UO_413 (O_413,N_2707,N_2359);
nor UO_414 (O_414,N_2840,N_2731);
xnor UO_415 (O_415,N_2857,N_2684);
nand UO_416 (O_416,N_2847,N_2551);
or UO_417 (O_417,N_2972,N_2872);
nor UO_418 (O_418,N_2616,N_2388);
or UO_419 (O_419,N_2279,N_2827);
and UO_420 (O_420,N_2868,N_2724);
nand UO_421 (O_421,N_2923,N_2864);
nand UO_422 (O_422,N_2618,N_2591);
or UO_423 (O_423,N_2519,N_2655);
or UO_424 (O_424,N_2855,N_2926);
or UO_425 (O_425,N_2739,N_2536);
nor UO_426 (O_426,N_2275,N_2802);
xor UO_427 (O_427,N_2335,N_2947);
nand UO_428 (O_428,N_2914,N_2427);
nand UO_429 (O_429,N_2754,N_2321);
nand UO_430 (O_430,N_2303,N_2754);
nor UO_431 (O_431,N_2442,N_2966);
nand UO_432 (O_432,N_2836,N_2398);
and UO_433 (O_433,N_2724,N_2915);
nand UO_434 (O_434,N_2531,N_2404);
and UO_435 (O_435,N_2439,N_2479);
xnor UO_436 (O_436,N_2362,N_2478);
nand UO_437 (O_437,N_2362,N_2280);
xnor UO_438 (O_438,N_2729,N_2407);
and UO_439 (O_439,N_2867,N_2509);
nand UO_440 (O_440,N_2293,N_2546);
xnor UO_441 (O_441,N_2451,N_2701);
or UO_442 (O_442,N_2775,N_2617);
or UO_443 (O_443,N_2818,N_2289);
nand UO_444 (O_444,N_2596,N_2875);
or UO_445 (O_445,N_2583,N_2862);
or UO_446 (O_446,N_2776,N_2744);
and UO_447 (O_447,N_2837,N_2652);
or UO_448 (O_448,N_2263,N_2606);
or UO_449 (O_449,N_2521,N_2779);
nor UO_450 (O_450,N_2336,N_2797);
nand UO_451 (O_451,N_2604,N_2888);
or UO_452 (O_452,N_2529,N_2283);
or UO_453 (O_453,N_2777,N_2737);
nor UO_454 (O_454,N_2252,N_2886);
nor UO_455 (O_455,N_2461,N_2839);
nor UO_456 (O_456,N_2685,N_2376);
or UO_457 (O_457,N_2773,N_2409);
and UO_458 (O_458,N_2683,N_2387);
or UO_459 (O_459,N_2524,N_2344);
xor UO_460 (O_460,N_2456,N_2516);
or UO_461 (O_461,N_2720,N_2860);
nor UO_462 (O_462,N_2820,N_2437);
nand UO_463 (O_463,N_2686,N_2490);
nor UO_464 (O_464,N_2431,N_2803);
and UO_465 (O_465,N_2993,N_2807);
or UO_466 (O_466,N_2970,N_2459);
and UO_467 (O_467,N_2890,N_2288);
xor UO_468 (O_468,N_2602,N_2695);
nand UO_469 (O_469,N_2309,N_2976);
or UO_470 (O_470,N_2846,N_2432);
nor UO_471 (O_471,N_2599,N_2650);
and UO_472 (O_472,N_2815,N_2886);
or UO_473 (O_473,N_2545,N_2821);
and UO_474 (O_474,N_2542,N_2989);
nand UO_475 (O_475,N_2411,N_2458);
xor UO_476 (O_476,N_2796,N_2763);
nor UO_477 (O_477,N_2514,N_2661);
or UO_478 (O_478,N_2746,N_2540);
nand UO_479 (O_479,N_2999,N_2426);
or UO_480 (O_480,N_2780,N_2823);
nor UO_481 (O_481,N_2940,N_2643);
and UO_482 (O_482,N_2672,N_2927);
nor UO_483 (O_483,N_2746,N_2376);
xnor UO_484 (O_484,N_2335,N_2587);
and UO_485 (O_485,N_2833,N_2567);
nor UO_486 (O_486,N_2696,N_2925);
xor UO_487 (O_487,N_2920,N_2866);
and UO_488 (O_488,N_2316,N_2385);
and UO_489 (O_489,N_2799,N_2734);
and UO_490 (O_490,N_2847,N_2408);
xnor UO_491 (O_491,N_2368,N_2316);
xnor UO_492 (O_492,N_2357,N_2843);
nand UO_493 (O_493,N_2591,N_2543);
nand UO_494 (O_494,N_2460,N_2879);
xor UO_495 (O_495,N_2853,N_2266);
nand UO_496 (O_496,N_2862,N_2799);
nand UO_497 (O_497,N_2793,N_2616);
nor UO_498 (O_498,N_2971,N_2426);
nor UO_499 (O_499,N_2478,N_2604);
endmodule