module basic_1500_15000_2000_5_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_1379,In_69);
xnor U1 (N_1,In_527,In_1235);
nand U2 (N_2,In_498,In_605);
and U3 (N_3,In_1486,In_396);
and U4 (N_4,In_1373,In_613);
xor U5 (N_5,In_583,In_102);
nor U6 (N_6,In_1176,In_129);
nand U7 (N_7,In_1179,In_1416);
nand U8 (N_8,In_1439,In_543);
nand U9 (N_9,In_382,In_112);
and U10 (N_10,In_323,In_161);
and U11 (N_11,In_1436,In_966);
xnor U12 (N_12,In_876,In_1071);
xnor U13 (N_13,In_1277,In_1341);
or U14 (N_14,In_264,In_1150);
or U15 (N_15,In_655,In_89);
nor U16 (N_16,In_813,In_680);
nor U17 (N_17,In_776,In_615);
nor U18 (N_18,In_1295,In_1493);
nand U19 (N_19,In_872,In_538);
xnor U20 (N_20,In_1230,In_1136);
nand U21 (N_21,In_3,In_1325);
nand U22 (N_22,In_1220,In_120);
nor U23 (N_23,In_25,In_508);
xor U24 (N_24,In_104,In_434);
nand U25 (N_25,In_1080,In_1424);
and U26 (N_26,In_331,In_414);
nor U27 (N_27,In_113,In_98);
and U28 (N_28,In_1246,In_921);
or U29 (N_29,In_1254,In_1134);
nor U30 (N_30,In_1426,In_16);
xnor U31 (N_31,In_864,In_784);
or U32 (N_32,In_941,In_79);
or U33 (N_33,In_875,In_729);
and U34 (N_34,In_494,In_339);
and U35 (N_35,In_347,In_656);
nor U36 (N_36,In_74,In_562);
or U37 (N_37,In_885,In_37);
or U38 (N_38,In_1252,In_85);
nand U39 (N_39,In_1314,In_91);
xnor U40 (N_40,In_393,In_915);
or U41 (N_41,In_24,In_1137);
nor U42 (N_42,In_294,In_989);
nor U43 (N_43,In_933,In_718);
or U44 (N_44,In_447,In_327);
xnor U45 (N_45,In_1035,In_883);
nor U46 (N_46,In_525,In_381);
nand U47 (N_47,In_287,In_379);
or U48 (N_48,In_421,In_82);
xor U49 (N_49,In_1072,In_212);
and U50 (N_50,In_131,In_843);
xor U51 (N_51,In_118,In_1093);
xor U52 (N_52,In_550,In_953);
xor U53 (N_53,In_756,In_217);
xnor U54 (N_54,In_874,In_366);
xor U55 (N_55,In_315,In_1343);
xor U56 (N_56,In_677,In_942);
nor U57 (N_57,In_495,In_1479);
xnor U58 (N_58,In_1050,In_894);
or U59 (N_59,In_493,In_1124);
xnor U60 (N_60,In_1132,In_140);
xor U61 (N_61,In_260,In_1);
and U62 (N_62,In_920,In_554);
nor U63 (N_63,In_1077,In_956);
nor U64 (N_64,In_174,In_1318);
and U65 (N_65,In_1172,In_461);
and U66 (N_66,In_302,In_736);
or U67 (N_67,In_547,In_1247);
nor U68 (N_68,In_61,In_1346);
and U69 (N_69,In_1362,In_292);
nand U70 (N_70,In_1123,In_1096);
and U71 (N_71,In_619,In_1218);
nor U72 (N_72,In_228,In_505);
nor U73 (N_73,In_881,In_452);
nand U74 (N_74,In_130,In_1265);
and U75 (N_75,In_202,In_775);
or U76 (N_76,In_857,In_1461);
or U77 (N_77,In_1088,In_93);
or U78 (N_78,In_1180,In_1065);
xor U79 (N_79,In_1239,In_719);
or U80 (N_80,In_1487,In_1342);
and U81 (N_81,In_1385,In_594);
xor U82 (N_82,In_501,In_357);
nand U83 (N_83,In_1192,In_904);
nand U84 (N_84,In_1356,In_472);
xor U85 (N_85,In_1270,In_463);
and U86 (N_86,In_132,In_208);
nor U87 (N_87,In_721,In_570);
and U88 (N_88,In_485,In_895);
nor U89 (N_89,In_53,In_225);
nand U90 (N_90,In_1238,In_1293);
nand U91 (N_91,In_459,In_1211);
and U92 (N_92,In_976,In_1001);
or U93 (N_93,In_1083,In_1060);
and U94 (N_94,In_181,In_281);
and U95 (N_95,In_585,In_175);
nor U96 (N_96,In_936,In_401);
nand U97 (N_97,In_1047,In_246);
xor U98 (N_98,In_710,In_725);
nand U99 (N_99,In_738,In_33);
xor U100 (N_100,In_866,In_320);
xnor U101 (N_101,In_1483,In_67);
nor U102 (N_102,In_362,In_1010);
and U103 (N_103,In_1127,In_180);
nand U104 (N_104,In_1168,In_1320);
nor U105 (N_105,In_18,In_854);
or U106 (N_106,In_961,In_1111);
nor U107 (N_107,In_1337,In_1430);
and U108 (N_108,In_985,In_26);
nand U109 (N_109,In_1437,In_949);
or U110 (N_110,In_253,In_1361);
nor U111 (N_111,In_340,In_659);
or U112 (N_112,In_124,In_963);
nor U113 (N_113,In_544,In_1175);
and U114 (N_114,In_645,In_255);
nand U115 (N_115,In_648,In_449);
nand U116 (N_116,In_766,In_1038);
xor U117 (N_117,In_1201,In_984);
nor U118 (N_118,In_154,In_616);
xnor U119 (N_119,In_43,In_1082);
and U120 (N_120,In_643,In_336);
nor U121 (N_121,In_1100,In_1339);
and U122 (N_122,In_912,In_137);
nor U123 (N_123,In_333,In_1131);
nor U124 (N_124,In_141,In_1244);
xor U125 (N_125,In_670,In_57);
and U126 (N_126,In_997,In_350);
and U127 (N_127,In_1499,In_1425);
xnor U128 (N_128,In_60,In_898);
nand U129 (N_129,In_666,In_1377);
or U130 (N_130,In_1026,In_884);
and U131 (N_131,In_1161,In_367);
and U132 (N_132,In_455,In_54);
nor U133 (N_133,In_924,In_664);
or U134 (N_134,In_669,In_236);
nand U135 (N_135,In_480,In_391);
and U136 (N_136,In_624,In_599);
nand U137 (N_137,In_1368,In_1121);
nand U138 (N_138,In_709,In_1186);
nand U139 (N_139,In_853,In_553);
and U140 (N_140,In_1145,In_1352);
nor U141 (N_141,In_325,In_94);
nand U142 (N_142,In_1375,In_116);
nor U143 (N_143,In_15,In_297);
or U144 (N_144,In_633,In_178);
xnor U145 (N_145,In_798,In_1153);
nand U146 (N_146,In_801,In_380);
or U147 (N_147,In_986,In_695);
nor U148 (N_148,In_1338,In_127);
or U149 (N_149,In_841,In_460);
xnor U150 (N_150,In_417,In_1280);
xnor U151 (N_151,In_652,In_1159);
or U152 (N_152,In_261,In_692);
xnor U153 (N_153,In_809,In_360);
nand U154 (N_154,In_800,In_1422);
and U155 (N_155,In_681,In_403);
nand U156 (N_156,In_309,In_1248);
xor U157 (N_157,In_906,In_319);
or U158 (N_158,In_1146,In_958);
xnor U159 (N_159,In_375,In_560);
nor U160 (N_160,In_1363,In_63);
nor U161 (N_161,In_201,In_774);
and U162 (N_162,In_722,In_780);
nand U163 (N_163,In_858,In_687);
nand U164 (N_164,In_1365,In_926);
or U165 (N_165,In_183,In_781);
nor U166 (N_166,In_303,In_541);
nor U167 (N_167,In_213,In_152);
nand U168 (N_168,In_269,In_579);
and U169 (N_169,In_646,In_611);
xnor U170 (N_170,In_272,In_373);
xnor U171 (N_171,In_828,In_1216);
nor U172 (N_172,In_662,In_405);
nor U173 (N_173,In_757,In_456);
and U174 (N_174,In_172,In_1308);
nand U175 (N_175,In_1200,In_804);
or U176 (N_176,In_1196,In_660);
xor U177 (N_177,In_1138,In_270);
xor U178 (N_178,In_1470,In_932);
nand U179 (N_179,In_1183,In_789);
or U180 (N_180,In_1473,In_374);
nor U181 (N_181,In_531,In_816);
nor U182 (N_182,In_87,In_209);
nor U183 (N_183,In_1208,In_1344);
and U184 (N_184,In_1433,In_1116);
xnor U185 (N_185,In_983,In_995);
or U186 (N_186,In_330,In_160);
nand U187 (N_187,In_610,In_1335);
nand U188 (N_188,In_622,In_337);
or U189 (N_189,In_890,In_1130);
and U190 (N_190,In_1369,In_23);
nor U191 (N_191,In_517,In_909);
nor U192 (N_192,In_1484,In_1383);
or U193 (N_193,In_36,In_574);
nor U194 (N_194,In_1034,In_310);
and U195 (N_195,In_497,In_850);
xor U196 (N_196,In_163,In_749);
and U197 (N_197,In_1427,In_1163);
and U198 (N_198,In_451,In_307);
or U199 (N_199,In_1017,In_1125);
xor U200 (N_200,In_1207,In_1348);
and U201 (N_201,In_457,In_9);
or U202 (N_202,In_1106,In_1197);
nand U203 (N_203,In_1154,In_305);
and U204 (N_204,In_298,In_1457);
nor U205 (N_205,In_833,In_106);
or U206 (N_206,In_454,In_58);
xnor U207 (N_207,In_195,In_601);
nor U208 (N_208,In_1405,In_603);
nand U209 (N_209,In_415,In_581);
or U210 (N_210,In_1476,In_1110);
xor U211 (N_211,In_475,In_723);
xnor U212 (N_212,In_2,In_299);
nor U213 (N_213,In_1070,In_296);
and U214 (N_214,In_1412,In_188);
xnor U215 (N_215,In_1222,In_338);
and U216 (N_216,In_952,In_72);
or U217 (N_217,In_737,In_190);
nor U218 (N_218,In_1284,In_392);
nand U219 (N_219,In_462,In_1241);
and U220 (N_220,In_638,In_68);
and U221 (N_221,In_714,In_470);
xor U222 (N_222,In_930,In_772);
and U223 (N_223,In_1276,In_1481);
or U224 (N_224,In_522,In_675);
xor U225 (N_225,In_1205,In_978);
nand U226 (N_226,In_4,In_1313);
nand U227 (N_227,In_706,In_1144);
nor U228 (N_228,In_777,In_363);
or U229 (N_229,In_618,In_1296);
nor U230 (N_230,In_632,In_1090);
nor U231 (N_231,In_1115,In_1003);
nor U232 (N_232,In_1456,In_623);
nor U233 (N_233,In_487,In_1203);
and U234 (N_234,In_1251,In_827);
nand U235 (N_235,In_234,In_369);
xnor U236 (N_236,In_28,In_1267);
nand U237 (N_237,In_1016,In_192);
or U238 (N_238,In_621,In_489);
or U239 (N_239,In_387,In_849);
and U240 (N_240,In_1051,In_177);
and U241 (N_241,In_734,In_386);
nor U242 (N_242,In_1140,In_1444);
nand U243 (N_243,In_385,In_1411);
xnor U244 (N_244,In_1025,In_464);
xor U245 (N_245,In_661,In_771);
nand U246 (N_246,In_604,In_1471);
xnor U247 (N_247,In_1264,In_759);
nor U248 (N_248,In_262,In_304);
nor U249 (N_249,In_1262,In_1185);
and U250 (N_250,In_1067,In_240);
nand U251 (N_251,In_589,In_1294);
and U252 (N_252,In_1452,In_1249);
and U253 (N_253,In_397,In_101);
and U254 (N_254,In_948,In_561);
nor U255 (N_255,In_38,In_1128);
or U256 (N_256,In_96,In_939);
nor U257 (N_257,In_1255,In_239);
nor U258 (N_258,In_207,In_1417);
and U259 (N_259,In_916,In_1334);
and U260 (N_260,In_640,In_524);
or U261 (N_261,In_1189,In_846);
nor U262 (N_262,In_162,In_422);
xor U263 (N_263,In_861,In_990);
nor U264 (N_264,In_440,In_888);
xor U265 (N_265,In_1206,In_291);
nand U266 (N_266,In_918,In_1434);
or U267 (N_267,In_1122,In_697);
nor U268 (N_268,In_1061,In_443);
xor U269 (N_269,In_1005,In_206);
and U270 (N_270,In_991,In_488);
xnor U271 (N_271,In_1399,In_842);
or U272 (N_272,In_994,In_1073);
xnor U273 (N_273,In_83,In_548);
nor U274 (N_274,In_587,In_755);
or U275 (N_275,In_823,In_1391);
or U276 (N_276,In_769,In_627);
and U277 (N_277,In_50,In_1059);
nor U278 (N_278,In_1287,In_103);
nor U279 (N_279,In_1234,In_165);
xnor U280 (N_280,In_1143,In_418);
nor U281 (N_281,In_753,In_1466);
or U282 (N_282,In_537,In_796);
nor U283 (N_283,In_713,In_532);
nand U284 (N_284,In_1432,In_536);
nand U285 (N_285,In_892,In_150);
xnor U286 (N_286,In_1289,In_256);
nor U287 (N_287,In_609,In_1020);
nor U288 (N_288,In_840,In_1209);
xor U289 (N_289,In_1319,In_215);
xnor U290 (N_290,In_773,In_811);
nor U291 (N_291,In_726,In_1086);
or U292 (N_292,In_1162,In_1429);
and U293 (N_293,In_1353,In_241);
nor U294 (N_294,In_1190,In_896);
nand U295 (N_295,In_1006,In_1312);
xnor U296 (N_296,In_22,In_526);
nor U297 (N_297,In_266,In_179);
nand U298 (N_298,In_221,In_716);
xor U299 (N_299,In_17,In_573);
or U300 (N_300,In_1045,In_1064);
xor U301 (N_301,In_1400,In_1236);
and U302 (N_302,In_1039,In_248);
xnor U303 (N_303,In_1253,In_446);
nand U304 (N_304,In_81,In_184);
and U305 (N_305,In_1380,In_778);
nand U306 (N_306,In_598,In_378);
xnor U307 (N_307,In_1152,In_793);
xnor U308 (N_308,In_84,In_637);
nor U309 (N_309,In_923,In_1087);
nand U310 (N_310,In_332,In_176);
xnor U311 (N_311,In_683,In_1199);
nor U312 (N_312,In_308,In_1257);
nor U313 (N_313,In_419,In_634);
or U314 (N_314,In_913,In_1066);
xor U315 (N_315,In_569,In_1103);
and U316 (N_316,In_186,In_114);
xnor U317 (N_317,In_566,In_1081);
nand U318 (N_318,In_820,In_1445);
nand U319 (N_319,In_824,In_62);
nor U320 (N_320,In_329,In_671);
nor U321 (N_321,In_762,In_530);
or U322 (N_322,In_1193,In_1488);
nor U323 (N_323,In_1024,In_476);
xor U324 (N_324,In_149,In_490);
and U325 (N_325,In_252,In_168);
nor U326 (N_326,In_1108,In_169);
or U327 (N_327,In_258,In_1043);
xor U328 (N_328,In_1421,In_425);
and U329 (N_329,In_1160,In_491);
or U330 (N_330,In_712,In_1158);
and U331 (N_331,In_826,In_1302);
xnor U332 (N_332,In_1403,In_125);
and U333 (N_333,In_1079,In_1184);
and U334 (N_334,In_502,In_156);
nand U335 (N_335,In_705,In_1482);
or U336 (N_336,In_878,In_321);
nand U337 (N_337,In_703,In_159);
xor U338 (N_338,In_1221,In_732);
and U339 (N_339,In_1340,In_819);
xnor U340 (N_340,In_432,In_636);
and U341 (N_341,In_746,In_914);
nand U342 (N_342,In_1177,In_458);
and U343 (N_343,In_650,In_284);
and U344 (N_344,In_1229,In_1101);
nand U345 (N_345,In_1157,In_792);
nor U346 (N_346,In_468,In_1298);
nor U347 (N_347,In_977,In_441);
or U348 (N_348,In_1098,In_35);
and U349 (N_349,In_1495,In_552);
and U350 (N_350,In_1357,In_1392);
and U351 (N_351,In_171,In_748);
or U352 (N_352,In_1360,In_313);
or U353 (N_353,In_1114,In_56);
xor U354 (N_354,In_1394,In_410);
or U355 (N_355,In_249,In_343);
nand U356 (N_356,In_871,In_1268);
and U357 (N_357,In_273,In_741);
nor U358 (N_358,In_880,In_1015);
or U359 (N_359,In_473,In_563);
xor U360 (N_360,In_227,In_1478);
xor U361 (N_361,In_1069,In_251);
nand U362 (N_362,In_514,In_1149);
nor U363 (N_363,In_1260,In_980);
nand U364 (N_364,In_1291,In_546);
xnor U365 (N_365,In_1396,In_197);
and U366 (N_366,In_657,In_973);
nand U367 (N_367,In_1008,In_533);
xnor U368 (N_368,In_334,In_770);
or U369 (N_369,In_198,In_608);
or U370 (N_370,In_1347,In_7);
and U371 (N_371,In_797,In_1300);
or U372 (N_372,In_1258,In_223);
nor U373 (N_373,In_1057,In_612);
or U374 (N_374,In_1384,In_1414);
and U375 (N_375,In_1063,In_1333);
or U376 (N_376,In_1261,In_88);
and U377 (N_377,In_1272,In_1395);
nand U378 (N_378,In_499,In_582);
and U379 (N_379,In_1389,In_504);
and U380 (N_380,In_979,In_1386);
nor U381 (N_381,In_496,In_510);
or U382 (N_382,In_694,In_153);
nand U383 (N_383,In_76,In_1387);
or U384 (N_384,In_607,In_1075);
xnor U385 (N_385,In_651,In_1309);
nor U386 (N_386,In_1037,In_122);
or U387 (N_387,In_1311,In_1465);
or U388 (N_388,In_513,In_803);
nand U389 (N_389,In_500,In_629);
nand U390 (N_390,In_768,In_617);
nor U391 (N_391,In_998,In_193);
and U392 (N_392,In_220,In_21);
nand U393 (N_393,In_14,In_146);
and U394 (N_394,In_735,In_1243);
xor U395 (N_395,In_49,In_1329);
or U396 (N_396,In_1382,In_730);
and U397 (N_397,In_1388,In_185);
and U398 (N_398,In_205,In_1018);
nor U399 (N_399,In_1288,In_571);
xnor U400 (N_400,In_389,In_812);
xor U401 (N_401,In_1301,In_328);
xnor U402 (N_402,In_1279,In_77);
nand U403 (N_403,In_747,In_388);
nand U404 (N_404,In_1012,In_271);
or U405 (N_405,In_862,In_400);
xor U406 (N_406,In_663,In_863);
or U407 (N_407,In_602,In_760);
nand U408 (N_408,In_349,In_565);
nand U409 (N_409,In_1350,In_344);
xnor U410 (N_410,In_967,In_191);
or U411 (N_411,In_1058,In_1195);
nand U412 (N_412,In_635,In_1376);
and U413 (N_413,In_1171,In_1032);
nor U414 (N_414,In_1002,In_1477);
or U415 (N_415,In_242,In_229);
nand U416 (N_416,In_1419,In_1402);
and U417 (N_417,In_71,In_1092);
or U418 (N_418,In_352,In_1263);
nor U419 (N_419,In_224,In_1286);
nor U420 (N_420,In_406,In_1151);
nor U421 (N_421,In_1490,In_844);
and U422 (N_422,In_1463,In_951);
nor U423 (N_423,In_625,In_1046);
and U424 (N_424,In_428,In_549);
nor U425 (N_425,In_1271,In_64);
nor U426 (N_426,In_128,In_216);
nand U427 (N_427,In_744,In_1155);
nand U428 (N_428,In_86,In_518);
nor U429 (N_429,In_483,In_586);
nand U430 (N_430,In_6,In_1187);
xnor U431 (N_431,In_851,In_852);
nand U432 (N_432,In_1278,In_679);
nand U433 (N_433,In_1226,In_593);
nor U434 (N_434,In_1297,In_80);
nand U435 (N_435,In_938,In_1282);
nand U436 (N_436,In_1366,In_658);
xnor U437 (N_437,In_359,In_210);
and U438 (N_438,In_151,In_779);
or U439 (N_439,In_364,In_200);
or U440 (N_440,In_799,In_982);
nand U441 (N_441,In_268,In_384);
or U442 (N_442,In_420,In_109);
nor U443 (N_443,In_427,In_742);
and U444 (N_444,In_503,In_545);
nand U445 (N_445,In_1215,In_996);
or U446 (N_446,In_641,In_477);
xnor U447 (N_447,In_647,In_761);
or U448 (N_448,In_520,In_596);
xor U449 (N_449,In_147,In_48);
and U450 (N_450,In_653,In_1011);
xnor U451 (N_451,In_1242,In_1364);
nor U452 (N_452,In_1213,In_678);
xor U453 (N_453,In_435,In_399);
nand U454 (N_454,In_1450,In_311);
and U455 (N_455,In_971,In_654);
and U456 (N_456,In_821,In_740);
nor U457 (N_457,In_430,In_968);
xor U458 (N_458,In_959,In_155);
and U459 (N_459,In_764,In_572);
xnor U460 (N_460,In_506,In_444);
nand U461 (N_461,In_219,In_232);
and U462 (N_462,In_577,In_211);
and U463 (N_463,In_845,In_542);
xnor U464 (N_464,In_752,In_351);
and U465 (N_465,In_40,In_838);
and U466 (N_466,In_1469,In_1304);
nand U467 (N_467,In_829,In_372);
and U468 (N_468,In_471,In_237);
and U469 (N_469,In_383,In_288);
nand U470 (N_470,In_717,In_1095);
and U471 (N_471,In_1173,In_1397);
or U472 (N_472,In_962,In_1191);
and U473 (N_473,In_196,In_275);
nand U474 (N_474,In_1290,In_47);
nor U475 (N_475,In_157,In_1167);
and U476 (N_476,In_889,In_935);
and U477 (N_477,In_767,In_1409);
xor U478 (N_478,In_204,In_1423);
nor U479 (N_479,In_230,In_317);
or U480 (N_480,In_278,In_1028);
nor U481 (N_481,In_345,In_521);
xnor U482 (N_482,In_606,In_831);
nor U483 (N_483,In_39,In_631);
nand U484 (N_484,In_139,In_535);
xnor U485 (N_485,In_1310,In_1109);
or U486 (N_486,In_672,In_390);
xor U487 (N_487,In_1240,In_0);
or U488 (N_488,In_1198,In_1299);
and U489 (N_489,In_931,In_203);
xnor U490 (N_490,In_859,In_1156);
xnor U491 (N_491,In_754,In_873);
xnor U492 (N_492,In_97,In_1303);
and U493 (N_493,In_368,In_282);
xnor U494 (N_494,In_90,In_1042);
or U495 (N_495,In_274,In_733);
and U496 (N_496,In_466,In_1458);
nand U497 (N_497,In_250,In_1390);
or U498 (N_498,In_233,In_1358);
or U499 (N_499,In_30,In_1327);
xnor U500 (N_500,In_865,In_353);
xor U501 (N_501,In_1027,In_1345);
nand U502 (N_502,In_361,In_1354);
and U503 (N_503,In_1472,In_782);
and U504 (N_504,In_167,In_1322);
or U505 (N_505,In_907,In_126);
and U506 (N_506,In_1381,In_1462);
nor U507 (N_507,In_925,In_887);
and U508 (N_508,In_988,In_45);
nor U509 (N_509,In_115,In_13);
xor U510 (N_510,In_173,In_1494);
and U511 (N_511,In_34,In_1164);
nand U512 (N_512,In_136,In_293);
and U513 (N_513,In_19,In_590);
or U514 (N_514,In_1148,In_954);
nand U515 (N_515,In_1099,In_51);
xnor U516 (N_516,In_856,In_52);
nor U517 (N_517,In_99,In_1074);
nand U518 (N_518,In_992,In_1321);
nand U519 (N_519,In_642,In_684);
nor U520 (N_520,In_591,In_1371);
or U521 (N_521,In_1275,In_512);
xnor U522 (N_522,In_927,In_1431);
and U523 (N_523,In_699,In_515);
or U524 (N_524,In_1440,In_370);
and U525 (N_525,In_704,In_1496);
nand U526 (N_526,In_398,In_1367);
xor U527 (N_527,In_1459,In_969);
and U528 (N_528,In_1355,In_1474);
or U529 (N_529,In_588,In_981);
xor U530 (N_530,In_720,In_1492);
xor U531 (N_531,In_905,In_668);
and U532 (N_532,In_1330,In_715);
xor U533 (N_533,In_688,In_326);
nor U534 (N_534,In_1428,In_194);
nor U535 (N_535,In_133,In_947);
or U536 (N_536,In_1004,In_848);
xnor U537 (N_537,In_453,In_1378);
nand U538 (N_538,In_1233,In_170);
xor U539 (N_539,In_1336,In_1040);
nand U540 (N_540,In_965,In_100);
xor U541 (N_541,In_649,In_791);
or U542 (N_542,In_1129,In_839);
or U543 (N_543,In_867,In_1019);
and U544 (N_544,In_354,In_711);
xor U545 (N_545,In_1491,In_1225);
or U546 (N_546,In_1133,In_869);
nand U547 (N_547,In_832,In_402);
nand U548 (N_548,In_1178,In_745);
and U549 (N_549,In_199,In_1105);
xnor U550 (N_550,In_794,In_847);
xnor U551 (N_551,In_1166,In_231);
and U552 (N_552,In_1307,In_835);
nand U553 (N_553,In_407,In_92);
xor U554 (N_554,In_987,In_1078);
nor U555 (N_555,In_1169,In_807);
and U556 (N_556,In_1374,In_324);
nand U557 (N_557,In_1447,In_119);
or U558 (N_558,In_908,In_928);
nand U559 (N_559,In_117,In_439);
nand U560 (N_560,In_423,In_283);
nor U561 (N_561,In_1489,In_897);
nand U562 (N_562,In_802,In_600);
nand U563 (N_563,In_1041,In_482);
and U564 (N_564,In_817,In_335);
and U565 (N_565,In_408,In_1269);
or U566 (N_566,In_1250,In_576);
nand U567 (N_567,In_1316,In_1455);
nand U568 (N_568,In_960,In_1104);
and U569 (N_569,In_416,In_786);
nor U570 (N_570,In_486,In_42);
and U571 (N_571,In_1210,In_243);
or U572 (N_572,In_810,In_580);
or U573 (N_573,In_1049,In_690);
nor U574 (N_574,In_265,In_424);
nor U575 (N_575,In_20,In_893);
or U576 (N_576,In_882,In_346);
nand U577 (N_577,In_11,In_289);
nand U578 (N_578,In_1062,In_1435);
nor U579 (N_579,In_1231,In_696);
xor U580 (N_580,In_1135,In_999);
nand U581 (N_581,In_479,In_1259);
nand U582 (N_582,In_1285,In_1054);
and U583 (N_583,In_121,In_134);
xor U584 (N_584,In_860,In_693);
and U585 (N_585,In_164,In_944);
xor U586 (N_586,In_1056,In_993);
nand U587 (N_587,In_1076,In_1204);
or U588 (N_588,In_1443,In_280);
nor U589 (N_589,In_342,In_708);
xor U590 (N_590,In_1438,In_682);
or U591 (N_591,In_1256,In_433);
xnor U592 (N_592,In_934,In_822);
nor U593 (N_593,In_1449,In_138);
nor U594 (N_594,In_259,In_1181);
and U595 (N_595,In_787,In_575);
nor U596 (N_596,In_465,In_247);
nand U597 (N_597,In_628,In_65);
nand U598 (N_598,In_111,In_891);
xnor U599 (N_599,In_1141,In_673);
nand U600 (N_600,In_492,In_1227);
nor U601 (N_601,In_1009,In_551);
nor U602 (N_602,In_957,In_442);
xnor U603 (N_603,In_1464,In_1317);
nand U604 (N_604,In_946,In_371);
and U605 (N_605,In_1283,In_66);
nand U606 (N_606,In_1351,In_144);
nor U607 (N_607,In_244,In_970);
xnor U608 (N_608,In_877,In_739);
or U609 (N_609,In_306,In_1044);
or U610 (N_610,In_1188,In_1023);
and U611 (N_611,In_1237,In_855);
nand U612 (N_612,In_724,In_8);
and U613 (N_613,In_1013,In_751);
nor U614 (N_614,In_795,In_376);
or U615 (N_615,In_187,In_1117);
nor U616 (N_616,In_899,In_1091);
or U617 (N_617,In_945,In_301);
and U618 (N_618,In_356,In_701);
and U619 (N_619,In_377,In_1442);
nor U620 (N_620,In_1460,In_676);
nor U621 (N_621,In_1030,In_691);
nand U622 (N_622,In_974,In_1147);
xnor U623 (N_623,In_1052,In_507);
nor U624 (N_624,In_474,In_437);
xor U625 (N_625,In_10,In_630);
nand U626 (N_626,In_917,In_409);
nor U627 (N_627,In_105,In_886);
and U628 (N_628,In_758,In_59);
xnor U629 (N_629,In_1107,In_922);
and U630 (N_630,In_1331,In_1410);
or U631 (N_631,In_300,In_700);
or U632 (N_632,In_818,In_529);
nand U633 (N_633,In_355,In_785);
nor U634 (N_634,In_1393,In_808);
xnor U635 (N_635,In_1332,In_1055);
or U636 (N_636,In_950,In_1126);
xnor U637 (N_637,In_257,In_1033);
xnor U638 (N_638,In_557,In_1228);
xor U639 (N_639,In_41,In_394);
xnor U640 (N_640,In_511,In_44);
xor U641 (N_641,In_1475,In_1468);
nor U642 (N_642,In_834,In_592);
nand U643 (N_643,In_1021,In_1113);
nand U644 (N_644,In_1407,In_900);
nor U645 (N_645,In_1323,In_1142);
and U646 (N_646,In_1182,In_469);
and U647 (N_647,In_290,In_825);
or U648 (N_648,In_1170,In_245);
and U649 (N_649,In_166,In_254);
nand U650 (N_650,In_1454,In_1029);
nand U651 (N_651,In_1446,In_1084);
and U652 (N_652,In_1401,In_235);
xor U653 (N_653,In_75,In_467);
or U654 (N_654,In_830,In_727);
nand U655 (N_655,In_584,In_919);
and U656 (N_656,In_214,In_1217);
xnor U657 (N_657,In_814,In_1418);
nor U658 (N_658,In_667,In_1036);
nand U659 (N_659,In_226,In_1120);
or U660 (N_660,In_1370,In_32);
and U661 (N_661,In_322,In_626);
xor U662 (N_662,In_478,In_55);
and U663 (N_663,In_1408,In_411);
xor U664 (N_664,In_910,In_1219);
and U665 (N_665,In_731,In_1485);
or U666 (N_666,In_27,In_837);
xnor U667 (N_667,In_1031,In_78);
nor U668 (N_668,In_448,In_1328);
or U669 (N_669,In_1118,In_218);
nand U670 (N_670,In_1324,In_312);
nor U671 (N_671,In_1413,In_1224);
nand U672 (N_672,In_1014,In_564);
nor U673 (N_673,In_29,In_689);
nand U674 (N_674,In_445,In_285);
xnor U675 (N_675,In_110,In_901);
or U676 (N_676,In_1451,In_528);
xnor U677 (N_677,In_686,In_805);
xnor U678 (N_678,In_158,In_943);
and U679 (N_679,In_1112,In_836);
or U680 (N_680,In_70,In_578);
xor U681 (N_681,In_1406,In_404);
nand U682 (N_682,In_1048,In_1273);
xnor U683 (N_683,In_238,In_1085);
nor U684 (N_684,In_143,In_426);
nand U685 (N_685,In_107,In_222);
nand U686 (N_686,In_1119,In_595);
nand U687 (N_687,In_964,In_559);
nor U688 (N_688,In_358,In_815);
nor U689 (N_689,In_1000,In_263);
and U690 (N_690,In_509,In_412);
and U691 (N_691,In_556,In_1398);
or U692 (N_692,In_314,In_614);
and U693 (N_693,In_1281,In_879);
or U694 (N_694,In_665,In_702);
or U695 (N_695,In_277,In_1214);
xor U696 (N_696,In_1497,In_558);
nand U697 (N_697,In_431,In_1326);
nor U698 (N_698,In_365,In_911);
nand U699 (N_699,In_728,In_318);
nand U700 (N_700,In_1139,In_620);
or U701 (N_701,In_685,In_123);
nor U702 (N_702,In_267,In_142);
xnor U703 (N_703,In_1467,In_750);
xnor U704 (N_704,In_450,In_108);
nor U705 (N_705,In_148,In_940);
and U706 (N_706,In_972,In_348);
xor U707 (N_707,In_436,In_1349);
nand U708 (N_708,In_189,In_698);
xor U709 (N_709,In_540,In_1305);
nor U710 (N_710,In_1194,In_279);
and U711 (N_711,In_539,In_1202);
or U712 (N_712,In_806,In_1053);
and U713 (N_713,In_1266,In_674);
xor U714 (N_714,In_73,In_868);
or U715 (N_715,In_429,In_765);
nand U716 (N_716,In_567,In_276);
or U717 (N_717,In_286,In_1089);
and U718 (N_718,In_1022,In_1453);
nor U719 (N_719,In_95,In_1448);
and U720 (N_720,In_145,In_31);
or U721 (N_721,In_1404,In_135);
and U722 (N_722,In_903,In_182);
or U723 (N_723,In_788,In_1102);
nor U724 (N_724,In_484,In_1232);
or U725 (N_725,In_1315,In_5);
nand U726 (N_726,In_1441,In_763);
nand U727 (N_727,In_1165,In_975);
nand U728 (N_728,In_1498,In_707);
xnor U729 (N_729,In_395,In_1274);
nand U730 (N_730,In_597,In_1007);
xor U731 (N_731,In_1292,In_12);
or U732 (N_732,In_644,In_295);
xor U733 (N_733,In_955,In_1094);
and U734 (N_734,In_639,In_1306);
or U735 (N_735,In_743,In_519);
nor U736 (N_736,In_516,In_46);
nand U737 (N_737,In_1174,In_438);
nor U738 (N_738,In_1223,In_523);
and U739 (N_739,In_555,In_1245);
nor U740 (N_740,In_481,In_1212);
nor U741 (N_741,In_870,In_316);
nor U742 (N_742,In_341,In_929);
xor U743 (N_743,In_937,In_1068);
nand U744 (N_744,In_1097,In_1415);
or U745 (N_745,In_534,In_902);
nand U746 (N_746,In_783,In_568);
and U747 (N_747,In_1372,In_1480);
xnor U748 (N_748,In_790,In_413);
or U749 (N_749,In_1420,In_1359);
and U750 (N_750,In_1480,In_255);
nand U751 (N_751,In_235,In_538);
nor U752 (N_752,In_1069,In_1058);
xnor U753 (N_753,In_345,In_132);
xor U754 (N_754,In_292,In_576);
and U755 (N_755,In_1495,In_917);
nand U756 (N_756,In_1252,In_1481);
nor U757 (N_757,In_156,In_300);
nand U758 (N_758,In_385,In_669);
and U759 (N_759,In_1482,In_1417);
nor U760 (N_760,In_1172,In_953);
xnor U761 (N_761,In_274,In_898);
or U762 (N_762,In_1032,In_1300);
and U763 (N_763,In_334,In_1278);
and U764 (N_764,In_101,In_544);
xnor U765 (N_765,In_527,In_59);
or U766 (N_766,In_170,In_838);
xor U767 (N_767,In_529,In_269);
or U768 (N_768,In_830,In_112);
xnor U769 (N_769,In_1106,In_1300);
xor U770 (N_770,In_1283,In_922);
nand U771 (N_771,In_651,In_934);
xnor U772 (N_772,In_521,In_532);
and U773 (N_773,In_963,In_832);
xnor U774 (N_774,In_1378,In_743);
or U775 (N_775,In_834,In_1372);
xnor U776 (N_776,In_828,In_525);
or U777 (N_777,In_711,In_1321);
nand U778 (N_778,In_548,In_12);
xor U779 (N_779,In_895,In_84);
and U780 (N_780,In_216,In_790);
and U781 (N_781,In_1487,In_348);
xor U782 (N_782,In_767,In_1015);
and U783 (N_783,In_337,In_441);
and U784 (N_784,In_170,In_28);
or U785 (N_785,In_303,In_424);
or U786 (N_786,In_317,In_1244);
and U787 (N_787,In_592,In_62);
nor U788 (N_788,In_470,In_489);
and U789 (N_789,In_233,In_134);
or U790 (N_790,In_654,In_1275);
nor U791 (N_791,In_848,In_1480);
nor U792 (N_792,In_658,In_972);
and U793 (N_793,In_996,In_1306);
nand U794 (N_794,In_222,In_725);
nor U795 (N_795,In_646,In_1177);
and U796 (N_796,In_1252,In_1078);
nor U797 (N_797,In_1438,In_1263);
and U798 (N_798,In_1195,In_872);
nor U799 (N_799,In_710,In_702);
nand U800 (N_800,In_228,In_1200);
xor U801 (N_801,In_188,In_1185);
xor U802 (N_802,In_1499,In_1094);
nand U803 (N_803,In_978,In_502);
nand U804 (N_804,In_468,In_188);
or U805 (N_805,In_198,In_980);
or U806 (N_806,In_1326,In_609);
or U807 (N_807,In_1408,In_757);
nor U808 (N_808,In_1136,In_668);
xnor U809 (N_809,In_977,In_160);
or U810 (N_810,In_747,In_1064);
nand U811 (N_811,In_251,In_664);
and U812 (N_812,In_1200,In_128);
or U813 (N_813,In_1135,In_756);
nand U814 (N_814,In_1213,In_1070);
and U815 (N_815,In_621,In_749);
xnor U816 (N_816,In_78,In_322);
and U817 (N_817,In_1362,In_1337);
or U818 (N_818,In_192,In_865);
nand U819 (N_819,In_83,In_825);
and U820 (N_820,In_423,In_921);
and U821 (N_821,In_495,In_655);
and U822 (N_822,In_1068,In_83);
or U823 (N_823,In_374,In_206);
or U824 (N_824,In_1190,In_156);
nand U825 (N_825,In_461,In_557);
nand U826 (N_826,In_800,In_1471);
xnor U827 (N_827,In_14,In_1267);
nor U828 (N_828,In_1152,In_1038);
xor U829 (N_829,In_397,In_596);
and U830 (N_830,In_1228,In_396);
nor U831 (N_831,In_1450,In_1492);
nand U832 (N_832,In_244,In_23);
nor U833 (N_833,In_800,In_1147);
xor U834 (N_834,In_243,In_1100);
nand U835 (N_835,In_1003,In_928);
or U836 (N_836,In_1477,In_75);
nor U837 (N_837,In_260,In_216);
nand U838 (N_838,In_307,In_1072);
nand U839 (N_839,In_92,In_1320);
nor U840 (N_840,In_794,In_232);
and U841 (N_841,In_614,In_1390);
nand U842 (N_842,In_59,In_1160);
nand U843 (N_843,In_31,In_476);
nor U844 (N_844,In_725,In_87);
nand U845 (N_845,In_1425,In_833);
nor U846 (N_846,In_292,In_415);
and U847 (N_847,In_1299,In_1260);
xor U848 (N_848,In_146,In_302);
nor U849 (N_849,In_1267,In_1228);
or U850 (N_850,In_993,In_725);
or U851 (N_851,In_1066,In_1044);
nand U852 (N_852,In_588,In_1424);
and U853 (N_853,In_1126,In_587);
and U854 (N_854,In_758,In_1398);
or U855 (N_855,In_547,In_455);
nor U856 (N_856,In_1223,In_1313);
nand U857 (N_857,In_1268,In_1352);
or U858 (N_858,In_677,In_1319);
nor U859 (N_859,In_159,In_1046);
nand U860 (N_860,In_466,In_198);
nand U861 (N_861,In_243,In_1413);
nor U862 (N_862,In_391,In_1033);
nor U863 (N_863,In_598,In_421);
nand U864 (N_864,In_533,In_1346);
xor U865 (N_865,In_316,In_1432);
or U866 (N_866,In_301,In_560);
or U867 (N_867,In_1315,In_755);
or U868 (N_868,In_1068,In_1285);
nand U869 (N_869,In_1041,In_965);
and U870 (N_870,In_1413,In_1339);
or U871 (N_871,In_1045,In_1121);
nand U872 (N_872,In_865,In_77);
nand U873 (N_873,In_1170,In_464);
xnor U874 (N_874,In_1181,In_18);
xnor U875 (N_875,In_960,In_556);
nand U876 (N_876,In_360,In_846);
nor U877 (N_877,In_1111,In_771);
nand U878 (N_878,In_60,In_572);
xnor U879 (N_879,In_943,In_1028);
nand U880 (N_880,In_1194,In_702);
and U881 (N_881,In_657,In_669);
nor U882 (N_882,In_257,In_910);
xnor U883 (N_883,In_924,In_1484);
nand U884 (N_884,In_1152,In_406);
or U885 (N_885,In_1214,In_901);
nand U886 (N_886,In_1236,In_742);
or U887 (N_887,In_1376,In_1279);
and U888 (N_888,In_469,In_319);
and U889 (N_889,In_169,In_1081);
and U890 (N_890,In_629,In_1188);
nand U891 (N_891,In_1353,In_633);
xnor U892 (N_892,In_381,In_204);
nor U893 (N_893,In_1040,In_714);
nand U894 (N_894,In_149,In_1241);
nand U895 (N_895,In_496,In_1155);
nor U896 (N_896,In_209,In_1109);
and U897 (N_897,In_352,In_1328);
or U898 (N_898,In_1058,In_1205);
nand U899 (N_899,In_482,In_667);
or U900 (N_900,In_595,In_1491);
and U901 (N_901,In_1283,In_1144);
xnor U902 (N_902,In_652,In_1494);
xor U903 (N_903,In_1397,In_1455);
and U904 (N_904,In_398,In_78);
or U905 (N_905,In_140,In_819);
or U906 (N_906,In_403,In_832);
xor U907 (N_907,In_386,In_1060);
xnor U908 (N_908,In_1368,In_1355);
nand U909 (N_909,In_1123,In_1363);
nor U910 (N_910,In_1474,In_796);
or U911 (N_911,In_94,In_164);
nand U912 (N_912,In_1387,In_182);
nand U913 (N_913,In_973,In_1160);
nor U914 (N_914,In_204,In_361);
and U915 (N_915,In_1167,In_60);
xnor U916 (N_916,In_843,In_887);
xor U917 (N_917,In_659,In_440);
or U918 (N_918,In_464,In_890);
nand U919 (N_919,In_1358,In_1051);
nand U920 (N_920,In_1154,In_679);
and U921 (N_921,In_1180,In_747);
nor U922 (N_922,In_765,In_255);
or U923 (N_923,In_1336,In_1082);
xor U924 (N_924,In_250,In_62);
nand U925 (N_925,In_173,In_648);
and U926 (N_926,In_547,In_422);
nor U927 (N_927,In_384,In_748);
xnor U928 (N_928,In_1422,In_349);
xnor U929 (N_929,In_572,In_1458);
or U930 (N_930,In_17,In_498);
nor U931 (N_931,In_1332,In_1095);
and U932 (N_932,In_401,In_895);
and U933 (N_933,In_904,In_150);
nor U934 (N_934,In_249,In_1256);
or U935 (N_935,In_1038,In_475);
xor U936 (N_936,In_167,In_26);
nor U937 (N_937,In_1357,In_1476);
or U938 (N_938,In_556,In_1174);
or U939 (N_939,In_1019,In_1135);
xnor U940 (N_940,In_1345,In_1484);
and U941 (N_941,In_1119,In_743);
nand U942 (N_942,In_881,In_1390);
nand U943 (N_943,In_1457,In_1358);
nand U944 (N_944,In_1056,In_167);
and U945 (N_945,In_275,In_106);
xor U946 (N_946,In_1466,In_1207);
xnor U947 (N_947,In_841,In_87);
or U948 (N_948,In_55,In_362);
nor U949 (N_949,In_1438,In_562);
xor U950 (N_950,In_1142,In_34);
nor U951 (N_951,In_817,In_1438);
nor U952 (N_952,In_1241,In_321);
and U953 (N_953,In_1096,In_478);
nor U954 (N_954,In_280,In_1402);
or U955 (N_955,In_1023,In_32);
nor U956 (N_956,In_1283,In_452);
or U957 (N_957,In_1115,In_479);
nor U958 (N_958,In_88,In_61);
or U959 (N_959,In_496,In_438);
and U960 (N_960,In_1098,In_413);
and U961 (N_961,In_1496,In_1247);
or U962 (N_962,In_904,In_558);
and U963 (N_963,In_70,In_843);
xnor U964 (N_964,In_1469,In_1471);
nor U965 (N_965,In_331,In_870);
nor U966 (N_966,In_1314,In_776);
nor U967 (N_967,In_1203,In_1419);
and U968 (N_968,In_705,In_847);
or U969 (N_969,In_831,In_399);
or U970 (N_970,In_606,In_1089);
nand U971 (N_971,In_875,In_1095);
xor U972 (N_972,In_1058,In_803);
nor U973 (N_973,In_415,In_1453);
nand U974 (N_974,In_1450,In_771);
xnor U975 (N_975,In_193,In_265);
and U976 (N_976,In_910,In_471);
and U977 (N_977,In_595,In_594);
nand U978 (N_978,In_615,In_1493);
nand U979 (N_979,In_110,In_858);
xnor U980 (N_980,In_2,In_53);
xnor U981 (N_981,In_1141,In_1173);
and U982 (N_982,In_1189,In_688);
xnor U983 (N_983,In_729,In_789);
or U984 (N_984,In_1266,In_1138);
and U985 (N_985,In_732,In_1095);
and U986 (N_986,In_336,In_1407);
or U987 (N_987,In_428,In_946);
nand U988 (N_988,In_770,In_809);
or U989 (N_989,In_1083,In_1319);
and U990 (N_990,In_1341,In_1217);
nor U991 (N_991,In_363,In_385);
or U992 (N_992,In_902,In_1124);
xor U993 (N_993,In_192,In_1339);
or U994 (N_994,In_644,In_1491);
xnor U995 (N_995,In_789,In_1325);
nand U996 (N_996,In_1021,In_905);
or U997 (N_997,In_810,In_386);
or U998 (N_998,In_1369,In_756);
or U999 (N_999,In_1368,In_547);
nand U1000 (N_1000,In_1409,In_921);
or U1001 (N_1001,In_434,In_396);
nand U1002 (N_1002,In_350,In_1200);
or U1003 (N_1003,In_942,In_1066);
nor U1004 (N_1004,In_765,In_395);
and U1005 (N_1005,In_1031,In_675);
xnor U1006 (N_1006,In_197,In_760);
nand U1007 (N_1007,In_1148,In_628);
and U1008 (N_1008,In_912,In_483);
and U1009 (N_1009,In_1342,In_765);
nand U1010 (N_1010,In_301,In_908);
xnor U1011 (N_1011,In_533,In_33);
xor U1012 (N_1012,In_850,In_915);
or U1013 (N_1013,In_350,In_930);
or U1014 (N_1014,In_1273,In_251);
xor U1015 (N_1015,In_1388,In_524);
xor U1016 (N_1016,In_322,In_1137);
and U1017 (N_1017,In_554,In_240);
and U1018 (N_1018,In_1126,In_1104);
xnor U1019 (N_1019,In_744,In_806);
xnor U1020 (N_1020,In_1301,In_1368);
xnor U1021 (N_1021,In_462,In_220);
or U1022 (N_1022,In_541,In_644);
nor U1023 (N_1023,In_1488,In_491);
or U1024 (N_1024,In_1315,In_402);
and U1025 (N_1025,In_1140,In_909);
or U1026 (N_1026,In_1495,In_233);
xnor U1027 (N_1027,In_631,In_1434);
xor U1028 (N_1028,In_757,In_902);
and U1029 (N_1029,In_1105,In_410);
or U1030 (N_1030,In_1203,In_1243);
nand U1031 (N_1031,In_1316,In_989);
xor U1032 (N_1032,In_1406,In_1385);
nor U1033 (N_1033,In_643,In_1431);
nor U1034 (N_1034,In_124,In_101);
nor U1035 (N_1035,In_216,In_1423);
or U1036 (N_1036,In_670,In_1312);
xnor U1037 (N_1037,In_439,In_685);
or U1038 (N_1038,In_86,In_851);
xnor U1039 (N_1039,In_1110,In_1402);
xnor U1040 (N_1040,In_1062,In_180);
and U1041 (N_1041,In_626,In_1451);
or U1042 (N_1042,In_556,In_664);
nor U1043 (N_1043,In_345,In_1139);
nand U1044 (N_1044,In_1335,In_215);
or U1045 (N_1045,In_462,In_235);
or U1046 (N_1046,In_629,In_204);
nand U1047 (N_1047,In_248,In_535);
and U1048 (N_1048,In_1126,In_210);
or U1049 (N_1049,In_317,In_797);
or U1050 (N_1050,In_1381,In_61);
xnor U1051 (N_1051,In_828,In_139);
nand U1052 (N_1052,In_880,In_1499);
nand U1053 (N_1053,In_1457,In_1361);
and U1054 (N_1054,In_155,In_1411);
nor U1055 (N_1055,In_1290,In_837);
nand U1056 (N_1056,In_1109,In_762);
or U1057 (N_1057,In_1338,In_851);
nor U1058 (N_1058,In_836,In_1252);
xnor U1059 (N_1059,In_768,In_475);
and U1060 (N_1060,In_1422,In_1293);
xor U1061 (N_1061,In_192,In_46);
nand U1062 (N_1062,In_658,In_140);
nor U1063 (N_1063,In_4,In_1040);
nand U1064 (N_1064,In_1407,In_542);
nand U1065 (N_1065,In_1111,In_725);
xnor U1066 (N_1066,In_282,In_1028);
nand U1067 (N_1067,In_706,In_198);
nor U1068 (N_1068,In_180,In_1122);
nand U1069 (N_1069,In_1428,In_1184);
or U1070 (N_1070,In_838,In_1138);
nor U1071 (N_1071,In_345,In_1098);
or U1072 (N_1072,In_724,In_559);
nand U1073 (N_1073,In_612,In_228);
nand U1074 (N_1074,In_25,In_1237);
and U1075 (N_1075,In_1160,In_57);
and U1076 (N_1076,In_387,In_379);
xnor U1077 (N_1077,In_566,In_1008);
nor U1078 (N_1078,In_765,In_59);
or U1079 (N_1079,In_637,In_1369);
and U1080 (N_1080,In_791,In_1138);
and U1081 (N_1081,In_654,In_70);
xor U1082 (N_1082,In_631,In_472);
nand U1083 (N_1083,In_66,In_1318);
or U1084 (N_1084,In_739,In_597);
xor U1085 (N_1085,In_669,In_1438);
and U1086 (N_1086,In_649,In_984);
or U1087 (N_1087,In_598,In_968);
nand U1088 (N_1088,In_1415,In_3);
xor U1089 (N_1089,In_610,In_1140);
nand U1090 (N_1090,In_1303,In_655);
nand U1091 (N_1091,In_397,In_159);
or U1092 (N_1092,In_1020,In_1280);
or U1093 (N_1093,In_932,In_621);
nand U1094 (N_1094,In_1496,In_1145);
nand U1095 (N_1095,In_1387,In_558);
nor U1096 (N_1096,In_1057,In_1192);
nand U1097 (N_1097,In_955,In_802);
and U1098 (N_1098,In_1474,In_429);
nand U1099 (N_1099,In_106,In_168);
nor U1100 (N_1100,In_1284,In_183);
and U1101 (N_1101,In_1266,In_114);
nor U1102 (N_1102,In_345,In_856);
xnor U1103 (N_1103,In_199,In_1492);
or U1104 (N_1104,In_1279,In_584);
nand U1105 (N_1105,In_395,In_490);
or U1106 (N_1106,In_1177,In_218);
nand U1107 (N_1107,In_1189,In_512);
xnor U1108 (N_1108,In_358,In_1135);
and U1109 (N_1109,In_725,In_31);
nand U1110 (N_1110,In_907,In_673);
xor U1111 (N_1111,In_1310,In_1308);
nand U1112 (N_1112,In_1377,In_1054);
xnor U1113 (N_1113,In_184,In_1235);
or U1114 (N_1114,In_1487,In_1255);
or U1115 (N_1115,In_492,In_487);
nand U1116 (N_1116,In_1186,In_504);
nand U1117 (N_1117,In_641,In_388);
nand U1118 (N_1118,In_179,In_849);
nand U1119 (N_1119,In_727,In_1081);
or U1120 (N_1120,In_420,In_1445);
or U1121 (N_1121,In_676,In_181);
or U1122 (N_1122,In_385,In_354);
xnor U1123 (N_1123,In_746,In_116);
nand U1124 (N_1124,In_629,In_539);
or U1125 (N_1125,In_1188,In_1311);
nor U1126 (N_1126,In_668,In_1138);
or U1127 (N_1127,In_1322,In_760);
nor U1128 (N_1128,In_52,In_1432);
or U1129 (N_1129,In_1162,In_1325);
and U1130 (N_1130,In_122,In_334);
or U1131 (N_1131,In_665,In_865);
or U1132 (N_1132,In_511,In_567);
and U1133 (N_1133,In_1344,In_375);
nand U1134 (N_1134,In_757,In_556);
nand U1135 (N_1135,In_950,In_1475);
xor U1136 (N_1136,In_406,In_95);
and U1137 (N_1137,In_1453,In_468);
xnor U1138 (N_1138,In_9,In_359);
and U1139 (N_1139,In_461,In_555);
nor U1140 (N_1140,In_435,In_1153);
or U1141 (N_1141,In_776,In_343);
xor U1142 (N_1142,In_160,In_1313);
xor U1143 (N_1143,In_1432,In_415);
xnor U1144 (N_1144,In_1030,In_54);
xor U1145 (N_1145,In_786,In_1051);
nor U1146 (N_1146,In_11,In_83);
nor U1147 (N_1147,In_1017,In_511);
xnor U1148 (N_1148,In_1454,In_1461);
nor U1149 (N_1149,In_180,In_1353);
or U1150 (N_1150,In_1385,In_360);
and U1151 (N_1151,In_959,In_1146);
nor U1152 (N_1152,In_1097,In_585);
nand U1153 (N_1153,In_848,In_390);
nand U1154 (N_1154,In_116,In_721);
or U1155 (N_1155,In_770,In_1400);
xor U1156 (N_1156,In_745,In_999);
xnor U1157 (N_1157,In_1074,In_85);
xor U1158 (N_1158,In_1163,In_1355);
nand U1159 (N_1159,In_278,In_353);
nor U1160 (N_1160,In_838,In_1267);
nor U1161 (N_1161,In_981,In_357);
nor U1162 (N_1162,In_814,In_1069);
nand U1163 (N_1163,In_237,In_663);
and U1164 (N_1164,In_402,In_856);
nor U1165 (N_1165,In_1455,In_79);
xnor U1166 (N_1166,In_1315,In_1269);
nor U1167 (N_1167,In_499,In_1170);
nor U1168 (N_1168,In_1064,In_829);
and U1169 (N_1169,In_76,In_1250);
or U1170 (N_1170,In_1029,In_568);
or U1171 (N_1171,In_247,In_1302);
nand U1172 (N_1172,In_362,In_50);
xor U1173 (N_1173,In_95,In_343);
nor U1174 (N_1174,In_64,In_1396);
nand U1175 (N_1175,In_1287,In_88);
nand U1176 (N_1176,In_1169,In_1302);
or U1177 (N_1177,In_635,In_176);
or U1178 (N_1178,In_365,In_1375);
xor U1179 (N_1179,In_597,In_38);
nand U1180 (N_1180,In_974,In_129);
and U1181 (N_1181,In_77,In_1112);
or U1182 (N_1182,In_447,In_1021);
nor U1183 (N_1183,In_568,In_83);
nand U1184 (N_1184,In_314,In_951);
xor U1185 (N_1185,In_648,In_627);
or U1186 (N_1186,In_1492,In_1152);
xor U1187 (N_1187,In_1243,In_1076);
and U1188 (N_1188,In_1197,In_100);
nor U1189 (N_1189,In_842,In_1302);
nand U1190 (N_1190,In_1363,In_837);
and U1191 (N_1191,In_1197,In_179);
xor U1192 (N_1192,In_135,In_1176);
xnor U1193 (N_1193,In_1464,In_174);
xor U1194 (N_1194,In_1234,In_284);
nor U1195 (N_1195,In_1260,In_312);
xnor U1196 (N_1196,In_29,In_735);
or U1197 (N_1197,In_714,In_1404);
nand U1198 (N_1198,In_916,In_197);
nand U1199 (N_1199,In_830,In_1288);
or U1200 (N_1200,In_420,In_391);
xnor U1201 (N_1201,In_83,In_250);
and U1202 (N_1202,In_30,In_921);
or U1203 (N_1203,In_1377,In_726);
or U1204 (N_1204,In_1058,In_793);
and U1205 (N_1205,In_1287,In_681);
nor U1206 (N_1206,In_1162,In_1493);
and U1207 (N_1207,In_1219,In_234);
and U1208 (N_1208,In_447,In_1358);
nand U1209 (N_1209,In_1315,In_1021);
or U1210 (N_1210,In_608,In_461);
nand U1211 (N_1211,In_226,In_1367);
nand U1212 (N_1212,In_1067,In_1287);
nor U1213 (N_1213,In_606,In_1041);
nand U1214 (N_1214,In_149,In_548);
xnor U1215 (N_1215,In_1032,In_236);
and U1216 (N_1216,In_695,In_1060);
and U1217 (N_1217,In_921,In_475);
and U1218 (N_1218,In_1032,In_882);
and U1219 (N_1219,In_1237,In_1102);
xnor U1220 (N_1220,In_297,In_615);
nand U1221 (N_1221,In_136,In_432);
and U1222 (N_1222,In_290,In_774);
nor U1223 (N_1223,In_947,In_211);
xor U1224 (N_1224,In_599,In_113);
or U1225 (N_1225,In_702,In_622);
xor U1226 (N_1226,In_255,In_868);
nand U1227 (N_1227,In_1213,In_165);
xor U1228 (N_1228,In_35,In_436);
or U1229 (N_1229,In_1298,In_239);
or U1230 (N_1230,In_299,In_1269);
and U1231 (N_1231,In_672,In_1273);
nand U1232 (N_1232,In_782,In_458);
nor U1233 (N_1233,In_158,In_1295);
or U1234 (N_1234,In_1166,In_63);
or U1235 (N_1235,In_1192,In_332);
nor U1236 (N_1236,In_211,In_1342);
nor U1237 (N_1237,In_36,In_369);
nor U1238 (N_1238,In_153,In_1303);
nand U1239 (N_1239,In_553,In_940);
xor U1240 (N_1240,In_480,In_1471);
nand U1241 (N_1241,In_460,In_998);
nor U1242 (N_1242,In_933,In_888);
or U1243 (N_1243,In_24,In_153);
nor U1244 (N_1244,In_98,In_1284);
nand U1245 (N_1245,In_844,In_1413);
nor U1246 (N_1246,In_715,In_1220);
nand U1247 (N_1247,In_98,In_49);
or U1248 (N_1248,In_822,In_337);
or U1249 (N_1249,In_1303,In_281);
nand U1250 (N_1250,In_145,In_650);
xor U1251 (N_1251,In_1408,In_980);
nor U1252 (N_1252,In_1116,In_530);
and U1253 (N_1253,In_166,In_595);
nor U1254 (N_1254,In_773,In_358);
nand U1255 (N_1255,In_262,In_979);
nor U1256 (N_1256,In_1109,In_880);
xnor U1257 (N_1257,In_934,In_898);
or U1258 (N_1258,In_598,In_217);
xor U1259 (N_1259,In_1444,In_240);
and U1260 (N_1260,In_1191,In_881);
or U1261 (N_1261,In_1054,In_718);
or U1262 (N_1262,In_247,In_1349);
and U1263 (N_1263,In_1222,In_1159);
and U1264 (N_1264,In_0,In_310);
xnor U1265 (N_1265,In_244,In_716);
xor U1266 (N_1266,In_1081,In_1478);
nor U1267 (N_1267,In_1098,In_589);
and U1268 (N_1268,In_977,In_827);
nand U1269 (N_1269,In_926,In_210);
and U1270 (N_1270,In_617,In_1216);
nand U1271 (N_1271,In_926,In_1486);
or U1272 (N_1272,In_1310,In_1174);
nor U1273 (N_1273,In_1352,In_1096);
or U1274 (N_1274,In_1316,In_744);
nand U1275 (N_1275,In_90,In_295);
nand U1276 (N_1276,In_1210,In_399);
xnor U1277 (N_1277,In_259,In_197);
xor U1278 (N_1278,In_1198,In_319);
nor U1279 (N_1279,In_494,In_1016);
nor U1280 (N_1280,In_732,In_1456);
xor U1281 (N_1281,In_837,In_496);
nand U1282 (N_1282,In_634,In_475);
nor U1283 (N_1283,In_758,In_1154);
or U1284 (N_1284,In_893,In_121);
or U1285 (N_1285,In_292,In_879);
and U1286 (N_1286,In_266,In_427);
nor U1287 (N_1287,In_37,In_332);
and U1288 (N_1288,In_822,In_1365);
and U1289 (N_1289,In_672,In_1200);
and U1290 (N_1290,In_105,In_421);
or U1291 (N_1291,In_1004,In_865);
xor U1292 (N_1292,In_1300,In_1124);
or U1293 (N_1293,In_979,In_873);
xnor U1294 (N_1294,In_647,In_427);
nor U1295 (N_1295,In_1052,In_1476);
and U1296 (N_1296,In_936,In_1268);
nor U1297 (N_1297,In_1453,In_1289);
or U1298 (N_1298,In_433,In_894);
nand U1299 (N_1299,In_119,In_63);
or U1300 (N_1300,In_222,In_585);
or U1301 (N_1301,In_1247,In_1364);
or U1302 (N_1302,In_100,In_449);
nand U1303 (N_1303,In_787,In_764);
nand U1304 (N_1304,In_1454,In_142);
nor U1305 (N_1305,In_1053,In_669);
xnor U1306 (N_1306,In_271,In_122);
and U1307 (N_1307,In_616,In_251);
nand U1308 (N_1308,In_1018,In_292);
nand U1309 (N_1309,In_1480,In_422);
or U1310 (N_1310,In_401,In_190);
nor U1311 (N_1311,In_92,In_613);
nor U1312 (N_1312,In_657,In_295);
and U1313 (N_1313,In_1134,In_524);
and U1314 (N_1314,In_927,In_598);
and U1315 (N_1315,In_549,In_249);
nand U1316 (N_1316,In_1387,In_406);
nor U1317 (N_1317,In_814,In_847);
xnor U1318 (N_1318,In_1123,In_293);
and U1319 (N_1319,In_1128,In_421);
nor U1320 (N_1320,In_798,In_982);
nor U1321 (N_1321,In_155,In_711);
or U1322 (N_1322,In_1160,In_877);
xor U1323 (N_1323,In_383,In_281);
nand U1324 (N_1324,In_683,In_397);
xor U1325 (N_1325,In_1224,In_598);
or U1326 (N_1326,In_515,In_1344);
nand U1327 (N_1327,In_1007,In_1177);
nand U1328 (N_1328,In_1343,In_45);
nor U1329 (N_1329,In_1027,In_794);
and U1330 (N_1330,In_447,In_830);
or U1331 (N_1331,In_584,In_1322);
nand U1332 (N_1332,In_850,In_86);
xor U1333 (N_1333,In_1459,In_1257);
nand U1334 (N_1334,In_812,In_1228);
and U1335 (N_1335,In_589,In_620);
xor U1336 (N_1336,In_1324,In_728);
or U1337 (N_1337,In_424,In_1450);
xor U1338 (N_1338,In_197,In_789);
nand U1339 (N_1339,In_1422,In_1489);
and U1340 (N_1340,In_1496,In_823);
xnor U1341 (N_1341,In_322,In_340);
and U1342 (N_1342,In_1046,In_1347);
and U1343 (N_1343,In_1060,In_1099);
or U1344 (N_1344,In_526,In_1164);
or U1345 (N_1345,In_865,In_959);
nor U1346 (N_1346,In_976,In_582);
and U1347 (N_1347,In_1136,In_73);
and U1348 (N_1348,In_1458,In_867);
nor U1349 (N_1349,In_1097,In_1182);
or U1350 (N_1350,In_58,In_1274);
nor U1351 (N_1351,In_912,In_478);
or U1352 (N_1352,In_1418,In_575);
and U1353 (N_1353,In_190,In_371);
nand U1354 (N_1354,In_1351,In_333);
and U1355 (N_1355,In_1047,In_1059);
nand U1356 (N_1356,In_111,In_205);
xnor U1357 (N_1357,In_1368,In_1064);
nand U1358 (N_1358,In_920,In_146);
nand U1359 (N_1359,In_12,In_977);
nand U1360 (N_1360,In_219,In_94);
nor U1361 (N_1361,In_991,In_330);
xor U1362 (N_1362,In_343,In_1194);
nor U1363 (N_1363,In_45,In_1394);
xor U1364 (N_1364,In_220,In_820);
xor U1365 (N_1365,In_1308,In_1396);
nand U1366 (N_1366,In_209,In_752);
nand U1367 (N_1367,In_807,In_1396);
nor U1368 (N_1368,In_1310,In_1255);
and U1369 (N_1369,In_731,In_1360);
and U1370 (N_1370,In_231,In_865);
xor U1371 (N_1371,In_417,In_624);
xor U1372 (N_1372,In_794,In_1323);
or U1373 (N_1373,In_293,In_836);
and U1374 (N_1374,In_284,In_296);
nor U1375 (N_1375,In_919,In_1338);
nor U1376 (N_1376,In_878,In_375);
and U1377 (N_1377,In_377,In_310);
xor U1378 (N_1378,In_26,In_954);
xnor U1379 (N_1379,In_405,In_849);
or U1380 (N_1380,In_1292,In_591);
and U1381 (N_1381,In_980,In_1361);
nand U1382 (N_1382,In_17,In_1058);
and U1383 (N_1383,In_1256,In_1074);
xnor U1384 (N_1384,In_1447,In_1210);
nor U1385 (N_1385,In_573,In_247);
xor U1386 (N_1386,In_1397,In_357);
nand U1387 (N_1387,In_1031,In_772);
nand U1388 (N_1388,In_843,In_1210);
nor U1389 (N_1389,In_867,In_662);
and U1390 (N_1390,In_613,In_781);
or U1391 (N_1391,In_179,In_544);
or U1392 (N_1392,In_9,In_181);
nor U1393 (N_1393,In_364,In_850);
and U1394 (N_1394,In_109,In_1086);
and U1395 (N_1395,In_228,In_480);
nand U1396 (N_1396,In_174,In_558);
xor U1397 (N_1397,In_848,In_1086);
or U1398 (N_1398,In_24,In_279);
and U1399 (N_1399,In_593,In_289);
and U1400 (N_1400,In_894,In_1047);
xnor U1401 (N_1401,In_430,In_1320);
xor U1402 (N_1402,In_1426,In_420);
or U1403 (N_1403,In_461,In_504);
and U1404 (N_1404,In_928,In_674);
nand U1405 (N_1405,In_1446,In_898);
nand U1406 (N_1406,In_47,In_526);
and U1407 (N_1407,In_314,In_550);
or U1408 (N_1408,In_1316,In_983);
xnor U1409 (N_1409,In_78,In_242);
xor U1410 (N_1410,In_1360,In_387);
or U1411 (N_1411,In_421,In_766);
nand U1412 (N_1412,In_156,In_827);
nor U1413 (N_1413,In_356,In_480);
or U1414 (N_1414,In_1037,In_1242);
nor U1415 (N_1415,In_822,In_1206);
nand U1416 (N_1416,In_1280,In_1123);
xnor U1417 (N_1417,In_898,In_163);
nand U1418 (N_1418,In_1019,In_1013);
nand U1419 (N_1419,In_213,In_257);
nand U1420 (N_1420,In_91,In_1284);
and U1421 (N_1421,In_918,In_780);
and U1422 (N_1422,In_250,In_467);
or U1423 (N_1423,In_519,In_814);
or U1424 (N_1424,In_600,In_1074);
xnor U1425 (N_1425,In_6,In_946);
xnor U1426 (N_1426,In_1452,In_167);
xor U1427 (N_1427,In_156,In_833);
nor U1428 (N_1428,In_97,In_569);
nor U1429 (N_1429,In_729,In_773);
nand U1430 (N_1430,In_1470,In_1147);
nand U1431 (N_1431,In_5,In_130);
or U1432 (N_1432,In_307,In_982);
nand U1433 (N_1433,In_437,In_336);
and U1434 (N_1434,In_196,In_187);
nand U1435 (N_1435,In_596,In_1203);
nand U1436 (N_1436,In_596,In_1268);
nor U1437 (N_1437,In_267,In_187);
and U1438 (N_1438,In_926,In_61);
or U1439 (N_1439,In_598,In_1050);
nand U1440 (N_1440,In_1095,In_1097);
and U1441 (N_1441,In_215,In_893);
nor U1442 (N_1442,In_1079,In_913);
nor U1443 (N_1443,In_964,In_1272);
nor U1444 (N_1444,In_4,In_227);
nand U1445 (N_1445,In_866,In_619);
nor U1446 (N_1446,In_15,In_788);
or U1447 (N_1447,In_395,In_413);
and U1448 (N_1448,In_791,In_1401);
xor U1449 (N_1449,In_1214,In_898);
nand U1450 (N_1450,In_355,In_1218);
and U1451 (N_1451,In_1158,In_915);
or U1452 (N_1452,In_870,In_845);
nand U1453 (N_1453,In_1366,In_871);
or U1454 (N_1454,In_454,In_146);
xnor U1455 (N_1455,In_1306,In_594);
xor U1456 (N_1456,In_611,In_378);
or U1457 (N_1457,In_1114,In_1402);
xor U1458 (N_1458,In_829,In_1340);
nor U1459 (N_1459,In_1390,In_1248);
nor U1460 (N_1460,In_1361,In_351);
nand U1461 (N_1461,In_430,In_1495);
xor U1462 (N_1462,In_989,In_225);
nor U1463 (N_1463,In_305,In_152);
nand U1464 (N_1464,In_392,In_1432);
nand U1465 (N_1465,In_345,In_1328);
nor U1466 (N_1466,In_1032,In_852);
nor U1467 (N_1467,In_450,In_691);
nand U1468 (N_1468,In_602,In_1110);
or U1469 (N_1469,In_688,In_794);
or U1470 (N_1470,In_1328,In_644);
and U1471 (N_1471,In_243,In_220);
nor U1472 (N_1472,In_890,In_460);
nor U1473 (N_1473,In_769,In_545);
xnor U1474 (N_1474,In_708,In_733);
or U1475 (N_1475,In_359,In_844);
xor U1476 (N_1476,In_304,In_827);
nand U1477 (N_1477,In_630,In_460);
xor U1478 (N_1478,In_472,In_1455);
and U1479 (N_1479,In_1155,In_516);
xnor U1480 (N_1480,In_766,In_1363);
or U1481 (N_1481,In_369,In_1247);
and U1482 (N_1482,In_1421,In_738);
and U1483 (N_1483,In_216,In_1144);
xor U1484 (N_1484,In_318,In_171);
nand U1485 (N_1485,In_139,In_860);
and U1486 (N_1486,In_1211,In_1166);
or U1487 (N_1487,In_691,In_429);
xnor U1488 (N_1488,In_190,In_38);
nor U1489 (N_1489,In_359,In_428);
and U1490 (N_1490,In_422,In_1468);
or U1491 (N_1491,In_743,In_256);
xnor U1492 (N_1492,In_1444,In_290);
nor U1493 (N_1493,In_288,In_106);
nand U1494 (N_1494,In_1183,In_1454);
nand U1495 (N_1495,In_604,In_1070);
nor U1496 (N_1496,In_274,In_1021);
or U1497 (N_1497,In_247,In_1362);
nand U1498 (N_1498,In_1089,In_172);
or U1499 (N_1499,In_1077,In_469);
nor U1500 (N_1500,In_74,In_2);
xnor U1501 (N_1501,In_27,In_327);
nor U1502 (N_1502,In_1310,In_1378);
xor U1503 (N_1503,In_13,In_929);
and U1504 (N_1504,In_184,In_921);
or U1505 (N_1505,In_349,In_210);
and U1506 (N_1506,In_105,In_980);
nor U1507 (N_1507,In_202,In_1099);
or U1508 (N_1508,In_1432,In_814);
nand U1509 (N_1509,In_439,In_863);
and U1510 (N_1510,In_558,In_1008);
and U1511 (N_1511,In_2,In_705);
and U1512 (N_1512,In_978,In_955);
or U1513 (N_1513,In_214,In_731);
and U1514 (N_1514,In_1201,In_1134);
or U1515 (N_1515,In_944,In_927);
xor U1516 (N_1516,In_146,In_445);
and U1517 (N_1517,In_648,In_199);
or U1518 (N_1518,In_1215,In_1235);
xor U1519 (N_1519,In_888,In_453);
and U1520 (N_1520,In_631,In_77);
nor U1521 (N_1521,In_100,In_546);
nor U1522 (N_1522,In_735,In_344);
nor U1523 (N_1523,In_917,In_52);
xnor U1524 (N_1524,In_1070,In_469);
nand U1525 (N_1525,In_116,In_211);
and U1526 (N_1526,In_962,In_1396);
nor U1527 (N_1527,In_137,In_716);
or U1528 (N_1528,In_1100,In_1481);
and U1529 (N_1529,In_803,In_789);
and U1530 (N_1530,In_108,In_492);
and U1531 (N_1531,In_2,In_902);
xnor U1532 (N_1532,In_1237,In_1455);
nor U1533 (N_1533,In_1139,In_1305);
or U1534 (N_1534,In_1094,In_206);
nor U1535 (N_1535,In_891,In_1349);
or U1536 (N_1536,In_457,In_474);
nand U1537 (N_1537,In_1105,In_1125);
and U1538 (N_1538,In_459,In_689);
nand U1539 (N_1539,In_705,In_753);
and U1540 (N_1540,In_1250,In_840);
nand U1541 (N_1541,In_1140,In_1232);
xor U1542 (N_1542,In_120,In_934);
nand U1543 (N_1543,In_1081,In_932);
and U1544 (N_1544,In_57,In_1296);
and U1545 (N_1545,In_534,In_1355);
nand U1546 (N_1546,In_1326,In_572);
or U1547 (N_1547,In_1028,In_488);
nor U1548 (N_1548,In_659,In_580);
xnor U1549 (N_1549,In_1105,In_192);
nor U1550 (N_1550,In_877,In_1493);
nand U1551 (N_1551,In_376,In_339);
nor U1552 (N_1552,In_610,In_1163);
nand U1553 (N_1553,In_689,In_1185);
or U1554 (N_1554,In_951,In_817);
nor U1555 (N_1555,In_1292,In_800);
or U1556 (N_1556,In_1441,In_980);
or U1557 (N_1557,In_252,In_190);
or U1558 (N_1558,In_760,In_351);
xnor U1559 (N_1559,In_1345,In_681);
nor U1560 (N_1560,In_117,In_504);
nor U1561 (N_1561,In_238,In_535);
and U1562 (N_1562,In_866,In_366);
or U1563 (N_1563,In_1341,In_1409);
xor U1564 (N_1564,In_1190,In_233);
or U1565 (N_1565,In_722,In_1112);
and U1566 (N_1566,In_723,In_775);
xnor U1567 (N_1567,In_1212,In_1110);
xnor U1568 (N_1568,In_941,In_75);
and U1569 (N_1569,In_451,In_1113);
and U1570 (N_1570,In_552,In_1277);
or U1571 (N_1571,In_26,In_1063);
nand U1572 (N_1572,In_75,In_1266);
nand U1573 (N_1573,In_413,In_295);
nand U1574 (N_1574,In_332,In_1379);
xnor U1575 (N_1575,In_298,In_582);
nand U1576 (N_1576,In_694,In_1372);
nand U1577 (N_1577,In_1063,In_596);
and U1578 (N_1578,In_1240,In_271);
and U1579 (N_1579,In_1219,In_213);
xor U1580 (N_1580,In_846,In_56);
xnor U1581 (N_1581,In_618,In_955);
and U1582 (N_1582,In_266,In_348);
nor U1583 (N_1583,In_58,In_1425);
and U1584 (N_1584,In_1324,In_145);
nor U1585 (N_1585,In_958,In_939);
or U1586 (N_1586,In_542,In_875);
nand U1587 (N_1587,In_954,In_319);
nand U1588 (N_1588,In_290,In_201);
nor U1589 (N_1589,In_1259,In_924);
nand U1590 (N_1590,In_586,In_1289);
and U1591 (N_1591,In_549,In_902);
nor U1592 (N_1592,In_164,In_224);
nand U1593 (N_1593,In_1466,In_809);
or U1594 (N_1594,In_241,In_274);
nor U1595 (N_1595,In_1499,In_912);
nor U1596 (N_1596,In_684,In_285);
nand U1597 (N_1597,In_650,In_1189);
or U1598 (N_1598,In_63,In_993);
nor U1599 (N_1599,In_625,In_1002);
nand U1600 (N_1600,In_614,In_942);
or U1601 (N_1601,In_776,In_546);
and U1602 (N_1602,In_1312,In_589);
nand U1603 (N_1603,In_817,In_309);
and U1604 (N_1604,In_1141,In_258);
nand U1605 (N_1605,In_889,In_386);
nand U1606 (N_1606,In_1159,In_971);
and U1607 (N_1607,In_425,In_801);
or U1608 (N_1608,In_1424,In_130);
and U1609 (N_1609,In_399,In_172);
nor U1610 (N_1610,In_9,In_942);
and U1611 (N_1611,In_785,In_3);
or U1612 (N_1612,In_1142,In_1133);
or U1613 (N_1613,In_370,In_1350);
xnor U1614 (N_1614,In_899,In_1209);
nor U1615 (N_1615,In_790,In_791);
nor U1616 (N_1616,In_1478,In_744);
nor U1617 (N_1617,In_197,In_365);
nand U1618 (N_1618,In_250,In_1226);
and U1619 (N_1619,In_653,In_889);
nor U1620 (N_1620,In_5,In_1484);
xor U1621 (N_1621,In_1147,In_200);
nor U1622 (N_1622,In_699,In_959);
and U1623 (N_1623,In_281,In_553);
nor U1624 (N_1624,In_973,In_431);
nand U1625 (N_1625,In_690,In_788);
or U1626 (N_1626,In_462,In_1393);
nor U1627 (N_1627,In_818,In_1286);
nor U1628 (N_1628,In_1027,In_1418);
xor U1629 (N_1629,In_922,In_532);
nand U1630 (N_1630,In_1197,In_333);
xor U1631 (N_1631,In_1134,In_321);
nand U1632 (N_1632,In_189,In_1308);
or U1633 (N_1633,In_1226,In_841);
or U1634 (N_1634,In_224,In_1383);
and U1635 (N_1635,In_1321,In_1140);
or U1636 (N_1636,In_1402,In_622);
and U1637 (N_1637,In_465,In_36);
xor U1638 (N_1638,In_1337,In_1189);
nand U1639 (N_1639,In_517,In_343);
nand U1640 (N_1640,In_391,In_692);
or U1641 (N_1641,In_252,In_1437);
or U1642 (N_1642,In_896,In_1096);
or U1643 (N_1643,In_1268,In_112);
nor U1644 (N_1644,In_1188,In_1403);
or U1645 (N_1645,In_356,In_100);
nor U1646 (N_1646,In_455,In_17);
and U1647 (N_1647,In_1020,In_138);
nor U1648 (N_1648,In_1084,In_699);
xnor U1649 (N_1649,In_870,In_109);
or U1650 (N_1650,In_186,In_53);
nor U1651 (N_1651,In_649,In_244);
nor U1652 (N_1652,In_239,In_1002);
nor U1653 (N_1653,In_1025,In_1408);
xor U1654 (N_1654,In_176,In_389);
xor U1655 (N_1655,In_1115,In_662);
nor U1656 (N_1656,In_412,In_1482);
or U1657 (N_1657,In_949,In_535);
and U1658 (N_1658,In_335,In_675);
nand U1659 (N_1659,In_903,In_703);
xor U1660 (N_1660,In_1432,In_279);
or U1661 (N_1661,In_304,In_815);
nor U1662 (N_1662,In_653,In_397);
nand U1663 (N_1663,In_532,In_1150);
nor U1664 (N_1664,In_184,In_1460);
or U1665 (N_1665,In_1468,In_1487);
or U1666 (N_1666,In_227,In_1102);
nor U1667 (N_1667,In_147,In_1064);
or U1668 (N_1668,In_107,In_164);
nor U1669 (N_1669,In_1358,In_820);
and U1670 (N_1670,In_1373,In_1102);
and U1671 (N_1671,In_1377,In_1287);
nor U1672 (N_1672,In_869,In_415);
nand U1673 (N_1673,In_1481,In_1394);
xnor U1674 (N_1674,In_164,In_616);
nand U1675 (N_1675,In_631,In_611);
xor U1676 (N_1676,In_1038,In_1225);
and U1677 (N_1677,In_129,In_890);
nand U1678 (N_1678,In_67,In_337);
and U1679 (N_1679,In_340,In_1371);
nand U1680 (N_1680,In_169,In_890);
and U1681 (N_1681,In_1409,In_1146);
or U1682 (N_1682,In_1207,In_648);
nor U1683 (N_1683,In_810,In_655);
and U1684 (N_1684,In_213,In_414);
xnor U1685 (N_1685,In_1435,In_606);
and U1686 (N_1686,In_736,In_25);
xnor U1687 (N_1687,In_1076,In_1227);
nor U1688 (N_1688,In_466,In_382);
and U1689 (N_1689,In_1359,In_1391);
or U1690 (N_1690,In_758,In_1365);
or U1691 (N_1691,In_629,In_465);
nand U1692 (N_1692,In_692,In_1006);
nor U1693 (N_1693,In_743,In_464);
nor U1694 (N_1694,In_669,In_838);
nand U1695 (N_1695,In_829,In_232);
nand U1696 (N_1696,In_1035,In_713);
xnor U1697 (N_1697,In_442,In_453);
and U1698 (N_1698,In_368,In_1436);
nand U1699 (N_1699,In_1452,In_399);
and U1700 (N_1700,In_1434,In_219);
nand U1701 (N_1701,In_114,In_222);
and U1702 (N_1702,In_148,In_298);
or U1703 (N_1703,In_282,In_990);
nor U1704 (N_1704,In_1165,In_561);
xor U1705 (N_1705,In_165,In_265);
or U1706 (N_1706,In_912,In_337);
nand U1707 (N_1707,In_249,In_1242);
nor U1708 (N_1708,In_917,In_145);
xnor U1709 (N_1709,In_1385,In_520);
nor U1710 (N_1710,In_511,In_1351);
nor U1711 (N_1711,In_489,In_1017);
and U1712 (N_1712,In_1279,In_573);
and U1713 (N_1713,In_583,In_1389);
nor U1714 (N_1714,In_456,In_1015);
xor U1715 (N_1715,In_1383,In_811);
or U1716 (N_1716,In_1411,In_1389);
xnor U1717 (N_1717,In_603,In_1365);
or U1718 (N_1718,In_256,In_462);
nor U1719 (N_1719,In_1126,In_1072);
and U1720 (N_1720,In_865,In_82);
nand U1721 (N_1721,In_1482,In_932);
or U1722 (N_1722,In_87,In_642);
nor U1723 (N_1723,In_1007,In_1468);
or U1724 (N_1724,In_880,In_1026);
nand U1725 (N_1725,In_544,In_345);
or U1726 (N_1726,In_507,In_94);
nand U1727 (N_1727,In_513,In_355);
or U1728 (N_1728,In_1358,In_810);
nor U1729 (N_1729,In_1314,In_544);
and U1730 (N_1730,In_1343,In_1166);
xor U1731 (N_1731,In_399,In_495);
or U1732 (N_1732,In_595,In_1393);
and U1733 (N_1733,In_488,In_125);
nor U1734 (N_1734,In_204,In_704);
xor U1735 (N_1735,In_708,In_442);
xor U1736 (N_1736,In_298,In_255);
and U1737 (N_1737,In_598,In_104);
or U1738 (N_1738,In_1466,In_1177);
or U1739 (N_1739,In_676,In_996);
or U1740 (N_1740,In_922,In_155);
and U1741 (N_1741,In_201,In_679);
or U1742 (N_1742,In_45,In_132);
nor U1743 (N_1743,In_1111,In_1278);
nor U1744 (N_1744,In_20,In_773);
and U1745 (N_1745,In_1401,In_318);
xnor U1746 (N_1746,In_663,In_453);
nand U1747 (N_1747,In_760,In_282);
nor U1748 (N_1748,In_480,In_708);
xnor U1749 (N_1749,In_460,In_1095);
nand U1750 (N_1750,In_230,In_518);
nand U1751 (N_1751,In_25,In_283);
nor U1752 (N_1752,In_1189,In_530);
nor U1753 (N_1753,In_855,In_1014);
and U1754 (N_1754,In_1397,In_720);
nor U1755 (N_1755,In_329,In_404);
nand U1756 (N_1756,In_1421,In_561);
and U1757 (N_1757,In_75,In_1255);
and U1758 (N_1758,In_288,In_1376);
nor U1759 (N_1759,In_12,In_485);
nor U1760 (N_1760,In_1235,In_358);
or U1761 (N_1761,In_358,In_93);
nor U1762 (N_1762,In_276,In_675);
or U1763 (N_1763,In_1356,In_1217);
or U1764 (N_1764,In_958,In_379);
nor U1765 (N_1765,In_167,In_469);
xor U1766 (N_1766,In_168,In_670);
and U1767 (N_1767,In_407,In_90);
nand U1768 (N_1768,In_59,In_72);
nor U1769 (N_1769,In_883,In_1061);
nand U1770 (N_1770,In_1323,In_1061);
xor U1771 (N_1771,In_162,In_748);
or U1772 (N_1772,In_80,In_268);
xnor U1773 (N_1773,In_209,In_415);
xor U1774 (N_1774,In_384,In_590);
nor U1775 (N_1775,In_361,In_1057);
nand U1776 (N_1776,In_1142,In_452);
nand U1777 (N_1777,In_146,In_900);
xor U1778 (N_1778,In_17,In_5);
nand U1779 (N_1779,In_507,In_79);
nand U1780 (N_1780,In_1350,In_231);
nand U1781 (N_1781,In_349,In_1129);
xor U1782 (N_1782,In_976,In_1201);
and U1783 (N_1783,In_72,In_534);
or U1784 (N_1784,In_710,In_870);
xnor U1785 (N_1785,In_1349,In_1430);
or U1786 (N_1786,In_669,In_758);
nand U1787 (N_1787,In_493,In_662);
or U1788 (N_1788,In_1076,In_566);
and U1789 (N_1789,In_1104,In_91);
and U1790 (N_1790,In_425,In_976);
xor U1791 (N_1791,In_919,In_897);
and U1792 (N_1792,In_298,In_1314);
nand U1793 (N_1793,In_721,In_269);
xnor U1794 (N_1794,In_636,In_684);
nor U1795 (N_1795,In_1298,In_1301);
or U1796 (N_1796,In_1223,In_599);
or U1797 (N_1797,In_352,In_744);
xor U1798 (N_1798,In_780,In_634);
nand U1799 (N_1799,In_1236,In_1363);
nor U1800 (N_1800,In_595,In_428);
or U1801 (N_1801,In_758,In_1474);
and U1802 (N_1802,In_918,In_604);
or U1803 (N_1803,In_284,In_527);
or U1804 (N_1804,In_210,In_1325);
or U1805 (N_1805,In_1357,In_1407);
or U1806 (N_1806,In_489,In_500);
nand U1807 (N_1807,In_1373,In_1406);
nor U1808 (N_1808,In_608,In_602);
or U1809 (N_1809,In_602,In_219);
and U1810 (N_1810,In_928,In_537);
nand U1811 (N_1811,In_1127,In_669);
nand U1812 (N_1812,In_443,In_1482);
or U1813 (N_1813,In_11,In_467);
and U1814 (N_1814,In_477,In_793);
or U1815 (N_1815,In_1332,In_442);
or U1816 (N_1816,In_247,In_1233);
nor U1817 (N_1817,In_541,In_486);
and U1818 (N_1818,In_900,In_996);
nand U1819 (N_1819,In_786,In_300);
xnor U1820 (N_1820,In_295,In_237);
or U1821 (N_1821,In_757,In_1222);
and U1822 (N_1822,In_328,In_1237);
nor U1823 (N_1823,In_1187,In_161);
or U1824 (N_1824,In_315,In_402);
nor U1825 (N_1825,In_1487,In_503);
nor U1826 (N_1826,In_667,In_94);
nor U1827 (N_1827,In_407,In_250);
xnor U1828 (N_1828,In_498,In_262);
nand U1829 (N_1829,In_116,In_907);
or U1830 (N_1830,In_1465,In_573);
or U1831 (N_1831,In_809,In_1293);
or U1832 (N_1832,In_215,In_370);
or U1833 (N_1833,In_728,In_1271);
or U1834 (N_1834,In_255,In_1220);
nand U1835 (N_1835,In_136,In_693);
and U1836 (N_1836,In_1245,In_948);
or U1837 (N_1837,In_1454,In_936);
or U1838 (N_1838,In_865,In_1063);
nor U1839 (N_1839,In_210,In_675);
or U1840 (N_1840,In_1061,In_583);
nor U1841 (N_1841,In_27,In_276);
or U1842 (N_1842,In_1238,In_1340);
xnor U1843 (N_1843,In_1476,In_1227);
and U1844 (N_1844,In_256,In_846);
xor U1845 (N_1845,In_653,In_1085);
nand U1846 (N_1846,In_1352,In_388);
nor U1847 (N_1847,In_1400,In_608);
or U1848 (N_1848,In_276,In_202);
nor U1849 (N_1849,In_1266,In_193);
nand U1850 (N_1850,In_576,In_1249);
nand U1851 (N_1851,In_1489,In_1320);
xnor U1852 (N_1852,In_969,In_173);
nand U1853 (N_1853,In_141,In_1055);
nand U1854 (N_1854,In_375,In_70);
nand U1855 (N_1855,In_861,In_641);
nand U1856 (N_1856,In_800,In_1300);
nor U1857 (N_1857,In_720,In_1412);
or U1858 (N_1858,In_1310,In_41);
and U1859 (N_1859,In_680,In_971);
nand U1860 (N_1860,In_661,In_584);
nand U1861 (N_1861,In_1482,In_309);
and U1862 (N_1862,In_1328,In_35);
nor U1863 (N_1863,In_499,In_349);
nand U1864 (N_1864,In_787,In_158);
and U1865 (N_1865,In_1160,In_319);
and U1866 (N_1866,In_1251,In_845);
nor U1867 (N_1867,In_1111,In_246);
and U1868 (N_1868,In_574,In_815);
xnor U1869 (N_1869,In_381,In_1029);
nand U1870 (N_1870,In_775,In_497);
and U1871 (N_1871,In_384,In_174);
or U1872 (N_1872,In_355,In_194);
nand U1873 (N_1873,In_427,In_1143);
nor U1874 (N_1874,In_1015,In_337);
nand U1875 (N_1875,In_1408,In_964);
nand U1876 (N_1876,In_470,In_1464);
xor U1877 (N_1877,In_400,In_176);
and U1878 (N_1878,In_1032,In_1400);
nor U1879 (N_1879,In_1067,In_476);
or U1880 (N_1880,In_646,In_16);
xor U1881 (N_1881,In_1279,In_104);
xnor U1882 (N_1882,In_918,In_310);
nand U1883 (N_1883,In_466,In_1211);
xor U1884 (N_1884,In_383,In_1054);
nand U1885 (N_1885,In_330,In_74);
xnor U1886 (N_1886,In_503,In_348);
and U1887 (N_1887,In_1037,In_503);
nand U1888 (N_1888,In_660,In_1199);
and U1889 (N_1889,In_457,In_695);
nor U1890 (N_1890,In_1411,In_729);
xor U1891 (N_1891,In_1311,In_1364);
nor U1892 (N_1892,In_1097,In_942);
nand U1893 (N_1893,In_1113,In_1401);
and U1894 (N_1894,In_456,In_1398);
nand U1895 (N_1895,In_1452,In_1045);
or U1896 (N_1896,In_25,In_449);
xnor U1897 (N_1897,In_166,In_146);
or U1898 (N_1898,In_1126,In_516);
and U1899 (N_1899,In_1147,In_547);
xnor U1900 (N_1900,In_643,In_404);
nor U1901 (N_1901,In_397,In_686);
and U1902 (N_1902,In_691,In_585);
nand U1903 (N_1903,In_5,In_874);
or U1904 (N_1904,In_1319,In_1003);
and U1905 (N_1905,In_781,In_95);
nor U1906 (N_1906,In_288,In_505);
nor U1907 (N_1907,In_575,In_520);
or U1908 (N_1908,In_1181,In_824);
xnor U1909 (N_1909,In_302,In_269);
or U1910 (N_1910,In_511,In_340);
xor U1911 (N_1911,In_296,In_775);
xnor U1912 (N_1912,In_1255,In_698);
nor U1913 (N_1913,In_911,In_929);
nor U1914 (N_1914,In_1203,In_758);
xor U1915 (N_1915,In_799,In_89);
and U1916 (N_1916,In_1113,In_323);
and U1917 (N_1917,In_1304,In_1233);
or U1918 (N_1918,In_641,In_1148);
or U1919 (N_1919,In_1477,In_1149);
nor U1920 (N_1920,In_1038,In_456);
xor U1921 (N_1921,In_561,In_1493);
nand U1922 (N_1922,In_58,In_615);
and U1923 (N_1923,In_519,In_1075);
and U1924 (N_1924,In_51,In_1372);
and U1925 (N_1925,In_911,In_204);
or U1926 (N_1926,In_1093,In_569);
xor U1927 (N_1927,In_145,In_497);
nor U1928 (N_1928,In_946,In_202);
nor U1929 (N_1929,In_589,In_295);
or U1930 (N_1930,In_1180,In_957);
and U1931 (N_1931,In_323,In_691);
and U1932 (N_1932,In_200,In_1294);
nand U1933 (N_1933,In_12,In_1499);
nor U1934 (N_1934,In_717,In_932);
nand U1935 (N_1935,In_471,In_900);
xnor U1936 (N_1936,In_542,In_1355);
nand U1937 (N_1937,In_688,In_59);
or U1938 (N_1938,In_1318,In_1198);
and U1939 (N_1939,In_404,In_38);
and U1940 (N_1940,In_535,In_798);
xor U1941 (N_1941,In_1076,In_1455);
xnor U1942 (N_1942,In_512,In_921);
or U1943 (N_1943,In_405,In_1350);
and U1944 (N_1944,In_1258,In_1422);
nand U1945 (N_1945,In_266,In_806);
or U1946 (N_1946,In_735,In_1185);
xnor U1947 (N_1947,In_1095,In_924);
nand U1948 (N_1948,In_148,In_760);
and U1949 (N_1949,In_357,In_816);
nand U1950 (N_1950,In_806,In_10);
nand U1951 (N_1951,In_307,In_297);
nand U1952 (N_1952,In_949,In_1364);
nor U1953 (N_1953,In_1090,In_51);
and U1954 (N_1954,In_388,In_937);
nand U1955 (N_1955,In_115,In_371);
xor U1956 (N_1956,In_1210,In_790);
and U1957 (N_1957,In_1236,In_417);
nor U1958 (N_1958,In_1172,In_413);
nand U1959 (N_1959,In_764,In_297);
and U1960 (N_1960,In_402,In_472);
nand U1961 (N_1961,In_1090,In_264);
nand U1962 (N_1962,In_1411,In_1105);
xnor U1963 (N_1963,In_160,In_990);
or U1964 (N_1964,In_1141,In_1203);
and U1965 (N_1965,In_257,In_400);
xnor U1966 (N_1966,In_488,In_495);
nand U1967 (N_1967,In_780,In_1426);
or U1968 (N_1968,In_881,In_1134);
and U1969 (N_1969,In_1248,In_897);
nor U1970 (N_1970,In_1376,In_675);
or U1971 (N_1971,In_1100,In_1394);
nand U1972 (N_1972,In_363,In_1025);
nor U1973 (N_1973,In_1182,In_118);
nor U1974 (N_1974,In_761,In_715);
and U1975 (N_1975,In_1300,In_132);
or U1976 (N_1976,In_1075,In_494);
nor U1977 (N_1977,In_1239,In_1324);
nor U1978 (N_1978,In_178,In_272);
nand U1979 (N_1979,In_199,In_1074);
and U1980 (N_1980,In_950,In_1355);
nor U1981 (N_1981,In_1084,In_754);
and U1982 (N_1982,In_365,In_1306);
nor U1983 (N_1983,In_1401,In_64);
or U1984 (N_1984,In_482,In_1225);
or U1985 (N_1985,In_699,In_1149);
or U1986 (N_1986,In_723,In_482);
and U1987 (N_1987,In_254,In_446);
nor U1988 (N_1988,In_626,In_835);
nand U1989 (N_1989,In_1249,In_274);
or U1990 (N_1990,In_672,In_1159);
and U1991 (N_1991,In_1077,In_414);
nand U1992 (N_1992,In_1135,In_56);
nand U1993 (N_1993,In_562,In_1284);
and U1994 (N_1994,In_1440,In_722);
and U1995 (N_1995,In_945,In_594);
and U1996 (N_1996,In_1418,In_330);
nor U1997 (N_1997,In_315,In_1449);
nand U1998 (N_1998,In_1065,In_1106);
and U1999 (N_1999,In_1295,In_32);
nor U2000 (N_2000,In_1018,In_847);
xnor U2001 (N_2001,In_804,In_280);
and U2002 (N_2002,In_243,In_1225);
nor U2003 (N_2003,In_1460,In_984);
xor U2004 (N_2004,In_701,In_886);
xnor U2005 (N_2005,In_344,In_533);
nor U2006 (N_2006,In_894,In_1065);
nand U2007 (N_2007,In_395,In_365);
nand U2008 (N_2008,In_964,In_531);
or U2009 (N_2009,In_602,In_1080);
nand U2010 (N_2010,In_719,In_904);
nand U2011 (N_2011,In_1145,In_1031);
nand U2012 (N_2012,In_112,In_1303);
nand U2013 (N_2013,In_955,In_718);
nor U2014 (N_2014,In_1492,In_453);
xor U2015 (N_2015,In_857,In_652);
or U2016 (N_2016,In_181,In_157);
xnor U2017 (N_2017,In_322,In_254);
nand U2018 (N_2018,In_159,In_963);
and U2019 (N_2019,In_694,In_896);
and U2020 (N_2020,In_763,In_161);
nor U2021 (N_2021,In_342,In_679);
nor U2022 (N_2022,In_1363,In_903);
nor U2023 (N_2023,In_90,In_1161);
xnor U2024 (N_2024,In_319,In_758);
xor U2025 (N_2025,In_1422,In_729);
or U2026 (N_2026,In_1481,In_635);
or U2027 (N_2027,In_587,In_1425);
and U2028 (N_2028,In_845,In_150);
or U2029 (N_2029,In_1260,In_1098);
nor U2030 (N_2030,In_1381,In_147);
or U2031 (N_2031,In_907,In_620);
xnor U2032 (N_2032,In_1498,In_1412);
xor U2033 (N_2033,In_1398,In_1082);
or U2034 (N_2034,In_80,In_988);
or U2035 (N_2035,In_1210,In_646);
or U2036 (N_2036,In_1322,In_6);
nor U2037 (N_2037,In_573,In_59);
and U2038 (N_2038,In_987,In_392);
or U2039 (N_2039,In_97,In_475);
and U2040 (N_2040,In_357,In_933);
nand U2041 (N_2041,In_1298,In_1044);
nand U2042 (N_2042,In_870,In_1405);
nand U2043 (N_2043,In_727,In_123);
or U2044 (N_2044,In_911,In_117);
xor U2045 (N_2045,In_1382,In_347);
xnor U2046 (N_2046,In_1193,In_1086);
nor U2047 (N_2047,In_1117,In_589);
xnor U2048 (N_2048,In_1030,In_1322);
and U2049 (N_2049,In_891,In_418);
or U2050 (N_2050,In_182,In_1252);
xnor U2051 (N_2051,In_71,In_652);
xnor U2052 (N_2052,In_1385,In_245);
xnor U2053 (N_2053,In_420,In_253);
nand U2054 (N_2054,In_1389,In_220);
and U2055 (N_2055,In_679,In_1120);
xnor U2056 (N_2056,In_1065,In_589);
xnor U2057 (N_2057,In_47,In_225);
xor U2058 (N_2058,In_99,In_674);
nor U2059 (N_2059,In_64,In_332);
nand U2060 (N_2060,In_943,In_444);
nand U2061 (N_2061,In_331,In_511);
and U2062 (N_2062,In_502,In_1150);
and U2063 (N_2063,In_288,In_3);
nor U2064 (N_2064,In_610,In_419);
or U2065 (N_2065,In_146,In_829);
and U2066 (N_2066,In_269,In_147);
xor U2067 (N_2067,In_1373,In_965);
and U2068 (N_2068,In_530,In_522);
and U2069 (N_2069,In_34,In_240);
nand U2070 (N_2070,In_941,In_951);
nor U2071 (N_2071,In_689,In_609);
xnor U2072 (N_2072,In_934,In_393);
or U2073 (N_2073,In_1489,In_773);
and U2074 (N_2074,In_579,In_1184);
or U2075 (N_2075,In_714,In_1438);
nor U2076 (N_2076,In_1020,In_1302);
nand U2077 (N_2077,In_366,In_602);
nand U2078 (N_2078,In_28,In_1414);
and U2079 (N_2079,In_100,In_105);
or U2080 (N_2080,In_669,In_303);
nand U2081 (N_2081,In_132,In_148);
and U2082 (N_2082,In_217,In_1114);
and U2083 (N_2083,In_606,In_896);
and U2084 (N_2084,In_1187,In_127);
xor U2085 (N_2085,In_951,In_1219);
xor U2086 (N_2086,In_282,In_616);
and U2087 (N_2087,In_1427,In_412);
and U2088 (N_2088,In_627,In_1094);
or U2089 (N_2089,In_620,In_550);
nand U2090 (N_2090,In_1352,In_1199);
nor U2091 (N_2091,In_79,In_96);
and U2092 (N_2092,In_292,In_299);
nor U2093 (N_2093,In_833,In_948);
or U2094 (N_2094,In_1053,In_992);
nand U2095 (N_2095,In_759,In_329);
and U2096 (N_2096,In_495,In_1408);
xnor U2097 (N_2097,In_533,In_835);
nor U2098 (N_2098,In_1438,In_1160);
nor U2099 (N_2099,In_340,In_1158);
or U2100 (N_2100,In_1132,In_1229);
xor U2101 (N_2101,In_167,In_417);
nor U2102 (N_2102,In_1307,In_1373);
or U2103 (N_2103,In_474,In_962);
or U2104 (N_2104,In_772,In_1450);
nand U2105 (N_2105,In_168,In_506);
nor U2106 (N_2106,In_558,In_432);
and U2107 (N_2107,In_1151,In_998);
and U2108 (N_2108,In_891,In_175);
xor U2109 (N_2109,In_456,In_167);
nor U2110 (N_2110,In_290,In_1477);
or U2111 (N_2111,In_876,In_615);
xnor U2112 (N_2112,In_526,In_260);
nor U2113 (N_2113,In_1026,In_150);
nor U2114 (N_2114,In_176,In_883);
xor U2115 (N_2115,In_1082,In_294);
xnor U2116 (N_2116,In_1385,In_569);
and U2117 (N_2117,In_168,In_913);
and U2118 (N_2118,In_736,In_986);
or U2119 (N_2119,In_824,In_1389);
or U2120 (N_2120,In_802,In_85);
nand U2121 (N_2121,In_555,In_524);
or U2122 (N_2122,In_164,In_1269);
nand U2123 (N_2123,In_643,In_690);
nor U2124 (N_2124,In_466,In_21);
nor U2125 (N_2125,In_661,In_454);
or U2126 (N_2126,In_275,In_1015);
and U2127 (N_2127,In_1101,In_764);
or U2128 (N_2128,In_263,In_605);
nor U2129 (N_2129,In_236,In_39);
or U2130 (N_2130,In_904,In_115);
and U2131 (N_2131,In_864,In_156);
nor U2132 (N_2132,In_558,In_1489);
or U2133 (N_2133,In_323,In_783);
or U2134 (N_2134,In_1301,In_607);
nor U2135 (N_2135,In_1239,In_979);
nand U2136 (N_2136,In_1161,In_707);
xnor U2137 (N_2137,In_399,In_1351);
nand U2138 (N_2138,In_1390,In_1097);
xor U2139 (N_2139,In_775,In_934);
or U2140 (N_2140,In_1375,In_591);
nand U2141 (N_2141,In_79,In_805);
or U2142 (N_2142,In_424,In_1009);
xor U2143 (N_2143,In_807,In_1332);
nand U2144 (N_2144,In_617,In_1177);
nor U2145 (N_2145,In_71,In_926);
or U2146 (N_2146,In_184,In_1122);
nand U2147 (N_2147,In_912,In_1472);
nand U2148 (N_2148,In_363,In_709);
nor U2149 (N_2149,In_133,In_943);
nand U2150 (N_2150,In_354,In_958);
and U2151 (N_2151,In_1499,In_209);
nand U2152 (N_2152,In_127,In_392);
xor U2153 (N_2153,In_714,In_364);
xnor U2154 (N_2154,In_1475,In_918);
or U2155 (N_2155,In_910,In_628);
and U2156 (N_2156,In_472,In_905);
xnor U2157 (N_2157,In_221,In_1376);
nand U2158 (N_2158,In_1027,In_148);
nor U2159 (N_2159,In_1189,In_1181);
or U2160 (N_2160,In_60,In_391);
and U2161 (N_2161,In_1136,In_1376);
xnor U2162 (N_2162,In_709,In_728);
nand U2163 (N_2163,In_346,In_268);
and U2164 (N_2164,In_841,In_1293);
xor U2165 (N_2165,In_803,In_684);
xor U2166 (N_2166,In_1098,In_1);
or U2167 (N_2167,In_976,In_1431);
nand U2168 (N_2168,In_14,In_536);
and U2169 (N_2169,In_632,In_691);
and U2170 (N_2170,In_1015,In_335);
and U2171 (N_2171,In_115,In_1471);
and U2172 (N_2172,In_1245,In_313);
nand U2173 (N_2173,In_1189,In_1400);
nand U2174 (N_2174,In_1242,In_773);
nor U2175 (N_2175,In_623,In_605);
nand U2176 (N_2176,In_1263,In_1049);
and U2177 (N_2177,In_1467,In_258);
or U2178 (N_2178,In_1344,In_500);
nor U2179 (N_2179,In_601,In_734);
nor U2180 (N_2180,In_1029,In_391);
nor U2181 (N_2181,In_549,In_1164);
and U2182 (N_2182,In_852,In_948);
nand U2183 (N_2183,In_775,In_491);
nand U2184 (N_2184,In_683,In_646);
xnor U2185 (N_2185,In_660,In_438);
xor U2186 (N_2186,In_1085,In_937);
and U2187 (N_2187,In_426,In_343);
nand U2188 (N_2188,In_1411,In_159);
and U2189 (N_2189,In_794,In_775);
and U2190 (N_2190,In_342,In_556);
nand U2191 (N_2191,In_120,In_573);
nor U2192 (N_2192,In_1211,In_316);
nand U2193 (N_2193,In_934,In_1023);
nand U2194 (N_2194,In_1005,In_518);
or U2195 (N_2195,In_537,In_328);
and U2196 (N_2196,In_275,In_1267);
and U2197 (N_2197,In_1192,In_456);
xnor U2198 (N_2198,In_1072,In_1129);
and U2199 (N_2199,In_1146,In_1441);
xnor U2200 (N_2200,In_657,In_663);
and U2201 (N_2201,In_1028,In_519);
nand U2202 (N_2202,In_859,In_1399);
xor U2203 (N_2203,In_1031,In_1194);
nand U2204 (N_2204,In_937,In_1360);
nor U2205 (N_2205,In_1304,In_1279);
or U2206 (N_2206,In_1073,In_731);
xor U2207 (N_2207,In_587,In_445);
nor U2208 (N_2208,In_773,In_431);
nand U2209 (N_2209,In_214,In_596);
and U2210 (N_2210,In_1221,In_705);
nand U2211 (N_2211,In_316,In_90);
and U2212 (N_2212,In_67,In_1367);
and U2213 (N_2213,In_558,In_805);
xnor U2214 (N_2214,In_386,In_404);
or U2215 (N_2215,In_54,In_1098);
nor U2216 (N_2216,In_928,In_921);
and U2217 (N_2217,In_476,In_843);
nand U2218 (N_2218,In_1329,In_121);
xor U2219 (N_2219,In_1133,In_595);
nand U2220 (N_2220,In_1485,In_320);
nand U2221 (N_2221,In_473,In_1036);
and U2222 (N_2222,In_729,In_361);
nand U2223 (N_2223,In_707,In_469);
nor U2224 (N_2224,In_521,In_1330);
and U2225 (N_2225,In_606,In_736);
and U2226 (N_2226,In_601,In_579);
xnor U2227 (N_2227,In_431,In_1109);
nor U2228 (N_2228,In_1471,In_303);
nand U2229 (N_2229,In_1207,In_455);
nand U2230 (N_2230,In_253,In_995);
and U2231 (N_2231,In_26,In_475);
nand U2232 (N_2232,In_897,In_926);
nand U2233 (N_2233,In_1095,In_630);
and U2234 (N_2234,In_38,In_1285);
or U2235 (N_2235,In_484,In_435);
nor U2236 (N_2236,In_1208,In_526);
nor U2237 (N_2237,In_38,In_836);
nand U2238 (N_2238,In_1105,In_1235);
nand U2239 (N_2239,In_267,In_505);
nand U2240 (N_2240,In_1258,In_1037);
nand U2241 (N_2241,In_257,In_252);
nand U2242 (N_2242,In_96,In_1270);
or U2243 (N_2243,In_118,In_563);
xnor U2244 (N_2244,In_1341,In_942);
or U2245 (N_2245,In_419,In_720);
and U2246 (N_2246,In_1024,In_1023);
xor U2247 (N_2247,In_400,In_989);
nand U2248 (N_2248,In_630,In_964);
nand U2249 (N_2249,In_823,In_1418);
and U2250 (N_2250,In_1106,In_1236);
xor U2251 (N_2251,In_920,In_1128);
or U2252 (N_2252,In_1320,In_942);
or U2253 (N_2253,In_704,In_838);
xor U2254 (N_2254,In_956,In_892);
xor U2255 (N_2255,In_206,In_549);
xor U2256 (N_2256,In_1004,In_507);
and U2257 (N_2257,In_673,In_933);
xnor U2258 (N_2258,In_454,In_1203);
nand U2259 (N_2259,In_201,In_1003);
and U2260 (N_2260,In_1022,In_1374);
and U2261 (N_2261,In_485,In_241);
and U2262 (N_2262,In_487,In_259);
xor U2263 (N_2263,In_464,In_577);
nand U2264 (N_2264,In_1180,In_1058);
and U2265 (N_2265,In_1141,In_578);
nor U2266 (N_2266,In_503,In_703);
nand U2267 (N_2267,In_10,In_38);
nand U2268 (N_2268,In_183,In_1296);
nor U2269 (N_2269,In_200,In_872);
and U2270 (N_2270,In_1044,In_1153);
nand U2271 (N_2271,In_866,In_1069);
and U2272 (N_2272,In_1449,In_286);
nor U2273 (N_2273,In_1071,In_1246);
nor U2274 (N_2274,In_781,In_394);
nor U2275 (N_2275,In_348,In_161);
or U2276 (N_2276,In_144,In_1195);
and U2277 (N_2277,In_21,In_1475);
or U2278 (N_2278,In_367,In_447);
nand U2279 (N_2279,In_36,In_780);
or U2280 (N_2280,In_1212,In_332);
nor U2281 (N_2281,In_156,In_163);
nor U2282 (N_2282,In_407,In_240);
nor U2283 (N_2283,In_148,In_622);
or U2284 (N_2284,In_495,In_677);
and U2285 (N_2285,In_1142,In_563);
xor U2286 (N_2286,In_1108,In_259);
nand U2287 (N_2287,In_355,In_1264);
nor U2288 (N_2288,In_1017,In_545);
nand U2289 (N_2289,In_1382,In_1031);
or U2290 (N_2290,In_271,In_32);
or U2291 (N_2291,In_542,In_384);
xor U2292 (N_2292,In_367,In_847);
xnor U2293 (N_2293,In_1343,In_89);
xor U2294 (N_2294,In_36,In_772);
and U2295 (N_2295,In_8,In_326);
and U2296 (N_2296,In_1338,In_743);
nor U2297 (N_2297,In_466,In_728);
nand U2298 (N_2298,In_669,In_1441);
nand U2299 (N_2299,In_163,In_1120);
nand U2300 (N_2300,In_1301,In_311);
and U2301 (N_2301,In_357,In_1347);
nand U2302 (N_2302,In_1034,In_449);
or U2303 (N_2303,In_352,In_765);
xor U2304 (N_2304,In_34,In_1283);
nand U2305 (N_2305,In_695,In_134);
nor U2306 (N_2306,In_127,In_796);
nor U2307 (N_2307,In_1407,In_140);
and U2308 (N_2308,In_708,In_1003);
nand U2309 (N_2309,In_495,In_628);
nor U2310 (N_2310,In_1281,In_458);
nor U2311 (N_2311,In_131,In_156);
xnor U2312 (N_2312,In_1128,In_1292);
or U2313 (N_2313,In_1171,In_456);
xnor U2314 (N_2314,In_309,In_930);
nor U2315 (N_2315,In_379,In_1283);
and U2316 (N_2316,In_1470,In_30);
or U2317 (N_2317,In_740,In_570);
or U2318 (N_2318,In_1169,In_104);
nand U2319 (N_2319,In_1258,In_1036);
xor U2320 (N_2320,In_790,In_910);
and U2321 (N_2321,In_718,In_647);
xnor U2322 (N_2322,In_759,In_100);
nor U2323 (N_2323,In_1367,In_936);
xor U2324 (N_2324,In_1146,In_119);
nand U2325 (N_2325,In_957,In_502);
nand U2326 (N_2326,In_825,In_1080);
nor U2327 (N_2327,In_886,In_245);
or U2328 (N_2328,In_491,In_1123);
xor U2329 (N_2329,In_1216,In_1366);
or U2330 (N_2330,In_1156,In_1076);
nand U2331 (N_2331,In_178,In_705);
xor U2332 (N_2332,In_299,In_925);
nor U2333 (N_2333,In_337,In_340);
nor U2334 (N_2334,In_1403,In_790);
and U2335 (N_2335,In_1220,In_1225);
xor U2336 (N_2336,In_757,In_1429);
or U2337 (N_2337,In_147,In_124);
xnor U2338 (N_2338,In_1417,In_762);
and U2339 (N_2339,In_782,In_1328);
nor U2340 (N_2340,In_858,In_831);
xor U2341 (N_2341,In_888,In_552);
and U2342 (N_2342,In_588,In_448);
or U2343 (N_2343,In_349,In_67);
xnor U2344 (N_2344,In_1053,In_1176);
and U2345 (N_2345,In_284,In_335);
xor U2346 (N_2346,In_1241,In_709);
nor U2347 (N_2347,In_418,In_430);
or U2348 (N_2348,In_688,In_120);
and U2349 (N_2349,In_725,In_1266);
xnor U2350 (N_2350,In_24,In_1080);
nand U2351 (N_2351,In_882,In_868);
or U2352 (N_2352,In_526,In_1171);
and U2353 (N_2353,In_578,In_430);
or U2354 (N_2354,In_1116,In_441);
nor U2355 (N_2355,In_88,In_8);
nand U2356 (N_2356,In_471,In_664);
nor U2357 (N_2357,In_1450,In_1006);
and U2358 (N_2358,In_878,In_522);
xnor U2359 (N_2359,In_326,In_512);
and U2360 (N_2360,In_832,In_45);
nand U2361 (N_2361,In_1333,In_1054);
nand U2362 (N_2362,In_1275,In_22);
or U2363 (N_2363,In_843,In_724);
and U2364 (N_2364,In_279,In_1023);
xnor U2365 (N_2365,In_1238,In_692);
nor U2366 (N_2366,In_1358,In_1120);
nor U2367 (N_2367,In_161,In_462);
and U2368 (N_2368,In_1382,In_1105);
nor U2369 (N_2369,In_1217,In_511);
nand U2370 (N_2370,In_73,In_1252);
nor U2371 (N_2371,In_596,In_158);
nand U2372 (N_2372,In_656,In_605);
nor U2373 (N_2373,In_566,In_1114);
or U2374 (N_2374,In_251,In_1339);
nand U2375 (N_2375,In_749,In_641);
nand U2376 (N_2376,In_1184,In_1102);
or U2377 (N_2377,In_158,In_940);
xor U2378 (N_2378,In_385,In_247);
and U2379 (N_2379,In_90,In_1337);
xor U2380 (N_2380,In_974,In_1472);
nand U2381 (N_2381,In_1477,In_279);
or U2382 (N_2382,In_1148,In_1);
or U2383 (N_2383,In_1491,In_1402);
nand U2384 (N_2384,In_180,In_764);
or U2385 (N_2385,In_1144,In_7);
xor U2386 (N_2386,In_759,In_1440);
nor U2387 (N_2387,In_832,In_690);
nor U2388 (N_2388,In_1306,In_1173);
xnor U2389 (N_2389,In_997,In_182);
or U2390 (N_2390,In_686,In_633);
nand U2391 (N_2391,In_616,In_1276);
nor U2392 (N_2392,In_2,In_279);
nor U2393 (N_2393,In_171,In_1096);
or U2394 (N_2394,In_388,In_357);
xnor U2395 (N_2395,In_456,In_1415);
nand U2396 (N_2396,In_1234,In_1323);
and U2397 (N_2397,In_498,In_842);
nand U2398 (N_2398,In_782,In_586);
nor U2399 (N_2399,In_738,In_298);
or U2400 (N_2400,In_1490,In_523);
and U2401 (N_2401,In_1262,In_518);
nor U2402 (N_2402,In_1160,In_208);
xor U2403 (N_2403,In_1402,In_1385);
xor U2404 (N_2404,In_626,In_64);
xor U2405 (N_2405,In_999,In_159);
and U2406 (N_2406,In_1443,In_1269);
and U2407 (N_2407,In_1317,In_1258);
nand U2408 (N_2408,In_1381,In_1488);
or U2409 (N_2409,In_1249,In_1482);
nor U2410 (N_2410,In_650,In_1023);
xor U2411 (N_2411,In_1374,In_888);
and U2412 (N_2412,In_781,In_499);
or U2413 (N_2413,In_1405,In_4);
or U2414 (N_2414,In_225,In_956);
nor U2415 (N_2415,In_422,In_948);
nand U2416 (N_2416,In_1406,In_1469);
nor U2417 (N_2417,In_1000,In_1284);
nor U2418 (N_2418,In_1490,In_1448);
nand U2419 (N_2419,In_206,In_1250);
nor U2420 (N_2420,In_92,In_51);
or U2421 (N_2421,In_1350,In_1399);
nor U2422 (N_2422,In_107,In_761);
or U2423 (N_2423,In_800,In_330);
or U2424 (N_2424,In_1191,In_985);
nor U2425 (N_2425,In_787,In_689);
and U2426 (N_2426,In_1457,In_371);
or U2427 (N_2427,In_1326,In_139);
xor U2428 (N_2428,In_494,In_484);
or U2429 (N_2429,In_810,In_1198);
xnor U2430 (N_2430,In_123,In_1203);
and U2431 (N_2431,In_51,In_305);
nand U2432 (N_2432,In_428,In_451);
or U2433 (N_2433,In_940,In_515);
or U2434 (N_2434,In_880,In_788);
and U2435 (N_2435,In_543,In_123);
nor U2436 (N_2436,In_1078,In_786);
nand U2437 (N_2437,In_986,In_530);
nand U2438 (N_2438,In_1187,In_737);
or U2439 (N_2439,In_246,In_327);
nor U2440 (N_2440,In_370,In_47);
nand U2441 (N_2441,In_280,In_920);
and U2442 (N_2442,In_533,In_807);
or U2443 (N_2443,In_340,In_688);
or U2444 (N_2444,In_423,In_492);
nand U2445 (N_2445,In_106,In_603);
nor U2446 (N_2446,In_5,In_8);
and U2447 (N_2447,In_140,In_345);
xor U2448 (N_2448,In_205,In_1003);
nor U2449 (N_2449,In_1249,In_804);
and U2450 (N_2450,In_1095,In_726);
xnor U2451 (N_2451,In_773,In_658);
or U2452 (N_2452,In_135,In_1407);
nand U2453 (N_2453,In_1494,In_1020);
xnor U2454 (N_2454,In_981,In_1178);
nor U2455 (N_2455,In_338,In_1275);
or U2456 (N_2456,In_992,In_710);
or U2457 (N_2457,In_1059,In_210);
nand U2458 (N_2458,In_1435,In_342);
xor U2459 (N_2459,In_1325,In_1139);
nor U2460 (N_2460,In_323,In_432);
and U2461 (N_2461,In_253,In_131);
or U2462 (N_2462,In_931,In_779);
and U2463 (N_2463,In_898,In_869);
nand U2464 (N_2464,In_381,In_277);
xor U2465 (N_2465,In_392,In_469);
nand U2466 (N_2466,In_104,In_642);
xor U2467 (N_2467,In_1022,In_1345);
nor U2468 (N_2468,In_413,In_1202);
nor U2469 (N_2469,In_1066,In_73);
or U2470 (N_2470,In_1162,In_669);
nand U2471 (N_2471,In_557,In_1063);
or U2472 (N_2472,In_560,In_976);
or U2473 (N_2473,In_80,In_953);
and U2474 (N_2474,In_322,In_780);
nor U2475 (N_2475,In_1334,In_565);
nand U2476 (N_2476,In_293,In_1267);
nand U2477 (N_2477,In_169,In_797);
and U2478 (N_2478,In_531,In_873);
nor U2479 (N_2479,In_265,In_1091);
nand U2480 (N_2480,In_690,In_436);
or U2481 (N_2481,In_1039,In_1352);
nor U2482 (N_2482,In_1129,In_437);
nand U2483 (N_2483,In_417,In_577);
xor U2484 (N_2484,In_1063,In_706);
xnor U2485 (N_2485,In_329,In_1478);
and U2486 (N_2486,In_346,In_217);
nor U2487 (N_2487,In_998,In_1189);
nand U2488 (N_2488,In_530,In_1163);
nand U2489 (N_2489,In_700,In_1109);
xor U2490 (N_2490,In_1282,In_351);
or U2491 (N_2491,In_635,In_1035);
nor U2492 (N_2492,In_1286,In_117);
or U2493 (N_2493,In_1301,In_1058);
and U2494 (N_2494,In_371,In_1114);
xnor U2495 (N_2495,In_359,In_1076);
nor U2496 (N_2496,In_634,In_662);
and U2497 (N_2497,In_268,In_1069);
or U2498 (N_2498,In_1080,In_691);
or U2499 (N_2499,In_865,In_741);
xor U2500 (N_2500,In_163,In_1013);
nand U2501 (N_2501,In_1490,In_151);
xnor U2502 (N_2502,In_1230,In_1427);
xnor U2503 (N_2503,In_995,In_529);
nor U2504 (N_2504,In_1464,In_1336);
nor U2505 (N_2505,In_399,In_681);
and U2506 (N_2506,In_1008,In_896);
and U2507 (N_2507,In_880,In_1454);
and U2508 (N_2508,In_1323,In_348);
nand U2509 (N_2509,In_608,In_344);
and U2510 (N_2510,In_521,In_1113);
and U2511 (N_2511,In_460,In_1061);
nor U2512 (N_2512,In_942,In_1400);
nand U2513 (N_2513,In_355,In_389);
and U2514 (N_2514,In_1220,In_1262);
and U2515 (N_2515,In_982,In_335);
nor U2516 (N_2516,In_908,In_1195);
nand U2517 (N_2517,In_74,In_1440);
nor U2518 (N_2518,In_461,In_614);
xor U2519 (N_2519,In_148,In_801);
and U2520 (N_2520,In_1343,In_1);
xnor U2521 (N_2521,In_1304,In_1447);
and U2522 (N_2522,In_293,In_142);
and U2523 (N_2523,In_1020,In_1203);
and U2524 (N_2524,In_109,In_1181);
and U2525 (N_2525,In_1298,In_42);
xnor U2526 (N_2526,In_99,In_1032);
xor U2527 (N_2527,In_654,In_313);
and U2528 (N_2528,In_615,In_1116);
and U2529 (N_2529,In_372,In_861);
and U2530 (N_2530,In_1189,In_492);
xor U2531 (N_2531,In_1094,In_750);
nand U2532 (N_2532,In_600,In_89);
xnor U2533 (N_2533,In_1485,In_1117);
or U2534 (N_2534,In_812,In_482);
nor U2535 (N_2535,In_824,In_1362);
and U2536 (N_2536,In_463,In_1155);
nor U2537 (N_2537,In_1261,In_1285);
nand U2538 (N_2538,In_250,In_1147);
nand U2539 (N_2539,In_1076,In_834);
nand U2540 (N_2540,In_751,In_1029);
and U2541 (N_2541,In_1457,In_1229);
nor U2542 (N_2542,In_355,In_946);
nor U2543 (N_2543,In_1060,In_208);
or U2544 (N_2544,In_1293,In_427);
and U2545 (N_2545,In_14,In_1170);
nand U2546 (N_2546,In_1271,In_1492);
nor U2547 (N_2547,In_688,In_1122);
xor U2548 (N_2548,In_1326,In_1484);
or U2549 (N_2549,In_775,In_405);
xnor U2550 (N_2550,In_38,In_750);
or U2551 (N_2551,In_1093,In_424);
and U2552 (N_2552,In_449,In_1430);
and U2553 (N_2553,In_423,In_1267);
xnor U2554 (N_2554,In_605,In_472);
xnor U2555 (N_2555,In_607,In_791);
nand U2556 (N_2556,In_1415,In_1052);
nand U2557 (N_2557,In_395,In_565);
or U2558 (N_2558,In_95,In_777);
nor U2559 (N_2559,In_548,In_476);
nand U2560 (N_2560,In_910,In_807);
or U2561 (N_2561,In_997,In_291);
and U2562 (N_2562,In_679,In_1360);
and U2563 (N_2563,In_27,In_1042);
and U2564 (N_2564,In_711,In_959);
nand U2565 (N_2565,In_1299,In_860);
nand U2566 (N_2566,In_444,In_335);
or U2567 (N_2567,In_22,In_6);
nor U2568 (N_2568,In_1201,In_1173);
nor U2569 (N_2569,In_1090,In_1337);
xor U2570 (N_2570,In_213,In_1053);
and U2571 (N_2571,In_1059,In_203);
nor U2572 (N_2572,In_505,In_911);
xnor U2573 (N_2573,In_1092,In_104);
and U2574 (N_2574,In_723,In_967);
and U2575 (N_2575,In_905,In_188);
xnor U2576 (N_2576,In_1479,In_205);
and U2577 (N_2577,In_714,In_1314);
xor U2578 (N_2578,In_409,In_273);
and U2579 (N_2579,In_1437,In_166);
nand U2580 (N_2580,In_684,In_9);
nor U2581 (N_2581,In_1106,In_359);
xor U2582 (N_2582,In_1062,In_1057);
or U2583 (N_2583,In_899,In_753);
nor U2584 (N_2584,In_1281,In_513);
xnor U2585 (N_2585,In_89,In_737);
and U2586 (N_2586,In_1185,In_31);
nand U2587 (N_2587,In_43,In_1143);
nor U2588 (N_2588,In_1246,In_1010);
and U2589 (N_2589,In_577,In_225);
and U2590 (N_2590,In_757,In_1421);
xor U2591 (N_2591,In_820,In_1317);
xor U2592 (N_2592,In_1102,In_929);
xnor U2593 (N_2593,In_1211,In_564);
and U2594 (N_2594,In_1336,In_1194);
xnor U2595 (N_2595,In_1267,In_302);
xnor U2596 (N_2596,In_353,In_1015);
xnor U2597 (N_2597,In_723,In_1147);
nor U2598 (N_2598,In_666,In_906);
xnor U2599 (N_2599,In_455,In_301);
nand U2600 (N_2600,In_518,In_646);
or U2601 (N_2601,In_357,In_785);
nor U2602 (N_2602,In_49,In_32);
or U2603 (N_2603,In_1123,In_642);
xor U2604 (N_2604,In_1292,In_865);
nor U2605 (N_2605,In_471,In_353);
and U2606 (N_2606,In_808,In_1452);
or U2607 (N_2607,In_420,In_1051);
nand U2608 (N_2608,In_659,In_657);
or U2609 (N_2609,In_1046,In_1119);
nor U2610 (N_2610,In_741,In_638);
nor U2611 (N_2611,In_845,In_365);
nor U2612 (N_2612,In_437,In_529);
nand U2613 (N_2613,In_1234,In_135);
nand U2614 (N_2614,In_575,In_733);
xor U2615 (N_2615,In_567,In_1250);
nand U2616 (N_2616,In_1258,In_411);
or U2617 (N_2617,In_889,In_333);
or U2618 (N_2618,In_136,In_321);
or U2619 (N_2619,In_422,In_1064);
or U2620 (N_2620,In_733,In_428);
nor U2621 (N_2621,In_311,In_210);
and U2622 (N_2622,In_1256,In_432);
nor U2623 (N_2623,In_607,In_903);
or U2624 (N_2624,In_524,In_336);
xor U2625 (N_2625,In_1310,In_631);
or U2626 (N_2626,In_475,In_32);
or U2627 (N_2627,In_993,In_932);
and U2628 (N_2628,In_930,In_1126);
nor U2629 (N_2629,In_485,In_902);
or U2630 (N_2630,In_1197,In_840);
nor U2631 (N_2631,In_1268,In_511);
nor U2632 (N_2632,In_899,In_1428);
xor U2633 (N_2633,In_313,In_1204);
nand U2634 (N_2634,In_1151,In_242);
nor U2635 (N_2635,In_402,In_508);
or U2636 (N_2636,In_611,In_730);
and U2637 (N_2637,In_369,In_579);
or U2638 (N_2638,In_377,In_511);
xnor U2639 (N_2639,In_985,In_1181);
xnor U2640 (N_2640,In_424,In_295);
nand U2641 (N_2641,In_820,In_172);
and U2642 (N_2642,In_573,In_454);
and U2643 (N_2643,In_1435,In_396);
or U2644 (N_2644,In_874,In_528);
or U2645 (N_2645,In_131,In_303);
xor U2646 (N_2646,In_455,In_526);
xor U2647 (N_2647,In_1047,In_1184);
xnor U2648 (N_2648,In_719,In_374);
nand U2649 (N_2649,In_29,In_398);
nor U2650 (N_2650,In_692,In_401);
nand U2651 (N_2651,In_312,In_1024);
and U2652 (N_2652,In_975,In_1202);
and U2653 (N_2653,In_382,In_1241);
nor U2654 (N_2654,In_785,In_244);
nand U2655 (N_2655,In_576,In_1246);
or U2656 (N_2656,In_871,In_1267);
or U2657 (N_2657,In_133,In_373);
or U2658 (N_2658,In_585,In_1454);
nand U2659 (N_2659,In_1195,In_683);
or U2660 (N_2660,In_54,In_1247);
xnor U2661 (N_2661,In_13,In_1117);
nand U2662 (N_2662,In_10,In_113);
or U2663 (N_2663,In_736,In_141);
or U2664 (N_2664,In_1306,In_232);
xnor U2665 (N_2665,In_18,In_1141);
nand U2666 (N_2666,In_840,In_1389);
nor U2667 (N_2667,In_705,In_94);
and U2668 (N_2668,In_1466,In_1190);
xnor U2669 (N_2669,In_783,In_1459);
or U2670 (N_2670,In_719,In_591);
and U2671 (N_2671,In_46,In_753);
or U2672 (N_2672,In_157,In_424);
nand U2673 (N_2673,In_924,In_593);
nand U2674 (N_2674,In_174,In_84);
nand U2675 (N_2675,In_225,In_1410);
nand U2676 (N_2676,In_1469,In_959);
or U2677 (N_2677,In_1203,In_248);
and U2678 (N_2678,In_439,In_665);
nor U2679 (N_2679,In_233,In_473);
or U2680 (N_2680,In_44,In_1056);
or U2681 (N_2681,In_647,In_516);
nor U2682 (N_2682,In_576,In_1488);
nand U2683 (N_2683,In_570,In_187);
xor U2684 (N_2684,In_1452,In_372);
and U2685 (N_2685,In_398,In_644);
xnor U2686 (N_2686,In_752,In_1350);
and U2687 (N_2687,In_397,In_1437);
nor U2688 (N_2688,In_937,In_1234);
xnor U2689 (N_2689,In_382,In_943);
nor U2690 (N_2690,In_662,In_1016);
nand U2691 (N_2691,In_1085,In_1274);
nor U2692 (N_2692,In_329,In_803);
nor U2693 (N_2693,In_7,In_312);
nor U2694 (N_2694,In_549,In_52);
and U2695 (N_2695,In_78,In_695);
xnor U2696 (N_2696,In_414,In_1437);
and U2697 (N_2697,In_1060,In_1432);
nand U2698 (N_2698,In_1021,In_1235);
nor U2699 (N_2699,In_321,In_841);
or U2700 (N_2700,In_66,In_735);
nand U2701 (N_2701,In_911,In_1185);
nor U2702 (N_2702,In_15,In_1313);
or U2703 (N_2703,In_933,In_842);
xor U2704 (N_2704,In_1057,In_5);
or U2705 (N_2705,In_772,In_1467);
nor U2706 (N_2706,In_305,In_235);
or U2707 (N_2707,In_1413,In_394);
and U2708 (N_2708,In_1214,In_143);
xor U2709 (N_2709,In_585,In_875);
or U2710 (N_2710,In_859,In_1229);
nand U2711 (N_2711,In_624,In_292);
xor U2712 (N_2712,In_1227,In_454);
and U2713 (N_2713,In_409,In_747);
or U2714 (N_2714,In_254,In_859);
and U2715 (N_2715,In_1349,In_1376);
nand U2716 (N_2716,In_675,In_378);
or U2717 (N_2717,In_1282,In_1269);
nor U2718 (N_2718,In_1059,In_744);
nor U2719 (N_2719,In_177,In_1144);
and U2720 (N_2720,In_1172,In_46);
or U2721 (N_2721,In_1211,In_483);
xor U2722 (N_2722,In_90,In_810);
or U2723 (N_2723,In_621,In_235);
and U2724 (N_2724,In_7,In_579);
nor U2725 (N_2725,In_1277,In_829);
nor U2726 (N_2726,In_658,In_25);
or U2727 (N_2727,In_1444,In_220);
nor U2728 (N_2728,In_1374,In_438);
xnor U2729 (N_2729,In_493,In_1246);
nand U2730 (N_2730,In_833,In_351);
nor U2731 (N_2731,In_1336,In_798);
xnor U2732 (N_2732,In_1052,In_281);
nand U2733 (N_2733,In_470,In_1224);
and U2734 (N_2734,In_1255,In_741);
nand U2735 (N_2735,In_183,In_683);
nand U2736 (N_2736,In_32,In_374);
and U2737 (N_2737,In_1184,In_1243);
or U2738 (N_2738,In_1104,In_265);
and U2739 (N_2739,In_705,In_1011);
xnor U2740 (N_2740,In_799,In_5);
nor U2741 (N_2741,In_1123,In_1214);
and U2742 (N_2742,In_285,In_359);
xnor U2743 (N_2743,In_580,In_547);
and U2744 (N_2744,In_1492,In_328);
nor U2745 (N_2745,In_1369,In_847);
or U2746 (N_2746,In_21,In_379);
xor U2747 (N_2747,In_254,In_1376);
nand U2748 (N_2748,In_683,In_1358);
or U2749 (N_2749,In_186,In_1315);
nand U2750 (N_2750,In_451,In_251);
and U2751 (N_2751,In_1419,In_1047);
or U2752 (N_2752,In_1232,In_1383);
nand U2753 (N_2753,In_1326,In_922);
or U2754 (N_2754,In_23,In_356);
and U2755 (N_2755,In_353,In_690);
nand U2756 (N_2756,In_276,In_1378);
xnor U2757 (N_2757,In_1300,In_1089);
and U2758 (N_2758,In_829,In_456);
xor U2759 (N_2759,In_672,In_1368);
nand U2760 (N_2760,In_144,In_523);
xor U2761 (N_2761,In_1301,In_1477);
or U2762 (N_2762,In_1059,In_965);
nand U2763 (N_2763,In_826,In_814);
nor U2764 (N_2764,In_205,In_1457);
and U2765 (N_2765,In_1467,In_908);
nor U2766 (N_2766,In_519,In_366);
xor U2767 (N_2767,In_790,In_1414);
or U2768 (N_2768,In_194,In_1266);
xnor U2769 (N_2769,In_222,In_775);
nand U2770 (N_2770,In_752,In_498);
or U2771 (N_2771,In_589,In_657);
and U2772 (N_2772,In_332,In_956);
nor U2773 (N_2773,In_348,In_1010);
and U2774 (N_2774,In_1045,In_978);
nor U2775 (N_2775,In_492,In_1357);
xnor U2776 (N_2776,In_385,In_270);
and U2777 (N_2777,In_737,In_690);
xor U2778 (N_2778,In_952,In_222);
and U2779 (N_2779,In_920,In_442);
xnor U2780 (N_2780,In_285,In_391);
xor U2781 (N_2781,In_1470,In_1395);
and U2782 (N_2782,In_1191,In_344);
nor U2783 (N_2783,In_665,In_596);
xnor U2784 (N_2784,In_510,In_65);
or U2785 (N_2785,In_340,In_1437);
nor U2786 (N_2786,In_461,In_331);
xor U2787 (N_2787,In_661,In_1169);
nor U2788 (N_2788,In_269,In_667);
nor U2789 (N_2789,In_519,In_972);
or U2790 (N_2790,In_1092,In_554);
or U2791 (N_2791,In_239,In_1353);
or U2792 (N_2792,In_1003,In_1259);
nand U2793 (N_2793,In_942,In_791);
and U2794 (N_2794,In_1237,In_985);
and U2795 (N_2795,In_1306,In_759);
and U2796 (N_2796,In_1001,In_1401);
nor U2797 (N_2797,In_625,In_1028);
nand U2798 (N_2798,In_1122,In_914);
xor U2799 (N_2799,In_1259,In_564);
nor U2800 (N_2800,In_1270,In_458);
nor U2801 (N_2801,In_1041,In_737);
xnor U2802 (N_2802,In_998,In_356);
xor U2803 (N_2803,In_246,In_217);
nor U2804 (N_2804,In_457,In_1125);
and U2805 (N_2805,In_99,In_676);
or U2806 (N_2806,In_1291,In_1315);
nor U2807 (N_2807,In_798,In_586);
and U2808 (N_2808,In_525,In_190);
or U2809 (N_2809,In_93,In_1412);
or U2810 (N_2810,In_896,In_605);
nor U2811 (N_2811,In_1034,In_1372);
nor U2812 (N_2812,In_477,In_1036);
or U2813 (N_2813,In_277,In_285);
or U2814 (N_2814,In_1473,In_30);
xnor U2815 (N_2815,In_556,In_655);
and U2816 (N_2816,In_1487,In_1308);
nand U2817 (N_2817,In_544,In_1446);
xor U2818 (N_2818,In_1220,In_12);
and U2819 (N_2819,In_530,In_1035);
nand U2820 (N_2820,In_956,In_1046);
xor U2821 (N_2821,In_1344,In_625);
or U2822 (N_2822,In_935,In_1220);
nor U2823 (N_2823,In_530,In_425);
or U2824 (N_2824,In_864,In_1106);
nand U2825 (N_2825,In_258,In_414);
or U2826 (N_2826,In_409,In_589);
nand U2827 (N_2827,In_1142,In_527);
nand U2828 (N_2828,In_446,In_244);
xnor U2829 (N_2829,In_409,In_114);
xor U2830 (N_2830,In_720,In_966);
nor U2831 (N_2831,In_142,In_996);
and U2832 (N_2832,In_964,In_1230);
nor U2833 (N_2833,In_603,In_1295);
nand U2834 (N_2834,In_88,In_886);
or U2835 (N_2835,In_205,In_545);
and U2836 (N_2836,In_876,In_381);
xnor U2837 (N_2837,In_880,In_562);
nand U2838 (N_2838,In_1258,In_709);
nand U2839 (N_2839,In_1340,In_297);
nand U2840 (N_2840,In_1221,In_257);
or U2841 (N_2841,In_1406,In_1490);
nand U2842 (N_2842,In_1280,In_285);
or U2843 (N_2843,In_1210,In_598);
nand U2844 (N_2844,In_509,In_1489);
xor U2845 (N_2845,In_701,In_1315);
or U2846 (N_2846,In_1021,In_453);
nand U2847 (N_2847,In_943,In_1049);
xnor U2848 (N_2848,In_669,In_117);
or U2849 (N_2849,In_117,In_950);
or U2850 (N_2850,In_1096,In_1284);
nor U2851 (N_2851,In_232,In_107);
or U2852 (N_2852,In_1320,In_289);
nand U2853 (N_2853,In_1273,In_896);
and U2854 (N_2854,In_89,In_230);
or U2855 (N_2855,In_656,In_267);
xor U2856 (N_2856,In_1296,In_695);
xor U2857 (N_2857,In_958,In_1035);
nor U2858 (N_2858,In_437,In_841);
or U2859 (N_2859,In_1178,In_309);
xnor U2860 (N_2860,In_115,In_48);
nor U2861 (N_2861,In_63,In_663);
and U2862 (N_2862,In_474,In_898);
and U2863 (N_2863,In_550,In_1185);
nor U2864 (N_2864,In_1069,In_1057);
or U2865 (N_2865,In_999,In_1406);
nand U2866 (N_2866,In_1412,In_473);
nor U2867 (N_2867,In_1392,In_1332);
nor U2868 (N_2868,In_1285,In_499);
nor U2869 (N_2869,In_860,In_1468);
or U2870 (N_2870,In_1083,In_1328);
and U2871 (N_2871,In_788,In_743);
or U2872 (N_2872,In_1199,In_1224);
nor U2873 (N_2873,In_948,In_372);
nor U2874 (N_2874,In_501,In_980);
nand U2875 (N_2875,In_700,In_920);
nand U2876 (N_2876,In_130,In_1057);
and U2877 (N_2877,In_734,In_1181);
nor U2878 (N_2878,In_1464,In_647);
nor U2879 (N_2879,In_1443,In_1181);
and U2880 (N_2880,In_505,In_1050);
nor U2881 (N_2881,In_782,In_1111);
nor U2882 (N_2882,In_48,In_1272);
nor U2883 (N_2883,In_892,In_174);
nor U2884 (N_2884,In_1384,In_1289);
nand U2885 (N_2885,In_837,In_1398);
nand U2886 (N_2886,In_159,In_677);
xor U2887 (N_2887,In_713,In_1311);
nor U2888 (N_2888,In_313,In_881);
nand U2889 (N_2889,In_828,In_980);
xnor U2890 (N_2890,In_652,In_1346);
and U2891 (N_2891,In_767,In_183);
xor U2892 (N_2892,In_1299,In_208);
xor U2893 (N_2893,In_1004,In_1072);
nand U2894 (N_2894,In_547,In_261);
or U2895 (N_2895,In_930,In_964);
or U2896 (N_2896,In_837,In_627);
and U2897 (N_2897,In_696,In_654);
xnor U2898 (N_2898,In_154,In_259);
nand U2899 (N_2899,In_474,In_1014);
xor U2900 (N_2900,In_83,In_1149);
nand U2901 (N_2901,In_1149,In_1342);
nor U2902 (N_2902,In_1118,In_684);
nor U2903 (N_2903,In_1380,In_276);
nor U2904 (N_2904,In_1194,In_1234);
nor U2905 (N_2905,In_178,In_630);
nor U2906 (N_2906,In_686,In_1078);
xnor U2907 (N_2907,In_712,In_1190);
xor U2908 (N_2908,In_981,In_1443);
and U2909 (N_2909,In_1295,In_626);
and U2910 (N_2910,In_158,In_162);
and U2911 (N_2911,In_116,In_92);
nand U2912 (N_2912,In_717,In_1098);
or U2913 (N_2913,In_118,In_440);
and U2914 (N_2914,In_1412,In_687);
xnor U2915 (N_2915,In_1261,In_34);
nor U2916 (N_2916,In_1251,In_454);
xnor U2917 (N_2917,In_296,In_188);
nand U2918 (N_2918,In_1269,In_923);
nor U2919 (N_2919,In_970,In_973);
or U2920 (N_2920,In_1305,In_806);
nor U2921 (N_2921,In_154,In_1095);
and U2922 (N_2922,In_623,In_1151);
and U2923 (N_2923,In_839,In_1356);
xnor U2924 (N_2924,In_1120,In_1031);
and U2925 (N_2925,In_1476,In_214);
and U2926 (N_2926,In_1004,In_584);
nand U2927 (N_2927,In_940,In_530);
or U2928 (N_2928,In_91,In_1382);
xnor U2929 (N_2929,In_81,In_1029);
xor U2930 (N_2930,In_123,In_448);
nand U2931 (N_2931,In_1289,In_370);
or U2932 (N_2932,In_377,In_1413);
or U2933 (N_2933,In_636,In_726);
xor U2934 (N_2934,In_1414,In_702);
and U2935 (N_2935,In_870,In_279);
and U2936 (N_2936,In_435,In_885);
nor U2937 (N_2937,In_1053,In_1251);
xor U2938 (N_2938,In_196,In_1017);
or U2939 (N_2939,In_252,In_1198);
and U2940 (N_2940,In_250,In_1032);
xnor U2941 (N_2941,In_1171,In_745);
nand U2942 (N_2942,In_868,In_1167);
and U2943 (N_2943,In_1113,In_682);
or U2944 (N_2944,In_426,In_587);
nand U2945 (N_2945,In_1085,In_661);
nand U2946 (N_2946,In_1041,In_470);
nor U2947 (N_2947,In_508,In_604);
xor U2948 (N_2948,In_1310,In_853);
xor U2949 (N_2949,In_449,In_292);
or U2950 (N_2950,In_453,In_1375);
or U2951 (N_2951,In_1360,In_35);
nand U2952 (N_2952,In_26,In_267);
xnor U2953 (N_2953,In_1425,In_851);
or U2954 (N_2954,In_311,In_1039);
nand U2955 (N_2955,In_1383,In_541);
xor U2956 (N_2956,In_1028,In_638);
or U2957 (N_2957,In_1457,In_1128);
or U2958 (N_2958,In_1199,In_529);
or U2959 (N_2959,In_333,In_421);
and U2960 (N_2960,In_70,In_185);
or U2961 (N_2961,In_508,In_243);
xnor U2962 (N_2962,In_437,In_1205);
or U2963 (N_2963,In_669,In_1492);
nand U2964 (N_2964,In_246,In_936);
nand U2965 (N_2965,In_877,In_380);
nand U2966 (N_2966,In_284,In_902);
nor U2967 (N_2967,In_263,In_626);
xor U2968 (N_2968,In_381,In_362);
or U2969 (N_2969,In_511,In_502);
and U2970 (N_2970,In_851,In_745);
and U2971 (N_2971,In_821,In_1068);
or U2972 (N_2972,In_997,In_1033);
xor U2973 (N_2973,In_1494,In_83);
and U2974 (N_2974,In_1497,In_1350);
nand U2975 (N_2975,In_627,In_383);
or U2976 (N_2976,In_884,In_990);
xor U2977 (N_2977,In_419,In_162);
nand U2978 (N_2978,In_1487,In_73);
nor U2979 (N_2979,In_841,In_150);
xnor U2980 (N_2980,In_1160,In_804);
and U2981 (N_2981,In_798,In_1463);
or U2982 (N_2982,In_404,In_1268);
nand U2983 (N_2983,In_720,In_866);
and U2984 (N_2984,In_945,In_496);
xnor U2985 (N_2985,In_1446,In_605);
nand U2986 (N_2986,In_225,In_515);
and U2987 (N_2987,In_523,In_1289);
xnor U2988 (N_2988,In_754,In_569);
and U2989 (N_2989,In_1290,In_291);
nor U2990 (N_2990,In_116,In_597);
and U2991 (N_2991,In_751,In_1305);
nor U2992 (N_2992,In_1472,In_415);
or U2993 (N_2993,In_963,In_143);
nor U2994 (N_2994,In_1451,In_1172);
or U2995 (N_2995,In_852,In_38);
xnor U2996 (N_2996,In_1452,In_672);
nor U2997 (N_2997,In_1058,In_666);
xnor U2998 (N_2998,In_1292,In_907);
nor U2999 (N_2999,In_573,In_941);
xor U3000 (N_3000,N_2364,N_2624);
or U3001 (N_3001,N_1062,N_2811);
xnor U3002 (N_3002,N_1301,N_2787);
or U3003 (N_3003,N_2599,N_1431);
nor U3004 (N_3004,N_1468,N_636);
or U3005 (N_3005,N_325,N_1181);
nor U3006 (N_3006,N_2637,N_603);
nand U3007 (N_3007,N_1269,N_1905);
and U3008 (N_3008,N_2050,N_1873);
and U3009 (N_3009,N_1049,N_654);
or U3010 (N_3010,N_132,N_1047);
or U3011 (N_3011,N_77,N_2259);
nor U3012 (N_3012,N_2576,N_1566);
and U3013 (N_3013,N_2081,N_1337);
xnor U3014 (N_3014,N_430,N_204);
nor U3015 (N_3015,N_2759,N_2210);
and U3016 (N_3016,N_2310,N_1563);
xor U3017 (N_3017,N_2694,N_352);
or U3018 (N_3018,N_1981,N_1282);
or U3019 (N_3019,N_1613,N_1536);
xor U3020 (N_3020,N_2837,N_1291);
and U3021 (N_3021,N_2418,N_1073);
xor U3022 (N_3022,N_1950,N_2286);
xor U3023 (N_3023,N_874,N_2332);
or U3024 (N_3024,N_793,N_2345);
nor U3025 (N_3025,N_2497,N_766);
xor U3026 (N_3026,N_833,N_539);
xor U3027 (N_3027,N_131,N_1874);
or U3028 (N_3028,N_2243,N_1026);
or U3029 (N_3029,N_155,N_2900);
nor U3030 (N_3030,N_2778,N_2049);
nor U3031 (N_3031,N_1076,N_1609);
or U3032 (N_3032,N_2375,N_414);
nand U3033 (N_3033,N_2663,N_1196);
or U3034 (N_3034,N_473,N_973);
nand U3035 (N_3035,N_1817,N_241);
nand U3036 (N_3036,N_2311,N_2282);
nand U3037 (N_3037,N_715,N_1596);
or U3038 (N_3038,N_836,N_2630);
nor U3039 (N_3039,N_1651,N_2413);
or U3040 (N_3040,N_537,N_2247);
or U3041 (N_3041,N_996,N_1346);
or U3042 (N_3042,N_1370,N_1868);
and U3043 (N_3043,N_908,N_2161);
and U3044 (N_3044,N_1006,N_997);
and U3045 (N_3045,N_2910,N_984);
xnor U3046 (N_3046,N_2668,N_2367);
nand U3047 (N_3047,N_1013,N_2258);
and U3048 (N_3048,N_449,N_1998);
xor U3049 (N_3049,N_2277,N_2543);
and U3050 (N_3050,N_1512,N_413);
nor U3051 (N_3051,N_2231,N_2516);
nor U3052 (N_3052,N_1434,N_2276);
nand U3053 (N_3053,N_144,N_557);
or U3054 (N_3054,N_2262,N_274);
nor U3055 (N_3055,N_1132,N_1862);
xor U3056 (N_3056,N_804,N_2739);
nand U3057 (N_3057,N_1825,N_2303);
and U3058 (N_3058,N_2388,N_145);
nor U3059 (N_3059,N_2365,N_1005);
and U3060 (N_3060,N_978,N_2132);
or U3061 (N_3061,N_444,N_1360);
xnor U3062 (N_3062,N_2895,N_2675);
xnor U3063 (N_3063,N_2008,N_1284);
xnor U3064 (N_3064,N_1451,N_2963);
nor U3065 (N_3065,N_681,N_2875);
or U3066 (N_3066,N_1593,N_2436);
nand U3067 (N_3067,N_1273,N_1015);
xor U3068 (N_3068,N_2631,N_2201);
nor U3069 (N_3069,N_2944,N_1656);
or U3070 (N_3070,N_1888,N_2325);
nand U3071 (N_3071,N_1163,N_1653);
or U3072 (N_3072,N_2239,N_2851);
xnor U3073 (N_3073,N_1352,N_545);
nor U3074 (N_3074,N_1587,N_1716);
or U3075 (N_3075,N_2578,N_2348);
and U3076 (N_3076,N_1632,N_1810);
or U3077 (N_3077,N_2241,N_1329);
nor U3078 (N_3078,N_2990,N_2584);
nor U3079 (N_3079,N_2738,N_775);
xnor U3080 (N_3080,N_2858,N_811);
or U3081 (N_3081,N_2087,N_2406);
nor U3082 (N_3082,N_1080,N_907);
nand U3083 (N_3083,N_939,N_948);
or U3084 (N_3084,N_253,N_1782);
and U3085 (N_3085,N_2692,N_2942);
xnor U3086 (N_3086,N_1664,N_2586);
or U3087 (N_3087,N_675,N_2888);
xnor U3088 (N_3088,N_2653,N_1933);
nor U3089 (N_3089,N_2076,N_2472);
nand U3090 (N_3090,N_2456,N_1991);
or U3091 (N_3091,N_612,N_930);
and U3092 (N_3092,N_1537,N_1693);
and U3093 (N_3093,N_0,N_937);
nor U3094 (N_3094,N_1450,N_2080);
and U3095 (N_3095,N_812,N_34);
and U3096 (N_3096,N_1750,N_2545);
nor U3097 (N_3097,N_938,N_2131);
nor U3098 (N_3098,N_584,N_2526);
nand U3099 (N_3099,N_2866,N_1731);
and U3100 (N_3100,N_1378,N_1619);
xnor U3101 (N_3101,N_1505,N_1361);
or U3102 (N_3102,N_1897,N_1938);
nand U3103 (N_3103,N_260,N_336);
and U3104 (N_3104,N_1177,N_1463);
nor U3105 (N_3105,N_363,N_1447);
xor U3106 (N_3106,N_236,N_1719);
nand U3107 (N_3107,N_1717,N_1151);
xor U3108 (N_3108,N_983,N_747);
or U3109 (N_3109,N_1327,N_882);
nand U3110 (N_3110,N_2434,N_101);
and U3111 (N_3111,N_1105,N_1866);
or U3112 (N_3112,N_492,N_29);
nand U3113 (N_3113,N_1338,N_2224);
nand U3114 (N_3114,N_2640,N_374);
and U3115 (N_3115,N_2916,N_2063);
nand U3116 (N_3116,N_900,N_1009);
xnor U3117 (N_3117,N_1645,N_921);
nand U3118 (N_3118,N_2533,N_1698);
or U3119 (N_3119,N_895,N_1966);
nor U3120 (N_3120,N_1445,N_1772);
nand U3121 (N_3121,N_2819,N_849);
or U3122 (N_3122,N_1024,N_2935);
nor U3123 (N_3123,N_2902,N_623);
or U3124 (N_3124,N_1002,N_1161);
or U3125 (N_3125,N_2240,N_1584);
or U3126 (N_3126,N_224,N_2335);
and U3127 (N_3127,N_661,N_1977);
xnor U3128 (N_3128,N_1150,N_1108);
nand U3129 (N_3129,N_2883,N_2821);
and U3130 (N_3130,N_1003,N_110);
xor U3131 (N_3131,N_49,N_980);
nor U3132 (N_3132,N_2357,N_2577);
or U3133 (N_3133,N_1285,N_2251);
and U3134 (N_3134,N_2220,N_510);
xnor U3135 (N_3135,N_1236,N_2481);
and U3136 (N_3136,N_1046,N_2018);
and U3137 (N_3137,N_2077,N_749);
xor U3138 (N_3138,N_2905,N_318);
nand U3139 (N_3139,N_861,N_472);
and U3140 (N_3140,N_69,N_72);
nand U3141 (N_3141,N_1552,N_659);
or U3142 (N_3142,N_474,N_91);
and U3143 (N_3143,N_2029,N_560);
xnor U3144 (N_3144,N_2728,N_2130);
nand U3145 (N_3145,N_2295,N_656);
and U3146 (N_3146,N_421,N_1303);
or U3147 (N_3147,N_1854,N_2451);
nand U3148 (N_3148,N_1482,N_150);
or U3149 (N_3149,N_1790,N_2322);
nand U3150 (N_3150,N_1959,N_807);
nor U3151 (N_3151,N_1328,N_2566);
and U3152 (N_3152,N_1785,N_156);
nand U3153 (N_3153,N_169,N_1570);
or U3154 (N_3154,N_2670,N_962);
or U3155 (N_3155,N_1559,N_329);
nor U3156 (N_3156,N_736,N_166);
nor U3157 (N_3157,N_1092,N_1100);
xnor U3158 (N_3158,N_2094,N_203);
and U3159 (N_3159,N_1947,N_1680);
nand U3160 (N_3160,N_2710,N_279);
xor U3161 (N_3161,N_1562,N_196);
and U3162 (N_3162,N_1836,N_2312);
and U3163 (N_3163,N_2391,N_290);
xor U3164 (N_3164,N_323,N_1531);
nor U3165 (N_3165,N_1783,N_1377);
or U3166 (N_3166,N_885,N_614);
and U3167 (N_3167,N_2891,N_1726);
nand U3168 (N_3168,N_2736,N_1744);
or U3169 (N_3169,N_696,N_558);
or U3170 (N_3170,N_2560,N_1052);
xor U3171 (N_3171,N_1247,N_870);
xor U3172 (N_3172,N_167,N_338);
nor U3173 (N_3173,N_229,N_2849);
nor U3174 (N_3174,N_2880,N_1391);
nor U3175 (N_3175,N_2832,N_1980);
or U3176 (N_3176,N_129,N_2989);
nor U3177 (N_3177,N_1425,N_2124);
xor U3178 (N_3178,N_1703,N_2721);
and U3179 (N_3179,N_1637,N_918);
nor U3180 (N_3180,N_963,N_2030);
nor U3181 (N_3181,N_1676,N_852);
or U3182 (N_3182,N_238,N_187);
xor U3183 (N_3183,N_2592,N_2917);
nand U3184 (N_3184,N_1701,N_118);
xnor U3185 (N_3185,N_2643,N_476);
xor U3186 (N_3186,N_124,N_1223);
xor U3187 (N_3187,N_563,N_867);
nand U3188 (N_3188,N_506,N_662);
and U3189 (N_3189,N_2152,N_1294);
nand U3190 (N_3190,N_810,N_1452);
nor U3191 (N_3191,N_1381,N_1398);
xnor U3192 (N_3192,N_746,N_1979);
xnor U3193 (N_3193,N_1758,N_134);
xnor U3194 (N_3194,N_1277,N_1458);
nand U3195 (N_3195,N_1925,N_2625);
xnor U3196 (N_3196,N_2137,N_2458);
nand U3197 (N_3197,N_68,N_517);
and U3198 (N_3198,N_1475,N_1626);
nand U3199 (N_3199,N_1513,N_2818);
nor U3200 (N_3200,N_1364,N_546);
and U3201 (N_3201,N_718,N_1509);
xnor U3202 (N_3202,N_291,N_2657);
xnor U3203 (N_3203,N_1521,N_1226);
and U3204 (N_3204,N_720,N_19);
and U3205 (N_3205,N_1467,N_360);
xor U3206 (N_3206,N_2198,N_1295);
xor U3207 (N_3207,N_647,N_1323);
or U3208 (N_3208,N_1876,N_582);
nor U3209 (N_3209,N_1834,N_1707);
nor U3210 (N_3210,N_1160,N_1274);
or U3211 (N_3211,N_1634,N_934);
nor U3212 (N_3212,N_2001,N_1554);
nor U3213 (N_3213,N_1685,N_2429);
nand U3214 (N_3214,N_1743,N_2428);
and U3215 (N_3215,N_2278,N_2998);
nand U3216 (N_3216,N_1188,N_1110);
or U3217 (N_3217,N_2279,N_2177);
and U3218 (N_3218,N_1179,N_1963);
and U3219 (N_3219,N_2219,N_2767);
or U3220 (N_3220,N_2857,N_579);
xnor U3221 (N_3221,N_240,N_1881);
nor U3222 (N_3222,N_2816,N_298);
and U3223 (N_3223,N_2508,N_742);
nand U3224 (N_3224,N_2695,N_768);
and U3225 (N_3225,N_1212,N_1692);
nand U3226 (N_3226,N_864,N_445);
nand U3227 (N_3227,N_442,N_1837);
or U3228 (N_3228,N_2542,N_1912);
and U3229 (N_3229,N_95,N_2708);
and U3230 (N_3230,N_1745,N_572);
xnor U3231 (N_3231,N_2300,N_998);
nand U3232 (N_3232,N_1215,N_763);
nand U3233 (N_3233,N_2506,N_1879);
nor U3234 (N_3234,N_2366,N_25);
or U3235 (N_3235,N_2515,N_1671);
xnor U3236 (N_3236,N_2459,N_2709);
or U3237 (N_3237,N_2043,N_2985);
nand U3238 (N_3238,N_2476,N_188);
nand U3239 (N_3239,N_932,N_1638);
nor U3240 (N_3240,N_691,N_11);
or U3241 (N_3241,N_799,N_1522);
or U3242 (N_3242,N_1846,N_692);
and U3243 (N_3243,N_2536,N_2394);
and U3244 (N_3244,N_2652,N_2889);
nor U3245 (N_3245,N_1845,N_2314);
xnor U3246 (N_3246,N_1826,N_2794);
or U3247 (N_3247,N_1889,N_2575);
and U3248 (N_3248,N_2997,N_1043);
or U3249 (N_3249,N_2800,N_2133);
or U3250 (N_3250,N_708,N_1017);
or U3251 (N_3251,N_1548,N_1036);
nor U3252 (N_3252,N_1812,N_2809);
and U3253 (N_3253,N_2119,N_2184);
xor U3254 (N_3254,N_1891,N_1436);
nor U3255 (N_3255,N_1048,N_780);
nand U3256 (N_3256,N_941,N_2150);
nand U3257 (N_3257,N_2923,N_1034);
nand U3258 (N_3258,N_586,N_2981);
xnor U3259 (N_3259,N_1771,N_1582);
or U3260 (N_3260,N_2071,N_898);
and U3261 (N_3261,N_1464,N_2101);
or U3262 (N_3262,N_2272,N_803);
xnor U3263 (N_3263,N_2127,N_1984);
nand U3264 (N_3264,N_2423,N_2339);
or U3265 (N_3265,N_109,N_827);
xor U3266 (N_3266,N_1838,N_2301);
xnor U3267 (N_3267,N_2091,N_1121);
nand U3268 (N_3268,N_1324,N_2323);
nor U3269 (N_3269,N_757,N_1890);
nand U3270 (N_3270,N_1604,N_548);
and U3271 (N_3271,N_2245,N_2912);
nand U3272 (N_3272,N_218,N_1350);
or U3273 (N_3273,N_1202,N_308);
xor U3274 (N_3274,N_503,N_2052);
and U3275 (N_3275,N_24,N_295);
nor U3276 (N_3276,N_1694,N_2382);
nand U3277 (N_3277,N_967,N_2975);
nand U3278 (N_3278,N_1305,N_1008);
xor U3279 (N_3279,N_819,N_159);
nand U3280 (N_3280,N_2765,N_2209);
nand U3281 (N_3281,N_1710,N_434);
or U3282 (N_3282,N_2825,N_2351);
nand U3283 (N_3283,N_2878,N_2215);
or U3284 (N_3284,N_634,N_773);
and U3285 (N_3285,N_464,N_1753);
xor U3286 (N_3286,N_1166,N_147);
or U3287 (N_3287,N_1820,N_890);
and U3288 (N_3288,N_1037,N_1066);
or U3289 (N_3289,N_470,N_1715);
and U3290 (N_3290,N_956,N_562);
and U3291 (N_3291,N_2532,N_1589);
and U3292 (N_3292,N_2984,N_1235);
and U3293 (N_3293,N_1614,N_1799);
nand U3294 (N_3294,N_912,N_1886);
xor U3295 (N_3295,N_2117,N_1767);
or U3296 (N_3296,N_287,N_423);
and U3297 (N_3297,N_2733,N_82);
nor U3298 (N_3298,N_1298,N_2267);
nand U3299 (N_3299,N_754,N_100);
and U3300 (N_3300,N_1786,N_1978);
nand U3301 (N_3301,N_2467,N_1416);
and U3302 (N_3302,N_2791,N_41);
xnor U3303 (N_3303,N_349,N_2664);
or U3304 (N_3304,N_893,N_1276);
xnor U3305 (N_3305,N_1387,N_2494);
and U3306 (N_3306,N_1293,N_1004);
nor U3307 (N_3307,N_2945,N_1631);
or U3308 (N_3308,N_972,N_1109);
nor U3309 (N_3309,N_2349,N_1059);
and U3310 (N_3310,N_2783,N_2088);
or U3311 (N_3311,N_1677,N_2387);
and U3312 (N_3312,N_629,N_2569);
nand U3313 (N_3313,N_2069,N_1090);
nand U3314 (N_3314,N_1155,N_2606);
nor U3315 (N_3315,N_2060,N_632);
and U3316 (N_3316,N_142,N_2737);
nand U3317 (N_3317,N_2174,N_2141);
nor U3318 (N_3318,N_797,N_2971);
or U3319 (N_3319,N_304,N_2824);
xnor U3320 (N_3320,N_2949,N_2462);
and U3321 (N_3321,N_2405,N_1571);
nand U3322 (N_3322,N_2954,N_1126);
nand U3323 (N_3323,N_354,N_407);
xor U3324 (N_3324,N_2919,N_745);
and U3325 (N_3325,N_378,N_1779);
or U3326 (N_3326,N_249,N_478);
xnor U3327 (N_3327,N_1896,N_1898);
nand U3328 (N_3328,N_2730,N_99);
xor U3329 (N_3329,N_2774,N_2498);
or U3330 (N_3330,N_1757,N_1164);
xor U3331 (N_3331,N_488,N_751);
nor U3332 (N_3332,N_504,N_2877);
or U3333 (N_3333,N_1870,N_2143);
nor U3334 (N_3334,N_1479,N_471);
or U3335 (N_3335,N_2768,N_1099);
nor U3336 (N_3336,N_2823,N_1471);
and U3337 (N_3337,N_2014,N_2659);
nor U3338 (N_3338,N_2622,N_2126);
nor U3339 (N_3339,N_197,N_831);
nand U3340 (N_3340,N_243,N_1818);
nor U3341 (N_3341,N_313,N_834);
and U3342 (N_3342,N_1374,N_1203);
nor U3343 (N_3343,N_2782,N_2772);
or U3344 (N_3344,N_657,N_735);
and U3345 (N_3345,N_905,N_1987);
or U3346 (N_3346,N_271,N_2781);
nand U3347 (N_3347,N_2621,N_2750);
xor U3348 (N_3348,N_711,N_987);
nand U3349 (N_3349,N_2792,N_2333);
or U3350 (N_3350,N_2068,N_141);
xnor U3351 (N_3351,N_2978,N_1275);
and U3352 (N_3352,N_200,N_2414);
xnor U3353 (N_3353,N_1228,N_642);
nor U3354 (N_3354,N_2899,N_2965);
xor U3355 (N_3355,N_2847,N_2072);
or U3356 (N_3356,N_2714,N_2612);
xor U3357 (N_3357,N_2745,N_521);
or U3358 (N_3358,N_1515,N_1601);
or U3359 (N_3359,N_2031,N_2956);
or U3360 (N_3360,N_1413,N_722);
and U3361 (N_3361,N_565,N_192);
xnor U3362 (N_3362,N_880,N_1764);
nand U3363 (N_3363,N_276,N_981);
and U3364 (N_3364,N_1127,N_961);
xnor U3365 (N_3365,N_1201,N_1832);
or U3366 (N_3366,N_2962,N_1496);
xnor U3367 (N_3367,N_2761,N_952);
nor U3368 (N_3368,N_1107,N_126);
nor U3369 (N_3369,N_2672,N_1678);
nand U3370 (N_3370,N_1053,N_2921);
xor U3371 (N_3371,N_1233,N_2249);
xor U3372 (N_3372,N_2802,N_2273);
or U3373 (N_3373,N_319,N_2488);
nor U3374 (N_3374,N_252,N_2070);
nand U3375 (N_3375,N_2535,N_1712);
nor U3376 (N_3376,N_2810,N_1089);
or U3377 (N_3377,N_2013,N_705);
nand U3378 (N_3378,N_2884,N_1894);
nand U3379 (N_3379,N_2109,N_28);
and U3380 (N_3380,N_1795,N_168);
nand U3381 (N_3381,N_515,N_1390);
and U3382 (N_3382,N_270,N_2951);
and U3383 (N_3383,N_1306,N_222);
and U3384 (N_3384,N_2192,N_2107);
or U3385 (N_3385,N_2696,N_2324);
nand U3386 (N_3386,N_1939,N_2521);
xnor U3387 (N_3387,N_2281,N_1935);
or U3388 (N_3388,N_1639,N_2399);
or U3389 (N_3389,N_2960,N_486);
nand U3390 (N_3390,N_412,N_2505);
nor U3391 (N_3391,N_2235,N_2541);
nor U3392 (N_3392,N_876,N_2635);
xor U3393 (N_3393,N_1518,N_424);
xnor U3394 (N_3394,N_501,N_97);
xor U3395 (N_3395,N_945,N_399);
nor U3396 (N_3396,N_50,N_2595);
nand U3397 (N_3397,N_160,N_1794);
nand U3398 (N_3398,N_2534,N_2716);
nor U3399 (N_3399,N_346,N_112);
nand U3400 (N_3400,N_543,N_1180);
and U3401 (N_3401,N_410,N_1621);
nand U3402 (N_3402,N_267,N_2105);
xor U3403 (N_3403,N_2051,N_863);
nand U3404 (N_3404,N_2118,N_2442);
and U3405 (N_3405,N_601,N_2552);
nand U3406 (N_3406,N_2667,N_2510);
nand U3407 (N_3407,N_2142,N_456);
nor U3408 (N_3408,N_1516,N_1994);
and U3409 (N_3409,N_1594,N_739);
or U3410 (N_3410,N_2855,N_2961);
nand U3411 (N_3411,N_703,N_2529);
or U3412 (N_3412,N_625,N_630);
xor U3413 (N_3413,N_2826,N_1281);
nand U3414 (N_3414,N_2045,N_1895);
xor U3415 (N_3415,N_1194,N_390);
and U3416 (N_3416,N_48,N_246);
nand U3417 (N_3417,N_850,N_1529);
and U3418 (N_3418,N_1386,N_469);
xor U3419 (N_3419,N_2615,N_608);
and U3420 (N_3420,N_2844,N_949);
xnor U3421 (N_3421,N_2502,N_1357);
nor U3422 (N_3422,N_2645,N_2618);
nand U3423 (N_3423,N_1462,N_1747);
and U3424 (N_3424,N_358,N_2073);
nor U3425 (N_3425,N_261,N_2334);
nor U3426 (N_3426,N_1565,N_440);
nor U3427 (N_3427,N_993,N_302);
and U3428 (N_3428,N_965,N_2934);
nor U3429 (N_3429,N_2331,N_2634);
xnor U3430 (N_3430,N_225,N_646);
and U3431 (N_3431,N_2041,N_1214);
xnor U3432 (N_3432,N_2138,N_960);
nor U3433 (N_3433,N_2330,N_2165);
xnor U3434 (N_3434,N_1261,N_2197);
or U3435 (N_3435,N_2540,N_2892);
nand U3436 (N_3436,N_1469,N_2389);
xnor U3437 (N_3437,N_578,N_2248);
or U3438 (N_3438,N_1579,N_93);
nand U3439 (N_3439,N_928,N_1455);
nand U3440 (N_3440,N_2589,N_536);
or U3441 (N_3441,N_1941,N_633);
and U3442 (N_3442,N_1259,N_1229);
nand U3443 (N_3443,N_2038,N_2449);
and U3444 (N_3444,N_2565,N_2773);
and U3445 (N_3445,N_2553,N_36);
or U3446 (N_3446,N_2607,N_1474);
xor U3447 (N_3447,N_63,N_1489);
or U3448 (N_3448,N_2438,N_214);
or U3449 (N_3449,N_2003,N_1945);
or U3450 (N_3450,N_2355,N_458);
or U3451 (N_3451,N_724,N_208);
nor U3452 (N_3452,N_1333,N_695);
or U3453 (N_3453,N_289,N_726);
nor U3454 (N_3454,N_2676,N_1511);
nand U3455 (N_3455,N_1924,N_2901);
nor U3456 (N_3456,N_2724,N_1849);
nor U3457 (N_3457,N_835,N_2839);
xor U3458 (N_3458,N_2100,N_163);
and U3459 (N_3459,N_1453,N_250);
nand U3460 (N_3460,N_610,N_334);
nand U3461 (N_3461,N_600,N_1213);
or U3462 (N_3462,N_2308,N_1128);
or U3463 (N_3463,N_1191,N_2102);
or U3464 (N_3464,N_2830,N_2946);
and U3465 (N_3465,N_1646,N_1953);
nor U3466 (N_3466,N_817,N_326);
nand U3467 (N_3467,N_499,N_1220);
and U3468 (N_3468,N_1465,N_1131);
and U3469 (N_3469,N_1063,N_771);
nor U3470 (N_3470,N_1476,N_2715);
or U3471 (N_3471,N_2950,N_1407);
or U3472 (N_3472,N_1877,N_1486);
nor U3473 (N_3473,N_2316,N_2200);
nand U3474 (N_3474,N_830,N_1354);
nor U3475 (N_3475,N_1084,N_1936);
and U3476 (N_3476,N_2170,N_678);
xnor U3477 (N_3477,N_483,N_1777);
nand U3478 (N_3478,N_1755,N_2354);
nor U3479 (N_3479,N_1492,N_628);
and U3480 (N_3480,N_2591,N_712);
xor U3481 (N_3481,N_2964,N_2120);
and U3482 (N_3482,N_2854,N_2948);
or U3483 (N_3483,N_756,N_2583);
nor U3484 (N_3484,N_2993,N_2865);
nor U3485 (N_3485,N_10,N_688);
xnor U3486 (N_3486,N_1665,N_2374);
and U3487 (N_3487,N_2400,N_1330);
xnor U3488 (N_3488,N_2194,N_903);
nor U3489 (N_3489,N_1061,N_577);
nor U3490 (N_3490,N_2769,N_2539);
xnor U3491 (N_3491,N_1730,N_2597);
xor U3492 (N_3492,N_2940,N_89);
and U3493 (N_3493,N_1136,N_1580);
or U3494 (N_3494,N_2358,N_185);
xor U3495 (N_3495,N_1216,N_121);
nor U3496 (N_3496,N_299,N_1265);
xnor U3497 (N_3497,N_1137,N_2550);
nand U3498 (N_3498,N_2042,N_2157);
nand U3499 (N_3499,N_1542,N_462);
nand U3500 (N_3500,N_787,N_944);
or U3501 (N_3501,N_2493,N_940);
nor U3502 (N_3502,N_2776,N_1397);
nor U3503 (N_3503,N_1908,N_2268);
xor U3504 (N_3504,N_2690,N_1882);
xnor U3505 (N_3505,N_2315,N_2833);
nor U3506 (N_3506,N_2605,N_359);
nor U3507 (N_3507,N_2914,N_87);
xnor U3508 (N_3508,N_2288,N_832);
nand U3509 (N_3509,N_1674,N_2766);
and U3510 (N_3510,N_1075,N_2135);
xnor U3511 (N_3511,N_2430,N_664);
or U3512 (N_3512,N_1588,N_123);
nand U3513 (N_3513,N_845,N_130);
and U3514 (N_3514,N_1060,N_306);
nor U3515 (N_3515,N_602,N_538);
and U3516 (N_3516,N_1050,N_1219);
or U3517 (N_3517,N_1724,N_1493);
and U3518 (N_3518,N_674,N_1727);
nand U3519 (N_3519,N_2204,N_165);
nor U3520 (N_3520,N_1993,N_1734);
xnor U3521 (N_3521,N_2551,N_971);
and U3522 (N_3522,N_1130,N_2205);
nand U3523 (N_3523,N_1389,N_233);
and U3524 (N_3524,N_1172,N_1720);
or U3525 (N_3525,N_15,N_1932);
xnor U3526 (N_3526,N_2499,N_2372);
nor U3527 (N_3527,N_2376,N_822);
nor U3528 (N_3528,N_786,N_669);
nor U3529 (N_3529,N_2466,N_2343);
or U3530 (N_3530,N_618,N_1182);
and U3531 (N_3531,N_620,N_774);
xnor U3532 (N_3532,N_1417,N_668);
and U3533 (N_3533,N_1789,N_2626);
or U3534 (N_3534,N_2326,N_1982);
nor U3535 (N_3535,N_569,N_286);
xor U3536 (N_3536,N_1934,N_1158);
nor U3537 (N_3537,N_40,N_2427);
and U3538 (N_3538,N_2074,N_1242);
and U3539 (N_3539,N_2318,N_2214);
nor U3540 (N_3540,N_2178,N_1197);
nand U3541 (N_3541,N_2937,N_1507);
or U3542 (N_3542,N_2420,N_826);
nand U3543 (N_3543,N_2717,N_721);
nand U3544 (N_3544,N_62,N_331);
xnor U3545 (N_3545,N_1831,N_2688);
nand U3546 (N_3546,N_909,N_2411);
or U3547 (N_3547,N_593,N_855);
nand U3548 (N_3548,N_272,N_2144);
xnor U3549 (N_3549,N_247,N_1111);
or U3550 (N_3550,N_2460,N_1207);
and U3551 (N_3551,N_2448,N_1841);
or U3552 (N_3552,N_322,N_1320);
nor U3553 (N_3553,N_2876,N_764);
nor U3554 (N_3554,N_2232,N_2815);
and U3555 (N_3555,N_1114,N_1906);
xnor U3556 (N_3556,N_2004,N_1134);
nor U3557 (N_3557,N_2095,N_133);
xnor U3558 (N_3558,N_5,N_1414);
and U3559 (N_3559,N_931,N_617);
xnor U3560 (N_3560,N_2554,N_1221);
nand U3561 (N_3561,N_258,N_1018);
nor U3562 (N_3562,N_1940,N_1774);
and U3563 (N_3563,N_524,N_2629);
nand U3564 (N_3564,N_1970,N_92);
or U3565 (N_3565,N_999,N_119);
xor U3566 (N_3566,N_613,N_2202);
or U3567 (N_3567,N_666,N_886);
and U3568 (N_3568,N_991,N_658);
xnor U3569 (N_3569,N_1098,N_540);
and U3570 (N_3570,N_1178,N_2253);
xnor U3571 (N_3571,N_770,N_1667);
nand U3572 (N_3572,N_311,N_806);
or U3573 (N_3573,N_1553,N_840);
nor U3574 (N_3574,N_1550,N_1809);
nand U3575 (N_3575,N_2187,N_1278);
nand U3576 (N_3576,N_2544,N_1104);
or U3577 (N_3577,N_990,N_73);
nor U3578 (N_3578,N_1917,N_561);
or U3579 (N_3579,N_541,N_2886);
xnor U3580 (N_3580,N_2190,N_2644);
xnor U3581 (N_3581,N_2299,N_2168);
and U3582 (N_3582,N_2431,N_177);
nand U3583 (N_3583,N_1741,N_2482);
and U3584 (N_3584,N_2799,N_815);
and U3585 (N_3585,N_2154,N_1851);
or U3586 (N_3586,N_1106,N_2968);
and U3587 (N_3587,N_1392,N_877);
and U3588 (N_3588,N_1502,N_47);
or U3589 (N_3589,N_761,N_157);
and U3590 (N_3590,N_441,N_1200);
nand U3591 (N_3591,N_1538,N_2681);
and U3592 (N_3592,N_730,N_534);
or U3593 (N_3593,N_2564,N_2371);
or U3594 (N_3594,N_2735,N_2795);
or U3595 (N_3595,N_2838,N_6);
or U3596 (N_3596,N_2033,N_2939);
nor U3597 (N_3597,N_2931,N_682);
and U3598 (N_3598,N_1051,N_1395);
or U3599 (N_3599,N_959,N_2537);
nor U3600 (N_3600,N_1926,N_2729);
or U3601 (N_3601,N_2404,N_1603);
xor U3602 (N_3602,N_172,N_1367);
and U3603 (N_3603,N_2369,N_495);
or U3604 (N_3604,N_748,N_2140);
nor U3605 (N_3605,N_957,N_1319);
nor U3606 (N_3606,N_2022,N_1763);
nor U3607 (N_3607,N_1349,N_467);
xor U3608 (N_3608,N_2054,N_1690);
or U3609 (N_3609,N_958,N_741);
or U3610 (N_3610,N_704,N_1251);
xnor U3611 (N_3611,N_368,N_425);
nand U3612 (N_3612,N_1288,N_2379);
nand U3613 (N_3613,N_1776,N_1400);
xnor U3614 (N_3614,N_2421,N_1487);
nand U3615 (N_3615,N_1661,N_2148);
xnor U3616 (N_3616,N_357,N_535);
or U3617 (N_3617,N_18,N_1903);
nor U3618 (N_3618,N_2758,N_1740);
nand U3619 (N_3619,N_2867,N_2479);
or U3620 (N_3620,N_1206,N_1861);
or U3621 (N_3621,N_753,N_2518);
and U3622 (N_3622,N_285,N_714);
xnor U3623 (N_3623,N_1737,N_1919);
and U3624 (N_3624,N_255,N_2613);
and U3625 (N_3625,N_2337,N_1321);
or U3626 (N_3626,N_550,N_1956);
nand U3627 (N_3627,N_1650,N_643);
or U3628 (N_3628,N_2848,N_450);
or U3629 (N_3629,N_388,N_1765);
xor U3630 (N_3630,N_1709,N_923);
or U3631 (N_3631,N_2083,N_2872);
or U3632 (N_3632,N_175,N_523);
or U3633 (N_3633,N_369,N_401);
nand U3634 (N_3634,N_237,N_883);
nor U3635 (N_3635,N_989,N_1444);
xor U3636 (N_3636,N_427,N_316);
and U3637 (N_3637,N_1813,N_1954);
xnor U3638 (N_3638,N_2955,N_954);
xor U3639 (N_3639,N_1686,N_1103);
and U3640 (N_3640,N_2620,N_2925);
nand U3641 (N_3641,N_2410,N_111);
nand U3642 (N_3642,N_1618,N_1913);
or U3643 (N_3643,N_2727,N_1);
and U3644 (N_3644,N_2477,N_1573);
and U3645 (N_3645,N_2103,N_344);
xnor U3646 (N_3646,N_2959,N_1714);
and U3647 (N_3647,N_2058,N_750);
nand U3648 (N_3648,N_1840,N_2378);
nand U3649 (N_3649,N_280,N_1892);
nand U3650 (N_3650,N_1992,N_1844);
nor U3651 (N_3651,N_1517,N_1949);
nor U3652 (N_3652,N_1723,N_297);
and U3653 (N_3653,N_2291,N_1366);
or U3654 (N_3654,N_60,N_2034);
xnor U3655 (N_3655,N_2164,N_1124);
or U3656 (N_3656,N_404,N_1438);
nor U3657 (N_3657,N_235,N_2760);
nor U3658 (N_3658,N_1218,N_2317);
and U3659 (N_3659,N_697,N_1722);
or U3660 (N_3660,N_2520,N_65);
nor U3661 (N_3661,N_2596,N_994);
nor U3662 (N_3662,N_1426,N_2927);
xnor U3663 (N_3663,N_428,N_729);
and U3664 (N_3664,N_1410,N_2362);
nor U3665 (N_3665,N_398,N_1499);
and U3666 (N_3666,N_307,N_312);
xnor U3667 (N_3667,N_1435,N_1183);
or U3668 (N_3668,N_446,N_2044);
and U3669 (N_3669,N_2465,N_1423);
and U3670 (N_3670,N_2116,N_772);
xnor U3671 (N_3671,N_635,N_1101);
nand U3672 (N_3672,N_665,N_872);
xor U3673 (N_3673,N_2627,N_1616);
and U3674 (N_3674,N_1732,N_2556);
xor U3675 (N_3675,N_2790,N_17);
nor U3676 (N_3676,N_785,N_2723);
nand U3677 (N_3677,N_2697,N_1307);
and U3678 (N_3678,N_2037,N_1815);
xor U3679 (N_3679,N_640,N_310);
nand U3680 (N_3680,N_1788,N_1628);
nand U3681 (N_3681,N_341,N_2751);
and U3682 (N_3682,N_345,N_140);
nor U3683 (N_3683,N_2294,N_1598);
xor U3684 (N_3684,N_2475,N_529);
and U3685 (N_3685,N_1252,N_2402);
and U3686 (N_3686,N_1909,N_1199);
nor U3687 (N_3687,N_2384,N_556);
and U3688 (N_3688,N_1021,N_2039);
xnor U3689 (N_3689,N_942,N_1869);
xnor U3690 (N_3690,N_1768,N_479);
xnor U3691 (N_3691,N_881,N_955);
and U3692 (N_3692,N_936,N_1055);
and U3693 (N_3693,N_2779,N_1205);
nand U3694 (N_3694,N_1256,N_2305);
nor U3695 (N_3695,N_406,N_2725);
and U3696 (N_3696,N_1454,N_2856);
nand U3697 (N_3697,N_862,N_1793);
and U3698 (N_3698,N_220,N_1736);
nor U3699 (N_3699,N_777,N_278);
nor U3700 (N_3700,N_842,N_1687);
nor U3701 (N_3701,N_2233,N_1569);
or U3702 (N_3702,N_671,N_2911);
nor U3703 (N_3703,N_1369,N_1187);
xor U3704 (N_3704,N_2988,N_590);
and U3705 (N_3705,N_542,N_1914);
or U3706 (N_3706,N_2682,N_2489);
or U3707 (N_3707,N_396,N_1971);
nor U3708 (N_3708,N_320,N_2762);
or U3709 (N_3709,N_44,N_1696);
and U3710 (N_3710,N_30,N_227);
nor U3711 (N_3711,N_230,N_1415);
or U3712 (N_3712,N_205,N_1280);
and U3713 (N_3713,N_2179,N_2416);
and U3714 (N_3714,N_2417,N_1154);
nand U3715 (N_3715,N_1557,N_638);
xnor U3716 (N_3716,N_1466,N_327);
xor U3717 (N_3717,N_639,N_1605);
and U3718 (N_3718,N_2383,N_1976);
or U3719 (N_3719,N_1930,N_1931);
nor U3720 (N_3720,N_824,N_2065);
nor U3721 (N_3721,N_2673,N_254);
xor U3722 (N_3722,N_2234,N_1902);
nor U3723 (N_3723,N_2503,N_1962);
or U3724 (N_3724,N_2352,N_2026);
nand U3725 (N_3725,N_2099,N_2032);
and U3726 (N_3726,N_1032,N_2941);
nand U3727 (N_3727,N_2012,N_2195);
xnor U3728 (N_3728,N_1302,N_2639);
nor U3729 (N_3729,N_599,N_2992);
or U3730 (N_3730,N_1612,N_1057);
and U3731 (N_3731,N_699,N_2704);
nand U3732 (N_3732,N_2808,N_1960);
and U3733 (N_3733,N_2495,N_2859);
or U3734 (N_3734,N_1983,N_108);
nand U3735 (N_3735,N_1097,N_1640);
and U3736 (N_3736,N_294,N_210);
nand U3737 (N_3737,N_1490,N_911);
nor U3738 (N_3738,N_792,N_2982);
nand U3739 (N_3739,N_2307,N_888);
xnor U3740 (N_3740,N_2678,N_21);
or U3741 (N_3741,N_371,N_1478);
nand U3742 (N_3742,N_216,N_2079);
or U3743 (N_3743,N_380,N_333);
or U3744 (N_3744,N_892,N_1042);
nor U3745 (N_3745,N_790,N_782);
and U3746 (N_3746,N_1617,N_1315);
and U3747 (N_3747,N_2530,N_1999);
nand U3748 (N_3748,N_2401,N_1430);
xor U3749 (N_3749,N_2698,N_181);
and U3750 (N_3750,N_2199,N_370);
xnor U3751 (N_3751,N_2828,N_1530);
or U3752 (N_3752,N_182,N_207);
and U3753 (N_3753,N_106,N_816);
xor U3754 (N_3754,N_234,N_2222);
and U3755 (N_3755,N_1761,N_2601);
nor U3756 (N_3756,N_1232,N_1473);
nand U3757 (N_3757,N_694,N_1697);
and U3758 (N_3758,N_626,N_784);
xor U3759 (N_3759,N_1923,N_1850);
xor U3760 (N_3760,N_1428,N_2868);
or U3761 (N_3761,N_2784,N_2221);
or U3762 (N_3762,N_513,N_796);
nor U3763 (N_3763,N_1065,N_1523);
xor U3764 (N_3764,N_1822,N_411);
nand U3765 (N_3765,N_2006,N_2587);
nor U3766 (N_3766,N_571,N_2881);
xor U3767 (N_3767,N_161,N_583);
xnor U3768 (N_3768,N_2979,N_1916);
nand U3769 (N_3769,N_2756,N_1079);
or U3770 (N_3770,N_2064,N_314);
nor U3771 (N_3771,N_498,N_2468);
or U3772 (N_3772,N_2061,N_2994);
or U3773 (N_3773,N_2611,N_1289);
nand U3774 (N_3774,N_2425,N_783);
or U3775 (N_3775,N_223,N_1244);
nand U3776 (N_3776,N_460,N_2078);
xor U3777 (N_3777,N_1250,N_2522);
nand U3778 (N_3778,N_2129,N_2089);
or U3779 (N_3779,N_2549,N_1572);
nand U3780 (N_3780,N_321,N_1495);
xor U3781 (N_3781,N_2632,N_1855);
nor U3782 (N_3782,N_1967,N_2843);
or U3783 (N_3783,N_1498,N_2424);
or U3784 (N_3784,N_2570,N_1691);
nand U3785 (N_3785,N_1973,N_1733);
nand U3786 (N_3786,N_727,N_2112);
or U3787 (N_3787,N_1070,N_2722);
xor U3788 (N_3788,N_248,N_151);
nand U3789 (N_3789,N_2206,N_1025);
and U3790 (N_3790,N_1332,N_2338);
or U3791 (N_3791,N_1297,N_979);
nor U3792 (N_3792,N_392,N_1706);
nor U3793 (N_3793,N_2742,N_2125);
nand U3794 (N_3794,N_1225,N_1807);
or U3795 (N_3795,N_2397,N_353);
nor U3796 (N_3796,N_1746,N_1827);
or U3797 (N_3797,N_2585,N_2002);
nor U3798 (N_3798,N_525,N_1673);
nor U3799 (N_3799,N_573,N_1290);
xnor U3800 (N_3800,N_2134,N_776);
or U3801 (N_3801,N_2677,N_1491);
nor U3802 (N_3802,N_1133,N_74);
nand U3803 (N_3803,N_2594,N_1738);
nand U3804 (N_3804,N_1760,N_2732);
nor U3805 (N_3805,N_1682,N_364);
and U3806 (N_3806,N_1396,N_422);
or U3807 (N_3807,N_1045,N_1568);
or U3808 (N_3808,N_1424,N_2336);
or U3809 (N_3809,N_1144,N_317);
and U3810 (N_3810,N_137,N_690);
xnor U3811 (N_3811,N_1857,N_574);
nor U3812 (N_3812,N_1853,N_324);
nor U3813 (N_3813,N_2974,N_891);
and U3814 (N_3814,N_1729,N_379);
or U3815 (N_3815,N_2514,N_1901);
nand U3816 (N_3816,N_1759,N_2313);
nand U3817 (N_3817,N_1519,N_2563);
nor U3818 (N_3818,N_305,N_2996);
or U3819 (N_3819,N_1358,N_2193);
or U3820 (N_3820,N_2813,N_2680);
and U3821 (N_3821,N_2864,N_275);
nor U3822 (N_3822,N_239,N_107);
xor U3823 (N_3823,N_1088,N_731);
nor U3824 (N_3824,N_1600,N_982);
or U3825 (N_3825,N_454,N_343);
or U3826 (N_3826,N_1376,N_2158);
xor U3827 (N_3827,N_2342,N_553);
nor U3828 (N_3828,N_527,N_385);
nand U3829 (N_3829,N_2952,N_1659);
xor U3830 (N_3830,N_1602,N_180);
nor U3831 (N_3831,N_115,N_38);
and U3832 (N_3832,N_206,N_2185);
nand U3833 (N_3833,N_2007,N_2067);
or U3834 (N_3834,N_1549,N_1068);
or U3835 (N_3835,N_1186,N_2173);
and U3836 (N_3836,N_2171,N_2237);
or U3837 (N_3837,N_2356,N_2501);
nand U3838 (N_3838,N_1711,N_1770);
nand U3839 (N_3839,N_1944,N_2111);
nand U3840 (N_3840,N_2785,N_789);
nand U3841 (N_3841,N_1120,N_355);
and U3842 (N_3842,N_2344,N_740);
or U3843 (N_3843,N_1393,N_1928);
xor U3844 (N_3844,N_86,N_1402);
nor U3845 (N_3845,N_1975,N_27);
and U3846 (N_3846,N_2435,N_2986);
or U3847 (N_3847,N_1146,N_8);
nor U3848 (N_3848,N_365,N_2040);
or U3849 (N_3849,N_76,N_1116);
nand U3850 (N_3850,N_1208,N_125);
or U3851 (N_3851,N_947,N_2097);
nor U3852 (N_3852,N_847,N_2293);
and U3853 (N_3853,N_2419,N_1985);
nor U3854 (N_3854,N_2230,N_2835);
or U3855 (N_3855,N_2500,N_102);
nor U3856 (N_3856,N_779,N_1751);
xnor U3857 (N_3857,N_2770,N_2056);
xnor U3858 (N_3858,N_186,N_1607);
or U3859 (N_3859,N_96,N_2092);
xor U3860 (N_3860,N_1227,N_554);
xor U3861 (N_3861,N_597,N_935);
or U3862 (N_3862,N_1429,N_88);
and U3863 (N_3863,N_1558,N_1461);
xnor U3864 (N_3864,N_2803,N_2590);
xnor U3865 (N_3865,N_2487,N_337);
or U3866 (N_3866,N_1668,N_2182);
nor U3867 (N_3867,N_1514,N_866);
nand U3868 (N_3868,N_844,N_995);
or U3869 (N_3869,N_1713,N_2658);
and U3870 (N_3870,N_2236,N_2801);
or U3871 (N_3871,N_1769,N_1125);
or U3872 (N_3872,N_1500,N_814);
xnor U3873 (N_3873,N_1762,N_933);
nor U3874 (N_3874,N_209,N_381);
nor U3875 (N_3875,N_512,N_1778);
nand U3876 (N_3876,N_1418,N_61);
and U3877 (N_3877,N_778,N_2852);
and U3878 (N_3878,N_332,N_1595);
or U3879 (N_3879,N_173,N_2845);
nand U3880 (N_3880,N_383,N_1331);
or U3881 (N_3881,N_284,N_2450);
nand U3882 (N_3882,N_701,N_2452);
xor U3883 (N_3883,N_673,N_356);
xnor U3884 (N_3884,N_226,N_841);
nor U3885 (N_3885,N_418,N_1681);
nand U3886 (N_3886,N_1546,N_2180);
or U3887 (N_3887,N_1910,N_1148);
nand U3888 (N_3888,N_1044,N_350);
xnor U3889 (N_3889,N_2159,N_976);
or U3890 (N_3890,N_1082,N_2650);
nand U3891 (N_3891,N_2350,N_1404);
nand U3892 (N_3892,N_195,N_596);
xor U3893 (N_3893,N_1907,N_1094);
nor U3894 (N_3894,N_292,N_1344);
nand U3895 (N_3895,N_2020,N_2377);
and U3896 (N_3896,N_2457,N_1011);
or U3897 (N_3897,N_502,N_2225);
xnor U3898 (N_3898,N_1633,N_190);
and U3899 (N_3899,N_16,N_2804);
nor U3900 (N_3900,N_1420,N_1380);
nor U3901 (N_3901,N_2807,N_522);
nand U3902 (N_3902,N_2647,N_2380);
and U3903 (N_3903,N_566,N_2147);
xnor U3904 (N_3904,N_2274,N_1958);
and U3905 (N_3905,N_1411,N_1040);
xor U3906 (N_3906,N_1362,N_437);
nand U3907 (N_3907,N_2145,N_1684);
xor U3908 (N_3908,N_1142,N_1567);
nand U3909 (N_3909,N_1666,N_1883);
and U3910 (N_3910,N_1368,N_1016);
or U3911 (N_3911,N_679,N_1672);
nand U3912 (N_3912,N_1627,N_2207);
or U3913 (N_3913,N_426,N_2266);
or U3914 (N_3914,N_551,N_2713);
nand U3915 (N_3915,N_20,N_2217);
xnor U3916 (N_3916,N_443,N_2568);
and U3917 (N_3917,N_829,N_257);
nand U3918 (N_3918,N_342,N_598);
or U3919 (N_3919,N_2524,N_2991);
and U3920 (N_3920,N_1915,N_2246);
and U3921 (N_3921,N_2211,N_1798);
nand U3922 (N_3922,N_919,N_2208);
xor U3923 (N_3923,N_2936,N_2555);
or U3924 (N_3924,N_14,N_2598);
or U3925 (N_3925,N_1829,N_348);
nor U3926 (N_3926,N_416,N_135);
and U3927 (N_3927,N_975,N_2407);
xnor U3928 (N_3928,N_146,N_37);
nor U3929 (N_3929,N_1145,N_262);
nand U3930 (N_3930,N_1784,N_974);
xor U3931 (N_3931,N_2608,N_2188);
nor U3932 (N_3932,N_526,N_415);
nor U3933 (N_3933,N_2229,N_1773);
and U3934 (N_3934,N_1335,N_494);
nand U3935 (N_3935,N_1198,N_1835);
and U3936 (N_3936,N_2662,N_1102);
nor U3937 (N_3937,N_2562,N_2046);
nand U3938 (N_3938,N_906,N_859);
nor U3939 (N_3939,N_794,N_1961);
xnor U3940 (N_3940,N_1842,N_2085);
nor U3941 (N_3941,N_1279,N_2169);
or U3942 (N_3942,N_1308,N_2822);
or U3943 (N_3943,N_493,N_2390);
or U3944 (N_3944,N_174,N_283);
and U3945 (N_3945,N_2602,N_1441);
nand U3946 (N_3946,N_1823,N_1442);
nor U3947 (N_3947,N_51,N_1590);
nor U3948 (N_3948,N_1547,N_1336);
xor U3949 (N_3949,N_1384,N_2983);
nor U3950 (N_3950,N_2977,N_650);
nand U3951 (N_3951,N_966,N_1222);
and U3952 (N_3952,N_2353,N_2918);
xor U3953 (N_3953,N_1351,N_1578);
nand U3954 (N_3954,N_264,N_1532);
or U3955 (N_3955,N_1270,N_1752);
nand U3956 (N_3956,N_2122,N_2957);
nand U3957 (N_3957,N_738,N_2718);
nand U3958 (N_3958,N_951,N_2669);
nor U3959 (N_3959,N_1041,N_2151);
nor U3960 (N_3960,N_2920,N_839);
nor U3961 (N_3961,N_1147,N_1211);
or U3962 (N_3962,N_328,N_375);
nand U3963 (N_3963,N_925,N_1623);
nor U3964 (N_3964,N_2943,N_245);
and U3965 (N_3965,N_677,N_1000);
or U3966 (N_3966,N_2474,N_2463);
nor U3967 (N_3967,N_183,N_1986);
nor U3968 (N_3968,N_1540,N_367);
or U3969 (N_3969,N_858,N_1964);
nand U3970 (N_3970,N_1093,N_1480);
xor U3971 (N_3971,N_801,N_1143);
or U3972 (N_3972,N_655,N_1373);
or U3973 (N_3973,N_709,N_497);
nor U3974 (N_3974,N_2084,N_1343);
and U3975 (N_3975,N_837,N_1067);
xnor U3976 (N_3976,N_1880,N_199);
and U3977 (N_3977,N_2252,N_2471);
nor U3978 (N_3978,N_2885,N_1528);
nand U3979 (N_3979,N_2036,N_1662);
xnor U3980 (N_3980,N_1875,N_2139);
xor U3981 (N_3981,N_1408,N_1510);
nor U3982 (N_3982,N_2298,N_138);
xor U3983 (N_3983,N_2666,N_828);
nor U3984 (N_3984,N_795,N_1663);
nand U3985 (N_3985,N_2455,N_920);
xnor U3986 (N_3986,N_114,N_2250);
nand U3987 (N_3987,N_2439,N_2511);
nand U3988 (N_3988,N_491,N_2128);
and U3989 (N_3989,N_179,N_723);
xor U3990 (N_3990,N_567,N_1575);
and U3991 (N_3991,N_448,N_1286);
and U3992 (N_3992,N_1353,N_1830);
xor U3993 (N_3993,N_439,N_1240);
xnor U3994 (N_3994,N_2363,N_2558);
xnor U3995 (N_3995,N_2528,N_1409);
and U3996 (N_3996,N_821,N_860);
and U3997 (N_3997,N_2,N_2053);
and U3998 (N_3998,N_2947,N_631);
xor U3999 (N_3999,N_2478,N_728);
nand U4000 (N_4000,N_2958,N_242);
nand U4001 (N_4001,N_309,N_594);
xnor U4002 (N_4002,N_1029,N_589);
xor U4003 (N_4003,N_781,N_1394);
or U4004 (N_4004,N_1245,N_1443);
and U4005 (N_4005,N_500,N_1168);
nand U4006 (N_4006,N_2812,N_84);
nor U4007 (N_4007,N_813,N_1630);
nor U4008 (N_4008,N_2797,N_1412);
xnor U4009 (N_4009,N_1283,N_466);
nor U4010 (N_4010,N_59,N_846);
nand U4011 (N_4011,N_259,N_2110);
xnor U4012 (N_4012,N_1990,N_2480);
and U4013 (N_4013,N_2913,N_698);
or U4014 (N_4014,N_587,N_244);
xor U4015 (N_4015,N_676,N_1139);
nor U4016 (N_4016,N_2746,N_901);
or U4017 (N_4017,N_2869,N_2385);
xnor U4018 (N_4018,N_2381,N_148);
or U4019 (N_4019,N_1372,N_922);
xnor U4020 (N_4020,N_2327,N_823);
nand U4021 (N_4021,N_2932,N_2280);
nand U4022 (N_4022,N_743,N_2600);
and U4023 (N_4023,N_395,N_1253);
xnor U4024 (N_4024,N_2304,N_397);
nand U4025 (N_4025,N_1255,N_624);
xor U4026 (N_4026,N_1058,N_1995);
xor U4027 (N_4027,N_609,N_2403);
nor U4028 (N_4028,N_2840,N_1313);
xor U4029 (N_4029,N_1754,N_531);
or U4030 (N_4030,N_969,N_436);
xnor U4031 (N_4031,N_373,N_1249);
and U4032 (N_4032,N_2396,N_1766);
nor U4033 (N_4033,N_85,N_1946);
nand U4034 (N_4034,N_868,N_1636);
nand U4035 (N_4035,N_2648,N_303);
nor U4036 (N_4036,N_1023,N_1030);
xnor U4037 (N_4037,N_1583,N_2703);
nand U4038 (N_4038,N_1022,N_2025);
and U4039 (N_4039,N_12,N_644);
nor U4040 (N_4040,N_1800,N_616);
nor U4041 (N_4041,N_2743,N_1176);
nand U4042 (N_4042,N_1867,N_1943);
or U4043 (N_4043,N_848,N_528);
or U4044 (N_4044,N_431,N_2661);
xor U4045 (N_4045,N_2453,N_854);
xnor U4046 (N_4046,N_1972,N_1878);
nand U4047 (N_4047,N_1814,N_193);
and U4048 (N_4048,N_1056,N_2930);
nor U4049 (N_4049,N_35,N_1260);
nand U4050 (N_4050,N_1643,N_2780);
xnor U4051 (N_4051,N_351,N_79);
or U4052 (N_4052,N_2433,N_1811);
nand U4053 (N_4053,N_1254,N_1501);
nand U4054 (N_4054,N_2512,N_2580);
nor U4055 (N_4055,N_1989,N_818);
nand U4056 (N_4056,N_2684,N_451);
xnor U4057 (N_4057,N_713,N_570);
or U4058 (N_4058,N_1456,N_2255);
xnor U4059 (N_4059,N_564,N_1184);
nand U4060 (N_4060,N_171,N_1311);
nor U4061 (N_4061,N_1185,N_2628);
and U4062 (N_4062,N_1433,N_2557);
or U4063 (N_4063,N_2805,N_2491);
nand U4064 (N_4064,N_7,N_1340);
xor U4065 (N_4065,N_977,N_2446);
nor U4066 (N_4066,N_2115,N_1739);
or U4067 (N_4067,N_2191,N_1209);
nand U4068 (N_4068,N_1718,N_1700);
nor U4069 (N_4069,N_1839,N_2260);
nand U4070 (N_4070,N_2755,N_2244);
xor U4071 (N_4071,N_273,N_158);
xnor U4072 (N_4072,N_2066,N_568);
and U4073 (N_4073,N_1020,N_2793);
xor U4074 (N_4074,N_878,N_2024);
nor U4075 (N_4075,N_2393,N_2098);
xor U4076 (N_4076,N_652,N_1033);
and U4077 (N_4077,N_2181,N_2720);
and U4078 (N_4078,N_1152,N_2538);
or U4079 (N_4079,N_592,N_477);
nand U4080 (N_4080,N_384,N_2646);
xnor U4081 (N_4081,N_1085,N_1610);
nand U4082 (N_4082,N_1652,N_621);
or U4083 (N_4083,N_2970,N_2186);
or U4084 (N_4084,N_1382,N_1091);
xnor U4085 (N_4085,N_576,N_544);
or U4086 (N_4086,N_2035,N_2806);
xnor U4087 (N_4087,N_1371,N_1267);
and U4088 (N_4088,N_2999,N_2361);
nor U4089 (N_4089,N_988,N_825);
nand U4090 (N_4090,N_1421,N_530);
and U4091 (N_4091,N_1472,N_1027);
xor U4092 (N_4092,N_2370,N_2796);
nor U4093 (N_4093,N_2016,N_1375);
xor U4094 (N_4094,N_55,N_219);
and U4095 (N_4095,N_2614,N_759);
xnor U4096 (N_4096,N_1688,N_1806);
nor U4097 (N_4097,N_667,N_838);
xor U4098 (N_4098,N_2062,N_1780);
nor U4099 (N_4099,N_2359,N_2966);
nor U4100 (N_4100,N_595,N_871);
or U4101 (N_4101,N_2203,N_1173);
or U4102 (N_4102,N_2683,N_2149);
and U4103 (N_4103,N_1484,N_465);
xnor U4104 (N_4104,N_1123,N_2242);
and U4105 (N_4105,N_879,N_447);
xor U4106 (N_4106,N_2009,N_152);
nor U4107 (N_4107,N_1543,N_2265);
or U4108 (N_4108,N_2705,N_1440);
nor U4109 (N_4109,N_1843,N_1248);
nand U4110 (N_4110,N_1001,N_2863);
or U4111 (N_4111,N_604,N_201);
nand U4112 (N_4112,N_1620,N_1644);
or U4113 (N_4113,N_1341,N_2167);
nor U4114 (N_4114,N_929,N_1141);
and U4115 (N_4115,N_23,N_400);
nor U4116 (N_4116,N_2581,N_2392);
and U4117 (N_4117,N_2582,N_555);
nand U4118 (N_4118,N_2834,N_1246);
and U4119 (N_4119,N_1921,N_1576);
nor U4120 (N_4120,N_549,N_2226);
or U4121 (N_4121,N_80,N_1864);
nor U4122 (N_4122,N_2814,N_798);
xnor U4123 (N_4123,N_429,N_1054);
nand U4124 (N_4124,N_1581,N_2441);
xor U4125 (N_4125,N_2509,N_1860);
xnor U4126 (N_4126,N_719,N_1488);
and U4127 (N_4127,N_149,N_2915);
nor U4128 (N_4128,N_453,N_432);
xor U4129 (N_4129,N_1629,N_2028);
nand U4130 (N_4130,N_2788,N_67);
nand U4131 (N_4131,N_1074,N_1314);
and U4132 (N_4132,N_217,N_2017);
or U4133 (N_4133,N_1525,N_2484);
or U4134 (N_4134,N_1175,N_1190);
and U4135 (N_4135,N_435,N_660);
and U4136 (N_4136,N_2862,N_2454);
nor U4137 (N_4137,N_496,N_505);
xnor U4138 (N_4138,N_2775,N_800);
nand U4139 (N_4139,N_2075,N_1195);
nor U4140 (N_4140,N_985,N_1904);
nand U4141 (N_4141,N_672,N_706);
xor U4142 (N_4142,N_1996,N_2000);
nand U4143 (N_4143,N_2604,N_2289);
nand U4144 (N_4144,N_1847,N_75);
and U4145 (N_4145,N_103,N_269);
and U4146 (N_4146,N_507,N_2752);
nor U4147 (N_4147,N_869,N_3);
nor U4148 (N_4148,N_2712,N_9);
or U4149 (N_4149,N_1899,N_1551);
xnor U4150 (N_4150,N_2496,N_26);
xnor U4151 (N_4151,N_128,N_2106);
nor U4152 (N_4152,N_2559,N_1243);
nand U4153 (N_4153,N_263,N_2665);
nand U4154 (N_4154,N_902,N_1670);
or U4155 (N_4155,N_178,N_1748);
or U4156 (N_4156,N_2113,N_1885);
nand U4157 (N_4157,N_2641,N_2275);
nand U4158 (N_4158,N_637,N_268);
nor U4159 (N_4159,N_2093,N_377);
or U4160 (N_4160,N_857,N_2574);
nor U4161 (N_4161,N_1300,N_1348);
or U4162 (N_4162,N_1171,N_765);
xnor U4163 (N_4163,N_2706,N_2504);
or U4164 (N_4164,N_1422,N_559);
xnor U4165 (N_4165,N_2469,N_1816);
xnor U4166 (N_4166,N_2711,N_2933);
nor U4167 (N_4167,N_689,N_2373);
and U4168 (N_4168,N_2284,N_2903);
nand U4169 (N_4169,N_1695,N_1007);
nor U4170 (N_4170,N_1437,N_32);
and U4171 (N_4171,N_1675,N_1457);
xor U4172 (N_4172,N_1038,N_1948);
nor U4173 (N_4173,N_2908,N_281);
xor U4174 (N_4174,N_153,N_2086);
nor U4175 (N_4175,N_408,N_2213);
xor U4176 (N_4176,N_484,N_1805);
xor U4177 (N_4177,N_64,N_433);
and U4178 (N_4178,N_1791,N_2757);
nor U4179 (N_4179,N_2395,N_802);
xor U4180 (N_4180,N_1268,N_1705);
xnor U4181 (N_4181,N_1599,N_508);
or U4182 (N_4182,N_1702,N_1911);
nor U4183 (N_4183,N_1821,N_452);
and U4184 (N_4184,N_2292,N_1230);
nor U4185 (N_4185,N_393,N_2777);
xor U4186 (N_4186,N_1641,N_1952);
and U4187 (N_4187,N_1561,N_143);
nand U4188 (N_4188,N_170,N_805);
and U4189 (N_4189,N_2907,N_211);
xor U4190 (N_4190,N_419,N_2005);
or U4191 (N_4191,N_202,N_2870);
and U4192 (N_4192,N_1608,N_1019);
nor U4193 (N_4193,N_1234,N_1856);
nand U4194 (N_4194,N_2691,N_2263);
xor U4195 (N_4195,N_389,N_808);
xnor U4196 (N_4196,N_1189,N_1615);
or U4197 (N_4197,N_1654,N_2257);
nand U4198 (N_4198,N_588,N_591);
nor U4199 (N_4199,N_1555,N_347);
nand U4200 (N_4200,N_1506,N_176);
nor U4201 (N_4201,N_725,N_2764);
or U4202 (N_4202,N_924,N_105);
or U4203 (N_4203,N_1893,N_1271);
or U4204 (N_4204,N_1527,N_1379);
and U4205 (N_4205,N_1942,N_2059);
nand U4206 (N_4206,N_702,N_90);
or U4207 (N_4207,N_1848,N_382);
nor U4208 (N_4208,N_968,N_2166);
xnor U4209 (N_4209,N_1401,N_2296);
nor U4210 (N_4210,N_1635,N_1149);
or U4211 (N_4211,N_1081,N_58);
or U4212 (N_4212,N_2649,N_1403);
and U4213 (N_4213,N_2754,N_184);
nand U4214 (N_4214,N_127,N_70);
and U4215 (N_4215,N_1192,N_767);
xnor U4216 (N_4216,N_2196,N_2398);
and U4217 (N_4217,N_2820,N_2786);
nand U4218 (N_4218,N_581,N_732);
and U4219 (N_4219,N_2928,N_1014);
nand U4220 (N_4220,N_897,N_215);
or U4221 (N_4221,N_2894,N_1231);
and U4222 (N_4222,N_1955,N_1035);
nand U4223 (N_4223,N_2654,N_198);
or U4224 (N_4224,N_1477,N_282);
nand U4225 (N_4225,N_2104,N_2519);
and U4226 (N_4226,N_2346,N_1406);
nor U4227 (N_4227,N_2671,N_361);
nor U4228 (N_4228,N_758,N_1119);
and U4229 (N_4229,N_2057,N_2287);
nor U4230 (N_4230,N_2969,N_627);
or U4231 (N_4231,N_1900,N_1968);
nor U4232 (N_4232,N_2753,N_2609);
nand U4233 (N_4233,N_2027,N_887);
nor U4234 (N_4234,N_1405,N_2836);
nand U4235 (N_4235,N_2464,N_1266);
nor U4236 (N_4236,N_520,N_532);
nor U4237 (N_4237,N_1039,N_191);
nand U4238 (N_4238,N_1556,N_39);
xor U4239 (N_4239,N_1585,N_651);
or U4240 (N_4240,N_1920,N_2929);
nor U4241 (N_4241,N_2189,N_733);
or U4242 (N_4242,N_744,N_2924);
or U4243 (N_4243,N_2096,N_1965);
or U4244 (N_4244,N_914,N_1156);
or U4245 (N_4245,N_1974,N_2973);
xnor U4246 (N_4246,N_2490,N_649);
and U4247 (N_4247,N_1657,N_256);
nand U4248 (N_4248,N_916,N_992);
nand U4249 (N_4249,N_1622,N_2492);
nand U4250 (N_4250,N_2023,N_2651);
nand U4251 (N_4251,N_2873,N_2523);
nand U4252 (N_4252,N_2747,N_680);
nand U4253 (N_4253,N_2525,N_2328);
nand U4254 (N_4254,N_2527,N_1997);
and U4255 (N_4255,N_212,N_514);
nor U4256 (N_4256,N_2321,N_2619);
or U4257 (N_4257,N_717,N_1272);
nor U4258 (N_4258,N_2642,N_2748);
nand U4259 (N_4259,N_116,N_580);
xor U4260 (N_4260,N_1312,N_1689);
xnor U4261 (N_4261,N_1824,N_2636);
xor U4262 (N_4262,N_2426,N_760);
xor U4263 (N_4263,N_2763,N_950);
xnor U4264 (N_4264,N_2271,N_716);
nor U4265 (N_4265,N_1808,N_1988);
nor U4266 (N_4266,N_1819,N_1802);
nand U4267 (N_4267,N_873,N_1481);
and U4268 (N_4268,N_1647,N_684);
nand U4269 (N_4269,N_402,N_1448);
xor U4270 (N_4270,N_2547,N_809);
nor U4271 (N_4271,N_1241,N_2227);
nand U4272 (N_4272,N_164,N_2485);
nand U4273 (N_4273,N_2408,N_277);
nand U4274 (N_4274,N_2882,N_2700);
nor U4275 (N_4275,N_154,N_1865);
xnor U4276 (N_4276,N_1708,N_1258);
xor U4277 (N_4277,N_700,N_2329);
nor U4278 (N_4278,N_113,N_1539);
nor U4279 (N_4279,N_2798,N_2010);
and U4280 (N_4280,N_2347,N_2473);
or U4281 (N_4281,N_1365,N_2309);
xor U4282 (N_4282,N_1309,N_46);
nand U4283 (N_4283,N_2270,N_927);
and U4284 (N_4284,N_820,N_1884);
nor U4285 (N_4285,N_2156,N_1797);
xor U4286 (N_4286,N_455,N_66);
or U4287 (N_4287,N_300,N_1887);
nor U4288 (N_4288,N_2789,N_1112);
and U4289 (N_4289,N_1167,N_1591);
xor U4290 (N_4290,N_2216,N_1072);
and U4291 (N_4291,N_1419,N_585);
nor U4292 (N_4292,N_1210,N_1299);
nor U4293 (N_4293,N_1449,N_606);
nor U4294 (N_4294,N_489,N_1334);
or U4295 (N_4295,N_78,N_1439);
xnor U4296 (N_4296,N_1096,N_2285);
nor U4297 (N_4297,N_2283,N_2846);
nand U4298 (N_4298,N_2909,N_2517);
or U4299 (N_4299,N_485,N_2297);
nand U4300 (N_4300,N_2926,N_2702);
nand U4301 (N_4301,N_946,N_1318);
nor U4302 (N_4302,N_1342,N_1792);
or U4303 (N_4303,N_851,N_2432);
and U4304 (N_4304,N_2980,N_2153);
nand U4305 (N_4305,N_710,N_1193);
or U4306 (N_4306,N_2853,N_1592);
xnor U4307 (N_4307,N_1586,N_970);
xnor U4308 (N_4308,N_1159,N_663);
xor U4309 (N_4309,N_1728,N_917);
and U4310 (N_4310,N_2588,N_2610);
nand U4311 (N_4311,N_2011,N_1316);
nor U4312 (N_4312,N_964,N_619);
or U4313 (N_4313,N_2412,N_853);
nand U4314 (N_4314,N_1224,N_683);
or U4315 (N_4315,N_2731,N_2938);
nand U4316 (N_4316,N_120,N_1606);
or U4317 (N_4317,N_2386,N_645);
xor U4318 (N_4318,N_2123,N_2114);
nor U4319 (N_4319,N_1852,N_611);
xor U4320 (N_4320,N_293,N_915);
or U4321 (N_4321,N_894,N_1871);
or U4322 (N_4322,N_296,N_1957);
or U4323 (N_4323,N_417,N_2319);
or U4324 (N_4324,N_1239,N_1574);
nand U4325 (N_4325,N_1363,N_1028);
and U4326 (N_4326,N_2827,N_194);
nand U4327 (N_4327,N_1560,N_2548);
and U4328 (N_4328,N_1257,N_1660);
or U4329 (N_4329,N_2726,N_1508);
and U4330 (N_4330,N_2176,N_2976);
nand U4331 (N_4331,N_1138,N_2513);
nand U4332 (N_4332,N_1742,N_394);
and U4333 (N_4333,N_1922,N_1095);
or U4334 (N_4334,N_1725,N_2686);
and U4335 (N_4335,N_533,N_189);
nand U4336 (N_4336,N_641,N_136);
or U4337 (N_4337,N_2967,N_1359);
or U4338 (N_4338,N_1756,N_2871);
nand U4339 (N_4339,N_2146,N_1648);
or U4340 (N_4340,N_2567,N_1927);
or U4341 (N_4341,N_1937,N_1356);
and U4342 (N_4342,N_2687,N_2685);
xnor U4343 (N_4343,N_83,N_843);
xnor U4344 (N_4344,N_1470,N_139);
and U4345 (N_4345,N_2701,N_1086);
xnor U4346 (N_4346,N_1544,N_372);
nand U4347 (N_4347,N_1238,N_2341);
nand U4348 (N_4348,N_98,N_1625);
xor U4349 (N_4349,N_913,N_884);
and U4350 (N_4350,N_2320,N_2048);
and U4351 (N_4351,N_1534,N_2638);
or U4352 (N_4352,N_2579,N_2019);
xor U4353 (N_4353,N_376,N_788);
or U4354 (N_4354,N_1031,N_2616);
nor U4355 (N_4355,N_552,N_2693);
and U4356 (N_4356,N_605,N_475);
nand U4357 (N_4357,N_2771,N_2893);
xor U4358 (N_4358,N_2633,N_1735);
nor U4359 (N_4359,N_1597,N_1951);
nor U4360 (N_4360,N_22,N_221);
xnor U4361 (N_4361,N_707,N_330);
nand U4362 (N_4362,N_622,N_1427);
xnor U4363 (N_4363,N_2269,N_1483);
nand U4364 (N_4364,N_2995,N_2415);
xor U4365 (N_4365,N_1069,N_1064);
nand U4366 (N_4366,N_693,N_899);
nor U4367 (N_4367,N_2850,N_1929);
nor U4368 (N_4368,N_1749,N_1801);
xor U4369 (N_4369,N_391,N_482);
nor U4370 (N_4370,N_2603,N_1153);
xor U4371 (N_4371,N_516,N_1170);
xor U4372 (N_4372,N_2531,N_1535);
and U4373 (N_4373,N_575,N_737);
and U4374 (N_4374,N_1858,N_162);
xnor U4375 (N_4375,N_1262,N_463);
nand U4376 (N_4376,N_387,N_94);
and U4377 (N_4377,N_2254,N_2904);
and U4378 (N_4378,N_1833,N_2223);
nor U4379 (N_4379,N_2368,N_2655);
and U4380 (N_4380,N_2015,N_607);
and U4381 (N_4381,N_1494,N_653);
nand U4382 (N_4382,N_2055,N_1649);
xor U4383 (N_4383,N_2571,N_1165);
and U4384 (N_4384,N_547,N_2656);
nand U4385 (N_4385,N_2699,N_2573);
and U4386 (N_4386,N_670,N_2444);
nor U4387 (N_4387,N_2261,N_33);
and U4388 (N_4388,N_1264,N_2817);
xor U4389 (N_4389,N_1485,N_266);
xnor U4390 (N_4390,N_686,N_2674);
nand U4391 (N_4391,N_265,N_2264);
or U4392 (N_4392,N_232,N_1699);
or U4393 (N_4393,N_1310,N_1122);
xor U4394 (N_4394,N_2447,N_509);
xnor U4395 (N_4395,N_2306,N_2719);
xnor U4396 (N_4396,N_2749,N_1010);
and U4397 (N_4397,N_2163,N_865);
nand U4398 (N_4398,N_2689,N_288);
or U4399 (N_4399,N_1388,N_1658);
nor U4400 (N_4400,N_45,N_490);
or U4401 (N_4401,N_519,N_1642);
xor U4402 (N_4402,N_1217,N_1669);
or U4403 (N_4403,N_1775,N_2340);
nor U4404 (N_4404,N_54,N_420);
and U4405 (N_4405,N_943,N_2906);
and U4406 (N_4406,N_228,N_2861);
nor U4407 (N_4407,N_2360,N_386);
xnor U4408 (N_4408,N_2740,N_1129);
nand U4409 (N_4409,N_122,N_926);
xnor U4410 (N_4410,N_762,N_1524);
and U4411 (N_4411,N_2256,N_1460);
nand U4412 (N_4412,N_468,N_648);
and U4413 (N_4413,N_1432,N_896);
xnor U4414 (N_4414,N_1325,N_511);
or U4415 (N_4415,N_1787,N_1577);
nand U4416 (N_4416,N_457,N_1804);
nand U4417 (N_4417,N_1796,N_1781);
and U4418 (N_4418,N_2470,N_2741);
nand U4419 (N_4419,N_1541,N_1140);
and U4420 (N_4420,N_1347,N_1087);
nand U4421 (N_4421,N_1169,N_1459);
nand U4422 (N_4422,N_2422,N_2160);
nand U4423 (N_4423,N_2443,N_2121);
xnor U4424 (N_4424,N_2660,N_1117);
nor U4425 (N_4425,N_251,N_2507);
and U4426 (N_4426,N_2953,N_2483);
nor U4427 (N_4427,N_2021,N_52);
nand U4428 (N_4428,N_1263,N_1679);
nor U4429 (N_4429,N_2212,N_2898);
nor U4430 (N_4430,N_43,N_1237);
xor U4431 (N_4431,N_2896,N_366);
nand U4432 (N_4432,N_2302,N_362);
xnor U4433 (N_4433,N_231,N_1497);
and U4434 (N_4434,N_2486,N_1115);
or U4435 (N_4435,N_910,N_2082);
and U4436 (N_4436,N_1083,N_2572);
and U4437 (N_4437,N_2162,N_117);
or U4438 (N_4438,N_518,N_2136);
and U4439 (N_4439,N_875,N_459);
xnor U4440 (N_4440,N_1162,N_755);
or U4441 (N_4441,N_2409,N_2290);
nor U4442 (N_4442,N_1504,N_1355);
or U4443 (N_4443,N_2987,N_2440);
xor U4444 (N_4444,N_1828,N_1918);
and U4445 (N_4445,N_2874,N_1655);
or U4446 (N_4446,N_2461,N_2593);
nand U4447 (N_4447,N_1157,N_1296);
nor U4448 (N_4448,N_2623,N_1339);
or U4449 (N_4449,N_2922,N_2546);
and U4450 (N_4450,N_1078,N_1704);
nor U4451 (N_4451,N_1292,N_2172);
nor U4452 (N_4452,N_1287,N_1385);
and U4453 (N_4453,N_315,N_2679);
nor U4454 (N_4454,N_2228,N_2175);
nand U4455 (N_4455,N_409,N_2090);
xor U4456 (N_4456,N_1326,N_1446);
nand U4457 (N_4457,N_1520,N_2829);
nand U4458 (N_4458,N_752,N_2890);
xor U4459 (N_4459,N_31,N_2561);
and U4460 (N_4460,N_2744,N_1503);
or U4461 (N_4461,N_213,N_1071);
nor U4462 (N_4462,N_1012,N_480);
nand U4463 (N_4463,N_2238,N_1304);
and U4464 (N_4464,N_53,N_461);
nand U4465 (N_4465,N_1545,N_335);
or U4466 (N_4466,N_2841,N_1611);
nor U4467 (N_4467,N_1803,N_734);
nand U4468 (N_4468,N_2734,N_986);
xor U4469 (N_4469,N_1345,N_904);
nor U4470 (N_4470,N_687,N_889);
xor U4471 (N_4471,N_1683,N_2831);
or U4472 (N_4472,N_487,N_2707);
nor U4473 (N_4473,N_56,N_769);
nor U4474 (N_4474,N_2108,N_42);
or U4475 (N_4475,N_1174,N_13);
xnor U4476 (N_4476,N_1113,N_403);
nor U4477 (N_4477,N_1383,N_481);
nor U4478 (N_4478,N_2617,N_1118);
xnor U4479 (N_4479,N_791,N_1322);
and U4480 (N_4480,N_2047,N_1863);
or U4481 (N_4481,N_685,N_438);
nor U4482 (N_4482,N_81,N_1204);
nor U4483 (N_4483,N_2445,N_301);
nand U4484 (N_4484,N_615,N_2218);
nand U4485 (N_4485,N_2860,N_57);
or U4486 (N_4486,N_1399,N_1317);
nand U4487 (N_4487,N_1859,N_2897);
nor U4488 (N_4488,N_4,N_1872);
nor U4489 (N_4489,N_339,N_71);
xor U4490 (N_4490,N_2437,N_1135);
nand U4491 (N_4491,N_2155,N_2972);
and U4492 (N_4492,N_1624,N_2887);
and U4493 (N_4493,N_1526,N_1533);
and U4494 (N_4494,N_953,N_1721);
nor U4495 (N_4495,N_856,N_1077);
and U4496 (N_4496,N_1564,N_2842);
and U4497 (N_4497,N_340,N_405);
and U4498 (N_4498,N_104,N_1969);
nand U4499 (N_4499,N_2183,N_2879);
and U4500 (N_4500,N_2443,N_1847);
or U4501 (N_4501,N_2178,N_1450);
xor U4502 (N_4502,N_1999,N_2236);
nand U4503 (N_4503,N_1101,N_1755);
nand U4504 (N_4504,N_2358,N_2988);
xor U4505 (N_4505,N_768,N_1706);
and U4506 (N_4506,N_744,N_952);
or U4507 (N_4507,N_2305,N_2496);
or U4508 (N_4508,N_2438,N_1147);
nand U4509 (N_4509,N_553,N_2295);
xor U4510 (N_4510,N_1871,N_1546);
and U4511 (N_4511,N_1847,N_2238);
or U4512 (N_4512,N_809,N_2159);
and U4513 (N_4513,N_981,N_1919);
or U4514 (N_4514,N_152,N_605);
nor U4515 (N_4515,N_2754,N_551);
xor U4516 (N_4516,N_1563,N_218);
or U4517 (N_4517,N_1686,N_333);
and U4518 (N_4518,N_35,N_1823);
and U4519 (N_4519,N_2336,N_1699);
nor U4520 (N_4520,N_118,N_1049);
nand U4521 (N_4521,N_859,N_780);
or U4522 (N_4522,N_2447,N_1257);
nor U4523 (N_4523,N_1894,N_2707);
or U4524 (N_4524,N_2451,N_2953);
and U4525 (N_4525,N_2686,N_1829);
nand U4526 (N_4526,N_1702,N_1093);
xnor U4527 (N_4527,N_2819,N_974);
nand U4528 (N_4528,N_164,N_311);
nor U4529 (N_4529,N_1340,N_1050);
nand U4530 (N_4530,N_1032,N_2079);
and U4531 (N_4531,N_1742,N_886);
or U4532 (N_4532,N_2976,N_1448);
and U4533 (N_4533,N_782,N_1201);
and U4534 (N_4534,N_2652,N_2650);
or U4535 (N_4535,N_2637,N_1716);
nand U4536 (N_4536,N_653,N_1480);
nand U4537 (N_4537,N_197,N_1797);
or U4538 (N_4538,N_247,N_896);
nand U4539 (N_4539,N_452,N_210);
and U4540 (N_4540,N_1484,N_2878);
nand U4541 (N_4541,N_590,N_1928);
nor U4542 (N_4542,N_691,N_1631);
or U4543 (N_4543,N_1871,N_1285);
xor U4544 (N_4544,N_1070,N_2657);
or U4545 (N_4545,N_1912,N_2236);
and U4546 (N_4546,N_2736,N_1571);
or U4547 (N_4547,N_768,N_1800);
xor U4548 (N_4548,N_1385,N_1711);
and U4549 (N_4549,N_399,N_2833);
and U4550 (N_4550,N_1757,N_1819);
nand U4551 (N_4551,N_2813,N_2487);
xnor U4552 (N_4552,N_823,N_766);
xor U4553 (N_4553,N_860,N_2875);
nand U4554 (N_4554,N_273,N_2559);
xnor U4555 (N_4555,N_1166,N_2093);
or U4556 (N_4556,N_1184,N_2877);
nor U4557 (N_4557,N_2916,N_2069);
xor U4558 (N_4558,N_2937,N_1558);
xnor U4559 (N_4559,N_410,N_2649);
nor U4560 (N_4560,N_1458,N_904);
and U4561 (N_4561,N_250,N_1816);
and U4562 (N_4562,N_484,N_2095);
xnor U4563 (N_4563,N_650,N_1213);
and U4564 (N_4564,N_2682,N_1736);
or U4565 (N_4565,N_1449,N_301);
and U4566 (N_4566,N_2890,N_1411);
or U4567 (N_4567,N_1673,N_1886);
xnor U4568 (N_4568,N_2899,N_160);
or U4569 (N_4569,N_680,N_1597);
nor U4570 (N_4570,N_810,N_2198);
and U4571 (N_4571,N_1564,N_1267);
nor U4572 (N_4572,N_1312,N_1411);
xor U4573 (N_4573,N_1141,N_454);
and U4574 (N_4574,N_2815,N_1850);
nand U4575 (N_4575,N_2869,N_1470);
nand U4576 (N_4576,N_379,N_2311);
or U4577 (N_4577,N_1009,N_101);
xnor U4578 (N_4578,N_1575,N_1937);
and U4579 (N_4579,N_2317,N_1316);
nand U4580 (N_4580,N_1903,N_1642);
or U4581 (N_4581,N_1084,N_824);
nor U4582 (N_4582,N_2959,N_856);
nand U4583 (N_4583,N_2482,N_2094);
or U4584 (N_4584,N_424,N_2801);
nand U4585 (N_4585,N_2477,N_2872);
nor U4586 (N_4586,N_142,N_492);
and U4587 (N_4587,N_2367,N_963);
and U4588 (N_4588,N_2082,N_1560);
nor U4589 (N_4589,N_448,N_80);
nand U4590 (N_4590,N_510,N_1426);
xnor U4591 (N_4591,N_1879,N_2692);
xor U4592 (N_4592,N_142,N_1631);
nand U4593 (N_4593,N_2717,N_30);
or U4594 (N_4594,N_35,N_2189);
and U4595 (N_4595,N_723,N_2026);
or U4596 (N_4596,N_2067,N_1821);
or U4597 (N_4597,N_1006,N_2185);
or U4598 (N_4598,N_670,N_1193);
nor U4599 (N_4599,N_1414,N_605);
nand U4600 (N_4600,N_1950,N_2067);
nand U4601 (N_4601,N_1840,N_2417);
nor U4602 (N_4602,N_429,N_2819);
xor U4603 (N_4603,N_1999,N_2588);
or U4604 (N_4604,N_1774,N_897);
and U4605 (N_4605,N_1628,N_2349);
nor U4606 (N_4606,N_1442,N_1060);
nor U4607 (N_4607,N_2034,N_1310);
xnor U4608 (N_4608,N_1528,N_2169);
or U4609 (N_4609,N_1123,N_1599);
nor U4610 (N_4610,N_2686,N_1798);
xor U4611 (N_4611,N_1893,N_1607);
nand U4612 (N_4612,N_452,N_342);
nor U4613 (N_4613,N_368,N_997);
and U4614 (N_4614,N_2693,N_2035);
nor U4615 (N_4615,N_707,N_2759);
xnor U4616 (N_4616,N_794,N_1076);
or U4617 (N_4617,N_1896,N_1018);
and U4618 (N_4618,N_2339,N_2029);
and U4619 (N_4619,N_1669,N_1947);
nor U4620 (N_4620,N_169,N_441);
xor U4621 (N_4621,N_228,N_1732);
or U4622 (N_4622,N_2745,N_466);
and U4623 (N_4623,N_2236,N_1197);
nand U4624 (N_4624,N_2944,N_1367);
xnor U4625 (N_4625,N_1778,N_82);
nand U4626 (N_4626,N_2080,N_903);
nand U4627 (N_4627,N_1937,N_2841);
or U4628 (N_4628,N_2975,N_185);
nand U4629 (N_4629,N_1617,N_641);
or U4630 (N_4630,N_2661,N_1896);
nand U4631 (N_4631,N_2082,N_2294);
xnor U4632 (N_4632,N_1695,N_116);
nand U4633 (N_4633,N_2342,N_1899);
xor U4634 (N_4634,N_1577,N_2869);
and U4635 (N_4635,N_2745,N_534);
and U4636 (N_4636,N_1624,N_502);
nand U4637 (N_4637,N_902,N_2981);
nor U4638 (N_4638,N_309,N_442);
xnor U4639 (N_4639,N_899,N_1038);
nor U4640 (N_4640,N_123,N_2972);
nor U4641 (N_4641,N_2170,N_415);
xnor U4642 (N_4642,N_1565,N_2887);
nand U4643 (N_4643,N_2040,N_84);
nor U4644 (N_4644,N_2216,N_1620);
and U4645 (N_4645,N_1527,N_2407);
nand U4646 (N_4646,N_682,N_1318);
and U4647 (N_4647,N_1277,N_1687);
xnor U4648 (N_4648,N_786,N_2042);
or U4649 (N_4649,N_316,N_2223);
nand U4650 (N_4650,N_390,N_1344);
and U4651 (N_4651,N_1713,N_11);
or U4652 (N_4652,N_1867,N_1185);
nor U4653 (N_4653,N_1678,N_2000);
xor U4654 (N_4654,N_2429,N_1182);
xor U4655 (N_4655,N_1640,N_10);
nand U4656 (N_4656,N_2200,N_2873);
nand U4657 (N_4657,N_2766,N_192);
and U4658 (N_4658,N_2831,N_2280);
xor U4659 (N_4659,N_417,N_566);
xor U4660 (N_4660,N_1418,N_986);
and U4661 (N_4661,N_640,N_1632);
xnor U4662 (N_4662,N_1163,N_1134);
nand U4663 (N_4663,N_1032,N_1026);
xnor U4664 (N_4664,N_1192,N_1768);
and U4665 (N_4665,N_1806,N_517);
nand U4666 (N_4666,N_387,N_183);
xnor U4667 (N_4667,N_92,N_2747);
and U4668 (N_4668,N_1115,N_2363);
and U4669 (N_4669,N_1080,N_2740);
nand U4670 (N_4670,N_188,N_110);
xor U4671 (N_4671,N_2916,N_2030);
nor U4672 (N_4672,N_926,N_1391);
nor U4673 (N_4673,N_830,N_316);
nand U4674 (N_4674,N_2416,N_369);
or U4675 (N_4675,N_1098,N_94);
or U4676 (N_4676,N_577,N_2325);
nand U4677 (N_4677,N_2495,N_1398);
and U4678 (N_4678,N_131,N_691);
and U4679 (N_4679,N_581,N_2870);
and U4680 (N_4680,N_2808,N_682);
xnor U4681 (N_4681,N_1243,N_2664);
or U4682 (N_4682,N_440,N_1875);
nor U4683 (N_4683,N_2274,N_2003);
nand U4684 (N_4684,N_1650,N_365);
nand U4685 (N_4685,N_1706,N_2384);
xor U4686 (N_4686,N_1959,N_1349);
nor U4687 (N_4687,N_1866,N_2479);
and U4688 (N_4688,N_729,N_682);
nor U4689 (N_4689,N_745,N_2622);
xor U4690 (N_4690,N_2840,N_1139);
xnor U4691 (N_4691,N_2946,N_2351);
or U4692 (N_4692,N_2408,N_1634);
xor U4693 (N_4693,N_1571,N_519);
and U4694 (N_4694,N_2300,N_2268);
xnor U4695 (N_4695,N_2965,N_979);
xnor U4696 (N_4696,N_1479,N_2846);
or U4697 (N_4697,N_638,N_643);
and U4698 (N_4698,N_1754,N_1596);
xnor U4699 (N_4699,N_2577,N_2559);
xnor U4700 (N_4700,N_326,N_2921);
and U4701 (N_4701,N_1918,N_2400);
xor U4702 (N_4702,N_1267,N_1831);
nand U4703 (N_4703,N_821,N_160);
nor U4704 (N_4704,N_2903,N_2537);
xor U4705 (N_4705,N_1277,N_1249);
and U4706 (N_4706,N_2427,N_15);
nor U4707 (N_4707,N_1649,N_2143);
and U4708 (N_4708,N_1946,N_364);
or U4709 (N_4709,N_2301,N_609);
nand U4710 (N_4710,N_2452,N_1902);
and U4711 (N_4711,N_1104,N_2024);
and U4712 (N_4712,N_2254,N_1989);
nand U4713 (N_4713,N_1368,N_2464);
nor U4714 (N_4714,N_1196,N_2277);
and U4715 (N_4715,N_1960,N_2842);
or U4716 (N_4716,N_1998,N_2638);
and U4717 (N_4717,N_890,N_2278);
nand U4718 (N_4718,N_434,N_2083);
nand U4719 (N_4719,N_1229,N_1104);
nand U4720 (N_4720,N_2570,N_2175);
or U4721 (N_4721,N_1655,N_1944);
xnor U4722 (N_4722,N_764,N_1777);
and U4723 (N_4723,N_995,N_136);
and U4724 (N_4724,N_1940,N_782);
xor U4725 (N_4725,N_2783,N_24);
nand U4726 (N_4726,N_554,N_2686);
nand U4727 (N_4727,N_1690,N_2710);
and U4728 (N_4728,N_336,N_117);
xnor U4729 (N_4729,N_1812,N_1418);
nand U4730 (N_4730,N_896,N_2729);
and U4731 (N_4731,N_2262,N_1480);
nor U4732 (N_4732,N_2499,N_2857);
nand U4733 (N_4733,N_2674,N_762);
xor U4734 (N_4734,N_803,N_604);
or U4735 (N_4735,N_2850,N_2067);
nand U4736 (N_4736,N_1961,N_59);
nor U4737 (N_4737,N_2002,N_2402);
nor U4738 (N_4738,N_874,N_2522);
nand U4739 (N_4739,N_2091,N_1846);
xnor U4740 (N_4740,N_1802,N_2817);
or U4741 (N_4741,N_645,N_1848);
xor U4742 (N_4742,N_2599,N_2165);
or U4743 (N_4743,N_2955,N_194);
xnor U4744 (N_4744,N_2267,N_1528);
or U4745 (N_4745,N_1902,N_1702);
nor U4746 (N_4746,N_595,N_1540);
and U4747 (N_4747,N_1182,N_2912);
nor U4748 (N_4748,N_78,N_346);
nor U4749 (N_4749,N_2874,N_1026);
or U4750 (N_4750,N_2656,N_1051);
or U4751 (N_4751,N_2858,N_322);
and U4752 (N_4752,N_2269,N_2310);
xor U4753 (N_4753,N_387,N_831);
nand U4754 (N_4754,N_567,N_2836);
nor U4755 (N_4755,N_2728,N_2428);
and U4756 (N_4756,N_665,N_2314);
and U4757 (N_4757,N_927,N_1549);
nand U4758 (N_4758,N_2927,N_947);
nand U4759 (N_4759,N_2483,N_1786);
nor U4760 (N_4760,N_206,N_640);
and U4761 (N_4761,N_2312,N_2016);
nor U4762 (N_4762,N_1928,N_1808);
and U4763 (N_4763,N_2838,N_189);
xor U4764 (N_4764,N_1891,N_2628);
xor U4765 (N_4765,N_888,N_2393);
or U4766 (N_4766,N_2588,N_260);
nor U4767 (N_4767,N_1817,N_2874);
or U4768 (N_4768,N_690,N_284);
or U4769 (N_4769,N_497,N_1326);
nor U4770 (N_4770,N_2602,N_306);
or U4771 (N_4771,N_2024,N_2595);
and U4772 (N_4772,N_2977,N_2802);
xnor U4773 (N_4773,N_1192,N_1257);
xnor U4774 (N_4774,N_2183,N_542);
nand U4775 (N_4775,N_2603,N_1132);
or U4776 (N_4776,N_2588,N_2884);
or U4777 (N_4777,N_1040,N_321);
or U4778 (N_4778,N_1383,N_475);
nor U4779 (N_4779,N_2709,N_1407);
or U4780 (N_4780,N_1906,N_2115);
or U4781 (N_4781,N_2850,N_2018);
xnor U4782 (N_4782,N_1866,N_2095);
nor U4783 (N_4783,N_360,N_1081);
xnor U4784 (N_4784,N_2118,N_1449);
xnor U4785 (N_4785,N_1227,N_149);
xor U4786 (N_4786,N_2341,N_2510);
xor U4787 (N_4787,N_2885,N_1180);
nor U4788 (N_4788,N_1170,N_2596);
xor U4789 (N_4789,N_1892,N_1319);
or U4790 (N_4790,N_994,N_64);
nor U4791 (N_4791,N_2222,N_274);
and U4792 (N_4792,N_1911,N_2353);
nor U4793 (N_4793,N_2061,N_1329);
xnor U4794 (N_4794,N_220,N_2438);
and U4795 (N_4795,N_2047,N_1654);
nor U4796 (N_4796,N_1976,N_636);
or U4797 (N_4797,N_748,N_674);
nand U4798 (N_4798,N_2173,N_1755);
nand U4799 (N_4799,N_2132,N_2724);
and U4800 (N_4800,N_11,N_2501);
nor U4801 (N_4801,N_577,N_1496);
nor U4802 (N_4802,N_1965,N_1772);
nand U4803 (N_4803,N_639,N_2901);
xnor U4804 (N_4804,N_1244,N_2135);
nor U4805 (N_4805,N_1575,N_2589);
and U4806 (N_4806,N_1008,N_2444);
xor U4807 (N_4807,N_924,N_1647);
nor U4808 (N_4808,N_1087,N_2801);
or U4809 (N_4809,N_861,N_280);
nor U4810 (N_4810,N_1104,N_709);
and U4811 (N_4811,N_151,N_2094);
nand U4812 (N_4812,N_143,N_2060);
or U4813 (N_4813,N_1706,N_559);
or U4814 (N_4814,N_1642,N_2081);
xnor U4815 (N_4815,N_857,N_1146);
nor U4816 (N_4816,N_1904,N_1016);
xor U4817 (N_4817,N_71,N_2456);
xnor U4818 (N_4818,N_1102,N_1147);
xnor U4819 (N_4819,N_2176,N_60);
xor U4820 (N_4820,N_1734,N_2519);
nand U4821 (N_4821,N_2334,N_1052);
xnor U4822 (N_4822,N_763,N_327);
nor U4823 (N_4823,N_1408,N_2474);
nand U4824 (N_4824,N_1538,N_2436);
xor U4825 (N_4825,N_257,N_2861);
xor U4826 (N_4826,N_2715,N_2960);
nand U4827 (N_4827,N_1390,N_2189);
xnor U4828 (N_4828,N_2546,N_442);
nor U4829 (N_4829,N_537,N_1757);
and U4830 (N_4830,N_2363,N_2209);
and U4831 (N_4831,N_2104,N_1665);
nor U4832 (N_4832,N_2760,N_1911);
xnor U4833 (N_4833,N_2116,N_2986);
nor U4834 (N_4834,N_866,N_958);
or U4835 (N_4835,N_2883,N_2416);
and U4836 (N_4836,N_425,N_1179);
nand U4837 (N_4837,N_2430,N_2981);
nand U4838 (N_4838,N_2855,N_2965);
nand U4839 (N_4839,N_1227,N_2232);
nor U4840 (N_4840,N_2371,N_426);
xor U4841 (N_4841,N_2305,N_2379);
xor U4842 (N_4842,N_2228,N_2433);
nand U4843 (N_4843,N_268,N_425);
and U4844 (N_4844,N_258,N_2735);
xnor U4845 (N_4845,N_211,N_2477);
xnor U4846 (N_4846,N_2191,N_1044);
and U4847 (N_4847,N_438,N_1798);
and U4848 (N_4848,N_717,N_1082);
nand U4849 (N_4849,N_489,N_2984);
and U4850 (N_4850,N_1646,N_2951);
nand U4851 (N_4851,N_1177,N_1376);
and U4852 (N_4852,N_1499,N_1163);
and U4853 (N_4853,N_1802,N_864);
and U4854 (N_4854,N_2474,N_1319);
or U4855 (N_4855,N_204,N_1126);
or U4856 (N_4856,N_2850,N_248);
or U4857 (N_4857,N_494,N_423);
nor U4858 (N_4858,N_560,N_2774);
and U4859 (N_4859,N_2563,N_1130);
nand U4860 (N_4860,N_1139,N_2107);
nor U4861 (N_4861,N_2039,N_905);
and U4862 (N_4862,N_105,N_2144);
nor U4863 (N_4863,N_2211,N_316);
nand U4864 (N_4864,N_805,N_865);
or U4865 (N_4865,N_1728,N_2826);
nor U4866 (N_4866,N_929,N_2889);
or U4867 (N_4867,N_1188,N_1007);
or U4868 (N_4868,N_2009,N_344);
or U4869 (N_4869,N_1418,N_885);
and U4870 (N_4870,N_1054,N_2658);
or U4871 (N_4871,N_1810,N_1024);
xnor U4872 (N_4872,N_1880,N_2142);
nor U4873 (N_4873,N_151,N_2716);
nand U4874 (N_4874,N_1400,N_370);
or U4875 (N_4875,N_1851,N_519);
and U4876 (N_4876,N_2066,N_2310);
xnor U4877 (N_4877,N_1734,N_1223);
xnor U4878 (N_4878,N_975,N_2107);
nand U4879 (N_4879,N_1696,N_361);
nand U4880 (N_4880,N_654,N_55);
or U4881 (N_4881,N_1313,N_1834);
and U4882 (N_4882,N_2468,N_2818);
nand U4883 (N_4883,N_503,N_2495);
nor U4884 (N_4884,N_2966,N_89);
nand U4885 (N_4885,N_2393,N_1331);
and U4886 (N_4886,N_2965,N_1756);
nand U4887 (N_4887,N_1959,N_1033);
xnor U4888 (N_4888,N_2885,N_1772);
nand U4889 (N_4889,N_339,N_1132);
or U4890 (N_4890,N_1057,N_242);
xor U4891 (N_4891,N_2258,N_637);
nand U4892 (N_4892,N_2624,N_1271);
or U4893 (N_4893,N_2368,N_2116);
nor U4894 (N_4894,N_1307,N_1448);
nand U4895 (N_4895,N_2929,N_2478);
xor U4896 (N_4896,N_1657,N_2046);
and U4897 (N_4897,N_2762,N_2774);
or U4898 (N_4898,N_101,N_1539);
nor U4899 (N_4899,N_1572,N_2132);
xor U4900 (N_4900,N_18,N_762);
nor U4901 (N_4901,N_352,N_1779);
nand U4902 (N_4902,N_57,N_2243);
and U4903 (N_4903,N_1361,N_2345);
nor U4904 (N_4904,N_841,N_2662);
nand U4905 (N_4905,N_2013,N_897);
nor U4906 (N_4906,N_1869,N_2346);
nor U4907 (N_4907,N_627,N_2658);
or U4908 (N_4908,N_960,N_1391);
nor U4909 (N_4909,N_2047,N_2610);
nand U4910 (N_4910,N_2906,N_247);
nor U4911 (N_4911,N_2135,N_470);
or U4912 (N_4912,N_496,N_2220);
nor U4913 (N_4913,N_1499,N_1466);
xor U4914 (N_4914,N_2098,N_2299);
nor U4915 (N_4915,N_1486,N_1918);
xor U4916 (N_4916,N_1818,N_965);
and U4917 (N_4917,N_805,N_1529);
xor U4918 (N_4918,N_2416,N_1275);
nor U4919 (N_4919,N_1278,N_2690);
and U4920 (N_4920,N_840,N_2209);
xnor U4921 (N_4921,N_1,N_2885);
nor U4922 (N_4922,N_2243,N_537);
nand U4923 (N_4923,N_270,N_2363);
nor U4924 (N_4924,N_376,N_2519);
or U4925 (N_4925,N_2635,N_1917);
and U4926 (N_4926,N_830,N_1322);
nor U4927 (N_4927,N_1884,N_2175);
or U4928 (N_4928,N_1000,N_2097);
or U4929 (N_4929,N_381,N_102);
xnor U4930 (N_4930,N_1115,N_1818);
or U4931 (N_4931,N_2373,N_1406);
nor U4932 (N_4932,N_710,N_1468);
nand U4933 (N_4933,N_1667,N_920);
nor U4934 (N_4934,N_303,N_606);
nand U4935 (N_4935,N_1824,N_1077);
and U4936 (N_4936,N_2347,N_2464);
nand U4937 (N_4937,N_598,N_2088);
nand U4938 (N_4938,N_2167,N_545);
nor U4939 (N_4939,N_2796,N_516);
nor U4940 (N_4940,N_1159,N_627);
or U4941 (N_4941,N_411,N_2313);
and U4942 (N_4942,N_2273,N_1511);
or U4943 (N_4943,N_2866,N_2086);
or U4944 (N_4944,N_984,N_1825);
nand U4945 (N_4945,N_437,N_697);
and U4946 (N_4946,N_214,N_1118);
nor U4947 (N_4947,N_1180,N_336);
xnor U4948 (N_4948,N_1432,N_1896);
xor U4949 (N_4949,N_1904,N_2014);
nand U4950 (N_4950,N_2454,N_738);
xor U4951 (N_4951,N_2147,N_2631);
and U4952 (N_4952,N_2263,N_116);
and U4953 (N_4953,N_2471,N_1832);
and U4954 (N_4954,N_637,N_2175);
and U4955 (N_4955,N_1291,N_2420);
xnor U4956 (N_4956,N_27,N_2258);
xor U4957 (N_4957,N_1398,N_2558);
or U4958 (N_4958,N_1214,N_2825);
nor U4959 (N_4959,N_1522,N_1855);
and U4960 (N_4960,N_2315,N_516);
nor U4961 (N_4961,N_2861,N_97);
nor U4962 (N_4962,N_2852,N_396);
nand U4963 (N_4963,N_2182,N_2012);
nor U4964 (N_4964,N_1400,N_2400);
nor U4965 (N_4965,N_1304,N_1651);
or U4966 (N_4966,N_1619,N_1404);
nand U4967 (N_4967,N_1379,N_1700);
xnor U4968 (N_4968,N_2363,N_1180);
and U4969 (N_4969,N_1003,N_15);
and U4970 (N_4970,N_583,N_1413);
xnor U4971 (N_4971,N_575,N_2335);
or U4972 (N_4972,N_1619,N_1417);
nor U4973 (N_4973,N_1679,N_2769);
and U4974 (N_4974,N_1476,N_2334);
xor U4975 (N_4975,N_478,N_1445);
nand U4976 (N_4976,N_2487,N_489);
xor U4977 (N_4977,N_572,N_1556);
and U4978 (N_4978,N_1183,N_455);
or U4979 (N_4979,N_2232,N_695);
nand U4980 (N_4980,N_1702,N_2789);
nor U4981 (N_4981,N_2987,N_1994);
or U4982 (N_4982,N_1944,N_537);
and U4983 (N_4983,N_1627,N_1518);
and U4984 (N_4984,N_2470,N_2083);
nor U4985 (N_4985,N_2897,N_1215);
or U4986 (N_4986,N_1446,N_1730);
and U4987 (N_4987,N_560,N_714);
and U4988 (N_4988,N_1128,N_1717);
and U4989 (N_4989,N_2536,N_1100);
xor U4990 (N_4990,N_142,N_1915);
nor U4991 (N_4991,N_819,N_1801);
or U4992 (N_4992,N_1759,N_1802);
xor U4993 (N_4993,N_2321,N_2722);
or U4994 (N_4994,N_1203,N_2817);
nand U4995 (N_4995,N_1548,N_1642);
and U4996 (N_4996,N_502,N_1243);
or U4997 (N_4997,N_745,N_800);
and U4998 (N_4998,N_1125,N_1296);
and U4999 (N_4999,N_182,N_119);
xor U5000 (N_5000,N_2224,N_752);
xor U5001 (N_5001,N_1774,N_1642);
xnor U5002 (N_5002,N_113,N_2572);
or U5003 (N_5003,N_1487,N_677);
xnor U5004 (N_5004,N_561,N_2366);
or U5005 (N_5005,N_1121,N_423);
or U5006 (N_5006,N_768,N_2464);
nand U5007 (N_5007,N_2107,N_1430);
xnor U5008 (N_5008,N_1446,N_2750);
nand U5009 (N_5009,N_2794,N_851);
nand U5010 (N_5010,N_1950,N_2412);
nor U5011 (N_5011,N_1539,N_2223);
nand U5012 (N_5012,N_320,N_259);
or U5013 (N_5013,N_866,N_2400);
and U5014 (N_5014,N_2306,N_537);
or U5015 (N_5015,N_18,N_1734);
nor U5016 (N_5016,N_2661,N_2813);
or U5017 (N_5017,N_1996,N_1112);
nand U5018 (N_5018,N_1630,N_279);
nor U5019 (N_5019,N_768,N_2219);
nand U5020 (N_5020,N_229,N_2781);
or U5021 (N_5021,N_1869,N_1773);
nand U5022 (N_5022,N_1370,N_1419);
and U5023 (N_5023,N_2531,N_620);
and U5024 (N_5024,N_130,N_128);
or U5025 (N_5025,N_764,N_2525);
or U5026 (N_5026,N_2860,N_45);
xor U5027 (N_5027,N_1284,N_1604);
and U5028 (N_5028,N_60,N_2990);
nor U5029 (N_5029,N_734,N_2644);
xnor U5030 (N_5030,N_1905,N_1189);
xnor U5031 (N_5031,N_1621,N_1913);
nand U5032 (N_5032,N_1156,N_2292);
and U5033 (N_5033,N_2151,N_1050);
nand U5034 (N_5034,N_1401,N_650);
and U5035 (N_5035,N_356,N_2030);
or U5036 (N_5036,N_1892,N_826);
xor U5037 (N_5037,N_723,N_4);
xor U5038 (N_5038,N_937,N_849);
nor U5039 (N_5039,N_1671,N_2092);
xnor U5040 (N_5040,N_171,N_2324);
xor U5041 (N_5041,N_1324,N_495);
and U5042 (N_5042,N_1801,N_1215);
xor U5043 (N_5043,N_762,N_2849);
nand U5044 (N_5044,N_733,N_2440);
nor U5045 (N_5045,N_810,N_11);
and U5046 (N_5046,N_1127,N_977);
nor U5047 (N_5047,N_1500,N_2062);
xnor U5048 (N_5048,N_2150,N_1556);
and U5049 (N_5049,N_109,N_2534);
xor U5050 (N_5050,N_356,N_1767);
and U5051 (N_5051,N_649,N_147);
nand U5052 (N_5052,N_2936,N_633);
nand U5053 (N_5053,N_1952,N_1155);
nand U5054 (N_5054,N_1986,N_2437);
and U5055 (N_5055,N_1536,N_747);
nand U5056 (N_5056,N_90,N_2275);
xor U5057 (N_5057,N_1375,N_514);
and U5058 (N_5058,N_2167,N_1161);
and U5059 (N_5059,N_343,N_912);
nor U5060 (N_5060,N_947,N_985);
nand U5061 (N_5061,N_2416,N_956);
xor U5062 (N_5062,N_2180,N_1624);
nor U5063 (N_5063,N_100,N_1759);
xnor U5064 (N_5064,N_146,N_444);
or U5065 (N_5065,N_2395,N_2076);
or U5066 (N_5066,N_942,N_2033);
and U5067 (N_5067,N_2199,N_2325);
or U5068 (N_5068,N_1627,N_1160);
nor U5069 (N_5069,N_2059,N_2650);
nor U5070 (N_5070,N_1913,N_766);
or U5071 (N_5071,N_2792,N_1924);
and U5072 (N_5072,N_41,N_322);
or U5073 (N_5073,N_1581,N_1441);
xor U5074 (N_5074,N_1285,N_724);
nand U5075 (N_5075,N_1853,N_1419);
nand U5076 (N_5076,N_2055,N_1620);
and U5077 (N_5077,N_1239,N_1924);
nand U5078 (N_5078,N_2835,N_1123);
and U5079 (N_5079,N_2230,N_937);
nand U5080 (N_5080,N_1873,N_438);
nand U5081 (N_5081,N_1005,N_450);
or U5082 (N_5082,N_1025,N_1295);
xor U5083 (N_5083,N_1263,N_1383);
or U5084 (N_5084,N_1752,N_584);
and U5085 (N_5085,N_91,N_730);
and U5086 (N_5086,N_2549,N_2096);
or U5087 (N_5087,N_343,N_2596);
or U5088 (N_5088,N_980,N_584);
nand U5089 (N_5089,N_2810,N_1436);
xor U5090 (N_5090,N_2954,N_1850);
nor U5091 (N_5091,N_2228,N_173);
and U5092 (N_5092,N_162,N_987);
or U5093 (N_5093,N_1391,N_2875);
xor U5094 (N_5094,N_1706,N_343);
nor U5095 (N_5095,N_1415,N_1758);
nand U5096 (N_5096,N_2194,N_1315);
nand U5097 (N_5097,N_975,N_524);
or U5098 (N_5098,N_2519,N_2662);
nand U5099 (N_5099,N_1955,N_903);
and U5100 (N_5100,N_2278,N_356);
xnor U5101 (N_5101,N_103,N_1570);
xnor U5102 (N_5102,N_2192,N_38);
nor U5103 (N_5103,N_1458,N_2564);
xnor U5104 (N_5104,N_2888,N_235);
xor U5105 (N_5105,N_1367,N_1881);
and U5106 (N_5106,N_9,N_218);
nand U5107 (N_5107,N_543,N_165);
or U5108 (N_5108,N_1646,N_2878);
nor U5109 (N_5109,N_1668,N_1101);
or U5110 (N_5110,N_992,N_400);
xor U5111 (N_5111,N_2988,N_2497);
or U5112 (N_5112,N_1664,N_1643);
and U5113 (N_5113,N_368,N_1501);
and U5114 (N_5114,N_1385,N_1034);
and U5115 (N_5115,N_1560,N_2921);
nand U5116 (N_5116,N_2639,N_1116);
xnor U5117 (N_5117,N_2918,N_1871);
nand U5118 (N_5118,N_1684,N_2014);
nand U5119 (N_5119,N_842,N_2105);
and U5120 (N_5120,N_2474,N_1127);
nand U5121 (N_5121,N_1161,N_1977);
nand U5122 (N_5122,N_652,N_2015);
nand U5123 (N_5123,N_1317,N_837);
xnor U5124 (N_5124,N_397,N_1341);
xnor U5125 (N_5125,N_1117,N_1768);
or U5126 (N_5126,N_1434,N_2177);
xor U5127 (N_5127,N_725,N_24);
xnor U5128 (N_5128,N_1145,N_1261);
and U5129 (N_5129,N_143,N_2943);
xnor U5130 (N_5130,N_1250,N_613);
xor U5131 (N_5131,N_1041,N_990);
or U5132 (N_5132,N_797,N_1880);
and U5133 (N_5133,N_27,N_1598);
xnor U5134 (N_5134,N_106,N_1067);
xnor U5135 (N_5135,N_1558,N_152);
nor U5136 (N_5136,N_2204,N_783);
nor U5137 (N_5137,N_1277,N_2665);
or U5138 (N_5138,N_1652,N_644);
nand U5139 (N_5139,N_1905,N_1144);
nor U5140 (N_5140,N_130,N_1149);
xor U5141 (N_5141,N_700,N_305);
and U5142 (N_5142,N_2594,N_490);
and U5143 (N_5143,N_1692,N_1029);
and U5144 (N_5144,N_2953,N_1019);
or U5145 (N_5145,N_1952,N_1242);
nor U5146 (N_5146,N_1986,N_792);
nor U5147 (N_5147,N_2572,N_1562);
and U5148 (N_5148,N_891,N_1982);
xor U5149 (N_5149,N_1714,N_223);
xor U5150 (N_5150,N_441,N_748);
nand U5151 (N_5151,N_2231,N_2916);
or U5152 (N_5152,N_1811,N_2867);
nand U5153 (N_5153,N_2457,N_2326);
xnor U5154 (N_5154,N_284,N_2245);
or U5155 (N_5155,N_2760,N_2685);
nand U5156 (N_5156,N_2980,N_2412);
and U5157 (N_5157,N_1674,N_773);
and U5158 (N_5158,N_1194,N_519);
and U5159 (N_5159,N_1097,N_1174);
and U5160 (N_5160,N_1089,N_704);
nand U5161 (N_5161,N_2110,N_559);
or U5162 (N_5162,N_2356,N_2752);
xnor U5163 (N_5163,N_214,N_416);
xor U5164 (N_5164,N_2527,N_555);
and U5165 (N_5165,N_2636,N_1110);
xor U5166 (N_5166,N_1295,N_246);
nor U5167 (N_5167,N_1536,N_1709);
nand U5168 (N_5168,N_2116,N_1290);
xor U5169 (N_5169,N_1743,N_1082);
xnor U5170 (N_5170,N_831,N_1239);
xnor U5171 (N_5171,N_114,N_965);
or U5172 (N_5172,N_562,N_2346);
nor U5173 (N_5173,N_2912,N_883);
nor U5174 (N_5174,N_1237,N_117);
or U5175 (N_5175,N_2114,N_2534);
and U5176 (N_5176,N_2822,N_507);
and U5177 (N_5177,N_1501,N_1749);
or U5178 (N_5178,N_2293,N_666);
nand U5179 (N_5179,N_2214,N_1004);
nand U5180 (N_5180,N_309,N_397);
xor U5181 (N_5181,N_1046,N_834);
nand U5182 (N_5182,N_2831,N_1801);
nor U5183 (N_5183,N_119,N_1814);
or U5184 (N_5184,N_2656,N_2050);
xor U5185 (N_5185,N_1036,N_163);
and U5186 (N_5186,N_396,N_2956);
xor U5187 (N_5187,N_613,N_440);
xnor U5188 (N_5188,N_1738,N_1162);
nor U5189 (N_5189,N_2788,N_2551);
nor U5190 (N_5190,N_1546,N_1966);
and U5191 (N_5191,N_2820,N_18);
nor U5192 (N_5192,N_893,N_16);
xnor U5193 (N_5193,N_946,N_941);
and U5194 (N_5194,N_867,N_1459);
nand U5195 (N_5195,N_1410,N_1662);
nand U5196 (N_5196,N_2268,N_2699);
or U5197 (N_5197,N_1648,N_1962);
nand U5198 (N_5198,N_1811,N_2883);
nor U5199 (N_5199,N_1368,N_2654);
or U5200 (N_5200,N_1639,N_1390);
and U5201 (N_5201,N_1124,N_1795);
nand U5202 (N_5202,N_246,N_486);
or U5203 (N_5203,N_2812,N_687);
nand U5204 (N_5204,N_2697,N_2733);
nor U5205 (N_5205,N_1095,N_913);
and U5206 (N_5206,N_1933,N_255);
xor U5207 (N_5207,N_2743,N_329);
nand U5208 (N_5208,N_213,N_2127);
or U5209 (N_5209,N_363,N_2988);
or U5210 (N_5210,N_1267,N_726);
nor U5211 (N_5211,N_896,N_930);
nand U5212 (N_5212,N_685,N_522);
nand U5213 (N_5213,N_1370,N_218);
nor U5214 (N_5214,N_1450,N_636);
nor U5215 (N_5215,N_1571,N_2898);
and U5216 (N_5216,N_635,N_1895);
nor U5217 (N_5217,N_2812,N_1070);
and U5218 (N_5218,N_2885,N_2224);
nand U5219 (N_5219,N_1937,N_903);
or U5220 (N_5220,N_372,N_1044);
nor U5221 (N_5221,N_718,N_743);
nand U5222 (N_5222,N_214,N_2170);
or U5223 (N_5223,N_1141,N_1534);
or U5224 (N_5224,N_1358,N_936);
or U5225 (N_5225,N_734,N_2695);
or U5226 (N_5226,N_2452,N_2435);
and U5227 (N_5227,N_661,N_1601);
and U5228 (N_5228,N_2802,N_2504);
xnor U5229 (N_5229,N_1914,N_2957);
nor U5230 (N_5230,N_2,N_1268);
or U5231 (N_5231,N_2759,N_2140);
and U5232 (N_5232,N_1592,N_2024);
nor U5233 (N_5233,N_2432,N_2330);
nand U5234 (N_5234,N_217,N_464);
and U5235 (N_5235,N_878,N_2385);
and U5236 (N_5236,N_1304,N_1121);
and U5237 (N_5237,N_455,N_662);
xor U5238 (N_5238,N_1815,N_1859);
or U5239 (N_5239,N_469,N_2731);
and U5240 (N_5240,N_678,N_2590);
or U5241 (N_5241,N_694,N_1789);
nand U5242 (N_5242,N_2787,N_2031);
nor U5243 (N_5243,N_1855,N_771);
and U5244 (N_5244,N_1149,N_2757);
nor U5245 (N_5245,N_2193,N_2318);
xor U5246 (N_5246,N_2017,N_2171);
nor U5247 (N_5247,N_39,N_913);
nand U5248 (N_5248,N_985,N_2379);
or U5249 (N_5249,N_2414,N_1099);
xnor U5250 (N_5250,N_2508,N_527);
nand U5251 (N_5251,N_373,N_451);
and U5252 (N_5252,N_2966,N_1535);
or U5253 (N_5253,N_2582,N_698);
nor U5254 (N_5254,N_331,N_2881);
xor U5255 (N_5255,N_87,N_1611);
xnor U5256 (N_5256,N_137,N_229);
nand U5257 (N_5257,N_1864,N_2228);
or U5258 (N_5258,N_2358,N_1429);
or U5259 (N_5259,N_2630,N_1124);
xnor U5260 (N_5260,N_1755,N_246);
nor U5261 (N_5261,N_427,N_2386);
and U5262 (N_5262,N_2692,N_844);
or U5263 (N_5263,N_1051,N_2502);
or U5264 (N_5264,N_1461,N_291);
and U5265 (N_5265,N_1442,N_1825);
or U5266 (N_5266,N_651,N_2123);
or U5267 (N_5267,N_102,N_2665);
nor U5268 (N_5268,N_1036,N_1541);
nand U5269 (N_5269,N_954,N_685);
nand U5270 (N_5270,N_2546,N_609);
nor U5271 (N_5271,N_2092,N_655);
xor U5272 (N_5272,N_1208,N_457);
and U5273 (N_5273,N_1284,N_1330);
nor U5274 (N_5274,N_2682,N_2158);
xor U5275 (N_5275,N_585,N_314);
or U5276 (N_5276,N_266,N_1527);
and U5277 (N_5277,N_2422,N_955);
or U5278 (N_5278,N_903,N_2716);
and U5279 (N_5279,N_2625,N_1682);
xnor U5280 (N_5280,N_2997,N_1579);
xnor U5281 (N_5281,N_1191,N_2515);
or U5282 (N_5282,N_1966,N_763);
and U5283 (N_5283,N_617,N_2769);
xor U5284 (N_5284,N_1864,N_2971);
and U5285 (N_5285,N_72,N_523);
nand U5286 (N_5286,N_560,N_2237);
xnor U5287 (N_5287,N_191,N_2109);
or U5288 (N_5288,N_2628,N_1626);
and U5289 (N_5289,N_755,N_2818);
nor U5290 (N_5290,N_1440,N_1516);
and U5291 (N_5291,N_141,N_489);
xnor U5292 (N_5292,N_2996,N_1781);
or U5293 (N_5293,N_998,N_2458);
nor U5294 (N_5294,N_1306,N_2408);
nand U5295 (N_5295,N_2821,N_2517);
and U5296 (N_5296,N_888,N_283);
nor U5297 (N_5297,N_1530,N_1411);
nor U5298 (N_5298,N_1339,N_1559);
or U5299 (N_5299,N_242,N_1012);
nand U5300 (N_5300,N_2779,N_2687);
xor U5301 (N_5301,N_1367,N_2044);
nand U5302 (N_5302,N_1920,N_1612);
xor U5303 (N_5303,N_2781,N_1742);
xor U5304 (N_5304,N_2166,N_2637);
and U5305 (N_5305,N_967,N_2371);
nand U5306 (N_5306,N_2754,N_884);
xor U5307 (N_5307,N_306,N_56);
and U5308 (N_5308,N_1255,N_1032);
and U5309 (N_5309,N_1750,N_681);
xor U5310 (N_5310,N_367,N_434);
and U5311 (N_5311,N_922,N_2950);
and U5312 (N_5312,N_2387,N_1235);
or U5313 (N_5313,N_2038,N_55);
or U5314 (N_5314,N_2168,N_2099);
or U5315 (N_5315,N_290,N_2125);
nor U5316 (N_5316,N_2378,N_746);
or U5317 (N_5317,N_2745,N_982);
xnor U5318 (N_5318,N_1038,N_1144);
nand U5319 (N_5319,N_303,N_1727);
nand U5320 (N_5320,N_258,N_2772);
xor U5321 (N_5321,N_660,N_1073);
and U5322 (N_5322,N_478,N_1252);
or U5323 (N_5323,N_2924,N_1607);
and U5324 (N_5324,N_1822,N_1603);
nand U5325 (N_5325,N_2717,N_1669);
xnor U5326 (N_5326,N_514,N_1544);
nand U5327 (N_5327,N_1054,N_65);
or U5328 (N_5328,N_2734,N_222);
and U5329 (N_5329,N_2973,N_315);
or U5330 (N_5330,N_2302,N_1016);
and U5331 (N_5331,N_547,N_2510);
nor U5332 (N_5332,N_936,N_1154);
and U5333 (N_5333,N_1514,N_2814);
and U5334 (N_5334,N_633,N_87);
xnor U5335 (N_5335,N_1898,N_1388);
and U5336 (N_5336,N_35,N_364);
or U5337 (N_5337,N_2754,N_500);
or U5338 (N_5338,N_1841,N_1930);
or U5339 (N_5339,N_2781,N_1083);
nand U5340 (N_5340,N_1580,N_896);
and U5341 (N_5341,N_1090,N_385);
and U5342 (N_5342,N_1769,N_2706);
and U5343 (N_5343,N_2638,N_1592);
and U5344 (N_5344,N_1833,N_1788);
or U5345 (N_5345,N_2403,N_1996);
or U5346 (N_5346,N_314,N_1885);
nor U5347 (N_5347,N_856,N_2192);
nor U5348 (N_5348,N_312,N_2278);
and U5349 (N_5349,N_1470,N_1378);
xnor U5350 (N_5350,N_1594,N_176);
nor U5351 (N_5351,N_1510,N_1237);
nand U5352 (N_5352,N_866,N_335);
xnor U5353 (N_5353,N_2989,N_2872);
xnor U5354 (N_5354,N_1313,N_1786);
or U5355 (N_5355,N_2827,N_2156);
or U5356 (N_5356,N_351,N_306);
xor U5357 (N_5357,N_2563,N_1426);
and U5358 (N_5358,N_241,N_290);
nor U5359 (N_5359,N_1318,N_2630);
or U5360 (N_5360,N_922,N_428);
nor U5361 (N_5361,N_1424,N_620);
nand U5362 (N_5362,N_1106,N_2487);
and U5363 (N_5363,N_1401,N_2020);
xor U5364 (N_5364,N_674,N_51);
nand U5365 (N_5365,N_1844,N_1102);
or U5366 (N_5366,N_2625,N_1121);
and U5367 (N_5367,N_1808,N_1600);
nor U5368 (N_5368,N_2262,N_2508);
nor U5369 (N_5369,N_502,N_1093);
and U5370 (N_5370,N_835,N_13);
xnor U5371 (N_5371,N_699,N_1049);
nor U5372 (N_5372,N_2749,N_334);
or U5373 (N_5373,N_31,N_1056);
and U5374 (N_5374,N_1260,N_1271);
xnor U5375 (N_5375,N_822,N_2172);
nor U5376 (N_5376,N_1851,N_1498);
or U5377 (N_5377,N_167,N_1591);
xor U5378 (N_5378,N_566,N_2564);
nor U5379 (N_5379,N_641,N_415);
nor U5380 (N_5380,N_236,N_1783);
nor U5381 (N_5381,N_844,N_1587);
xor U5382 (N_5382,N_1146,N_2243);
and U5383 (N_5383,N_1962,N_1390);
nand U5384 (N_5384,N_873,N_2434);
and U5385 (N_5385,N_850,N_1000);
xor U5386 (N_5386,N_622,N_739);
nand U5387 (N_5387,N_595,N_970);
or U5388 (N_5388,N_2614,N_1553);
and U5389 (N_5389,N_2210,N_1498);
nor U5390 (N_5390,N_1027,N_1646);
nor U5391 (N_5391,N_1858,N_606);
or U5392 (N_5392,N_216,N_1718);
nand U5393 (N_5393,N_1152,N_2962);
xor U5394 (N_5394,N_1027,N_98);
xnor U5395 (N_5395,N_2874,N_1734);
nand U5396 (N_5396,N_2555,N_2760);
and U5397 (N_5397,N_795,N_737);
or U5398 (N_5398,N_1794,N_155);
nor U5399 (N_5399,N_2388,N_985);
xor U5400 (N_5400,N_2948,N_1953);
nand U5401 (N_5401,N_1509,N_1799);
nand U5402 (N_5402,N_851,N_873);
and U5403 (N_5403,N_2351,N_2713);
xnor U5404 (N_5404,N_2942,N_898);
nor U5405 (N_5405,N_86,N_1079);
nand U5406 (N_5406,N_2108,N_835);
xnor U5407 (N_5407,N_2431,N_43);
and U5408 (N_5408,N_1740,N_1809);
or U5409 (N_5409,N_918,N_1372);
nor U5410 (N_5410,N_2974,N_763);
or U5411 (N_5411,N_1397,N_1737);
xnor U5412 (N_5412,N_61,N_757);
nor U5413 (N_5413,N_1272,N_2276);
nor U5414 (N_5414,N_2432,N_1150);
xor U5415 (N_5415,N_2313,N_1570);
nand U5416 (N_5416,N_817,N_2167);
nor U5417 (N_5417,N_2997,N_569);
xnor U5418 (N_5418,N_2052,N_1153);
nand U5419 (N_5419,N_2139,N_2198);
nor U5420 (N_5420,N_235,N_1105);
nand U5421 (N_5421,N_2818,N_1221);
xor U5422 (N_5422,N_606,N_2390);
or U5423 (N_5423,N_1480,N_2505);
and U5424 (N_5424,N_2640,N_991);
and U5425 (N_5425,N_145,N_60);
xnor U5426 (N_5426,N_2570,N_1304);
nand U5427 (N_5427,N_1134,N_2845);
nor U5428 (N_5428,N_2022,N_2935);
nor U5429 (N_5429,N_502,N_1546);
xor U5430 (N_5430,N_1316,N_446);
xor U5431 (N_5431,N_1068,N_2718);
or U5432 (N_5432,N_2883,N_2291);
nor U5433 (N_5433,N_1295,N_1339);
and U5434 (N_5434,N_851,N_2809);
or U5435 (N_5435,N_650,N_2376);
nand U5436 (N_5436,N_423,N_932);
nor U5437 (N_5437,N_365,N_1326);
nand U5438 (N_5438,N_2822,N_1723);
xnor U5439 (N_5439,N_2094,N_2790);
nor U5440 (N_5440,N_515,N_2431);
nor U5441 (N_5441,N_2566,N_2588);
nor U5442 (N_5442,N_676,N_1480);
or U5443 (N_5443,N_1293,N_556);
nand U5444 (N_5444,N_983,N_1560);
and U5445 (N_5445,N_2321,N_1856);
or U5446 (N_5446,N_2403,N_1370);
xnor U5447 (N_5447,N_2731,N_1582);
or U5448 (N_5448,N_1516,N_290);
and U5449 (N_5449,N_2778,N_2115);
nand U5450 (N_5450,N_1723,N_575);
and U5451 (N_5451,N_2305,N_1914);
nand U5452 (N_5452,N_2159,N_1290);
nand U5453 (N_5453,N_2673,N_1526);
or U5454 (N_5454,N_1256,N_2977);
xor U5455 (N_5455,N_1642,N_319);
nand U5456 (N_5456,N_30,N_48);
xnor U5457 (N_5457,N_188,N_1385);
nor U5458 (N_5458,N_2393,N_2983);
or U5459 (N_5459,N_181,N_2613);
nand U5460 (N_5460,N_1313,N_2071);
and U5461 (N_5461,N_1038,N_2383);
or U5462 (N_5462,N_2029,N_843);
nand U5463 (N_5463,N_1982,N_523);
nor U5464 (N_5464,N_591,N_633);
nor U5465 (N_5465,N_245,N_1779);
and U5466 (N_5466,N_1384,N_2659);
and U5467 (N_5467,N_2962,N_2731);
nand U5468 (N_5468,N_2130,N_2622);
and U5469 (N_5469,N_1044,N_1311);
xor U5470 (N_5470,N_337,N_732);
xor U5471 (N_5471,N_1230,N_1923);
nand U5472 (N_5472,N_2604,N_2886);
nor U5473 (N_5473,N_35,N_2459);
and U5474 (N_5474,N_289,N_2409);
or U5475 (N_5475,N_2014,N_2434);
nor U5476 (N_5476,N_567,N_2695);
nor U5477 (N_5477,N_303,N_1986);
nand U5478 (N_5478,N_1241,N_2039);
or U5479 (N_5479,N_2384,N_1068);
nor U5480 (N_5480,N_1444,N_1016);
nor U5481 (N_5481,N_979,N_3);
and U5482 (N_5482,N_2267,N_746);
nand U5483 (N_5483,N_347,N_2255);
nor U5484 (N_5484,N_1668,N_2984);
nand U5485 (N_5485,N_300,N_1361);
and U5486 (N_5486,N_1830,N_578);
nor U5487 (N_5487,N_1215,N_1305);
xnor U5488 (N_5488,N_380,N_2945);
or U5489 (N_5489,N_1856,N_1541);
xnor U5490 (N_5490,N_131,N_2239);
and U5491 (N_5491,N_2830,N_536);
nor U5492 (N_5492,N_869,N_2751);
nand U5493 (N_5493,N_2383,N_683);
xor U5494 (N_5494,N_1472,N_1432);
and U5495 (N_5495,N_861,N_2545);
and U5496 (N_5496,N_2974,N_880);
nor U5497 (N_5497,N_1569,N_2404);
nor U5498 (N_5498,N_1229,N_2769);
and U5499 (N_5499,N_170,N_454);
or U5500 (N_5500,N_2751,N_1922);
or U5501 (N_5501,N_1018,N_1125);
nand U5502 (N_5502,N_1837,N_138);
nand U5503 (N_5503,N_389,N_1662);
nor U5504 (N_5504,N_643,N_1966);
nor U5505 (N_5505,N_2080,N_132);
or U5506 (N_5506,N_1905,N_576);
and U5507 (N_5507,N_676,N_1490);
nor U5508 (N_5508,N_143,N_1679);
xnor U5509 (N_5509,N_1316,N_1448);
and U5510 (N_5510,N_1490,N_1428);
or U5511 (N_5511,N_2355,N_1732);
nand U5512 (N_5512,N_1885,N_319);
nor U5513 (N_5513,N_912,N_1556);
xor U5514 (N_5514,N_2987,N_1781);
nand U5515 (N_5515,N_2375,N_2555);
or U5516 (N_5516,N_28,N_2845);
nand U5517 (N_5517,N_2270,N_1461);
nand U5518 (N_5518,N_1681,N_1443);
and U5519 (N_5519,N_2061,N_1043);
nand U5520 (N_5520,N_927,N_662);
nor U5521 (N_5521,N_727,N_2931);
nor U5522 (N_5522,N_1285,N_423);
nand U5523 (N_5523,N_156,N_2646);
or U5524 (N_5524,N_991,N_1770);
nand U5525 (N_5525,N_1390,N_1075);
and U5526 (N_5526,N_1982,N_1211);
nand U5527 (N_5527,N_2708,N_1397);
and U5528 (N_5528,N_129,N_569);
nor U5529 (N_5529,N_2245,N_2738);
or U5530 (N_5530,N_2561,N_1942);
and U5531 (N_5531,N_2721,N_1632);
nand U5532 (N_5532,N_1760,N_541);
and U5533 (N_5533,N_1495,N_2976);
nor U5534 (N_5534,N_1204,N_92);
nor U5535 (N_5535,N_441,N_1511);
and U5536 (N_5536,N_2898,N_2252);
and U5537 (N_5537,N_1457,N_2932);
or U5538 (N_5538,N_2340,N_699);
or U5539 (N_5539,N_987,N_1979);
nor U5540 (N_5540,N_1779,N_1031);
or U5541 (N_5541,N_1092,N_2279);
and U5542 (N_5542,N_2479,N_2918);
or U5543 (N_5543,N_1367,N_2442);
and U5544 (N_5544,N_1726,N_1380);
and U5545 (N_5545,N_1147,N_924);
nand U5546 (N_5546,N_2217,N_843);
xnor U5547 (N_5547,N_128,N_207);
nand U5548 (N_5548,N_1666,N_517);
nor U5549 (N_5549,N_1501,N_78);
nor U5550 (N_5550,N_352,N_1219);
xor U5551 (N_5551,N_2114,N_2134);
or U5552 (N_5552,N_2591,N_2337);
and U5553 (N_5553,N_2576,N_702);
and U5554 (N_5554,N_2496,N_1062);
xnor U5555 (N_5555,N_286,N_211);
nor U5556 (N_5556,N_1048,N_1824);
xnor U5557 (N_5557,N_2765,N_2572);
xor U5558 (N_5558,N_939,N_1673);
or U5559 (N_5559,N_903,N_1662);
and U5560 (N_5560,N_2637,N_2549);
nand U5561 (N_5561,N_2491,N_137);
nor U5562 (N_5562,N_1305,N_2446);
and U5563 (N_5563,N_927,N_1845);
or U5564 (N_5564,N_2493,N_1299);
or U5565 (N_5565,N_17,N_1297);
xor U5566 (N_5566,N_1021,N_250);
nand U5567 (N_5567,N_2212,N_2669);
or U5568 (N_5568,N_1169,N_923);
xor U5569 (N_5569,N_12,N_2061);
nand U5570 (N_5570,N_694,N_1368);
nor U5571 (N_5571,N_854,N_2979);
and U5572 (N_5572,N_2659,N_494);
nor U5573 (N_5573,N_1601,N_1106);
nor U5574 (N_5574,N_2769,N_1301);
nand U5575 (N_5575,N_1216,N_1102);
nand U5576 (N_5576,N_154,N_577);
nor U5577 (N_5577,N_2410,N_2979);
xor U5578 (N_5578,N_2556,N_1374);
or U5579 (N_5579,N_1579,N_622);
nor U5580 (N_5580,N_2284,N_805);
and U5581 (N_5581,N_2156,N_826);
or U5582 (N_5582,N_1178,N_2549);
xnor U5583 (N_5583,N_1204,N_2777);
xnor U5584 (N_5584,N_990,N_499);
nor U5585 (N_5585,N_412,N_510);
or U5586 (N_5586,N_2157,N_2385);
or U5587 (N_5587,N_356,N_3);
and U5588 (N_5588,N_2125,N_1549);
and U5589 (N_5589,N_2952,N_862);
nor U5590 (N_5590,N_2401,N_412);
xnor U5591 (N_5591,N_918,N_540);
and U5592 (N_5592,N_2260,N_2582);
and U5593 (N_5593,N_1273,N_1294);
or U5594 (N_5594,N_775,N_2229);
and U5595 (N_5595,N_527,N_2941);
nand U5596 (N_5596,N_2550,N_1821);
and U5597 (N_5597,N_2634,N_1679);
and U5598 (N_5598,N_1428,N_2861);
and U5599 (N_5599,N_1072,N_1911);
or U5600 (N_5600,N_2356,N_1176);
nor U5601 (N_5601,N_2916,N_2088);
or U5602 (N_5602,N_2487,N_469);
or U5603 (N_5603,N_1129,N_2778);
nand U5604 (N_5604,N_2203,N_1533);
xnor U5605 (N_5605,N_1993,N_609);
or U5606 (N_5606,N_1661,N_388);
nor U5607 (N_5607,N_1390,N_2757);
and U5608 (N_5608,N_709,N_2700);
nor U5609 (N_5609,N_2988,N_2605);
nor U5610 (N_5610,N_1782,N_816);
nand U5611 (N_5611,N_377,N_1639);
xnor U5612 (N_5612,N_2818,N_1509);
nand U5613 (N_5613,N_2402,N_1375);
nand U5614 (N_5614,N_256,N_1377);
and U5615 (N_5615,N_2993,N_636);
and U5616 (N_5616,N_1915,N_37);
and U5617 (N_5617,N_989,N_2794);
or U5618 (N_5618,N_2527,N_1515);
and U5619 (N_5619,N_2869,N_513);
nor U5620 (N_5620,N_80,N_713);
and U5621 (N_5621,N_1618,N_2285);
xor U5622 (N_5622,N_18,N_936);
nand U5623 (N_5623,N_587,N_2159);
xnor U5624 (N_5624,N_1542,N_759);
xnor U5625 (N_5625,N_2611,N_2632);
and U5626 (N_5626,N_2750,N_54);
nor U5627 (N_5627,N_1740,N_141);
and U5628 (N_5628,N_29,N_121);
nor U5629 (N_5629,N_2756,N_1885);
or U5630 (N_5630,N_1971,N_1271);
nand U5631 (N_5631,N_51,N_940);
xnor U5632 (N_5632,N_1931,N_2559);
nor U5633 (N_5633,N_1441,N_1379);
and U5634 (N_5634,N_1729,N_1449);
nand U5635 (N_5635,N_701,N_1435);
nand U5636 (N_5636,N_2071,N_428);
nor U5637 (N_5637,N_2113,N_835);
or U5638 (N_5638,N_626,N_2632);
nand U5639 (N_5639,N_1155,N_514);
xor U5640 (N_5640,N_365,N_1928);
nand U5641 (N_5641,N_1756,N_2123);
or U5642 (N_5642,N_410,N_1650);
xor U5643 (N_5643,N_1397,N_2608);
or U5644 (N_5644,N_2276,N_1057);
and U5645 (N_5645,N_2788,N_2181);
nand U5646 (N_5646,N_1973,N_2805);
or U5647 (N_5647,N_96,N_1410);
xnor U5648 (N_5648,N_2159,N_2043);
and U5649 (N_5649,N_2456,N_1456);
xnor U5650 (N_5650,N_2890,N_410);
or U5651 (N_5651,N_508,N_2280);
nand U5652 (N_5652,N_1565,N_1490);
or U5653 (N_5653,N_361,N_1214);
or U5654 (N_5654,N_1008,N_2133);
or U5655 (N_5655,N_478,N_294);
or U5656 (N_5656,N_1814,N_2674);
nand U5657 (N_5657,N_1910,N_2791);
xnor U5658 (N_5658,N_484,N_2392);
or U5659 (N_5659,N_1982,N_1282);
or U5660 (N_5660,N_2885,N_988);
nand U5661 (N_5661,N_724,N_2910);
nor U5662 (N_5662,N_81,N_2650);
nand U5663 (N_5663,N_2455,N_2587);
nand U5664 (N_5664,N_1646,N_576);
nand U5665 (N_5665,N_1439,N_781);
and U5666 (N_5666,N_1294,N_133);
nand U5667 (N_5667,N_2821,N_2180);
xnor U5668 (N_5668,N_1031,N_2524);
nand U5669 (N_5669,N_779,N_1811);
xor U5670 (N_5670,N_596,N_1280);
nor U5671 (N_5671,N_515,N_536);
or U5672 (N_5672,N_2202,N_2332);
and U5673 (N_5673,N_364,N_1266);
nor U5674 (N_5674,N_2041,N_1427);
or U5675 (N_5675,N_2641,N_654);
nand U5676 (N_5676,N_845,N_2377);
and U5677 (N_5677,N_2401,N_2269);
and U5678 (N_5678,N_2272,N_534);
or U5679 (N_5679,N_2185,N_1490);
or U5680 (N_5680,N_178,N_2200);
nand U5681 (N_5681,N_936,N_1988);
and U5682 (N_5682,N_1742,N_81);
nand U5683 (N_5683,N_695,N_1933);
nand U5684 (N_5684,N_880,N_6);
xnor U5685 (N_5685,N_805,N_2687);
or U5686 (N_5686,N_629,N_1279);
xor U5687 (N_5687,N_2290,N_1183);
and U5688 (N_5688,N_2430,N_1098);
or U5689 (N_5689,N_2296,N_1731);
and U5690 (N_5690,N_653,N_2313);
xor U5691 (N_5691,N_144,N_563);
or U5692 (N_5692,N_2538,N_969);
nand U5693 (N_5693,N_1582,N_2195);
or U5694 (N_5694,N_1602,N_502);
xnor U5695 (N_5695,N_374,N_1058);
and U5696 (N_5696,N_2326,N_2214);
and U5697 (N_5697,N_1048,N_2980);
or U5698 (N_5698,N_1652,N_1391);
xnor U5699 (N_5699,N_425,N_2634);
nand U5700 (N_5700,N_2014,N_1913);
nor U5701 (N_5701,N_2122,N_1231);
nor U5702 (N_5702,N_1552,N_2591);
and U5703 (N_5703,N_2455,N_2956);
nand U5704 (N_5704,N_2484,N_2019);
and U5705 (N_5705,N_1547,N_904);
and U5706 (N_5706,N_1825,N_746);
and U5707 (N_5707,N_80,N_617);
nand U5708 (N_5708,N_23,N_2715);
xnor U5709 (N_5709,N_561,N_1841);
nand U5710 (N_5710,N_688,N_92);
xnor U5711 (N_5711,N_2655,N_2316);
nand U5712 (N_5712,N_2734,N_447);
or U5713 (N_5713,N_2725,N_1857);
or U5714 (N_5714,N_1681,N_1680);
xnor U5715 (N_5715,N_280,N_2235);
nor U5716 (N_5716,N_2945,N_725);
and U5717 (N_5717,N_2336,N_1792);
xor U5718 (N_5718,N_1121,N_1640);
xor U5719 (N_5719,N_1613,N_142);
or U5720 (N_5720,N_1815,N_170);
xnor U5721 (N_5721,N_165,N_1590);
nand U5722 (N_5722,N_2270,N_2480);
nor U5723 (N_5723,N_905,N_2288);
xor U5724 (N_5724,N_1700,N_781);
or U5725 (N_5725,N_2280,N_712);
nand U5726 (N_5726,N_287,N_1568);
xnor U5727 (N_5727,N_1980,N_416);
xnor U5728 (N_5728,N_2148,N_396);
and U5729 (N_5729,N_2416,N_2918);
or U5730 (N_5730,N_723,N_109);
nor U5731 (N_5731,N_2656,N_1606);
and U5732 (N_5732,N_2362,N_1102);
nand U5733 (N_5733,N_185,N_2429);
nand U5734 (N_5734,N_2242,N_1464);
and U5735 (N_5735,N_1342,N_1423);
xnor U5736 (N_5736,N_1968,N_2447);
xnor U5737 (N_5737,N_696,N_315);
or U5738 (N_5738,N_999,N_182);
nor U5739 (N_5739,N_2284,N_2485);
nor U5740 (N_5740,N_834,N_807);
xnor U5741 (N_5741,N_1895,N_1973);
and U5742 (N_5742,N_2605,N_2415);
xor U5743 (N_5743,N_2130,N_887);
and U5744 (N_5744,N_2815,N_2064);
nor U5745 (N_5745,N_1501,N_1181);
and U5746 (N_5746,N_638,N_2780);
xor U5747 (N_5747,N_1716,N_1779);
and U5748 (N_5748,N_142,N_2138);
nor U5749 (N_5749,N_880,N_1319);
and U5750 (N_5750,N_779,N_2077);
xnor U5751 (N_5751,N_2282,N_2636);
nor U5752 (N_5752,N_562,N_675);
nor U5753 (N_5753,N_618,N_797);
nand U5754 (N_5754,N_2352,N_1707);
nor U5755 (N_5755,N_2375,N_23);
and U5756 (N_5756,N_913,N_1304);
or U5757 (N_5757,N_690,N_2650);
xor U5758 (N_5758,N_2982,N_2168);
and U5759 (N_5759,N_607,N_1967);
xor U5760 (N_5760,N_1094,N_1058);
and U5761 (N_5761,N_306,N_1945);
nand U5762 (N_5762,N_289,N_1709);
and U5763 (N_5763,N_2391,N_2741);
nand U5764 (N_5764,N_1546,N_806);
or U5765 (N_5765,N_580,N_1131);
nand U5766 (N_5766,N_459,N_2397);
nor U5767 (N_5767,N_2311,N_1865);
nor U5768 (N_5768,N_2577,N_1980);
xor U5769 (N_5769,N_2498,N_2654);
nand U5770 (N_5770,N_2047,N_1764);
nand U5771 (N_5771,N_2480,N_2375);
or U5772 (N_5772,N_2328,N_1760);
xor U5773 (N_5773,N_2780,N_1153);
and U5774 (N_5774,N_2759,N_2170);
xnor U5775 (N_5775,N_2618,N_436);
nand U5776 (N_5776,N_776,N_2041);
or U5777 (N_5777,N_816,N_2793);
and U5778 (N_5778,N_2051,N_746);
or U5779 (N_5779,N_589,N_2825);
xnor U5780 (N_5780,N_2850,N_1279);
xnor U5781 (N_5781,N_2508,N_1350);
and U5782 (N_5782,N_2216,N_2444);
or U5783 (N_5783,N_1772,N_442);
nor U5784 (N_5784,N_44,N_1775);
and U5785 (N_5785,N_889,N_2084);
xnor U5786 (N_5786,N_727,N_867);
and U5787 (N_5787,N_839,N_2161);
nor U5788 (N_5788,N_455,N_2206);
nand U5789 (N_5789,N_1188,N_1832);
xor U5790 (N_5790,N_1576,N_2492);
and U5791 (N_5791,N_690,N_752);
xnor U5792 (N_5792,N_2929,N_1913);
or U5793 (N_5793,N_795,N_153);
and U5794 (N_5794,N_2122,N_1720);
xor U5795 (N_5795,N_2367,N_2618);
xor U5796 (N_5796,N_2303,N_1505);
xor U5797 (N_5797,N_477,N_123);
nand U5798 (N_5798,N_1933,N_2740);
and U5799 (N_5799,N_1555,N_1522);
xor U5800 (N_5800,N_1275,N_730);
and U5801 (N_5801,N_327,N_1224);
xor U5802 (N_5802,N_1862,N_2757);
nand U5803 (N_5803,N_2819,N_1388);
and U5804 (N_5804,N_723,N_1020);
nand U5805 (N_5805,N_1235,N_878);
nor U5806 (N_5806,N_2028,N_2310);
nand U5807 (N_5807,N_923,N_628);
xor U5808 (N_5808,N_281,N_2111);
nand U5809 (N_5809,N_317,N_589);
nor U5810 (N_5810,N_203,N_1548);
xor U5811 (N_5811,N_2390,N_1303);
nor U5812 (N_5812,N_2897,N_2950);
and U5813 (N_5813,N_1951,N_1843);
nor U5814 (N_5814,N_1225,N_1641);
or U5815 (N_5815,N_1022,N_1044);
nor U5816 (N_5816,N_1632,N_62);
xnor U5817 (N_5817,N_668,N_1333);
or U5818 (N_5818,N_2436,N_1832);
xor U5819 (N_5819,N_2227,N_1810);
and U5820 (N_5820,N_1852,N_2040);
or U5821 (N_5821,N_1279,N_1493);
xor U5822 (N_5822,N_2849,N_2091);
nand U5823 (N_5823,N_415,N_2071);
nor U5824 (N_5824,N_2852,N_1331);
nor U5825 (N_5825,N_170,N_694);
nor U5826 (N_5826,N_203,N_332);
nand U5827 (N_5827,N_1869,N_2392);
or U5828 (N_5828,N_2857,N_157);
xor U5829 (N_5829,N_1102,N_2689);
and U5830 (N_5830,N_2728,N_2643);
xor U5831 (N_5831,N_2482,N_2102);
nor U5832 (N_5832,N_898,N_493);
nor U5833 (N_5833,N_2836,N_407);
nor U5834 (N_5834,N_2971,N_119);
or U5835 (N_5835,N_855,N_250);
and U5836 (N_5836,N_2854,N_1808);
and U5837 (N_5837,N_284,N_2238);
nor U5838 (N_5838,N_437,N_1945);
nand U5839 (N_5839,N_523,N_1263);
and U5840 (N_5840,N_1914,N_372);
nand U5841 (N_5841,N_328,N_292);
or U5842 (N_5842,N_2236,N_41);
nand U5843 (N_5843,N_85,N_2178);
and U5844 (N_5844,N_2247,N_1813);
nand U5845 (N_5845,N_2354,N_2212);
or U5846 (N_5846,N_712,N_305);
xnor U5847 (N_5847,N_401,N_1910);
xnor U5848 (N_5848,N_2417,N_2232);
nor U5849 (N_5849,N_1273,N_2765);
or U5850 (N_5850,N_1228,N_43);
xor U5851 (N_5851,N_1703,N_2954);
xor U5852 (N_5852,N_962,N_625);
xnor U5853 (N_5853,N_1399,N_2776);
and U5854 (N_5854,N_52,N_840);
nand U5855 (N_5855,N_1869,N_2223);
xor U5856 (N_5856,N_1338,N_1360);
xor U5857 (N_5857,N_2323,N_1530);
or U5858 (N_5858,N_483,N_2559);
xor U5859 (N_5859,N_634,N_2959);
or U5860 (N_5860,N_1655,N_1333);
or U5861 (N_5861,N_291,N_1401);
xnor U5862 (N_5862,N_1413,N_2955);
xor U5863 (N_5863,N_2073,N_1465);
nor U5864 (N_5864,N_617,N_391);
xor U5865 (N_5865,N_2090,N_1282);
nand U5866 (N_5866,N_98,N_1718);
or U5867 (N_5867,N_2139,N_62);
nor U5868 (N_5868,N_1381,N_2896);
or U5869 (N_5869,N_74,N_1840);
or U5870 (N_5870,N_609,N_2764);
or U5871 (N_5871,N_358,N_851);
or U5872 (N_5872,N_2282,N_1184);
or U5873 (N_5873,N_2894,N_1563);
nor U5874 (N_5874,N_902,N_1187);
nor U5875 (N_5875,N_2045,N_616);
nand U5876 (N_5876,N_2128,N_2962);
or U5877 (N_5877,N_686,N_1722);
nand U5878 (N_5878,N_2889,N_2372);
nor U5879 (N_5879,N_2750,N_2105);
xnor U5880 (N_5880,N_2233,N_1631);
and U5881 (N_5881,N_1505,N_871);
or U5882 (N_5882,N_1123,N_215);
nor U5883 (N_5883,N_635,N_2964);
nand U5884 (N_5884,N_1732,N_1556);
or U5885 (N_5885,N_800,N_2712);
and U5886 (N_5886,N_2289,N_125);
xor U5887 (N_5887,N_257,N_2145);
and U5888 (N_5888,N_2890,N_933);
xnor U5889 (N_5889,N_135,N_867);
nor U5890 (N_5890,N_2272,N_1260);
nand U5891 (N_5891,N_726,N_2706);
nor U5892 (N_5892,N_638,N_2375);
and U5893 (N_5893,N_903,N_1201);
nor U5894 (N_5894,N_1081,N_1772);
and U5895 (N_5895,N_1800,N_1808);
nand U5896 (N_5896,N_562,N_1693);
xnor U5897 (N_5897,N_2422,N_318);
xor U5898 (N_5898,N_2958,N_2976);
xnor U5899 (N_5899,N_2055,N_2497);
or U5900 (N_5900,N_874,N_504);
or U5901 (N_5901,N_440,N_2479);
xor U5902 (N_5902,N_2876,N_811);
or U5903 (N_5903,N_2097,N_1935);
nor U5904 (N_5904,N_1185,N_35);
or U5905 (N_5905,N_1637,N_341);
xor U5906 (N_5906,N_1077,N_866);
nand U5907 (N_5907,N_587,N_2247);
and U5908 (N_5908,N_1708,N_286);
or U5909 (N_5909,N_1469,N_1390);
or U5910 (N_5910,N_1820,N_2750);
nand U5911 (N_5911,N_95,N_2692);
nand U5912 (N_5912,N_99,N_1529);
nand U5913 (N_5913,N_1413,N_455);
xor U5914 (N_5914,N_2814,N_843);
nand U5915 (N_5915,N_2155,N_1948);
and U5916 (N_5916,N_1151,N_340);
or U5917 (N_5917,N_1243,N_10);
nor U5918 (N_5918,N_2528,N_1371);
xnor U5919 (N_5919,N_1702,N_797);
nand U5920 (N_5920,N_2212,N_1479);
and U5921 (N_5921,N_807,N_2006);
nand U5922 (N_5922,N_2955,N_308);
nand U5923 (N_5923,N_2723,N_1635);
and U5924 (N_5924,N_810,N_1792);
and U5925 (N_5925,N_2372,N_2911);
nor U5926 (N_5926,N_2910,N_2404);
xnor U5927 (N_5927,N_1458,N_2176);
or U5928 (N_5928,N_1039,N_1516);
or U5929 (N_5929,N_640,N_192);
or U5930 (N_5930,N_1674,N_977);
nor U5931 (N_5931,N_1546,N_2197);
xnor U5932 (N_5932,N_2108,N_1822);
xnor U5933 (N_5933,N_1974,N_2719);
nand U5934 (N_5934,N_972,N_714);
and U5935 (N_5935,N_966,N_147);
xnor U5936 (N_5936,N_495,N_1682);
xnor U5937 (N_5937,N_1319,N_2901);
nor U5938 (N_5938,N_2972,N_2275);
or U5939 (N_5939,N_1697,N_329);
nand U5940 (N_5940,N_1495,N_733);
or U5941 (N_5941,N_416,N_1091);
nor U5942 (N_5942,N_2596,N_889);
nor U5943 (N_5943,N_2313,N_1475);
or U5944 (N_5944,N_415,N_1908);
and U5945 (N_5945,N_495,N_1517);
or U5946 (N_5946,N_2623,N_2741);
and U5947 (N_5947,N_711,N_1902);
or U5948 (N_5948,N_2314,N_1593);
and U5949 (N_5949,N_326,N_417);
nor U5950 (N_5950,N_431,N_1217);
nor U5951 (N_5951,N_953,N_2197);
or U5952 (N_5952,N_728,N_214);
xnor U5953 (N_5953,N_436,N_1762);
nor U5954 (N_5954,N_854,N_1960);
and U5955 (N_5955,N_738,N_1111);
nand U5956 (N_5956,N_551,N_1399);
or U5957 (N_5957,N_228,N_2037);
xnor U5958 (N_5958,N_410,N_2634);
or U5959 (N_5959,N_1615,N_2761);
xnor U5960 (N_5960,N_2985,N_1793);
and U5961 (N_5961,N_1675,N_1483);
nor U5962 (N_5962,N_2500,N_1678);
nor U5963 (N_5963,N_1928,N_664);
and U5964 (N_5964,N_1651,N_1491);
xor U5965 (N_5965,N_1639,N_1165);
xor U5966 (N_5966,N_2627,N_347);
nand U5967 (N_5967,N_24,N_1062);
xnor U5968 (N_5968,N_2555,N_325);
xnor U5969 (N_5969,N_1185,N_1212);
nor U5970 (N_5970,N_2287,N_2454);
nand U5971 (N_5971,N_2308,N_1612);
or U5972 (N_5972,N_1923,N_1075);
nor U5973 (N_5973,N_475,N_1725);
xnor U5974 (N_5974,N_1861,N_2580);
xnor U5975 (N_5975,N_2292,N_414);
and U5976 (N_5976,N_496,N_2373);
nand U5977 (N_5977,N_1162,N_1761);
nand U5978 (N_5978,N_1068,N_2320);
or U5979 (N_5979,N_107,N_1564);
nand U5980 (N_5980,N_2542,N_489);
xor U5981 (N_5981,N_1953,N_990);
and U5982 (N_5982,N_461,N_2291);
nor U5983 (N_5983,N_1880,N_1432);
xor U5984 (N_5984,N_2780,N_2046);
and U5985 (N_5985,N_1753,N_1145);
nand U5986 (N_5986,N_1192,N_1175);
or U5987 (N_5987,N_2421,N_229);
or U5988 (N_5988,N_1903,N_1828);
nand U5989 (N_5989,N_1032,N_1088);
xor U5990 (N_5990,N_297,N_677);
or U5991 (N_5991,N_2886,N_2510);
and U5992 (N_5992,N_2985,N_73);
xnor U5993 (N_5993,N_1906,N_2474);
and U5994 (N_5994,N_2940,N_1343);
and U5995 (N_5995,N_1500,N_2658);
xnor U5996 (N_5996,N_2432,N_1454);
and U5997 (N_5997,N_1108,N_328);
xor U5998 (N_5998,N_152,N_2);
and U5999 (N_5999,N_1437,N_2562);
nand U6000 (N_6000,N_4911,N_3755);
nor U6001 (N_6001,N_3221,N_5197);
nand U6002 (N_6002,N_3013,N_3108);
xor U6003 (N_6003,N_4376,N_3361);
xor U6004 (N_6004,N_3910,N_3200);
and U6005 (N_6005,N_4561,N_4651);
and U6006 (N_6006,N_5876,N_5302);
nor U6007 (N_6007,N_3263,N_3109);
and U6008 (N_6008,N_4889,N_3416);
nor U6009 (N_6009,N_4163,N_5211);
xnor U6010 (N_6010,N_3867,N_4224);
or U6011 (N_6011,N_4565,N_5405);
or U6012 (N_6012,N_5261,N_5766);
or U6013 (N_6013,N_5137,N_5916);
or U6014 (N_6014,N_4257,N_5143);
nor U6015 (N_6015,N_4299,N_3826);
nor U6016 (N_6016,N_4689,N_3336);
and U6017 (N_6017,N_3815,N_5582);
and U6018 (N_6018,N_4191,N_4789);
nor U6019 (N_6019,N_5037,N_5740);
nor U6020 (N_6020,N_3187,N_3603);
xnor U6021 (N_6021,N_5927,N_4141);
or U6022 (N_6022,N_4560,N_5016);
xnor U6023 (N_6023,N_5159,N_3299);
xnor U6024 (N_6024,N_3433,N_5433);
nor U6025 (N_6025,N_5899,N_4883);
nand U6026 (N_6026,N_3553,N_3337);
or U6027 (N_6027,N_5798,N_4764);
xnor U6028 (N_6028,N_4851,N_3092);
xor U6029 (N_6029,N_4281,N_4748);
nor U6030 (N_6030,N_3848,N_4431);
nor U6031 (N_6031,N_5608,N_5650);
nand U6032 (N_6032,N_3794,N_4924);
or U6033 (N_6033,N_4276,N_4821);
and U6034 (N_6034,N_5204,N_4065);
nor U6035 (N_6035,N_4912,N_4763);
nand U6036 (N_6036,N_4036,N_4966);
or U6037 (N_6037,N_4765,N_5780);
xnor U6038 (N_6038,N_4363,N_3659);
and U6039 (N_6039,N_5555,N_3342);
nor U6040 (N_6040,N_5304,N_3766);
xnor U6041 (N_6041,N_3206,N_4578);
nor U6042 (N_6042,N_4867,N_4421);
or U6043 (N_6043,N_4980,N_4156);
xor U6044 (N_6044,N_4109,N_3960);
nand U6045 (N_6045,N_4270,N_5799);
xor U6046 (N_6046,N_5332,N_4770);
nor U6047 (N_6047,N_3096,N_5420);
nand U6048 (N_6048,N_3690,N_5535);
nor U6049 (N_6049,N_3721,N_4467);
nor U6050 (N_6050,N_3512,N_5826);
xor U6051 (N_6051,N_3945,N_3437);
nand U6052 (N_6052,N_4468,N_5196);
and U6053 (N_6053,N_5586,N_3630);
xnor U6054 (N_6054,N_3606,N_3104);
nor U6055 (N_6055,N_5371,N_3385);
nor U6056 (N_6056,N_5096,N_5794);
nor U6057 (N_6057,N_4498,N_4871);
nor U6058 (N_6058,N_4197,N_3199);
and U6059 (N_6059,N_5845,N_3073);
and U6060 (N_6060,N_5522,N_4564);
or U6061 (N_6061,N_4427,N_4027);
and U6062 (N_6062,N_3389,N_4370);
xnor U6063 (N_6063,N_3579,N_4590);
nand U6064 (N_6064,N_5620,N_3856);
xnor U6065 (N_6065,N_4635,N_3773);
xor U6066 (N_6066,N_4339,N_5451);
or U6067 (N_6067,N_5083,N_3452);
or U6068 (N_6068,N_4486,N_5355);
nor U6069 (N_6069,N_5984,N_4664);
or U6070 (N_6070,N_4182,N_4799);
or U6071 (N_6071,N_4325,N_5807);
nor U6072 (N_6072,N_5413,N_5682);
or U6073 (N_6073,N_3418,N_4668);
or U6074 (N_6074,N_5047,N_4108);
xor U6075 (N_6075,N_5452,N_5442);
nor U6076 (N_6076,N_4541,N_5503);
xor U6077 (N_6077,N_3032,N_4020);
nor U6078 (N_6078,N_4682,N_4804);
xnor U6079 (N_6079,N_3338,N_5931);
or U6080 (N_6080,N_5365,N_5394);
or U6081 (N_6081,N_5026,N_3818);
or U6082 (N_6082,N_3154,N_4750);
xor U6083 (N_6083,N_5078,N_5817);
nand U6084 (N_6084,N_5696,N_3636);
nand U6085 (N_6085,N_5119,N_5932);
nor U6086 (N_6086,N_5590,N_3303);
or U6087 (N_6087,N_3965,N_3800);
nand U6088 (N_6088,N_4920,N_5943);
or U6089 (N_6089,N_3106,N_3666);
or U6090 (N_6090,N_3901,N_3069);
nand U6091 (N_6091,N_3001,N_3130);
xnor U6092 (N_6092,N_5004,N_4003);
nor U6093 (N_6093,N_4524,N_4934);
xor U6094 (N_6094,N_5157,N_3870);
and U6095 (N_6095,N_4698,N_4674);
and U6096 (N_6096,N_4795,N_5972);
or U6097 (N_6097,N_3396,N_5208);
and U6098 (N_6098,N_5066,N_3862);
nor U6099 (N_6099,N_4387,N_4093);
and U6100 (N_6100,N_4885,N_5360);
nor U6101 (N_6101,N_5444,N_3838);
nand U6102 (N_6102,N_5864,N_5021);
and U6103 (N_6103,N_5154,N_3267);
nand U6104 (N_6104,N_3033,N_3426);
xor U6105 (N_6105,N_3458,N_3384);
xnor U6106 (N_6106,N_5253,N_5954);
and U6107 (N_6107,N_3562,N_5112);
and U6108 (N_6108,N_3400,N_3688);
nand U6109 (N_6109,N_3621,N_4522);
nor U6110 (N_6110,N_4017,N_3607);
xor U6111 (N_6111,N_3289,N_5121);
nor U6112 (N_6112,N_3691,N_3209);
and U6113 (N_6113,N_3140,N_4619);
and U6114 (N_6114,N_5041,N_5431);
or U6115 (N_6115,N_5426,N_3467);
nand U6116 (N_6116,N_4814,N_3242);
xor U6117 (N_6117,N_5067,N_5500);
nor U6118 (N_6118,N_3778,N_3518);
xnor U6119 (N_6119,N_5311,N_4329);
and U6120 (N_6120,N_5013,N_5249);
nor U6121 (N_6121,N_3550,N_3834);
or U6122 (N_6122,N_3872,N_4807);
nand U6123 (N_6123,N_4075,N_5569);
and U6124 (N_6124,N_4741,N_3596);
xnor U6125 (N_6125,N_5028,N_5467);
nand U6126 (N_6126,N_3932,N_4260);
and U6127 (N_6127,N_4049,N_3650);
or U6128 (N_6128,N_4350,N_4353);
xnor U6129 (N_6129,N_5147,N_3668);
nor U6130 (N_6130,N_4235,N_4459);
nor U6131 (N_6131,N_4263,N_4729);
nand U6132 (N_6132,N_4756,N_3419);
xor U6133 (N_6133,N_5510,N_4837);
xnor U6134 (N_6134,N_4688,N_3733);
and U6135 (N_6135,N_5161,N_4731);
nor U6136 (N_6136,N_3064,N_5215);
or U6137 (N_6137,N_4480,N_4212);
or U6138 (N_6138,N_3495,N_5148);
and U6139 (N_6139,N_4220,N_3785);
and U6140 (N_6140,N_5802,N_3328);
nand U6141 (N_6141,N_4011,N_5629);
xnor U6142 (N_6142,N_3016,N_5448);
and U6143 (N_6143,N_5070,N_4818);
nand U6144 (N_6144,N_3178,N_3643);
and U6145 (N_6145,N_4057,N_4357);
or U6146 (N_6146,N_4776,N_3448);
xor U6147 (N_6147,N_4061,N_3849);
xor U6148 (N_6148,N_5377,N_5344);
nand U6149 (N_6149,N_3955,N_5842);
and U6150 (N_6150,N_3174,N_5949);
or U6151 (N_6151,N_3601,N_4392);
nor U6152 (N_6152,N_3158,N_5293);
and U6153 (N_6153,N_3594,N_4405);
and U6154 (N_6154,N_3739,N_4097);
and U6155 (N_6155,N_3922,N_5662);
nand U6156 (N_6156,N_5717,N_5664);
xor U6157 (N_6157,N_5468,N_4333);
and U6158 (N_6158,N_5481,N_4830);
and U6159 (N_6159,N_3217,N_4058);
xnor U6160 (N_6160,N_4247,N_3115);
and U6161 (N_6161,N_5556,N_4323);
nand U6162 (N_6162,N_4110,N_4437);
nand U6163 (N_6163,N_3205,N_4589);
nand U6164 (N_6164,N_5553,N_3625);
nor U6165 (N_6165,N_3789,N_4724);
and U6166 (N_6166,N_4899,N_4308);
nand U6167 (N_6167,N_3368,N_4418);
nand U6168 (N_6168,N_3142,N_4569);
and U6169 (N_6169,N_4793,N_4375);
or U6170 (N_6170,N_3908,N_4155);
nand U6171 (N_6171,N_5554,N_4746);
nor U6172 (N_6172,N_4879,N_4643);
or U6173 (N_6173,N_4391,N_5635);
and U6174 (N_6174,N_4131,N_4219);
xor U6175 (N_6175,N_4164,N_4601);
or U6176 (N_6176,N_4424,N_5750);
xnor U6177 (N_6177,N_4877,N_3191);
nor U6178 (N_6178,N_4379,N_5689);
xor U6179 (N_6179,N_4300,N_5808);
xnor U6180 (N_6180,N_4021,N_5517);
nor U6181 (N_6181,N_5713,N_5513);
xnor U6182 (N_6182,N_3276,N_5795);
nand U6183 (N_6183,N_5001,N_5505);
nor U6184 (N_6184,N_5823,N_5552);
nand U6185 (N_6185,N_4287,N_5834);
and U6186 (N_6186,N_3207,N_3624);
or U6187 (N_6187,N_3160,N_4126);
xnor U6188 (N_6188,N_4827,N_4211);
xor U6189 (N_6189,N_5474,N_4785);
nand U6190 (N_6190,N_5109,N_5429);
nand U6191 (N_6191,N_3439,N_3372);
and U6192 (N_6192,N_5188,N_5372);
nand U6193 (N_6193,N_5130,N_4367);
nor U6194 (N_6194,N_5787,N_5090);
nand U6195 (N_6195,N_4996,N_5935);
or U6196 (N_6196,N_3176,N_5829);
xor U6197 (N_6197,N_4646,N_4332);
and U6198 (N_6198,N_5461,N_4727);
nand U6199 (N_6199,N_3296,N_4227);
and U6200 (N_6200,N_5515,N_3044);
xor U6201 (N_6201,N_3480,N_4628);
nand U6202 (N_6202,N_4918,N_5348);
nand U6203 (N_6203,N_5407,N_4185);
or U6204 (N_6204,N_3939,N_5134);
nor U6205 (N_6205,N_3216,N_4404);
xnor U6206 (N_6206,N_3612,N_3376);
or U6207 (N_6207,N_4811,N_4758);
nor U6208 (N_6208,N_4695,N_5031);
and U6209 (N_6209,N_3557,N_5640);
nor U6210 (N_6210,N_3099,N_4686);
xnor U6211 (N_6211,N_5909,N_3737);
nand U6212 (N_6212,N_4351,N_4501);
xor U6213 (N_6213,N_3757,N_5368);
xnor U6214 (N_6214,N_4993,N_5987);
xnor U6215 (N_6215,N_5851,N_5404);
or U6216 (N_6216,N_5944,N_4342);
nand U6217 (N_6217,N_4166,N_4473);
nor U6218 (N_6218,N_3724,N_4624);
xnor U6219 (N_6219,N_5256,N_4816);
nor U6220 (N_6220,N_3846,N_3884);
or U6221 (N_6221,N_4749,N_4513);
and U6222 (N_6222,N_5310,N_5095);
nand U6223 (N_6223,N_3483,N_5173);
xnor U6224 (N_6224,N_4666,N_4389);
xor U6225 (N_6225,N_3473,N_5709);
nor U6226 (N_6226,N_3365,N_3608);
xor U6227 (N_6227,N_5698,N_5647);
xor U6228 (N_6228,N_3320,N_4396);
xnor U6229 (N_6229,N_4484,N_3532);
nor U6230 (N_6230,N_4687,N_5265);
nor U6231 (N_6231,N_5945,N_5369);
or U6232 (N_6232,N_4562,N_5989);
xnor U6233 (N_6233,N_4998,N_5006);
nor U6234 (N_6234,N_4834,N_5880);
xnor U6235 (N_6235,N_5122,N_5781);
xnor U6236 (N_6236,N_3037,N_5334);
xnor U6237 (N_6237,N_5184,N_3719);
nor U6238 (N_6238,N_4436,N_5558);
xnor U6239 (N_6239,N_5491,N_3683);
nand U6240 (N_6240,N_4496,N_3502);
and U6241 (N_6241,N_5030,N_5991);
nor U6242 (N_6242,N_4667,N_4990);
nor U6243 (N_6243,N_4554,N_5094);
nand U6244 (N_6244,N_3589,N_3215);
xnor U6245 (N_6245,N_3172,N_4923);
nand U6246 (N_6246,N_5570,N_3475);
nand U6247 (N_6247,N_4576,N_3904);
and U6248 (N_6248,N_3315,N_4095);
nand U6249 (N_6249,N_4665,N_5782);
xor U6250 (N_6250,N_4159,N_4302);
nor U6251 (N_6251,N_4237,N_4747);
and U6252 (N_6252,N_4754,N_3580);
nand U6253 (N_6253,N_3049,N_4435);
or U6254 (N_6254,N_3253,N_4451);
and U6255 (N_6255,N_3568,N_5020);
or U6256 (N_6256,N_3841,N_5349);
nor U6257 (N_6257,N_4937,N_3201);
nand U6258 (N_6258,N_3806,N_3722);
or U6259 (N_6259,N_4411,N_5146);
and U6260 (N_6260,N_5470,N_3959);
xor U6261 (N_6261,N_4605,N_3819);
xor U6262 (N_6262,N_5283,N_5193);
or U6263 (N_6263,N_4661,N_3428);
nand U6264 (N_6264,N_5600,N_5721);
or U6265 (N_6265,N_3648,N_5425);
nand U6266 (N_6266,N_3723,N_4177);
nand U6267 (N_6267,N_5391,N_4705);
nor U6268 (N_6268,N_4832,N_3449);
or U6269 (N_6269,N_5800,N_3551);
nor U6270 (N_6270,N_3190,N_5406);
xor U6271 (N_6271,N_5303,N_5353);
nor U6272 (N_6272,N_4419,N_3879);
and U6273 (N_6273,N_5496,N_5938);
nand U6274 (N_6274,N_3339,N_5035);
nand U6275 (N_6275,N_5018,N_3358);
nor U6276 (N_6276,N_3827,N_5596);
xnor U6277 (N_6277,N_3656,N_4654);
nand U6278 (N_6278,N_3516,N_4847);
and U6279 (N_6279,N_5678,N_3117);
and U6280 (N_6280,N_3796,N_3335);
nand U6281 (N_6281,N_4297,N_3671);
nor U6282 (N_6282,N_5207,N_3219);
or U6283 (N_6283,N_3284,N_3229);
nor U6284 (N_6284,N_5317,N_5174);
nand U6285 (N_6285,N_5409,N_5463);
or U6286 (N_6286,N_4952,N_3103);
nor U6287 (N_6287,N_3503,N_5988);
nand U6288 (N_6288,N_5063,N_5268);
xnor U6289 (N_6289,N_3768,N_3052);
or U6290 (N_6290,N_5271,N_5234);
nand U6291 (N_6291,N_5309,N_5040);
and U6292 (N_6292,N_3405,N_4153);
or U6293 (N_6293,N_3735,N_5730);
and U6294 (N_6294,N_5354,N_3840);
and U6295 (N_6295,N_5770,N_4478);
and U6296 (N_6296,N_5551,N_4091);
xnor U6297 (N_6297,N_5301,N_3062);
xnor U6298 (N_6298,N_5290,N_5612);
nand U6299 (N_6299,N_5755,N_4213);
xnor U6300 (N_6300,N_4571,N_4417);
or U6301 (N_6301,N_5285,N_5670);
nor U6302 (N_6302,N_4259,N_4098);
xor U6303 (N_6303,N_3005,N_5076);
nor U6304 (N_6304,N_4870,N_3110);
nand U6305 (N_6305,N_3708,N_3598);
nor U6306 (N_6306,N_3414,N_3902);
and U6307 (N_6307,N_3756,N_4981);
xor U6308 (N_6308,N_5905,N_5761);
xor U6309 (N_6309,N_4113,N_5904);
nor U6310 (N_6310,N_3639,N_5350);
and U6311 (N_6311,N_5531,N_3009);
or U6312 (N_6312,N_3992,N_5925);
nor U6313 (N_6313,N_3260,N_4187);
xor U6314 (N_6314,N_5424,N_3194);
nand U6315 (N_6315,N_3162,N_5875);
xnor U6316 (N_6316,N_5902,N_4111);
nand U6317 (N_6317,N_3318,N_4127);
or U6318 (N_6318,N_4640,N_3905);
or U6319 (N_6319,N_5549,N_5435);
and U6320 (N_6320,N_5291,N_5890);
nand U6321 (N_6321,N_3933,N_4780);
and U6322 (N_6322,N_4005,N_4439);
or U6323 (N_6323,N_3442,N_4454);
xor U6324 (N_6324,N_3541,N_4201);
or U6325 (N_6325,N_4248,N_4186);
and U6326 (N_6326,N_3181,N_4775);
and U6327 (N_6327,N_4502,N_3593);
nor U6328 (N_6328,N_5888,N_3821);
or U6329 (N_6329,N_3258,N_4519);
nand U6330 (N_6330,N_3151,N_3810);
xnor U6331 (N_6331,N_4778,N_3564);
or U6332 (N_6332,N_4495,N_4946);
xnor U6333 (N_6333,N_5710,N_3374);
or U6334 (N_6334,N_5366,N_3943);
nor U6335 (N_6335,N_3696,N_3015);
xnor U6336 (N_6336,N_3897,N_3007);
nor U6337 (N_6337,N_3295,N_4782);
or U6338 (N_6338,N_3802,N_3980);
nor U6339 (N_6339,N_3380,N_3168);
and U6340 (N_6340,N_5385,N_4253);
nor U6341 (N_6341,N_3710,N_3393);
or U6342 (N_6342,N_3245,N_3540);
nand U6343 (N_6343,N_5323,N_3399);
or U6344 (N_6344,N_5788,N_4528);
and U6345 (N_6345,N_3198,N_3997);
or U6346 (N_6346,N_5685,N_5158);
or U6347 (N_6347,N_3128,N_5477);
and U6348 (N_6348,N_4773,N_4986);
nor U6349 (N_6349,N_3978,N_3485);
and U6350 (N_6350,N_4526,N_4032);
and U6351 (N_6351,N_5509,N_3326);
nand U6352 (N_6352,N_3192,N_4004);
nand U6353 (N_6353,N_4115,N_4099);
nand U6354 (N_6354,N_3610,N_3252);
or U6355 (N_6355,N_5745,N_3985);
or U6356 (N_6356,N_4568,N_4898);
and U6357 (N_6357,N_3177,N_5928);
or U6358 (N_6358,N_5815,N_3213);
and U6359 (N_6359,N_3188,N_3238);
and U6360 (N_6360,N_4195,N_5053);
and U6361 (N_6361,N_5979,N_3514);
or U6362 (N_6362,N_4653,N_4888);
nand U6363 (N_6363,N_5728,N_5460);
and U6364 (N_6364,N_4139,N_5639);
xnor U6365 (N_6365,N_3930,N_5275);
or U6366 (N_6366,N_3774,N_4178);
nand U6367 (N_6367,N_5400,N_4401);
nor U6368 (N_6368,N_3169,N_5218);
and U6369 (N_6369,N_5908,N_4138);
and U6370 (N_6370,N_4050,N_3051);
nand U6371 (N_6371,N_5512,N_5055);
nor U6372 (N_6372,N_4073,N_4397);
nand U6373 (N_6373,N_5810,N_5277);
nand U6374 (N_6374,N_5432,N_4002);
nand U6375 (N_6375,N_4771,N_5912);
xnor U6376 (N_6376,N_3752,N_3196);
or U6377 (N_6377,N_3406,N_4380);
xnor U6378 (N_6378,N_4162,N_3411);
and U6379 (N_6379,N_4712,N_4107);
xnor U6380 (N_6380,N_5584,N_3956);
or U6381 (N_6381,N_4685,N_5965);
or U6382 (N_6382,N_5416,N_4823);
or U6383 (N_6383,N_4225,N_3011);
nand U6384 (N_6384,N_5466,N_5085);
and U6385 (N_6385,N_4916,N_3617);
and U6386 (N_6386,N_4149,N_5205);
nor U6387 (N_6387,N_3547,N_4266);
and U6388 (N_6388,N_4913,N_5648);
or U6389 (N_6389,N_4557,N_5926);
or U6390 (N_6390,N_3570,N_3434);
nor U6391 (N_6391,N_5162,N_4544);
xor U6392 (N_6392,N_3701,N_3695);
xnor U6393 (N_6393,N_3059,N_5669);
nor U6394 (N_6394,N_3046,N_5410);
xnor U6395 (N_6395,N_4381,N_4919);
and U6396 (N_6396,N_5417,N_4446);
nand U6397 (N_6397,N_3455,N_5191);
or U6398 (N_6398,N_5897,N_3272);
and U6399 (N_6399,N_5024,N_4445);
and U6400 (N_6400,N_3446,N_5089);
or U6401 (N_6401,N_4040,N_3750);
or U6402 (N_6402,N_3298,N_4671);
and U6403 (N_6403,N_5540,N_4356);
nand U6404 (N_6404,N_3890,N_5626);
nor U6405 (N_6405,N_5748,N_4696);
or U6406 (N_6406,N_5005,N_5113);
or U6407 (N_6407,N_5797,N_3764);
nand U6408 (N_6408,N_4849,N_5386);
and U6409 (N_6409,N_5746,N_4080);
nor U6410 (N_6410,N_3889,N_3310);
or U6411 (N_6411,N_3432,N_4701);
nor U6412 (N_6412,N_3983,N_5610);
and U6413 (N_6413,N_4931,N_3039);
and U6414 (N_6414,N_3609,N_3864);
or U6415 (N_6415,N_5098,N_5950);
or U6416 (N_6416,N_5454,N_5176);
or U6417 (N_6417,N_4752,N_5217);
nor U6418 (N_6418,N_3835,N_5573);
nor U6419 (N_6419,N_3929,N_5325);
xor U6420 (N_6420,N_5257,N_3831);
nand U6421 (N_6421,N_4147,N_3792);
or U6422 (N_6422,N_4489,N_5796);
or U6423 (N_6423,N_5064,N_4124);
xor U6424 (N_6424,N_4079,N_5776);
and U6425 (N_6425,N_5525,N_4045);
xnor U6426 (N_6426,N_3599,N_3588);
and U6427 (N_6427,N_5264,N_5145);
nor U6428 (N_6428,N_4599,N_3071);
and U6429 (N_6429,N_5084,N_5223);
nor U6430 (N_6430,N_5869,N_3918);
xor U6431 (N_6431,N_3304,N_5895);
nand U6432 (N_6432,N_3105,N_5900);
nor U6433 (N_6433,N_5952,N_4796);
nand U6434 (N_6434,N_4648,N_5252);
or U6435 (N_6435,N_5266,N_4317);
nor U6436 (N_6436,N_3886,N_3692);
or U6437 (N_6437,N_3996,N_3012);
xor U6438 (N_6438,N_4670,N_5116);
and U6439 (N_6439,N_4878,N_4662);
nand U6440 (N_6440,N_3873,N_5998);
xor U6441 (N_6441,N_3543,N_5199);
nor U6442 (N_6442,N_3490,N_5069);
nand U6443 (N_6443,N_3984,N_3002);
xor U6444 (N_6444,N_3824,N_5248);
and U6445 (N_6445,N_3732,N_4230);
or U6446 (N_6446,N_4861,N_3133);
xnor U6447 (N_6447,N_3288,N_3409);
nand U6448 (N_6448,N_4615,N_3189);
or U6449 (N_6449,N_4609,N_3808);
or U6450 (N_6450,N_5544,N_5194);
and U6451 (N_6451,N_3534,N_3280);
and U6452 (N_6452,N_4290,N_5486);
xnor U6453 (N_6453,N_5080,N_5738);
nand U6454 (N_6454,N_5521,N_5251);
or U6455 (N_6455,N_4365,N_5446);
nor U6456 (N_6456,N_3447,N_3454);
or U6457 (N_6457,N_3424,N_5753);
and U6458 (N_6458,N_4518,N_4797);
or U6459 (N_6459,N_3210,N_3070);
or U6460 (N_6460,N_5818,N_4304);
and U6461 (N_6461,N_5907,N_5367);
xor U6462 (N_6462,N_4621,N_4344);
nor U6463 (N_6463,N_3363,N_3644);
nor U6464 (N_6464,N_5806,N_4769);
and U6465 (N_6465,N_3146,N_4450);
and U6466 (N_6466,N_4865,N_5627);
xor U6467 (N_6467,N_5281,N_4608);
nor U6468 (N_6468,N_3026,N_3567);
nand U6469 (N_6469,N_5092,N_4974);
nand U6470 (N_6470,N_5995,N_4134);
and U6471 (N_6471,N_5229,N_5307);
or U6472 (N_6472,N_3771,N_5767);
nand U6473 (N_6473,N_3672,N_5680);
and U6474 (N_6474,N_3573,N_4265);
and U6475 (N_6475,N_3687,N_3079);
nor U6476 (N_6476,N_4786,N_4140);
or U6477 (N_6477,N_5983,N_3173);
nor U6478 (N_6478,N_4105,N_4991);
nand U6479 (N_6479,N_4530,N_3472);
xnor U6480 (N_6480,N_4305,N_4409);
nor U6481 (N_6481,N_4638,N_5102);
xor U6482 (N_6482,N_5529,N_3973);
nor U6483 (N_6483,N_3230,N_4825);
and U6484 (N_6484,N_5338,N_4790);
or U6485 (N_6485,N_3751,N_4470);
xnor U6486 (N_6486,N_4887,N_5502);
or U6487 (N_6487,N_4517,N_5499);
nand U6488 (N_6488,N_4412,N_5288);
nor U6489 (N_6489,N_5674,N_4348);
nand U6490 (N_6490,N_5624,N_3144);
xnor U6491 (N_6491,N_4977,N_3231);
nand U6492 (N_6492,N_5032,N_3837);
and U6493 (N_6493,N_4965,N_3663);
or U6494 (N_6494,N_5528,N_4172);
or U6495 (N_6495,N_5661,N_5050);
nand U6496 (N_6496,N_5622,N_4456);
nand U6497 (N_6497,N_3065,N_3271);
nor U6498 (N_6498,N_4236,N_5286);
or U6499 (N_6499,N_3090,N_3379);
or U6500 (N_6500,N_3697,N_4700);
or U6501 (N_6501,N_5656,N_3050);
or U6502 (N_6502,N_4655,N_4895);
and U6503 (N_6503,N_4994,N_5560);
and U6504 (N_6504,N_4926,N_5472);
nand U6505 (N_6505,N_4369,N_5227);
or U6506 (N_6506,N_5246,N_3297);
xnor U6507 (N_6507,N_4941,N_5414);
nand U6508 (N_6508,N_3360,N_4836);
nand U6509 (N_6509,N_5884,N_5827);
nand U6510 (N_6510,N_3854,N_5343);
nand U6511 (N_6511,N_4360,N_4047);
nor U6512 (N_6512,N_4805,N_4945);
and U6513 (N_6513,N_3619,N_3102);
and U6514 (N_6514,N_3075,N_5445);
nand U6515 (N_6515,N_5120,N_4326);
xnor U6516 (N_6516,N_3239,N_5002);
nand U6517 (N_6517,N_4713,N_4892);
and U6518 (N_6518,N_5930,N_4692);
nand U6519 (N_6519,N_4168,N_5581);
nor U6520 (N_6520,N_5777,N_4269);
and U6521 (N_6521,N_4720,N_3072);
nand U6522 (N_6522,N_5592,N_4129);
and U6523 (N_6523,N_3963,N_4857);
nand U6524 (N_6524,N_3018,N_3505);
nor U6525 (N_6525,N_5376,N_5314);
and U6526 (N_6526,N_5219,N_4928);
nor U6527 (N_6527,N_4844,N_3497);
and U6528 (N_6528,N_3971,N_5003);
or U6529 (N_6529,N_3830,N_3370);
and U6530 (N_6530,N_3132,N_3909);
nand U6531 (N_6531,N_5398,N_5744);
and U6532 (N_6532,N_3208,N_4053);
xnor U6533 (N_6533,N_3127,N_5103);
nand U6534 (N_6534,N_3123,N_4715);
xnor U6535 (N_6535,N_3255,N_5480);
xor U6536 (N_6536,N_5572,N_3354);
nand U6537 (N_6537,N_5361,N_3839);
nor U6538 (N_6538,N_3633,N_5957);
xnor U6539 (N_6539,N_5720,N_5287);
nand U6540 (N_6540,N_4132,N_5599);
nor U6541 (N_6541,N_3008,N_3522);
or U6542 (N_6542,N_3163,N_4206);
and U6543 (N_6543,N_3262,N_4262);
nor U6544 (N_6544,N_4798,N_5563);
or U6545 (N_6545,N_3866,N_5847);
nor U6546 (N_6546,N_4971,N_3076);
and U6547 (N_6547,N_4901,N_4074);
and U6548 (N_6548,N_5866,N_3402);
xnor U6549 (N_6549,N_5898,N_5604);
nor U6550 (N_6550,N_3499,N_5852);
nor U6551 (N_6551,N_4322,N_5272);
or U6552 (N_6552,N_4534,N_5541);
xnor U6553 (N_6553,N_4022,N_5783);
and U6554 (N_6554,N_4420,N_3727);
nand U6555 (N_6555,N_5008,N_5437);
or U6556 (N_6556,N_3235,N_3887);
and U6557 (N_6557,N_3150,N_3894);
or U6558 (N_6558,N_3538,N_4398);
nor U6559 (N_6559,N_4846,N_3638);
xnor U6560 (N_6560,N_3627,N_3999);
and U6561 (N_6561,N_4694,N_5542);
nand U6562 (N_6562,N_3703,N_5319);
nand U6563 (N_6563,N_3082,N_4423);
and U6564 (N_6564,N_5862,N_3811);
or U6565 (N_6565,N_3595,N_5537);
or U6566 (N_6566,N_3138,N_4595);
xnor U6567 (N_6567,N_3647,N_4644);
nor U6568 (N_6568,N_4951,N_5792);
xnor U6569 (N_6569,N_3003,N_4603);
nand U6570 (N_6570,N_4160,N_5785);
and U6571 (N_6571,N_5059,N_5363);
and U6572 (N_6572,N_4866,N_4580);
and U6573 (N_6573,N_4154,N_5733);
nand U6574 (N_6574,N_3685,N_5881);
xor U6575 (N_6575,N_3022,N_3974);
xnor U6576 (N_6576,N_3741,N_3319);
and U6577 (N_6577,N_5007,N_5887);
or U6578 (N_6578,N_5603,N_4908);
or U6579 (N_6579,N_4531,N_4232);
or U6580 (N_6580,N_5142,N_5643);
and U6581 (N_6581,N_4552,N_3545);
or U6582 (N_6582,N_3078,N_3620);
xnor U6583 (N_6583,N_4399,N_4018);
nand U6584 (N_6584,N_3249,N_4950);
and U6585 (N_6585,N_4516,N_3184);
nand U6586 (N_6586,N_4960,N_3662);
nor U6587 (N_6587,N_4649,N_4944);
nand U6588 (N_6588,N_3883,N_4347);
xnor U6589 (N_6589,N_5953,N_5330);
nor U6590 (N_6590,N_3250,N_5816);
and U6591 (N_6591,N_3118,N_5835);
nor U6592 (N_6592,N_3674,N_4947);
nand U6593 (N_6593,N_5380,N_5663);
or U6594 (N_6594,N_4082,N_4463);
or U6595 (N_6595,N_5919,N_4550);
nand U6596 (N_6596,N_3544,N_3845);
nor U6597 (N_6597,N_5846,N_3738);
and U6598 (N_6598,N_5789,N_5981);
nand U6599 (N_6599,N_5975,N_5729);
nand U6600 (N_6600,N_3470,N_5839);
or U6601 (N_6601,N_3730,N_4485);
nor U6602 (N_6602,N_4476,N_3256);
or U6603 (N_6603,N_4567,N_5786);
or U6604 (N_6604,N_4242,N_3097);
nor U6605 (N_6605,N_3582,N_4511);
nand U6606 (N_6606,N_5676,N_4469);
nor U6607 (N_6607,N_5168,N_4313);
xnor U6608 (N_6608,N_4432,N_5045);
or U6609 (N_6609,N_3847,N_3420);
nor U6610 (N_6610,N_5861,N_4210);
xor U6611 (N_6611,N_3585,N_5688);
and U6612 (N_6612,N_4874,N_4940);
or U6613 (N_6613,N_5236,N_3681);
nor U6614 (N_6614,N_4540,N_3031);
and U6615 (N_6615,N_4383,N_3976);
xnor U6616 (N_6616,N_5300,N_4145);
xnor U6617 (N_6617,N_5014,N_4964);
and U6618 (N_6618,N_3491,N_5044);
nor U6619 (N_6619,N_4779,N_5160);
nand U6620 (N_6620,N_5614,N_3006);
or U6621 (N_6621,N_3836,N_3471);
nand U6622 (N_6622,N_4483,N_5595);
or U6623 (N_6623,N_5660,N_3356);
nor U6624 (N_6624,N_3248,N_3654);
nand U6625 (N_6625,N_5634,N_4092);
and U6626 (N_6626,N_4613,N_4566);
nand U6627 (N_6627,N_3226,N_3350);
or U6628 (N_6628,N_5779,N_5822);
or U6629 (N_6629,N_5126,N_4295);
or U6630 (N_6630,N_3042,N_3972);
or U6631 (N_6631,N_3227,N_4106);
nand U6632 (N_6632,N_5172,N_5628);
xor U6633 (N_6633,N_4767,N_3548);
nand U6634 (N_6634,N_3660,N_4725);
xor U6635 (N_6635,N_3359,N_3019);
nor U6636 (N_6636,N_3149,N_5993);
xor U6637 (N_6637,N_3587,N_4774);
nor U6638 (N_6638,N_3391,N_4772);
and U6639 (N_6639,N_4673,N_3048);
or U6640 (N_6640,N_5255,N_5233);
and U6641 (N_6641,N_3709,N_5370);
xor U6642 (N_6642,N_3367,N_4975);
or U6643 (N_6643,N_4978,N_3694);
or U6644 (N_6644,N_5469,N_4007);
nor U6645 (N_6645,N_5418,N_4890);
and U6646 (N_6646,N_3726,N_5894);
xor U6647 (N_6647,N_4925,N_3101);
nand U6648 (N_6648,N_4294,N_5872);
nor U6649 (N_6649,N_3241,N_5732);
and U6650 (N_6650,N_5388,N_3425);
and U6651 (N_6651,N_4144,N_4592);
nand U6652 (N_6652,N_4548,N_3852);
or U6653 (N_6653,N_3917,N_4598);
and U6654 (N_6654,N_5478,N_5479);
or U6655 (N_6655,N_3124,N_4216);
xor U6656 (N_6656,N_4240,N_5038);
and U6657 (N_6657,N_5011,N_5495);
or U6658 (N_6658,N_3094,N_3493);
or U6659 (N_6659,N_4198,N_4553);
xor U6660 (N_6660,N_5153,N_5315);
and U6661 (N_6661,N_5805,N_5985);
or U6662 (N_6662,N_5775,N_5606);
and U6663 (N_6663,N_3961,N_5440);
or U6664 (N_6664,N_5830,N_4067);
nor U6665 (N_6665,N_3832,N_5657);
and U6666 (N_6666,N_3185,N_5803);
nand U6667 (N_6667,N_3334,N_4320);
nor U6668 (N_6668,N_4193,N_4634);
and U6669 (N_6669,N_5850,N_5118);
xor U6670 (N_6670,N_3640,N_5441);
or U6671 (N_6671,N_3622,N_5029);
and U6672 (N_6672,N_3004,N_5675);
or U6673 (N_6673,N_4133,N_4037);
and U6674 (N_6674,N_3237,N_3556);
nand U6675 (N_6675,N_4374,N_3055);
or U6676 (N_6676,N_4026,N_5642);
and U6677 (N_6677,N_3618,N_3398);
nand U6678 (N_6678,N_5757,N_5773);
and U6679 (N_6679,N_5258,N_4708);
or U6680 (N_6680,N_3408,N_3182);
nand U6681 (N_6681,N_5390,N_5838);
and U6682 (N_6682,N_3829,N_5532);
xor U6683 (N_6683,N_4217,N_4508);
and U6684 (N_6684,N_5986,N_3317);
and U6685 (N_6685,N_5690,N_5771);
nand U6686 (N_6686,N_5763,N_4481);
nand U6687 (N_6687,N_3364,N_4403);
or U6688 (N_6688,N_5228,N_3214);
xnor U6689 (N_6689,N_5171,N_3068);
and U6690 (N_6690,N_5305,N_5976);
xor U6691 (N_6691,N_4428,N_3027);
and U6692 (N_6692,N_4330,N_3958);
nor U6693 (N_6693,N_4479,N_5978);
or U6694 (N_6694,N_4104,N_3487);
xnor U6695 (N_6695,N_5279,N_3159);
nand U6696 (N_6696,N_5086,N_3628);
nand U6697 (N_6697,N_5071,N_3665);
xor U6698 (N_6698,N_3651,N_3949);
or U6699 (N_6699,N_3330,N_4303);
and U6700 (N_6700,N_4868,N_3047);
xor U6701 (N_6701,N_4917,N_5187);
nor U6702 (N_6702,N_3197,N_5566);
nor U6703 (N_6703,N_3488,N_3855);
nor U6704 (N_6704,N_5179,N_3913);
or U6705 (N_6705,N_3179,N_3085);
and U6706 (N_6706,N_3584,N_4954);
xor U6707 (N_6707,N_5828,N_3028);
nor U6708 (N_6708,N_4135,N_5523);
xor U6709 (N_6709,N_5762,N_4228);
and U6710 (N_6710,N_3698,N_3747);
or U6711 (N_6711,N_5088,N_5632);
nand U6712 (N_6712,N_4028,N_3634);
and U6713 (N_6713,N_4448,N_5557);
nor U6714 (N_6714,N_4963,N_5097);
nor U6715 (N_6715,N_4334,N_3803);
or U6716 (N_6716,N_4143,N_3469);
nand U6717 (N_6717,N_4354,N_5677);
or U6718 (N_6718,N_4167,N_3378);
or U6719 (N_6719,N_5170,N_4038);
xnor U6720 (N_6720,N_3860,N_4543);
nand U6721 (N_6721,N_3677,N_5585);
xor U6722 (N_6722,N_3083,N_4051);
nand U6723 (N_6723,N_5920,N_3161);
and U6724 (N_6724,N_3931,N_4475);
or U6725 (N_6725,N_3034,N_5222);
xor U6726 (N_6726,N_5081,N_3842);
nand U6727 (N_6727,N_5843,N_5804);
and U6728 (N_6728,N_5963,N_3877);
xnor U6729 (N_6729,N_4062,N_3035);
nand U6730 (N_6730,N_3798,N_5449);
and U6731 (N_6731,N_5213,N_4284);
xnor U6732 (N_6732,N_4070,N_4364);
nand U6733 (N_6733,N_5743,N_5110);
nand U6734 (N_6734,N_4386,N_4324);
xor U6735 (N_6735,N_3928,N_4393);
or U6736 (N_6736,N_5623,N_5646);
or U6737 (N_6737,N_4985,N_3575);
and U6738 (N_6738,N_5588,N_4999);
nor U6739 (N_6739,N_5243,N_5747);
nor U6740 (N_6740,N_5752,N_5793);
or U6741 (N_6741,N_5383,N_3987);
or U6742 (N_6742,N_4792,N_5577);
nand U6743 (N_6743,N_4610,N_3331);
xor U6744 (N_6744,N_3729,N_5242);
and U6745 (N_6745,N_5093,N_5990);
nor U6746 (N_6746,N_3944,N_5575);
xnor U6747 (N_6747,N_4581,N_4939);
nor U6748 (N_6748,N_4681,N_5699);
nand U6749 (N_6749,N_5231,N_3228);
xnor U6750 (N_6750,N_3220,N_4542);
xnor U6751 (N_6751,N_3581,N_3371);
nand U6752 (N_6752,N_3463,N_4535);
nor U6753 (N_6753,N_3074,N_4340);
nor U6754 (N_6754,N_5206,N_5117);
or U6755 (N_6755,N_5051,N_5289);
nand U6756 (N_6756,N_4622,N_5630);
or U6757 (N_6757,N_4935,N_4068);
and U6758 (N_6758,N_4152,N_5333);
nor U6759 (N_6759,N_3950,N_4848);
and U6760 (N_6760,N_4440,N_3134);
xnor U6761 (N_6761,N_4251,N_5061);
and U6762 (N_6762,N_5882,N_4967);
nor U6763 (N_6763,N_3868,N_4791);
or U6764 (N_6764,N_4243,N_3693);
xnor U6765 (N_6765,N_4717,N_5597);
xnor U6766 (N_6766,N_5924,N_5389);
nand U6767 (N_6767,N_4315,N_4137);
xor U6768 (N_6768,N_4781,N_5401);
nor U6769 (N_6769,N_4229,N_4088);
and U6770 (N_6770,N_3014,N_4096);
xor U6771 (N_6771,N_5631,N_3707);
or U6772 (N_6772,N_5649,N_5378);
and U6773 (N_6773,N_3574,N_3308);
nor U6774 (N_6774,N_4310,N_5459);
or U6775 (N_6775,N_4840,N_3896);
or U6776 (N_6776,N_4632,N_3743);
nor U6777 (N_6777,N_3565,N_5959);
nor U6778 (N_6778,N_4740,N_3443);
nand U6779 (N_6779,N_4161,N_3940);
xor U6780 (N_6780,N_5561,N_3533);
xor U6781 (N_6781,N_3116,N_4490);
or U6782 (N_6782,N_4884,N_4757);
and U6783 (N_6783,N_4094,N_3347);
and U6784 (N_6784,N_4721,N_5520);
or U6785 (N_6785,N_3286,N_3770);
or U6786 (N_6786,N_5106,N_3948);
xor U6787 (N_6787,N_4184,N_5210);
nor U6788 (N_6788,N_4845,N_5621);
or U6789 (N_6789,N_5443,N_5356);
and U6790 (N_6790,N_5605,N_3966);
nand U6791 (N_6791,N_4255,N_5485);
xnor U6792 (N_6792,N_4669,N_4071);
nand U6793 (N_6793,N_3285,N_4841);
and U6794 (N_6794,N_4171,N_5591);
and U6795 (N_6795,N_4142,N_5465);
nor U6796 (N_6796,N_3641,N_4100);
or U6797 (N_6797,N_4116,N_3119);
nor U6798 (N_6798,N_4711,N_3462);
or U6799 (N_6799,N_3925,N_5175);
or U6800 (N_6800,N_4222,N_4869);
xnor U6801 (N_6801,N_4415,N_3592);
xnor U6802 (N_6802,N_3791,N_3273);
xnor U6803 (N_6803,N_5273,N_3456);
nor U6804 (N_6804,N_5964,N_3281);
xor U6805 (N_6805,N_5751,N_3761);
and U6806 (N_6806,N_5711,N_5999);
and U6807 (N_6807,N_5704,N_5982);
xor U6808 (N_6808,N_4000,N_3436);
or U6809 (N_6809,N_3322,N_5165);
or U6810 (N_6810,N_4810,N_5824);
nand U6811 (N_6811,N_3947,N_5203);
and U6812 (N_6812,N_3468,N_5896);
xnor U6813 (N_6813,N_3613,N_4559);
xor U6814 (N_6814,N_5671,N_3404);
xnor U6815 (N_6815,N_4812,N_4044);
and U6816 (N_6816,N_3713,N_3851);
nor U6817 (N_6817,N_4413,N_5419);
xnor U6818 (N_6818,N_3478,N_5618);
nand U6819 (N_6819,N_4549,N_3136);
xnor U6820 (N_6820,N_5961,N_4956);
nor U6821 (N_6821,N_5225,N_4600);
or U6822 (N_6822,N_3711,N_3900);
or U6823 (N_6823,N_5316,N_3871);
nand U6824 (N_6824,N_4642,N_4808);
or U6825 (N_6825,N_3427,N_3125);
or U6826 (N_6826,N_4394,N_3646);
nand U6827 (N_6827,N_5655,N_3091);
and U6828 (N_6828,N_5833,N_3734);
or U6829 (N_6829,N_5966,N_4352);
and U6830 (N_6830,N_5854,N_5318);
nand U6831 (N_6831,N_3387,N_3680);
and U6832 (N_6832,N_5321,N_5455);
xnor U6833 (N_6833,N_4267,N_5166);
xnor U6834 (N_6834,N_3989,N_5209);
nor U6835 (N_6835,N_4165,N_5673);
nor U6836 (N_6836,N_4979,N_4819);
xnor U6837 (N_6837,N_5903,N_5644);
xor U6838 (N_6838,N_5259,N_5942);
nor U6839 (N_6839,N_3982,N_5428);
nor U6840 (N_6840,N_3498,N_5705);
or U6841 (N_6841,N_4783,N_5458);
and U6842 (N_6842,N_4982,N_4244);
nor U6843 (N_6843,N_5579,N_3290);
nand U6844 (N_6844,N_3885,N_4761);
or U6845 (N_6845,N_4278,N_4932);
nor U6846 (N_6846,N_3788,N_4146);
nor U6847 (N_6847,N_5156,N_5539);
and U6848 (N_6848,N_3998,N_5269);
xnor U6849 (N_6849,N_5619,N_3535);
and U6850 (N_6850,N_4472,N_4361);
xor U6851 (N_6851,N_5589,N_5077);
or U6852 (N_6852,N_5115,N_4449);
xor U6853 (N_6853,N_4922,N_4123);
nand U6854 (N_6854,N_5832,N_3193);
nor U6855 (N_6855,N_4112,N_5347);
or U6856 (N_6856,N_5123,N_3496);
xnor U6857 (N_6857,N_3268,N_3429);
or U6858 (N_6858,N_5237,N_4637);
nor U6859 (N_6859,N_4042,N_4988);
nor U6860 (N_6860,N_5504,N_4730);
and U6861 (N_6861,N_4886,N_5128);
nand U6862 (N_6862,N_5186,N_3807);
or U6863 (N_6863,N_5494,N_3500);
and U6864 (N_6864,N_5087,N_4509);
xor U6865 (N_6865,N_4272,N_4471);
and U6866 (N_6866,N_3484,N_4506);
nor U6867 (N_6867,N_5645,N_4938);
and U6868 (N_6868,N_5278,N_4118);
nor U6869 (N_6869,N_4008,N_3403);
nor U6870 (N_6870,N_3525,N_5214);
xnor U6871 (N_6871,N_4366,N_4572);
nor U6872 (N_6872,N_5543,N_5860);
nor U6873 (N_6873,N_4343,N_4130);
nand U6874 (N_6874,N_3390,N_4824);
xnor U6875 (N_6875,N_3345,N_4030);
xor U6876 (N_6876,N_4525,N_3444);
xnor U6877 (N_6877,N_4076,N_3355);
nor U6878 (N_6878,N_5450,N_3962);
or U6879 (N_6879,N_3968,N_3569);
xor U6880 (N_6880,N_4202,N_4829);
and U6881 (N_6881,N_3919,N_3912);
xor U6882 (N_6882,N_3431,N_3899);
nand U6883 (N_6883,N_5958,N_3563);
nand U6884 (N_6884,N_3986,N_3137);
and U6885 (N_6885,N_4959,N_4349);
and U6886 (N_6886,N_4537,N_4894);
nor U6887 (N_6887,N_5402,N_4151);
or U6888 (N_6888,N_3520,N_3517);
and U6889 (N_6889,N_3111,N_4809);
or U6890 (N_6890,N_4009,N_5488);
or U6891 (N_6891,N_4577,N_5056);
xor U6892 (N_6892,N_4574,N_3513);
nand U6893 (N_6893,N_5507,N_4529);
or U6894 (N_6894,N_3718,N_5346);
nand U6895 (N_6895,N_4400,N_4046);
and U6896 (N_6896,N_5107,N_5980);
nand U6897 (N_6897,N_4555,N_3795);
and U6898 (N_6898,N_3875,N_5867);
and U6899 (N_6899,N_5012,N_4903);
xnor U6900 (N_6900,N_4016,N_3170);
or U6901 (N_6901,N_5326,N_3141);
xnor U6902 (N_6902,N_5082,N_5731);
nand U6903 (N_6903,N_4858,N_3357);
and U6904 (N_6904,N_3853,N_3352);
or U6905 (N_6905,N_3951,N_4072);
and U6906 (N_6906,N_5396,N_3509);
nand U6907 (N_6907,N_3464,N_5167);
nor U6908 (N_6908,N_3820,N_3508);
or U6909 (N_6909,N_5100,N_5819);
xor U6910 (N_6910,N_5941,N_3775);
nand U6911 (N_6911,N_5534,N_4128);
xor U6912 (N_6912,N_4189,N_5801);
and U6913 (N_6913,N_3977,N_4914);
and U6914 (N_6914,N_4385,N_3457);
nor U6915 (N_6915,N_4538,N_4558);
or U6916 (N_6916,N_3486,N_5456);
or U6917 (N_6917,N_3812,N_5735);
nand U6918 (N_6918,N_5482,N_4921);
nor U6919 (N_6919,N_5034,N_5967);
and U6920 (N_6920,N_3926,N_5345);
nor U6921 (N_6921,N_5422,N_3546);
nand U6922 (N_6922,N_4274,N_4943);
and U6923 (N_6923,N_4103,N_4461);
xor U6924 (N_6924,N_5393,N_5879);
nand U6925 (N_6925,N_5739,N_4170);
xor U6926 (N_6926,N_5889,N_5436);
nor U6927 (N_6927,N_3952,N_3941);
nor U6928 (N_6928,N_5150,N_3279);
or U6929 (N_6929,N_4205,N_5598);
and U6930 (N_6930,N_3777,N_5855);
nand U6931 (N_6931,N_5727,N_3523);
xnor U6932 (N_6932,N_4289,N_4657);
xor U6933 (N_6933,N_5033,N_3754);
xor U6934 (N_6934,N_3725,N_4672);
and U6935 (N_6935,N_5140,N_4196);
nand U6936 (N_6936,N_3257,N_4784);
nand U6937 (N_6937,N_5977,N_5741);
xnor U6938 (N_6938,N_4716,N_5151);
xor U6939 (N_6939,N_4208,N_3131);
xnor U6940 (N_6940,N_5364,N_3611);
and U6941 (N_6941,N_3501,N_3301);
xor U6942 (N_6942,N_3164,N_4194);
and U6943 (N_6943,N_4880,N_5858);
nor U6944 (N_6944,N_3882,N_5929);
and U6945 (N_6945,N_5742,N_4234);
xor U6946 (N_6946,N_3657,N_4286);
or U6947 (N_6947,N_5381,N_4697);
xnor U6948 (N_6948,N_3410,N_5820);
or U6949 (N_6949,N_4579,N_3053);
nand U6950 (N_6950,N_5636,N_4355);
nand U6951 (N_6951,N_4444,N_5571);
nand U6952 (N_6952,N_4906,N_3474);
xor U6953 (N_6953,N_5357,N_4718);
and U6954 (N_6954,N_3935,N_3043);
nor U6955 (N_6955,N_3669,N_3597);
nor U6956 (N_6956,N_4794,N_5715);
nand U6957 (N_6957,N_4709,N_5439);
nand U6958 (N_6958,N_5892,N_4710);
and U6959 (N_6959,N_4684,N_3504);
nor U6960 (N_6960,N_5758,N_4318);
xor U6961 (N_6961,N_5601,N_4086);
nor U6962 (N_6962,N_5877,N_4390);
or U6963 (N_6963,N_3616,N_4972);
nand U6964 (N_6964,N_3045,N_4745);
nand U6965 (N_6965,N_3843,N_3507);
nand U6966 (N_6966,N_4545,N_4173);
nor U6967 (N_6967,N_5791,N_5638);
and U6968 (N_6968,N_3246,N_5760);
or U6969 (N_6969,N_3080,N_5497);
xor U6970 (N_6970,N_4034,N_3994);
or U6971 (N_6971,N_4504,N_4588);
xor U6972 (N_6972,N_3305,N_5239);
or U6973 (N_6973,N_3089,N_3302);
and U6974 (N_6974,N_4677,N_5423);
xor U6975 (N_6975,N_5901,N_3635);
xnor U6976 (N_6976,N_4815,N_3086);
or U6977 (N_6977,N_4268,N_3183);
or U6978 (N_6978,N_4551,N_4025);
nor U6979 (N_6979,N_3270,N_3706);
and U6980 (N_6980,N_4382,N_5133);
or U6981 (N_6981,N_3081,N_3526);
xor U6982 (N_6982,N_3122,N_5853);
nand U6983 (N_6983,N_5250,N_5493);
and U6984 (N_6984,N_5282,N_4407);
xnor U6985 (N_6985,N_3529,N_5637);
nor U6986 (N_6986,N_3343,N_5384);
or U6987 (N_6987,N_4203,N_3023);
or U6988 (N_6988,N_4371,N_5152);
nand U6989 (N_6989,N_4618,N_4059);
xnor U6990 (N_6990,N_3388,N_5968);
nand U6991 (N_6991,N_5609,N_5594);
or U6992 (N_6992,N_5336,N_4043);
nor U6993 (N_6993,N_5292,N_3717);
xnor U6994 (N_6994,N_3736,N_4188);
and U6995 (N_6995,N_5136,N_4199);
nor U6996 (N_6996,N_5939,N_5593);
or U6997 (N_6997,N_4491,N_3519);
nand U6998 (N_6998,N_3275,N_3967);
and U6999 (N_6999,N_3898,N_5578);
xor U7000 (N_7000,N_4341,N_3938);
nand U7001 (N_7001,N_4575,N_5238);
or U7002 (N_7002,N_4948,N_3934);
nand U7003 (N_7003,N_5178,N_4973);
or U7004 (N_7004,N_4447,N_3763);
or U7005 (N_7005,N_3661,N_3891);
xnor U7006 (N_7006,N_3600,N_3783);
and U7007 (N_7007,N_4582,N_4054);
and U7008 (N_7008,N_5049,N_5408);
and U7009 (N_7009,N_4293,N_3166);
nand U7010 (N_7010,N_5790,N_4862);
xor U7011 (N_7011,N_3038,N_3605);
and U7012 (N_7012,N_4298,N_4855);
nand U7013 (N_7013,N_3521,N_4744);
xor U7014 (N_7014,N_4319,N_3591);
nand U7015 (N_7015,N_3740,N_4233);
or U7016 (N_7016,N_5224,N_5580);
or U7017 (N_7017,N_5036,N_5778);
nor U7018 (N_7018,N_4378,N_4826);
nand U7019 (N_7019,N_4055,N_4680);
xnor U7020 (N_7020,N_5057,N_4828);
nand U7021 (N_7021,N_5043,N_3058);
nand U7022 (N_7022,N_3292,N_3892);
nor U7023 (N_7023,N_3844,N_5857);
or U7024 (N_7024,N_4547,N_5473);
xor U7025 (N_7025,N_3155,N_5765);
nand U7026 (N_7026,N_4949,N_4961);
nor U7027 (N_7027,N_4282,N_3095);
nand U7028 (N_7028,N_5583,N_5104);
xor U7029 (N_7029,N_4312,N_3712);
nor U7030 (N_7030,N_5155,N_5471);
nand U7031 (N_7031,N_4064,N_5719);
nor U7032 (N_7032,N_3383,N_3776);
or U7033 (N_7033,N_4013,N_3036);
or U7034 (N_7034,N_5073,N_4306);
xnor U7035 (N_7035,N_5695,N_3156);
or U7036 (N_7036,N_4597,N_4623);
nor U7037 (N_7037,N_4214,N_5324);
or U7038 (N_7038,N_4006,N_5859);
and U7039 (N_7039,N_4813,N_3460);
or U7040 (N_7040,N_5917,N_4585);
and U7041 (N_7041,N_3157,N_5075);
nor U7042 (N_7042,N_3139,N_4762);
and U7043 (N_7043,N_5681,N_3351);
nor U7044 (N_7044,N_3911,N_4650);
and U7045 (N_7045,N_4583,N_3658);
nor U7046 (N_7046,N_4556,N_5723);
and U7047 (N_7047,N_3816,N_3135);
nand U7048 (N_7048,N_3247,N_3057);
nand U7049 (N_7049,N_5726,N_3307);
or U7050 (N_7050,N_3440,N_5652);
or U7051 (N_7051,N_5836,N_4881);
nand U7052 (N_7052,N_4090,N_3340);
nand U7053 (N_7053,N_3804,N_4148);
xnor U7054 (N_7054,N_3283,N_4492);
nand U7055 (N_7055,N_3552,N_4122);
xor U7056 (N_7056,N_3878,N_3536);
nand U7057 (N_7057,N_5200,N_5772);
and U7058 (N_7058,N_4150,N_4714);
and U7059 (N_7059,N_4641,N_4052);
nor U7060 (N_7060,N_4311,N_4245);
nor U7061 (N_7061,N_3924,N_4309);
nand U7062 (N_7062,N_3664,N_3466);
or U7063 (N_7063,N_5559,N_5022);
and U7064 (N_7064,N_5015,N_5501);
nor U7065 (N_7065,N_4751,N_3936);
nand U7066 (N_7066,N_5475,N_5462);
and U7067 (N_7067,N_3784,N_3293);
nand U7068 (N_7068,N_3772,N_4584);
xor U7069 (N_7069,N_3957,N_4969);
or U7070 (N_7070,N_5997,N_4493);
and U7071 (N_7071,N_5873,N_4121);
and U7072 (N_7072,N_5848,N_3675);
xor U7073 (N_7073,N_3549,N_5352);
or U7074 (N_7074,N_3441,N_3054);
nand U7075 (N_7075,N_5245,N_5722);
nand U7076 (N_7076,N_4893,N_5027);
nand U7077 (N_7077,N_4942,N_4256);
nor U7078 (N_7078,N_5091,N_5487);
nand U7079 (N_7079,N_4652,N_5617);
nand U7080 (N_7080,N_3254,N_3790);
nor U7081 (N_7081,N_5994,N_5641);
or U7082 (N_7082,N_4102,N_3126);
and U7083 (N_7083,N_4627,N_3020);
and U7084 (N_7084,N_3341,N_5039);
and U7085 (N_7085,N_4169,N_5276);
or U7086 (N_7086,N_5546,N_4438);
and U7087 (N_7087,N_4433,N_4001);
or U7088 (N_7088,N_4464,N_3222);
or U7089 (N_7089,N_5574,N_3765);
nand U7090 (N_7090,N_4119,N_3107);
or U7091 (N_7091,N_3061,N_3715);
or U7092 (N_7092,N_5241,N_5921);
or U7093 (N_7093,N_3857,N_3578);
xnor U7094 (N_7094,N_5962,N_3964);
nand U7095 (N_7095,N_4277,N_5923);
and U7096 (N_7096,N_5940,N_4358);
nand U7097 (N_7097,N_3705,N_5296);
or U7098 (N_7098,N_4726,N_3348);
xnor U7099 (N_7099,N_3314,N_4728);
xor U7100 (N_7100,N_4968,N_4395);
nand U7101 (N_7101,N_3278,N_5125);
nand U7102 (N_7102,N_4788,N_3572);
nor U7103 (N_7103,N_4853,N_3067);
or U7104 (N_7104,N_4859,N_3714);
nand U7105 (N_7105,N_3782,N_4180);
nand U7106 (N_7106,N_3797,N_4683);
nand U7107 (N_7107,N_5506,N_3143);
nand U7108 (N_7108,N_3528,N_5749);
nor U7109 (N_7109,N_5538,N_4630);
nor U7110 (N_7110,N_4831,N_5438);
nand U7111 (N_7111,N_4285,N_3165);
and U7112 (N_7112,N_4593,N_4563);
nand U7113 (N_7113,N_5124,N_4573);
xnor U7114 (N_7114,N_3264,N_3203);
nand U7115 (N_7115,N_4453,N_3494);
or U7116 (N_7116,N_3554,N_3025);
or U7117 (N_7117,N_3459,N_5351);
nor U7118 (N_7118,N_4087,N_3993);
xor U7119 (N_7119,N_3731,N_4570);
nand U7120 (N_7120,N_5373,N_3325);
or U7121 (N_7121,N_4801,N_5484);
nor U7122 (N_7122,N_4704,N_5737);
xor U7123 (N_7123,N_3979,N_3401);
xnor U7124 (N_7124,N_5403,N_5457);
xnor U7125 (N_7125,N_4839,N_4029);
xnor U7126 (N_7126,N_5362,N_5411);
and U7127 (N_7127,N_4015,N_4690);
nor U7128 (N_7128,N_4069,N_4500);
xor U7129 (N_7129,N_3742,N_4457);
xor U7130 (N_7130,N_4930,N_4803);
or U7131 (N_7131,N_3799,N_5625);
and U7132 (N_7132,N_3539,N_3040);
nand U7133 (N_7133,N_4915,N_3623);
nor U7134 (N_7134,N_5933,N_4620);
xnor U7135 (N_7135,N_3323,N_4957);
nand U7136 (N_7136,N_5048,N_3329);
xnor U7137 (N_7137,N_3779,N_5725);
xor U7138 (N_7138,N_3234,N_4465);
nand U7139 (N_7139,N_3029,N_5131);
or U7140 (N_7140,N_5177,N_5530);
xnor U7141 (N_7141,N_3180,N_5611);
xnor U7142 (N_7142,N_3515,N_5498);
and U7143 (N_7143,N_3916,N_4882);
nor U7144 (N_7144,N_4209,N_5516);
or U7145 (N_7145,N_4402,N_5254);
nor U7146 (N_7146,N_5870,N_5399);
nor U7147 (N_7147,N_5545,N_5335);
and U7148 (N_7148,N_5821,N_4636);
nor U7149 (N_7149,N_3880,N_5375);
and U7150 (N_7150,N_3823,N_5754);
and U7151 (N_7151,N_5340,N_4460);
and U7152 (N_7152,N_5840,N_4676);
nor U7153 (N_7153,N_4625,N_3700);
or U7154 (N_7154,N_4307,N_5914);
or U7155 (N_7155,N_3858,N_4586);
nand U7156 (N_7156,N_4604,N_4958);
nor U7157 (N_7157,N_4514,N_4179);
nand U7158 (N_7158,N_3531,N_4338);
xnor U7159 (N_7159,N_3087,N_3828);
and U7160 (N_7160,N_3626,N_3346);
or U7161 (N_7161,N_3202,N_4362);
or U7162 (N_7162,N_4510,N_5651);
nor U7163 (N_7163,N_3537,N_4301);
xnor U7164 (N_7164,N_4239,N_5065);
and U7165 (N_7165,N_5079,N_3991);
nand U7166 (N_7166,N_5910,N_5686);
and U7167 (N_7167,N_3313,N_3914);
xnor U7168 (N_7168,N_3375,N_3954);
and U7169 (N_7169,N_3895,N_3793);
xor U7170 (N_7170,N_4458,N_4426);
nand U7171 (N_7171,N_5814,N_4466);
xnor U7172 (N_7172,N_3814,N_3822);
nor U7173 (N_7173,N_4523,N_3394);
and U7174 (N_7174,N_3689,N_5010);
nor U7175 (N_7175,N_4842,N_5337);
or U7176 (N_7176,N_5464,N_5382);
nand U7177 (N_7177,N_5138,N_5135);
nor U7178 (N_7178,N_4085,N_4346);
nor U7179 (N_7179,N_5232,N_5616);
nand U7180 (N_7180,N_3309,N_3558);
or U7181 (N_7181,N_5180,N_4835);
xor U7182 (N_7182,N_3559,N_3937);
and U7183 (N_7183,N_4633,N_3642);
nand U7184 (N_7184,N_5576,N_4101);
or U7185 (N_7185,N_4238,N_4328);
nand U7186 (N_7186,N_5706,N_4907);
nand U7187 (N_7187,N_4250,N_5769);
nor U7188 (N_7188,N_4010,N_4041);
nand U7189 (N_7189,N_3653,N_4616);
and U7190 (N_7190,N_5331,N_4546);
nor U7191 (N_7191,N_5841,N_5141);
and U7192 (N_7192,N_4158,N_3746);
or U7193 (N_7193,N_5955,N_3218);
nor U7194 (N_7194,N_4806,N_4117);
xnor U7195 (N_7195,N_4345,N_4494);
nand U7196 (N_7196,N_4656,N_4331);
nor U7197 (N_7197,N_5240,N_5322);
xor U7198 (N_7198,N_4192,N_5518);
nor U7199 (N_7199,N_5192,N_4425);
or U7200 (N_7200,N_5181,N_4336);
nor U7201 (N_7201,N_4321,N_3686);
and U7202 (N_7202,N_3477,N_3749);
or U7203 (N_7203,N_5868,N_3066);
nor U7204 (N_7204,N_4658,N_4737);
or U7205 (N_7205,N_3236,N_5262);
and U7206 (N_7206,N_5911,N_5212);
nor U7207 (N_7207,N_3637,N_3204);
xnor U7208 (N_7208,N_3767,N_5492);
nor U7209 (N_7209,N_5244,N_5427);
xor U7210 (N_7210,N_5313,N_5511);
and U7211 (N_7211,N_5550,N_5956);
and U7212 (N_7212,N_5665,N_3476);
nand U7213 (N_7213,N_5514,N_4442);
xnor U7214 (N_7214,N_5298,N_3942);
and U7215 (N_7215,N_3825,N_3787);
nand U7216 (N_7216,N_5489,N_4639);
and U7217 (N_7217,N_5046,N_3438);
nand U7218 (N_7218,N_5891,N_5216);
or U7219 (N_7219,N_3244,N_3287);
and U7220 (N_7220,N_5700,N_3555);
and U7221 (N_7221,N_3645,N_3786);
nor U7222 (N_7222,N_5062,N_4970);
or U7223 (N_7223,N_5415,N_4702);
or U7224 (N_7224,N_3212,N_3881);
nor U7225 (N_7225,N_5329,N_5374);
xnor U7226 (N_7226,N_4900,N_4031);
xor U7227 (N_7227,N_4962,N_5948);
xnor U7228 (N_7228,N_4843,N_3571);
and U7229 (N_7229,N_3602,N_5295);
xor U7230 (N_7230,N_5659,N_3453);
nor U7231 (N_7231,N_4902,N_3833);
or U7232 (N_7232,N_3353,N_3332);
xor U7233 (N_7233,N_4733,N_4800);
nor U7234 (N_7234,N_5718,N_3682);
and U7235 (N_7235,N_5768,N_3063);
or U7236 (N_7236,N_5547,N_5692);
xnor U7237 (N_7237,N_3673,N_5863);
nand U7238 (N_7238,N_5000,N_4896);
and U7239 (N_7239,N_5068,N_4678);
xnor U7240 (N_7240,N_3506,N_4434);
nor U7241 (N_7241,N_3586,N_5195);
and U7242 (N_7242,N_3333,N_5837);
nor U7243 (N_7243,N_3077,N_5267);
nor U7244 (N_7244,N_4384,N_3265);
nand U7245 (N_7245,N_3461,N_4241);
nand U7246 (N_7246,N_3465,N_5883);
or U7247 (N_7247,N_4254,N_4035);
or U7248 (N_7248,N_3223,N_5885);
nor U7249 (N_7249,N_4699,N_4125);
and U7250 (N_7250,N_4631,N_4992);
nor U7251 (N_7251,N_5058,N_3720);
and U7252 (N_7252,N_3492,N_3632);
xnor U7253 (N_7253,N_5263,N_3988);
nor U7254 (N_7254,N_5865,N_5654);
xnor U7255 (N_7255,N_3530,N_3649);
xnor U7256 (N_7256,N_5679,N_5328);
nor U7257 (N_7257,N_4174,N_4499);
xnor U7258 (N_7258,N_5653,N_3859);
xnor U7259 (N_7259,N_4231,N_4768);
or U7260 (N_7260,N_3366,N_5312);
and U7261 (N_7261,N_3211,N_4462);
xnor U7262 (N_7262,N_3527,N_5568);
nand U7263 (N_7263,N_4864,N_5724);
and U7264 (N_7264,N_3423,N_5913);
nor U7265 (N_7265,N_5886,N_5825);
and U7266 (N_7266,N_5712,N_3021);
and U7267 (N_7267,N_5284,N_3716);
nand U7268 (N_7268,N_4337,N_5716);
xnor U7269 (N_7269,N_4327,N_5691);
and U7270 (N_7270,N_4136,N_4377);
nor U7271 (N_7271,N_3953,N_5734);
xor U7272 (N_7272,N_5190,N_3024);
xor U7273 (N_7273,N_5607,N_3524);
and U7274 (N_7274,N_4512,N_4264);
nand U7275 (N_7275,N_3148,N_4703);
nand U7276 (N_7276,N_3678,N_4441);
nand U7277 (N_7277,N_5784,N_3129);
nor U7278 (N_7278,N_3277,N_3728);
nor U7279 (N_7279,N_4359,N_5072);
xnor U7280 (N_7280,N_3274,N_3813);
nor U7281 (N_7281,N_5144,N_4288);
and U7282 (N_7282,N_3300,N_5708);
or U7283 (N_7283,N_3147,N_5937);
xor U7284 (N_7284,N_3758,N_5526);
nand U7285 (N_7285,N_3923,N_5992);
or U7286 (N_7286,N_5759,N_4611);
and U7287 (N_7287,N_3990,N_3369);
or U7288 (N_7288,N_3604,N_3153);
xnor U7289 (N_7289,N_5260,N_5936);
xor U7290 (N_7290,N_3655,N_5453);
nor U7291 (N_7291,N_5694,N_3056);
nor U7292 (N_7292,N_5764,N_4497);
xor U7293 (N_7293,N_3017,N_4372);
or U7294 (N_7294,N_4927,N_5202);
nor U7295 (N_7295,N_4820,N_4989);
nor U7296 (N_7296,N_3395,N_3224);
or U7297 (N_7297,N_3702,N_3511);
xor U7298 (N_7298,N_5274,N_4221);
xor U7299 (N_7299,N_5658,N_5099);
or U7300 (N_7300,N_4190,N_3760);
nand U7301 (N_7301,N_5970,N_5874);
nor U7302 (N_7302,N_3576,N_4296);
xnor U7303 (N_7303,N_3084,N_4503);
nand U7304 (N_7304,N_5060,N_5114);
nor U7305 (N_7305,N_5412,N_4976);
xnor U7306 (N_7306,N_4200,N_5666);
nand U7307 (N_7307,N_4617,N_4024);
nor U7308 (N_7308,N_5844,N_4838);
nor U7309 (N_7309,N_4742,N_4414);
and U7310 (N_7310,N_5221,N_3479);
nand U7311 (N_7311,N_4406,N_3392);
or U7312 (N_7312,N_4258,N_3510);
nor U7313 (N_7313,N_3920,N_4872);
and U7314 (N_7314,N_3000,N_4474);
and U7315 (N_7315,N_5025,N_5548);
and U7316 (N_7316,N_3542,N_5127);
nand U7317 (N_7317,N_4455,N_5306);
nand U7318 (N_7318,N_5297,N_5490);
or U7319 (N_7319,N_3112,N_3676);
nor U7320 (N_7320,N_4273,N_3240);
xnor U7321 (N_7321,N_3407,N_4753);
nor U7322 (N_7322,N_5947,N_4261);
or U7323 (N_7323,N_4995,N_4594);
nor U7324 (N_7324,N_3907,N_5341);
and U7325 (N_7325,N_3780,N_4607);
or U7326 (N_7326,N_4738,N_3195);
nor U7327 (N_7327,N_3817,N_3652);
nor U7328 (N_7328,N_5308,N_3888);
nand U7329 (N_7329,N_5871,N_3995);
xnor U7330 (N_7330,N_5201,N_5774);
and U7331 (N_7331,N_4732,N_5707);
nor U7332 (N_7332,N_4120,N_3417);
nor U7333 (N_7333,N_5220,N_5587);
nor U7334 (N_7334,N_3327,N_3748);
nor U7335 (N_7335,N_3753,N_5052);
and U7336 (N_7336,N_5519,N_5633);
and U7337 (N_7337,N_4719,N_3906);
and U7338 (N_7338,N_5971,N_5960);
nor U7339 (N_7339,N_4706,N_4487);
xor U7340 (N_7340,N_3415,N_4089);
nor U7341 (N_7341,N_3781,N_5969);
nand U7342 (N_7342,N_5687,N_4536);
or U7343 (N_7343,N_4019,N_5893);
nand U7344 (N_7344,N_4157,N_5565);
xnor U7345 (N_7345,N_5074,N_3577);
xor U7346 (N_7346,N_4039,N_5164);
nor U7347 (N_7347,N_5527,N_4707);
nor U7348 (N_7348,N_5139,N_3362);
xor U7349 (N_7349,N_4953,N_5736);
and U7350 (N_7350,N_3259,N_4854);
nor U7351 (N_7351,N_3382,N_5430);
xor U7352 (N_7352,N_3373,N_3667);
nor U7353 (N_7353,N_4279,N_5395);
and U7354 (N_7354,N_4955,N_3381);
nand U7355 (N_7355,N_3450,N_4691);
nor U7356 (N_7356,N_3088,N_3927);
and U7357 (N_7357,N_5294,N_3970);
nand U7358 (N_7358,N_4817,N_5230);
xnor U7359 (N_7359,N_3294,N_3261);
and U7360 (N_7360,N_4204,N_3629);
nor U7361 (N_7361,N_4755,N_4929);
nand U7362 (N_7362,N_5226,N_3422);
xor U7363 (N_7363,N_5615,N_3481);
or U7364 (N_7364,N_3861,N_4207);
nand U7365 (N_7365,N_5567,N_3745);
nor U7366 (N_7366,N_3186,N_5129);
nand U7367 (N_7367,N_4675,N_4997);
nor U7368 (N_7368,N_3614,N_3113);
or U7369 (N_7369,N_4443,N_4875);
nor U7370 (N_7370,N_3762,N_3489);
nor U7371 (N_7371,N_4314,N_4368);
or U7372 (N_7372,N_5533,N_4897);
nor U7373 (N_7373,N_4936,N_4078);
or U7374 (N_7374,N_4983,N_3266);
or U7375 (N_7375,N_4275,N_5023);
nor U7376 (N_7376,N_4521,N_3615);
and U7377 (N_7377,N_4373,N_4612);
xor U7378 (N_7378,N_5327,N_5132);
nor U7379 (N_7379,N_3349,N_4060);
and U7380 (N_7380,N_3311,N_4223);
nor U7381 (N_7381,N_4802,N_3631);
xor U7382 (N_7382,N_5974,N_5183);
and U7383 (N_7383,N_4292,N_4723);
and U7384 (N_7384,N_5169,N_3435);
or U7385 (N_7385,N_4452,N_4679);
nor U7386 (N_7386,N_3421,N_4176);
and U7387 (N_7387,N_4822,N_5149);
xnor U7388 (N_7388,N_4736,N_4833);
xor U7389 (N_7389,N_5101,N_4663);
nor U7390 (N_7390,N_4246,N_4876);
nand U7391 (N_7391,N_4909,N_4587);
nor U7392 (N_7392,N_3041,N_5701);
xnor U7393 (N_7393,N_4408,N_5247);
nor U7394 (N_7394,N_4183,N_3098);
or U7395 (N_7395,N_4477,N_4429);
or U7396 (N_7396,N_4083,N_4023);
and U7397 (N_7397,N_5198,N_3093);
and U7398 (N_7398,N_3850,N_3225);
xor U7399 (N_7399,N_4505,N_4081);
and U7400 (N_7400,N_5270,N_3915);
xor U7401 (N_7401,N_3946,N_4249);
xor U7402 (N_7402,N_5812,N_3893);
or U7403 (N_7403,N_5054,N_5320);
nand U7404 (N_7404,N_4175,N_5483);
and U7405 (N_7405,N_4722,N_4777);
and U7406 (N_7406,N_4520,N_5693);
or U7407 (N_7407,N_5359,N_4760);
nor U7408 (N_7408,N_5756,N_5811);
nand U7409 (N_7409,N_3060,N_4850);
nor U7410 (N_7410,N_4647,N_3413);
nor U7411 (N_7411,N_4591,N_5697);
nand U7412 (N_7412,N_3445,N_4533);
or U7413 (N_7413,N_3100,N_3583);
nor U7414 (N_7414,N_4659,N_3121);
nor U7415 (N_7415,N_3874,N_3759);
or U7416 (N_7416,N_5922,N_5668);
nand U7417 (N_7417,N_4614,N_4410);
xor U7418 (N_7418,N_5878,N_5397);
nor U7419 (N_7419,N_4933,N_5019);
and U7420 (N_7420,N_5042,N_4335);
nand U7421 (N_7421,N_5996,N_3863);
or U7422 (N_7422,N_5564,N_4048);
xnor U7423 (N_7423,N_5299,N_4482);
nand U7424 (N_7424,N_5536,N_4787);
or U7425 (N_7425,N_5508,N_4606);
nor U7426 (N_7426,N_3232,N_3167);
xor U7427 (N_7427,N_5421,N_4283);
and U7428 (N_7428,N_3175,N_4527);
nand U7429 (N_7429,N_4660,N_4084);
nor U7430 (N_7430,N_4602,N_4077);
xnor U7431 (N_7431,N_3560,N_4873);
or U7432 (N_7432,N_5702,N_3312);
and U7433 (N_7433,N_5339,N_5163);
and U7434 (N_7434,N_4271,N_4056);
or U7435 (N_7435,N_5856,N_3397);
xor U7436 (N_7436,N_4539,N_5562);
xor U7437 (N_7437,N_3699,N_3451);
or U7438 (N_7438,N_3152,N_5809);
xnor U7439 (N_7439,N_4626,N_5849);
xor U7440 (N_7440,N_3010,N_4735);
xnor U7441 (N_7441,N_5946,N_5476);
or U7442 (N_7442,N_5703,N_4515);
nand U7443 (N_7443,N_3744,N_5973);
nand U7444 (N_7444,N_3412,N_3876);
xnor U7445 (N_7445,N_3679,N_3590);
nand U7446 (N_7446,N_3769,N_5280);
nor U7447 (N_7447,N_5683,N_5524);
nor U7448 (N_7448,N_3377,N_4693);
nor U7449 (N_7449,N_3114,N_3306);
nand U7450 (N_7450,N_5358,N_4181);
and U7451 (N_7451,N_5105,N_3251);
nand U7452 (N_7452,N_4226,N_4218);
xor U7453 (N_7453,N_4860,N_3805);
xor U7454 (N_7454,N_3030,N_3566);
or U7455 (N_7455,N_5613,N_3975);
xor U7456 (N_7456,N_4280,N_5379);
and U7457 (N_7457,N_3386,N_5684);
nor U7458 (N_7458,N_4904,N_4905);
xor U7459 (N_7459,N_5813,N_4852);
xor U7460 (N_7460,N_5831,N_4252);
xnor U7461 (N_7461,N_4984,N_3869);
xor U7462 (N_7462,N_4910,N_3809);
nor U7463 (N_7463,N_3684,N_3969);
nand U7464 (N_7464,N_4645,N_4987);
nor U7465 (N_7465,N_4488,N_4734);
xnor U7466 (N_7466,N_4422,N_4766);
or U7467 (N_7467,N_5342,N_5951);
or U7468 (N_7468,N_3269,N_5108);
xor U7469 (N_7469,N_4507,N_5934);
xnor U7470 (N_7470,N_4759,N_4891);
and U7471 (N_7471,N_5915,N_5906);
xor U7472 (N_7472,N_5182,N_5189);
xor U7473 (N_7473,N_3482,N_5714);
nand U7474 (N_7474,N_4012,N_3981);
xor U7475 (N_7475,N_3171,N_4316);
nor U7476 (N_7476,N_4863,N_4596);
nand U7477 (N_7477,N_5235,N_3903);
nand U7478 (N_7478,N_4739,N_3670);
or U7479 (N_7479,N_5185,N_4388);
and U7480 (N_7480,N_4291,N_3704);
nand U7481 (N_7481,N_4856,N_4532);
xor U7482 (N_7482,N_5017,N_3561);
nor U7483 (N_7483,N_5672,N_4430);
nor U7484 (N_7484,N_4743,N_3321);
xor U7485 (N_7485,N_5918,N_3120);
nand U7486 (N_7486,N_5009,N_3145);
xor U7487 (N_7487,N_3233,N_3430);
or U7488 (N_7488,N_4114,N_5602);
nand U7489 (N_7489,N_3243,N_5392);
xnor U7490 (N_7490,N_4066,N_3344);
nand U7491 (N_7491,N_3282,N_3921);
and U7492 (N_7492,N_3324,N_4033);
nor U7493 (N_7493,N_4416,N_5387);
and U7494 (N_7494,N_3291,N_5111);
nand U7495 (N_7495,N_4215,N_3865);
or U7496 (N_7496,N_5667,N_3801);
nand U7497 (N_7497,N_4629,N_5447);
nand U7498 (N_7498,N_5434,N_3316);
nand U7499 (N_7499,N_4063,N_4014);
nand U7500 (N_7500,N_3109,N_3236);
and U7501 (N_7501,N_5948,N_4736);
xor U7502 (N_7502,N_4986,N_5566);
xnor U7503 (N_7503,N_5139,N_5674);
xnor U7504 (N_7504,N_4011,N_5166);
and U7505 (N_7505,N_3481,N_3344);
and U7506 (N_7506,N_5948,N_3613);
or U7507 (N_7507,N_4527,N_4602);
or U7508 (N_7508,N_5154,N_3013);
xnor U7509 (N_7509,N_5954,N_4981);
nand U7510 (N_7510,N_4531,N_4191);
and U7511 (N_7511,N_5964,N_4143);
xnor U7512 (N_7512,N_5628,N_4444);
xnor U7513 (N_7513,N_4658,N_4601);
and U7514 (N_7514,N_4676,N_4461);
and U7515 (N_7515,N_5994,N_5242);
or U7516 (N_7516,N_3332,N_5595);
and U7517 (N_7517,N_5762,N_5565);
nor U7518 (N_7518,N_3929,N_4528);
nand U7519 (N_7519,N_3498,N_3436);
xor U7520 (N_7520,N_5968,N_5223);
nand U7521 (N_7521,N_5156,N_3975);
or U7522 (N_7522,N_4980,N_5885);
nor U7523 (N_7523,N_3687,N_3751);
or U7524 (N_7524,N_4325,N_3460);
xnor U7525 (N_7525,N_3413,N_4503);
and U7526 (N_7526,N_3620,N_5915);
and U7527 (N_7527,N_4791,N_5682);
and U7528 (N_7528,N_4965,N_5651);
nand U7529 (N_7529,N_4301,N_5817);
nor U7530 (N_7530,N_4176,N_3091);
or U7531 (N_7531,N_3062,N_4218);
nor U7532 (N_7532,N_3334,N_5141);
or U7533 (N_7533,N_5470,N_5720);
xor U7534 (N_7534,N_3214,N_4511);
xor U7535 (N_7535,N_3644,N_3775);
nand U7536 (N_7536,N_3250,N_3561);
and U7537 (N_7537,N_5262,N_4954);
and U7538 (N_7538,N_3953,N_5763);
and U7539 (N_7539,N_5561,N_4107);
and U7540 (N_7540,N_3146,N_3391);
or U7541 (N_7541,N_3955,N_3421);
nand U7542 (N_7542,N_5151,N_3248);
xor U7543 (N_7543,N_5860,N_3521);
and U7544 (N_7544,N_4174,N_5532);
and U7545 (N_7545,N_4702,N_3755);
nor U7546 (N_7546,N_5655,N_5163);
and U7547 (N_7547,N_4320,N_4599);
or U7548 (N_7548,N_3214,N_4712);
nor U7549 (N_7549,N_5293,N_4326);
nor U7550 (N_7550,N_5908,N_3721);
nand U7551 (N_7551,N_4631,N_5663);
nor U7552 (N_7552,N_5822,N_5043);
and U7553 (N_7553,N_4183,N_3420);
nor U7554 (N_7554,N_4896,N_5781);
nor U7555 (N_7555,N_5999,N_4487);
or U7556 (N_7556,N_5882,N_3471);
nand U7557 (N_7557,N_5233,N_3862);
nand U7558 (N_7558,N_5453,N_5166);
nor U7559 (N_7559,N_3370,N_4251);
or U7560 (N_7560,N_3962,N_5272);
nor U7561 (N_7561,N_4005,N_3161);
and U7562 (N_7562,N_4064,N_3844);
xnor U7563 (N_7563,N_3591,N_5682);
xnor U7564 (N_7564,N_4220,N_4242);
xor U7565 (N_7565,N_3868,N_5127);
nand U7566 (N_7566,N_5048,N_3224);
nor U7567 (N_7567,N_4080,N_5230);
nor U7568 (N_7568,N_5336,N_5952);
nand U7569 (N_7569,N_4787,N_4951);
and U7570 (N_7570,N_4640,N_4955);
nor U7571 (N_7571,N_5840,N_4039);
xor U7572 (N_7572,N_3977,N_4697);
xor U7573 (N_7573,N_3224,N_5590);
nand U7574 (N_7574,N_5975,N_3754);
and U7575 (N_7575,N_3835,N_5518);
xor U7576 (N_7576,N_3102,N_3284);
or U7577 (N_7577,N_3209,N_3717);
nor U7578 (N_7578,N_5760,N_4997);
nand U7579 (N_7579,N_4358,N_4128);
and U7580 (N_7580,N_3596,N_3060);
and U7581 (N_7581,N_3118,N_5997);
and U7582 (N_7582,N_3372,N_4865);
nor U7583 (N_7583,N_3739,N_4822);
or U7584 (N_7584,N_5902,N_5228);
and U7585 (N_7585,N_5259,N_4344);
nor U7586 (N_7586,N_3370,N_4141);
and U7587 (N_7587,N_4647,N_3049);
and U7588 (N_7588,N_4989,N_4849);
nor U7589 (N_7589,N_5223,N_3734);
and U7590 (N_7590,N_5387,N_3397);
nor U7591 (N_7591,N_4821,N_4995);
nor U7592 (N_7592,N_5230,N_3105);
or U7593 (N_7593,N_5864,N_3930);
nor U7594 (N_7594,N_4066,N_4239);
or U7595 (N_7595,N_5091,N_3384);
xnor U7596 (N_7596,N_4769,N_3862);
nand U7597 (N_7597,N_3014,N_5748);
and U7598 (N_7598,N_4056,N_4310);
and U7599 (N_7599,N_3844,N_4164);
xnor U7600 (N_7600,N_3920,N_5668);
and U7601 (N_7601,N_5220,N_3832);
or U7602 (N_7602,N_5796,N_5950);
xor U7603 (N_7603,N_5547,N_4913);
or U7604 (N_7604,N_5276,N_3594);
and U7605 (N_7605,N_4616,N_4725);
and U7606 (N_7606,N_4550,N_5435);
xor U7607 (N_7607,N_4895,N_3047);
and U7608 (N_7608,N_4080,N_3033);
nor U7609 (N_7609,N_3212,N_4677);
nand U7610 (N_7610,N_4615,N_4743);
nor U7611 (N_7611,N_4932,N_5659);
nor U7612 (N_7612,N_5694,N_5867);
nor U7613 (N_7613,N_5972,N_3953);
and U7614 (N_7614,N_4668,N_3581);
nor U7615 (N_7615,N_3348,N_5505);
xor U7616 (N_7616,N_4057,N_4059);
xnor U7617 (N_7617,N_3500,N_5471);
and U7618 (N_7618,N_3485,N_4634);
and U7619 (N_7619,N_5718,N_3200);
or U7620 (N_7620,N_3517,N_5215);
xor U7621 (N_7621,N_4610,N_4080);
or U7622 (N_7622,N_3277,N_4381);
or U7623 (N_7623,N_3920,N_4771);
nand U7624 (N_7624,N_3262,N_5652);
nor U7625 (N_7625,N_4808,N_4734);
nand U7626 (N_7626,N_4722,N_3162);
xnor U7627 (N_7627,N_4525,N_3930);
nand U7628 (N_7628,N_4010,N_5103);
xnor U7629 (N_7629,N_4979,N_3093);
nand U7630 (N_7630,N_3077,N_4401);
xor U7631 (N_7631,N_3364,N_3626);
and U7632 (N_7632,N_4064,N_5214);
or U7633 (N_7633,N_3683,N_3165);
or U7634 (N_7634,N_5019,N_4504);
or U7635 (N_7635,N_5420,N_4752);
or U7636 (N_7636,N_4527,N_5520);
or U7637 (N_7637,N_3327,N_5822);
or U7638 (N_7638,N_4093,N_5046);
nand U7639 (N_7639,N_5322,N_5164);
xor U7640 (N_7640,N_4821,N_5976);
nand U7641 (N_7641,N_5995,N_3669);
or U7642 (N_7642,N_5718,N_3425);
nand U7643 (N_7643,N_5127,N_4788);
nand U7644 (N_7644,N_4228,N_3662);
or U7645 (N_7645,N_4210,N_5868);
nand U7646 (N_7646,N_3269,N_4775);
nand U7647 (N_7647,N_4576,N_3475);
nand U7648 (N_7648,N_5718,N_5192);
nand U7649 (N_7649,N_5485,N_4363);
nand U7650 (N_7650,N_3404,N_3853);
or U7651 (N_7651,N_4171,N_3854);
nand U7652 (N_7652,N_3393,N_3311);
or U7653 (N_7653,N_4871,N_4018);
nor U7654 (N_7654,N_4529,N_5287);
xnor U7655 (N_7655,N_4591,N_3978);
and U7656 (N_7656,N_5049,N_3542);
or U7657 (N_7657,N_5934,N_3904);
nor U7658 (N_7658,N_3171,N_3832);
or U7659 (N_7659,N_4453,N_4621);
or U7660 (N_7660,N_4132,N_5280);
nand U7661 (N_7661,N_5080,N_3240);
or U7662 (N_7662,N_4844,N_5847);
or U7663 (N_7663,N_4905,N_4873);
xnor U7664 (N_7664,N_5645,N_3679);
xnor U7665 (N_7665,N_4880,N_3739);
or U7666 (N_7666,N_3072,N_4286);
nand U7667 (N_7667,N_3651,N_4885);
and U7668 (N_7668,N_3516,N_4839);
xor U7669 (N_7669,N_4667,N_4122);
nor U7670 (N_7670,N_3441,N_3521);
and U7671 (N_7671,N_5495,N_5761);
xor U7672 (N_7672,N_5903,N_4113);
nor U7673 (N_7673,N_4721,N_3133);
nand U7674 (N_7674,N_5483,N_3321);
nor U7675 (N_7675,N_5794,N_4924);
nor U7676 (N_7676,N_3017,N_4973);
and U7677 (N_7677,N_5742,N_5249);
and U7678 (N_7678,N_3262,N_5464);
or U7679 (N_7679,N_3313,N_5433);
and U7680 (N_7680,N_5144,N_5838);
or U7681 (N_7681,N_5065,N_5740);
nand U7682 (N_7682,N_5338,N_5857);
nand U7683 (N_7683,N_4418,N_5403);
and U7684 (N_7684,N_4378,N_5042);
nand U7685 (N_7685,N_4576,N_4252);
and U7686 (N_7686,N_3352,N_3903);
and U7687 (N_7687,N_3549,N_5710);
xnor U7688 (N_7688,N_3318,N_4727);
nor U7689 (N_7689,N_3802,N_5157);
and U7690 (N_7690,N_3953,N_3557);
xor U7691 (N_7691,N_5112,N_4061);
nor U7692 (N_7692,N_5995,N_3846);
or U7693 (N_7693,N_4944,N_4714);
and U7694 (N_7694,N_3736,N_4065);
nor U7695 (N_7695,N_4955,N_4545);
nor U7696 (N_7696,N_4200,N_4692);
xor U7697 (N_7697,N_3918,N_4846);
nor U7698 (N_7698,N_4919,N_4296);
xnor U7699 (N_7699,N_3941,N_3354);
nor U7700 (N_7700,N_5901,N_3650);
xnor U7701 (N_7701,N_5867,N_3343);
and U7702 (N_7702,N_4177,N_3226);
nor U7703 (N_7703,N_5114,N_4508);
xnor U7704 (N_7704,N_5349,N_4703);
and U7705 (N_7705,N_3371,N_3771);
nand U7706 (N_7706,N_4973,N_5838);
nand U7707 (N_7707,N_5213,N_4670);
xor U7708 (N_7708,N_3403,N_3023);
nand U7709 (N_7709,N_4858,N_3931);
and U7710 (N_7710,N_4026,N_3436);
and U7711 (N_7711,N_4614,N_5800);
xor U7712 (N_7712,N_4932,N_3943);
or U7713 (N_7713,N_4947,N_5288);
or U7714 (N_7714,N_4615,N_5774);
nor U7715 (N_7715,N_5990,N_3169);
nand U7716 (N_7716,N_3161,N_4794);
xnor U7717 (N_7717,N_3152,N_4403);
and U7718 (N_7718,N_5291,N_5913);
nor U7719 (N_7719,N_4230,N_4241);
xnor U7720 (N_7720,N_4502,N_5118);
nor U7721 (N_7721,N_5897,N_4840);
nand U7722 (N_7722,N_4006,N_3059);
or U7723 (N_7723,N_3386,N_3219);
xor U7724 (N_7724,N_3063,N_5042);
nor U7725 (N_7725,N_4219,N_4329);
xor U7726 (N_7726,N_3463,N_5381);
or U7727 (N_7727,N_3644,N_4249);
xnor U7728 (N_7728,N_4637,N_3304);
nand U7729 (N_7729,N_4644,N_3899);
nor U7730 (N_7730,N_4734,N_5267);
and U7731 (N_7731,N_4154,N_3965);
nor U7732 (N_7732,N_3652,N_5871);
nor U7733 (N_7733,N_5412,N_4257);
and U7734 (N_7734,N_4670,N_5167);
xnor U7735 (N_7735,N_4096,N_5168);
nor U7736 (N_7736,N_3202,N_3275);
xor U7737 (N_7737,N_5492,N_5679);
or U7738 (N_7738,N_3700,N_5692);
or U7739 (N_7739,N_4931,N_4541);
and U7740 (N_7740,N_4533,N_3299);
and U7741 (N_7741,N_5890,N_4658);
xnor U7742 (N_7742,N_3370,N_4008);
nor U7743 (N_7743,N_3524,N_5658);
nand U7744 (N_7744,N_4674,N_4280);
xnor U7745 (N_7745,N_4356,N_5729);
xor U7746 (N_7746,N_5671,N_5937);
nand U7747 (N_7747,N_5763,N_3100);
or U7748 (N_7748,N_3998,N_4081);
nand U7749 (N_7749,N_3587,N_4944);
or U7750 (N_7750,N_5165,N_3479);
nor U7751 (N_7751,N_4318,N_3592);
or U7752 (N_7752,N_4835,N_4153);
xnor U7753 (N_7753,N_5891,N_3403);
or U7754 (N_7754,N_3298,N_5959);
and U7755 (N_7755,N_4640,N_4776);
nor U7756 (N_7756,N_4789,N_5643);
nor U7757 (N_7757,N_4626,N_5545);
or U7758 (N_7758,N_3765,N_4183);
nand U7759 (N_7759,N_3219,N_4311);
or U7760 (N_7760,N_4228,N_3522);
xor U7761 (N_7761,N_3438,N_3423);
xor U7762 (N_7762,N_4227,N_5342);
nor U7763 (N_7763,N_3606,N_4269);
and U7764 (N_7764,N_3201,N_4266);
or U7765 (N_7765,N_4005,N_4262);
xnor U7766 (N_7766,N_5836,N_4247);
and U7767 (N_7767,N_4480,N_4812);
or U7768 (N_7768,N_3729,N_4077);
and U7769 (N_7769,N_3824,N_3540);
and U7770 (N_7770,N_5219,N_5207);
nand U7771 (N_7771,N_3914,N_3147);
or U7772 (N_7772,N_5404,N_3638);
and U7773 (N_7773,N_3097,N_5665);
nor U7774 (N_7774,N_3672,N_4056);
xnor U7775 (N_7775,N_5896,N_3148);
nand U7776 (N_7776,N_4519,N_3227);
and U7777 (N_7777,N_5091,N_3313);
xor U7778 (N_7778,N_5609,N_4806);
nor U7779 (N_7779,N_5000,N_4004);
or U7780 (N_7780,N_4536,N_3263);
nand U7781 (N_7781,N_4036,N_3427);
xor U7782 (N_7782,N_5829,N_3894);
and U7783 (N_7783,N_3158,N_4856);
and U7784 (N_7784,N_3200,N_5052);
nor U7785 (N_7785,N_4628,N_4162);
nor U7786 (N_7786,N_3495,N_4751);
nor U7787 (N_7787,N_3390,N_4980);
or U7788 (N_7788,N_4329,N_4059);
xnor U7789 (N_7789,N_4405,N_3059);
nand U7790 (N_7790,N_4272,N_5365);
nand U7791 (N_7791,N_5206,N_3606);
nor U7792 (N_7792,N_3985,N_5167);
xor U7793 (N_7793,N_3715,N_3423);
nor U7794 (N_7794,N_4267,N_5905);
xnor U7795 (N_7795,N_4113,N_3801);
and U7796 (N_7796,N_5507,N_4757);
and U7797 (N_7797,N_5017,N_4808);
xnor U7798 (N_7798,N_3590,N_4423);
nand U7799 (N_7799,N_3467,N_5213);
or U7800 (N_7800,N_3800,N_5516);
nand U7801 (N_7801,N_5152,N_3986);
nor U7802 (N_7802,N_5597,N_3193);
xnor U7803 (N_7803,N_4105,N_3737);
xnor U7804 (N_7804,N_5007,N_4950);
or U7805 (N_7805,N_4785,N_4379);
nor U7806 (N_7806,N_5118,N_3987);
or U7807 (N_7807,N_5143,N_3943);
nand U7808 (N_7808,N_4263,N_5411);
xor U7809 (N_7809,N_3158,N_5600);
nand U7810 (N_7810,N_5883,N_4369);
nor U7811 (N_7811,N_3013,N_3255);
nand U7812 (N_7812,N_4280,N_4013);
nor U7813 (N_7813,N_3158,N_4421);
or U7814 (N_7814,N_5182,N_3778);
and U7815 (N_7815,N_3339,N_5778);
and U7816 (N_7816,N_5067,N_5863);
and U7817 (N_7817,N_5130,N_5648);
nand U7818 (N_7818,N_4218,N_3024);
or U7819 (N_7819,N_5571,N_5527);
nand U7820 (N_7820,N_5065,N_5175);
and U7821 (N_7821,N_5586,N_4401);
and U7822 (N_7822,N_3255,N_5203);
nand U7823 (N_7823,N_5714,N_4656);
xor U7824 (N_7824,N_3837,N_3207);
xor U7825 (N_7825,N_5699,N_4951);
nor U7826 (N_7826,N_5752,N_4029);
and U7827 (N_7827,N_5620,N_3479);
nor U7828 (N_7828,N_4936,N_4929);
and U7829 (N_7829,N_4155,N_3843);
or U7830 (N_7830,N_4531,N_3250);
nor U7831 (N_7831,N_5473,N_4999);
and U7832 (N_7832,N_5181,N_3642);
nand U7833 (N_7833,N_4963,N_3440);
xor U7834 (N_7834,N_4921,N_4585);
nand U7835 (N_7835,N_3073,N_3653);
or U7836 (N_7836,N_3625,N_4721);
xor U7837 (N_7837,N_3768,N_5825);
nor U7838 (N_7838,N_5204,N_4025);
or U7839 (N_7839,N_3088,N_5750);
or U7840 (N_7840,N_3469,N_3016);
nand U7841 (N_7841,N_4810,N_5644);
xor U7842 (N_7842,N_5305,N_4697);
nor U7843 (N_7843,N_5743,N_5589);
nand U7844 (N_7844,N_3914,N_4869);
and U7845 (N_7845,N_3821,N_4397);
xor U7846 (N_7846,N_4851,N_3096);
nand U7847 (N_7847,N_3398,N_4616);
xor U7848 (N_7848,N_4698,N_5253);
xnor U7849 (N_7849,N_3813,N_4791);
or U7850 (N_7850,N_3953,N_4969);
xnor U7851 (N_7851,N_4000,N_3531);
or U7852 (N_7852,N_5240,N_5610);
nor U7853 (N_7853,N_5802,N_3306);
nand U7854 (N_7854,N_4091,N_5110);
or U7855 (N_7855,N_5579,N_4298);
nor U7856 (N_7856,N_4791,N_5229);
and U7857 (N_7857,N_3410,N_5319);
nor U7858 (N_7858,N_5039,N_4397);
nor U7859 (N_7859,N_5782,N_5911);
and U7860 (N_7860,N_3378,N_5973);
nor U7861 (N_7861,N_5371,N_3759);
or U7862 (N_7862,N_5702,N_5586);
nor U7863 (N_7863,N_5440,N_3518);
nor U7864 (N_7864,N_5663,N_3094);
nor U7865 (N_7865,N_3465,N_3340);
and U7866 (N_7866,N_5025,N_5330);
xor U7867 (N_7867,N_3270,N_4896);
and U7868 (N_7868,N_4097,N_3850);
xor U7869 (N_7869,N_4448,N_5894);
xnor U7870 (N_7870,N_3432,N_5839);
or U7871 (N_7871,N_4639,N_4468);
nor U7872 (N_7872,N_5438,N_5108);
or U7873 (N_7873,N_5325,N_5854);
nor U7874 (N_7874,N_5125,N_4985);
and U7875 (N_7875,N_3864,N_3512);
xor U7876 (N_7876,N_4532,N_5373);
xor U7877 (N_7877,N_3651,N_4449);
or U7878 (N_7878,N_4830,N_3574);
and U7879 (N_7879,N_4181,N_5161);
nor U7880 (N_7880,N_5904,N_5668);
nor U7881 (N_7881,N_5470,N_5461);
and U7882 (N_7882,N_5983,N_5937);
nor U7883 (N_7883,N_4817,N_4139);
or U7884 (N_7884,N_4621,N_3183);
and U7885 (N_7885,N_5380,N_3212);
nor U7886 (N_7886,N_3169,N_5173);
xnor U7887 (N_7887,N_3129,N_5419);
and U7888 (N_7888,N_4979,N_5660);
or U7889 (N_7889,N_5809,N_5582);
nand U7890 (N_7890,N_3725,N_3208);
xnor U7891 (N_7891,N_3246,N_4811);
or U7892 (N_7892,N_4322,N_3948);
xnor U7893 (N_7893,N_4037,N_3430);
xnor U7894 (N_7894,N_4940,N_5870);
nor U7895 (N_7895,N_5556,N_3948);
or U7896 (N_7896,N_5670,N_3997);
and U7897 (N_7897,N_3990,N_3442);
nand U7898 (N_7898,N_5541,N_5843);
and U7899 (N_7899,N_3576,N_4277);
and U7900 (N_7900,N_5041,N_5895);
nor U7901 (N_7901,N_4027,N_3473);
or U7902 (N_7902,N_4845,N_4839);
nor U7903 (N_7903,N_5448,N_3879);
nand U7904 (N_7904,N_4607,N_3726);
and U7905 (N_7905,N_5538,N_5125);
or U7906 (N_7906,N_5592,N_4281);
and U7907 (N_7907,N_4248,N_4732);
nor U7908 (N_7908,N_4092,N_4437);
and U7909 (N_7909,N_4924,N_5008);
nand U7910 (N_7910,N_3834,N_3719);
nor U7911 (N_7911,N_3263,N_4041);
xnor U7912 (N_7912,N_3747,N_5412);
xor U7913 (N_7913,N_4166,N_3209);
or U7914 (N_7914,N_3260,N_4256);
nor U7915 (N_7915,N_4762,N_5056);
and U7916 (N_7916,N_5929,N_5869);
nand U7917 (N_7917,N_5517,N_5008);
nand U7918 (N_7918,N_4496,N_5371);
or U7919 (N_7919,N_4769,N_5183);
nor U7920 (N_7920,N_5525,N_3372);
nand U7921 (N_7921,N_3382,N_5589);
xnor U7922 (N_7922,N_3672,N_5251);
nor U7923 (N_7923,N_5377,N_3630);
xnor U7924 (N_7924,N_3134,N_5640);
xor U7925 (N_7925,N_5014,N_4113);
xnor U7926 (N_7926,N_5700,N_3395);
and U7927 (N_7927,N_4640,N_5285);
nand U7928 (N_7928,N_4269,N_3584);
or U7929 (N_7929,N_5222,N_4914);
xor U7930 (N_7930,N_3130,N_4110);
nor U7931 (N_7931,N_4391,N_4067);
nand U7932 (N_7932,N_5926,N_5265);
or U7933 (N_7933,N_5368,N_5859);
and U7934 (N_7934,N_3557,N_3176);
xnor U7935 (N_7935,N_3715,N_3222);
nand U7936 (N_7936,N_4836,N_3778);
nor U7937 (N_7937,N_3776,N_5148);
nand U7938 (N_7938,N_4408,N_3276);
nor U7939 (N_7939,N_4465,N_3338);
nand U7940 (N_7940,N_4084,N_4326);
or U7941 (N_7941,N_4783,N_4662);
or U7942 (N_7942,N_3783,N_4560);
and U7943 (N_7943,N_5114,N_5992);
and U7944 (N_7944,N_4639,N_5512);
or U7945 (N_7945,N_4902,N_4949);
nor U7946 (N_7946,N_5345,N_4009);
nor U7947 (N_7947,N_5539,N_5627);
nor U7948 (N_7948,N_4117,N_4573);
and U7949 (N_7949,N_3288,N_3888);
and U7950 (N_7950,N_5297,N_4735);
xor U7951 (N_7951,N_3794,N_5178);
nand U7952 (N_7952,N_3049,N_3746);
xnor U7953 (N_7953,N_3540,N_4935);
nand U7954 (N_7954,N_3358,N_3123);
nand U7955 (N_7955,N_5888,N_5791);
and U7956 (N_7956,N_4742,N_5638);
or U7957 (N_7957,N_5565,N_3418);
nand U7958 (N_7958,N_4564,N_4988);
and U7959 (N_7959,N_5930,N_5034);
nor U7960 (N_7960,N_5435,N_3034);
nor U7961 (N_7961,N_3462,N_3949);
nand U7962 (N_7962,N_4107,N_4629);
nand U7963 (N_7963,N_5094,N_3673);
nand U7964 (N_7964,N_5646,N_5297);
nor U7965 (N_7965,N_3983,N_4568);
nand U7966 (N_7966,N_3725,N_5615);
xor U7967 (N_7967,N_4376,N_5340);
nand U7968 (N_7968,N_5984,N_3051);
nor U7969 (N_7969,N_5543,N_3842);
and U7970 (N_7970,N_3207,N_3628);
and U7971 (N_7971,N_4259,N_5681);
xor U7972 (N_7972,N_3732,N_5507);
or U7973 (N_7973,N_5151,N_5059);
and U7974 (N_7974,N_4505,N_3387);
xnor U7975 (N_7975,N_3959,N_4459);
xnor U7976 (N_7976,N_4170,N_5760);
nand U7977 (N_7977,N_5090,N_3110);
and U7978 (N_7978,N_4829,N_4238);
nor U7979 (N_7979,N_3689,N_3356);
xor U7980 (N_7980,N_5632,N_3074);
nor U7981 (N_7981,N_3728,N_4355);
nand U7982 (N_7982,N_3196,N_3050);
or U7983 (N_7983,N_4451,N_4619);
or U7984 (N_7984,N_3634,N_5441);
nand U7985 (N_7985,N_4253,N_3545);
and U7986 (N_7986,N_5113,N_4797);
nor U7987 (N_7987,N_4064,N_5858);
and U7988 (N_7988,N_4724,N_4438);
nand U7989 (N_7989,N_4977,N_5035);
xnor U7990 (N_7990,N_5712,N_5627);
nor U7991 (N_7991,N_3457,N_4379);
nor U7992 (N_7992,N_4561,N_5292);
xnor U7993 (N_7993,N_5029,N_4220);
xor U7994 (N_7994,N_4291,N_4976);
and U7995 (N_7995,N_5896,N_4493);
xor U7996 (N_7996,N_5592,N_3012);
nand U7997 (N_7997,N_5731,N_5335);
or U7998 (N_7998,N_5517,N_5428);
and U7999 (N_7999,N_4415,N_4932);
nand U8000 (N_8000,N_4023,N_5275);
xor U8001 (N_8001,N_4320,N_3951);
xor U8002 (N_8002,N_5766,N_3524);
or U8003 (N_8003,N_4277,N_4310);
or U8004 (N_8004,N_5164,N_5014);
and U8005 (N_8005,N_5727,N_4467);
nor U8006 (N_8006,N_4978,N_5478);
xnor U8007 (N_8007,N_3267,N_4498);
nand U8008 (N_8008,N_5571,N_3267);
xor U8009 (N_8009,N_4191,N_5133);
nor U8010 (N_8010,N_5211,N_4641);
or U8011 (N_8011,N_3435,N_4504);
nor U8012 (N_8012,N_4809,N_5079);
nand U8013 (N_8013,N_4188,N_4382);
xnor U8014 (N_8014,N_4858,N_4686);
or U8015 (N_8015,N_3142,N_4745);
or U8016 (N_8016,N_3814,N_3954);
nand U8017 (N_8017,N_5892,N_4818);
nand U8018 (N_8018,N_5904,N_5135);
nand U8019 (N_8019,N_3837,N_3657);
nand U8020 (N_8020,N_3264,N_3488);
nor U8021 (N_8021,N_4800,N_3961);
or U8022 (N_8022,N_5414,N_5805);
and U8023 (N_8023,N_4682,N_3097);
xnor U8024 (N_8024,N_4434,N_5162);
xnor U8025 (N_8025,N_5074,N_3716);
nor U8026 (N_8026,N_3796,N_4861);
nor U8027 (N_8027,N_4286,N_3766);
xnor U8028 (N_8028,N_4846,N_5891);
or U8029 (N_8029,N_5983,N_3940);
nand U8030 (N_8030,N_3914,N_5493);
xor U8031 (N_8031,N_3487,N_4863);
or U8032 (N_8032,N_3586,N_5443);
nor U8033 (N_8033,N_5742,N_3292);
and U8034 (N_8034,N_5676,N_3663);
nand U8035 (N_8035,N_4427,N_5947);
nor U8036 (N_8036,N_4706,N_5686);
and U8037 (N_8037,N_4059,N_3362);
nand U8038 (N_8038,N_4668,N_4785);
nor U8039 (N_8039,N_4841,N_5534);
xor U8040 (N_8040,N_5677,N_4933);
xor U8041 (N_8041,N_3785,N_3541);
nor U8042 (N_8042,N_3573,N_4254);
nor U8043 (N_8043,N_4926,N_3390);
nand U8044 (N_8044,N_4848,N_4565);
and U8045 (N_8045,N_4352,N_5420);
or U8046 (N_8046,N_5949,N_3810);
nand U8047 (N_8047,N_3924,N_3649);
nand U8048 (N_8048,N_5500,N_5184);
and U8049 (N_8049,N_3699,N_5429);
or U8050 (N_8050,N_3328,N_4763);
nor U8051 (N_8051,N_5697,N_3264);
or U8052 (N_8052,N_5244,N_5885);
or U8053 (N_8053,N_3270,N_3632);
nor U8054 (N_8054,N_5780,N_3344);
nand U8055 (N_8055,N_5465,N_3248);
nand U8056 (N_8056,N_3228,N_5816);
nand U8057 (N_8057,N_3087,N_5809);
nand U8058 (N_8058,N_3709,N_3034);
nand U8059 (N_8059,N_5252,N_3436);
nor U8060 (N_8060,N_3871,N_5063);
or U8061 (N_8061,N_3144,N_4770);
and U8062 (N_8062,N_5293,N_5205);
or U8063 (N_8063,N_5322,N_4825);
nor U8064 (N_8064,N_4257,N_5388);
xnor U8065 (N_8065,N_5463,N_3796);
or U8066 (N_8066,N_4143,N_3664);
nand U8067 (N_8067,N_4311,N_4594);
xnor U8068 (N_8068,N_5740,N_5364);
xor U8069 (N_8069,N_3026,N_5258);
nor U8070 (N_8070,N_4992,N_3746);
or U8071 (N_8071,N_4474,N_5907);
nor U8072 (N_8072,N_4187,N_5756);
xnor U8073 (N_8073,N_4249,N_3365);
and U8074 (N_8074,N_4909,N_5192);
and U8075 (N_8075,N_3725,N_3155);
or U8076 (N_8076,N_5109,N_3914);
and U8077 (N_8077,N_3383,N_3824);
nand U8078 (N_8078,N_5365,N_4318);
xnor U8079 (N_8079,N_4909,N_3400);
or U8080 (N_8080,N_4020,N_4988);
or U8081 (N_8081,N_3477,N_4338);
nand U8082 (N_8082,N_4968,N_3707);
nand U8083 (N_8083,N_3515,N_3690);
nand U8084 (N_8084,N_3078,N_5051);
or U8085 (N_8085,N_4748,N_4365);
and U8086 (N_8086,N_3832,N_4789);
and U8087 (N_8087,N_5245,N_3661);
and U8088 (N_8088,N_4961,N_4484);
xnor U8089 (N_8089,N_5510,N_5173);
or U8090 (N_8090,N_3651,N_5204);
xor U8091 (N_8091,N_5143,N_5528);
xnor U8092 (N_8092,N_5240,N_4558);
and U8093 (N_8093,N_3058,N_5886);
xnor U8094 (N_8094,N_5947,N_4113);
nor U8095 (N_8095,N_3625,N_4480);
nand U8096 (N_8096,N_5816,N_4730);
nand U8097 (N_8097,N_4598,N_5321);
xor U8098 (N_8098,N_4661,N_4363);
xor U8099 (N_8099,N_4940,N_3932);
xor U8100 (N_8100,N_5581,N_5724);
or U8101 (N_8101,N_3662,N_5998);
nor U8102 (N_8102,N_3552,N_3920);
xor U8103 (N_8103,N_5486,N_5267);
xor U8104 (N_8104,N_3295,N_4189);
and U8105 (N_8105,N_4321,N_3975);
or U8106 (N_8106,N_3105,N_3780);
or U8107 (N_8107,N_4180,N_4185);
and U8108 (N_8108,N_3005,N_3557);
or U8109 (N_8109,N_4407,N_3264);
and U8110 (N_8110,N_3113,N_5788);
nor U8111 (N_8111,N_3612,N_4801);
xor U8112 (N_8112,N_5001,N_4016);
nand U8113 (N_8113,N_4278,N_5656);
nor U8114 (N_8114,N_3911,N_3806);
nand U8115 (N_8115,N_5211,N_5055);
and U8116 (N_8116,N_4537,N_5110);
or U8117 (N_8117,N_5649,N_4276);
nor U8118 (N_8118,N_3166,N_4959);
nor U8119 (N_8119,N_4742,N_5946);
nor U8120 (N_8120,N_3638,N_5725);
xnor U8121 (N_8121,N_5122,N_4018);
nand U8122 (N_8122,N_4938,N_4411);
nand U8123 (N_8123,N_3903,N_5157);
nor U8124 (N_8124,N_3358,N_4132);
and U8125 (N_8125,N_3831,N_5041);
nor U8126 (N_8126,N_3533,N_3829);
and U8127 (N_8127,N_5551,N_4092);
nor U8128 (N_8128,N_4973,N_4625);
xor U8129 (N_8129,N_4262,N_3186);
and U8130 (N_8130,N_5612,N_3258);
or U8131 (N_8131,N_4419,N_5363);
or U8132 (N_8132,N_5916,N_5104);
nand U8133 (N_8133,N_5530,N_5795);
nor U8134 (N_8134,N_3497,N_5711);
and U8135 (N_8135,N_3734,N_5158);
and U8136 (N_8136,N_3326,N_5498);
nor U8137 (N_8137,N_3156,N_4146);
nand U8138 (N_8138,N_4781,N_5606);
or U8139 (N_8139,N_3668,N_3720);
xor U8140 (N_8140,N_5909,N_4114);
and U8141 (N_8141,N_3837,N_4570);
nand U8142 (N_8142,N_5315,N_3233);
and U8143 (N_8143,N_4605,N_5289);
nand U8144 (N_8144,N_5887,N_4708);
or U8145 (N_8145,N_5106,N_5187);
or U8146 (N_8146,N_4922,N_4768);
nor U8147 (N_8147,N_5043,N_5116);
xnor U8148 (N_8148,N_3767,N_4605);
nor U8149 (N_8149,N_4969,N_3975);
nor U8150 (N_8150,N_3539,N_5941);
xor U8151 (N_8151,N_4228,N_3324);
or U8152 (N_8152,N_3955,N_5418);
or U8153 (N_8153,N_3512,N_4766);
and U8154 (N_8154,N_4654,N_4289);
and U8155 (N_8155,N_4396,N_4908);
or U8156 (N_8156,N_3506,N_3252);
xnor U8157 (N_8157,N_5165,N_5869);
and U8158 (N_8158,N_4825,N_5059);
nor U8159 (N_8159,N_5878,N_4108);
nand U8160 (N_8160,N_3566,N_3848);
xor U8161 (N_8161,N_4909,N_5172);
or U8162 (N_8162,N_4909,N_4887);
xor U8163 (N_8163,N_3433,N_5777);
or U8164 (N_8164,N_5183,N_5625);
xnor U8165 (N_8165,N_5500,N_3377);
nand U8166 (N_8166,N_5602,N_3220);
nand U8167 (N_8167,N_3396,N_3206);
nor U8168 (N_8168,N_4541,N_3174);
nand U8169 (N_8169,N_4199,N_5776);
nor U8170 (N_8170,N_3913,N_5752);
or U8171 (N_8171,N_5820,N_5573);
xnor U8172 (N_8172,N_5974,N_4838);
and U8173 (N_8173,N_5834,N_3952);
and U8174 (N_8174,N_3311,N_3787);
or U8175 (N_8175,N_4970,N_3407);
xnor U8176 (N_8176,N_3773,N_5707);
xnor U8177 (N_8177,N_3770,N_5188);
xnor U8178 (N_8178,N_4691,N_4872);
and U8179 (N_8179,N_3540,N_3849);
and U8180 (N_8180,N_5084,N_4072);
and U8181 (N_8181,N_4816,N_4087);
and U8182 (N_8182,N_5097,N_5961);
nor U8183 (N_8183,N_5258,N_5800);
xnor U8184 (N_8184,N_5666,N_4195);
nor U8185 (N_8185,N_5254,N_3226);
nor U8186 (N_8186,N_4639,N_3475);
nand U8187 (N_8187,N_3160,N_3416);
and U8188 (N_8188,N_3123,N_3656);
xor U8189 (N_8189,N_5473,N_4484);
nor U8190 (N_8190,N_5410,N_5135);
or U8191 (N_8191,N_5797,N_4132);
or U8192 (N_8192,N_3847,N_4912);
or U8193 (N_8193,N_4224,N_5146);
and U8194 (N_8194,N_5575,N_3422);
or U8195 (N_8195,N_5801,N_4781);
nand U8196 (N_8196,N_5985,N_5097);
nand U8197 (N_8197,N_4162,N_5435);
nor U8198 (N_8198,N_5327,N_3094);
nor U8199 (N_8199,N_4349,N_4506);
and U8200 (N_8200,N_5633,N_5082);
and U8201 (N_8201,N_5670,N_3268);
or U8202 (N_8202,N_4249,N_3816);
or U8203 (N_8203,N_4324,N_5371);
xor U8204 (N_8204,N_3634,N_5035);
and U8205 (N_8205,N_4577,N_3616);
or U8206 (N_8206,N_4956,N_3645);
or U8207 (N_8207,N_4791,N_4572);
nor U8208 (N_8208,N_5684,N_5139);
or U8209 (N_8209,N_3842,N_3414);
or U8210 (N_8210,N_5248,N_4304);
xnor U8211 (N_8211,N_3791,N_4296);
and U8212 (N_8212,N_4400,N_5816);
xor U8213 (N_8213,N_3049,N_5223);
nor U8214 (N_8214,N_5201,N_5018);
or U8215 (N_8215,N_3275,N_4149);
nand U8216 (N_8216,N_3488,N_4847);
nor U8217 (N_8217,N_3441,N_4708);
or U8218 (N_8218,N_4377,N_3014);
nand U8219 (N_8219,N_3515,N_5446);
nor U8220 (N_8220,N_4698,N_4835);
or U8221 (N_8221,N_5278,N_3130);
and U8222 (N_8222,N_4780,N_5690);
nor U8223 (N_8223,N_4344,N_4249);
and U8224 (N_8224,N_5963,N_3984);
nand U8225 (N_8225,N_5633,N_3656);
or U8226 (N_8226,N_4066,N_5034);
or U8227 (N_8227,N_5281,N_5272);
and U8228 (N_8228,N_5268,N_5690);
nor U8229 (N_8229,N_5927,N_3095);
and U8230 (N_8230,N_4900,N_4190);
xnor U8231 (N_8231,N_4547,N_3009);
and U8232 (N_8232,N_4819,N_4696);
xnor U8233 (N_8233,N_5497,N_3975);
xnor U8234 (N_8234,N_4009,N_5273);
xnor U8235 (N_8235,N_3140,N_4055);
nand U8236 (N_8236,N_4387,N_4571);
xor U8237 (N_8237,N_3913,N_3121);
xor U8238 (N_8238,N_5875,N_3297);
and U8239 (N_8239,N_3885,N_4119);
and U8240 (N_8240,N_3880,N_4237);
nand U8241 (N_8241,N_3142,N_3866);
and U8242 (N_8242,N_4967,N_4529);
and U8243 (N_8243,N_4490,N_4562);
xnor U8244 (N_8244,N_3983,N_4821);
nand U8245 (N_8245,N_4140,N_4539);
nor U8246 (N_8246,N_4406,N_4812);
or U8247 (N_8247,N_3774,N_5591);
nor U8248 (N_8248,N_3906,N_4762);
and U8249 (N_8249,N_4469,N_5618);
xnor U8250 (N_8250,N_3101,N_3004);
and U8251 (N_8251,N_5440,N_3813);
xnor U8252 (N_8252,N_5250,N_5310);
nor U8253 (N_8253,N_5595,N_4104);
and U8254 (N_8254,N_3763,N_4414);
and U8255 (N_8255,N_5773,N_5165);
nor U8256 (N_8256,N_3341,N_5728);
and U8257 (N_8257,N_4837,N_3694);
and U8258 (N_8258,N_3099,N_4934);
xnor U8259 (N_8259,N_3015,N_3214);
nand U8260 (N_8260,N_5174,N_5996);
nor U8261 (N_8261,N_5373,N_4960);
nor U8262 (N_8262,N_3807,N_5136);
or U8263 (N_8263,N_3026,N_4823);
and U8264 (N_8264,N_4690,N_4149);
nand U8265 (N_8265,N_3418,N_5253);
and U8266 (N_8266,N_4688,N_3045);
xnor U8267 (N_8267,N_5757,N_4009);
xor U8268 (N_8268,N_4288,N_3495);
nand U8269 (N_8269,N_4411,N_5113);
or U8270 (N_8270,N_5982,N_4727);
nor U8271 (N_8271,N_4571,N_5373);
nand U8272 (N_8272,N_3380,N_3781);
or U8273 (N_8273,N_3487,N_3515);
and U8274 (N_8274,N_3668,N_4629);
or U8275 (N_8275,N_5785,N_4977);
xor U8276 (N_8276,N_4489,N_4281);
xor U8277 (N_8277,N_3778,N_3268);
nand U8278 (N_8278,N_5098,N_4266);
or U8279 (N_8279,N_4255,N_4793);
or U8280 (N_8280,N_4308,N_5136);
nand U8281 (N_8281,N_3721,N_3237);
and U8282 (N_8282,N_4925,N_3422);
and U8283 (N_8283,N_4889,N_5213);
nand U8284 (N_8284,N_4571,N_3363);
nor U8285 (N_8285,N_5742,N_3106);
nor U8286 (N_8286,N_4812,N_3010);
nand U8287 (N_8287,N_4536,N_3988);
xnor U8288 (N_8288,N_4336,N_4153);
nor U8289 (N_8289,N_4296,N_4845);
nor U8290 (N_8290,N_4971,N_3391);
and U8291 (N_8291,N_3656,N_5532);
and U8292 (N_8292,N_4927,N_3395);
nand U8293 (N_8293,N_5221,N_3803);
nand U8294 (N_8294,N_4806,N_4396);
xnor U8295 (N_8295,N_4880,N_3138);
and U8296 (N_8296,N_4791,N_4858);
nor U8297 (N_8297,N_4188,N_5294);
xnor U8298 (N_8298,N_4588,N_4946);
and U8299 (N_8299,N_5238,N_5562);
xor U8300 (N_8300,N_5886,N_5323);
and U8301 (N_8301,N_4812,N_3852);
xnor U8302 (N_8302,N_5846,N_4278);
xnor U8303 (N_8303,N_5929,N_5998);
nand U8304 (N_8304,N_5818,N_3496);
or U8305 (N_8305,N_3392,N_3723);
nor U8306 (N_8306,N_5823,N_5398);
and U8307 (N_8307,N_5397,N_4826);
nor U8308 (N_8308,N_3849,N_4068);
or U8309 (N_8309,N_4258,N_4329);
nand U8310 (N_8310,N_5803,N_5404);
xnor U8311 (N_8311,N_4387,N_5692);
nor U8312 (N_8312,N_3578,N_3662);
or U8313 (N_8313,N_4226,N_4153);
and U8314 (N_8314,N_4341,N_4011);
and U8315 (N_8315,N_4492,N_4974);
nand U8316 (N_8316,N_3315,N_3750);
and U8317 (N_8317,N_5245,N_5526);
and U8318 (N_8318,N_5191,N_5808);
or U8319 (N_8319,N_4376,N_3581);
and U8320 (N_8320,N_5356,N_3414);
nor U8321 (N_8321,N_4355,N_5491);
or U8322 (N_8322,N_5112,N_5295);
xnor U8323 (N_8323,N_5347,N_5220);
nand U8324 (N_8324,N_3836,N_4713);
and U8325 (N_8325,N_5258,N_5050);
xor U8326 (N_8326,N_4523,N_4290);
xnor U8327 (N_8327,N_3357,N_4611);
and U8328 (N_8328,N_3755,N_5340);
xor U8329 (N_8329,N_3061,N_5516);
or U8330 (N_8330,N_3896,N_3736);
and U8331 (N_8331,N_5866,N_4015);
nand U8332 (N_8332,N_4099,N_5090);
xnor U8333 (N_8333,N_5328,N_3714);
or U8334 (N_8334,N_4584,N_5577);
nor U8335 (N_8335,N_5301,N_5587);
nand U8336 (N_8336,N_4656,N_3715);
and U8337 (N_8337,N_3774,N_3721);
nand U8338 (N_8338,N_5254,N_4174);
nor U8339 (N_8339,N_3879,N_5326);
and U8340 (N_8340,N_5768,N_4847);
or U8341 (N_8341,N_3621,N_3387);
nand U8342 (N_8342,N_4904,N_4242);
or U8343 (N_8343,N_4824,N_4544);
nand U8344 (N_8344,N_4336,N_4474);
and U8345 (N_8345,N_5373,N_5372);
nand U8346 (N_8346,N_3009,N_3989);
and U8347 (N_8347,N_3646,N_5299);
or U8348 (N_8348,N_5081,N_4322);
nor U8349 (N_8349,N_4060,N_5146);
and U8350 (N_8350,N_5383,N_5296);
nand U8351 (N_8351,N_3108,N_3543);
and U8352 (N_8352,N_5597,N_4983);
or U8353 (N_8353,N_5261,N_5325);
or U8354 (N_8354,N_4676,N_4482);
and U8355 (N_8355,N_3890,N_4012);
nor U8356 (N_8356,N_4627,N_4427);
nand U8357 (N_8357,N_5285,N_3341);
nand U8358 (N_8358,N_4972,N_4204);
or U8359 (N_8359,N_4221,N_3960);
nor U8360 (N_8360,N_3935,N_4052);
or U8361 (N_8361,N_5318,N_3978);
nand U8362 (N_8362,N_3880,N_4777);
nand U8363 (N_8363,N_5443,N_4238);
nand U8364 (N_8364,N_5566,N_4591);
and U8365 (N_8365,N_5236,N_5111);
xor U8366 (N_8366,N_5624,N_3761);
nor U8367 (N_8367,N_5121,N_4621);
xnor U8368 (N_8368,N_3434,N_4353);
or U8369 (N_8369,N_3349,N_4837);
and U8370 (N_8370,N_4110,N_4946);
or U8371 (N_8371,N_4217,N_5521);
nor U8372 (N_8372,N_5252,N_3219);
nand U8373 (N_8373,N_5305,N_4497);
nor U8374 (N_8374,N_3731,N_5013);
nand U8375 (N_8375,N_5478,N_3166);
nand U8376 (N_8376,N_3472,N_3364);
nand U8377 (N_8377,N_5805,N_3831);
nor U8378 (N_8378,N_5998,N_5000);
xor U8379 (N_8379,N_5440,N_3436);
nor U8380 (N_8380,N_3374,N_4727);
or U8381 (N_8381,N_3778,N_4783);
or U8382 (N_8382,N_4379,N_5402);
xor U8383 (N_8383,N_4407,N_5608);
nor U8384 (N_8384,N_3367,N_3502);
nor U8385 (N_8385,N_5699,N_4278);
and U8386 (N_8386,N_3838,N_4760);
nor U8387 (N_8387,N_4621,N_5740);
and U8388 (N_8388,N_4181,N_4582);
nand U8389 (N_8389,N_5419,N_4614);
nor U8390 (N_8390,N_4566,N_5999);
and U8391 (N_8391,N_4529,N_4405);
nand U8392 (N_8392,N_5898,N_5032);
and U8393 (N_8393,N_5933,N_5849);
or U8394 (N_8394,N_4264,N_4826);
or U8395 (N_8395,N_5555,N_3546);
nor U8396 (N_8396,N_5838,N_5646);
xor U8397 (N_8397,N_5923,N_3434);
or U8398 (N_8398,N_4957,N_3608);
nand U8399 (N_8399,N_3077,N_4590);
xnor U8400 (N_8400,N_4900,N_3307);
or U8401 (N_8401,N_3071,N_4163);
and U8402 (N_8402,N_5862,N_3459);
or U8403 (N_8403,N_5793,N_3840);
xor U8404 (N_8404,N_4782,N_4984);
or U8405 (N_8405,N_3090,N_5431);
or U8406 (N_8406,N_3542,N_4782);
nor U8407 (N_8407,N_4398,N_5717);
nand U8408 (N_8408,N_5384,N_4366);
or U8409 (N_8409,N_4195,N_5291);
and U8410 (N_8410,N_4447,N_4185);
nand U8411 (N_8411,N_4885,N_4232);
or U8412 (N_8412,N_3306,N_5900);
or U8413 (N_8413,N_4833,N_3416);
and U8414 (N_8414,N_3888,N_4916);
nor U8415 (N_8415,N_5268,N_3089);
and U8416 (N_8416,N_4991,N_4988);
nor U8417 (N_8417,N_3008,N_3022);
or U8418 (N_8418,N_4587,N_3786);
or U8419 (N_8419,N_5165,N_4647);
and U8420 (N_8420,N_3958,N_4228);
nand U8421 (N_8421,N_3142,N_3219);
and U8422 (N_8422,N_4511,N_5254);
or U8423 (N_8423,N_3294,N_4409);
xor U8424 (N_8424,N_5189,N_5984);
xor U8425 (N_8425,N_4567,N_5565);
or U8426 (N_8426,N_3641,N_3957);
nor U8427 (N_8427,N_4249,N_4967);
nand U8428 (N_8428,N_4766,N_5050);
or U8429 (N_8429,N_3401,N_4488);
and U8430 (N_8430,N_4638,N_4166);
nand U8431 (N_8431,N_5883,N_3761);
nand U8432 (N_8432,N_3496,N_4770);
nand U8433 (N_8433,N_3607,N_5482);
and U8434 (N_8434,N_5416,N_3090);
nand U8435 (N_8435,N_3444,N_3293);
nand U8436 (N_8436,N_5885,N_4964);
and U8437 (N_8437,N_5242,N_4056);
xnor U8438 (N_8438,N_3531,N_3288);
or U8439 (N_8439,N_3045,N_3166);
or U8440 (N_8440,N_5752,N_4191);
or U8441 (N_8441,N_3659,N_3284);
or U8442 (N_8442,N_3717,N_5350);
nor U8443 (N_8443,N_3132,N_5716);
xnor U8444 (N_8444,N_4026,N_5494);
and U8445 (N_8445,N_4106,N_5834);
and U8446 (N_8446,N_3133,N_4800);
xnor U8447 (N_8447,N_3854,N_5639);
nand U8448 (N_8448,N_4801,N_5653);
xor U8449 (N_8449,N_5752,N_5421);
and U8450 (N_8450,N_4372,N_5682);
nor U8451 (N_8451,N_4236,N_5338);
xnor U8452 (N_8452,N_3176,N_4242);
or U8453 (N_8453,N_5269,N_4017);
nand U8454 (N_8454,N_3785,N_3540);
or U8455 (N_8455,N_5114,N_5793);
nor U8456 (N_8456,N_4425,N_3860);
or U8457 (N_8457,N_3969,N_5425);
nor U8458 (N_8458,N_5869,N_5855);
nor U8459 (N_8459,N_3930,N_4056);
xnor U8460 (N_8460,N_5815,N_4452);
and U8461 (N_8461,N_3874,N_3269);
nor U8462 (N_8462,N_3118,N_4518);
and U8463 (N_8463,N_5823,N_5720);
nor U8464 (N_8464,N_4456,N_3214);
or U8465 (N_8465,N_3748,N_3212);
or U8466 (N_8466,N_5749,N_4843);
nand U8467 (N_8467,N_5627,N_4526);
and U8468 (N_8468,N_3485,N_5756);
nor U8469 (N_8469,N_5734,N_5652);
nor U8470 (N_8470,N_3317,N_3710);
nand U8471 (N_8471,N_5130,N_5334);
or U8472 (N_8472,N_5744,N_4791);
and U8473 (N_8473,N_4579,N_3264);
nand U8474 (N_8474,N_3954,N_3064);
nand U8475 (N_8475,N_5006,N_3260);
xnor U8476 (N_8476,N_4196,N_5985);
and U8477 (N_8477,N_4233,N_5668);
xnor U8478 (N_8478,N_4262,N_5606);
and U8479 (N_8479,N_3379,N_5482);
nor U8480 (N_8480,N_4201,N_4259);
nand U8481 (N_8481,N_4597,N_4519);
xnor U8482 (N_8482,N_5065,N_3706);
or U8483 (N_8483,N_4377,N_4872);
nor U8484 (N_8484,N_5154,N_5265);
nor U8485 (N_8485,N_5353,N_3056);
or U8486 (N_8486,N_5315,N_5336);
nand U8487 (N_8487,N_4203,N_4103);
or U8488 (N_8488,N_5022,N_5371);
nor U8489 (N_8489,N_3280,N_4736);
xor U8490 (N_8490,N_3210,N_3983);
nand U8491 (N_8491,N_4375,N_4130);
and U8492 (N_8492,N_3098,N_5808);
or U8493 (N_8493,N_3408,N_4167);
xor U8494 (N_8494,N_3772,N_5706);
nor U8495 (N_8495,N_4607,N_5716);
and U8496 (N_8496,N_4229,N_4512);
xnor U8497 (N_8497,N_3688,N_5849);
xor U8498 (N_8498,N_3387,N_5348);
xnor U8499 (N_8499,N_3539,N_3242);
and U8500 (N_8500,N_5975,N_5433);
nor U8501 (N_8501,N_3335,N_4369);
or U8502 (N_8502,N_5203,N_3960);
nand U8503 (N_8503,N_3874,N_5656);
nor U8504 (N_8504,N_5692,N_4719);
nand U8505 (N_8505,N_4162,N_4576);
nor U8506 (N_8506,N_3004,N_5658);
or U8507 (N_8507,N_5443,N_5406);
xor U8508 (N_8508,N_3722,N_5909);
nor U8509 (N_8509,N_4556,N_3836);
nand U8510 (N_8510,N_3626,N_3290);
xor U8511 (N_8511,N_5004,N_5862);
or U8512 (N_8512,N_3291,N_4053);
nand U8513 (N_8513,N_4658,N_4341);
or U8514 (N_8514,N_5721,N_3165);
or U8515 (N_8515,N_4625,N_3875);
nand U8516 (N_8516,N_3784,N_3128);
nor U8517 (N_8517,N_5703,N_4819);
nor U8518 (N_8518,N_3937,N_5038);
xor U8519 (N_8519,N_5072,N_4098);
or U8520 (N_8520,N_4237,N_3783);
nand U8521 (N_8521,N_5478,N_5274);
nor U8522 (N_8522,N_5115,N_3728);
nor U8523 (N_8523,N_5392,N_5935);
or U8524 (N_8524,N_4283,N_4963);
xor U8525 (N_8525,N_3592,N_3296);
nor U8526 (N_8526,N_4174,N_3750);
xor U8527 (N_8527,N_5532,N_3718);
xnor U8528 (N_8528,N_5047,N_4541);
nor U8529 (N_8529,N_4185,N_3192);
nor U8530 (N_8530,N_4770,N_5041);
nor U8531 (N_8531,N_4648,N_3719);
xnor U8532 (N_8532,N_5990,N_3772);
or U8533 (N_8533,N_4913,N_4380);
nand U8534 (N_8534,N_3974,N_4475);
nor U8535 (N_8535,N_3227,N_4958);
xnor U8536 (N_8536,N_4313,N_3515);
or U8537 (N_8537,N_4889,N_5845);
nor U8538 (N_8538,N_5031,N_4259);
or U8539 (N_8539,N_4064,N_5675);
nor U8540 (N_8540,N_5534,N_4955);
nand U8541 (N_8541,N_5370,N_4682);
or U8542 (N_8542,N_3390,N_4552);
and U8543 (N_8543,N_3560,N_5654);
nor U8544 (N_8544,N_3677,N_5292);
xor U8545 (N_8545,N_4096,N_4793);
xor U8546 (N_8546,N_5277,N_4403);
nand U8547 (N_8547,N_4984,N_5147);
or U8548 (N_8548,N_4841,N_3822);
nand U8549 (N_8549,N_3076,N_5617);
nor U8550 (N_8550,N_5796,N_5973);
xor U8551 (N_8551,N_3184,N_4253);
nor U8552 (N_8552,N_3368,N_5843);
nand U8553 (N_8553,N_5788,N_5981);
or U8554 (N_8554,N_3945,N_4154);
xor U8555 (N_8555,N_4339,N_3976);
or U8556 (N_8556,N_4970,N_3738);
nand U8557 (N_8557,N_4314,N_5379);
and U8558 (N_8558,N_3669,N_5771);
and U8559 (N_8559,N_3126,N_3540);
nand U8560 (N_8560,N_3569,N_4262);
xnor U8561 (N_8561,N_5683,N_5210);
and U8562 (N_8562,N_5036,N_5978);
or U8563 (N_8563,N_4577,N_5570);
and U8564 (N_8564,N_3949,N_5883);
or U8565 (N_8565,N_4484,N_4912);
and U8566 (N_8566,N_5721,N_4064);
or U8567 (N_8567,N_4768,N_3801);
and U8568 (N_8568,N_4545,N_5044);
nor U8569 (N_8569,N_5800,N_4450);
and U8570 (N_8570,N_4346,N_3744);
nand U8571 (N_8571,N_5877,N_5848);
nor U8572 (N_8572,N_3696,N_3480);
or U8573 (N_8573,N_3809,N_3301);
and U8574 (N_8574,N_3033,N_4465);
or U8575 (N_8575,N_3616,N_4717);
xor U8576 (N_8576,N_4604,N_4740);
or U8577 (N_8577,N_3079,N_3683);
nand U8578 (N_8578,N_3826,N_5258);
and U8579 (N_8579,N_3193,N_5094);
and U8580 (N_8580,N_4174,N_4451);
nor U8581 (N_8581,N_4014,N_5693);
or U8582 (N_8582,N_3907,N_3668);
or U8583 (N_8583,N_5947,N_3123);
nor U8584 (N_8584,N_3216,N_5560);
nand U8585 (N_8585,N_4212,N_5144);
and U8586 (N_8586,N_3212,N_5911);
or U8587 (N_8587,N_3298,N_3792);
nor U8588 (N_8588,N_3813,N_5061);
xnor U8589 (N_8589,N_3404,N_5265);
and U8590 (N_8590,N_3030,N_5752);
xor U8591 (N_8591,N_3898,N_3759);
or U8592 (N_8592,N_4240,N_3120);
nand U8593 (N_8593,N_3420,N_4462);
xor U8594 (N_8594,N_3685,N_3932);
and U8595 (N_8595,N_5972,N_3722);
and U8596 (N_8596,N_5716,N_3554);
nand U8597 (N_8597,N_4983,N_4122);
or U8598 (N_8598,N_3129,N_5646);
nand U8599 (N_8599,N_5088,N_3463);
and U8600 (N_8600,N_4451,N_5082);
nor U8601 (N_8601,N_4704,N_5156);
and U8602 (N_8602,N_4477,N_3328);
and U8603 (N_8603,N_3034,N_5176);
or U8604 (N_8604,N_3077,N_5163);
nand U8605 (N_8605,N_4562,N_3783);
xor U8606 (N_8606,N_3623,N_5367);
xor U8607 (N_8607,N_5762,N_4429);
or U8608 (N_8608,N_4825,N_5421);
xnor U8609 (N_8609,N_3744,N_5669);
or U8610 (N_8610,N_5459,N_4209);
nand U8611 (N_8611,N_5689,N_5099);
nor U8612 (N_8612,N_5314,N_5282);
nand U8613 (N_8613,N_4561,N_3001);
nor U8614 (N_8614,N_3365,N_3499);
and U8615 (N_8615,N_4692,N_5270);
and U8616 (N_8616,N_5048,N_5240);
xnor U8617 (N_8617,N_5416,N_3754);
nor U8618 (N_8618,N_3515,N_3043);
nor U8619 (N_8619,N_5382,N_5366);
or U8620 (N_8620,N_3388,N_4787);
nor U8621 (N_8621,N_4247,N_4565);
and U8622 (N_8622,N_3614,N_4694);
nor U8623 (N_8623,N_5721,N_5667);
xor U8624 (N_8624,N_3370,N_5799);
nor U8625 (N_8625,N_4957,N_5693);
nand U8626 (N_8626,N_5830,N_5835);
or U8627 (N_8627,N_4589,N_3026);
nand U8628 (N_8628,N_5629,N_3578);
xor U8629 (N_8629,N_4577,N_4215);
and U8630 (N_8630,N_5479,N_5075);
or U8631 (N_8631,N_4352,N_4744);
nand U8632 (N_8632,N_4390,N_5604);
and U8633 (N_8633,N_3831,N_4561);
nand U8634 (N_8634,N_4517,N_3257);
or U8635 (N_8635,N_4310,N_5806);
xnor U8636 (N_8636,N_3002,N_5534);
xnor U8637 (N_8637,N_4159,N_3105);
xnor U8638 (N_8638,N_3095,N_5431);
and U8639 (N_8639,N_4031,N_4523);
and U8640 (N_8640,N_4108,N_3314);
or U8641 (N_8641,N_3191,N_4305);
and U8642 (N_8642,N_3645,N_4350);
or U8643 (N_8643,N_5515,N_4665);
nand U8644 (N_8644,N_5032,N_4414);
or U8645 (N_8645,N_5455,N_3557);
xnor U8646 (N_8646,N_4548,N_4054);
or U8647 (N_8647,N_5063,N_5358);
or U8648 (N_8648,N_3724,N_4135);
nor U8649 (N_8649,N_3652,N_5997);
or U8650 (N_8650,N_3913,N_3884);
nand U8651 (N_8651,N_4188,N_4640);
nor U8652 (N_8652,N_4752,N_3908);
nor U8653 (N_8653,N_5833,N_3820);
or U8654 (N_8654,N_4924,N_3143);
xnor U8655 (N_8655,N_4108,N_5831);
nor U8656 (N_8656,N_3673,N_4356);
nor U8657 (N_8657,N_3775,N_4544);
xor U8658 (N_8658,N_5662,N_3258);
nor U8659 (N_8659,N_4930,N_5927);
xnor U8660 (N_8660,N_5858,N_4845);
nor U8661 (N_8661,N_5311,N_4087);
nand U8662 (N_8662,N_3715,N_3099);
or U8663 (N_8663,N_5095,N_4757);
nand U8664 (N_8664,N_5141,N_4114);
and U8665 (N_8665,N_4837,N_4373);
and U8666 (N_8666,N_5869,N_4214);
nand U8667 (N_8667,N_4933,N_4031);
or U8668 (N_8668,N_3191,N_3461);
nor U8669 (N_8669,N_5408,N_5853);
and U8670 (N_8670,N_5881,N_4778);
and U8671 (N_8671,N_4739,N_5934);
or U8672 (N_8672,N_5133,N_4773);
or U8673 (N_8673,N_5246,N_4215);
and U8674 (N_8674,N_5496,N_3932);
or U8675 (N_8675,N_5109,N_3090);
xor U8676 (N_8676,N_5614,N_3182);
or U8677 (N_8677,N_5107,N_4089);
and U8678 (N_8678,N_3743,N_5370);
xor U8679 (N_8679,N_5466,N_4085);
nor U8680 (N_8680,N_5294,N_4085);
and U8681 (N_8681,N_3928,N_3517);
or U8682 (N_8682,N_3455,N_3288);
or U8683 (N_8683,N_3854,N_5698);
and U8684 (N_8684,N_5344,N_3982);
and U8685 (N_8685,N_3470,N_3893);
nand U8686 (N_8686,N_5933,N_4958);
xnor U8687 (N_8687,N_3288,N_5391);
xnor U8688 (N_8688,N_3347,N_5474);
nor U8689 (N_8689,N_5686,N_3595);
and U8690 (N_8690,N_4183,N_4671);
nor U8691 (N_8691,N_3928,N_4646);
xnor U8692 (N_8692,N_4264,N_3016);
nand U8693 (N_8693,N_3401,N_4737);
or U8694 (N_8694,N_4074,N_4965);
nand U8695 (N_8695,N_4767,N_3014);
or U8696 (N_8696,N_3743,N_4850);
or U8697 (N_8697,N_5950,N_4319);
xnor U8698 (N_8698,N_5844,N_4898);
nor U8699 (N_8699,N_5909,N_3312);
or U8700 (N_8700,N_5848,N_3654);
and U8701 (N_8701,N_3357,N_3540);
nand U8702 (N_8702,N_4953,N_5542);
and U8703 (N_8703,N_5951,N_5995);
nand U8704 (N_8704,N_4780,N_4121);
nand U8705 (N_8705,N_5350,N_3930);
and U8706 (N_8706,N_3430,N_3196);
nand U8707 (N_8707,N_5545,N_3166);
or U8708 (N_8708,N_3604,N_5535);
xnor U8709 (N_8709,N_5408,N_4675);
nor U8710 (N_8710,N_5397,N_5390);
xnor U8711 (N_8711,N_4659,N_5515);
or U8712 (N_8712,N_5604,N_5294);
xnor U8713 (N_8713,N_3753,N_3183);
and U8714 (N_8714,N_5793,N_3468);
xor U8715 (N_8715,N_4189,N_4014);
nand U8716 (N_8716,N_3413,N_4373);
nor U8717 (N_8717,N_5966,N_4191);
xor U8718 (N_8718,N_5147,N_3332);
nand U8719 (N_8719,N_3402,N_3385);
nor U8720 (N_8720,N_3646,N_3469);
xor U8721 (N_8721,N_4031,N_4833);
xor U8722 (N_8722,N_3268,N_5661);
nand U8723 (N_8723,N_3461,N_4871);
and U8724 (N_8724,N_5390,N_3386);
xor U8725 (N_8725,N_4103,N_4295);
xnor U8726 (N_8726,N_5672,N_5244);
nor U8727 (N_8727,N_4736,N_3997);
nor U8728 (N_8728,N_3193,N_3271);
xor U8729 (N_8729,N_4931,N_4847);
and U8730 (N_8730,N_4251,N_5365);
xnor U8731 (N_8731,N_4436,N_5454);
nor U8732 (N_8732,N_4964,N_3491);
nand U8733 (N_8733,N_4260,N_4902);
nor U8734 (N_8734,N_3015,N_3971);
xnor U8735 (N_8735,N_3649,N_3071);
nand U8736 (N_8736,N_3493,N_3292);
xor U8737 (N_8737,N_5433,N_3184);
nand U8738 (N_8738,N_3805,N_4854);
and U8739 (N_8739,N_5540,N_4084);
and U8740 (N_8740,N_5491,N_4268);
nor U8741 (N_8741,N_4639,N_5170);
xor U8742 (N_8742,N_3806,N_5161);
and U8743 (N_8743,N_3642,N_3358);
or U8744 (N_8744,N_5294,N_4939);
and U8745 (N_8745,N_4240,N_5592);
nor U8746 (N_8746,N_3309,N_5841);
xor U8747 (N_8747,N_4880,N_3333);
xnor U8748 (N_8748,N_4448,N_5481);
nor U8749 (N_8749,N_3099,N_4083);
xor U8750 (N_8750,N_3969,N_4379);
nand U8751 (N_8751,N_4480,N_5653);
nor U8752 (N_8752,N_3740,N_4836);
or U8753 (N_8753,N_4431,N_3487);
nor U8754 (N_8754,N_3329,N_3610);
xnor U8755 (N_8755,N_3285,N_5206);
xor U8756 (N_8756,N_3634,N_5791);
or U8757 (N_8757,N_3693,N_4686);
nand U8758 (N_8758,N_3566,N_5473);
nor U8759 (N_8759,N_3123,N_5198);
xor U8760 (N_8760,N_4201,N_5399);
and U8761 (N_8761,N_4241,N_4449);
xor U8762 (N_8762,N_5793,N_3061);
and U8763 (N_8763,N_4499,N_3420);
and U8764 (N_8764,N_5027,N_5098);
nand U8765 (N_8765,N_5594,N_5510);
or U8766 (N_8766,N_3220,N_5583);
or U8767 (N_8767,N_5601,N_3311);
or U8768 (N_8768,N_3299,N_5909);
nor U8769 (N_8769,N_5585,N_3197);
and U8770 (N_8770,N_3787,N_3432);
nor U8771 (N_8771,N_5037,N_3857);
nand U8772 (N_8772,N_5665,N_3676);
or U8773 (N_8773,N_4150,N_5406);
nand U8774 (N_8774,N_5465,N_4265);
nor U8775 (N_8775,N_5169,N_5549);
xor U8776 (N_8776,N_4901,N_3297);
and U8777 (N_8777,N_4734,N_4624);
nand U8778 (N_8778,N_3159,N_3794);
nand U8779 (N_8779,N_4922,N_5443);
nand U8780 (N_8780,N_3800,N_4080);
nand U8781 (N_8781,N_5157,N_5410);
and U8782 (N_8782,N_3423,N_5779);
or U8783 (N_8783,N_4547,N_3890);
or U8784 (N_8784,N_3922,N_4916);
nor U8785 (N_8785,N_5937,N_5860);
or U8786 (N_8786,N_3159,N_5450);
and U8787 (N_8787,N_4389,N_4595);
nor U8788 (N_8788,N_3780,N_5838);
xnor U8789 (N_8789,N_4913,N_4562);
nand U8790 (N_8790,N_3917,N_3447);
nand U8791 (N_8791,N_5016,N_4212);
nor U8792 (N_8792,N_3639,N_4115);
or U8793 (N_8793,N_3482,N_5671);
or U8794 (N_8794,N_3539,N_5986);
nor U8795 (N_8795,N_5991,N_3157);
and U8796 (N_8796,N_3360,N_4398);
nor U8797 (N_8797,N_3618,N_3600);
nor U8798 (N_8798,N_3998,N_5954);
nor U8799 (N_8799,N_3133,N_3819);
nor U8800 (N_8800,N_5381,N_4084);
nand U8801 (N_8801,N_5938,N_5787);
nor U8802 (N_8802,N_5687,N_5981);
or U8803 (N_8803,N_3894,N_4498);
nor U8804 (N_8804,N_4239,N_5273);
nand U8805 (N_8805,N_3506,N_4571);
xor U8806 (N_8806,N_3306,N_3425);
or U8807 (N_8807,N_4608,N_3476);
or U8808 (N_8808,N_5094,N_3389);
nor U8809 (N_8809,N_5112,N_3197);
or U8810 (N_8810,N_5529,N_3136);
nand U8811 (N_8811,N_3753,N_4268);
xor U8812 (N_8812,N_4261,N_5340);
and U8813 (N_8813,N_4318,N_4092);
nand U8814 (N_8814,N_3270,N_3398);
and U8815 (N_8815,N_4861,N_5071);
nor U8816 (N_8816,N_4927,N_4567);
or U8817 (N_8817,N_4324,N_5956);
and U8818 (N_8818,N_5662,N_5136);
nor U8819 (N_8819,N_4395,N_5401);
nor U8820 (N_8820,N_5692,N_5506);
xor U8821 (N_8821,N_4318,N_3357);
and U8822 (N_8822,N_5462,N_4024);
xnor U8823 (N_8823,N_3852,N_5674);
xor U8824 (N_8824,N_3651,N_4901);
or U8825 (N_8825,N_4893,N_3725);
and U8826 (N_8826,N_4717,N_3515);
xor U8827 (N_8827,N_5188,N_3304);
xor U8828 (N_8828,N_3186,N_4669);
xnor U8829 (N_8829,N_3471,N_5621);
and U8830 (N_8830,N_3797,N_3399);
nor U8831 (N_8831,N_5837,N_3462);
xnor U8832 (N_8832,N_3557,N_5973);
nor U8833 (N_8833,N_4462,N_3207);
nand U8834 (N_8834,N_4693,N_4356);
nor U8835 (N_8835,N_3193,N_4358);
nand U8836 (N_8836,N_5210,N_5620);
nand U8837 (N_8837,N_3987,N_4068);
or U8838 (N_8838,N_5215,N_3601);
and U8839 (N_8839,N_3053,N_5193);
or U8840 (N_8840,N_4431,N_3288);
nor U8841 (N_8841,N_4415,N_4116);
nand U8842 (N_8842,N_5321,N_4083);
or U8843 (N_8843,N_5695,N_4551);
nand U8844 (N_8844,N_3339,N_5423);
and U8845 (N_8845,N_5367,N_4506);
nor U8846 (N_8846,N_5320,N_3296);
or U8847 (N_8847,N_4907,N_3718);
nand U8848 (N_8848,N_5148,N_3824);
nand U8849 (N_8849,N_3600,N_3671);
xor U8850 (N_8850,N_5992,N_5013);
or U8851 (N_8851,N_4773,N_5355);
and U8852 (N_8852,N_3282,N_3156);
xor U8853 (N_8853,N_4032,N_4297);
nand U8854 (N_8854,N_4624,N_5683);
and U8855 (N_8855,N_5644,N_3956);
or U8856 (N_8856,N_3489,N_3924);
and U8857 (N_8857,N_3166,N_5537);
nor U8858 (N_8858,N_3820,N_3947);
nand U8859 (N_8859,N_5541,N_3748);
or U8860 (N_8860,N_5166,N_4746);
nand U8861 (N_8861,N_3490,N_4565);
nor U8862 (N_8862,N_5701,N_4656);
and U8863 (N_8863,N_4704,N_5975);
xor U8864 (N_8864,N_5585,N_5078);
nor U8865 (N_8865,N_4454,N_5140);
nor U8866 (N_8866,N_4899,N_5470);
or U8867 (N_8867,N_5656,N_3988);
xor U8868 (N_8868,N_5733,N_4611);
xnor U8869 (N_8869,N_5844,N_4042);
xnor U8870 (N_8870,N_4697,N_3399);
or U8871 (N_8871,N_3278,N_5177);
and U8872 (N_8872,N_5700,N_4237);
nand U8873 (N_8873,N_4233,N_3368);
and U8874 (N_8874,N_3757,N_3496);
and U8875 (N_8875,N_5986,N_4810);
nand U8876 (N_8876,N_4882,N_5237);
nand U8877 (N_8877,N_5042,N_4690);
and U8878 (N_8878,N_5424,N_3389);
xnor U8879 (N_8879,N_5321,N_5622);
or U8880 (N_8880,N_5518,N_3164);
nand U8881 (N_8881,N_4580,N_4295);
nor U8882 (N_8882,N_3014,N_5757);
or U8883 (N_8883,N_5858,N_5279);
nand U8884 (N_8884,N_3710,N_4715);
nor U8885 (N_8885,N_3666,N_5061);
or U8886 (N_8886,N_4524,N_5700);
and U8887 (N_8887,N_4324,N_4187);
and U8888 (N_8888,N_5377,N_3538);
or U8889 (N_8889,N_3420,N_3481);
or U8890 (N_8890,N_5372,N_3711);
nor U8891 (N_8891,N_5738,N_4362);
xnor U8892 (N_8892,N_5420,N_5196);
and U8893 (N_8893,N_4523,N_5993);
nand U8894 (N_8894,N_3173,N_4716);
nor U8895 (N_8895,N_4180,N_4049);
or U8896 (N_8896,N_4938,N_3246);
or U8897 (N_8897,N_5882,N_4884);
and U8898 (N_8898,N_5315,N_4415);
xnor U8899 (N_8899,N_4270,N_3486);
or U8900 (N_8900,N_5659,N_3145);
nor U8901 (N_8901,N_3209,N_5053);
xor U8902 (N_8902,N_3424,N_5538);
nand U8903 (N_8903,N_5181,N_4542);
xor U8904 (N_8904,N_5012,N_3978);
nand U8905 (N_8905,N_5887,N_3938);
and U8906 (N_8906,N_5459,N_5090);
xnor U8907 (N_8907,N_5583,N_5410);
nand U8908 (N_8908,N_5221,N_3721);
or U8909 (N_8909,N_4077,N_4933);
xor U8910 (N_8910,N_5945,N_5632);
nor U8911 (N_8911,N_5600,N_3951);
xnor U8912 (N_8912,N_3837,N_4355);
or U8913 (N_8913,N_4498,N_5839);
and U8914 (N_8914,N_4681,N_5602);
nor U8915 (N_8915,N_3510,N_4513);
and U8916 (N_8916,N_3960,N_5859);
nand U8917 (N_8917,N_4210,N_3069);
nor U8918 (N_8918,N_3081,N_3291);
or U8919 (N_8919,N_5418,N_4113);
and U8920 (N_8920,N_4942,N_4408);
nand U8921 (N_8921,N_3311,N_3559);
or U8922 (N_8922,N_5660,N_5250);
nand U8923 (N_8923,N_4965,N_5115);
xor U8924 (N_8924,N_4352,N_5957);
and U8925 (N_8925,N_4203,N_5710);
nand U8926 (N_8926,N_3604,N_3589);
nor U8927 (N_8927,N_4048,N_3408);
nand U8928 (N_8928,N_4472,N_5439);
or U8929 (N_8929,N_4773,N_3814);
nand U8930 (N_8930,N_5882,N_4958);
nand U8931 (N_8931,N_5174,N_5872);
nor U8932 (N_8932,N_3060,N_4370);
nor U8933 (N_8933,N_4910,N_3109);
nand U8934 (N_8934,N_4308,N_3222);
xnor U8935 (N_8935,N_4136,N_3744);
and U8936 (N_8936,N_3802,N_4836);
and U8937 (N_8937,N_4888,N_5811);
nor U8938 (N_8938,N_4873,N_3820);
nand U8939 (N_8939,N_4048,N_4153);
and U8940 (N_8940,N_5389,N_5308);
and U8941 (N_8941,N_4289,N_5056);
xor U8942 (N_8942,N_4420,N_5667);
xor U8943 (N_8943,N_4944,N_3562);
and U8944 (N_8944,N_3020,N_3387);
xor U8945 (N_8945,N_3685,N_3919);
xnor U8946 (N_8946,N_4113,N_3469);
and U8947 (N_8947,N_5952,N_3967);
and U8948 (N_8948,N_4927,N_4332);
or U8949 (N_8949,N_4738,N_4397);
xnor U8950 (N_8950,N_4965,N_4287);
nand U8951 (N_8951,N_4886,N_3598);
nor U8952 (N_8952,N_3883,N_5401);
and U8953 (N_8953,N_4972,N_5054);
xnor U8954 (N_8954,N_3212,N_5819);
or U8955 (N_8955,N_3232,N_5078);
and U8956 (N_8956,N_5984,N_5071);
nand U8957 (N_8957,N_5126,N_3656);
nor U8958 (N_8958,N_5630,N_3058);
nor U8959 (N_8959,N_3374,N_3802);
or U8960 (N_8960,N_3045,N_3161);
nor U8961 (N_8961,N_3399,N_3164);
and U8962 (N_8962,N_5918,N_3952);
or U8963 (N_8963,N_4975,N_3204);
xnor U8964 (N_8964,N_3454,N_4068);
xor U8965 (N_8965,N_5018,N_5652);
or U8966 (N_8966,N_5600,N_4632);
nor U8967 (N_8967,N_3818,N_5032);
xor U8968 (N_8968,N_4370,N_5069);
nor U8969 (N_8969,N_5767,N_3876);
nor U8970 (N_8970,N_3514,N_5752);
xnor U8971 (N_8971,N_3613,N_4172);
xnor U8972 (N_8972,N_4839,N_3843);
nor U8973 (N_8973,N_4343,N_3405);
nand U8974 (N_8974,N_3156,N_5009);
or U8975 (N_8975,N_4555,N_4553);
and U8976 (N_8976,N_4578,N_5433);
xnor U8977 (N_8977,N_4684,N_3468);
nor U8978 (N_8978,N_5730,N_3554);
nor U8979 (N_8979,N_3202,N_4152);
nor U8980 (N_8980,N_5382,N_4155);
xnor U8981 (N_8981,N_4361,N_3665);
nand U8982 (N_8982,N_5012,N_5937);
or U8983 (N_8983,N_3783,N_4510);
or U8984 (N_8984,N_3764,N_3873);
and U8985 (N_8985,N_4718,N_5790);
nor U8986 (N_8986,N_5215,N_3493);
nand U8987 (N_8987,N_3695,N_3395);
and U8988 (N_8988,N_4322,N_4406);
nor U8989 (N_8989,N_4266,N_3593);
nor U8990 (N_8990,N_5221,N_4833);
xor U8991 (N_8991,N_5967,N_5129);
nand U8992 (N_8992,N_5194,N_3758);
xor U8993 (N_8993,N_5189,N_3230);
xnor U8994 (N_8994,N_5259,N_5352);
or U8995 (N_8995,N_3480,N_5045);
nand U8996 (N_8996,N_5553,N_3345);
xor U8997 (N_8997,N_5077,N_5297);
or U8998 (N_8998,N_4301,N_5575);
nand U8999 (N_8999,N_5703,N_4343);
xor U9000 (N_9000,N_8404,N_7604);
nor U9001 (N_9001,N_6479,N_8273);
nor U9002 (N_9002,N_6346,N_8070);
nand U9003 (N_9003,N_7296,N_7939);
and U9004 (N_9004,N_7233,N_6339);
nor U9005 (N_9005,N_6644,N_6157);
or U9006 (N_9006,N_7986,N_7255);
or U9007 (N_9007,N_8945,N_8221);
and U9008 (N_9008,N_8819,N_8251);
or U9009 (N_9009,N_8242,N_8573);
nand U9010 (N_9010,N_8049,N_7334);
nor U9011 (N_9011,N_8328,N_6068);
xnor U9012 (N_9012,N_8399,N_7404);
and U9013 (N_9013,N_8772,N_6536);
nand U9014 (N_9014,N_7128,N_6015);
or U9015 (N_9015,N_6800,N_6091);
xor U9016 (N_9016,N_6863,N_6960);
nand U9017 (N_9017,N_6482,N_8548);
nor U9018 (N_9018,N_7639,N_8947);
nor U9019 (N_9019,N_6746,N_7187);
and U9020 (N_9020,N_8226,N_6999);
nor U9021 (N_9021,N_8732,N_7111);
and U9022 (N_9022,N_8874,N_6174);
xnor U9023 (N_9023,N_6309,N_8456);
xor U9024 (N_9024,N_8164,N_8295);
and U9025 (N_9025,N_7586,N_8030);
xnor U9026 (N_9026,N_6169,N_8855);
nor U9027 (N_9027,N_6350,N_8987);
or U9028 (N_9028,N_8312,N_7227);
nand U9029 (N_9029,N_8733,N_8095);
or U9030 (N_9030,N_8810,N_8009);
and U9031 (N_9031,N_8782,N_8002);
and U9032 (N_9032,N_6119,N_6601);
nand U9033 (N_9033,N_8254,N_7705);
nand U9034 (N_9034,N_7763,N_7168);
nand U9035 (N_9035,N_7571,N_7777);
nor U9036 (N_9036,N_8234,N_7938);
xor U9037 (N_9037,N_7865,N_7841);
or U9038 (N_9038,N_7288,N_7589);
nor U9039 (N_9039,N_6907,N_8672);
nor U9040 (N_9040,N_7207,N_8439);
nand U9041 (N_9041,N_6217,N_6668);
and U9042 (N_9042,N_6685,N_7023);
nor U9043 (N_9043,N_8657,N_7019);
or U9044 (N_9044,N_6300,N_8908);
nand U9045 (N_9045,N_6875,N_8899);
and U9046 (N_9046,N_6188,N_6964);
nand U9047 (N_9047,N_8122,N_8952);
xnor U9048 (N_9048,N_6653,N_8449);
xor U9049 (N_9049,N_6593,N_7521);
nand U9050 (N_9050,N_8724,N_6039);
nand U9051 (N_9051,N_7430,N_8541);
nand U9052 (N_9052,N_8005,N_8969);
xor U9053 (N_9053,N_6920,N_6265);
and U9054 (N_9054,N_7158,N_8338);
xor U9055 (N_9055,N_8118,N_7453);
or U9056 (N_9056,N_7951,N_8648);
or U9057 (N_9057,N_8434,N_6703);
and U9058 (N_9058,N_8068,N_8508);
and U9059 (N_9059,N_7578,N_7486);
or U9060 (N_9060,N_6697,N_8039);
nand U9061 (N_9061,N_8063,N_7648);
or U9062 (N_9062,N_7313,N_7029);
or U9063 (N_9063,N_8116,N_6180);
or U9064 (N_9064,N_7390,N_8527);
and U9065 (N_9065,N_7354,N_6911);
xnor U9066 (N_9066,N_7797,N_6430);
or U9067 (N_9067,N_7742,N_8773);
xor U9068 (N_9068,N_8781,N_8814);
nand U9069 (N_9069,N_6465,N_8942);
nand U9070 (N_9070,N_6834,N_8822);
xor U9071 (N_9071,N_7940,N_8110);
or U9072 (N_9072,N_6233,N_6542);
or U9073 (N_9073,N_8055,N_8883);
xnor U9074 (N_9074,N_6208,N_7009);
nand U9075 (N_9075,N_8484,N_6320);
nor U9076 (N_9076,N_6880,N_8085);
nand U9077 (N_9077,N_7934,N_7899);
or U9078 (N_9078,N_8971,N_6006);
and U9079 (N_9079,N_8139,N_8452);
and U9080 (N_9080,N_6105,N_6821);
or U9081 (N_9081,N_7320,N_7552);
or U9082 (N_9082,N_8424,N_8165);
nor U9083 (N_9083,N_7381,N_7593);
xnor U9084 (N_9084,N_8124,N_7646);
nor U9085 (N_9085,N_7045,N_7993);
or U9086 (N_9086,N_8436,N_7956);
and U9087 (N_9087,N_7916,N_8728);
or U9088 (N_9088,N_8785,N_8142);
or U9089 (N_9089,N_6059,N_6973);
nand U9090 (N_9090,N_8516,N_7941);
nor U9091 (N_9091,N_6066,N_6807);
nor U9092 (N_9092,N_8799,N_7670);
nor U9093 (N_9093,N_6134,N_8796);
and U9094 (N_9094,N_6355,N_6935);
and U9095 (N_9095,N_7640,N_8683);
nor U9096 (N_9096,N_7832,N_6824);
nor U9097 (N_9097,N_8358,N_8053);
or U9098 (N_9098,N_6885,N_7846);
nand U9099 (N_9099,N_6152,N_6822);
nor U9100 (N_9100,N_7905,N_7694);
or U9101 (N_9101,N_8830,N_7307);
xor U9102 (N_9102,N_8745,N_8504);
xor U9103 (N_9103,N_6285,N_8249);
or U9104 (N_9104,N_6596,N_8492);
or U9105 (N_9105,N_6184,N_7112);
nand U9106 (N_9106,N_7582,N_8612);
nor U9107 (N_9107,N_6253,N_8602);
xor U9108 (N_9108,N_7962,N_7321);
and U9109 (N_9109,N_8730,N_8911);
nor U9110 (N_9110,N_6416,N_8138);
nor U9111 (N_9111,N_8914,N_7871);
nor U9112 (N_9112,N_7231,N_8718);
xor U9113 (N_9113,N_8200,N_6996);
and U9114 (N_9114,N_8537,N_6149);
nand U9115 (N_9115,N_7125,N_6695);
xor U9116 (N_9116,N_6649,N_8647);
or U9117 (N_9117,N_6966,N_6295);
nor U9118 (N_9118,N_7740,N_6839);
nand U9119 (N_9119,N_8109,N_7926);
nand U9120 (N_9120,N_7588,N_7149);
and U9121 (N_9121,N_6938,N_8598);
nand U9122 (N_9122,N_6929,N_8052);
nand U9123 (N_9123,N_6014,N_6587);
nor U9124 (N_9124,N_8214,N_7503);
nand U9125 (N_9125,N_7650,N_7276);
nand U9126 (N_9126,N_6675,N_8089);
nor U9127 (N_9127,N_8862,N_6474);
xnor U9128 (N_9128,N_8276,N_8539);
or U9129 (N_9129,N_7386,N_8061);
or U9130 (N_9130,N_7081,N_6787);
or U9131 (N_9131,N_8681,N_6267);
nand U9132 (N_9132,N_8203,N_6958);
and U9133 (N_9133,N_8531,N_6426);
nand U9134 (N_9134,N_8778,N_6510);
and U9135 (N_9135,N_8075,N_8738);
and U9136 (N_9136,N_6343,N_7726);
nand U9137 (N_9137,N_7937,N_7765);
and U9138 (N_9138,N_8490,N_7062);
and U9139 (N_9139,N_6835,N_8210);
nor U9140 (N_9140,N_8524,N_7744);
and U9141 (N_9141,N_6572,N_7882);
and U9142 (N_9142,N_8169,N_6828);
xnor U9143 (N_9143,N_7867,N_8088);
or U9144 (N_9144,N_8589,N_8984);
nand U9145 (N_9145,N_8275,N_6256);
nor U9146 (N_9146,N_6759,N_7382);
and U9147 (N_9147,N_7718,N_8586);
and U9148 (N_9148,N_6901,N_7278);
nand U9149 (N_9149,N_7075,N_7105);
xnor U9150 (N_9150,N_6219,N_8595);
nand U9151 (N_9151,N_8507,N_7135);
nand U9152 (N_9152,N_8727,N_6705);
and U9153 (N_9153,N_6995,N_6225);
xnor U9154 (N_9154,N_7802,N_8430);
xnor U9155 (N_9155,N_7116,N_8550);
nand U9156 (N_9156,N_7847,N_6809);
or U9157 (N_9157,N_6077,N_6774);
nor U9158 (N_9158,N_7557,N_6769);
or U9159 (N_9159,N_8482,N_7725);
and U9160 (N_9160,N_6124,N_7051);
nor U9161 (N_9161,N_8438,N_8800);
nor U9162 (N_9162,N_8829,N_7374);
nor U9163 (N_9163,N_6406,N_6113);
and U9164 (N_9164,N_7040,N_6242);
nand U9165 (N_9165,N_6762,N_8175);
nor U9166 (N_9166,N_8685,N_6206);
or U9167 (N_9167,N_8188,N_6330);
and U9168 (N_9168,N_6715,N_7532);
xnor U9169 (N_9169,N_6467,N_7770);
nand U9170 (N_9170,N_7618,N_7540);
and U9171 (N_9171,N_8371,N_6965);
nor U9172 (N_9172,N_6001,N_8288);
nand U9173 (N_9173,N_7595,N_6879);
xnor U9174 (N_9174,N_7409,N_8036);
nand U9175 (N_9175,N_6148,N_6379);
and U9176 (N_9176,N_6031,N_6801);
nand U9177 (N_9177,N_8437,N_7336);
nand U9178 (N_9178,N_7814,N_7329);
or U9179 (N_9179,N_7999,N_6399);
xnor U9180 (N_9180,N_6045,N_6090);
and U9181 (N_9181,N_6266,N_7195);
xnor U9182 (N_9182,N_6236,N_6518);
and U9183 (N_9183,N_7903,N_7561);
nor U9184 (N_9184,N_7414,N_7308);
nor U9185 (N_9185,N_8154,N_8902);
nand U9186 (N_9186,N_6282,N_7964);
nor U9187 (N_9187,N_7746,N_6244);
nor U9188 (N_9188,N_7331,N_7043);
xor U9189 (N_9189,N_6700,N_7053);
nand U9190 (N_9190,N_7335,N_6509);
or U9191 (N_9191,N_6475,N_6020);
xnor U9192 (N_9192,N_7886,N_6251);
or U9193 (N_9193,N_7722,N_7470);
nand U9194 (N_9194,N_8852,N_7448);
or U9195 (N_9195,N_6261,N_6983);
nand U9196 (N_9196,N_6000,N_6449);
xor U9197 (N_9197,N_7574,N_8283);
or U9198 (N_9198,N_8755,N_8160);
nor U9199 (N_9199,N_7804,N_8267);
nor U9200 (N_9200,N_8513,N_7200);
and U9201 (N_9201,N_8082,N_6670);
and U9202 (N_9202,N_6733,N_8040);
and U9203 (N_9203,N_8306,N_6490);
nand U9204 (N_9204,N_8567,N_7018);
nor U9205 (N_9205,N_6210,N_8795);
nand U9206 (N_9206,N_7709,N_7151);
nand U9207 (N_9207,N_8624,N_6761);
nor U9208 (N_9208,N_6163,N_7041);
and U9209 (N_9209,N_8367,N_8467);
and U9210 (N_9210,N_8496,N_8059);
or U9211 (N_9211,N_7380,N_8475);
nand U9212 (N_9212,N_7910,N_7468);
xor U9213 (N_9213,N_6606,N_6940);
xor U9214 (N_9214,N_6257,N_6137);
or U9215 (N_9215,N_7267,N_7417);
nand U9216 (N_9216,N_8307,N_8754);
and U9217 (N_9217,N_6304,N_6293);
and U9218 (N_9218,N_7475,N_6928);
nand U9219 (N_9219,N_7680,N_8473);
nor U9220 (N_9220,N_7800,N_8892);
xor U9221 (N_9221,N_6401,N_7606);
xnor U9222 (N_9222,N_6894,N_8543);
and U9223 (N_9223,N_7114,N_8305);
nand U9224 (N_9224,N_7295,N_7172);
xnor U9225 (N_9225,N_7418,N_7849);
xnor U9226 (N_9226,N_8391,N_6364);
nor U9227 (N_9227,N_6856,N_7576);
and U9228 (N_9228,N_7790,N_8356);
and U9229 (N_9229,N_8860,N_7512);
and U9230 (N_9230,N_6892,N_7454);
nor U9231 (N_9231,N_8790,N_7368);
xnor U9232 (N_9232,N_7101,N_6888);
nand U9233 (N_9233,N_6029,N_8921);
and U9234 (N_9234,N_8000,N_7178);
nor U9235 (N_9235,N_6096,N_6146);
xor U9236 (N_9236,N_7658,N_8406);
and U9237 (N_9237,N_6042,N_7750);
xnor U9238 (N_9238,N_7667,N_8279);
or U9239 (N_9239,N_7154,N_7176);
and U9240 (N_9240,N_6511,N_7353);
nor U9241 (N_9241,N_7108,N_6906);
nand U9242 (N_9242,N_6579,N_6598);
nor U9243 (N_9243,N_7069,N_6602);
or U9244 (N_9244,N_8282,N_6594);
nand U9245 (N_9245,N_6589,N_6792);
nand U9246 (N_9246,N_6874,N_8613);
or U9247 (N_9247,N_6352,N_8823);
xor U9248 (N_9248,N_8857,N_6607);
nand U9249 (N_9249,N_8925,N_8615);
nand U9250 (N_9250,N_8466,N_8831);
nor U9251 (N_9251,N_8280,N_6757);
nand U9252 (N_9252,N_6680,N_6126);
nor U9253 (N_9253,N_6513,N_6179);
nand U9254 (N_9254,N_8007,N_7877);
nand U9255 (N_9255,N_7492,N_8509);
or U9256 (N_9256,N_7031,N_8532);
nand U9257 (N_9257,N_8032,N_8461);
and U9258 (N_9258,N_8669,N_7421);
xnor U9259 (N_9259,N_8020,N_8815);
and U9260 (N_9260,N_6424,N_6993);
and U9261 (N_9261,N_7309,N_6333);
nor U9262 (N_9262,N_7921,N_8723);
and U9263 (N_9263,N_8670,N_7537);
nor U9264 (N_9264,N_8783,N_8652);
nor U9265 (N_9265,N_6610,N_8735);
xnor U9266 (N_9266,N_7021,N_8576);
nor U9267 (N_9267,N_6915,N_6443);
xnor U9268 (N_9268,N_6711,N_7326);
xor U9269 (N_9269,N_6563,N_8364);
xor U9270 (N_9270,N_8211,N_7579);
or U9271 (N_9271,N_8596,N_7690);
or U9272 (N_9272,N_7079,N_6141);
and U9273 (N_9273,N_7126,N_6478);
nand U9274 (N_9274,N_6538,N_6004);
and U9275 (N_9275,N_7050,N_8592);
and U9276 (N_9276,N_8471,N_8818);
xor U9277 (N_9277,N_6299,N_7767);
nand U9278 (N_9278,N_7619,N_7609);
or U9279 (N_9279,N_8177,N_7923);
nand U9280 (N_9280,N_7346,N_7303);
nor U9281 (N_9281,N_7237,N_6094);
or U9282 (N_9282,N_7403,N_7592);
or U9283 (N_9283,N_8972,N_8923);
nor U9284 (N_9284,N_6561,N_6858);
or U9285 (N_9285,N_7985,N_6963);
xor U9286 (N_9286,N_6489,N_6464);
and U9287 (N_9287,N_7584,N_7524);
and U9288 (N_9288,N_6952,N_8445);
nor U9289 (N_9289,N_8885,N_8850);
nand U9290 (N_9290,N_6506,N_6065);
xor U9291 (N_9291,N_8431,N_8083);
nand U9292 (N_9292,N_6483,N_6850);
and U9293 (N_9293,N_8714,N_8149);
nor U9294 (N_9294,N_7212,N_8137);
and U9295 (N_9295,N_7929,N_7664);
and U9296 (N_9296,N_6463,N_8583);
nand U9297 (N_9297,N_6576,N_6493);
and U9298 (N_9298,N_7645,N_8111);
xor U9299 (N_9299,N_7808,N_6220);
and U9300 (N_9300,N_8924,N_8983);
xor U9301 (N_9301,N_6375,N_6165);
nor U9302 (N_9302,N_8352,N_8131);
and U9303 (N_9303,N_8120,N_8243);
and U9304 (N_9304,N_8198,N_8540);
nor U9305 (N_9305,N_8928,N_6345);
xnor U9306 (N_9306,N_6784,N_8300);
or U9307 (N_9307,N_7906,N_7543);
and U9308 (N_9308,N_8065,N_8938);
nor U9309 (N_9309,N_7093,N_7189);
and U9310 (N_9310,N_8476,N_7091);
xnor U9311 (N_9311,N_6072,N_8396);
and U9312 (N_9312,N_8272,N_8562);
or U9313 (N_9313,N_7751,N_8581);
and U9314 (N_9314,N_7196,N_8003);
xor U9315 (N_9315,N_6055,N_7925);
or U9316 (N_9316,N_8486,N_7387);
and U9317 (N_9317,N_6433,N_6704);
xor U9318 (N_9318,N_8631,N_6458);
nand U9319 (N_9319,N_6497,N_8479);
and U9320 (N_9320,N_8290,N_7431);
xnor U9321 (N_9321,N_6767,N_7193);
xnor U9322 (N_9322,N_8824,N_7446);
and U9323 (N_9323,N_8186,N_7282);
nor U9324 (N_9324,N_7973,N_8552);
xor U9325 (N_9325,N_8423,N_6073);
and U9326 (N_9326,N_7566,N_7104);
and U9327 (N_9327,N_6505,N_7612);
xnor U9328 (N_9328,N_8538,N_8895);
xnor U9329 (N_9329,N_6970,N_7698);
or U9330 (N_9330,N_7523,N_6196);
nor U9331 (N_9331,N_6953,N_8671);
nor U9332 (N_9332,N_6980,N_7241);
nor U9333 (N_9333,N_7902,N_8788);
nand U9334 (N_9334,N_6779,N_8878);
and U9335 (N_9335,N_8098,N_8004);
or U9336 (N_9336,N_6337,N_6175);
and U9337 (N_9337,N_7780,N_7162);
xor U9338 (N_9338,N_7057,N_8215);
or U9339 (N_9339,N_7788,N_6041);
nand U9340 (N_9340,N_6764,N_6583);
nand U9341 (N_9341,N_6117,N_8843);
nand U9342 (N_9342,N_7030,N_8890);
nor U9343 (N_9343,N_7337,N_7560);
nand U9344 (N_9344,N_8978,N_7654);
xor U9345 (N_9345,N_8974,N_6531);
nor U9346 (N_9346,N_7263,N_8907);
nand U9347 (N_9347,N_6447,N_6612);
and U9348 (N_9348,N_8792,N_6325);
nand U9349 (N_9349,N_8667,N_8327);
xnor U9350 (N_9350,N_8889,N_8879);
nand U9351 (N_9351,N_8835,N_8603);
or U9352 (N_9352,N_7302,N_6440);
and U9353 (N_9353,N_7248,N_6177);
nor U9354 (N_9354,N_7946,N_6310);
nand U9355 (N_9355,N_8045,N_6867);
xor U9356 (N_9356,N_8303,N_7798);
xor U9357 (N_9357,N_6092,N_8150);
nand U9358 (N_9358,N_6789,N_6326);
nor U9359 (N_9359,N_7657,N_6183);
nand U9360 (N_9360,N_7223,N_8027);
nor U9361 (N_9361,N_8599,N_7357);
and U9362 (N_9362,N_8378,N_6771);
or U9363 (N_9363,N_7054,N_8698);
xnor U9364 (N_9364,N_7813,N_6414);
xor U9365 (N_9365,N_6569,N_7887);
xor U9366 (N_9366,N_6636,N_8238);
nand U9367 (N_9367,N_7465,N_8780);
or U9368 (N_9368,N_8740,N_8465);
xor U9369 (N_9369,N_8315,N_7674);
nand U9370 (N_9370,N_7686,N_6254);
or U9371 (N_9371,N_6381,N_6327);
nand U9372 (N_9372,N_7013,N_7365);
nor U9373 (N_9373,N_7539,N_7131);
nor U9374 (N_9374,N_7478,N_6150);
nand U9375 (N_9375,N_7433,N_7710);
nand U9376 (N_9376,N_6128,N_7506);
nor U9377 (N_9377,N_8304,N_6147);
and U9378 (N_9378,N_6156,N_6144);
xnor U9379 (N_9379,N_8750,N_8563);
nor U9380 (N_9380,N_6584,N_6336);
xor U9381 (N_9381,N_6232,N_7637);
nor U9382 (N_9382,N_7016,N_6398);
and U9383 (N_9383,N_8347,N_7316);
or U9384 (N_9384,N_8751,N_8334);
nand U9385 (N_9385,N_6080,N_8610);
or U9386 (N_9386,N_6246,N_8235);
nand U9387 (N_9387,N_6713,N_6408);
nand U9388 (N_9388,N_6903,N_6603);
nand U9389 (N_9389,N_7174,N_7119);
nand U9390 (N_9390,N_6298,N_6671);
nor U9391 (N_9391,N_6294,N_6585);
xnor U9392 (N_9392,N_6878,N_6061);
nor U9393 (N_9393,N_6145,N_8162);
xor U9394 (N_9394,N_8067,N_7161);
or U9395 (N_9395,N_8134,N_6853);
nand U9396 (N_9396,N_8208,N_8369);
nand U9397 (N_9397,N_6022,N_6659);
nor U9398 (N_9398,N_6614,N_7089);
nor U9399 (N_9399,N_8337,N_7972);
and U9400 (N_9400,N_7583,N_7864);
nand U9401 (N_9401,N_8517,N_7229);
and U9402 (N_9402,N_8093,N_8884);
and U9403 (N_9403,N_7152,N_8661);
nor U9404 (N_9404,N_6548,N_6496);
and U9405 (N_9405,N_8656,N_8264);
xor U9406 (N_9406,N_8555,N_7875);
and U9407 (N_9407,N_7602,N_6898);
nand U9408 (N_9408,N_6830,N_7971);
nor U9409 (N_9409,N_7274,N_6303);
nand U9410 (N_9410,N_6205,N_8444);
and U9411 (N_9411,N_6485,N_6812);
xnor U9412 (N_9412,N_8939,N_8016);
nor U9413 (N_9413,N_7236,N_8114);
nor U9414 (N_9414,N_7142,N_6854);
or U9415 (N_9415,N_8521,N_6925);
and U9416 (N_9416,N_8271,N_8340);
xor U9417 (N_9417,N_7530,N_7830);
nor U9418 (N_9418,N_8183,N_8918);
or U9419 (N_9419,N_8140,N_7772);
nor U9420 (N_9420,N_7377,N_8643);
and U9421 (N_9421,N_6544,N_6630);
nand U9422 (N_9422,N_8559,N_6744);
xor U9423 (N_9423,N_7113,N_6372);
nor U9424 (N_9424,N_7860,N_8828);
and U9425 (N_9425,N_8566,N_6388);
and U9426 (N_9426,N_8277,N_6095);
and U9427 (N_9427,N_8336,N_7100);
nor U9428 (N_9428,N_8190,N_8887);
nor U9429 (N_9429,N_6871,N_7033);
or U9430 (N_9430,N_8632,N_6605);
nand U9431 (N_9431,N_8064,N_6480);
or U9432 (N_9432,N_7476,N_7333);
nand U9433 (N_9433,N_8588,N_6632);
or U9434 (N_9434,N_6241,N_8979);
nand U9435 (N_9435,N_8460,N_6287);
nand U9436 (N_9436,N_8074,N_6487);
xnor U9437 (N_9437,N_7577,N_8342);
or U9438 (N_9438,N_8167,N_6560);
nor U9439 (N_9439,N_8833,N_6328);
nor U9440 (N_9440,N_8247,N_6491);
nand U9441 (N_9441,N_7145,N_6305);
xor U9442 (N_9442,N_7678,N_8017);
xor U9443 (N_9443,N_7968,N_6338);
xor U9444 (N_9444,N_8867,N_7220);
and U9445 (N_9445,N_7035,N_7146);
nand U9446 (N_9446,N_6516,N_8076);
nand U9447 (N_9447,N_6747,N_7496);
nand U9448 (N_9448,N_7436,N_6026);
xnor U9449 (N_9449,N_8260,N_7010);
nor U9450 (N_9450,N_7753,N_7181);
nand U9451 (N_9451,N_6005,N_6526);
nor U9452 (N_9452,N_7070,N_7652);
or U9453 (N_9453,N_6722,N_6191);
or U9454 (N_9454,N_7547,N_8443);
nand U9455 (N_9455,N_6488,N_7489);
nand U9456 (N_9456,N_8665,N_8712);
nand U9457 (N_9457,N_7055,N_8410);
nand U9458 (N_9458,N_6377,N_8620);
and U9459 (N_9459,N_7842,N_6826);
nand U9460 (N_9460,N_7078,N_6389);
or U9461 (N_9461,N_6840,N_6450);
nand U9462 (N_9462,N_6990,N_7262);
xnor U9463 (N_9463,N_7514,N_8392);
nand U9464 (N_9464,N_7952,N_8663);
xor U9465 (N_9465,N_8310,N_7242);
and U9466 (N_9466,N_7815,N_7721);
and U9467 (N_9467,N_6620,N_7001);
nor U9468 (N_9468,N_6720,N_7816);
or U9469 (N_9469,N_7568,N_6131);
nor U9470 (N_9470,N_7201,N_7919);
nor U9471 (N_9471,N_7520,N_7538);
xor U9472 (N_9472,N_7559,N_6278);
nor U9473 (N_9473,N_8511,N_7504);
xnor U9474 (N_9474,N_8881,N_6886);
nor U9475 (N_9475,N_6286,N_7301);
nor U9476 (N_9476,N_8988,N_6959);
nor U9477 (N_9477,N_7736,N_6737);
or U9478 (N_9478,N_6638,N_8816);
and U9479 (N_9479,N_7005,N_6679);
nor U9480 (N_9480,N_8909,N_8742);
and U9481 (N_9481,N_7717,N_7617);
or U9482 (N_9482,N_7693,N_7655);
or U9483 (N_9483,N_7319,N_6248);
xnor U9484 (N_9484,N_7856,N_6941);
nand U9485 (N_9485,N_6986,N_6766);
and U9486 (N_9486,N_8308,N_8989);
xnor U9487 (N_9487,N_7920,N_7039);
xor U9488 (N_9488,N_6321,N_8489);
xor U9489 (N_9489,N_7794,N_6899);
and U9490 (N_9490,N_6547,N_6260);
nor U9491 (N_9491,N_7199,N_6089);
and U9492 (N_9492,N_7924,N_6831);
xor U9493 (N_9493,N_7297,N_8692);
or U9494 (N_9494,N_8927,N_7310);
or U9495 (N_9495,N_7825,N_7868);
xnor U9496 (N_9496,N_6155,N_7542);
and U9497 (N_9497,N_7124,N_7515);
and U9498 (N_9498,N_8397,N_7188);
xor U9499 (N_9499,N_7712,N_6643);
and U9500 (N_9500,N_7186,N_6949);
nand U9501 (N_9501,N_7180,N_6311);
and U9502 (N_9502,N_8353,N_7396);
nor U9503 (N_9503,N_8031,N_6931);
xnor U9504 (N_9504,N_8985,N_8682);
or U9505 (N_9505,N_8807,N_7271);
xnor U9506 (N_9506,N_6167,N_7415);
xor U9507 (N_9507,N_7215,N_6689);
nand U9508 (N_9508,N_6577,N_8932);
nand U9509 (N_9509,N_6776,N_8941);
or U9510 (N_9510,N_6914,N_6347);
or U9511 (N_9511,N_6817,N_7743);
xnor U9512 (N_9512,N_8078,N_6658);
nand U9513 (N_9513,N_8536,N_6773);
nand U9514 (N_9514,N_7771,N_7732);
nand U9515 (N_9515,N_6275,N_6778);
nor U9516 (N_9516,N_7836,N_8679);
nand U9517 (N_9517,N_6234,N_7981);
or U9518 (N_9518,N_8132,N_7420);
and U9519 (N_9519,N_7058,N_6405);
and U9520 (N_9520,N_6151,N_8230);
xnor U9521 (N_9521,N_8877,N_7960);
xor U9522 (N_9522,N_6500,N_7389);
or U9523 (N_9523,N_8905,N_7672);
xnor U9524 (N_9524,N_7094,N_7775);
nand U9525 (N_9525,N_8777,N_7385);
xor U9526 (N_9526,N_8993,N_6035);
nand U9527 (N_9527,N_8638,N_8207);
or U9528 (N_9528,N_8051,N_7615);
xnor U9529 (N_9529,N_7338,N_8706);
nand U9530 (N_9530,N_7824,N_7697);
nand U9531 (N_9531,N_6553,N_8798);
or U9532 (N_9532,N_8866,N_7622);
nor U9533 (N_9533,N_6452,N_6739);
xnor U9534 (N_9534,N_7474,N_7580);
nand U9535 (N_9535,N_8646,N_8287);
xnor U9536 (N_9536,N_7266,N_8417);
or U9537 (N_9537,N_7422,N_7363);
xor U9538 (N_9538,N_7644,N_8936);
or U9539 (N_9539,N_7912,N_8113);
xor U9540 (N_9540,N_7757,N_8704);
or U9541 (N_9541,N_8299,N_6228);
nand U9542 (N_9542,N_7117,N_8359);
nor U9543 (N_9543,N_7799,N_7160);
xor U9544 (N_9544,N_6471,N_7388);
xnor U9545 (N_9545,N_8227,N_8035);
nand U9546 (N_9546,N_8191,N_8854);
nor U9547 (N_9547,N_7769,N_6650);
nor U9548 (N_9548,N_8351,N_6361);
xnor U9549 (N_9549,N_7240,N_6866);
or U9550 (N_9550,N_7293,N_6604);
nor U9551 (N_9551,N_8864,N_7412);
xnor U9552 (N_9552,N_8660,N_8454);
and U9553 (N_9553,N_8687,N_7025);
nand U9554 (N_9554,N_7256,N_6557);
or U9555 (N_9555,N_8033,N_8689);
and U9556 (N_9556,N_7272,N_6955);
nand U9557 (N_9557,N_7961,N_7438);
or U9558 (N_9558,N_6988,N_7965);
xnor U9559 (N_9559,N_7760,N_7947);
xor U9560 (N_9560,N_7783,N_8954);
and U9561 (N_9561,N_7411,N_8321);
and U9562 (N_9562,N_8117,N_8494);
nand U9563 (N_9563,N_7234,N_6799);
or U9564 (N_9564,N_8153,N_8320);
nor U9565 (N_9565,N_6905,N_8827);
nand U9566 (N_9566,N_7083,N_8505);
nor U9567 (N_9567,N_8518,N_8529);
nand U9568 (N_9568,N_7853,N_8270);
or U9569 (N_9569,N_6631,N_7419);
or U9570 (N_9570,N_7118,N_7148);
or U9571 (N_9571,N_6111,N_7216);
nand U9572 (N_9572,N_6539,N_7834);
xor U9573 (N_9573,N_7391,N_6841);
xnor U9574 (N_9574,N_6642,N_7059);
nand U9575 (N_9575,N_8130,N_7198);
nor U9576 (N_9576,N_6460,N_6815);
nor U9577 (N_9577,N_8313,N_7205);
or U9578 (N_9578,N_7888,N_6218);
xor U9579 (N_9579,N_7507,N_6373);
xor U9580 (N_9580,N_7564,N_6729);
xor U9581 (N_9581,N_7121,N_7074);
or U9582 (N_9582,N_8825,N_6763);
nor U9583 (N_9583,N_8876,N_8256);
nor U9584 (N_9584,N_6833,N_6067);
xor U9585 (N_9585,N_7779,N_7575);
and U9586 (N_9586,N_6566,N_6382);
nand U9587 (N_9587,N_6384,N_6616);
or U9588 (N_9588,N_7003,N_6076);
and U9589 (N_9589,N_7287,N_8481);
or U9590 (N_9590,N_7076,N_8753);
nand U9591 (N_9591,N_6573,N_8970);
nor U9592 (N_9592,N_6741,N_7298);
nand U9593 (N_9593,N_6340,N_8094);
and U9594 (N_9594,N_8694,N_6582);
nand U9595 (N_9595,N_8224,N_6088);
and U9596 (N_9596,N_6537,N_7635);
nand U9597 (N_9597,N_8642,N_6276);
or U9598 (N_9598,N_6502,N_6288);
nand U9599 (N_9599,N_6192,N_8253);
xor U9600 (N_9600,N_7456,N_6992);
and U9601 (N_9601,N_8549,N_7792);
or U9602 (N_9602,N_7008,N_7061);
xor U9603 (N_9603,N_8726,N_7232);
or U9604 (N_9604,N_7891,N_7373);
nor U9605 (N_9605,N_7581,N_6292);
and U9606 (N_9606,N_8699,N_6371);
or U9607 (N_9607,N_8209,N_6574);
nor U9608 (N_9608,N_6877,N_8805);
nor U9609 (N_9609,N_7976,N_7245);
and U9610 (N_9610,N_8419,N_8991);
nand U9611 (N_9611,N_8673,N_6810);
nand U9612 (N_9612,N_8178,N_8056);
xor U9613 (N_9613,N_7279,N_8963);
nor U9614 (N_9614,N_7687,N_6639);
nor U9615 (N_9615,N_8897,N_8844);
nor U9616 (N_9616,N_7330,N_7932);
and U9617 (N_9617,N_8943,N_6550);
nor U9618 (N_9618,N_8820,N_6565);
or U9619 (N_9619,N_8856,N_6492);
or U9620 (N_9620,N_7260,N_7970);
nor U9621 (N_9621,N_6429,N_7183);
xor U9622 (N_9622,N_8703,N_7787);
nand U9623 (N_9623,N_7845,N_8764);
nor U9624 (N_9624,N_8469,N_7410);
nand U9625 (N_9625,N_8144,N_6932);
nand U9626 (N_9626,N_7895,N_6770);
nor U9627 (N_9627,N_7681,N_7315);
or U9628 (N_9628,N_6062,N_7192);
xor U9629 (N_9629,N_7628,N_6392);
and U9630 (N_9630,N_7812,N_8355);
xnor U9631 (N_9631,N_6690,N_8361);
xnor U9632 (N_9632,N_7228,N_7805);
and U9633 (N_9633,N_6843,N_6608);
or U9634 (N_9634,N_7634,N_8668);
nor U9635 (N_9635,N_7861,N_6738);
nand U9636 (N_9636,N_6376,N_7706);
nor U9637 (N_9637,N_7509,N_6984);
nor U9638 (N_9638,N_8766,N_6423);
and U9639 (N_9639,N_8298,N_6805);
nor U9640 (N_9640,N_6417,N_6717);
or U9641 (N_9641,N_7884,N_6393);
nor U9642 (N_9642,N_6698,N_6472);
nor U9643 (N_9643,N_8433,N_8281);
and U9644 (N_9644,N_8557,N_7957);
or U9645 (N_9645,N_7731,N_7259);
nand U9646 (N_9646,N_6535,N_8330);
or U9647 (N_9647,N_6823,N_8803);
nand U9648 (N_9648,N_8578,N_7450);
and U9649 (N_9649,N_6551,N_8691);
xor U9650 (N_9650,N_6876,N_7169);
xor U9651 (N_9651,N_6135,N_7627);
nor U9652 (N_9652,N_7442,N_7343);
and U9653 (N_9653,N_7498,N_8092);
nand U9654 (N_9654,N_8977,N_7349);
xor U9655 (N_9655,N_7127,N_8213);
nand U9656 (N_9656,N_8530,N_6540);
nand U9657 (N_9657,N_8953,N_7892);
xor U9658 (N_9658,N_8245,N_7513);
or U9659 (N_9659,N_8804,N_7696);
nand U9660 (N_9660,N_8389,N_8870);
xor U9661 (N_9661,N_8769,N_7364);
and U9662 (N_9662,N_6057,N_7483);
and U9663 (N_9663,N_7708,N_7324);
xor U9664 (N_9664,N_6368,N_6190);
and U9665 (N_9665,N_7833,N_6613);
or U9666 (N_9666,N_7164,N_6317);
xnor U9667 (N_9667,N_7407,N_7129);
xor U9668 (N_9668,N_7633,N_6825);
xnor U9669 (N_9669,N_6954,N_7803);
xnor U9670 (N_9670,N_7729,N_8676);
nor U9671 (N_9671,N_8651,N_6193);
xnor U9672 (N_9672,N_7848,N_7028);
and U9673 (N_9673,N_8180,N_6229);
nor U9674 (N_9674,N_8405,N_8323);
or U9675 (N_9675,N_7268,N_7137);
nor U9676 (N_9676,N_8990,N_8655);
xnor U9677 (N_9677,N_6344,N_8107);
nor U9678 (N_9678,N_6178,N_8503);
or U9679 (N_9679,N_7764,N_6360);
nand U9680 (N_9680,N_6008,N_8457);
and U9681 (N_9681,N_7555,N_8108);
nand U9682 (N_9682,N_7567,N_8289);
and U9683 (N_9683,N_6978,N_8637);
or U9684 (N_9684,N_7429,N_6431);
and U9685 (N_9685,N_6806,N_7980);
nor U9686 (N_9686,N_7866,N_6665);
or U9687 (N_9687,N_7990,N_6442);
and U9688 (N_9688,N_6819,N_7345);
nor U9689 (N_9689,N_8400,N_7528);
nor U9690 (N_9690,N_8653,N_6312);
xnor U9691 (N_9691,N_7701,N_7323);
xnor U9692 (N_9692,N_8845,N_8863);
nor U9693 (N_9693,N_6921,N_8791);
and U9694 (N_9694,N_7194,N_6648);
and U9695 (N_9695,N_8961,N_7294);
and U9696 (N_9696,N_7713,N_7840);
nand U9697 (N_9697,N_8992,N_6221);
and U9698 (N_9698,N_6897,N_7098);
and U9699 (N_9699,N_6793,N_7210);
nor U9700 (N_9700,N_7894,N_7774);
nor U9701 (N_9701,N_6852,N_7434);
or U9702 (N_9702,N_7402,N_8919);
nand U9703 (N_9703,N_6263,N_7641);
or U9704 (N_9704,N_6227,N_6358);
xnor U9705 (N_9705,N_7165,N_7631);
nand U9706 (N_9706,N_7510,N_8028);
nor U9707 (N_9707,N_6494,N_7546);
nand U9708 (N_9708,N_8341,N_6071);
xnor U9709 (N_9709,N_6855,N_8789);
nor U9710 (N_9710,N_8440,N_8693);
nor U9711 (N_9711,N_7066,N_7109);
nand U9712 (N_9712,N_7747,N_8395);
nor U9713 (N_9713,N_7254,N_6455);
and U9714 (N_9714,N_8101,N_6979);
nor U9715 (N_9715,N_6176,N_8317);
xnor U9716 (N_9716,N_6297,N_7443);
and U9717 (N_9717,N_7469,N_7688);
xnor U9718 (N_9718,N_6619,N_8960);
nor U9719 (N_9719,N_8565,N_6435);
nor U9720 (N_9720,N_8244,N_8384);
nor U9721 (N_9721,N_6237,N_6290);
and U9722 (N_9722,N_6075,N_7273);
xor U9723 (N_9723,N_6944,N_6198);
or U9724 (N_9724,N_7289,N_7325);
or U9725 (N_9725,N_8628,N_8266);
xor U9726 (N_9726,N_6116,N_8090);
or U9727 (N_9727,N_7208,N_7873);
or U9728 (N_9728,N_8520,N_6633);
nor U9729 (N_9729,N_7044,N_7684);
nor U9730 (N_9730,N_8808,N_8797);
or U9731 (N_9731,N_8184,N_6058);
and U9732 (N_9732,N_6837,N_6924);
or U9733 (N_9733,N_7449,N_7632);
xor U9734 (N_9734,N_6827,N_6971);
nor U9735 (N_9735,N_8627,N_7277);
nor U9736 (N_9736,N_7064,N_8293);
and U9737 (N_9737,N_7077,N_6054);
and U9738 (N_9738,N_6081,N_8459);
nand U9739 (N_9739,N_8201,N_8836);
and U9740 (N_9740,N_8707,N_8898);
nand U9741 (N_9741,N_7917,N_8577);
nor U9742 (N_9742,N_6628,N_7497);
or U9743 (N_9743,N_7572,N_8634);
nand U9744 (N_9744,N_6813,N_8708);
nor U9745 (N_9745,N_8848,N_8394);
nand U9746 (N_9746,N_8502,N_6567);
and U9747 (N_9747,N_6786,N_7974);
or U9748 (N_9748,N_6820,N_6100);
nor U9749 (N_9749,N_6238,N_6661);
and U9750 (N_9750,N_7206,N_7682);
xor U9751 (N_9751,N_8420,N_6755);
nor U9752 (N_9752,N_8901,N_8366);
or U9753 (N_9753,N_7616,N_7505);
and U9754 (N_9754,N_7317,N_8463);
nand U9755 (N_9755,N_6597,N_6279);
xor U9756 (N_9756,N_8127,N_8956);
xnor U9757 (N_9757,N_6136,N_6568);
nor U9758 (N_9758,N_7351,N_6975);
nor U9759 (N_9759,N_7928,N_8741);
xor U9760 (N_9760,N_8121,N_7494);
and U9761 (N_9761,N_8084,N_8023);
and U9762 (N_9762,N_7702,N_7073);
or U9763 (N_9763,N_7874,N_6887);
xnor U9764 (N_9764,N_7328,N_6790);
and U9765 (N_9765,N_6701,N_8401);
nor U9766 (N_9766,N_8455,N_7857);
or U9767 (N_9767,N_6063,N_8760);
xnor U9768 (N_9768,N_8239,N_8594);
and U9769 (N_9769,N_7662,N_7369);
nand U9770 (N_9770,N_7544,N_8206);
xor U9771 (N_9771,N_7367,N_7809);
xnor U9772 (N_9772,N_8622,N_7484);
nand U9773 (N_9773,N_8858,N_8386);
xor U9774 (N_9774,N_7378,N_7099);
nand U9775 (N_9775,N_7379,N_6437);
nand U9776 (N_9776,N_8967,N_6037);
or U9777 (N_9777,N_6331,N_7909);
and U9778 (N_9778,N_7977,N_8675);
or U9779 (N_9779,N_8379,N_8222);
xor U9780 (N_9780,N_8192,N_7230);
and U9781 (N_9781,N_8172,N_6224);
or U9782 (N_9782,N_8677,N_6469);
nor U9783 (N_9783,N_6873,N_8115);
nor U9784 (N_9784,N_6348,N_8846);
and U9785 (N_9785,N_8348,N_7837);
nor U9786 (N_9786,N_7318,N_7948);
and U9787 (N_9787,N_6515,N_6552);
nand U9788 (N_9788,N_7585,N_8717);
or U9789 (N_9789,N_8995,N_8106);
and U9790 (N_9790,N_8837,N_8817);
nand U9791 (N_9791,N_8570,N_8709);
nor U9792 (N_9792,N_6441,N_7123);
nor U9793 (N_9793,N_7102,N_8126);
xor U9794 (N_9794,N_7413,N_6160);
xor U9795 (N_9795,N_6865,N_8297);
nor U9796 (N_9796,N_8073,N_7455);
xnor U9797 (N_9797,N_7140,N_6484);
xnor U9798 (N_9798,N_6599,N_6981);
xnor U9799 (N_9799,N_7994,N_7945);
nand U9800 (N_9800,N_7024,N_8077);
xnor U9801 (N_9801,N_8787,N_8640);
nor U9802 (N_9802,N_8146,N_8618);
and U9803 (N_9803,N_6087,N_6798);
and U9804 (N_9804,N_7653,N_8523);
nor U9805 (N_9805,N_7911,N_8813);
or U9806 (N_9806,N_8324,N_7487);
nor U9807 (N_9807,N_8758,N_6622);
nor U9808 (N_9808,N_6592,N_7608);
xnor U9809 (N_9809,N_6968,N_8333);
xor U9810 (N_9810,N_8841,N_6504);
xnor U9811 (N_9811,N_8498,N_8861);
nand U9812 (N_9812,N_7243,N_6765);
nor U9813 (N_9813,N_6942,N_7372);
or U9814 (N_9814,N_8335,N_6101);
and U9815 (N_9815,N_8161,N_8409);
nor U9816 (N_9816,N_7679,N_7988);
nand U9817 (N_9817,N_6258,N_6872);
and U9818 (N_9818,N_7471,N_6663);
nand U9819 (N_9819,N_6950,N_6315);
xor U9820 (N_9820,N_6772,N_8980);
nor U9821 (N_9821,N_6943,N_8951);
nand U9822 (N_9822,N_6913,N_7522);
nor U9823 (N_9823,N_6754,N_6272);
xor U9824 (N_9824,N_6752,N_6794);
nand U9825 (N_9825,N_8382,N_7768);
and U9826 (N_9826,N_6154,N_8286);
xor U9827 (N_9827,N_7225,N_7397);
or U9828 (N_9828,N_7870,N_7340);
or U9829 (N_9829,N_6127,N_8512);
and U9830 (N_9830,N_6166,N_6555);
or U9831 (N_9831,N_7536,N_7950);
and U9832 (N_9832,N_8584,N_7036);
and U9833 (N_9833,N_8179,N_7133);
and U9834 (N_9834,N_8166,N_6781);
or U9835 (N_9835,N_6994,N_6291);
and U9836 (N_9836,N_7156,N_8725);
nor U9837 (N_9837,N_7499,N_6882);
nand U9838 (N_9838,N_7405,N_6323);
xnor U9839 (N_9839,N_6571,N_7534);
nand U9840 (N_9840,N_7224,N_8684);
or U9841 (N_9841,N_7171,N_8339);
nor U9842 (N_9842,N_8946,N_6412);
and U9843 (N_9843,N_8331,N_6222);
or U9844 (N_9844,N_6432,N_6207);
and U9845 (N_9845,N_8920,N_6987);
xor U9846 (N_9846,N_7984,N_7011);
or U9847 (N_9847,N_6070,N_8765);
nor U9848 (N_9848,N_7292,N_8719);
nand U9849 (N_9849,N_8875,N_6669);
or U9850 (N_9850,N_6378,N_6621);
or U9851 (N_9851,N_6123,N_7656);
and U9852 (N_9852,N_7006,N_7838);
or U9853 (N_9853,N_7918,N_6473);
or U9854 (N_9854,N_7426,N_7776);
and U9855 (N_9855,N_6335,N_7529);
and U9856 (N_9856,N_8241,N_7822);
nand U9857 (N_9857,N_8233,N_7179);
or U9858 (N_9858,N_8533,N_7827);
nand U9859 (N_9859,N_6354,N_6098);
xor U9860 (N_9860,N_6033,N_8006);
nand U9861 (N_9861,N_6301,N_8976);
or U9862 (N_9862,N_6780,N_6532);
xnor U9863 (N_9863,N_6477,N_7675);
nand U9864 (N_9864,N_6420,N_8219);
nor U9865 (N_9865,N_8365,N_8014);
or U9866 (N_9866,N_6027,N_7545);
xor U9867 (N_9867,N_6724,N_8141);
nand U9868 (N_9868,N_8880,N_6499);
nand U9869 (N_9869,N_7533,N_8526);
xnor U9870 (N_9870,N_7752,N_8545);
nor U9871 (N_9871,N_8387,N_6060);
xnor U9872 (N_9872,N_8955,N_6677);
nand U9873 (N_9873,N_6939,N_8022);
or U9874 (N_9874,N_8701,N_6250);
and U9875 (N_9875,N_7823,N_7042);
nor U9876 (N_9876,N_6170,N_6341);
xnor U9877 (N_9877,N_6588,N_6674);
xnor U9878 (N_9878,N_8500,N_8157);
nand U9879 (N_9879,N_8403,N_8362);
xnor U9880 (N_9880,N_8659,N_7935);
xnor U9881 (N_9881,N_7563,N_8413);
and U9882 (N_9882,N_8412,N_6777);
nor U9883 (N_9883,N_8480,N_6947);
and U9884 (N_9884,N_7943,N_8900);
nand U9885 (N_9885,N_6546,N_6507);
nor U9886 (N_9886,N_7573,N_6446);
and U9887 (N_9887,N_7197,N_7348);
nand U9888 (N_9888,N_6749,N_6107);
xor U9889 (N_9889,N_6554,N_8318);
and U9890 (N_9890,N_7643,N_7789);
xnor U9891 (N_9891,N_6403,N_8350);
xnor U9892 (N_9892,N_6590,N_6140);
xnor U9893 (N_9893,N_8906,N_6991);
nor U9894 (N_9894,N_7778,N_6397);
nor U9895 (N_9895,N_6164,N_8737);
and U9896 (N_9896,N_6402,N_8933);
nor U9897 (N_9897,N_6693,N_7477);
or U9898 (N_9898,N_8407,N_6891);
and U9899 (N_9899,N_6896,N_8937);
nand U9900 (N_9900,N_6349,N_6367);
nand U9901 (N_9901,N_6656,N_6314);
or U9902 (N_9902,N_8301,N_7601);
nor U9903 (N_9903,N_7550,N_6726);
or U9904 (N_9904,N_7737,N_8636);
xnor U9905 (N_9905,N_7649,N_8958);
or U9906 (N_9906,N_6721,N_8393);
nand U9907 (N_9907,N_6019,N_8994);
and U9908 (N_9908,N_8291,N_7110);
or U9909 (N_9909,N_8722,N_7314);
nand U9910 (N_9910,N_8853,N_6427);
or U9911 (N_9911,N_8102,N_8756);
or U9912 (N_9912,N_7138,N_7896);
or U9913 (N_9913,N_6667,N_8194);
or U9914 (N_9914,N_7458,N_8931);
nor U9915 (N_9915,N_8284,N_8212);
nand U9916 (N_9916,N_7460,N_7614);
xor U9917 (N_9917,N_6086,N_7147);
nand U9918 (N_9918,N_7922,N_6889);
and U9919 (N_9919,N_7663,N_7034);
nand U9920 (N_9920,N_6919,N_8158);
xor U9921 (N_9921,N_8381,N_8182);
and U9922 (N_9922,N_7949,N_6936);
nor U9923 (N_9923,N_6010,N_6386);
and U9924 (N_9924,N_7668,N_6106);
nor U9925 (N_9925,N_6374,N_8081);
and U9926 (N_9926,N_7084,N_8811);
xnor U9927 (N_9927,N_8054,N_8499);
or U9928 (N_9928,N_6112,N_6069);
and U9929 (N_9929,N_7253,N_8470);
and U9930 (N_9930,N_8849,N_7275);
xnor U9931 (N_9931,N_8997,N_6387);
nor U9932 (N_9932,N_8585,N_8294);
or U9933 (N_9933,N_7375,N_6273);
nor U9934 (N_9934,N_6049,N_7281);
xnor U9935 (N_9935,N_8119,N_7209);
nor U9936 (N_9936,N_7955,N_7959);
and U9937 (N_9937,N_8982,N_6280);
nor U9938 (N_9938,N_8826,N_8973);
xnor U9939 (N_9939,N_8525,N_7095);
and U9940 (N_9940,N_7488,N_6791);
or U9941 (N_9941,N_7989,N_8202);
nand U9942 (N_9942,N_8913,N_6064);
or U9943 (N_9943,N_6428,N_6047);
and U9944 (N_9944,N_6760,N_8590);
nand U9945 (N_9945,N_8185,N_6209);
nor U9946 (N_9946,N_7068,N_8561);
nand U9947 (N_9947,N_7611,N_7511);
or U9948 (N_9948,N_8148,N_8037);
and U9949 (N_9949,N_6723,N_7355);
xnor U9950 (N_9950,N_7967,N_6409);
xor U9951 (N_9951,N_8432,N_8872);
nand U9952 (N_9952,N_8176,N_8926);
and U9953 (N_9953,N_6422,N_8123);
xor U9954 (N_9954,N_7482,N_8232);
or U9955 (N_9955,N_7370,N_8551);
nor U9956 (N_9956,N_7286,N_7020);
and U9957 (N_9957,N_7673,N_8446);
or U9958 (N_9958,N_8060,N_6640);
or U9959 (N_9959,N_7191,N_8163);
or U9960 (N_9960,N_8173,N_8569);
nand U9961 (N_9961,N_6732,N_8746);
or U9962 (N_9962,N_6951,N_6758);
nand U9963 (N_9963,N_8047,N_8891);
nor U9964 (N_9964,N_6052,N_6407);
xnor U9965 (N_9965,N_6586,N_8058);
or U9966 (N_9966,N_6534,N_8731);
xor U9967 (N_9967,N_8375,N_7872);
xnor U9968 (N_9968,N_6525,N_7327);
nor U9969 (N_9969,N_7360,N_7120);
and U9970 (N_9970,N_8959,N_8859);
xor U9971 (N_9971,N_8493,N_7090);
and U9972 (N_9972,N_8228,N_6933);
nand U9973 (N_9973,N_8601,N_7786);
and U9974 (N_9974,N_7807,N_6074);
and U9975 (N_9975,N_8842,N_8246);
nand U9976 (N_9976,N_6696,N_6082);
nor U9977 (N_9977,N_6818,N_6719);
xor U9978 (N_9978,N_8448,N_7596);
and U9979 (N_9979,N_7835,N_7167);
and U9980 (N_9980,N_7843,N_8802);
or U9981 (N_9981,N_8217,N_7184);
xnor U9982 (N_9982,N_7218,N_8147);
or U9983 (N_9983,N_7214,N_8840);
nand U9984 (N_9984,N_6862,N_6881);
nand U9985 (N_9985,N_7395,N_7562);
xor U9986 (N_9986,N_7213,N_6211);
nand U9987 (N_9987,N_7982,N_7502);
and U9988 (N_9988,N_8012,N_8453);
or U9989 (N_9989,N_6296,N_6390);
or U9990 (N_9990,N_7699,N_8666);
and U9991 (N_9991,N_8274,N_8026);
nor U9992 (N_9992,N_7432,N_7852);
or U9993 (N_9993,N_6120,N_6411);
xnor U9994 (N_9994,N_8729,N_6842);
and U9995 (N_9995,N_8248,N_8639);
and U9996 (N_9996,N_7508,N_7211);
xnor U9997 (N_9997,N_7927,N_6556);
nand U9998 (N_9998,N_6625,N_7285);
nor U9999 (N_9999,N_6421,N_8547);
and U10000 (N_10000,N_7844,N_6439);
nor U10001 (N_10001,N_7423,N_6890);
nor U10002 (N_10002,N_8650,N_7610);
xor U10003 (N_10003,N_8558,N_7383);
and U10004 (N_10004,N_6974,N_6844);
nand U10005 (N_10005,N_6247,N_8105);
or U10006 (N_10006,N_8057,N_8767);
xor U10007 (N_10007,N_8635,N_8574);
xnor U10008 (N_10008,N_8368,N_6934);
nand U10009 (N_10009,N_8411,N_7629);
and U10010 (N_10010,N_6676,N_7855);
and U10011 (N_10011,N_6153,N_6673);
xor U10012 (N_10012,N_6083,N_6797);
nand U10013 (N_10013,N_6731,N_8776);
nand U10014 (N_10014,N_8644,N_7600);
and U10015 (N_10015,N_8104,N_6097);
xnor U10016 (N_10016,N_8903,N_8296);
and U10017 (N_10017,N_6618,N_8623);
xnor U10018 (N_10018,N_7092,N_8664);
xnor U10019 (N_10019,N_7002,N_6391);
and U10020 (N_10020,N_7669,N_6215);
nor U10021 (N_10021,N_6775,N_6269);
nand U10022 (N_10022,N_6351,N_6796);
nand U10023 (N_10023,N_6032,N_7879);
xor U10024 (N_10024,N_7027,N_6591);
xor U10025 (N_10025,N_7264,N_6716);
nand U10026 (N_10026,N_8501,N_6486);
and U10027 (N_10027,N_8839,N_8948);
nor U10028 (N_10028,N_7913,N_6945);
nor U10029 (N_10029,N_6158,N_8616);
xor U10030 (N_10030,N_8302,N_8633);
nand U10031 (N_10031,N_8218,N_8688);
xor U10032 (N_10032,N_6527,N_7936);
or U10033 (N_10033,N_6654,N_7106);
xnor U10034 (N_10034,N_8779,N_7202);
or U10035 (N_10035,N_7526,N_6118);
and U10036 (N_10036,N_6040,N_7480);
or U10037 (N_10037,N_6028,N_8690);
or U10038 (N_10038,N_6634,N_7141);
nor U10039 (N_10039,N_8168,N_7306);
xor U10040 (N_10040,N_6342,N_8886);
nor U10041 (N_10041,N_7408,N_7659);
xor U10042 (N_10042,N_8125,N_6687);
nor U10043 (N_10043,N_8621,N_7347);
nor U10044 (N_10044,N_8962,N_6735);
nand U10045 (N_10045,N_7048,N_8882);
nor U10046 (N_10046,N_7143,N_8629);
and U10047 (N_10047,N_8152,N_7716);
and U10048 (N_10048,N_6200,N_8388);
or U10049 (N_10049,N_7569,N_7554);
or U10050 (N_10050,N_6143,N_6910);
nor U10051 (N_10051,N_6025,N_6559);
and U10052 (N_10052,N_7914,N_7890);
or U10053 (N_10053,N_8174,N_7130);
and U10054 (N_10054,N_8560,N_7666);
nand U10055 (N_10055,N_8380,N_7150);
nor U10056 (N_10056,N_7996,N_8422);
nand U10057 (N_10057,N_7551,N_7818);
nand U10058 (N_10058,N_8332,N_8237);
nor U10059 (N_10059,N_7185,N_8506);
nand U10060 (N_10060,N_7107,N_7361);
xor U10061 (N_10061,N_6672,N_8447);
nand U10062 (N_10062,N_7052,N_8292);
xor U10063 (N_10063,N_8752,N_8832);
and U10064 (N_10064,N_7088,N_6804);
or U10065 (N_10065,N_6750,N_8794);
nand U10066 (N_10066,N_7441,N_8252);
xor U10067 (N_10067,N_8564,N_6734);
and U10068 (N_10068,N_6926,N_6223);
xor U10069 (N_10069,N_7762,N_8259);
nor U10070 (N_10070,N_6139,N_7014);
nand U10071 (N_10071,N_6365,N_6404);
nor U10072 (N_10072,N_7122,N_7817);
or U10073 (N_10073,N_6307,N_6845);
or U10074 (N_10074,N_6909,N_6453);
xor U10075 (N_10075,N_8021,N_8888);
nor U10076 (N_10076,N_7017,N_7247);
nor U10077 (N_10077,N_7352,N_6313);
or U10078 (N_10078,N_7638,N_6629);
nand U10079 (N_10079,N_7071,N_6457);
nand U10080 (N_10080,N_6363,N_6937);
nor U10081 (N_10081,N_8087,N_6162);
or U10082 (N_10082,N_7425,N_7881);
or U10083 (N_10083,N_6255,N_6519);
nand U10084 (N_10084,N_6595,N_8774);
nor U10085 (N_10085,N_7392,N_8649);
nor U10086 (N_10086,N_7738,N_6289);
or U10087 (N_10087,N_6635,N_6016);
or U10088 (N_10088,N_8042,N_7525);
and U10089 (N_10089,N_8944,N_7784);
xor U10090 (N_10090,N_6121,N_6520);
xnor U10091 (N_10091,N_7715,N_7284);
nor U10092 (N_10092,N_7829,N_8697);
or U10093 (N_10093,N_7007,N_7975);
nor U10094 (N_10094,N_7516,N_8225);
nor U10095 (N_10095,N_7217,N_7683);
and U10096 (N_10096,N_8749,N_7692);
and U10097 (N_10097,N_6549,N_6002);
nor U10098 (N_10098,N_8223,N_7821);
nand U10099 (N_10099,N_8528,N_8763);
xnor U10100 (N_10100,N_7219,N_8069);
or U10101 (N_10101,N_8702,N_6243);
or U10102 (N_10102,N_6611,N_7791);
and U10103 (N_10103,N_8968,N_6130);
nor U10104 (N_10104,N_6785,N_6385);
or U10105 (N_10105,N_7037,N_8491);
nor U10106 (N_10106,N_7793,N_6922);
nand U10107 (N_10107,N_7876,N_7362);
or U10108 (N_10108,N_6495,N_6109);
xor U10109 (N_10109,N_8205,N_8893);
xor U10110 (N_10110,N_6847,N_7144);
nand U10111 (N_10111,N_6962,N_6306);
and U10112 (N_10112,N_6977,N_7859);
and U10113 (N_10113,N_6528,N_8099);
and U10114 (N_10114,N_8710,N_8775);
nor U10115 (N_10115,N_8736,N_8606);
xor U10116 (N_10116,N_8641,N_8451);
and U10117 (N_10117,N_6262,N_7987);
or U10118 (N_10118,N_8345,N_8159);
nand U10119 (N_10119,N_8171,N_6989);
nand U10120 (N_10120,N_7930,N_8519);
and U10121 (N_10121,N_7820,N_7739);
or U10122 (N_10122,N_8376,N_8869);
xnor U10123 (N_10123,N_7464,N_8495);
nor U10124 (N_10124,N_6864,N_7481);
nand U10125 (N_10125,N_6930,N_7398);
xnor U10126 (N_10126,N_6459,N_6860);
or U10127 (N_10127,N_6728,N_6541);
nor U10128 (N_10128,N_8268,N_8464);
nand U10129 (N_10129,N_7339,N_7851);
and U10130 (N_10130,N_6836,N_8739);
or U10131 (N_10131,N_6036,N_7134);
nand U10132 (N_10132,N_6110,N_6181);
or U10133 (N_10133,N_8609,N_7749);
or U10134 (N_10134,N_8263,N_6957);
xnor U10135 (N_10135,N_8043,N_6912);
nor U10136 (N_10136,N_7558,N_6617);
nor U10137 (N_10137,N_6099,N_7304);
xnor U10138 (N_10138,N_7745,N_6908);
nand U10139 (N_10139,N_7953,N_6003);
nand U10140 (N_10140,N_7136,N_8197);
and U10141 (N_10141,N_6104,N_8319);
nand U10142 (N_10142,N_7332,N_7163);
nand U10143 (N_10143,N_6946,N_7621);
xor U10144 (N_10144,N_7495,N_6159);
or U10145 (N_10145,N_7252,N_6578);
or U10146 (N_10146,N_6011,N_6383);
nor U10147 (N_10147,N_6084,N_8600);
nor U10148 (N_10148,N_6413,N_6829);
nand U10149 (N_10149,N_7399,N_6647);
nand U10150 (N_10150,N_6956,N_6664);
nand U10151 (N_10151,N_8580,N_7491);
and U10152 (N_10152,N_8743,N_7898);
and U10153 (N_10153,N_7356,N_6883);
or U10154 (N_10154,N_6740,N_7944);
or U10155 (N_10155,N_8674,N_7394);
and U10156 (N_10156,N_7300,N_7155);
or U10157 (N_10157,N_8838,N_8019);
nor U10158 (N_10158,N_6425,N_8812);
nor U10159 (N_10159,N_8917,N_7685);
nor U10160 (N_10160,N_8930,N_6575);
xor U10161 (N_10161,N_7261,N_8196);
nand U10162 (N_10162,N_6699,N_8572);
and U10163 (N_10163,N_6395,N_8442);
nand U10164 (N_10164,N_8258,N_7642);
nor U10165 (N_10165,N_6727,N_8257);
nor U10166 (N_10166,N_6462,N_7754);
nor U10167 (N_10167,N_7072,N_6756);
or U10168 (N_10168,N_8128,N_7933);
or U10169 (N_10169,N_8136,N_7773);
and U10170 (N_10170,N_8510,N_7623);
nand U10171 (N_10171,N_7097,N_6362);
nor U10172 (N_10172,N_7979,N_7598);
and U10173 (N_10173,N_8383,N_7756);
xnor U10174 (N_10174,N_8062,N_7153);
nor U10175 (N_10175,N_8143,N_7660);
xnor U10176 (N_10176,N_8091,N_6195);
nor U10177 (N_10177,N_6318,N_6017);
or U10178 (N_10178,N_6470,N_7344);
and U10179 (N_10179,N_7531,N_7591);
xnor U10180 (N_10180,N_8398,N_8678);
nor U10181 (N_10181,N_7819,N_8129);
or U10182 (N_10182,N_7203,N_7741);
nor U10183 (N_10183,N_7517,N_8311);
and U10184 (N_10184,N_7893,N_6712);
xor U10185 (N_10185,N_7026,N_7400);
nor U10186 (N_10186,N_6203,N_7613);
nor U10187 (N_10187,N_8957,N_8086);
nor U10188 (N_10188,N_7587,N_7258);
nor U10189 (N_10189,N_8662,N_8587);
or U10190 (N_10190,N_6419,N_8189);
and U10191 (N_10191,N_7553,N_6708);
or U10192 (N_10192,N_6694,N_6508);
or U10193 (N_10193,N_7445,N_8011);
nand U10194 (N_10194,N_7594,N_8255);
or U10195 (N_10195,N_7416,N_6562);
nor U10196 (N_10196,N_6861,N_7661);
nand U10197 (N_10197,N_7785,N_6893);
or U10198 (N_10198,N_8071,N_7358);
nor U10199 (N_10199,N_8231,N_7424);
and U10200 (N_10200,N_6216,N_7590);
or U10201 (N_10201,N_8611,N_8579);
nand U10202 (N_10202,N_7485,N_6369);
or U10203 (N_10203,N_7992,N_6846);
xor U10204 (N_10204,N_6615,N_6048);
nand U10205 (N_10205,N_6691,N_8614);
or U10206 (N_10206,N_6284,N_7556);
or U10207 (N_10207,N_8713,N_7795);
xor U10208 (N_10208,N_8801,N_6816);
or U10209 (N_10209,N_8771,N_7863);
xnor U10210 (N_10210,N_8605,N_8762);
nor U10211 (N_10211,N_8535,N_7730);
xnor U10212 (N_10212,N_8097,N_8044);
nand U10213 (N_10213,N_6895,N_8001);
and U10214 (N_10214,N_6021,N_7599);
nand U10215 (N_10215,N_6782,N_7463);
nand U10216 (N_10216,N_6768,N_8770);
nor U10217 (N_10217,N_6194,N_7651);
nand U10218 (N_10218,N_8145,N_6231);
xnor U10219 (N_10219,N_8544,N_8744);
nand U10220 (N_10220,N_7004,N_8155);
nand U10221 (N_10221,N_8066,N_7060);
nor U10222 (N_10222,N_7467,N_6214);
and U10223 (N_10223,N_7630,N_7406);
or U10224 (N_10224,N_7473,N_7322);
nor U10225 (N_10225,N_6115,N_7761);
xor U10226 (N_10226,N_8426,N_6239);
nand U10227 (N_10227,N_6415,N_7811);
xnor U10228 (N_10228,N_7493,N_7733);
nand U10229 (N_10229,N_8048,N_8133);
and U10230 (N_10230,N_8096,N_8285);
or U10231 (N_10231,N_6917,N_6396);
or U10232 (N_10232,N_6524,N_8322);
nor U10233 (N_10233,N_7139,N_8597);
or U10234 (N_10234,N_7435,N_6370);
nor U10235 (N_10235,N_8363,N_6030);
xnor U10236 (N_10236,N_7997,N_6523);
or U10237 (N_10237,N_8193,N_8170);
xnor U10238 (N_10238,N_8996,N_6138);
and U10239 (N_10239,N_8010,N_8416);
xor U10240 (N_10240,N_7067,N_7257);
and U10241 (N_10241,N_7714,N_6581);
and U10242 (N_10242,N_7607,N_6743);
and U10243 (N_10243,N_7440,N_8806);
and U10244 (N_10244,N_6624,N_6503);
nand U10245 (N_10245,N_7689,N_6832);
and U10246 (N_10246,N_6102,N_8269);
or U10247 (N_10247,N_8871,N_8575);
nand U10248 (N_10248,N_6481,N_6900);
and U10249 (N_10249,N_7182,N_6129);
and U10250 (N_10250,N_8038,N_6249);
and U10251 (N_10251,N_8934,N_6454);
and U10252 (N_10252,N_8236,N_6870);
nor U10253 (N_10253,N_8721,N_8626);
nor U10254 (N_10254,N_7087,N_8402);
or U10255 (N_10255,N_7269,N_8630);
nand U10256 (N_10256,N_7625,N_7204);
nand U10257 (N_10257,N_7490,N_7707);
nor U10258 (N_10258,N_8408,N_7056);
nand U10259 (N_10259,N_7359,N_6501);
or U10260 (N_10260,N_8716,N_6707);
nor U10261 (N_10261,N_6264,N_7978);
or U10262 (N_10262,N_7782,N_7570);
and U10263 (N_10263,N_7447,N_6512);
and U10264 (N_10264,N_6053,N_7728);
xor U10265 (N_10265,N_6356,N_6125);
and U10266 (N_10266,N_8553,N_6666);
nand U10267 (N_10267,N_6122,N_6982);
and U10268 (N_10268,N_6366,N_6627);
or U10269 (N_10269,N_8896,N_6808);
or U10270 (N_10270,N_6009,N_8216);
xor U10271 (N_10271,N_8975,N_6626);
nand U10272 (N_10272,N_6600,N_6093);
xnor U10273 (N_10273,N_7647,N_7393);
and U10274 (N_10274,N_6702,N_8904);
nor U10275 (N_10275,N_6142,N_8761);
or U10276 (N_10276,N_6660,N_8617);
nand U10277 (N_10277,N_6838,N_7235);
and U10278 (N_10278,N_8607,N_7519);
xnor U10279 (N_10279,N_6972,N_7597);
and U10280 (N_10280,N_7854,N_7096);
xor U10281 (N_10281,N_8024,N_6132);
or U10282 (N_10282,N_6182,N_8514);
nor U10283 (N_10283,N_7244,N_6357);
xnor U10284 (N_10284,N_7000,N_8472);
or U10285 (N_10285,N_8385,N_8013);
nand U10286 (N_10286,N_8658,N_7942);
xnor U10287 (N_10287,N_6332,N_6133);
or U10288 (N_10288,N_8326,N_7720);
nand U10289 (N_10289,N_7624,N_7724);
xor U10290 (N_10290,N_6230,N_7371);
or U10291 (N_10291,N_8112,N_7080);
or U10292 (N_10292,N_6359,N_6745);
or U10293 (N_10293,N_8343,N_8204);
or U10294 (N_10294,N_6410,N_7366);
xnor U10295 (N_10295,N_8314,N_8793);
or U10296 (N_10296,N_8229,N_8240);
and U10297 (N_10297,N_7472,N_8034);
or U10298 (N_10298,N_7897,N_7880);
nand U10299 (N_10299,N_7901,N_6783);
xor U10300 (N_10300,N_6609,N_6085);
nand U10301 (N_10301,N_7085,N_7265);
or U10302 (N_10302,N_8418,N_7889);
xor U10303 (N_10303,N_7222,N_6709);
and U10304 (N_10304,N_8711,N_6199);
nand U10305 (N_10305,N_7312,N_7527);
nand U10306 (N_10306,N_8964,N_8571);
or U10307 (N_10307,N_8497,N_7676);
nor U10308 (N_10308,N_8757,N_6187);
and U10309 (N_10309,N_8025,N_7270);
and U10310 (N_10310,N_8374,N_6302);
xor U10311 (N_10311,N_6013,N_7170);
and U10312 (N_10312,N_7915,N_8415);
nand U10313 (N_10313,N_7781,N_7565);
xnor U10314 (N_10314,N_7479,N_6204);
nand U10315 (N_10315,N_8390,N_8485);
xnor U10316 (N_10316,N_8344,N_8734);
and U10317 (N_10317,N_7869,N_6688);
nor U10318 (N_10318,N_8786,N_7457);
nand U10319 (N_10319,N_6171,N_7839);
or U10320 (N_10320,N_8018,N_7704);
or U10321 (N_10321,N_8784,N_6023);
or U10322 (N_10322,N_7401,N_6436);
nor U10323 (N_10323,N_6322,N_6213);
nand U10324 (N_10324,N_7291,N_8966);
and U10325 (N_10325,N_7626,N_7991);
xor U10326 (N_10326,N_7734,N_8261);
nor U10327 (N_10327,N_6461,N_6245);
nand U10328 (N_10328,N_8072,N_6018);
and U10329 (N_10329,N_7462,N_8425);
nor U10330 (N_10330,N_6655,N_6530);
and U10331 (N_10331,N_7452,N_8748);
nor U10332 (N_10332,N_6274,N_7015);
or U10333 (N_10333,N_7451,N_6859);
xnor U10334 (N_10334,N_6451,N_7350);
nand U10335 (N_10335,N_6646,N_8821);
and U10336 (N_10336,N_6570,N_6564);
nor U10337 (N_10337,N_7691,N_7046);
or U10338 (N_10338,N_6788,N_7758);
nor U10339 (N_10339,N_6212,N_8619);
or U10340 (N_10340,N_6078,N_8029);
nand U10341 (N_10341,N_8654,N_8487);
and U10342 (N_10342,N_6651,N_7883);
nand U10343 (N_10343,N_7723,N_6706);
xnor U10344 (N_10344,N_6730,N_7801);
nand U10345 (N_10345,N_6038,N_8357);
xor U10346 (N_10346,N_7115,N_8477);
or U10347 (N_10347,N_6849,N_8591);
nand U10348 (N_10348,N_8768,N_6498);
nor U10349 (N_10349,N_6438,N_6533);
and U10350 (N_10350,N_6108,N_7459);
nand U10351 (N_10351,N_6418,N_7900);
xor U10352 (N_10352,N_7998,N_6725);
xor U10353 (N_10353,N_7700,N_7063);
nand U10354 (N_10354,N_8329,N_8156);
xnor U10355 (N_10355,N_8940,N_7246);
and U10356 (N_10356,N_6904,N_6869);
and U10357 (N_10357,N_8715,N_8346);
nand U10358 (N_10358,N_6448,N_6923);
or U10359 (N_10359,N_7549,N_7755);
nand U10360 (N_10360,N_7427,N_7958);
nand U10361 (N_10361,N_7103,N_6916);
and U10362 (N_10362,N_6168,N_7966);
nor U10363 (N_10363,N_6814,N_7541);
nand U10364 (N_10364,N_7735,N_6802);
and U10365 (N_10365,N_6985,N_7850);
nand U10366 (N_10366,N_8912,N_6444);
nand U10367 (N_10367,N_7132,N_6380);
xnor U10368 (N_10368,N_8705,N_7086);
nor U10369 (N_10369,N_7636,N_7796);
nor U10370 (N_10370,N_7461,N_7239);
nor U10371 (N_10371,N_8429,N_7862);
or U10372 (N_10372,N_6517,N_6927);
nand U10373 (N_10373,N_6811,N_8474);
or U10374 (N_10374,N_6277,N_6051);
or U10375 (N_10375,N_6268,N_6545);
nand U10376 (N_10376,N_8103,N_6969);
nor U10377 (N_10377,N_6851,N_8910);
or U10378 (N_10378,N_8534,N_7695);
nor U10379 (N_10379,N_7766,N_6400);
nand U10380 (N_10380,N_7166,N_8354);
nor U10381 (N_10381,N_6173,N_7065);
and U10382 (N_10382,N_7603,N_8680);
and U10383 (N_10383,N_8582,N_8435);
or U10384 (N_10384,N_6514,N_7500);
nor U10385 (N_10385,N_6645,N_7466);
nor U10386 (N_10386,N_6466,N_8041);
or U10387 (N_10387,N_7175,N_7159);
nor U10388 (N_10388,N_7047,N_7826);
nor U10389 (N_10389,N_8151,N_6201);
nand U10390 (N_10390,N_7904,N_6652);
nand U10391 (N_10391,N_8441,N_6434);
nor U10392 (N_10392,N_6103,N_7828);
nand U10393 (N_10393,N_7250,N_8250);
nand U10394 (N_10394,N_7878,N_6902);
nand U10395 (N_10395,N_6114,N_8046);
and U10396 (N_10396,N_7885,N_8080);
or U10397 (N_10397,N_8593,N_6998);
and U10398 (N_10398,N_8050,N_7384);
nand U10399 (N_10399,N_7501,N_8916);
nand U10400 (N_10400,N_6884,N_6012);
or U10401 (N_10401,N_6948,N_6580);
xnor U10402 (N_10402,N_6681,N_6308);
and U10403 (N_10403,N_7810,N_8759);
or U10404 (N_10404,N_8195,N_6456);
nor U10405 (N_10405,N_8468,N_7444);
and U10406 (N_10406,N_6657,N_7858);
nor U10407 (N_10407,N_7038,N_7439);
and U10408 (N_10408,N_6710,N_8949);
xnor U10409 (N_10409,N_6334,N_8100);
or U10410 (N_10410,N_8556,N_8372);
and U10411 (N_10411,N_8414,N_8428);
xnor U10412 (N_10412,N_6637,N_8998);
or U10413 (N_10413,N_7931,N_7719);
nor U10414 (N_10414,N_8349,N_7831);
nor U10415 (N_10415,N_6050,N_8522);
nand U10416 (N_10416,N_6529,N_8488);
and U10417 (N_10417,N_6161,N_6662);
or U10418 (N_10418,N_8181,N_7157);
xor U10419 (N_10419,N_8868,N_8999);
nand U10420 (N_10420,N_6961,N_6044);
nand U10421 (N_10421,N_8421,N_6034);
xor U10422 (N_10422,N_6189,N_6918);
or U10423 (N_10423,N_7703,N_6748);
xor U10424 (N_10424,N_7173,N_6270);
nor U10425 (N_10425,N_7221,N_8608);
and U10426 (N_10426,N_6623,N_6684);
nand U10427 (N_10427,N_8747,N_7022);
nor U10428 (N_10428,N_7665,N_6714);
xor U10429 (N_10429,N_6240,N_7305);
nor U10430 (N_10430,N_6718,N_6468);
xor U10431 (N_10431,N_6641,N_8458);
and U10432 (N_10432,N_8981,N_7311);
xor U10433 (N_10433,N_7190,N_7341);
or U10434 (N_10434,N_8809,N_7995);
nand U10435 (N_10435,N_8686,N_6521);
xnor U10436 (N_10436,N_7290,N_8986);
nand U10437 (N_10437,N_8373,N_8625);
and U10438 (N_10438,N_8700,N_8262);
nor U10439 (N_10439,N_8546,N_8645);
nand U10440 (N_10440,N_6394,N_7620);
and U10441 (N_10441,N_8316,N_6329);
nor U10442 (N_10442,N_7428,N_6046);
nand U10443 (N_10443,N_8950,N_8873);
nor U10444 (N_10444,N_6056,N_7280);
and U10445 (N_10445,N_7548,N_8199);
nor U10446 (N_10446,N_7908,N_8265);
nand U10447 (N_10447,N_8360,N_6742);
or U10448 (N_10448,N_7376,N_6283);
nor U10449 (N_10449,N_8450,N_8865);
nor U10450 (N_10450,N_7082,N_7806);
or U10451 (N_10451,N_6235,N_7049);
and U10452 (N_10452,N_6185,N_6172);
xor U10453 (N_10453,N_6736,N_6271);
and U10454 (N_10454,N_6324,N_8079);
nand U10455 (N_10455,N_8462,N_8542);
nor U10456 (N_10456,N_6997,N_6319);
and U10457 (N_10457,N_6678,N_6558);
xnor U10458 (N_10458,N_7605,N_6686);
and U10459 (N_10459,N_8377,N_6316);
xor U10460 (N_10460,N_6197,N_7535);
or U10461 (N_10461,N_6682,N_7671);
nand U10462 (N_10462,N_6692,N_6079);
nor U10463 (N_10463,N_6683,N_7299);
nand U10464 (N_10464,N_8187,N_7963);
nand U10465 (N_10465,N_6751,N_7251);
and U10466 (N_10466,N_8015,N_8695);
or U10467 (N_10467,N_8915,N_7437);
or U10468 (N_10468,N_7342,N_6024);
nand U10469 (N_10469,N_6857,N_8309);
and U10470 (N_10470,N_8696,N_7012);
xnor U10471 (N_10471,N_6976,N_6252);
nand U10472 (N_10472,N_8427,N_6281);
or U10473 (N_10473,N_7759,N_8847);
or U10474 (N_10474,N_8834,N_8515);
nand U10475 (N_10475,N_7249,N_6803);
nand U10476 (N_10476,N_8554,N_7518);
xor U10477 (N_10477,N_7983,N_7283);
nand U10478 (N_10478,N_8135,N_8965);
nor U10479 (N_10479,N_7748,N_8568);
or U10480 (N_10480,N_8008,N_6967);
or U10481 (N_10481,N_6868,N_8478);
or U10482 (N_10482,N_6226,N_7032);
nand U10483 (N_10483,N_8604,N_7177);
nor U10484 (N_10484,N_8278,N_8370);
nand U10485 (N_10485,N_6848,N_6795);
or U10486 (N_10486,N_8325,N_8720);
and U10487 (N_10487,N_7677,N_7969);
nor U10488 (N_10488,N_6202,N_6543);
or U10489 (N_10489,N_8929,N_6259);
nor U10490 (N_10490,N_6522,N_8922);
xor U10491 (N_10491,N_7238,N_7711);
or U10492 (N_10492,N_6186,N_7727);
xnor U10493 (N_10493,N_7954,N_7907);
nor U10494 (N_10494,N_6043,N_6476);
xor U10495 (N_10495,N_6445,N_8483);
nor U10496 (N_10496,N_8935,N_8894);
nand U10497 (N_10497,N_6753,N_8220);
and U10498 (N_10498,N_6353,N_6007);
nor U10499 (N_10499,N_8851,N_7226);
nor U10500 (N_10500,N_7459,N_7461);
nor U10501 (N_10501,N_8674,N_8701);
or U10502 (N_10502,N_6970,N_7721);
and U10503 (N_10503,N_8900,N_8893);
xor U10504 (N_10504,N_8467,N_8761);
xnor U10505 (N_10505,N_8292,N_8209);
nand U10506 (N_10506,N_7437,N_8673);
and U10507 (N_10507,N_7620,N_7876);
and U10508 (N_10508,N_6762,N_7585);
nand U10509 (N_10509,N_7180,N_8804);
nor U10510 (N_10510,N_7755,N_7303);
xor U10511 (N_10511,N_8184,N_6186);
and U10512 (N_10512,N_6974,N_8360);
nand U10513 (N_10513,N_8775,N_8025);
nand U10514 (N_10514,N_8993,N_8847);
and U10515 (N_10515,N_7616,N_6536);
xnor U10516 (N_10516,N_6579,N_8302);
or U10517 (N_10517,N_7647,N_7165);
and U10518 (N_10518,N_7897,N_8261);
nand U10519 (N_10519,N_8109,N_8565);
nor U10520 (N_10520,N_7479,N_6791);
and U10521 (N_10521,N_7974,N_6339);
nor U10522 (N_10522,N_8686,N_6910);
nand U10523 (N_10523,N_7674,N_6361);
nor U10524 (N_10524,N_6361,N_8089);
nor U10525 (N_10525,N_8292,N_7960);
or U10526 (N_10526,N_7571,N_6320);
and U10527 (N_10527,N_6523,N_7604);
xnor U10528 (N_10528,N_7892,N_8059);
or U10529 (N_10529,N_7913,N_6430);
and U10530 (N_10530,N_6513,N_8464);
or U10531 (N_10531,N_8907,N_6604);
or U10532 (N_10532,N_8910,N_8961);
or U10533 (N_10533,N_6924,N_8205);
or U10534 (N_10534,N_8076,N_6850);
or U10535 (N_10535,N_7630,N_7787);
and U10536 (N_10536,N_8514,N_8461);
nand U10537 (N_10537,N_6902,N_8451);
nand U10538 (N_10538,N_6606,N_6056);
and U10539 (N_10539,N_6353,N_6086);
nor U10540 (N_10540,N_7508,N_7227);
nand U10541 (N_10541,N_8802,N_8697);
nand U10542 (N_10542,N_7732,N_8657);
and U10543 (N_10543,N_6436,N_6518);
and U10544 (N_10544,N_8974,N_6298);
and U10545 (N_10545,N_6621,N_8851);
nand U10546 (N_10546,N_8636,N_6160);
nor U10547 (N_10547,N_6617,N_6101);
xor U10548 (N_10548,N_8989,N_7893);
nand U10549 (N_10549,N_8073,N_8609);
and U10550 (N_10550,N_6785,N_7239);
nor U10551 (N_10551,N_6786,N_7105);
xor U10552 (N_10552,N_6639,N_7470);
and U10553 (N_10553,N_7182,N_6500);
and U10554 (N_10554,N_7187,N_7690);
or U10555 (N_10555,N_8915,N_7160);
nand U10556 (N_10556,N_8924,N_8722);
or U10557 (N_10557,N_8074,N_6884);
and U10558 (N_10558,N_8134,N_6698);
nand U10559 (N_10559,N_7273,N_7342);
nor U10560 (N_10560,N_7510,N_8004);
nand U10561 (N_10561,N_6397,N_8880);
nor U10562 (N_10562,N_8594,N_8495);
nor U10563 (N_10563,N_8208,N_8639);
xor U10564 (N_10564,N_8777,N_8494);
xnor U10565 (N_10565,N_8872,N_7599);
xnor U10566 (N_10566,N_8740,N_8242);
nand U10567 (N_10567,N_7439,N_8028);
nor U10568 (N_10568,N_8724,N_8502);
and U10569 (N_10569,N_7214,N_7390);
nand U10570 (N_10570,N_6711,N_6571);
xnor U10571 (N_10571,N_8746,N_6132);
nand U10572 (N_10572,N_7677,N_7560);
xor U10573 (N_10573,N_6943,N_7768);
or U10574 (N_10574,N_6303,N_7732);
and U10575 (N_10575,N_6540,N_6911);
and U10576 (N_10576,N_7731,N_8799);
nor U10577 (N_10577,N_7654,N_7605);
xor U10578 (N_10578,N_7011,N_7811);
nor U10579 (N_10579,N_7844,N_8504);
nor U10580 (N_10580,N_7674,N_6620);
nor U10581 (N_10581,N_6216,N_6799);
nor U10582 (N_10582,N_8949,N_7577);
or U10583 (N_10583,N_6744,N_8476);
or U10584 (N_10584,N_7211,N_8498);
nand U10585 (N_10585,N_6916,N_6730);
nor U10586 (N_10586,N_6239,N_7986);
xnor U10587 (N_10587,N_8839,N_6588);
nand U10588 (N_10588,N_7126,N_7258);
and U10589 (N_10589,N_8571,N_6573);
nand U10590 (N_10590,N_7709,N_6552);
nor U10591 (N_10591,N_7651,N_8919);
xnor U10592 (N_10592,N_6550,N_8638);
xor U10593 (N_10593,N_8131,N_6058);
and U10594 (N_10594,N_6064,N_6462);
nor U10595 (N_10595,N_6340,N_6387);
and U10596 (N_10596,N_6973,N_7989);
and U10597 (N_10597,N_6050,N_8260);
and U10598 (N_10598,N_6515,N_6811);
or U10599 (N_10599,N_6556,N_7891);
nor U10600 (N_10600,N_6072,N_8657);
or U10601 (N_10601,N_8001,N_6625);
nor U10602 (N_10602,N_6275,N_6796);
nand U10603 (N_10603,N_7128,N_7620);
xnor U10604 (N_10604,N_8790,N_6256);
or U10605 (N_10605,N_7020,N_8733);
and U10606 (N_10606,N_7849,N_8734);
or U10607 (N_10607,N_7486,N_6699);
xnor U10608 (N_10608,N_7207,N_8782);
nor U10609 (N_10609,N_8459,N_6601);
nand U10610 (N_10610,N_6783,N_7092);
nand U10611 (N_10611,N_8453,N_6033);
nor U10612 (N_10612,N_8818,N_8437);
xnor U10613 (N_10613,N_6542,N_7648);
or U10614 (N_10614,N_7547,N_7615);
xnor U10615 (N_10615,N_8351,N_8868);
and U10616 (N_10616,N_8207,N_6802);
nand U10617 (N_10617,N_6669,N_7437);
and U10618 (N_10618,N_7015,N_8826);
xnor U10619 (N_10619,N_7798,N_7915);
nor U10620 (N_10620,N_6327,N_8429);
nand U10621 (N_10621,N_8360,N_7978);
nand U10622 (N_10622,N_6079,N_7200);
or U10623 (N_10623,N_7748,N_8124);
and U10624 (N_10624,N_8523,N_6242);
xor U10625 (N_10625,N_6729,N_8292);
nand U10626 (N_10626,N_6610,N_6121);
and U10627 (N_10627,N_6149,N_6701);
xor U10628 (N_10628,N_7290,N_6237);
nand U10629 (N_10629,N_6245,N_6237);
xnor U10630 (N_10630,N_7049,N_7592);
xnor U10631 (N_10631,N_6333,N_7939);
xnor U10632 (N_10632,N_8381,N_8342);
xnor U10633 (N_10633,N_7325,N_6314);
xnor U10634 (N_10634,N_6709,N_6319);
nor U10635 (N_10635,N_8821,N_7380);
or U10636 (N_10636,N_6701,N_8443);
nor U10637 (N_10637,N_6566,N_8990);
and U10638 (N_10638,N_8231,N_8022);
nand U10639 (N_10639,N_7262,N_8256);
xnor U10640 (N_10640,N_7247,N_7089);
and U10641 (N_10641,N_8038,N_6606);
or U10642 (N_10642,N_8051,N_7218);
or U10643 (N_10643,N_7321,N_7181);
and U10644 (N_10644,N_7850,N_7371);
nor U10645 (N_10645,N_8706,N_8087);
nand U10646 (N_10646,N_6031,N_7481);
and U10647 (N_10647,N_7304,N_8307);
xnor U10648 (N_10648,N_7821,N_6823);
or U10649 (N_10649,N_8951,N_7293);
xnor U10650 (N_10650,N_7304,N_6747);
xnor U10651 (N_10651,N_8882,N_8747);
and U10652 (N_10652,N_8643,N_6312);
and U10653 (N_10653,N_8989,N_6880);
nand U10654 (N_10654,N_6352,N_6843);
or U10655 (N_10655,N_6917,N_7542);
xor U10656 (N_10656,N_8307,N_8523);
nand U10657 (N_10657,N_7452,N_6738);
and U10658 (N_10658,N_7317,N_8616);
or U10659 (N_10659,N_7377,N_7841);
nand U10660 (N_10660,N_7222,N_7735);
xnor U10661 (N_10661,N_8144,N_7465);
xor U10662 (N_10662,N_7717,N_8908);
xnor U10663 (N_10663,N_6822,N_6427);
and U10664 (N_10664,N_6610,N_7622);
nor U10665 (N_10665,N_6766,N_8463);
or U10666 (N_10666,N_8980,N_6494);
nand U10667 (N_10667,N_8202,N_6510);
nor U10668 (N_10668,N_6720,N_7095);
or U10669 (N_10669,N_6849,N_6587);
nand U10670 (N_10670,N_8050,N_7403);
or U10671 (N_10671,N_8547,N_7714);
and U10672 (N_10672,N_8728,N_7537);
xnor U10673 (N_10673,N_6790,N_8327);
xnor U10674 (N_10674,N_8256,N_7334);
nor U10675 (N_10675,N_6782,N_7812);
and U10676 (N_10676,N_6437,N_8385);
nor U10677 (N_10677,N_6105,N_6487);
or U10678 (N_10678,N_6005,N_8364);
xor U10679 (N_10679,N_8088,N_8696);
or U10680 (N_10680,N_7026,N_6813);
xor U10681 (N_10681,N_6776,N_8842);
or U10682 (N_10682,N_7624,N_6191);
or U10683 (N_10683,N_6798,N_7028);
nor U10684 (N_10684,N_6848,N_8794);
or U10685 (N_10685,N_8123,N_6106);
nand U10686 (N_10686,N_6423,N_6440);
nor U10687 (N_10687,N_7712,N_8758);
or U10688 (N_10688,N_7755,N_6301);
nand U10689 (N_10689,N_7412,N_6465);
and U10690 (N_10690,N_7629,N_8898);
and U10691 (N_10691,N_7220,N_6557);
and U10692 (N_10692,N_8047,N_8235);
nor U10693 (N_10693,N_8183,N_7116);
nand U10694 (N_10694,N_7307,N_6057);
and U10695 (N_10695,N_8979,N_6700);
or U10696 (N_10696,N_6300,N_7450);
or U10697 (N_10697,N_8127,N_8506);
nor U10698 (N_10698,N_6556,N_7714);
and U10699 (N_10699,N_7318,N_8430);
and U10700 (N_10700,N_7642,N_6034);
and U10701 (N_10701,N_7961,N_6938);
xnor U10702 (N_10702,N_8234,N_6700);
xor U10703 (N_10703,N_6183,N_8328);
or U10704 (N_10704,N_6848,N_6287);
xnor U10705 (N_10705,N_7011,N_8144);
xnor U10706 (N_10706,N_6252,N_8402);
or U10707 (N_10707,N_8584,N_7836);
and U10708 (N_10708,N_8269,N_6892);
or U10709 (N_10709,N_7570,N_6691);
nor U10710 (N_10710,N_6561,N_7779);
and U10711 (N_10711,N_6727,N_7042);
nor U10712 (N_10712,N_6569,N_6555);
nand U10713 (N_10713,N_8034,N_8899);
xor U10714 (N_10714,N_7098,N_8410);
nor U10715 (N_10715,N_8472,N_8441);
or U10716 (N_10716,N_6363,N_8580);
nand U10717 (N_10717,N_7348,N_7324);
xor U10718 (N_10718,N_6991,N_6496);
nor U10719 (N_10719,N_8369,N_7078);
or U10720 (N_10720,N_8199,N_8243);
or U10721 (N_10721,N_7042,N_8987);
and U10722 (N_10722,N_7855,N_6791);
or U10723 (N_10723,N_6489,N_6847);
nor U10724 (N_10724,N_6810,N_6923);
nor U10725 (N_10725,N_7691,N_8441);
nor U10726 (N_10726,N_6469,N_7677);
nand U10727 (N_10727,N_6118,N_8879);
nand U10728 (N_10728,N_7870,N_8677);
xnor U10729 (N_10729,N_8866,N_6538);
and U10730 (N_10730,N_7411,N_7347);
xnor U10731 (N_10731,N_6728,N_6842);
or U10732 (N_10732,N_6930,N_6527);
and U10733 (N_10733,N_6973,N_6278);
and U10734 (N_10734,N_6486,N_6290);
or U10735 (N_10735,N_7781,N_6779);
nor U10736 (N_10736,N_7345,N_8169);
nand U10737 (N_10737,N_8859,N_6965);
xor U10738 (N_10738,N_8875,N_7022);
nand U10739 (N_10739,N_6880,N_6769);
or U10740 (N_10740,N_6375,N_8563);
and U10741 (N_10741,N_7016,N_8882);
or U10742 (N_10742,N_7111,N_6036);
and U10743 (N_10743,N_8902,N_7938);
xor U10744 (N_10744,N_8356,N_8855);
nand U10745 (N_10745,N_7611,N_6942);
nand U10746 (N_10746,N_8836,N_8026);
xor U10747 (N_10747,N_6444,N_7341);
nand U10748 (N_10748,N_7098,N_6735);
or U10749 (N_10749,N_6099,N_8291);
or U10750 (N_10750,N_6199,N_8084);
nand U10751 (N_10751,N_8409,N_6071);
and U10752 (N_10752,N_8433,N_6180);
nand U10753 (N_10753,N_6578,N_7527);
xor U10754 (N_10754,N_6452,N_6703);
xnor U10755 (N_10755,N_6091,N_7543);
nand U10756 (N_10756,N_7785,N_6100);
and U10757 (N_10757,N_6613,N_6154);
nor U10758 (N_10758,N_6896,N_6980);
nand U10759 (N_10759,N_7069,N_6179);
nor U10760 (N_10760,N_6774,N_7957);
nand U10761 (N_10761,N_6091,N_8663);
nor U10762 (N_10762,N_7282,N_7662);
or U10763 (N_10763,N_8136,N_6337);
nor U10764 (N_10764,N_8995,N_8475);
nor U10765 (N_10765,N_7742,N_7133);
or U10766 (N_10766,N_7616,N_8618);
xor U10767 (N_10767,N_8490,N_7092);
and U10768 (N_10768,N_6756,N_6986);
nand U10769 (N_10769,N_7265,N_8349);
or U10770 (N_10770,N_6708,N_7241);
nand U10771 (N_10771,N_7671,N_6360);
nor U10772 (N_10772,N_6536,N_8793);
nor U10773 (N_10773,N_6693,N_8448);
xor U10774 (N_10774,N_7503,N_6356);
nand U10775 (N_10775,N_6138,N_8907);
or U10776 (N_10776,N_6599,N_7695);
nand U10777 (N_10777,N_8144,N_7733);
or U10778 (N_10778,N_8541,N_8335);
and U10779 (N_10779,N_7383,N_7023);
nor U10780 (N_10780,N_6940,N_7722);
or U10781 (N_10781,N_7956,N_6508);
nand U10782 (N_10782,N_8237,N_8704);
or U10783 (N_10783,N_8303,N_8410);
nor U10784 (N_10784,N_7302,N_6612);
nor U10785 (N_10785,N_8739,N_7306);
nand U10786 (N_10786,N_8978,N_7274);
xnor U10787 (N_10787,N_8715,N_6988);
nand U10788 (N_10788,N_7145,N_7311);
and U10789 (N_10789,N_6149,N_8577);
or U10790 (N_10790,N_6404,N_7496);
nor U10791 (N_10791,N_8486,N_8699);
or U10792 (N_10792,N_6172,N_7662);
and U10793 (N_10793,N_8712,N_8954);
and U10794 (N_10794,N_7129,N_7370);
or U10795 (N_10795,N_8963,N_8130);
nand U10796 (N_10796,N_6109,N_7194);
or U10797 (N_10797,N_7576,N_7150);
xnor U10798 (N_10798,N_6858,N_6323);
xnor U10799 (N_10799,N_8207,N_6129);
nand U10800 (N_10800,N_7875,N_7362);
xnor U10801 (N_10801,N_8025,N_8977);
nor U10802 (N_10802,N_6733,N_6312);
nor U10803 (N_10803,N_6106,N_8613);
nor U10804 (N_10804,N_8214,N_6664);
and U10805 (N_10805,N_6499,N_8015);
and U10806 (N_10806,N_8122,N_7032);
xor U10807 (N_10807,N_7152,N_8116);
xor U10808 (N_10808,N_6039,N_8603);
nand U10809 (N_10809,N_7618,N_8175);
xor U10810 (N_10810,N_6981,N_6540);
and U10811 (N_10811,N_8356,N_8214);
nand U10812 (N_10812,N_7736,N_7727);
nor U10813 (N_10813,N_6819,N_8413);
or U10814 (N_10814,N_8072,N_8567);
nand U10815 (N_10815,N_6219,N_6444);
and U10816 (N_10816,N_8757,N_8893);
nand U10817 (N_10817,N_7651,N_7565);
xnor U10818 (N_10818,N_8703,N_6687);
xnor U10819 (N_10819,N_6839,N_6277);
and U10820 (N_10820,N_7914,N_8050);
or U10821 (N_10821,N_6690,N_7070);
nand U10822 (N_10822,N_8154,N_6187);
nand U10823 (N_10823,N_6158,N_6795);
or U10824 (N_10824,N_7031,N_8257);
xnor U10825 (N_10825,N_6397,N_8463);
nor U10826 (N_10826,N_8509,N_7080);
nand U10827 (N_10827,N_6603,N_8066);
nor U10828 (N_10828,N_6871,N_6686);
xnor U10829 (N_10829,N_8914,N_6974);
nand U10830 (N_10830,N_8900,N_8929);
nor U10831 (N_10831,N_7421,N_6945);
and U10832 (N_10832,N_7142,N_8768);
or U10833 (N_10833,N_7061,N_8139);
or U10834 (N_10834,N_6123,N_8454);
nand U10835 (N_10835,N_8805,N_8756);
and U10836 (N_10836,N_7084,N_8500);
xnor U10837 (N_10837,N_6313,N_6267);
or U10838 (N_10838,N_8836,N_7518);
or U10839 (N_10839,N_7623,N_7988);
or U10840 (N_10840,N_8988,N_8090);
nand U10841 (N_10841,N_7332,N_7533);
nand U10842 (N_10842,N_6705,N_8026);
nor U10843 (N_10843,N_6530,N_7980);
or U10844 (N_10844,N_6068,N_7112);
nor U10845 (N_10845,N_8392,N_6499);
nor U10846 (N_10846,N_6680,N_7201);
and U10847 (N_10847,N_7189,N_6076);
xnor U10848 (N_10848,N_8754,N_7551);
xor U10849 (N_10849,N_8482,N_6818);
or U10850 (N_10850,N_8410,N_7750);
or U10851 (N_10851,N_8255,N_7451);
nand U10852 (N_10852,N_6767,N_8938);
nor U10853 (N_10853,N_8316,N_8272);
nor U10854 (N_10854,N_6483,N_7447);
or U10855 (N_10855,N_8150,N_6393);
nand U10856 (N_10856,N_8576,N_6785);
nor U10857 (N_10857,N_6396,N_8365);
xor U10858 (N_10858,N_8826,N_8575);
nor U10859 (N_10859,N_7538,N_7904);
xor U10860 (N_10860,N_6979,N_7147);
xor U10861 (N_10861,N_7951,N_7045);
nand U10862 (N_10862,N_8273,N_8640);
or U10863 (N_10863,N_6332,N_6511);
and U10864 (N_10864,N_8005,N_6712);
and U10865 (N_10865,N_6378,N_6401);
and U10866 (N_10866,N_8427,N_8336);
and U10867 (N_10867,N_7907,N_6260);
xor U10868 (N_10868,N_8975,N_8360);
and U10869 (N_10869,N_7773,N_7744);
and U10870 (N_10870,N_8752,N_8052);
nor U10871 (N_10871,N_7836,N_7710);
or U10872 (N_10872,N_6440,N_6752);
nor U10873 (N_10873,N_7345,N_6835);
or U10874 (N_10874,N_8396,N_7236);
nand U10875 (N_10875,N_6755,N_8363);
and U10876 (N_10876,N_6680,N_7640);
or U10877 (N_10877,N_7480,N_7752);
xor U10878 (N_10878,N_8207,N_6603);
or U10879 (N_10879,N_6864,N_6524);
nor U10880 (N_10880,N_7499,N_7619);
nor U10881 (N_10881,N_7639,N_6989);
nand U10882 (N_10882,N_8019,N_7340);
nand U10883 (N_10883,N_7800,N_8594);
or U10884 (N_10884,N_7151,N_6708);
nor U10885 (N_10885,N_7406,N_6953);
xor U10886 (N_10886,N_7468,N_7926);
xor U10887 (N_10887,N_7035,N_8449);
nand U10888 (N_10888,N_8735,N_7723);
nand U10889 (N_10889,N_7730,N_8217);
and U10890 (N_10890,N_7430,N_6590);
nor U10891 (N_10891,N_6953,N_6003);
and U10892 (N_10892,N_8818,N_6966);
nor U10893 (N_10893,N_8313,N_8868);
xor U10894 (N_10894,N_8034,N_7143);
or U10895 (N_10895,N_6545,N_7987);
or U10896 (N_10896,N_6908,N_8903);
or U10897 (N_10897,N_7991,N_6212);
or U10898 (N_10898,N_8271,N_6010);
nor U10899 (N_10899,N_7088,N_8706);
and U10900 (N_10900,N_8154,N_8965);
xnor U10901 (N_10901,N_6757,N_8643);
or U10902 (N_10902,N_6435,N_7748);
nand U10903 (N_10903,N_6574,N_6676);
nand U10904 (N_10904,N_7595,N_6372);
xnor U10905 (N_10905,N_7827,N_7614);
or U10906 (N_10906,N_7169,N_8355);
nand U10907 (N_10907,N_6580,N_6264);
and U10908 (N_10908,N_7712,N_7347);
and U10909 (N_10909,N_7681,N_8386);
xor U10910 (N_10910,N_6816,N_6046);
and U10911 (N_10911,N_8041,N_6139);
or U10912 (N_10912,N_8423,N_7460);
or U10913 (N_10913,N_8290,N_7308);
xnor U10914 (N_10914,N_7016,N_8583);
xor U10915 (N_10915,N_8695,N_8172);
xor U10916 (N_10916,N_6503,N_7099);
nand U10917 (N_10917,N_7129,N_6886);
xor U10918 (N_10918,N_6233,N_7429);
or U10919 (N_10919,N_6200,N_7179);
or U10920 (N_10920,N_8075,N_6636);
nand U10921 (N_10921,N_7913,N_6135);
and U10922 (N_10922,N_8055,N_6102);
nand U10923 (N_10923,N_7005,N_8895);
and U10924 (N_10924,N_8596,N_6916);
nand U10925 (N_10925,N_6918,N_7834);
xnor U10926 (N_10926,N_7642,N_6425);
and U10927 (N_10927,N_8748,N_8938);
xor U10928 (N_10928,N_8336,N_6170);
or U10929 (N_10929,N_8938,N_6115);
or U10930 (N_10930,N_6955,N_8521);
nor U10931 (N_10931,N_8468,N_6034);
and U10932 (N_10932,N_8402,N_6347);
or U10933 (N_10933,N_6602,N_6471);
or U10934 (N_10934,N_8239,N_6957);
and U10935 (N_10935,N_7955,N_8998);
nand U10936 (N_10936,N_8183,N_7452);
xor U10937 (N_10937,N_7410,N_6663);
xor U10938 (N_10938,N_7839,N_8111);
and U10939 (N_10939,N_8044,N_7979);
nand U10940 (N_10940,N_8015,N_8918);
nor U10941 (N_10941,N_8880,N_7989);
or U10942 (N_10942,N_8103,N_7669);
nor U10943 (N_10943,N_7692,N_8570);
and U10944 (N_10944,N_7250,N_7130);
or U10945 (N_10945,N_8741,N_8925);
nand U10946 (N_10946,N_6268,N_6200);
nand U10947 (N_10947,N_7456,N_6423);
xor U10948 (N_10948,N_8110,N_8824);
nand U10949 (N_10949,N_7919,N_8363);
and U10950 (N_10950,N_8641,N_7871);
and U10951 (N_10951,N_8988,N_8061);
xor U10952 (N_10952,N_8645,N_8475);
xnor U10953 (N_10953,N_7051,N_7888);
and U10954 (N_10954,N_6679,N_7710);
and U10955 (N_10955,N_6556,N_8595);
and U10956 (N_10956,N_8036,N_7912);
xor U10957 (N_10957,N_8979,N_6609);
nor U10958 (N_10958,N_6088,N_6095);
xor U10959 (N_10959,N_6859,N_8434);
or U10960 (N_10960,N_6070,N_8871);
nor U10961 (N_10961,N_8770,N_8094);
xnor U10962 (N_10962,N_7958,N_7660);
nand U10963 (N_10963,N_6128,N_8330);
and U10964 (N_10964,N_6279,N_7636);
and U10965 (N_10965,N_6820,N_8000);
and U10966 (N_10966,N_7097,N_6645);
nand U10967 (N_10967,N_7877,N_8140);
xor U10968 (N_10968,N_7157,N_7332);
or U10969 (N_10969,N_6538,N_7075);
nand U10970 (N_10970,N_8829,N_8969);
or U10971 (N_10971,N_7284,N_6801);
nor U10972 (N_10972,N_8326,N_8022);
nand U10973 (N_10973,N_6752,N_7585);
nor U10974 (N_10974,N_7699,N_7107);
xnor U10975 (N_10975,N_7197,N_7941);
and U10976 (N_10976,N_8896,N_6811);
nor U10977 (N_10977,N_8530,N_8710);
nand U10978 (N_10978,N_7277,N_7984);
or U10979 (N_10979,N_6541,N_8582);
or U10980 (N_10980,N_8606,N_8151);
nand U10981 (N_10981,N_6800,N_8013);
and U10982 (N_10982,N_7191,N_7197);
nand U10983 (N_10983,N_8088,N_8057);
xnor U10984 (N_10984,N_6261,N_6989);
xnor U10985 (N_10985,N_6790,N_7862);
nand U10986 (N_10986,N_6187,N_7271);
and U10987 (N_10987,N_7056,N_7905);
xnor U10988 (N_10988,N_8297,N_7308);
and U10989 (N_10989,N_8529,N_6934);
or U10990 (N_10990,N_7018,N_7625);
and U10991 (N_10991,N_6983,N_6247);
xor U10992 (N_10992,N_7243,N_7099);
nor U10993 (N_10993,N_6696,N_7254);
nor U10994 (N_10994,N_7366,N_6973);
and U10995 (N_10995,N_6167,N_7452);
nor U10996 (N_10996,N_7224,N_7273);
nor U10997 (N_10997,N_8777,N_8851);
or U10998 (N_10998,N_7455,N_7735);
nand U10999 (N_10999,N_8974,N_6052);
or U11000 (N_11000,N_7844,N_6452);
xor U11001 (N_11001,N_7285,N_8066);
xnor U11002 (N_11002,N_7871,N_6517);
and U11003 (N_11003,N_6538,N_6607);
nor U11004 (N_11004,N_8946,N_8168);
xor U11005 (N_11005,N_7150,N_6959);
xor U11006 (N_11006,N_8521,N_8545);
nor U11007 (N_11007,N_8334,N_7804);
nor U11008 (N_11008,N_7300,N_8031);
nand U11009 (N_11009,N_8175,N_8860);
nor U11010 (N_11010,N_8590,N_6513);
and U11011 (N_11011,N_7157,N_8536);
nor U11012 (N_11012,N_8763,N_6306);
and U11013 (N_11013,N_7940,N_8625);
xnor U11014 (N_11014,N_8384,N_6461);
and U11015 (N_11015,N_8657,N_7194);
nor U11016 (N_11016,N_8679,N_8642);
nor U11017 (N_11017,N_7695,N_8790);
nand U11018 (N_11018,N_6521,N_6643);
or U11019 (N_11019,N_7561,N_8017);
nand U11020 (N_11020,N_8676,N_6186);
nand U11021 (N_11021,N_6700,N_6791);
nor U11022 (N_11022,N_7473,N_8943);
and U11023 (N_11023,N_7405,N_6213);
nor U11024 (N_11024,N_8293,N_6680);
nand U11025 (N_11025,N_7777,N_6283);
xor U11026 (N_11026,N_8472,N_8718);
xor U11027 (N_11027,N_7111,N_6403);
xnor U11028 (N_11028,N_6127,N_7278);
xor U11029 (N_11029,N_8481,N_6473);
nand U11030 (N_11030,N_8229,N_8443);
or U11031 (N_11031,N_8508,N_8472);
and U11032 (N_11032,N_8183,N_8567);
nand U11033 (N_11033,N_6922,N_8052);
nand U11034 (N_11034,N_6344,N_8817);
or U11035 (N_11035,N_7796,N_6891);
or U11036 (N_11036,N_6213,N_7751);
nand U11037 (N_11037,N_8463,N_8620);
or U11038 (N_11038,N_6142,N_8585);
nor U11039 (N_11039,N_7555,N_8122);
and U11040 (N_11040,N_6864,N_7507);
nand U11041 (N_11041,N_8077,N_6128);
xnor U11042 (N_11042,N_6731,N_6676);
or U11043 (N_11043,N_6524,N_8032);
nor U11044 (N_11044,N_6390,N_6236);
or U11045 (N_11045,N_7774,N_8854);
nor U11046 (N_11046,N_6453,N_7874);
and U11047 (N_11047,N_7785,N_8521);
nand U11048 (N_11048,N_6961,N_6668);
or U11049 (N_11049,N_7753,N_7920);
and U11050 (N_11050,N_7622,N_6715);
nand U11051 (N_11051,N_8131,N_8004);
nand U11052 (N_11052,N_8842,N_7187);
xor U11053 (N_11053,N_8943,N_8100);
and U11054 (N_11054,N_8225,N_7835);
nor U11055 (N_11055,N_6974,N_7017);
nand U11056 (N_11056,N_6528,N_8100);
and U11057 (N_11057,N_7235,N_6468);
and U11058 (N_11058,N_7056,N_6132);
nand U11059 (N_11059,N_8384,N_8366);
nand U11060 (N_11060,N_7702,N_6062);
xor U11061 (N_11061,N_8183,N_6626);
xor U11062 (N_11062,N_7747,N_8940);
nand U11063 (N_11063,N_8415,N_8904);
nand U11064 (N_11064,N_7374,N_8620);
xnor U11065 (N_11065,N_7910,N_8216);
and U11066 (N_11066,N_6838,N_8313);
xor U11067 (N_11067,N_6852,N_8451);
and U11068 (N_11068,N_8172,N_8311);
nand U11069 (N_11069,N_6255,N_6887);
xnor U11070 (N_11070,N_6406,N_6252);
or U11071 (N_11071,N_8432,N_7248);
nand U11072 (N_11072,N_6849,N_7363);
nand U11073 (N_11073,N_7865,N_8799);
xnor U11074 (N_11074,N_8315,N_8654);
nor U11075 (N_11075,N_7678,N_6782);
or U11076 (N_11076,N_6254,N_8123);
and U11077 (N_11077,N_6735,N_6678);
and U11078 (N_11078,N_7146,N_7980);
or U11079 (N_11079,N_8291,N_6417);
or U11080 (N_11080,N_8803,N_7711);
xnor U11081 (N_11081,N_6275,N_7447);
nand U11082 (N_11082,N_6809,N_7636);
xnor U11083 (N_11083,N_6325,N_6408);
and U11084 (N_11084,N_8917,N_7883);
or U11085 (N_11085,N_8454,N_7318);
nand U11086 (N_11086,N_8157,N_6988);
nor U11087 (N_11087,N_7743,N_7829);
nand U11088 (N_11088,N_8828,N_7300);
or U11089 (N_11089,N_8460,N_7118);
xnor U11090 (N_11090,N_7251,N_7494);
or U11091 (N_11091,N_7956,N_7113);
nand U11092 (N_11092,N_7056,N_8223);
nor U11093 (N_11093,N_7219,N_7785);
nand U11094 (N_11094,N_7977,N_6810);
xnor U11095 (N_11095,N_6368,N_7207);
nor U11096 (N_11096,N_7667,N_8834);
or U11097 (N_11097,N_6768,N_6998);
nor U11098 (N_11098,N_7259,N_8929);
nor U11099 (N_11099,N_8671,N_6356);
and U11100 (N_11100,N_7493,N_6420);
and U11101 (N_11101,N_8581,N_8347);
xor U11102 (N_11102,N_6522,N_6532);
xor U11103 (N_11103,N_8455,N_7000);
nand U11104 (N_11104,N_7587,N_6632);
or U11105 (N_11105,N_6433,N_7264);
and U11106 (N_11106,N_6626,N_6427);
and U11107 (N_11107,N_6536,N_8467);
and U11108 (N_11108,N_7405,N_8445);
nand U11109 (N_11109,N_6151,N_7601);
xor U11110 (N_11110,N_6833,N_8193);
or U11111 (N_11111,N_7872,N_8534);
nand U11112 (N_11112,N_6295,N_6278);
or U11113 (N_11113,N_7295,N_8202);
and U11114 (N_11114,N_8444,N_8928);
xor U11115 (N_11115,N_6983,N_7731);
and U11116 (N_11116,N_8686,N_8038);
nor U11117 (N_11117,N_7912,N_6450);
nand U11118 (N_11118,N_6425,N_7482);
and U11119 (N_11119,N_8625,N_8531);
or U11120 (N_11120,N_6799,N_8007);
and U11121 (N_11121,N_6291,N_6764);
xor U11122 (N_11122,N_8561,N_7257);
and U11123 (N_11123,N_8855,N_8881);
nand U11124 (N_11124,N_6429,N_7145);
and U11125 (N_11125,N_8204,N_6924);
and U11126 (N_11126,N_7616,N_8511);
xor U11127 (N_11127,N_8195,N_6352);
xnor U11128 (N_11128,N_6943,N_8889);
and U11129 (N_11129,N_7136,N_7768);
or U11130 (N_11130,N_7037,N_6533);
nor U11131 (N_11131,N_6669,N_6140);
xnor U11132 (N_11132,N_8519,N_8081);
nand U11133 (N_11133,N_7456,N_7553);
xnor U11134 (N_11134,N_6288,N_8632);
or U11135 (N_11135,N_6226,N_6058);
xnor U11136 (N_11136,N_7284,N_6201);
or U11137 (N_11137,N_7095,N_7879);
xnor U11138 (N_11138,N_6970,N_8293);
nand U11139 (N_11139,N_7321,N_6799);
and U11140 (N_11140,N_6583,N_6427);
xor U11141 (N_11141,N_7735,N_6182);
nor U11142 (N_11142,N_6837,N_6398);
xor U11143 (N_11143,N_8870,N_8494);
or U11144 (N_11144,N_6342,N_7426);
nor U11145 (N_11145,N_7435,N_8311);
nor U11146 (N_11146,N_7411,N_6331);
xnor U11147 (N_11147,N_8875,N_6207);
nor U11148 (N_11148,N_6994,N_7412);
xnor U11149 (N_11149,N_7015,N_6498);
nor U11150 (N_11150,N_7389,N_7274);
nor U11151 (N_11151,N_6802,N_6511);
nor U11152 (N_11152,N_6843,N_6362);
xor U11153 (N_11153,N_8365,N_8662);
and U11154 (N_11154,N_8612,N_8386);
xnor U11155 (N_11155,N_6631,N_8651);
or U11156 (N_11156,N_6789,N_7227);
and U11157 (N_11157,N_7918,N_7478);
nor U11158 (N_11158,N_8969,N_7782);
nor U11159 (N_11159,N_7431,N_7922);
or U11160 (N_11160,N_7834,N_8660);
nor U11161 (N_11161,N_7951,N_7051);
xor U11162 (N_11162,N_6239,N_6761);
and U11163 (N_11163,N_7346,N_8808);
nor U11164 (N_11164,N_8664,N_6498);
nor U11165 (N_11165,N_6625,N_7355);
xnor U11166 (N_11166,N_6463,N_8627);
xor U11167 (N_11167,N_7154,N_8873);
nand U11168 (N_11168,N_6905,N_7602);
or U11169 (N_11169,N_7777,N_8319);
nor U11170 (N_11170,N_8818,N_6856);
and U11171 (N_11171,N_6328,N_7062);
or U11172 (N_11172,N_7695,N_7386);
nand U11173 (N_11173,N_6305,N_7061);
or U11174 (N_11174,N_7378,N_6519);
xnor U11175 (N_11175,N_7101,N_6053);
nor U11176 (N_11176,N_6002,N_7616);
or U11177 (N_11177,N_6992,N_8975);
and U11178 (N_11178,N_6020,N_6946);
xnor U11179 (N_11179,N_6382,N_6332);
xor U11180 (N_11180,N_8961,N_8056);
nand U11181 (N_11181,N_7801,N_6086);
and U11182 (N_11182,N_7531,N_6259);
xnor U11183 (N_11183,N_8996,N_8657);
xor U11184 (N_11184,N_6669,N_7284);
nand U11185 (N_11185,N_7336,N_8920);
nand U11186 (N_11186,N_6808,N_8402);
nor U11187 (N_11187,N_7733,N_8405);
and U11188 (N_11188,N_8872,N_8673);
and U11189 (N_11189,N_7104,N_8182);
or U11190 (N_11190,N_7394,N_7669);
nor U11191 (N_11191,N_7994,N_8248);
or U11192 (N_11192,N_6099,N_7695);
and U11193 (N_11193,N_7460,N_8571);
nand U11194 (N_11194,N_6731,N_8526);
xnor U11195 (N_11195,N_6132,N_8323);
and U11196 (N_11196,N_8148,N_6968);
or U11197 (N_11197,N_8445,N_6363);
nand U11198 (N_11198,N_8081,N_6806);
nor U11199 (N_11199,N_7050,N_8545);
xnor U11200 (N_11200,N_6085,N_6611);
and U11201 (N_11201,N_8660,N_6835);
xnor U11202 (N_11202,N_6679,N_6166);
and U11203 (N_11203,N_7626,N_8694);
nand U11204 (N_11204,N_8330,N_8894);
xor U11205 (N_11205,N_6478,N_7306);
xor U11206 (N_11206,N_7059,N_7210);
or U11207 (N_11207,N_8610,N_7604);
xor U11208 (N_11208,N_7485,N_8493);
nand U11209 (N_11209,N_7164,N_6306);
nand U11210 (N_11210,N_8012,N_6427);
and U11211 (N_11211,N_6247,N_7178);
and U11212 (N_11212,N_6182,N_6425);
nor U11213 (N_11213,N_7235,N_8160);
nand U11214 (N_11214,N_6173,N_6101);
nor U11215 (N_11215,N_7853,N_6439);
and U11216 (N_11216,N_8332,N_7466);
nor U11217 (N_11217,N_8275,N_8367);
or U11218 (N_11218,N_8082,N_8594);
nand U11219 (N_11219,N_7067,N_8742);
or U11220 (N_11220,N_7980,N_7762);
nor U11221 (N_11221,N_7143,N_6338);
xnor U11222 (N_11222,N_7353,N_8459);
or U11223 (N_11223,N_8016,N_8346);
xor U11224 (N_11224,N_8198,N_7985);
nor U11225 (N_11225,N_8819,N_7931);
and U11226 (N_11226,N_7944,N_8465);
and U11227 (N_11227,N_6361,N_8068);
or U11228 (N_11228,N_6237,N_8778);
nor U11229 (N_11229,N_6690,N_8186);
and U11230 (N_11230,N_8366,N_8612);
and U11231 (N_11231,N_8933,N_7172);
or U11232 (N_11232,N_6385,N_8266);
nand U11233 (N_11233,N_6728,N_7758);
and U11234 (N_11234,N_7397,N_7713);
and U11235 (N_11235,N_6753,N_8841);
or U11236 (N_11236,N_6327,N_6473);
xnor U11237 (N_11237,N_6546,N_6982);
nor U11238 (N_11238,N_8286,N_6947);
xnor U11239 (N_11239,N_7883,N_7798);
and U11240 (N_11240,N_7549,N_6104);
and U11241 (N_11241,N_8286,N_7823);
nor U11242 (N_11242,N_8411,N_6184);
nor U11243 (N_11243,N_6332,N_8519);
and U11244 (N_11244,N_7056,N_7240);
xor U11245 (N_11245,N_7198,N_7183);
xnor U11246 (N_11246,N_6563,N_8804);
or U11247 (N_11247,N_6879,N_8913);
xnor U11248 (N_11248,N_8737,N_6591);
xnor U11249 (N_11249,N_7100,N_7860);
and U11250 (N_11250,N_8350,N_8359);
nand U11251 (N_11251,N_6627,N_7501);
or U11252 (N_11252,N_6990,N_6123);
and U11253 (N_11253,N_6750,N_8077);
and U11254 (N_11254,N_6677,N_8750);
nand U11255 (N_11255,N_8779,N_7096);
or U11256 (N_11256,N_8119,N_7075);
or U11257 (N_11257,N_6071,N_7016);
and U11258 (N_11258,N_8583,N_6719);
nand U11259 (N_11259,N_6128,N_7036);
nand U11260 (N_11260,N_7680,N_8878);
xor U11261 (N_11261,N_7646,N_7304);
xor U11262 (N_11262,N_6047,N_6985);
and U11263 (N_11263,N_7854,N_6910);
nand U11264 (N_11264,N_8266,N_7122);
and U11265 (N_11265,N_8832,N_7371);
nand U11266 (N_11266,N_6713,N_6133);
and U11267 (N_11267,N_7720,N_7051);
nor U11268 (N_11268,N_8611,N_7068);
and U11269 (N_11269,N_7742,N_8674);
nor U11270 (N_11270,N_7642,N_8282);
xnor U11271 (N_11271,N_6093,N_7320);
and U11272 (N_11272,N_8437,N_7248);
and U11273 (N_11273,N_7131,N_6643);
and U11274 (N_11274,N_7164,N_8468);
or U11275 (N_11275,N_8669,N_8041);
or U11276 (N_11276,N_8414,N_6498);
or U11277 (N_11277,N_7749,N_8696);
and U11278 (N_11278,N_8152,N_7289);
nand U11279 (N_11279,N_8645,N_8569);
xor U11280 (N_11280,N_8732,N_8501);
and U11281 (N_11281,N_8766,N_7124);
or U11282 (N_11282,N_8504,N_6388);
xnor U11283 (N_11283,N_7531,N_8332);
or U11284 (N_11284,N_6352,N_7517);
or U11285 (N_11285,N_8694,N_6998);
and U11286 (N_11286,N_7492,N_7543);
or U11287 (N_11287,N_8173,N_7262);
xnor U11288 (N_11288,N_8668,N_7777);
nor U11289 (N_11289,N_6683,N_7409);
and U11290 (N_11290,N_7408,N_8581);
and U11291 (N_11291,N_7125,N_8751);
xor U11292 (N_11292,N_6081,N_8092);
nor U11293 (N_11293,N_6211,N_8213);
nand U11294 (N_11294,N_8031,N_8532);
or U11295 (N_11295,N_7770,N_6094);
xnor U11296 (N_11296,N_7395,N_8850);
xor U11297 (N_11297,N_7901,N_8714);
nor U11298 (N_11298,N_7669,N_8131);
xnor U11299 (N_11299,N_8838,N_6991);
xor U11300 (N_11300,N_6784,N_6592);
or U11301 (N_11301,N_6526,N_7008);
nor U11302 (N_11302,N_6590,N_8160);
and U11303 (N_11303,N_8239,N_8118);
nor U11304 (N_11304,N_8097,N_7514);
and U11305 (N_11305,N_7462,N_8307);
nor U11306 (N_11306,N_8944,N_8059);
xnor U11307 (N_11307,N_7137,N_6761);
xor U11308 (N_11308,N_6625,N_8547);
nor U11309 (N_11309,N_6574,N_7563);
xor U11310 (N_11310,N_6461,N_8289);
nor U11311 (N_11311,N_6291,N_7399);
nor U11312 (N_11312,N_7003,N_6451);
nor U11313 (N_11313,N_8950,N_7822);
xnor U11314 (N_11314,N_7043,N_7819);
and U11315 (N_11315,N_6492,N_7922);
xnor U11316 (N_11316,N_6695,N_7819);
xnor U11317 (N_11317,N_7978,N_7937);
nand U11318 (N_11318,N_6783,N_7661);
nor U11319 (N_11319,N_8662,N_7160);
or U11320 (N_11320,N_6387,N_6641);
nor U11321 (N_11321,N_8990,N_7372);
xnor U11322 (N_11322,N_8963,N_6248);
and U11323 (N_11323,N_6658,N_6590);
or U11324 (N_11324,N_6048,N_7376);
and U11325 (N_11325,N_8532,N_6186);
nand U11326 (N_11326,N_6854,N_6108);
nor U11327 (N_11327,N_8201,N_8741);
and U11328 (N_11328,N_8789,N_7727);
xnor U11329 (N_11329,N_7209,N_7072);
xnor U11330 (N_11330,N_6943,N_8931);
nand U11331 (N_11331,N_8650,N_8629);
nand U11332 (N_11332,N_7499,N_6767);
and U11333 (N_11333,N_7436,N_6261);
nor U11334 (N_11334,N_6720,N_6178);
nor U11335 (N_11335,N_7093,N_8228);
xor U11336 (N_11336,N_7029,N_6895);
xor U11337 (N_11337,N_6800,N_8815);
nor U11338 (N_11338,N_8168,N_6911);
nand U11339 (N_11339,N_8993,N_8547);
xnor U11340 (N_11340,N_8407,N_6096);
nand U11341 (N_11341,N_8438,N_7172);
or U11342 (N_11342,N_6272,N_6393);
nor U11343 (N_11343,N_6647,N_8275);
and U11344 (N_11344,N_6878,N_8386);
nor U11345 (N_11345,N_6613,N_8677);
xnor U11346 (N_11346,N_8351,N_7097);
nand U11347 (N_11347,N_6113,N_8469);
nand U11348 (N_11348,N_7937,N_7532);
nor U11349 (N_11349,N_7364,N_6218);
xor U11350 (N_11350,N_6947,N_7322);
nand U11351 (N_11351,N_6796,N_6561);
xnor U11352 (N_11352,N_8152,N_8445);
xor U11353 (N_11353,N_6172,N_6596);
nor U11354 (N_11354,N_7521,N_6683);
and U11355 (N_11355,N_7072,N_8609);
or U11356 (N_11356,N_8916,N_7584);
nand U11357 (N_11357,N_6100,N_6317);
nor U11358 (N_11358,N_8116,N_7094);
nand U11359 (N_11359,N_6671,N_6689);
or U11360 (N_11360,N_6132,N_8774);
xnor U11361 (N_11361,N_6735,N_7638);
nand U11362 (N_11362,N_8064,N_8505);
nand U11363 (N_11363,N_8107,N_7023);
nand U11364 (N_11364,N_7485,N_6596);
or U11365 (N_11365,N_7717,N_7407);
or U11366 (N_11366,N_6115,N_6499);
and U11367 (N_11367,N_8354,N_7688);
nand U11368 (N_11368,N_6290,N_6852);
or U11369 (N_11369,N_7785,N_7128);
nor U11370 (N_11370,N_8380,N_6814);
nor U11371 (N_11371,N_7810,N_6354);
nor U11372 (N_11372,N_8542,N_6856);
or U11373 (N_11373,N_6840,N_8032);
nor U11374 (N_11374,N_6953,N_8571);
nor U11375 (N_11375,N_6749,N_6886);
and U11376 (N_11376,N_8318,N_7234);
nand U11377 (N_11377,N_8536,N_6147);
xnor U11378 (N_11378,N_8285,N_8602);
nor U11379 (N_11379,N_6885,N_7012);
or U11380 (N_11380,N_8529,N_8401);
or U11381 (N_11381,N_7737,N_8148);
or U11382 (N_11382,N_7094,N_6567);
xnor U11383 (N_11383,N_8454,N_7767);
or U11384 (N_11384,N_7259,N_8572);
nand U11385 (N_11385,N_8200,N_7995);
xor U11386 (N_11386,N_6297,N_8074);
or U11387 (N_11387,N_8552,N_7980);
nor U11388 (N_11388,N_8653,N_6504);
xnor U11389 (N_11389,N_6550,N_7222);
xnor U11390 (N_11390,N_6138,N_6043);
nand U11391 (N_11391,N_7186,N_6196);
and U11392 (N_11392,N_8765,N_6171);
nor U11393 (N_11393,N_8023,N_6126);
xor U11394 (N_11394,N_8049,N_6784);
and U11395 (N_11395,N_8501,N_7596);
and U11396 (N_11396,N_6710,N_6862);
and U11397 (N_11397,N_6500,N_6897);
nand U11398 (N_11398,N_6850,N_7814);
nand U11399 (N_11399,N_7333,N_6242);
or U11400 (N_11400,N_7561,N_6921);
xnor U11401 (N_11401,N_7954,N_8852);
or U11402 (N_11402,N_8357,N_8054);
nand U11403 (N_11403,N_7017,N_8770);
and U11404 (N_11404,N_6448,N_8378);
nand U11405 (N_11405,N_7154,N_6261);
nand U11406 (N_11406,N_8294,N_6671);
nor U11407 (N_11407,N_6131,N_7848);
xor U11408 (N_11408,N_7119,N_8712);
xnor U11409 (N_11409,N_6340,N_7162);
xnor U11410 (N_11410,N_8769,N_7354);
and U11411 (N_11411,N_8058,N_6911);
and U11412 (N_11412,N_7433,N_7908);
xor U11413 (N_11413,N_6477,N_7751);
nand U11414 (N_11414,N_8564,N_6244);
and U11415 (N_11415,N_8088,N_8199);
xor U11416 (N_11416,N_7561,N_8360);
or U11417 (N_11417,N_8666,N_8056);
nand U11418 (N_11418,N_8774,N_6044);
nand U11419 (N_11419,N_6520,N_6856);
xnor U11420 (N_11420,N_6983,N_8280);
or U11421 (N_11421,N_6396,N_7344);
nor U11422 (N_11422,N_6505,N_7727);
nor U11423 (N_11423,N_7662,N_6536);
nor U11424 (N_11424,N_7601,N_8611);
nand U11425 (N_11425,N_8748,N_8802);
and U11426 (N_11426,N_6856,N_6177);
nand U11427 (N_11427,N_8264,N_8641);
and U11428 (N_11428,N_8007,N_8521);
xnor U11429 (N_11429,N_8058,N_6976);
xnor U11430 (N_11430,N_6456,N_6925);
and U11431 (N_11431,N_6995,N_8355);
xnor U11432 (N_11432,N_7999,N_8503);
or U11433 (N_11433,N_6465,N_8197);
or U11434 (N_11434,N_7710,N_8155);
nand U11435 (N_11435,N_6602,N_6527);
nand U11436 (N_11436,N_6451,N_6226);
or U11437 (N_11437,N_7995,N_8276);
nand U11438 (N_11438,N_6569,N_6357);
nand U11439 (N_11439,N_7892,N_8111);
or U11440 (N_11440,N_7776,N_8158);
nand U11441 (N_11441,N_8625,N_8993);
or U11442 (N_11442,N_8585,N_8661);
nand U11443 (N_11443,N_6557,N_6110);
nand U11444 (N_11444,N_7029,N_7408);
nor U11445 (N_11445,N_8935,N_8399);
or U11446 (N_11446,N_8262,N_6672);
xor U11447 (N_11447,N_7495,N_8634);
or U11448 (N_11448,N_7365,N_6005);
xor U11449 (N_11449,N_8868,N_7892);
or U11450 (N_11450,N_6225,N_6915);
nand U11451 (N_11451,N_7105,N_7114);
nand U11452 (N_11452,N_7655,N_8367);
xnor U11453 (N_11453,N_7103,N_8690);
xor U11454 (N_11454,N_8837,N_8489);
nor U11455 (N_11455,N_7461,N_8977);
nor U11456 (N_11456,N_8276,N_6194);
xnor U11457 (N_11457,N_8454,N_6435);
nand U11458 (N_11458,N_7447,N_7557);
or U11459 (N_11459,N_8151,N_7649);
or U11460 (N_11460,N_6078,N_6657);
xnor U11461 (N_11461,N_6446,N_8257);
and U11462 (N_11462,N_8762,N_6801);
nand U11463 (N_11463,N_6045,N_7255);
or U11464 (N_11464,N_7654,N_8829);
or U11465 (N_11465,N_6297,N_6613);
xor U11466 (N_11466,N_7533,N_6166);
nand U11467 (N_11467,N_7158,N_6128);
nand U11468 (N_11468,N_6368,N_7927);
or U11469 (N_11469,N_7306,N_8703);
or U11470 (N_11470,N_7604,N_7897);
xor U11471 (N_11471,N_6201,N_8141);
or U11472 (N_11472,N_8961,N_7384);
xor U11473 (N_11473,N_8062,N_6001);
or U11474 (N_11474,N_8710,N_7179);
or U11475 (N_11475,N_7825,N_7193);
nand U11476 (N_11476,N_6663,N_7480);
nor U11477 (N_11477,N_8927,N_6881);
xnor U11478 (N_11478,N_6964,N_6290);
nand U11479 (N_11479,N_7323,N_6114);
nand U11480 (N_11480,N_8766,N_7431);
or U11481 (N_11481,N_8363,N_6034);
or U11482 (N_11482,N_8013,N_6547);
and U11483 (N_11483,N_6639,N_6848);
nand U11484 (N_11484,N_6577,N_8661);
or U11485 (N_11485,N_8079,N_7691);
nand U11486 (N_11486,N_7051,N_8196);
nand U11487 (N_11487,N_6415,N_8212);
nor U11488 (N_11488,N_7432,N_6259);
and U11489 (N_11489,N_8254,N_8641);
xor U11490 (N_11490,N_8997,N_8078);
or U11491 (N_11491,N_6998,N_7146);
nor U11492 (N_11492,N_7554,N_7480);
nor U11493 (N_11493,N_7263,N_6675);
nand U11494 (N_11494,N_8391,N_8581);
or U11495 (N_11495,N_7016,N_6373);
nor U11496 (N_11496,N_7847,N_8553);
and U11497 (N_11497,N_8245,N_6710);
nand U11498 (N_11498,N_8053,N_6107);
nor U11499 (N_11499,N_8769,N_6619);
xor U11500 (N_11500,N_7542,N_6264);
nor U11501 (N_11501,N_7823,N_6683);
or U11502 (N_11502,N_8572,N_8926);
xnor U11503 (N_11503,N_7270,N_8808);
xnor U11504 (N_11504,N_8699,N_7860);
nand U11505 (N_11505,N_7247,N_8572);
xnor U11506 (N_11506,N_7962,N_7161);
nand U11507 (N_11507,N_7695,N_7632);
or U11508 (N_11508,N_8772,N_6911);
xor U11509 (N_11509,N_7442,N_8874);
and U11510 (N_11510,N_6298,N_7027);
nand U11511 (N_11511,N_7897,N_7787);
nor U11512 (N_11512,N_8901,N_8783);
and U11513 (N_11513,N_6058,N_8120);
nand U11514 (N_11514,N_8898,N_8373);
nor U11515 (N_11515,N_8606,N_6768);
or U11516 (N_11516,N_7543,N_8766);
xnor U11517 (N_11517,N_6619,N_8229);
nand U11518 (N_11518,N_7291,N_8826);
nand U11519 (N_11519,N_7329,N_8528);
nor U11520 (N_11520,N_8353,N_6796);
nor U11521 (N_11521,N_8193,N_7527);
nor U11522 (N_11522,N_7616,N_6442);
nor U11523 (N_11523,N_8685,N_8050);
nand U11524 (N_11524,N_7951,N_6375);
xor U11525 (N_11525,N_8304,N_7608);
and U11526 (N_11526,N_6196,N_7072);
nand U11527 (N_11527,N_6736,N_8924);
xnor U11528 (N_11528,N_7420,N_8187);
nand U11529 (N_11529,N_8489,N_6473);
nor U11530 (N_11530,N_8842,N_8158);
nand U11531 (N_11531,N_8108,N_8037);
and U11532 (N_11532,N_8455,N_6555);
and U11533 (N_11533,N_8047,N_8258);
nand U11534 (N_11534,N_8898,N_8942);
and U11535 (N_11535,N_7347,N_7564);
nand U11536 (N_11536,N_7052,N_8101);
nor U11537 (N_11537,N_7848,N_8591);
xor U11538 (N_11538,N_8982,N_7062);
nor U11539 (N_11539,N_6880,N_6869);
nand U11540 (N_11540,N_6042,N_7197);
or U11541 (N_11541,N_8284,N_7474);
nor U11542 (N_11542,N_7272,N_6526);
nand U11543 (N_11543,N_8572,N_6961);
xnor U11544 (N_11544,N_6396,N_8247);
xnor U11545 (N_11545,N_7641,N_7074);
nor U11546 (N_11546,N_6551,N_8641);
xor U11547 (N_11547,N_8861,N_7036);
xnor U11548 (N_11548,N_7212,N_8011);
xor U11549 (N_11549,N_6714,N_8932);
nand U11550 (N_11550,N_6223,N_6828);
xor U11551 (N_11551,N_7539,N_8139);
or U11552 (N_11552,N_8485,N_7147);
or U11553 (N_11553,N_7846,N_7682);
or U11554 (N_11554,N_6438,N_6922);
xnor U11555 (N_11555,N_7059,N_7816);
or U11556 (N_11556,N_7806,N_7730);
and U11557 (N_11557,N_8289,N_8306);
or U11558 (N_11558,N_8592,N_7321);
nand U11559 (N_11559,N_8529,N_7024);
nand U11560 (N_11560,N_6608,N_7188);
or U11561 (N_11561,N_6649,N_6330);
nor U11562 (N_11562,N_6942,N_8421);
nor U11563 (N_11563,N_6763,N_6736);
xnor U11564 (N_11564,N_7365,N_8257);
xnor U11565 (N_11565,N_8764,N_6358);
nor U11566 (N_11566,N_8345,N_8440);
nor U11567 (N_11567,N_7238,N_7456);
or U11568 (N_11568,N_6070,N_7563);
xor U11569 (N_11569,N_7054,N_8410);
nor U11570 (N_11570,N_6020,N_6471);
nor U11571 (N_11571,N_8376,N_7715);
nor U11572 (N_11572,N_7684,N_8965);
or U11573 (N_11573,N_6315,N_6446);
nand U11574 (N_11574,N_6695,N_8198);
or U11575 (N_11575,N_8474,N_8435);
nand U11576 (N_11576,N_6803,N_8970);
xnor U11577 (N_11577,N_8411,N_7263);
nor U11578 (N_11578,N_8967,N_7077);
and U11579 (N_11579,N_7167,N_6368);
or U11580 (N_11580,N_6239,N_6070);
nor U11581 (N_11581,N_7328,N_7640);
or U11582 (N_11582,N_6928,N_6096);
and U11583 (N_11583,N_7282,N_8175);
or U11584 (N_11584,N_7633,N_6128);
xor U11585 (N_11585,N_8299,N_8006);
and U11586 (N_11586,N_6145,N_8702);
and U11587 (N_11587,N_6899,N_7298);
nand U11588 (N_11588,N_6090,N_8817);
xnor U11589 (N_11589,N_6585,N_8686);
and U11590 (N_11590,N_6150,N_8399);
xnor U11591 (N_11591,N_7246,N_7532);
nand U11592 (N_11592,N_6236,N_8451);
nor U11593 (N_11593,N_6535,N_8104);
xnor U11594 (N_11594,N_8508,N_6894);
and U11595 (N_11595,N_6159,N_7034);
nand U11596 (N_11596,N_8354,N_6853);
and U11597 (N_11597,N_7980,N_6628);
nand U11598 (N_11598,N_8857,N_6039);
nor U11599 (N_11599,N_6221,N_8975);
xor U11600 (N_11600,N_6023,N_6608);
nor U11601 (N_11601,N_7088,N_8453);
and U11602 (N_11602,N_7613,N_8290);
xor U11603 (N_11603,N_8535,N_8814);
nand U11604 (N_11604,N_8425,N_8645);
or U11605 (N_11605,N_8006,N_8247);
nor U11606 (N_11606,N_8268,N_6790);
nand U11607 (N_11607,N_6669,N_7945);
and U11608 (N_11608,N_6195,N_8412);
xor U11609 (N_11609,N_6979,N_6927);
xor U11610 (N_11610,N_6887,N_8209);
or U11611 (N_11611,N_8889,N_6799);
and U11612 (N_11612,N_8157,N_8546);
xor U11613 (N_11613,N_8712,N_6389);
and U11614 (N_11614,N_8670,N_7168);
nand U11615 (N_11615,N_7717,N_7689);
nor U11616 (N_11616,N_7356,N_6107);
and U11617 (N_11617,N_7081,N_8604);
or U11618 (N_11618,N_7764,N_6188);
or U11619 (N_11619,N_8859,N_8397);
nor U11620 (N_11620,N_6040,N_7820);
or U11621 (N_11621,N_8401,N_7919);
and U11622 (N_11622,N_8625,N_8881);
or U11623 (N_11623,N_6120,N_6919);
and U11624 (N_11624,N_6612,N_6074);
nor U11625 (N_11625,N_6011,N_7419);
nor U11626 (N_11626,N_8265,N_7586);
or U11627 (N_11627,N_6449,N_8666);
or U11628 (N_11628,N_8284,N_7947);
or U11629 (N_11629,N_8634,N_8946);
nand U11630 (N_11630,N_6985,N_7896);
nand U11631 (N_11631,N_8958,N_8468);
xor U11632 (N_11632,N_6511,N_6846);
nand U11633 (N_11633,N_7905,N_6296);
nand U11634 (N_11634,N_7441,N_7000);
xor U11635 (N_11635,N_6048,N_6808);
and U11636 (N_11636,N_8146,N_8557);
and U11637 (N_11637,N_7891,N_6849);
xnor U11638 (N_11638,N_7063,N_8252);
and U11639 (N_11639,N_7721,N_8774);
nor U11640 (N_11640,N_8457,N_8519);
xor U11641 (N_11641,N_7322,N_6856);
nor U11642 (N_11642,N_8177,N_6250);
xnor U11643 (N_11643,N_8088,N_8499);
and U11644 (N_11644,N_8010,N_8998);
or U11645 (N_11645,N_7723,N_7407);
and U11646 (N_11646,N_6193,N_7898);
or U11647 (N_11647,N_7619,N_7773);
xor U11648 (N_11648,N_6903,N_6766);
nand U11649 (N_11649,N_8672,N_8342);
nor U11650 (N_11650,N_8944,N_7499);
nor U11651 (N_11651,N_6755,N_6864);
nor U11652 (N_11652,N_8320,N_6118);
or U11653 (N_11653,N_8712,N_8190);
nor U11654 (N_11654,N_7168,N_6122);
and U11655 (N_11655,N_6456,N_7719);
nor U11656 (N_11656,N_8223,N_7157);
nor U11657 (N_11657,N_6319,N_7666);
xnor U11658 (N_11658,N_7231,N_6542);
nand U11659 (N_11659,N_6116,N_7965);
nor U11660 (N_11660,N_8363,N_8383);
or U11661 (N_11661,N_8445,N_8109);
or U11662 (N_11662,N_6658,N_6772);
nor U11663 (N_11663,N_8982,N_8368);
nand U11664 (N_11664,N_7733,N_6540);
or U11665 (N_11665,N_8516,N_8720);
nand U11666 (N_11666,N_6371,N_6458);
nand U11667 (N_11667,N_6577,N_7310);
nand U11668 (N_11668,N_6584,N_6696);
or U11669 (N_11669,N_8606,N_6315);
and U11670 (N_11670,N_6969,N_6332);
or U11671 (N_11671,N_7523,N_8025);
and U11672 (N_11672,N_6190,N_7281);
xor U11673 (N_11673,N_6593,N_7513);
and U11674 (N_11674,N_6047,N_6317);
nor U11675 (N_11675,N_7899,N_6096);
xor U11676 (N_11676,N_8192,N_6638);
and U11677 (N_11677,N_7572,N_7368);
nor U11678 (N_11678,N_6616,N_8181);
nand U11679 (N_11679,N_7566,N_6858);
or U11680 (N_11680,N_6538,N_8194);
nor U11681 (N_11681,N_6410,N_7569);
xor U11682 (N_11682,N_8400,N_6756);
nor U11683 (N_11683,N_7197,N_6541);
nand U11684 (N_11684,N_7964,N_7819);
nor U11685 (N_11685,N_6939,N_6957);
xnor U11686 (N_11686,N_8171,N_6690);
xnor U11687 (N_11687,N_6468,N_8907);
and U11688 (N_11688,N_7720,N_6998);
nor U11689 (N_11689,N_6508,N_8708);
nor U11690 (N_11690,N_6367,N_7594);
nand U11691 (N_11691,N_6088,N_8475);
or U11692 (N_11692,N_8034,N_7233);
nor U11693 (N_11693,N_6467,N_6283);
xnor U11694 (N_11694,N_8131,N_8297);
xor U11695 (N_11695,N_7287,N_8300);
or U11696 (N_11696,N_8974,N_8559);
nand U11697 (N_11697,N_7033,N_7603);
nor U11698 (N_11698,N_7005,N_6283);
nor U11699 (N_11699,N_7017,N_7058);
nor U11700 (N_11700,N_6404,N_7578);
nor U11701 (N_11701,N_8144,N_6970);
and U11702 (N_11702,N_8042,N_8928);
xnor U11703 (N_11703,N_6692,N_8726);
xnor U11704 (N_11704,N_8105,N_8920);
and U11705 (N_11705,N_6326,N_6746);
xor U11706 (N_11706,N_8401,N_7075);
xnor U11707 (N_11707,N_6303,N_8776);
xnor U11708 (N_11708,N_8202,N_7361);
or U11709 (N_11709,N_8530,N_6283);
xnor U11710 (N_11710,N_8676,N_6445);
and U11711 (N_11711,N_8885,N_8363);
and U11712 (N_11712,N_6220,N_7001);
and U11713 (N_11713,N_6010,N_6615);
nand U11714 (N_11714,N_6765,N_8496);
xor U11715 (N_11715,N_7242,N_8446);
and U11716 (N_11716,N_7204,N_6597);
nor U11717 (N_11717,N_6854,N_8011);
nor U11718 (N_11718,N_7611,N_7504);
nor U11719 (N_11719,N_6885,N_8157);
xnor U11720 (N_11720,N_8231,N_8634);
or U11721 (N_11721,N_6467,N_7009);
nand U11722 (N_11722,N_6101,N_7326);
nor U11723 (N_11723,N_7323,N_8307);
nor U11724 (N_11724,N_6643,N_7295);
nand U11725 (N_11725,N_6894,N_6203);
nand U11726 (N_11726,N_8811,N_6034);
or U11727 (N_11727,N_7794,N_7335);
nand U11728 (N_11728,N_8205,N_7361);
and U11729 (N_11729,N_8809,N_6815);
nor U11730 (N_11730,N_7290,N_6753);
xnor U11731 (N_11731,N_6371,N_7073);
or U11732 (N_11732,N_6920,N_7353);
nand U11733 (N_11733,N_8619,N_8827);
or U11734 (N_11734,N_8753,N_8308);
xor U11735 (N_11735,N_7078,N_6425);
nand U11736 (N_11736,N_8926,N_7283);
xnor U11737 (N_11737,N_7405,N_6324);
or U11738 (N_11738,N_7802,N_8274);
xor U11739 (N_11739,N_6289,N_8434);
or U11740 (N_11740,N_6713,N_6314);
and U11741 (N_11741,N_6893,N_6297);
and U11742 (N_11742,N_6544,N_8253);
nor U11743 (N_11743,N_6910,N_7286);
nor U11744 (N_11744,N_6857,N_8155);
nand U11745 (N_11745,N_6774,N_7695);
or U11746 (N_11746,N_6521,N_7008);
nand U11747 (N_11747,N_6158,N_7853);
xor U11748 (N_11748,N_8409,N_7134);
nor U11749 (N_11749,N_8641,N_6146);
xnor U11750 (N_11750,N_7233,N_6180);
xor U11751 (N_11751,N_7742,N_7626);
and U11752 (N_11752,N_8647,N_7924);
xor U11753 (N_11753,N_6570,N_6764);
and U11754 (N_11754,N_8400,N_6601);
nand U11755 (N_11755,N_6385,N_6564);
and U11756 (N_11756,N_8225,N_7174);
nor U11757 (N_11757,N_8134,N_7087);
nor U11758 (N_11758,N_6468,N_7385);
nor U11759 (N_11759,N_8745,N_6939);
nand U11760 (N_11760,N_7702,N_8060);
nand U11761 (N_11761,N_6375,N_8839);
and U11762 (N_11762,N_8482,N_6414);
nand U11763 (N_11763,N_8229,N_7755);
xnor U11764 (N_11764,N_6575,N_6665);
or U11765 (N_11765,N_7712,N_8144);
nand U11766 (N_11766,N_7161,N_7944);
xor U11767 (N_11767,N_6396,N_7104);
or U11768 (N_11768,N_6115,N_7109);
and U11769 (N_11769,N_6840,N_6948);
and U11770 (N_11770,N_8318,N_6353);
xnor U11771 (N_11771,N_6867,N_8876);
nand U11772 (N_11772,N_6110,N_7951);
xnor U11773 (N_11773,N_7268,N_8456);
nor U11774 (N_11774,N_7834,N_8263);
or U11775 (N_11775,N_8576,N_6766);
nand U11776 (N_11776,N_6005,N_8566);
xor U11777 (N_11777,N_8328,N_7597);
nand U11778 (N_11778,N_6200,N_7871);
nor U11779 (N_11779,N_7063,N_6230);
and U11780 (N_11780,N_8409,N_7173);
xor U11781 (N_11781,N_7977,N_7129);
nor U11782 (N_11782,N_6683,N_6982);
nand U11783 (N_11783,N_8539,N_6034);
xnor U11784 (N_11784,N_6598,N_8605);
and U11785 (N_11785,N_8170,N_6701);
xor U11786 (N_11786,N_6530,N_6520);
xnor U11787 (N_11787,N_7406,N_7681);
xor U11788 (N_11788,N_7518,N_8672);
or U11789 (N_11789,N_8480,N_8592);
nor U11790 (N_11790,N_6459,N_7053);
xor U11791 (N_11791,N_6101,N_6718);
or U11792 (N_11792,N_6983,N_7718);
xnor U11793 (N_11793,N_6557,N_8661);
nand U11794 (N_11794,N_8359,N_6920);
nand U11795 (N_11795,N_8974,N_6794);
xnor U11796 (N_11796,N_7349,N_7318);
and U11797 (N_11797,N_7440,N_6633);
and U11798 (N_11798,N_6140,N_6709);
nor U11799 (N_11799,N_8520,N_7571);
or U11800 (N_11800,N_7532,N_8586);
and U11801 (N_11801,N_7970,N_7913);
xnor U11802 (N_11802,N_8959,N_7704);
or U11803 (N_11803,N_8495,N_8664);
and U11804 (N_11804,N_7863,N_8748);
nand U11805 (N_11805,N_6470,N_6856);
or U11806 (N_11806,N_6216,N_8890);
and U11807 (N_11807,N_7937,N_7963);
nor U11808 (N_11808,N_6497,N_7758);
nand U11809 (N_11809,N_7827,N_6127);
xnor U11810 (N_11810,N_8202,N_6436);
and U11811 (N_11811,N_7519,N_6321);
nand U11812 (N_11812,N_8268,N_8000);
and U11813 (N_11813,N_8928,N_8567);
xor U11814 (N_11814,N_7981,N_6064);
xor U11815 (N_11815,N_7388,N_6193);
nand U11816 (N_11816,N_7389,N_7779);
nor U11817 (N_11817,N_8770,N_7963);
nor U11818 (N_11818,N_7334,N_6330);
nor U11819 (N_11819,N_6196,N_7078);
xnor U11820 (N_11820,N_7740,N_8573);
or U11821 (N_11821,N_7048,N_7586);
or U11822 (N_11822,N_6830,N_7350);
and U11823 (N_11823,N_6637,N_6636);
or U11824 (N_11824,N_6563,N_7863);
nor U11825 (N_11825,N_8933,N_8623);
xnor U11826 (N_11826,N_8565,N_6920);
nor U11827 (N_11827,N_8164,N_8687);
and U11828 (N_11828,N_6305,N_6909);
xor U11829 (N_11829,N_7976,N_8241);
or U11830 (N_11830,N_7561,N_8334);
xnor U11831 (N_11831,N_6829,N_6308);
xor U11832 (N_11832,N_6525,N_6200);
nor U11833 (N_11833,N_7757,N_8066);
nor U11834 (N_11834,N_6921,N_7133);
and U11835 (N_11835,N_7186,N_7946);
nand U11836 (N_11836,N_6682,N_6360);
xor U11837 (N_11837,N_8263,N_6550);
nor U11838 (N_11838,N_8372,N_7314);
nor U11839 (N_11839,N_8900,N_8746);
xor U11840 (N_11840,N_6288,N_6380);
nor U11841 (N_11841,N_8966,N_7023);
or U11842 (N_11842,N_8099,N_7439);
xor U11843 (N_11843,N_6749,N_8628);
and U11844 (N_11844,N_7806,N_7713);
and U11845 (N_11845,N_7774,N_6775);
nor U11846 (N_11846,N_7915,N_6465);
xnor U11847 (N_11847,N_7840,N_8797);
nand U11848 (N_11848,N_6942,N_8829);
or U11849 (N_11849,N_7731,N_6532);
nor U11850 (N_11850,N_8763,N_6462);
or U11851 (N_11851,N_7683,N_8132);
or U11852 (N_11852,N_7069,N_8032);
xnor U11853 (N_11853,N_6852,N_8902);
nand U11854 (N_11854,N_7688,N_6211);
and U11855 (N_11855,N_8611,N_8844);
xor U11856 (N_11856,N_8115,N_7568);
nand U11857 (N_11857,N_6129,N_6939);
or U11858 (N_11858,N_6761,N_7214);
xor U11859 (N_11859,N_8829,N_6317);
nand U11860 (N_11860,N_6955,N_8062);
nand U11861 (N_11861,N_8113,N_8352);
nand U11862 (N_11862,N_6861,N_7570);
nor U11863 (N_11863,N_8906,N_6423);
nor U11864 (N_11864,N_7610,N_7029);
and U11865 (N_11865,N_6935,N_8184);
nand U11866 (N_11866,N_8566,N_8003);
or U11867 (N_11867,N_6371,N_7176);
nor U11868 (N_11868,N_7791,N_8202);
or U11869 (N_11869,N_8177,N_7345);
or U11870 (N_11870,N_6307,N_8137);
and U11871 (N_11871,N_7204,N_6577);
nor U11872 (N_11872,N_7458,N_7822);
nand U11873 (N_11873,N_8123,N_8493);
and U11874 (N_11874,N_7697,N_8609);
nor U11875 (N_11875,N_8538,N_7998);
and U11876 (N_11876,N_6305,N_8401);
and U11877 (N_11877,N_6858,N_7013);
nand U11878 (N_11878,N_6274,N_6677);
and U11879 (N_11879,N_8527,N_6465);
xor U11880 (N_11880,N_7323,N_8702);
nand U11881 (N_11881,N_6498,N_7836);
nand U11882 (N_11882,N_6088,N_7097);
and U11883 (N_11883,N_7891,N_6419);
xnor U11884 (N_11884,N_6879,N_8894);
or U11885 (N_11885,N_7068,N_6469);
or U11886 (N_11886,N_8897,N_7476);
nor U11887 (N_11887,N_6464,N_6300);
nor U11888 (N_11888,N_6565,N_6334);
nor U11889 (N_11889,N_8271,N_8008);
and U11890 (N_11890,N_6778,N_6339);
xnor U11891 (N_11891,N_6543,N_8482);
and U11892 (N_11892,N_7634,N_8578);
xor U11893 (N_11893,N_8814,N_8083);
and U11894 (N_11894,N_6911,N_8027);
xnor U11895 (N_11895,N_8628,N_8726);
nor U11896 (N_11896,N_8688,N_8100);
xor U11897 (N_11897,N_7512,N_6855);
nor U11898 (N_11898,N_8849,N_6717);
xnor U11899 (N_11899,N_7669,N_7236);
xor U11900 (N_11900,N_8044,N_7256);
or U11901 (N_11901,N_8075,N_8735);
and U11902 (N_11902,N_7509,N_8572);
nor U11903 (N_11903,N_7255,N_8598);
nand U11904 (N_11904,N_8351,N_8651);
nand U11905 (N_11905,N_6684,N_8027);
nor U11906 (N_11906,N_7682,N_7607);
and U11907 (N_11907,N_7958,N_7461);
and U11908 (N_11908,N_6929,N_7176);
nor U11909 (N_11909,N_7370,N_8468);
nor U11910 (N_11910,N_6048,N_8124);
and U11911 (N_11911,N_6980,N_7385);
xor U11912 (N_11912,N_8473,N_8307);
or U11913 (N_11913,N_6765,N_8930);
nor U11914 (N_11914,N_7687,N_6177);
and U11915 (N_11915,N_6770,N_7808);
nor U11916 (N_11916,N_6821,N_6622);
nor U11917 (N_11917,N_6774,N_8407);
or U11918 (N_11918,N_7481,N_6817);
nor U11919 (N_11919,N_8459,N_8865);
nor U11920 (N_11920,N_6811,N_6345);
or U11921 (N_11921,N_7290,N_7706);
and U11922 (N_11922,N_6375,N_8101);
and U11923 (N_11923,N_7245,N_7476);
nor U11924 (N_11924,N_7524,N_7283);
and U11925 (N_11925,N_7583,N_8447);
nor U11926 (N_11926,N_8167,N_8162);
nand U11927 (N_11927,N_8941,N_6383);
nand U11928 (N_11928,N_6694,N_8439);
xnor U11929 (N_11929,N_7507,N_8906);
nor U11930 (N_11930,N_7553,N_6413);
and U11931 (N_11931,N_6775,N_6965);
nand U11932 (N_11932,N_8194,N_7737);
or U11933 (N_11933,N_7407,N_6819);
nand U11934 (N_11934,N_6193,N_8734);
and U11935 (N_11935,N_7764,N_8002);
xor U11936 (N_11936,N_8347,N_7567);
and U11937 (N_11937,N_8586,N_6578);
xor U11938 (N_11938,N_6660,N_6564);
and U11939 (N_11939,N_8442,N_6656);
and U11940 (N_11940,N_6646,N_7790);
xor U11941 (N_11941,N_8294,N_8825);
or U11942 (N_11942,N_8009,N_7358);
nand U11943 (N_11943,N_8244,N_7316);
xnor U11944 (N_11944,N_6349,N_7051);
or U11945 (N_11945,N_6265,N_7406);
nand U11946 (N_11946,N_6485,N_8676);
or U11947 (N_11947,N_7466,N_8535);
xor U11948 (N_11948,N_6024,N_6053);
nor U11949 (N_11949,N_7671,N_7250);
xor U11950 (N_11950,N_8436,N_8863);
or U11951 (N_11951,N_7866,N_7856);
or U11952 (N_11952,N_7417,N_7721);
nor U11953 (N_11953,N_8474,N_6221);
nor U11954 (N_11954,N_6157,N_8532);
or U11955 (N_11955,N_6944,N_6216);
and U11956 (N_11956,N_7981,N_6810);
xnor U11957 (N_11957,N_7941,N_8988);
or U11958 (N_11958,N_6209,N_7412);
nor U11959 (N_11959,N_8192,N_8410);
xor U11960 (N_11960,N_8416,N_8641);
and U11961 (N_11961,N_6309,N_6366);
nand U11962 (N_11962,N_7279,N_8399);
xor U11963 (N_11963,N_6977,N_8476);
nand U11964 (N_11964,N_8736,N_8941);
nand U11965 (N_11965,N_8276,N_8985);
xnor U11966 (N_11966,N_7937,N_8393);
nand U11967 (N_11967,N_8514,N_7458);
and U11968 (N_11968,N_7803,N_8124);
or U11969 (N_11969,N_8126,N_8548);
nor U11970 (N_11970,N_7060,N_6245);
or U11971 (N_11971,N_7409,N_6943);
and U11972 (N_11972,N_6701,N_6468);
nor U11973 (N_11973,N_8181,N_7806);
and U11974 (N_11974,N_7213,N_8414);
or U11975 (N_11975,N_6531,N_6684);
or U11976 (N_11976,N_7568,N_6829);
or U11977 (N_11977,N_7036,N_8567);
nor U11978 (N_11978,N_6545,N_6508);
xnor U11979 (N_11979,N_7829,N_7915);
xor U11980 (N_11980,N_7612,N_8517);
or U11981 (N_11981,N_7073,N_6986);
nor U11982 (N_11982,N_6407,N_6172);
xnor U11983 (N_11983,N_6441,N_7510);
and U11984 (N_11984,N_7137,N_8370);
nand U11985 (N_11985,N_8250,N_8396);
nand U11986 (N_11986,N_6019,N_8437);
nand U11987 (N_11987,N_6825,N_8821);
nor U11988 (N_11988,N_8761,N_7159);
nor U11989 (N_11989,N_6314,N_6714);
xor U11990 (N_11990,N_8843,N_7490);
xor U11991 (N_11991,N_8640,N_7318);
xor U11992 (N_11992,N_8948,N_7674);
nand U11993 (N_11993,N_7706,N_7774);
nand U11994 (N_11994,N_6421,N_8257);
and U11995 (N_11995,N_8686,N_6576);
nor U11996 (N_11996,N_8093,N_7264);
and U11997 (N_11997,N_6959,N_7419);
nand U11998 (N_11998,N_6535,N_6419);
nor U11999 (N_11999,N_7733,N_7358);
xor U12000 (N_12000,N_11737,N_10368);
xor U12001 (N_12001,N_11402,N_11827);
nand U12002 (N_12002,N_10586,N_10094);
xnor U12003 (N_12003,N_9267,N_9412);
or U12004 (N_12004,N_9999,N_11619);
nor U12005 (N_12005,N_10893,N_10501);
or U12006 (N_12006,N_10865,N_10287);
nand U12007 (N_12007,N_9151,N_10769);
or U12008 (N_12008,N_11865,N_10332);
nor U12009 (N_12009,N_9059,N_10993);
and U12010 (N_12010,N_10905,N_11064);
nand U12011 (N_12011,N_9260,N_9673);
nor U12012 (N_12012,N_10782,N_9062);
nor U12013 (N_12013,N_9503,N_9996);
nand U12014 (N_12014,N_9731,N_10852);
or U12015 (N_12015,N_11475,N_9700);
or U12016 (N_12016,N_10972,N_11647);
or U12017 (N_12017,N_9941,N_11766);
and U12018 (N_12018,N_10876,N_9956);
or U12019 (N_12019,N_10262,N_9159);
nor U12020 (N_12020,N_9210,N_11129);
xnor U12021 (N_12021,N_9255,N_11528);
nand U12022 (N_12022,N_10346,N_9202);
or U12023 (N_12023,N_10323,N_10173);
and U12024 (N_12024,N_10574,N_11880);
nor U12025 (N_12025,N_11909,N_11868);
xnor U12026 (N_12026,N_11059,N_9680);
and U12027 (N_12027,N_10577,N_9106);
nor U12028 (N_12028,N_11840,N_11327);
and U12029 (N_12029,N_9172,N_11613);
nor U12030 (N_12030,N_10082,N_9737);
nand U12031 (N_12031,N_10440,N_9660);
or U12032 (N_12032,N_11347,N_11163);
or U12033 (N_12033,N_10302,N_9063);
nand U12034 (N_12034,N_9735,N_11893);
and U12035 (N_12035,N_9857,N_11323);
and U12036 (N_12036,N_11663,N_9577);
xnor U12037 (N_12037,N_11911,N_9839);
or U12038 (N_12038,N_9187,N_11841);
and U12039 (N_12039,N_11174,N_11157);
nand U12040 (N_12040,N_10264,N_10595);
or U12041 (N_12041,N_11539,N_10295);
and U12042 (N_12042,N_10142,N_9155);
nand U12043 (N_12043,N_9301,N_10539);
nand U12044 (N_12044,N_11043,N_10158);
and U12045 (N_12045,N_10992,N_9642);
xnor U12046 (N_12046,N_11046,N_11125);
or U12047 (N_12047,N_10961,N_10982);
nor U12048 (N_12048,N_9471,N_10715);
xnor U12049 (N_12049,N_10114,N_10910);
xor U12050 (N_12050,N_9604,N_10144);
nor U12051 (N_12051,N_11874,N_9959);
nand U12052 (N_12052,N_9726,N_11141);
or U12053 (N_12053,N_11436,N_11366);
nor U12054 (N_12054,N_9665,N_9909);
and U12055 (N_12055,N_10472,N_10103);
xnor U12056 (N_12056,N_9979,N_10596);
nor U12057 (N_12057,N_9937,N_9876);
xor U12058 (N_12058,N_9512,N_11600);
xor U12059 (N_12059,N_10848,N_11115);
or U12060 (N_12060,N_10898,N_11314);
nand U12061 (N_12061,N_9685,N_9966);
or U12062 (N_12062,N_11920,N_11712);
nor U12063 (N_12063,N_11305,N_9372);
nor U12064 (N_12064,N_9991,N_10329);
nor U12065 (N_12065,N_9182,N_9021);
nand U12066 (N_12066,N_11717,N_11992);
and U12067 (N_12067,N_10489,N_11710);
nor U12068 (N_12068,N_9717,N_11888);
xnor U12069 (N_12069,N_10348,N_9205);
and U12070 (N_12070,N_10223,N_10627);
and U12071 (N_12071,N_10716,N_9124);
nor U12072 (N_12072,N_9747,N_11975);
nor U12073 (N_12073,N_11932,N_11867);
xor U12074 (N_12074,N_9249,N_11568);
xor U12075 (N_12075,N_10112,N_10268);
and U12076 (N_12076,N_11665,N_9510);
nor U12077 (N_12077,N_9366,N_10860);
xor U12078 (N_12078,N_11906,N_9513);
and U12079 (N_12079,N_11324,N_10592);
and U12080 (N_12080,N_11689,N_11538);
xnor U12081 (N_12081,N_9156,N_10617);
or U12082 (N_12082,N_10850,N_10817);
xor U12083 (N_12083,N_11554,N_11441);
and U12084 (N_12084,N_9905,N_10591);
or U12085 (N_12085,N_10823,N_10754);
nor U12086 (N_12086,N_9396,N_9800);
nand U12087 (N_12087,N_9086,N_9201);
nand U12088 (N_12088,N_11261,N_9600);
xor U12089 (N_12089,N_9364,N_9653);
or U12090 (N_12090,N_11733,N_9145);
or U12091 (N_12091,N_9089,N_10006);
nand U12092 (N_12092,N_11682,N_10784);
and U12093 (N_12093,N_9031,N_11887);
or U12094 (N_12094,N_9575,N_10189);
or U12095 (N_12095,N_10026,N_11702);
and U12096 (N_12096,N_9824,N_9949);
nand U12097 (N_12097,N_10689,N_10713);
and U12098 (N_12098,N_11716,N_9040);
xnor U12099 (N_12099,N_11462,N_10662);
xnor U12100 (N_12100,N_10120,N_10476);
xnor U12101 (N_12101,N_10305,N_10808);
and U12102 (N_12102,N_11839,N_9128);
nand U12103 (N_12103,N_9178,N_9231);
and U12104 (N_12104,N_9034,N_10971);
and U12105 (N_12105,N_10202,N_11098);
xnor U12106 (N_12106,N_9872,N_10360);
nand U12107 (N_12107,N_11916,N_10718);
nand U12108 (N_12108,N_9409,N_10275);
or U12109 (N_12109,N_9995,N_9079);
nand U12110 (N_12110,N_9353,N_10045);
or U12111 (N_12111,N_11580,N_10109);
nor U12112 (N_12112,N_11671,N_11859);
nor U12113 (N_12113,N_11995,N_10683);
nor U12114 (N_12114,N_11773,N_10075);
or U12115 (N_12115,N_11862,N_9015);
nand U12116 (N_12116,N_10767,N_10251);
nand U12117 (N_12117,N_11805,N_11257);
nor U12118 (N_12118,N_10786,N_10989);
and U12119 (N_12119,N_9678,N_11564);
or U12120 (N_12120,N_11715,N_9545);
nor U12121 (N_12121,N_11382,N_10804);
or U12122 (N_12122,N_9216,N_9593);
and U12123 (N_12123,N_11645,N_9313);
and U12124 (N_12124,N_10956,N_10722);
nand U12125 (N_12125,N_10690,N_9413);
nand U12126 (N_12126,N_9757,N_9865);
and U12127 (N_12127,N_9729,N_9931);
nor U12128 (N_12128,N_10326,N_10755);
nor U12129 (N_12129,N_10681,N_9098);
xnor U12130 (N_12130,N_10863,N_9190);
nand U12131 (N_12131,N_10918,N_9227);
xnor U12132 (N_12132,N_11807,N_10152);
nand U12133 (N_12133,N_10735,N_9226);
xor U12134 (N_12134,N_9212,N_9771);
or U12135 (N_12135,N_10449,N_11511);
or U12136 (N_12136,N_9035,N_10661);
and U12137 (N_12137,N_9228,N_11616);
nand U12138 (N_12138,N_10724,N_10694);
nor U12139 (N_12139,N_10952,N_11017);
or U12140 (N_12140,N_11131,N_11998);
and U12141 (N_12141,N_9773,N_11668);
nand U12142 (N_12142,N_10900,N_9103);
nor U12143 (N_12143,N_10698,N_10549);
nand U12144 (N_12144,N_10631,N_11588);
nor U12145 (N_12145,N_11074,N_9386);
and U12146 (N_12146,N_9361,N_10373);
or U12147 (N_12147,N_11806,N_10381);
nand U12148 (N_12148,N_10225,N_9567);
nor U12149 (N_12149,N_9169,N_10564);
and U12150 (N_12150,N_10639,N_9494);
or U12151 (N_12151,N_11765,N_10397);
and U12152 (N_12152,N_10442,N_10580);
or U12153 (N_12153,N_10944,N_9809);
xor U12154 (N_12154,N_11927,N_9390);
and U12155 (N_12155,N_11545,N_11727);
xnor U12156 (N_12156,N_9197,N_9463);
and U12157 (N_12157,N_9204,N_11006);
nor U12158 (N_12158,N_9767,N_9799);
or U12159 (N_12159,N_10936,N_10292);
nand U12160 (N_12160,N_10590,N_9990);
and U12161 (N_12161,N_11656,N_9482);
xnor U12162 (N_12162,N_9423,N_9874);
or U12163 (N_12163,N_9293,N_10392);
nor U12164 (N_12164,N_9427,N_10967);
and U12165 (N_12165,N_10078,N_10391);
or U12166 (N_12166,N_10061,N_9886);
nor U12167 (N_12167,N_10677,N_9417);
nand U12168 (N_12168,N_11453,N_10987);
or U12169 (N_12169,N_11465,N_10912);
and U12170 (N_12170,N_10390,N_10315);
and U12171 (N_12171,N_11073,N_9768);
and U12172 (N_12172,N_9582,N_11186);
and U12173 (N_12173,N_11735,N_9849);
or U12174 (N_12174,N_11358,N_11696);
and U12175 (N_12175,N_9324,N_11637);
and U12176 (N_12176,N_9272,N_9614);
nor U12177 (N_12177,N_9153,N_9064);
or U12178 (N_12178,N_10766,N_11774);
xor U12179 (N_12179,N_11572,N_10975);
xor U12180 (N_12180,N_10077,N_11375);
xor U12181 (N_12181,N_10899,N_10645);
or U12182 (N_12182,N_11171,N_10543);
and U12183 (N_12183,N_10603,N_10573);
nand U12184 (N_12184,N_9317,N_11329);
or U12185 (N_12185,N_9971,N_10976);
nor U12186 (N_12186,N_9517,N_9418);
xor U12187 (N_12187,N_11255,N_9043);
and U12188 (N_12188,N_11630,N_10664);
xor U12189 (N_12189,N_10949,N_9362);
nand U12190 (N_12190,N_11144,N_9442);
and U12191 (N_12191,N_10629,N_10818);
or U12192 (N_12192,N_9134,N_11274);
nand U12193 (N_12193,N_9536,N_10678);
and U12194 (N_12194,N_9623,N_10479);
or U12195 (N_12195,N_9848,N_9568);
nor U12196 (N_12196,N_9077,N_11151);
or U12197 (N_12197,N_11183,N_9573);
nand U12198 (N_12198,N_10088,N_10730);
nor U12199 (N_12199,N_10347,N_9852);
nor U12200 (N_12200,N_10418,N_10836);
and U12201 (N_12201,N_9903,N_10528);
and U12202 (N_12202,N_11557,N_10463);
or U12203 (N_12203,N_9123,N_9783);
nand U12204 (N_12204,N_9777,N_11933);
nand U12205 (N_12205,N_11275,N_9681);
nand U12206 (N_12206,N_10998,N_11757);
or U12207 (N_12207,N_10255,N_11793);
xnor U12208 (N_12208,N_10535,N_9053);
and U12209 (N_12209,N_10191,N_9118);
or U12210 (N_12210,N_9348,N_11348);
or U12211 (N_12211,N_11177,N_10922);
and U12212 (N_12212,N_9320,N_11626);
nor U12213 (N_12213,N_10113,N_10569);
nand U12214 (N_12214,N_11563,N_9472);
or U12215 (N_12215,N_11896,N_10762);
and U12216 (N_12216,N_10515,N_9920);
nand U12217 (N_12217,N_10869,N_10481);
nor U12218 (N_12218,N_10529,N_11155);
or U12219 (N_12219,N_9061,N_10499);
nand U12220 (N_12220,N_10085,N_9405);
nand U12221 (N_12221,N_11924,N_10599);
nand U12222 (N_12222,N_9758,N_9621);
nor U12223 (N_12223,N_9547,N_9752);
or U12224 (N_12224,N_9631,N_10155);
or U12225 (N_12225,N_10247,N_9051);
nor U12226 (N_12226,N_9778,N_9085);
nand U12227 (N_12227,N_11188,N_11761);
or U12228 (N_12228,N_9612,N_9071);
and U12229 (N_12229,N_9273,N_11479);
nand U12230 (N_12230,N_10525,N_9625);
or U12231 (N_12231,N_10376,N_11411);
or U12232 (N_12232,N_10246,N_10212);
nand U12233 (N_12233,N_10425,N_9684);
or U12234 (N_12234,N_9559,N_9963);
or U12235 (N_12235,N_10055,N_10053);
and U12236 (N_12236,N_11272,N_10278);
nor U12237 (N_12237,N_10636,N_9613);
nor U12238 (N_12238,N_11683,N_9521);
nand U12239 (N_12239,N_10140,N_10932);
or U12240 (N_12240,N_11142,N_11824);
nand U12241 (N_12241,N_11214,N_11590);
nand U12242 (N_12242,N_10706,N_10995);
and U12243 (N_12243,N_11136,N_9993);
nor U12244 (N_12244,N_9323,N_10897);
and U12245 (N_12245,N_11178,N_11181);
or U12246 (N_12246,N_9470,N_10427);
nand U12247 (N_12247,N_10907,N_11662);
or U12248 (N_12248,N_10163,N_11099);
nor U12249 (N_12249,N_9637,N_10190);
xor U12250 (N_12250,N_11037,N_9105);
nand U12251 (N_12251,N_11768,N_10024);
and U12252 (N_12252,N_10740,N_11578);
or U12253 (N_12253,N_11670,N_10195);
xnor U12254 (N_12254,N_11969,N_11176);
and U12255 (N_12255,N_11800,N_10530);
nand U12256 (N_12256,N_9798,N_11980);
nand U12257 (N_12257,N_9304,N_9232);
nor U12258 (N_12258,N_10902,N_11147);
xor U12259 (N_12259,N_11105,N_10619);
and U12260 (N_12260,N_9734,N_10999);
nand U12261 (N_12261,N_9251,N_10692);
and U12262 (N_12262,N_9942,N_9358);
or U12263 (N_12263,N_9017,N_11293);
and U12264 (N_12264,N_9452,N_11250);
nand U12265 (N_12265,N_11981,N_11222);
or U12266 (N_12266,N_10412,N_11675);
nor U12267 (N_12267,N_9893,N_10606);
and U12268 (N_12268,N_10948,N_10483);
or U12269 (N_12269,N_9380,N_9630);
xnor U12270 (N_12270,N_10203,N_11842);
or U12271 (N_12271,N_9627,N_10273);
nor U12272 (N_12272,N_9391,N_10791);
or U12273 (N_12273,N_9654,N_10903);
xor U12274 (N_12274,N_10333,N_11522);
nor U12275 (N_12275,N_11116,N_11446);
nor U12276 (N_12276,N_10915,N_11084);
xor U12277 (N_12277,N_10675,N_9538);
nor U12278 (N_12278,N_10423,N_10623);
xnor U12279 (N_12279,N_10695,N_10162);
nand U12280 (N_12280,N_11565,N_10759);
and U12281 (N_12281,N_10977,N_11336);
nor U12282 (N_12282,N_9708,N_11127);
or U12283 (N_12283,N_10316,N_9009);
xnor U12284 (N_12284,N_9264,N_11211);
or U12285 (N_12285,N_9050,N_11756);
nor U12286 (N_12286,N_10238,N_9461);
or U12287 (N_12287,N_9336,N_10039);
nand U12288 (N_12288,N_9531,N_9307);
nor U12289 (N_12289,N_9634,N_11118);
nor U12290 (N_12290,N_9200,N_10584);
nor U12291 (N_12291,N_11233,N_11412);
xnor U12292 (N_12292,N_11159,N_9352);
nand U12293 (N_12293,N_10781,N_10194);
and U12294 (N_12294,N_9180,N_9347);
nand U12295 (N_12295,N_9940,N_9042);
and U12296 (N_12296,N_10057,N_10856);
nor U12297 (N_12297,N_9422,N_11625);
nand U12298 (N_12298,N_10285,N_11471);
or U12299 (N_12299,N_11573,N_9952);
nand U12300 (N_12300,N_9793,N_10761);
or U12301 (N_12301,N_10044,N_9355);
xnor U12302 (N_12302,N_9132,N_11655);
or U12303 (N_12303,N_9481,N_10745);
nor U12304 (N_12304,N_9867,N_9663);
and U12305 (N_12305,N_9860,N_9584);
or U12306 (N_12306,N_11295,N_11648);
xnor U12307 (N_12307,N_11667,N_10701);
nor U12308 (N_12308,N_10974,N_10269);
or U12309 (N_12309,N_11100,N_9449);
xnor U12310 (N_12310,N_9898,N_11638);
nand U12311 (N_12311,N_10452,N_9306);
and U12312 (N_12312,N_9933,N_10254);
xnor U12313 (N_12313,N_9075,N_11569);
xor U12314 (N_12314,N_10557,N_11200);
nor U12315 (N_12315,N_11015,N_10825);
or U12316 (N_12316,N_10705,N_10841);
nor U12317 (N_12317,N_10032,N_9770);
nor U12318 (N_12318,N_10291,N_11606);
xnor U12319 (N_12319,N_9214,N_10231);
nor U12320 (N_12320,N_11967,N_10598);
and U12321 (N_12321,N_11432,N_9511);
nand U12322 (N_12322,N_11890,N_11399);
nor U12323 (N_12323,N_11044,N_11700);
and U12324 (N_12324,N_11621,N_11310);
or U12325 (N_12325,N_9961,N_9211);
nor U12326 (N_12326,N_10802,N_9149);
and U12327 (N_12327,N_11033,N_10406);
xnor U12328 (N_12328,N_9083,N_9540);
xnor U12329 (N_12329,N_10179,N_11820);
and U12330 (N_12330,N_9420,N_10828);
or U12331 (N_12331,N_11858,N_11658);
nand U12332 (N_12332,N_11540,N_11623);
and U12333 (N_12333,N_11734,N_11405);
nand U12334 (N_12334,N_11597,N_9407);
or U12335 (N_12335,N_11929,N_10983);
nand U12336 (N_12336,N_11976,N_9802);
nand U12337 (N_12337,N_10408,N_11930);
xor U12338 (N_12338,N_11102,N_11705);
nor U12339 (N_12339,N_9791,N_9912);
nor U12340 (N_12340,N_9426,N_11373);
nor U12341 (N_12341,N_10774,N_10493);
xor U12342 (N_12342,N_10356,N_10845);
nor U12343 (N_12343,N_10838,N_9645);
xnor U12344 (N_12344,N_9498,N_11473);
and U12345 (N_12345,N_10613,N_9274);
xnor U12346 (N_12346,N_11622,N_11204);
and U12347 (N_12347,N_11113,N_11771);
or U12348 (N_12348,N_10351,N_11352);
xnor U12349 (N_12349,N_9842,N_9827);
nor U12350 (N_12350,N_9240,N_10959);
nor U12351 (N_12351,N_10719,N_9938);
and U12352 (N_12352,N_11869,N_11928);
xor U12353 (N_12353,N_10296,N_9992);
and U12354 (N_12354,N_10357,N_11326);
or U12355 (N_12355,N_9004,N_9025);
and U12356 (N_12356,N_10785,N_10879);
and U12357 (N_12357,N_10693,N_10159);
nor U12358 (N_12358,N_11226,N_11476);
and U12359 (N_12359,N_10647,N_9090);
nor U12360 (N_12360,N_9732,N_11739);
and U12361 (N_12361,N_11139,N_10330);
xnor U12362 (N_12362,N_10510,N_11835);
xor U12363 (N_12363,N_11090,N_11227);
xor U12364 (N_12364,N_11986,N_9981);
nand U12365 (N_12365,N_10321,N_9252);
nor U12366 (N_12366,N_10393,N_9987);
or U12367 (N_12367,N_11532,N_11282);
xor U12368 (N_12368,N_9616,N_9601);
xor U12369 (N_12369,N_9344,N_11503);
and U12370 (N_12370,N_10562,N_11050);
xor U12371 (N_12371,N_10986,N_10455);
or U12372 (N_12372,N_11523,N_9280);
xor U12373 (N_12373,N_9977,N_9398);
and U12374 (N_12374,N_10753,N_11703);
nand U12375 (N_12375,N_11831,N_9581);
nand U12376 (N_12376,N_9177,N_10249);
nor U12377 (N_12377,N_10468,N_10593);
and U12378 (N_12378,N_11685,N_9147);
or U12379 (N_12379,N_10395,N_9488);
and U12380 (N_12380,N_10643,N_11978);
xor U12381 (N_12381,N_9333,N_11393);
and U12382 (N_12382,N_9588,N_11923);
nand U12383 (N_12383,N_9707,N_10301);
nor U12384 (N_12384,N_9733,N_11194);
or U12385 (N_12385,N_10712,N_9710);
and U12386 (N_12386,N_10178,N_9455);
nand U12387 (N_12387,N_11158,N_10386);
nand U12388 (N_12388,N_11866,N_11649);
nand U12389 (N_12389,N_9864,N_9594);
nor U12390 (N_12390,N_10950,N_11094);
xnor U12391 (N_12391,N_11801,N_9702);
nor U12392 (N_12392,N_11520,N_10670);
nor U12393 (N_12393,N_10906,N_11075);
nand U12394 (N_12394,N_10511,N_10589);
or U12395 (N_12395,N_11506,N_10908);
nand U12396 (N_12396,N_9254,N_11197);
and U12397 (N_12397,N_10957,N_11848);
and U12398 (N_12398,N_10064,N_10339);
and U12399 (N_12399,N_9524,N_11755);
xnor U12400 (N_12400,N_11990,N_10306);
nand U12401 (N_12401,N_10985,N_9571);
xnor U12402 (N_12402,N_9976,N_11660);
or U12403 (N_12403,N_9853,N_9057);
or U12404 (N_12404,N_9535,N_11857);
or U12405 (N_12405,N_10022,N_9024);
and U12406 (N_12406,N_10122,N_9003);
and U12407 (N_12407,N_10877,N_9823);
nand U12408 (N_12408,N_9465,N_10086);
or U12409 (N_12409,N_10208,N_11316);
or U12410 (N_12410,N_10235,N_9497);
and U12411 (N_12411,N_9000,N_11633);
xor U12412 (N_12412,N_9919,N_9329);
and U12413 (N_12413,N_9882,N_11172);
nor U12414 (N_12414,N_9556,N_10851);
nor U12415 (N_12415,N_10136,N_10568);
and U12416 (N_12416,N_9657,N_9739);
nor U12417 (N_12417,N_9428,N_10980);
xor U12418 (N_12418,N_9074,N_10146);
and U12419 (N_12419,N_9485,N_9394);
nand U12420 (N_12420,N_9238,N_11886);
nor U12421 (N_12421,N_11794,N_11844);
and U12422 (N_12422,N_9763,N_10538);
nand U12423 (N_12423,N_10696,N_9826);
xor U12424 (N_12424,N_11301,N_11979);
or U12425 (N_12425,N_11229,N_10074);
nor U12426 (N_12426,N_11270,N_11950);
xor U12427 (N_12427,N_9669,N_11235);
and U12428 (N_12428,N_11065,N_9878);
nand U12429 (N_12429,N_11669,N_9095);
nor U12430 (N_12430,N_11121,N_9456);
xnor U12431 (N_12431,N_11130,N_10419);
or U12432 (N_12432,N_9819,N_9048);
nor U12433 (N_12433,N_9244,N_9469);
nor U12434 (N_12434,N_9220,N_9140);
nand U12435 (N_12435,N_9821,N_9659);
xor U12436 (N_12436,N_11317,N_10261);
nand U12437 (N_12437,N_9300,N_9199);
and U12438 (N_12438,N_9125,N_11586);
nor U12439 (N_12439,N_9828,N_11832);
or U12440 (N_12440,N_11057,N_10720);
nor U12441 (N_12441,N_9687,N_11516);
nand U12442 (N_12442,N_11816,N_10253);
nand U12443 (N_12443,N_9871,N_9960);
nor U12444 (N_12444,N_11718,N_10855);
xor U12445 (N_12445,N_11743,N_9805);
nor U12446 (N_12446,N_10741,N_9602);
xor U12447 (N_12447,N_11818,N_10783);
and U12448 (N_12448,N_10625,N_11559);
nand U12449 (N_12449,N_10551,N_11991);
nand U12450 (N_12450,N_11398,N_9879);
nand U12451 (N_12451,N_11052,N_10721);
xor U12452 (N_12452,N_10129,N_11325);
xnor U12453 (N_12453,N_11591,N_10250);
nor U12454 (N_12454,N_10215,N_11104);
xor U12455 (N_12455,N_9213,N_10801);
and U12456 (N_12456,N_10388,N_11965);
xor U12457 (N_12457,N_10115,N_10007);
or U12458 (N_12458,N_11397,N_10990);
or U12459 (N_12459,N_9332,N_11396);
nand U12460 (N_12460,N_9989,N_10496);
and U12461 (N_12461,N_11984,N_10375);
and U12462 (N_12462,N_11322,N_10224);
or U12463 (N_12463,N_11461,N_11946);
nand U12464 (N_12464,N_10181,N_9387);
nand U12465 (N_12465,N_11456,N_11515);
and U12466 (N_12466,N_10776,N_9781);
nor U12467 (N_12467,N_9855,N_11791);
xor U12468 (N_12468,N_10954,N_9544);
or U12469 (N_12469,N_9723,N_9229);
or U12470 (N_12470,N_10338,N_9672);
xnor U12471 (N_12471,N_9667,N_9974);
and U12472 (N_12472,N_9837,N_9914);
or U12473 (N_12473,N_11983,N_9222);
xnor U12474 (N_12474,N_10450,N_11741);
xnor U12475 (N_12475,N_9859,N_9640);
and U12476 (N_12476,N_11497,N_10209);
and U12477 (N_12477,N_11241,N_9351);
and U12478 (N_12478,N_10916,N_10938);
or U12479 (N_12479,N_9972,N_10787);
nand U12480 (N_12480,N_11072,N_9755);
and U12481 (N_12481,N_11740,N_11627);
or U12482 (N_12482,N_10369,N_9840);
nor U12483 (N_12483,N_10708,N_11910);
or U12484 (N_12484,N_11302,N_11234);
xor U12485 (N_12485,N_11750,N_10884);
or U12486 (N_12486,N_10151,N_10428);
and U12487 (N_12487,N_9910,N_10260);
and U12488 (N_12488,N_9143,N_9373);
nor U12489 (N_12489,N_10409,N_10204);
and U12490 (N_12490,N_11931,N_11736);
or U12491 (N_12491,N_11319,N_9792);
nor U12492 (N_12492,N_10892,N_11510);
xnor U12493 (N_12493,N_10978,N_9985);
xnor U12494 (N_12494,N_11882,N_10180);
nor U12495 (N_12495,N_11639,N_11146);
xor U12496 (N_12496,N_11720,N_11369);
nand U12497 (N_12497,N_9858,N_10649);
nor U12498 (N_12498,N_10150,N_11679);
nor U12499 (N_12499,N_9760,N_10778);
nand U12500 (N_12500,N_11042,N_9656);
nand U12501 (N_12501,N_11289,N_9108);
nor U12502 (N_12502,N_9862,N_11894);
xnor U12503 (N_12503,N_9766,N_9850);
xor U12504 (N_12504,N_11789,N_10717);
nand U12505 (N_12505,N_11145,N_11798);
nor U12506 (N_12506,N_10005,N_10207);
and U12507 (N_12507,N_10199,N_10644);
xnor U12508 (N_12508,N_9701,N_10895);
nor U12509 (N_12509,N_10600,N_10399);
nand U12510 (N_12510,N_10447,N_9779);
or U12511 (N_12511,N_10458,N_9450);
or U12512 (N_12512,N_9424,N_10313);
and U12513 (N_12513,N_9318,N_9002);
and U12514 (N_12514,N_9276,N_11243);
or U12515 (N_12515,N_10751,N_9266);
xnor U12516 (N_12516,N_9484,N_10826);
nor U12517 (N_12517,N_9501,N_10737);
or U12518 (N_12518,N_9887,N_9745);
or U12519 (N_12519,N_11708,N_9709);
nand U12520 (N_12520,N_10821,N_11269);
xor U12521 (N_12521,N_9546,N_11232);
xnor U12522 (N_12522,N_9107,N_9343);
and U12523 (N_12523,N_9945,N_9237);
xnor U12524 (N_12524,N_9808,N_10228);
or U12525 (N_12525,N_9796,N_10023);
nand U12526 (N_12526,N_11300,N_9946);
nor U12527 (N_12527,N_9198,N_11407);
xor U12528 (N_12528,N_9831,N_10789);
and U12529 (N_12529,N_11362,N_11277);
xnor U12530 (N_12530,N_10844,N_9291);
or U12531 (N_12531,N_11230,N_9294);
xor U12532 (N_12532,N_9221,N_11484);
xor U12533 (N_12533,N_11408,N_11541);
nand U12534 (N_12534,N_9360,N_11926);
and U12535 (N_12535,N_9924,N_11507);
or U12536 (N_12536,N_10991,N_9639);
or U12537 (N_12537,N_9636,N_9176);
xnor U12538 (N_12538,N_10051,N_9529);
nor U12539 (N_12539,N_11355,N_10832);
or U12540 (N_12540,N_10544,N_10834);
nand U12541 (N_12541,N_11977,N_11889);
and U12542 (N_12542,N_11068,N_10536);
nor U12543 (N_12543,N_9045,N_11742);
or U12544 (N_12544,N_11337,N_11416);
nor U12545 (N_12545,N_11562,N_10211);
and U12546 (N_12546,N_11120,N_11086);
or U12547 (N_12547,N_9620,N_9346);
or U12548 (N_12548,N_9493,N_9587);
and U12549 (N_12549,N_10940,N_9440);
and U12550 (N_12550,N_9316,N_11137);
and U12551 (N_12551,N_10665,N_10581);
and U12552 (N_12552,N_10342,N_11304);
and U12553 (N_12553,N_11466,N_11834);
nand U12554 (N_12554,N_10018,N_11615);
or U12555 (N_12555,N_9219,N_10669);
and U12556 (N_12556,N_10049,N_9950);
xor U12557 (N_12557,N_9988,N_11108);
or U12558 (N_12558,N_11721,N_11029);
nor U12559 (N_12559,N_11031,N_10046);
nand U12560 (N_12560,N_11431,N_11095);
xor U12561 (N_12561,N_11486,N_9629);
and U12562 (N_12562,N_10547,N_9926);
nor U12563 (N_12563,N_9868,N_10572);
nand U12564 (N_12564,N_11917,N_10668);
nand U12565 (N_12565,N_9589,N_10080);
and U12566 (N_12566,N_11331,N_11542);
nand U12567 (N_12567,N_11501,N_9965);
nor U12568 (N_12568,N_9643,N_11674);
nand U12569 (N_12569,N_10579,N_11256);
nor U12570 (N_12570,N_10484,N_11328);
xor U12571 (N_12571,N_11769,N_10337);
or U12572 (N_12572,N_10359,N_10362);
or U12573 (N_12573,N_11262,N_9292);
nand U12574 (N_12574,N_10065,N_11829);
or U12575 (N_12575,N_10859,N_11001);
or U12576 (N_12576,N_11895,N_10711);
or U12577 (N_12577,N_11109,N_9081);
nand U12578 (N_12578,N_10355,N_10526);
nand U12579 (N_12579,N_11394,N_11608);
xnor U12580 (N_12580,N_11213,N_11164);
xor U12581 (N_12581,N_9036,N_9875);
or U12582 (N_12582,N_11598,N_9619);
nand U12583 (N_12583,N_11023,N_11258);
and U12584 (N_12584,N_11560,N_11852);
nand U12585 (N_12585,N_10100,N_10641);
and U12586 (N_12586,N_11838,N_9207);
nor U12587 (N_12587,N_10312,N_10098);
or U12588 (N_12588,N_11821,N_9110);
or U12589 (N_12589,N_10340,N_9148);
nand U12590 (N_12590,N_10833,N_9179);
nor U12591 (N_12591,N_11185,N_9113);
nand U12592 (N_12592,N_11504,N_9130);
nand U12593 (N_12593,N_10175,N_10125);
or U12594 (N_12594,N_10758,N_9167);
and U12595 (N_12595,N_9955,N_9998);
nor U12596 (N_12596,N_9431,N_11081);
nand U12597 (N_12597,N_11706,N_10068);
nand U12598 (N_12598,N_10035,N_9916);
nor U12599 (N_12599,N_11400,N_11076);
and U12600 (N_12600,N_9776,N_9296);
and U12601 (N_12601,N_11751,N_9127);
or U12602 (N_12602,N_11083,N_9135);
nor U12603 (N_12603,N_11103,N_9445);
and U12604 (N_12604,N_10276,N_11653);
xnor U12605 (N_12605,N_9927,N_9270);
and U12606 (N_12606,N_10843,N_11051);
nor U12607 (N_12607,N_11779,N_9530);
xor U12608 (N_12608,N_9901,N_9066);
or U12609 (N_12609,N_9632,N_11066);
and U12610 (N_12610,N_9129,N_10854);
and U12611 (N_12611,N_10929,N_9023);
xor U12612 (N_12612,N_9434,N_9235);
nor U12613 (N_12613,N_9012,N_10233);
or U12614 (N_12614,N_10660,N_9561);
xnor U12615 (N_12615,N_11711,N_11069);
nand U12616 (N_12616,N_9939,N_11485);
or U12617 (N_12617,N_9978,N_9131);
or U12618 (N_12618,N_9789,N_10968);
nand U12619 (N_12619,N_10614,N_9185);
xor U12620 (N_12620,N_10079,N_9038);
xor U12621 (N_12621,N_9406,N_9873);
nand U12622 (N_12622,N_9441,N_9746);
or U12623 (N_12623,N_10646,N_9404);
nor U12624 (N_12624,N_11960,N_11018);
nor U12625 (N_12625,N_9438,N_11643);
nor U12626 (N_12626,N_9818,N_11659);
nand U12627 (N_12627,N_10028,N_11438);
and U12628 (N_12628,N_10582,N_9402);
nor U12629 (N_12629,N_9263,N_11254);
and U12630 (N_12630,N_9285,N_9122);
or U12631 (N_12631,N_9870,N_10748);
or U12632 (N_12632,N_11149,N_10226);
xor U12633 (N_12633,N_11437,N_10763);
nor U12634 (N_12634,N_10453,N_11907);
nor U12635 (N_12635,N_10608,N_9502);
xor U12636 (N_12636,N_9562,N_11225);
nand U12637 (N_12637,N_11561,N_10001);
nand U12638 (N_12638,N_10004,N_9047);
and U12639 (N_12639,N_9753,N_11748);
nand U12640 (N_12640,N_10130,N_9383);
xor U12641 (N_12641,N_9807,N_11448);
nand U12642 (N_12642,N_10868,N_11672);
and U12643 (N_12643,N_9617,N_10605);
and U12644 (N_12644,N_10220,N_9415);
nor U12645 (N_12645,N_10182,N_9607);
or U12646 (N_12646,N_11551,N_10488);
nor U12647 (N_12647,N_10744,N_10890);
nor U12648 (N_12648,N_9881,N_11693);
and U12649 (N_12649,N_10042,N_9121);
nor U12650 (N_12650,N_10597,N_11731);
or U12651 (N_12651,N_9730,N_11007);
xnor U12652 (N_12652,N_10700,N_10602);
nor U12653 (N_12653,N_10421,N_11518);
and U12654 (N_12654,N_9311,N_11321);
xor U12655 (N_12655,N_9586,N_9369);
nand U12656 (N_12656,N_10941,N_10506);
nor U12657 (N_12657,N_10813,N_9835);
xnor U12658 (N_12658,N_10256,N_9574);
nand U12659 (N_12659,N_10410,N_11078);
and U12660 (N_12660,N_9934,N_11219);
and U12661 (N_12661,N_11878,N_9191);
xor U12662 (N_12662,N_11491,N_11935);
nor U12663 (N_12663,N_9774,N_11087);
nand U12664 (N_12664,N_11698,N_10609);
xnor U12665 (N_12665,N_9894,N_11134);
xnor U12666 (N_12666,N_10087,N_10354);
nand U12667 (N_12667,N_10658,N_10019);
nand U12668 (N_12668,N_11404,N_10198);
xnor U12669 (N_12669,N_9499,N_11810);
and U12670 (N_12670,N_10298,N_11215);
nor U12671 (N_12671,N_11775,N_11596);
or U12672 (N_12672,N_10252,N_11611);
or U12673 (N_12673,N_9688,N_10084);
nand U12674 (N_12674,N_11126,N_11414);
nor U12675 (N_12675,N_11420,N_11860);
and U12676 (N_12676,N_11447,N_9670);
and U12677 (N_12677,N_11368,N_10997);
and U12678 (N_12678,N_10523,N_11624);
or U12679 (N_12679,N_9305,N_10655);
nand U12680 (N_12680,N_10415,N_11025);
or U12681 (N_12681,N_11024,N_11828);
or U12682 (N_12682,N_9432,N_10628);
nand U12683 (N_12683,N_9345,N_11217);
nand U12684 (N_12684,N_9416,N_9705);
or U12685 (N_12685,N_10352,N_10725);
xnor U12686 (N_12686,N_9056,N_11035);
xnor U12687 (N_12687,N_9350,N_11216);
xnor U12688 (N_12688,N_9044,N_9608);
or U12689 (N_12689,N_9328,N_9271);
nor U12690 (N_12690,N_9635,N_9157);
xnor U12691 (N_12691,N_9314,N_9338);
or U12692 (N_12692,N_9339,N_11850);
or U12693 (N_12693,N_10265,N_9741);
and U12694 (N_12694,N_10404,N_11440);
or U12695 (N_12695,N_10994,N_9217);
nor U12696 (N_12696,N_10576,N_9473);
nand U12697 (N_12697,N_10402,N_11056);
and U12698 (N_12698,N_10030,N_11745);
nand U12699 (N_12699,N_10772,N_9929);
and U12700 (N_12700,N_11196,N_11026);
and U12701 (N_12701,N_11753,N_10206);
and U12702 (N_12702,N_10575,N_9738);
nand U12703 (N_12703,N_9389,N_11601);
nor U12704 (N_12704,N_10875,N_10861);
or U12705 (N_12705,N_11989,N_10107);
nor U12706 (N_12706,N_9014,N_9393);
xor U12707 (N_12707,N_9060,N_9166);
and U12708 (N_12708,N_9379,N_10881);
xnor U12709 (N_12709,N_9772,N_11166);
or U12710 (N_12710,N_10002,N_9321);
and U12711 (N_12711,N_11160,N_9967);
xnor U12712 (N_12712,N_11180,N_10210);
and U12713 (N_12713,N_11458,N_11020);
nand U12714 (N_12714,N_11856,N_9288);
or U12715 (N_12715,N_10437,N_10872);
xor U12716 (N_12716,N_9506,N_9368);
or U12717 (N_12717,N_10299,N_9563);
xnor U12718 (N_12718,N_10743,N_11237);
and U12719 (N_12719,N_9644,N_11439);
and U12720 (N_12720,N_10793,N_9651);
or U12721 (N_12721,N_11193,N_10334);
xnor U12722 (N_12722,N_10413,N_11354);
or U12723 (N_12723,N_11847,N_9786);
nand U12724 (N_12724,N_11592,N_11964);
nand U12725 (N_12725,N_10322,N_9088);
xor U12726 (N_12726,N_11636,N_10840);
or U12727 (N_12727,N_9419,N_10732);
nor U12728 (N_12728,N_11195,N_11101);
nor U12729 (N_12729,N_9740,N_11320);
or U12730 (N_12730,N_11027,N_9489);
or U12731 (N_12731,N_10697,N_10736);
and U12732 (N_12732,N_11032,N_9676);
and U12733 (N_12733,N_11008,N_11093);
or U12734 (N_12734,N_10684,N_11218);
xnor U12735 (N_12735,N_10411,N_9692);
and U12736 (N_12736,N_11266,N_11021);
or U12737 (N_12737,N_10556,N_9683);
nand U12738 (N_12738,N_10667,N_9281);
and U12739 (N_12739,N_9532,N_11822);
nor U12740 (N_12740,N_11372,N_10156);
nand U12741 (N_12741,N_11381,N_11455);
nor U12742 (N_12742,N_11948,N_11921);
and U12743 (N_12743,N_10911,N_10092);
or U12744 (N_12744,N_10749,N_9436);
nor U12745 (N_12745,N_10517,N_9628);
or U12746 (N_12746,N_10883,N_10277);
or U12747 (N_12747,N_10962,N_9505);
nor U12748 (N_12748,N_9504,N_11357);
xnor U12749 (N_12749,N_9475,N_10282);
nor U12750 (N_12750,N_11283,N_9541);
nand U12751 (N_12751,N_9164,N_10090);
xor U12752 (N_12752,N_9500,N_11576);
nand U12753 (N_12753,N_11954,N_9720);
nor U12754 (N_12754,N_9527,N_10227);
xnor U12755 (N_12755,N_11535,N_11553);
nand U12756 (N_12756,N_9958,N_10361);
nor U12757 (N_12757,N_10127,N_11962);
nand U12758 (N_12758,N_11005,N_11334);
and U12759 (N_12759,N_10846,N_9225);
or U12760 (N_12760,N_11190,N_10234);
nor U12761 (N_12761,N_10979,N_11434);
and U12762 (N_12762,N_11536,N_11688);
nand U12763 (N_12763,N_11409,N_10171);
xor U12764 (N_12764,N_10200,N_11786);
xor U12765 (N_12765,N_9566,N_11014);
nand U12766 (N_12766,N_11985,N_11422);
xnor U12767 (N_12767,N_11220,N_9282);
nor U12768 (N_12768,N_9453,N_10842);
or U12769 (N_12769,N_11268,N_9877);
and U12770 (N_12770,N_11898,N_10490);
or U12771 (N_12771,N_10060,N_11498);
xor U12772 (N_12772,N_11879,N_9005);
nand U12773 (N_12773,N_11517,N_11642);
xnor U12774 (N_12774,N_10102,N_11199);
or U12775 (N_12775,N_9880,N_9605);
and U12776 (N_12776,N_10524,N_9444);
xnor U12777 (N_12777,N_10503,N_11747);
nand U12778 (N_12778,N_9312,N_11430);
xor U12779 (N_12779,N_9904,N_10015);
or U12780 (N_12780,N_9165,N_9611);
or U12781 (N_12781,N_9215,N_10803);
xnor U12782 (N_12782,N_11264,N_10814);
nand U12783 (N_12783,N_9954,N_11079);
and U12784 (N_12784,N_11876,N_9365);
nand U12785 (N_12785,N_10010,N_9648);
or U12786 (N_12786,N_10792,N_11036);
and U12787 (N_12787,N_11961,N_11558);
and U12788 (N_12788,N_10430,N_11169);
and U12789 (N_12789,N_11817,N_10118);
and U12790 (N_12790,N_11963,N_11521);
or U12791 (N_12791,N_10003,N_10733);
and U12792 (N_12792,N_10300,N_11333);
and U12793 (N_12793,N_10746,N_10110);
or U12794 (N_12794,N_11132,N_10070);
and U12795 (N_12795,N_10314,N_9930);
nand U12796 (N_12796,N_9811,N_9248);
nand U12797 (N_12797,N_11604,N_10663);
and U12798 (N_12798,N_9697,N_9649);
and U12799 (N_12799,N_11492,N_9534);
xor U12800 (N_12800,N_10245,N_9957);
xor U12801 (N_12801,N_9902,N_9928);
or U12802 (N_12802,N_11210,N_10981);
xnor U12803 (N_12803,N_10350,N_9487);
xnor U12804 (N_12804,N_11010,N_11644);
or U12805 (N_12805,N_10960,N_11085);
xnor U12806 (N_12806,N_11206,N_9655);
xnor U12807 (N_12807,N_9539,N_9078);
and U12808 (N_12808,N_10920,N_11280);
and U12809 (N_12809,N_10521,N_11468);
and U12810 (N_12810,N_10487,N_9794);
nor U12811 (N_12811,N_10477,N_10494);
and U12812 (N_12812,N_9013,N_11278);
and U12813 (N_12813,N_10467,N_10239);
nor U12814 (N_12814,N_11242,N_10567);
and U12815 (N_12815,N_11004,N_11605);
nor U12816 (N_12816,N_11854,N_11170);
and U12817 (N_12817,N_10676,N_9973);
xor U12818 (N_12818,N_10289,N_9287);
and U12819 (N_12819,N_11238,N_9250);
nor U12820 (N_12820,N_11594,N_11285);
and U12821 (N_12821,N_10063,N_10089);
nand U12822 (N_12822,N_10327,N_10111);
or U12823 (N_12823,N_11488,N_10888);
nand U12824 (N_12824,N_11949,N_9111);
and U12825 (N_12825,N_10638,N_11449);
and U12826 (N_12826,N_10345,N_11915);
xor U12827 (N_12827,N_10218,N_11514);
nand U12828 (N_12828,N_9550,N_9410);
nand U12829 (N_12829,N_10138,N_11651);
nand U12830 (N_12830,N_10824,N_11942);
and U12831 (N_12831,N_9762,N_9883);
and U12832 (N_12832,N_11875,N_11150);
nor U12833 (N_12833,N_9782,N_11749);
and U12834 (N_12834,N_10723,N_9247);
and U12835 (N_12835,N_11661,N_10324);
nand U12836 (N_12836,N_11067,N_11038);
nor U12837 (N_12837,N_9552,N_9724);
and U12838 (N_12838,N_10270,N_11341);
nor U12839 (N_12839,N_10734,N_10095);
or U12840 (N_12840,N_11602,N_9467);
or U12841 (N_12841,N_11386,N_9962);
and U12842 (N_12842,N_9261,N_10474);
and U12843 (N_12843,N_10942,N_9764);
xor U12844 (N_12844,N_11135,N_9528);
nor U12845 (N_12845,N_11088,N_11919);
and U12846 (N_12846,N_9714,N_11138);
and U12847 (N_12847,N_11054,N_11003);
and U12848 (N_12848,N_10482,N_11451);
and U12849 (N_12849,N_10072,N_11389);
and U12850 (N_12850,N_10141,N_9579);
nand U12851 (N_12851,N_10027,N_10779);
xor U12852 (N_12852,N_9039,N_11764);
nor U12853 (N_12853,N_10885,N_11982);
nor U12854 (N_12854,N_9006,N_11599);
nand U12855 (N_12855,N_10012,N_9020);
nor U12856 (N_12856,N_10559,N_11843);
or U12857 (N_12857,N_10344,N_10214);
or U12858 (N_12858,N_9233,N_11759);
nor U12859 (N_12859,N_9668,N_9633);
nor U12860 (N_12860,N_9780,N_11092);
xor U12861 (N_12861,N_11244,N_9788);
xnor U12862 (N_12862,N_9994,N_11531);
nand U12863 (N_12863,N_10849,N_9268);
or U12864 (N_12864,N_10933,N_11934);
xnor U12865 (N_12865,N_10222,N_11585);
and U12866 (N_12866,N_9549,N_10176);
or U12867 (N_12867,N_11426,N_11678);
or U12868 (N_12868,N_10671,N_10632);
nor U12869 (N_12869,N_10328,N_10013);
xor U12870 (N_12870,N_9516,N_11478);
nand U12871 (N_12871,N_10796,N_10016);
or U12872 (N_12872,N_11053,N_11509);
nor U12873 (N_12873,N_9814,N_10552);
and U12874 (N_12874,N_11784,N_10157);
or U12875 (N_12875,N_9403,N_11676);
nor U12876 (N_12876,N_9496,N_11684);
nand U12877 (N_12877,N_11881,N_9283);
or U12878 (N_12878,N_10471,N_9486);
nor U12879 (N_12879,N_11951,N_11719);
nor U12880 (N_12880,N_9411,N_9430);
nor U12881 (N_12881,N_11294,N_9377);
and U12882 (N_12882,N_11427,N_11459);
nor U12883 (N_12883,N_10166,N_9895);
xnor U12884 (N_12884,N_9082,N_10454);
nand U12885 (N_12885,N_9367,N_9970);
and U12886 (N_12886,N_11813,N_9188);
nand U12887 (N_12887,N_10308,N_9560);
xnor U12888 (N_12888,N_10963,N_11738);
nor U12889 (N_12889,N_10691,N_10765);
xnor U12890 (N_12890,N_11251,N_11286);
nand U12891 (N_12891,N_9716,N_10290);
xnor U12892 (N_12892,N_9029,N_10637);
nand U12893 (N_12893,N_10434,N_11785);
nor U12894 (N_12894,N_11344,N_11987);
or U12895 (N_12895,N_10857,N_9290);
and U12896 (N_12896,N_9869,N_9162);
nand U12897 (N_12897,N_11425,N_9018);
xor U12898 (N_12898,N_9069,N_10913);
and U12899 (N_12899,N_10624,N_11128);
xor U12900 (N_12900,N_9184,N_10816);
nor U12901 (N_12901,N_10618,N_11959);
nor U12902 (N_12902,N_11746,N_10853);
xor U12903 (N_12903,N_9299,N_10121);
xor U12904 (N_12904,N_11855,N_9196);
nor U12905 (N_12905,N_11744,N_9829);
and U12906 (N_12906,N_10657,N_10076);
or U12907 (N_12907,N_10570,N_9590);
or U12908 (N_12908,N_10901,N_9342);
nand U12909 (N_12909,N_10835,N_10945);
nand U12910 (N_12910,N_11571,N_9181);
and U12911 (N_12911,N_11346,N_10988);
and U12912 (N_12912,N_11460,N_11885);
or U12913 (N_12913,N_10831,N_10545);
xnor U12914 (N_12914,N_11641,N_11383);
or U12915 (N_12915,N_9693,N_10699);
and U12916 (N_12916,N_10429,N_9690);
nand U12917 (N_12917,N_9548,N_10436);
nor U12918 (N_12918,N_9054,N_10919);
nand U12919 (N_12919,N_10183,N_10043);
xor U12920 (N_12920,N_9703,N_10040);
nor U12921 (N_12921,N_11593,N_10924);
and U12922 (N_12922,N_10871,N_11508);
and U12923 (N_12923,N_11287,N_10674);
or U12924 (N_12924,N_10738,N_11767);
xor U12925 (N_12925,N_9866,N_10052);
and U12926 (N_12926,N_10866,N_10174);
nand U12927 (N_12927,N_10507,N_10473);
nand U12928 (N_12928,N_11260,N_10777);
and U12929 (N_12929,N_11359,N_10727);
and U12930 (N_12930,N_9696,N_11699);
xnor U12931 (N_12931,N_9727,N_10143);
xor U12932 (N_12932,N_11363,N_9698);
or U12933 (N_12933,N_11096,N_11011);
and U12934 (N_12934,N_11002,N_11192);
xnor U12935 (N_12935,N_9790,N_9278);
nor U12936 (N_12936,N_10927,N_10304);
nand U12937 (N_12937,N_9357,N_10101);
nand U12938 (N_12938,N_11292,N_10147);
nor U12939 (N_12939,N_9921,N_9326);
nand U12940 (N_12940,N_9603,N_9349);
xor U12941 (N_12941,N_9421,N_10435);
xor U12942 (N_12942,N_11477,N_11245);
xnor U12943 (N_12943,N_11444,N_11529);
nand U12944 (N_12944,N_11570,N_10274);
nor U12945 (N_12945,N_11533,N_10492);
nand U12946 (N_12946,N_11823,N_11587);
xor U12947 (N_12947,N_9951,N_11947);
nand U12948 (N_12948,N_11861,N_10904);
or U12949 (N_12949,N_10648,N_11758);
nand U12950 (N_12950,N_10422,N_11958);
xor U12951 (N_12951,N_10672,N_9885);
nand U12952 (N_12952,N_10405,N_10566);
nand U12953 (N_12953,N_11423,N_10154);
and U12954 (N_12954,N_9569,N_9785);
nor U12955 (N_12955,N_9152,N_9997);
and U12956 (N_12956,N_11953,N_11870);
xnor U12957 (N_12957,N_10236,N_9514);
nand U12958 (N_12958,N_10242,N_11082);
and U12959 (N_12959,N_9892,N_9836);
nand U12960 (N_12960,N_11306,N_10232);
nand U12961 (N_12961,N_9119,N_11513);
nor U12962 (N_12962,N_10622,N_11296);
nor U12963 (N_12963,N_9209,N_9065);
nand U12964 (N_12964,N_9136,N_10820);
nor U12965 (N_12965,N_10955,N_9126);
and U12966 (N_12966,N_9968,N_9376);
nand U12967 (N_12967,N_9388,N_11997);
nand U12968 (N_12968,N_9666,N_9297);
or U12969 (N_12969,N_9055,N_10651);
or U12970 (N_12970,N_11349,N_11902);
nor U12971 (N_12971,N_9750,N_11311);
xor U12972 (N_12972,N_11377,N_11481);
and U12973 (N_12973,N_11332,N_9459);
xor U12974 (N_12974,N_11550,N_11781);
or U12975 (N_12975,N_10168,N_10378);
or U12976 (N_12976,N_10491,N_10534);
xnor U12977 (N_12977,N_9116,N_11628);
xor U12978 (N_12978,N_10134,N_10266);
and U12979 (N_12979,N_10128,N_9142);
xnor U12980 (N_12980,N_11620,N_10284);
nand U12981 (N_12981,N_9975,N_9558);
xor U12982 (N_12982,N_9585,N_10213);
nand U12983 (N_12983,N_11039,N_10800);
and U12984 (N_12984,N_9058,N_11966);
or U12985 (N_12985,N_10807,N_10372);
nor U12986 (N_12986,N_10319,N_11161);
and U12987 (N_12987,N_10219,N_10230);
or U12988 (N_12988,N_9918,N_10502);
or U12989 (N_12989,N_9032,N_10459);
or U12990 (N_12990,N_10259,N_9030);
nor U12991 (N_12991,N_11897,N_11041);
or U12992 (N_12992,N_9718,N_11077);
xnor U12993 (N_12993,N_11340,N_9592);
or U12994 (N_12994,N_9515,N_10640);
nand U12995 (N_12995,N_9622,N_11607);
nor U12996 (N_12996,N_10439,N_9446);
nand U12997 (N_12997,N_11208,N_11391);
nand U12998 (N_12998,N_11945,N_11070);
xor U12999 (N_12999,N_10073,N_11577);
nor U13000 (N_13000,N_10830,N_10750);
nor U13001 (N_13001,N_11016,N_11970);
nor U13002 (N_13002,N_9448,N_9097);
and U13003 (N_13003,N_10331,N_9443);
and U13004 (N_13004,N_9067,N_11635);
nor U13005 (N_13005,N_10578,N_9922);
or U13006 (N_13006,N_11308,N_9555);
nor U13007 (N_13007,N_9102,N_10293);
nand U13008 (N_13008,N_9094,N_9269);
nor U13009 (N_13009,N_9374,N_11153);
and U13010 (N_13010,N_10343,N_9392);
or U13011 (N_13011,N_10520,N_9141);
nand U13012 (N_13012,N_11061,N_11048);
xnor U13013 (N_13013,N_10161,N_9239);
nand U13014 (N_13014,N_10533,N_11640);
nor U13015 (N_13015,N_10460,N_11175);
xor U13016 (N_13016,N_10426,N_9457);
and U13017 (N_13017,N_11239,N_11315);
xor U13018 (N_13018,N_11788,N_11677);
or U13019 (N_13019,N_10553,N_9341);
nand U13020 (N_13020,N_9661,N_10185);
xnor U13021 (N_13021,N_10363,N_9378);
and U13022 (N_13022,N_9277,N_11891);
or U13023 (N_13023,N_10119,N_9597);
nor U13024 (N_13024,N_10135,N_9509);
nand U13025 (N_13025,N_10656,N_9598);
nand U13026 (N_13026,N_11298,N_11376);
nand U13027 (N_13027,N_11307,N_11106);
nor U13028 (N_13028,N_11168,N_9923);
xnor U13029 (N_13029,N_11695,N_10106);
and U13030 (N_13030,N_11546,N_10752);
nor U13031 (N_13031,N_10041,N_10882);
nand U13032 (N_13032,N_9906,N_11249);
or U13033 (N_13033,N_11450,N_11162);
or U13034 (N_13034,N_10267,N_9425);
nor U13035 (N_13035,N_10280,N_9932);
nand U13036 (N_13036,N_9578,N_10620);
or U13037 (N_13037,N_11803,N_9286);
nor U13038 (N_13038,N_10193,N_10133);
xnor U13039 (N_13039,N_10367,N_10031);
nand U13040 (N_13040,N_9715,N_11783);
or U13041 (N_13041,N_10448,N_11124);
nor U13042 (N_13042,N_10811,N_10237);
or U13043 (N_13043,N_9451,N_10635);
and U13044 (N_13044,N_10137,N_9624);
xnor U13045 (N_13045,N_11034,N_10531);
xor U13046 (N_13046,N_9236,N_10069);
nor U13047 (N_13047,N_9615,N_11714);
or U13048 (N_13048,N_9289,N_11378);
nand U13049 (N_13049,N_9695,N_9986);
nor U13050 (N_13050,N_9834,N_9076);
and U13051 (N_13051,N_11697,N_9144);
nor U13052 (N_13052,N_9911,N_11156);
nor U13053 (N_13053,N_9170,N_9899);
nand U13054 (N_13054,N_10780,N_11707);
nand U13055 (N_13055,N_11614,N_11548);
and U13056 (N_13056,N_11259,N_11811);
nor U13057 (N_13057,N_9679,N_11291);
and U13058 (N_13058,N_10398,N_11500);
xor U13059 (N_13059,N_10020,N_11330);
nand U13060 (N_13060,N_11752,N_11846);
xor U13061 (N_13061,N_11631,N_11730);
nor U13062 (N_13062,N_10205,N_9576);
nor U13063 (N_13063,N_9033,N_9856);
and U13064 (N_13064,N_10958,N_9087);
nand U13065 (N_13065,N_10432,N_11883);
nand U13066 (N_13066,N_9175,N_9253);
or U13067 (N_13067,N_10126,N_10921);
and U13068 (N_13068,N_9719,N_10887);
nand U13069 (N_13069,N_10894,N_9399);
nor U13070 (N_13070,N_9694,N_9889);
or U13071 (N_13071,N_10951,N_9308);
and U13072 (N_13072,N_9230,N_11071);
nand U13073 (N_13073,N_10417,N_11988);
or U13074 (N_13074,N_11552,N_11792);
xnor U13075 (N_13075,N_10548,N_11148);
nor U13076 (N_13076,N_10048,N_10047);
xor U13077 (N_13077,N_10058,N_11173);
nor U13078 (N_13078,N_9662,N_10462);
xnor U13079 (N_13079,N_11974,N_11912);
nor U13080 (N_13080,N_10288,N_9284);
nor U13081 (N_13081,N_10475,N_11830);
xnor U13082 (N_13082,N_10806,N_9580);
xnor U13083 (N_13083,N_10066,N_9984);
nor U13084 (N_13084,N_9599,N_11467);
nand U13085 (N_13085,N_10403,N_10400);
and U13086 (N_13086,N_9298,N_11288);
or U13087 (N_13087,N_9722,N_11815);
xnor U13088 (N_13088,N_9256,N_9553);
xnor U13089 (N_13089,N_9706,N_9721);
xnor U13090 (N_13090,N_10703,N_9072);
nand U13091 (N_13091,N_10445,N_10160);
xnor U13092 (N_13092,N_9223,N_9775);
nand U13093 (N_13093,N_11973,N_10819);
nand U13094 (N_13094,N_11826,N_9743);
nand U13095 (N_13095,N_9658,N_11335);
nand U13096 (N_13096,N_9749,N_10747);
or U13097 (N_13097,N_9109,N_9322);
or U13098 (N_13098,N_9841,N_10729);
or U13099 (N_13099,N_9897,N_9769);
or U13100 (N_13100,N_9310,N_10424);
or U13101 (N_13101,N_11123,N_11778);
nor U13102 (N_13102,N_10034,N_10380);
nor U13103 (N_13103,N_11547,N_10926);
or U13104 (N_13104,N_9689,N_9218);
or U13105 (N_13105,N_11309,N_11941);
xor U13106 (N_13106,N_9896,N_11231);
xnor U13107 (N_13107,N_9099,N_11212);
and U13108 (N_13108,N_11457,N_11603);
nand U13109 (N_13109,N_10809,N_10704);
or U13110 (N_13110,N_11884,N_10946);
nor U13111 (N_13111,N_10188,N_9832);
or U13112 (N_13112,N_9595,N_11454);
nor U13113 (N_13113,N_11360,N_11284);
nor U13114 (N_13114,N_11940,N_10874);
nand U13115 (N_13115,N_9331,N_11493);
xnor U13116 (N_13116,N_10630,N_10389);
nor U13117 (N_13117,N_9359,N_10497);
xnor U13118 (N_13118,N_11971,N_10486);
and U13119 (N_13119,N_11119,N_10033);
nor U13120 (N_13120,N_10197,N_11780);
and U13121 (N_13121,N_11167,N_9262);
and U13122 (N_13122,N_10770,N_11385);
nand U13123 (N_13123,N_11845,N_11502);
nand U13124 (N_13124,N_10056,N_11392);
or U13125 (N_13125,N_10607,N_9751);
nor U13126 (N_13126,N_10541,N_10594);
xor U13127 (N_13127,N_11111,N_10177);
nor U13128 (N_13128,N_9258,N_9699);
xnor U13129 (N_13129,N_11191,N_11387);
nor U13130 (N_13130,N_10878,N_11913);
or U13131 (N_13131,N_11804,N_11728);
xnor U13132 (N_13132,N_9947,N_10414);
xnor U13133 (N_13133,N_11202,N_9028);
xor U13134 (N_13134,N_9279,N_10371);
nor U13135 (N_13135,N_11080,N_9682);
nand U13136 (N_13136,N_10923,N_11595);
or U13137 (N_13137,N_10810,N_10666);
or U13138 (N_13138,N_10480,N_9460);
nand U13139 (N_13139,N_11418,N_11772);
xor U13140 (N_13140,N_9725,N_11140);
nand U13141 (N_13141,N_11634,N_11583);
nor U13142 (N_13142,N_10478,N_11030);
nor U13143 (N_13143,N_11534,N_10540);
nor U13144 (N_13144,N_9638,N_10798);
nor U13145 (N_13145,N_10864,N_9572);
nand U13146 (N_13146,N_11401,N_11726);
or U13147 (N_13147,N_11526,N_11790);
or U13148 (N_13148,N_11410,N_9565);
xor U13149 (N_13149,N_10466,N_10588);
or U13150 (N_13150,N_9171,N_11692);
and U13151 (N_13151,N_10099,N_11819);
xnor U13152 (N_13152,N_10546,N_9523);
nor U13153 (N_13153,N_11421,N_11617);
and U13154 (N_13154,N_11729,N_9816);
nand U13155 (N_13155,N_9761,N_11351);
nor U13156 (N_13156,N_9803,N_10431);
or U13157 (N_13157,N_10132,N_9011);
or U13158 (N_13158,N_10303,N_11110);
nor U13159 (N_13159,N_9820,N_9812);
or U13160 (N_13160,N_10017,N_10297);
nand U13161 (N_13161,N_10062,N_10317);
nor U13162 (N_13162,N_9983,N_9334);
nand U13163 (N_13163,N_11223,N_10728);
nor U13164 (N_13164,N_10310,N_11312);
xor U13165 (N_13165,N_11247,N_9943);
nor U13166 (N_13166,N_10984,N_10272);
nor U13167 (N_13167,N_9728,N_10123);
or U13168 (N_13168,N_11936,N_10091);
nand U13169 (N_13169,N_11303,N_9371);
and U13170 (N_13170,N_9520,N_11443);
xor U13171 (N_13171,N_10286,N_11379);
nor U13172 (N_13172,N_11487,N_9195);
nor U13173 (N_13173,N_9908,N_11925);
nor U13174 (N_13174,N_11994,N_9327);
xnor U13175 (N_13175,N_11776,N_11922);
nor U13176 (N_13176,N_10318,N_9464);
or U13177 (N_13177,N_11000,N_9257);
or U13178 (N_13178,N_11107,N_9795);
xor U13179 (N_13179,N_10021,N_11666);
and U13180 (N_13180,N_11429,N_11445);
nor U13181 (N_13181,N_11664,N_11361);
or U13182 (N_13182,N_9052,N_11143);
xor U13183 (N_13183,N_11474,N_11544);
xnor U13184 (N_13184,N_9093,N_11575);
and U13185 (N_13185,N_11089,N_9117);
and U13186 (N_13186,N_11763,N_9007);
nor U13187 (N_13187,N_10108,N_9797);
nor U13188 (N_13188,N_11632,N_9609);
nand U13189 (N_13189,N_10930,N_9491);
nand U13190 (N_13190,N_11777,N_10516);
or U13191 (N_13191,N_10827,N_11567);
xor U13192 (N_13192,N_10500,N_10294);
or U13193 (N_13193,N_10366,N_11796);
nand U13194 (N_13194,N_10495,N_9104);
nor U13195 (N_13195,N_10438,N_9026);
nor U13196 (N_13196,N_11184,N_11395);
xor U13197 (N_13197,N_10527,N_11713);
nor U13198 (N_13198,N_10935,N_9194);
nand U13199 (N_13199,N_9542,N_10867);
nor U13200 (N_13200,N_10358,N_9163);
nand U13201 (N_13201,N_9096,N_9861);
or U13202 (N_13202,N_11833,N_10407);
xnor U13203 (N_13203,N_9138,N_10554);
and U13204 (N_13204,N_9935,N_11864);
or U13205 (N_13205,N_11537,N_9526);
and U13206 (N_13206,N_10394,N_11345);
and U13207 (N_13207,N_11704,N_11364);
xor U13208 (N_13208,N_10457,N_9375);
and U13209 (N_13209,N_10686,N_10917);
nand U13210 (N_13210,N_10837,N_10610);
or U13211 (N_13211,N_10271,N_11472);
or U13212 (N_13212,N_9234,N_11681);
and U13213 (N_13213,N_11470,N_11589);
nor U13214 (N_13214,N_11901,N_9037);
nor U13215 (N_13215,N_9907,N_11944);
or U13216 (N_13216,N_10008,N_10243);
nor U13217 (N_13217,N_9677,N_10653);
xnor U13218 (N_13218,N_10059,N_11228);
and U13219 (N_13219,N_9408,N_11452);
nand U13220 (N_13220,N_9070,N_10889);
or U13221 (N_13221,N_9830,N_9474);
or U13222 (N_13222,N_11836,N_11221);
nor U13223 (N_13223,N_11956,N_11629);
nand U13224 (N_13224,N_10505,N_9046);
nor U13225 (N_13225,N_10731,N_9787);
and U13226 (N_13226,N_9641,N_11795);
or U13227 (N_13227,N_9208,N_11353);
and U13228 (N_13228,N_9647,N_10096);
nand U13229 (N_13229,N_9784,N_9477);
or U13230 (N_13230,N_11770,N_11428);
and U13231 (N_13231,N_9468,N_11028);
and U13232 (N_13232,N_10611,N_11290);
nand U13233 (N_13233,N_11837,N_9295);
nor U13234 (N_13234,N_11045,N_11782);
or U13235 (N_13235,N_11968,N_10522);
and U13236 (N_13236,N_9846,N_9822);
nor U13237 (N_13237,N_10470,N_9596);
nand U13238 (N_13238,N_10221,N_11374);
nor U13239 (N_13239,N_11701,N_10870);
xor U13240 (N_13240,N_11612,N_11646);
nor U13241 (N_13241,N_9458,N_9010);
or U13242 (N_13242,N_9150,N_9711);
nand U13243 (N_13243,N_9041,N_11318);
and U13244 (N_13244,N_11236,N_11342);
xor U13245 (N_13245,N_10465,N_10011);
xnor U13246 (N_13246,N_10931,N_9183);
nor U13247 (N_13247,N_11365,N_11581);
or U13248 (N_13248,N_10587,N_10139);
nand U13249 (N_13249,N_11265,N_9671);
nand U13250 (N_13250,N_11797,N_10886);
or U13251 (N_13251,N_11725,N_11505);
and U13252 (N_13252,N_10947,N_9847);
xor U13253 (N_13253,N_11122,N_9462);
and U13254 (N_13254,N_10335,N_10642);
nor U13255 (N_13255,N_11117,N_10970);
and U13256 (N_13256,N_9370,N_9900);
or U13257 (N_13257,N_9888,N_11957);
and U13258 (N_13258,N_11343,N_10508);
nor U13259 (N_13259,N_11182,N_10558);
and U13260 (N_13260,N_11722,N_11009);
nand U13261 (N_13261,N_10167,N_10518);
xor U13262 (N_13262,N_11905,N_9936);
xnor U13263 (N_13263,N_9833,N_11338);
nand U13264 (N_13264,N_11694,N_9092);
and U13265 (N_13265,N_10311,N_9851);
xnor U13266 (N_13266,N_10896,N_10192);
xor U13267 (N_13267,N_10229,N_9964);
nor U13268 (N_13268,N_9114,N_11566);
nor U13269 (N_13269,N_9168,N_10281);
nor U13270 (N_13270,N_10307,N_9810);
nor U13271 (N_13271,N_9275,N_9354);
and U13272 (N_13272,N_10196,N_9192);
nor U13273 (N_13273,N_9309,N_10469);
nor U13274 (N_13274,N_9193,N_11419);
or U13275 (N_13275,N_10621,N_10964);
xor U13276 (N_13276,N_9435,N_10679);
and U13277 (N_13277,N_10773,N_11209);
and U13278 (N_13278,N_10244,N_10757);
nand U13279 (N_13279,N_11022,N_11279);
nor U13280 (N_13280,N_10000,N_10839);
nand U13281 (N_13281,N_10050,N_11490);
nand U13282 (N_13282,N_10186,N_10514);
nand U13283 (N_13283,N_9027,N_11047);
nand U13284 (N_13284,N_9381,N_11825);
nand U13285 (N_13285,N_11496,N_9161);
xor U13286 (N_13286,N_10377,N_10365);
or U13287 (N_13287,N_9825,N_11812);
nand U13288 (N_13288,N_11680,N_9704);
xor U13289 (N_13289,N_9845,N_11556);
or U13290 (N_13290,N_10320,N_10153);
nor U13291 (N_13291,N_9817,N_10714);
nor U13292 (N_13292,N_10217,N_10036);
nand U13293 (N_13293,N_10148,N_10054);
nand U13294 (N_13294,N_10847,N_10105);
nand U13295 (N_13295,N_10943,N_10537);
nor U13296 (N_13296,N_11762,N_11914);
nor U13297 (N_13297,N_9507,N_9154);
and U13298 (N_13298,N_10498,N_10688);
nand U13299 (N_13299,N_9691,N_9564);
or U13300 (N_13300,N_10604,N_9982);
and U13301 (N_13301,N_11205,N_11271);
xnor U13302 (N_13302,N_11062,N_10726);
or U13303 (N_13303,N_9174,N_10925);
nor U13304 (N_13304,N_10756,N_9884);
and U13305 (N_13305,N_9675,N_10532);
xnor U13306 (N_13306,N_9913,N_10025);
nand U13307 (N_13307,N_11152,N_11339);
xnor U13308 (N_13308,N_11367,N_11787);
xor U13309 (N_13309,N_10788,N_9016);
or U13310 (N_13310,N_11494,N_9337);
nor U13311 (N_13311,N_10973,N_10353);
and U13312 (N_13312,N_11019,N_9890);
nor U13313 (N_13313,N_11527,N_11267);
or U13314 (N_13314,N_10485,N_9139);
nor U13315 (N_13315,N_11246,N_10873);
nand U13316 (N_13316,N_11060,N_11900);
nand U13317 (N_13317,N_10165,N_9490);
nand U13318 (N_13318,N_9815,N_10464);
xor U13319 (N_13319,N_11525,N_11207);
nand U13320 (N_13320,N_11424,N_10258);
nor U13321 (N_13321,N_9115,N_9173);
nor U13322 (N_13322,N_9980,N_10097);
and U13323 (N_13323,N_11657,N_10083);
or U13324 (N_13324,N_10822,N_9019);
or U13325 (N_13325,N_9242,N_9806);
nor U13326 (N_13326,N_9022,N_10382);
xnor U13327 (N_13327,N_11584,N_10349);
or U13328 (N_13328,N_11165,N_11918);
nand U13329 (N_13329,N_10169,N_11224);
xnor U13330 (N_13330,N_10009,N_10702);
xnor U13331 (N_13331,N_11904,N_9137);
or U13332 (N_13332,N_9112,N_11380);
nand U13333 (N_13333,N_9969,N_10965);
and U13334 (N_13334,N_9519,N_9742);
nand U13335 (N_13335,N_9925,N_10093);
nand U13336 (N_13336,N_9385,N_10634);
nand U13337 (N_13337,N_10038,N_11760);
or U13338 (N_13338,N_11938,N_10709);
nor U13339 (N_13339,N_11483,N_9765);
and U13340 (N_13340,N_11097,N_10561);
nor U13341 (N_13341,N_10612,N_9606);
and U13342 (N_13342,N_9340,N_10616);
and U13343 (N_13343,N_10862,N_9537);
nand U13344 (N_13344,N_9429,N_11198);
nor U13345 (N_13345,N_10037,N_11417);
and U13346 (N_13346,N_10650,N_11201);
nor U13347 (N_13347,N_11415,N_10673);
xor U13348 (N_13348,N_10815,N_9508);
and U13349 (N_13349,N_9049,N_9543);
and U13350 (N_13350,N_9008,N_11114);
and U13351 (N_13351,N_10739,N_10797);
nand U13352 (N_13352,N_9356,N_9756);
or U13353 (N_13353,N_10014,N_9259);
nor U13354 (N_13354,N_10441,N_9759);
nand U13355 (N_13355,N_10812,N_10659);
and U13356 (N_13356,N_11530,N_9146);
nand U13357 (N_13357,N_10170,N_10937);
nand U13358 (N_13358,N_9686,N_10504);
nand U13359 (N_13359,N_9748,N_10257);
nand U13360 (N_13360,N_9382,N_9953);
and U13361 (N_13361,N_10768,N_10550);
and U13362 (N_13362,N_11091,N_11574);
or U13363 (N_13363,N_11802,N_9712);
or U13364 (N_13364,N_9335,N_11390);
xnor U13365 (N_13365,N_9447,N_11686);
or U13366 (N_13366,N_11276,N_10184);
or U13367 (N_13367,N_10081,N_9551);
or U13368 (N_13368,N_10370,N_11799);
and U13369 (N_13369,N_10934,N_11482);
nand U13370 (N_13370,N_9674,N_9480);
or U13371 (N_13371,N_9101,N_9570);
or U13372 (N_13372,N_10283,N_10654);
and U13373 (N_13373,N_10341,N_9891);
nand U13374 (N_13374,N_9915,N_11313);
or U13375 (N_13375,N_9133,N_10914);
and U13376 (N_13376,N_10996,N_10149);
or U13377 (N_13377,N_9395,N_10401);
xnor U13378 (N_13378,N_11724,N_9080);
nand U13379 (N_13379,N_10216,N_9206);
xor U13380 (N_13380,N_9091,N_10117);
nand U13381 (N_13381,N_10794,N_11996);
or U13382 (N_13382,N_9224,N_11495);
or U13383 (N_13383,N_10633,N_9713);
and U13384 (N_13384,N_9948,N_11609);
nor U13385 (N_13385,N_9158,N_10240);
and U13386 (N_13386,N_10443,N_9917);
xor U13387 (N_13387,N_11903,N_9303);
xnor U13388 (N_13388,N_9610,N_10565);
nand U13389 (N_13389,N_10775,N_10446);
nor U13390 (N_13390,N_10953,N_9437);
or U13391 (N_13391,N_9330,N_11939);
or U13392 (N_13392,N_11555,N_9476);
or U13393 (N_13393,N_9838,N_11908);
nand U13394 (N_13394,N_9533,N_11723);
nor U13395 (N_13395,N_11524,N_10685);
xnor U13396 (N_13396,N_9483,N_10416);
nand U13397 (N_13397,N_9454,N_9001);
or U13398 (N_13398,N_11937,N_11610);
and U13399 (N_13399,N_10451,N_9844);
and U13400 (N_13400,N_9120,N_11442);
or U13401 (N_13401,N_10104,N_10387);
xor U13402 (N_13402,N_9466,N_11463);
or U13403 (N_13403,N_9944,N_10164);
nor U13404 (N_13404,N_9843,N_9100);
nand U13405 (N_13405,N_11480,N_10145);
xnor U13406 (N_13406,N_9246,N_11248);
xor U13407 (N_13407,N_11582,N_10374);
nand U13408 (N_13408,N_11403,N_9384);
nor U13409 (N_13409,N_10384,N_10601);
and U13410 (N_13410,N_11654,N_9325);
or U13411 (N_13411,N_9414,N_9189);
nor U13412 (N_13412,N_10707,N_10891);
nor U13413 (N_13413,N_10858,N_9245);
nor U13414 (N_13414,N_10742,N_10909);
and U13415 (N_13415,N_9068,N_9652);
xor U13416 (N_13416,N_11413,N_11112);
and U13417 (N_13417,N_9315,N_11709);
or U13418 (N_13418,N_11013,N_11808);
xnor U13419 (N_13419,N_10513,N_11252);
xor U13420 (N_13420,N_10583,N_10444);
xor U13421 (N_13421,N_10124,N_11187);
xor U13422 (N_13422,N_10969,N_9478);
nand U13423 (N_13423,N_11873,N_10116);
nor U13424 (N_13424,N_11273,N_9801);
nor U13425 (N_13425,N_11350,N_9186);
nand U13426 (N_13426,N_10805,N_10682);
or U13427 (N_13427,N_9646,N_9243);
and U13428 (N_13428,N_11464,N_11543);
nor U13429 (N_13429,N_11058,N_11691);
and U13430 (N_13430,N_10555,N_9626);
and U13431 (N_13431,N_11189,N_9525);
or U13432 (N_13432,N_10710,N_11299);
or U13433 (N_13433,N_10790,N_10071);
and U13434 (N_13434,N_11203,N_10172);
nand U13435 (N_13435,N_10263,N_9319);
or U13436 (N_13436,N_10560,N_10928);
nand U13437 (N_13437,N_11849,N_10325);
nand U13438 (N_13438,N_11877,N_11469);
nor U13439 (N_13439,N_10131,N_9591);
or U13440 (N_13440,N_9754,N_11972);
nor U13441 (N_13441,N_9302,N_11549);
nand U13442 (N_13442,N_11512,N_11863);
nand U13443 (N_13443,N_11579,N_10309);
xor U13444 (N_13444,N_9554,N_11049);
and U13445 (N_13445,N_11999,N_11690);
nor U13446 (N_13446,N_10760,N_11063);
or U13447 (N_13447,N_9401,N_10571);
nor U13448 (N_13448,N_11133,N_10652);
xor U13449 (N_13449,N_10336,N_11384);
and U13450 (N_13450,N_11433,N_9664);
xnor U13451 (N_13451,N_11943,N_10939);
nand U13452 (N_13452,N_10966,N_10456);
nor U13453 (N_13453,N_9203,N_11388);
xnor U13454 (N_13454,N_11154,N_11281);
xnor U13455 (N_13455,N_9618,N_10201);
nor U13456 (N_13456,N_9241,N_10379);
or U13457 (N_13457,N_9522,N_11618);
xor U13458 (N_13458,N_10764,N_11732);
or U13459 (N_13459,N_10799,N_10248);
xnor U13460 (N_13460,N_10687,N_10067);
and U13461 (N_13461,N_10187,N_10385);
and U13462 (N_13462,N_11297,N_9863);
nor U13463 (N_13463,N_10279,N_11809);
nand U13464 (N_13464,N_11371,N_10512);
nand U13465 (N_13465,N_10433,N_9479);
xnor U13466 (N_13466,N_9518,N_9439);
and U13467 (N_13467,N_11853,N_9363);
nand U13468 (N_13468,N_11871,N_11179);
xor U13469 (N_13469,N_11993,N_10364);
nand U13470 (N_13470,N_11489,N_9495);
nand U13471 (N_13471,N_11012,N_9583);
or U13472 (N_13472,N_11872,N_10509);
nor U13473 (N_13473,N_9744,N_10795);
nand U13474 (N_13474,N_10563,N_9492);
or U13475 (N_13475,N_9736,N_10420);
and U13476 (N_13476,N_11814,N_9650);
and U13477 (N_13477,N_11673,N_10771);
xor U13478 (N_13478,N_10519,N_10615);
xnor U13479 (N_13479,N_10241,N_11370);
and U13480 (N_13480,N_10029,N_11955);
nand U13481 (N_13481,N_9804,N_11406);
and U13482 (N_13482,N_10829,N_9557);
nand U13483 (N_13483,N_11040,N_10461);
and U13484 (N_13484,N_11652,N_11435);
xnor U13485 (N_13485,N_11356,N_10396);
nand U13486 (N_13486,N_10626,N_11851);
nand U13487 (N_13487,N_11499,N_11687);
or U13488 (N_13488,N_11263,N_11240);
xor U13489 (N_13489,N_11754,N_11650);
nand U13490 (N_13490,N_9813,N_10880);
or U13491 (N_13491,N_9084,N_11899);
and U13492 (N_13492,N_9433,N_10383);
xor U13493 (N_13493,N_11952,N_9160);
nand U13494 (N_13494,N_10585,N_10542);
nand U13495 (N_13495,N_11055,N_9854);
and U13496 (N_13496,N_10680,N_11253);
or U13497 (N_13497,N_9400,N_11519);
xnor U13498 (N_13498,N_9397,N_9073);
xnor U13499 (N_13499,N_11892,N_9265);
nor U13500 (N_13500,N_11578,N_10761);
nor U13501 (N_13501,N_9775,N_10917);
xnor U13502 (N_13502,N_9495,N_11779);
nand U13503 (N_13503,N_11138,N_10361);
nor U13504 (N_13504,N_10904,N_9982);
or U13505 (N_13505,N_10854,N_11605);
xor U13506 (N_13506,N_10803,N_9881);
nor U13507 (N_13507,N_10749,N_9891);
nand U13508 (N_13508,N_10867,N_10722);
or U13509 (N_13509,N_9988,N_9053);
and U13510 (N_13510,N_10447,N_9666);
and U13511 (N_13511,N_11248,N_11735);
and U13512 (N_13512,N_11554,N_10676);
and U13513 (N_13513,N_11387,N_11770);
nor U13514 (N_13514,N_11960,N_10407);
nand U13515 (N_13515,N_9561,N_9237);
nor U13516 (N_13516,N_10484,N_10641);
nand U13517 (N_13517,N_11682,N_11186);
and U13518 (N_13518,N_9081,N_11378);
xnor U13519 (N_13519,N_9098,N_11360);
nor U13520 (N_13520,N_9195,N_11284);
nor U13521 (N_13521,N_10093,N_11533);
or U13522 (N_13522,N_10420,N_10164);
or U13523 (N_13523,N_11532,N_11376);
nand U13524 (N_13524,N_9685,N_9148);
and U13525 (N_13525,N_9021,N_9787);
nor U13526 (N_13526,N_9797,N_10463);
and U13527 (N_13527,N_10106,N_11182);
or U13528 (N_13528,N_11727,N_9129);
and U13529 (N_13529,N_11144,N_10349);
and U13530 (N_13530,N_9840,N_11193);
and U13531 (N_13531,N_10926,N_11948);
xor U13532 (N_13532,N_9521,N_9305);
nor U13533 (N_13533,N_10021,N_11040);
nand U13534 (N_13534,N_11913,N_11597);
and U13535 (N_13535,N_11347,N_10051);
nand U13536 (N_13536,N_9156,N_9607);
xnor U13537 (N_13537,N_9337,N_9977);
or U13538 (N_13538,N_9158,N_9008);
and U13539 (N_13539,N_11961,N_10988);
or U13540 (N_13540,N_9442,N_11632);
xnor U13541 (N_13541,N_9143,N_11269);
or U13542 (N_13542,N_11358,N_9861);
or U13543 (N_13543,N_11519,N_11221);
and U13544 (N_13544,N_9013,N_11761);
xor U13545 (N_13545,N_9869,N_11539);
and U13546 (N_13546,N_9412,N_9152);
or U13547 (N_13547,N_11508,N_10491);
nand U13548 (N_13548,N_10601,N_11668);
nand U13549 (N_13549,N_9263,N_11585);
or U13550 (N_13550,N_11787,N_11593);
xor U13551 (N_13551,N_10840,N_10945);
xnor U13552 (N_13552,N_11770,N_10581);
nor U13553 (N_13553,N_10623,N_9244);
nor U13554 (N_13554,N_11673,N_11096);
nand U13555 (N_13555,N_10197,N_10310);
xnor U13556 (N_13556,N_10760,N_9210);
nand U13557 (N_13557,N_11478,N_9832);
and U13558 (N_13558,N_11450,N_11174);
nor U13559 (N_13559,N_10482,N_9586);
and U13560 (N_13560,N_10915,N_10008);
and U13561 (N_13561,N_11694,N_9688);
nor U13562 (N_13562,N_10778,N_11601);
xnor U13563 (N_13563,N_10861,N_11660);
nor U13564 (N_13564,N_11187,N_9214);
and U13565 (N_13565,N_10612,N_9071);
xnor U13566 (N_13566,N_9376,N_9832);
xor U13567 (N_13567,N_11431,N_10397);
xnor U13568 (N_13568,N_9790,N_10665);
xor U13569 (N_13569,N_11879,N_10140);
xnor U13570 (N_13570,N_10596,N_9400);
xor U13571 (N_13571,N_10018,N_11601);
nor U13572 (N_13572,N_9385,N_10283);
nor U13573 (N_13573,N_9713,N_11058);
and U13574 (N_13574,N_9111,N_10185);
nor U13575 (N_13575,N_9551,N_10207);
nor U13576 (N_13576,N_9705,N_9534);
nand U13577 (N_13577,N_9567,N_10199);
and U13578 (N_13578,N_10591,N_10378);
nand U13579 (N_13579,N_11502,N_10184);
nand U13580 (N_13580,N_10569,N_11911);
xor U13581 (N_13581,N_9927,N_10668);
and U13582 (N_13582,N_11113,N_9179);
xnor U13583 (N_13583,N_11774,N_9584);
nor U13584 (N_13584,N_9961,N_11693);
nand U13585 (N_13585,N_9379,N_9332);
xor U13586 (N_13586,N_11717,N_10678);
nand U13587 (N_13587,N_9756,N_10262);
nor U13588 (N_13588,N_10347,N_9424);
xor U13589 (N_13589,N_9622,N_11879);
nand U13590 (N_13590,N_11424,N_10046);
or U13591 (N_13591,N_9946,N_11037);
and U13592 (N_13592,N_11231,N_11342);
xnor U13593 (N_13593,N_11223,N_11922);
nor U13594 (N_13594,N_10349,N_10626);
and U13595 (N_13595,N_11627,N_11950);
or U13596 (N_13596,N_9500,N_9763);
xor U13597 (N_13597,N_9010,N_11216);
or U13598 (N_13598,N_11829,N_9015);
nor U13599 (N_13599,N_10023,N_9826);
nor U13600 (N_13600,N_9745,N_9683);
and U13601 (N_13601,N_9064,N_11258);
and U13602 (N_13602,N_11811,N_11984);
and U13603 (N_13603,N_9409,N_11846);
or U13604 (N_13604,N_9970,N_10255);
or U13605 (N_13605,N_10619,N_11315);
nand U13606 (N_13606,N_11304,N_9888);
xnor U13607 (N_13607,N_9578,N_11928);
nand U13608 (N_13608,N_11360,N_11032);
xnor U13609 (N_13609,N_10456,N_9872);
nand U13610 (N_13610,N_11879,N_11522);
xnor U13611 (N_13611,N_9329,N_11458);
or U13612 (N_13612,N_11916,N_11005);
xor U13613 (N_13613,N_10905,N_10067);
xnor U13614 (N_13614,N_9584,N_9430);
xnor U13615 (N_13615,N_11848,N_10952);
nor U13616 (N_13616,N_10139,N_11361);
and U13617 (N_13617,N_9410,N_10526);
or U13618 (N_13618,N_10392,N_11779);
xor U13619 (N_13619,N_10890,N_11793);
nand U13620 (N_13620,N_11205,N_11128);
nand U13621 (N_13621,N_10013,N_9344);
xor U13622 (N_13622,N_10431,N_9777);
xor U13623 (N_13623,N_11544,N_9664);
nand U13624 (N_13624,N_9105,N_10061);
nand U13625 (N_13625,N_11146,N_10180);
nor U13626 (N_13626,N_9737,N_11216);
or U13627 (N_13627,N_10374,N_11646);
nand U13628 (N_13628,N_10077,N_11568);
nand U13629 (N_13629,N_10826,N_9114);
nor U13630 (N_13630,N_10704,N_9216);
xor U13631 (N_13631,N_10786,N_10657);
xor U13632 (N_13632,N_11467,N_11460);
nor U13633 (N_13633,N_11986,N_9835);
nand U13634 (N_13634,N_11848,N_10288);
nand U13635 (N_13635,N_9251,N_9334);
or U13636 (N_13636,N_11894,N_11394);
or U13637 (N_13637,N_10711,N_9776);
and U13638 (N_13638,N_10578,N_10780);
nand U13639 (N_13639,N_9894,N_9022);
and U13640 (N_13640,N_11163,N_9666);
or U13641 (N_13641,N_9917,N_9266);
and U13642 (N_13642,N_11306,N_10035);
xor U13643 (N_13643,N_11019,N_9929);
or U13644 (N_13644,N_10545,N_9226);
or U13645 (N_13645,N_10250,N_10607);
and U13646 (N_13646,N_9505,N_10256);
nand U13647 (N_13647,N_11822,N_11739);
nand U13648 (N_13648,N_9951,N_10891);
or U13649 (N_13649,N_10287,N_11714);
or U13650 (N_13650,N_9747,N_10911);
or U13651 (N_13651,N_9463,N_9411);
nor U13652 (N_13652,N_9662,N_10915);
xnor U13653 (N_13653,N_11559,N_10732);
or U13654 (N_13654,N_9152,N_11935);
xnor U13655 (N_13655,N_9401,N_10643);
xor U13656 (N_13656,N_11428,N_9844);
or U13657 (N_13657,N_10374,N_11487);
nor U13658 (N_13658,N_9957,N_11256);
nor U13659 (N_13659,N_9936,N_10371);
xor U13660 (N_13660,N_9956,N_10269);
xor U13661 (N_13661,N_11572,N_9199);
nand U13662 (N_13662,N_10744,N_10434);
nand U13663 (N_13663,N_9501,N_11511);
nor U13664 (N_13664,N_9106,N_9913);
or U13665 (N_13665,N_10228,N_9266);
xor U13666 (N_13666,N_11902,N_11471);
or U13667 (N_13667,N_11036,N_11507);
nand U13668 (N_13668,N_9183,N_9564);
xor U13669 (N_13669,N_11811,N_9213);
and U13670 (N_13670,N_9639,N_11465);
and U13671 (N_13671,N_10636,N_9824);
xnor U13672 (N_13672,N_9138,N_11055);
nand U13673 (N_13673,N_10516,N_11968);
nor U13674 (N_13674,N_10653,N_9612);
nor U13675 (N_13675,N_10658,N_11480);
nor U13676 (N_13676,N_10794,N_9217);
nor U13677 (N_13677,N_9260,N_10690);
nand U13678 (N_13678,N_11225,N_10767);
or U13679 (N_13679,N_9242,N_11702);
and U13680 (N_13680,N_10653,N_11626);
xor U13681 (N_13681,N_9260,N_10606);
or U13682 (N_13682,N_10595,N_10706);
or U13683 (N_13683,N_11960,N_9648);
xor U13684 (N_13684,N_9683,N_9865);
nor U13685 (N_13685,N_10994,N_10423);
nor U13686 (N_13686,N_9685,N_9665);
xnor U13687 (N_13687,N_11879,N_10446);
xor U13688 (N_13688,N_9166,N_10163);
xnor U13689 (N_13689,N_9493,N_9262);
nor U13690 (N_13690,N_10585,N_11395);
xnor U13691 (N_13691,N_9934,N_11969);
xor U13692 (N_13692,N_9860,N_10558);
or U13693 (N_13693,N_9399,N_10770);
nor U13694 (N_13694,N_9743,N_10054);
and U13695 (N_13695,N_10805,N_10487);
and U13696 (N_13696,N_11544,N_10752);
and U13697 (N_13697,N_10010,N_10940);
nand U13698 (N_13698,N_9198,N_9919);
nor U13699 (N_13699,N_11452,N_11998);
xnor U13700 (N_13700,N_10309,N_10274);
nand U13701 (N_13701,N_9555,N_11868);
nand U13702 (N_13702,N_10904,N_11405);
xnor U13703 (N_13703,N_11386,N_11611);
nand U13704 (N_13704,N_9219,N_9168);
or U13705 (N_13705,N_10879,N_10424);
or U13706 (N_13706,N_11421,N_11678);
and U13707 (N_13707,N_11746,N_10257);
nand U13708 (N_13708,N_10258,N_11977);
nor U13709 (N_13709,N_9707,N_11439);
or U13710 (N_13710,N_11934,N_9787);
nand U13711 (N_13711,N_10762,N_11147);
nand U13712 (N_13712,N_11326,N_11181);
xnor U13713 (N_13713,N_9683,N_11202);
or U13714 (N_13714,N_11113,N_9471);
xnor U13715 (N_13715,N_10883,N_9258);
xor U13716 (N_13716,N_9452,N_10876);
and U13717 (N_13717,N_9033,N_10566);
or U13718 (N_13718,N_11514,N_10388);
nand U13719 (N_13719,N_11363,N_9250);
nor U13720 (N_13720,N_9813,N_9070);
xnor U13721 (N_13721,N_10208,N_10452);
nor U13722 (N_13722,N_10891,N_11658);
or U13723 (N_13723,N_9135,N_9921);
or U13724 (N_13724,N_11057,N_9072);
and U13725 (N_13725,N_11061,N_10286);
nand U13726 (N_13726,N_9161,N_9359);
nand U13727 (N_13727,N_10984,N_11483);
nand U13728 (N_13728,N_11915,N_10185);
nand U13729 (N_13729,N_9749,N_9926);
xnor U13730 (N_13730,N_10333,N_11556);
and U13731 (N_13731,N_11352,N_11485);
or U13732 (N_13732,N_9413,N_9367);
nand U13733 (N_13733,N_10895,N_10856);
nand U13734 (N_13734,N_9285,N_10836);
or U13735 (N_13735,N_11855,N_10620);
nor U13736 (N_13736,N_10662,N_11709);
nor U13737 (N_13737,N_11442,N_10776);
or U13738 (N_13738,N_9589,N_10760);
xnor U13739 (N_13739,N_10554,N_9880);
nor U13740 (N_13740,N_9024,N_9898);
or U13741 (N_13741,N_9679,N_10663);
nor U13742 (N_13742,N_9824,N_9491);
nand U13743 (N_13743,N_10143,N_11921);
xor U13744 (N_13744,N_11129,N_11937);
nand U13745 (N_13745,N_10352,N_10670);
and U13746 (N_13746,N_11529,N_10267);
nand U13747 (N_13747,N_9597,N_10468);
or U13748 (N_13748,N_10264,N_9534);
xnor U13749 (N_13749,N_11832,N_10013);
nor U13750 (N_13750,N_11609,N_10044);
or U13751 (N_13751,N_11310,N_9142);
and U13752 (N_13752,N_10928,N_10866);
xnor U13753 (N_13753,N_10765,N_10434);
nor U13754 (N_13754,N_11644,N_11891);
or U13755 (N_13755,N_10839,N_11557);
or U13756 (N_13756,N_9856,N_9291);
nand U13757 (N_13757,N_10569,N_9882);
or U13758 (N_13758,N_10332,N_11146);
or U13759 (N_13759,N_11390,N_9391);
and U13760 (N_13760,N_10139,N_10372);
nor U13761 (N_13761,N_10337,N_10589);
or U13762 (N_13762,N_10227,N_11658);
nor U13763 (N_13763,N_10568,N_11127);
and U13764 (N_13764,N_9498,N_10523);
and U13765 (N_13765,N_10160,N_11812);
nor U13766 (N_13766,N_10057,N_11398);
and U13767 (N_13767,N_11998,N_11240);
and U13768 (N_13768,N_11313,N_10863);
or U13769 (N_13769,N_10575,N_9766);
or U13770 (N_13770,N_11503,N_11456);
nand U13771 (N_13771,N_9106,N_9092);
xor U13772 (N_13772,N_10375,N_9394);
and U13773 (N_13773,N_11362,N_11201);
nor U13774 (N_13774,N_9580,N_9208);
nand U13775 (N_13775,N_10119,N_10769);
and U13776 (N_13776,N_11541,N_11085);
xor U13777 (N_13777,N_10336,N_9465);
and U13778 (N_13778,N_10986,N_11285);
nand U13779 (N_13779,N_11427,N_10395);
xnor U13780 (N_13780,N_10870,N_9028);
nor U13781 (N_13781,N_10780,N_9156);
nand U13782 (N_13782,N_9269,N_11678);
and U13783 (N_13783,N_11916,N_11840);
or U13784 (N_13784,N_10343,N_9599);
and U13785 (N_13785,N_11069,N_10587);
and U13786 (N_13786,N_10252,N_9266);
nand U13787 (N_13787,N_9806,N_10963);
or U13788 (N_13788,N_10942,N_11856);
or U13789 (N_13789,N_9942,N_10585);
nand U13790 (N_13790,N_10354,N_9893);
nand U13791 (N_13791,N_10724,N_9322);
xnor U13792 (N_13792,N_9906,N_10939);
nor U13793 (N_13793,N_11457,N_9328);
or U13794 (N_13794,N_11716,N_11142);
nand U13795 (N_13795,N_9539,N_9493);
or U13796 (N_13796,N_10015,N_10061);
and U13797 (N_13797,N_11683,N_10616);
xnor U13798 (N_13798,N_10949,N_9220);
and U13799 (N_13799,N_11980,N_9272);
xor U13800 (N_13800,N_10312,N_11466);
and U13801 (N_13801,N_9861,N_9197);
nand U13802 (N_13802,N_9953,N_10241);
or U13803 (N_13803,N_11823,N_9413);
nor U13804 (N_13804,N_9146,N_11125);
xor U13805 (N_13805,N_11070,N_11069);
or U13806 (N_13806,N_9897,N_9431);
or U13807 (N_13807,N_11783,N_9858);
nand U13808 (N_13808,N_9363,N_9848);
nand U13809 (N_13809,N_9153,N_11673);
nand U13810 (N_13810,N_9866,N_9145);
nor U13811 (N_13811,N_10184,N_9707);
nand U13812 (N_13812,N_11299,N_10343);
or U13813 (N_13813,N_11210,N_11915);
nor U13814 (N_13814,N_9684,N_10276);
nand U13815 (N_13815,N_9681,N_9417);
nand U13816 (N_13816,N_10406,N_9875);
nor U13817 (N_13817,N_11734,N_10564);
xnor U13818 (N_13818,N_9961,N_9838);
nand U13819 (N_13819,N_11804,N_9564);
nor U13820 (N_13820,N_10675,N_10147);
xor U13821 (N_13821,N_10276,N_10662);
and U13822 (N_13822,N_10924,N_11540);
nor U13823 (N_13823,N_10207,N_10077);
xnor U13824 (N_13824,N_11813,N_11139);
or U13825 (N_13825,N_10491,N_11515);
or U13826 (N_13826,N_10418,N_9967);
or U13827 (N_13827,N_11797,N_10567);
or U13828 (N_13828,N_11487,N_10678);
xor U13829 (N_13829,N_11597,N_11475);
and U13830 (N_13830,N_9762,N_10037);
or U13831 (N_13831,N_9117,N_10096);
or U13832 (N_13832,N_11169,N_10009);
or U13833 (N_13833,N_10579,N_10375);
nand U13834 (N_13834,N_10584,N_11146);
or U13835 (N_13835,N_9166,N_9778);
nand U13836 (N_13836,N_10010,N_9791);
nand U13837 (N_13837,N_10114,N_10763);
xnor U13838 (N_13838,N_9512,N_10549);
or U13839 (N_13839,N_9766,N_9609);
nand U13840 (N_13840,N_10627,N_11122);
nand U13841 (N_13841,N_9299,N_11795);
nor U13842 (N_13842,N_10297,N_10533);
xnor U13843 (N_13843,N_9571,N_10233);
nand U13844 (N_13844,N_9922,N_9759);
xnor U13845 (N_13845,N_11043,N_10818);
nor U13846 (N_13846,N_10946,N_10586);
or U13847 (N_13847,N_10065,N_10938);
and U13848 (N_13848,N_10403,N_10092);
nand U13849 (N_13849,N_11704,N_9416);
and U13850 (N_13850,N_11278,N_11043);
xor U13851 (N_13851,N_9513,N_9146);
nand U13852 (N_13852,N_11359,N_10972);
or U13853 (N_13853,N_10065,N_9769);
and U13854 (N_13854,N_10672,N_9863);
nor U13855 (N_13855,N_9068,N_10814);
nand U13856 (N_13856,N_9016,N_11465);
nor U13857 (N_13857,N_10496,N_9393);
nand U13858 (N_13858,N_10755,N_10471);
nor U13859 (N_13859,N_11147,N_9655);
xor U13860 (N_13860,N_11959,N_11439);
and U13861 (N_13861,N_9505,N_11182);
or U13862 (N_13862,N_11894,N_9151);
nor U13863 (N_13863,N_10716,N_10509);
and U13864 (N_13864,N_9631,N_10712);
and U13865 (N_13865,N_11348,N_11355);
nor U13866 (N_13866,N_10108,N_9207);
nand U13867 (N_13867,N_11797,N_9298);
and U13868 (N_13868,N_11228,N_9232);
and U13869 (N_13869,N_10327,N_10406);
or U13870 (N_13870,N_9996,N_10745);
or U13871 (N_13871,N_10231,N_11071);
and U13872 (N_13872,N_11972,N_10475);
nor U13873 (N_13873,N_9242,N_9793);
and U13874 (N_13874,N_11793,N_10144);
and U13875 (N_13875,N_10818,N_11193);
nor U13876 (N_13876,N_9799,N_9873);
and U13877 (N_13877,N_11979,N_11747);
nor U13878 (N_13878,N_10692,N_11067);
nand U13879 (N_13879,N_9753,N_9654);
and U13880 (N_13880,N_11816,N_9457);
and U13881 (N_13881,N_11706,N_11962);
and U13882 (N_13882,N_9972,N_9941);
or U13883 (N_13883,N_10203,N_9549);
or U13884 (N_13884,N_10628,N_11508);
nand U13885 (N_13885,N_10868,N_11612);
xnor U13886 (N_13886,N_9373,N_10504);
nor U13887 (N_13887,N_9421,N_11904);
nand U13888 (N_13888,N_9390,N_11802);
nand U13889 (N_13889,N_9982,N_9294);
or U13890 (N_13890,N_9573,N_10080);
nor U13891 (N_13891,N_9275,N_9861);
nand U13892 (N_13892,N_10967,N_11963);
xor U13893 (N_13893,N_10895,N_11029);
and U13894 (N_13894,N_10499,N_9466);
or U13895 (N_13895,N_11072,N_11689);
and U13896 (N_13896,N_11378,N_11426);
xnor U13897 (N_13897,N_11981,N_11185);
xor U13898 (N_13898,N_9478,N_9849);
nand U13899 (N_13899,N_11704,N_10851);
nor U13900 (N_13900,N_9082,N_10293);
or U13901 (N_13901,N_10207,N_9956);
xnor U13902 (N_13902,N_11581,N_11804);
xor U13903 (N_13903,N_10285,N_10554);
and U13904 (N_13904,N_10023,N_10674);
nor U13905 (N_13905,N_10124,N_10230);
nand U13906 (N_13906,N_10336,N_9520);
nand U13907 (N_13907,N_9332,N_9839);
nor U13908 (N_13908,N_9064,N_11667);
or U13909 (N_13909,N_9320,N_10992);
nor U13910 (N_13910,N_11200,N_11844);
or U13911 (N_13911,N_11135,N_10368);
or U13912 (N_13912,N_11930,N_9921);
or U13913 (N_13913,N_9304,N_11693);
or U13914 (N_13914,N_11324,N_9742);
xnor U13915 (N_13915,N_10103,N_10590);
nor U13916 (N_13916,N_9140,N_9868);
nor U13917 (N_13917,N_9614,N_11386);
xnor U13918 (N_13918,N_11205,N_9129);
xor U13919 (N_13919,N_11412,N_10243);
nand U13920 (N_13920,N_10877,N_10780);
nand U13921 (N_13921,N_11994,N_11262);
nor U13922 (N_13922,N_11264,N_10117);
nand U13923 (N_13923,N_10257,N_10940);
nor U13924 (N_13924,N_10082,N_9416);
or U13925 (N_13925,N_11408,N_11026);
or U13926 (N_13926,N_9072,N_10826);
nor U13927 (N_13927,N_9820,N_11779);
and U13928 (N_13928,N_9100,N_11907);
nand U13929 (N_13929,N_11580,N_9123);
nand U13930 (N_13930,N_10587,N_9767);
or U13931 (N_13931,N_9050,N_9726);
and U13932 (N_13932,N_9920,N_11069);
nand U13933 (N_13933,N_11511,N_11170);
nor U13934 (N_13934,N_9900,N_9845);
nor U13935 (N_13935,N_11018,N_9383);
xnor U13936 (N_13936,N_9919,N_9566);
or U13937 (N_13937,N_10439,N_9589);
nor U13938 (N_13938,N_10346,N_11747);
or U13939 (N_13939,N_9660,N_11777);
nand U13940 (N_13940,N_9408,N_11855);
xor U13941 (N_13941,N_9122,N_11027);
xnor U13942 (N_13942,N_9853,N_10466);
and U13943 (N_13943,N_9505,N_9266);
xnor U13944 (N_13944,N_11364,N_9109);
xor U13945 (N_13945,N_9002,N_10002);
nor U13946 (N_13946,N_10423,N_10519);
nor U13947 (N_13947,N_10004,N_9260);
nand U13948 (N_13948,N_10313,N_10091);
xor U13949 (N_13949,N_10641,N_10381);
and U13950 (N_13950,N_11730,N_11639);
xnor U13951 (N_13951,N_11283,N_11919);
nand U13952 (N_13952,N_9079,N_10814);
nor U13953 (N_13953,N_9539,N_9374);
or U13954 (N_13954,N_11910,N_11823);
and U13955 (N_13955,N_11731,N_9450);
nand U13956 (N_13956,N_10406,N_10083);
nand U13957 (N_13957,N_9037,N_9813);
nor U13958 (N_13958,N_10335,N_11028);
xnor U13959 (N_13959,N_10702,N_10193);
xor U13960 (N_13960,N_10297,N_9095);
nor U13961 (N_13961,N_9607,N_11865);
nand U13962 (N_13962,N_11214,N_10296);
xor U13963 (N_13963,N_9210,N_10032);
and U13964 (N_13964,N_9997,N_11133);
or U13965 (N_13965,N_9071,N_10035);
nor U13966 (N_13966,N_9746,N_11790);
xor U13967 (N_13967,N_10065,N_9654);
nor U13968 (N_13968,N_11688,N_10053);
xor U13969 (N_13969,N_9844,N_9625);
and U13970 (N_13970,N_11610,N_9112);
nand U13971 (N_13971,N_9287,N_11205);
or U13972 (N_13972,N_9644,N_9051);
nor U13973 (N_13973,N_9102,N_11399);
nor U13974 (N_13974,N_9540,N_11410);
nor U13975 (N_13975,N_11756,N_9161);
xnor U13976 (N_13976,N_9251,N_10622);
xor U13977 (N_13977,N_10157,N_9241);
nand U13978 (N_13978,N_9923,N_11265);
xor U13979 (N_13979,N_10220,N_11766);
nor U13980 (N_13980,N_9131,N_10389);
xor U13981 (N_13981,N_11358,N_11291);
and U13982 (N_13982,N_10023,N_11316);
xnor U13983 (N_13983,N_11733,N_10534);
nor U13984 (N_13984,N_10445,N_9190);
or U13985 (N_13985,N_11234,N_11805);
or U13986 (N_13986,N_9230,N_9021);
xnor U13987 (N_13987,N_9965,N_11899);
or U13988 (N_13988,N_11369,N_9486);
or U13989 (N_13989,N_11235,N_10021);
nand U13990 (N_13990,N_11791,N_10876);
or U13991 (N_13991,N_11914,N_9250);
and U13992 (N_13992,N_9421,N_9386);
nand U13993 (N_13993,N_9197,N_11624);
nand U13994 (N_13994,N_9659,N_11999);
nand U13995 (N_13995,N_10354,N_10353);
nor U13996 (N_13996,N_10388,N_10221);
and U13997 (N_13997,N_10044,N_10732);
and U13998 (N_13998,N_9161,N_9895);
and U13999 (N_13999,N_11912,N_9412);
nand U14000 (N_14000,N_11076,N_10790);
xor U14001 (N_14001,N_9303,N_9733);
and U14002 (N_14002,N_9796,N_11450);
xnor U14003 (N_14003,N_11444,N_9326);
nand U14004 (N_14004,N_11410,N_9710);
xnor U14005 (N_14005,N_9994,N_10712);
nand U14006 (N_14006,N_11840,N_10090);
nand U14007 (N_14007,N_9960,N_9375);
nand U14008 (N_14008,N_10711,N_10811);
xnor U14009 (N_14009,N_11841,N_11169);
nor U14010 (N_14010,N_10691,N_11017);
nor U14011 (N_14011,N_11219,N_9204);
nor U14012 (N_14012,N_11303,N_9376);
nor U14013 (N_14013,N_11709,N_9034);
nor U14014 (N_14014,N_11813,N_9787);
or U14015 (N_14015,N_9787,N_9537);
nor U14016 (N_14016,N_9157,N_9842);
xnor U14017 (N_14017,N_11008,N_10724);
nand U14018 (N_14018,N_10873,N_9286);
or U14019 (N_14019,N_11239,N_9731);
or U14020 (N_14020,N_10689,N_9037);
and U14021 (N_14021,N_11499,N_11405);
and U14022 (N_14022,N_9852,N_10640);
and U14023 (N_14023,N_11610,N_9907);
nor U14024 (N_14024,N_10457,N_10990);
and U14025 (N_14025,N_10277,N_9090);
nand U14026 (N_14026,N_9983,N_11039);
xor U14027 (N_14027,N_10049,N_10689);
xnor U14028 (N_14028,N_11393,N_11959);
nand U14029 (N_14029,N_10628,N_11352);
nand U14030 (N_14030,N_10349,N_10589);
or U14031 (N_14031,N_10264,N_9143);
xnor U14032 (N_14032,N_9409,N_11574);
nor U14033 (N_14033,N_10378,N_9612);
nand U14034 (N_14034,N_10412,N_10589);
or U14035 (N_14035,N_10321,N_9457);
xnor U14036 (N_14036,N_9418,N_10996);
and U14037 (N_14037,N_9271,N_9053);
or U14038 (N_14038,N_11783,N_9091);
xnor U14039 (N_14039,N_9346,N_11598);
and U14040 (N_14040,N_11850,N_10788);
and U14041 (N_14041,N_10738,N_11704);
and U14042 (N_14042,N_11512,N_10362);
or U14043 (N_14043,N_10783,N_11696);
xor U14044 (N_14044,N_11935,N_11613);
and U14045 (N_14045,N_11518,N_10732);
and U14046 (N_14046,N_11469,N_10413);
and U14047 (N_14047,N_11739,N_9872);
and U14048 (N_14048,N_9728,N_10227);
nand U14049 (N_14049,N_11099,N_10293);
xor U14050 (N_14050,N_9671,N_11672);
nand U14051 (N_14051,N_10231,N_9335);
nand U14052 (N_14052,N_10299,N_9812);
xnor U14053 (N_14053,N_10592,N_10142);
and U14054 (N_14054,N_11438,N_9702);
nand U14055 (N_14055,N_10269,N_9157);
nand U14056 (N_14056,N_10592,N_11726);
nor U14057 (N_14057,N_11896,N_11138);
nor U14058 (N_14058,N_9272,N_10799);
xnor U14059 (N_14059,N_9590,N_9255);
xnor U14060 (N_14060,N_9311,N_9931);
and U14061 (N_14061,N_9823,N_9811);
or U14062 (N_14062,N_9018,N_11235);
or U14063 (N_14063,N_9463,N_11434);
nand U14064 (N_14064,N_11407,N_9851);
nor U14065 (N_14065,N_9850,N_10274);
and U14066 (N_14066,N_11377,N_10836);
and U14067 (N_14067,N_10287,N_11721);
nand U14068 (N_14068,N_9653,N_9855);
nand U14069 (N_14069,N_9359,N_10955);
nand U14070 (N_14070,N_9580,N_9180);
xnor U14071 (N_14071,N_11978,N_11182);
and U14072 (N_14072,N_9166,N_10770);
nand U14073 (N_14073,N_11271,N_9828);
xnor U14074 (N_14074,N_10969,N_11811);
and U14075 (N_14075,N_9138,N_9563);
nor U14076 (N_14076,N_10956,N_11837);
nor U14077 (N_14077,N_11547,N_9073);
and U14078 (N_14078,N_9388,N_11920);
nand U14079 (N_14079,N_10686,N_11340);
nand U14080 (N_14080,N_10640,N_11173);
xor U14081 (N_14081,N_10536,N_9632);
nor U14082 (N_14082,N_10603,N_10810);
nor U14083 (N_14083,N_9164,N_11146);
nor U14084 (N_14084,N_10772,N_10717);
nor U14085 (N_14085,N_9066,N_11826);
nor U14086 (N_14086,N_9274,N_10588);
or U14087 (N_14087,N_9687,N_10070);
nand U14088 (N_14088,N_11222,N_10683);
and U14089 (N_14089,N_9489,N_11319);
or U14090 (N_14090,N_10209,N_9424);
nand U14091 (N_14091,N_10164,N_9117);
nand U14092 (N_14092,N_9327,N_11388);
and U14093 (N_14093,N_11244,N_9602);
and U14094 (N_14094,N_10897,N_9081);
and U14095 (N_14095,N_10848,N_10572);
xor U14096 (N_14096,N_11067,N_10300);
nand U14097 (N_14097,N_11684,N_11912);
nand U14098 (N_14098,N_9419,N_10552);
nand U14099 (N_14099,N_10299,N_10950);
or U14100 (N_14100,N_11149,N_9099);
nand U14101 (N_14101,N_10309,N_10729);
or U14102 (N_14102,N_11005,N_10691);
and U14103 (N_14103,N_10051,N_9578);
and U14104 (N_14104,N_11045,N_10370);
or U14105 (N_14105,N_10809,N_11923);
nor U14106 (N_14106,N_9228,N_9738);
and U14107 (N_14107,N_10894,N_11947);
and U14108 (N_14108,N_9419,N_9099);
xor U14109 (N_14109,N_9467,N_9836);
or U14110 (N_14110,N_11477,N_11735);
nand U14111 (N_14111,N_10717,N_11784);
xor U14112 (N_14112,N_10126,N_11122);
nor U14113 (N_14113,N_11448,N_9875);
or U14114 (N_14114,N_11326,N_9019);
or U14115 (N_14115,N_9241,N_9891);
nand U14116 (N_14116,N_10063,N_11788);
xnor U14117 (N_14117,N_10482,N_11626);
or U14118 (N_14118,N_9500,N_10526);
and U14119 (N_14119,N_9560,N_11437);
nand U14120 (N_14120,N_11473,N_10208);
nand U14121 (N_14121,N_9712,N_11423);
or U14122 (N_14122,N_9307,N_10138);
xnor U14123 (N_14123,N_10630,N_10313);
nor U14124 (N_14124,N_10744,N_11770);
nor U14125 (N_14125,N_9732,N_11197);
and U14126 (N_14126,N_10670,N_10622);
and U14127 (N_14127,N_9096,N_10404);
nor U14128 (N_14128,N_11339,N_10113);
xnor U14129 (N_14129,N_11104,N_11464);
xor U14130 (N_14130,N_11616,N_11714);
nor U14131 (N_14131,N_10117,N_10455);
and U14132 (N_14132,N_11693,N_10846);
and U14133 (N_14133,N_11180,N_9609);
nand U14134 (N_14134,N_9518,N_9104);
nor U14135 (N_14135,N_9840,N_10111);
nor U14136 (N_14136,N_9999,N_9489);
nor U14137 (N_14137,N_11076,N_11088);
nand U14138 (N_14138,N_11563,N_9017);
nand U14139 (N_14139,N_10204,N_11441);
or U14140 (N_14140,N_11626,N_10887);
or U14141 (N_14141,N_11562,N_10854);
or U14142 (N_14142,N_9585,N_10919);
nand U14143 (N_14143,N_9480,N_9069);
nand U14144 (N_14144,N_9174,N_9545);
nor U14145 (N_14145,N_11069,N_10185);
xor U14146 (N_14146,N_10011,N_10322);
nand U14147 (N_14147,N_9334,N_11806);
and U14148 (N_14148,N_9181,N_9422);
or U14149 (N_14149,N_10417,N_10156);
xnor U14150 (N_14150,N_9315,N_11064);
nor U14151 (N_14151,N_10562,N_9385);
or U14152 (N_14152,N_10352,N_9808);
or U14153 (N_14153,N_11156,N_11614);
or U14154 (N_14154,N_9883,N_11294);
xor U14155 (N_14155,N_10236,N_10884);
nor U14156 (N_14156,N_11359,N_9089);
nor U14157 (N_14157,N_10481,N_10633);
nor U14158 (N_14158,N_9238,N_9016);
xor U14159 (N_14159,N_10918,N_11240);
nor U14160 (N_14160,N_9474,N_9158);
xnor U14161 (N_14161,N_9700,N_10053);
xor U14162 (N_14162,N_10885,N_11871);
and U14163 (N_14163,N_9785,N_10629);
nor U14164 (N_14164,N_11145,N_10112);
nor U14165 (N_14165,N_9141,N_9866);
nand U14166 (N_14166,N_11858,N_9738);
or U14167 (N_14167,N_10832,N_10613);
xnor U14168 (N_14168,N_9315,N_9794);
nand U14169 (N_14169,N_9315,N_11266);
nor U14170 (N_14170,N_10156,N_11792);
or U14171 (N_14171,N_11292,N_11507);
nor U14172 (N_14172,N_9490,N_10414);
nor U14173 (N_14173,N_9870,N_9226);
and U14174 (N_14174,N_11599,N_10704);
xor U14175 (N_14175,N_10342,N_11692);
xor U14176 (N_14176,N_9337,N_11704);
nor U14177 (N_14177,N_10460,N_10812);
nor U14178 (N_14178,N_10712,N_11393);
nor U14179 (N_14179,N_9536,N_10620);
or U14180 (N_14180,N_9919,N_10359);
nor U14181 (N_14181,N_10359,N_10979);
nand U14182 (N_14182,N_10347,N_9853);
and U14183 (N_14183,N_11842,N_11650);
and U14184 (N_14184,N_10509,N_10404);
xor U14185 (N_14185,N_11675,N_10651);
or U14186 (N_14186,N_10583,N_10539);
nand U14187 (N_14187,N_10383,N_11595);
nor U14188 (N_14188,N_11601,N_11428);
nor U14189 (N_14189,N_10088,N_9619);
or U14190 (N_14190,N_9461,N_9556);
nand U14191 (N_14191,N_9695,N_11369);
nor U14192 (N_14192,N_9969,N_11736);
nand U14193 (N_14193,N_11663,N_9859);
or U14194 (N_14194,N_11625,N_11397);
nand U14195 (N_14195,N_11617,N_10334);
nand U14196 (N_14196,N_9808,N_9942);
nand U14197 (N_14197,N_11643,N_9848);
nand U14198 (N_14198,N_11522,N_9450);
and U14199 (N_14199,N_9339,N_9947);
nand U14200 (N_14200,N_10749,N_11873);
nand U14201 (N_14201,N_9879,N_11983);
xnor U14202 (N_14202,N_9861,N_10501);
or U14203 (N_14203,N_11332,N_10735);
or U14204 (N_14204,N_10106,N_9321);
and U14205 (N_14205,N_10480,N_11013);
xnor U14206 (N_14206,N_9770,N_11199);
or U14207 (N_14207,N_11227,N_11766);
and U14208 (N_14208,N_10542,N_10367);
nand U14209 (N_14209,N_10669,N_10640);
xor U14210 (N_14210,N_11256,N_9114);
xor U14211 (N_14211,N_11440,N_10689);
nand U14212 (N_14212,N_11794,N_9595);
and U14213 (N_14213,N_9350,N_11750);
nand U14214 (N_14214,N_11059,N_10232);
and U14215 (N_14215,N_10902,N_9437);
xor U14216 (N_14216,N_11665,N_11496);
xor U14217 (N_14217,N_9756,N_11363);
xor U14218 (N_14218,N_10814,N_10913);
xor U14219 (N_14219,N_9323,N_10787);
xor U14220 (N_14220,N_9928,N_11527);
and U14221 (N_14221,N_10659,N_9908);
and U14222 (N_14222,N_9864,N_9911);
or U14223 (N_14223,N_9824,N_9822);
and U14224 (N_14224,N_9087,N_9979);
and U14225 (N_14225,N_11092,N_9895);
nand U14226 (N_14226,N_10461,N_10343);
nor U14227 (N_14227,N_10410,N_9873);
nand U14228 (N_14228,N_9364,N_11121);
or U14229 (N_14229,N_11145,N_9917);
nor U14230 (N_14230,N_11859,N_10014);
nor U14231 (N_14231,N_11309,N_10456);
xor U14232 (N_14232,N_11379,N_9573);
nand U14233 (N_14233,N_10577,N_11576);
nand U14234 (N_14234,N_10504,N_11621);
nor U14235 (N_14235,N_10452,N_10221);
xor U14236 (N_14236,N_9003,N_9594);
and U14237 (N_14237,N_11387,N_10081);
nor U14238 (N_14238,N_9846,N_9244);
and U14239 (N_14239,N_11707,N_9020);
nor U14240 (N_14240,N_9989,N_11769);
or U14241 (N_14241,N_10524,N_9906);
nand U14242 (N_14242,N_11387,N_11732);
xnor U14243 (N_14243,N_11177,N_9668);
and U14244 (N_14244,N_11392,N_9446);
or U14245 (N_14245,N_11687,N_9066);
nor U14246 (N_14246,N_10470,N_9549);
or U14247 (N_14247,N_11946,N_11398);
nand U14248 (N_14248,N_10062,N_10522);
nor U14249 (N_14249,N_11819,N_11902);
nor U14250 (N_14250,N_11744,N_10951);
nor U14251 (N_14251,N_9035,N_11786);
and U14252 (N_14252,N_11392,N_10608);
and U14253 (N_14253,N_11708,N_11618);
xor U14254 (N_14254,N_10123,N_11492);
nand U14255 (N_14255,N_11369,N_9295);
nor U14256 (N_14256,N_11299,N_9615);
xnor U14257 (N_14257,N_10309,N_10620);
nor U14258 (N_14258,N_10015,N_9072);
xor U14259 (N_14259,N_11075,N_9104);
nand U14260 (N_14260,N_10571,N_11933);
xnor U14261 (N_14261,N_10050,N_10128);
xor U14262 (N_14262,N_10120,N_10470);
or U14263 (N_14263,N_11431,N_11425);
and U14264 (N_14264,N_10080,N_9305);
nor U14265 (N_14265,N_10691,N_11793);
nand U14266 (N_14266,N_9836,N_10866);
xnor U14267 (N_14267,N_9123,N_10982);
or U14268 (N_14268,N_9727,N_9056);
nor U14269 (N_14269,N_10627,N_11138);
nand U14270 (N_14270,N_10654,N_9711);
or U14271 (N_14271,N_9904,N_9206);
nor U14272 (N_14272,N_11562,N_9837);
xor U14273 (N_14273,N_9813,N_9571);
nand U14274 (N_14274,N_9541,N_10409);
and U14275 (N_14275,N_10407,N_11717);
xor U14276 (N_14276,N_10884,N_10160);
xnor U14277 (N_14277,N_9997,N_9327);
xor U14278 (N_14278,N_9167,N_10032);
nand U14279 (N_14279,N_11665,N_10135);
nor U14280 (N_14280,N_10386,N_11910);
nand U14281 (N_14281,N_11188,N_10748);
and U14282 (N_14282,N_9998,N_11300);
nand U14283 (N_14283,N_9417,N_11512);
and U14284 (N_14284,N_9643,N_11191);
or U14285 (N_14285,N_11761,N_11496);
nor U14286 (N_14286,N_10958,N_10451);
nor U14287 (N_14287,N_11256,N_10175);
nor U14288 (N_14288,N_9657,N_9871);
nor U14289 (N_14289,N_9603,N_11359);
nand U14290 (N_14290,N_9645,N_10690);
and U14291 (N_14291,N_9746,N_11436);
and U14292 (N_14292,N_11722,N_10607);
xor U14293 (N_14293,N_11467,N_11493);
xnor U14294 (N_14294,N_9119,N_11771);
nand U14295 (N_14295,N_9657,N_11635);
nor U14296 (N_14296,N_11881,N_10432);
and U14297 (N_14297,N_9170,N_10766);
nor U14298 (N_14298,N_11861,N_11929);
and U14299 (N_14299,N_11965,N_11990);
nor U14300 (N_14300,N_11824,N_10353);
nand U14301 (N_14301,N_9492,N_11319);
or U14302 (N_14302,N_10509,N_11224);
or U14303 (N_14303,N_9871,N_10482);
nor U14304 (N_14304,N_10426,N_10550);
and U14305 (N_14305,N_11113,N_9935);
or U14306 (N_14306,N_10694,N_10917);
or U14307 (N_14307,N_9863,N_9578);
or U14308 (N_14308,N_9086,N_9798);
nand U14309 (N_14309,N_9742,N_9723);
xnor U14310 (N_14310,N_10328,N_11699);
and U14311 (N_14311,N_9745,N_9049);
nor U14312 (N_14312,N_9069,N_11065);
nand U14313 (N_14313,N_10374,N_11489);
nor U14314 (N_14314,N_11371,N_11817);
xnor U14315 (N_14315,N_11124,N_9465);
xor U14316 (N_14316,N_11626,N_10014);
nor U14317 (N_14317,N_10751,N_11576);
or U14318 (N_14318,N_9907,N_11897);
and U14319 (N_14319,N_11735,N_10520);
or U14320 (N_14320,N_9564,N_11648);
xor U14321 (N_14321,N_10622,N_11520);
or U14322 (N_14322,N_11515,N_9752);
xnor U14323 (N_14323,N_9616,N_11294);
nand U14324 (N_14324,N_9731,N_11015);
or U14325 (N_14325,N_9951,N_11291);
xnor U14326 (N_14326,N_9179,N_11985);
nor U14327 (N_14327,N_9863,N_10224);
nand U14328 (N_14328,N_10330,N_9974);
nor U14329 (N_14329,N_9591,N_10076);
nand U14330 (N_14330,N_9923,N_9461);
and U14331 (N_14331,N_11371,N_11483);
and U14332 (N_14332,N_11483,N_11014);
xor U14333 (N_14333,N_9574,N_9908);
xor U14334 (N_14334,N_11750,N_9897);
nor U14335 (N_14335,N_10084,N_10533);
or U14336 (N_14336,N_9072,N_11332);
xnor U14337 (N_14337,N_11326,N_10388);
nand U14338 (N_14338,N_9086,N_10168);
and U14339 (N_14339,N_9675,N_10630);
nand U14340 (N_14340,N_10377,N_11625);
xnor U14341 (N_14341,N_9156,N_11554);
and U14342 (N_14342,N_10999,N_10143);
xnor U14343 (N_14343,N_11725,N_10649);
nor U14344 (N_14344,N_10460,N_11434);
and U14345 (N_14345,N_9353,N_10149);
nand U14346 (N_14346,N_11180,N_9451);
or U14347 (N_14347,N_10032,N_9778);
or U14348 (N_14348,N_11893,N_11638);
nand U14349 (N_14349,N_11821,N_9586);
nand U14350 (N_14350,N_9660,N_9152);
nor U14351 (N_14351,N_10123,N_10212);
and U14352 (N_14352,N_10105,N_11472);
nand U14353 (N_14353,N_10217,N_10329);
nor U14354 (N_14354,N_11560,N_9912);
and U14355 (N_14355,N_9594,N_9214);
or U14356 (N_14356,N_10512,N_10419);
or U14357 (N_14357,N_9655,N_11575);
xnor U14358 (N_14358,N_10407,N_10618);
xor U14359 (N_14359,N_10070,N_10768);
nand U14360 (N_14360,N_10152,N_10584);
nand U14361 (N_14361,N_10439,N_9066);
xor U14362 (N_14362,N_9137,N_9360);
xor U14363 (N_14363,N_11696,N_9491);
nand U14364 (N_14364,N_10000,N_11866);
and U14365 (N_14365,N_10659,N_10009);
or U14366 (N_14366,N_10731,N_9731);
nand U14367 (N_14367,N_10614,N_10087);
nand U14368 (N_14368,N_9953,N_11442);
xnor U14369 (N_14369,N_9479,N_11462);
or U14370 (N_14370,N_10986,N_9792);
nor U14371 (N_14371,N_11210,N_11195);
nor U14372 (N_14372,N_11738,N_10717);
and U14373 (N_14373,N_11906,N_9325);
nor U14374 (N_14374,N_9313,N_10368);
and U14375 (N_14375,N_9076,N_11919);
xor U14376 (N_14376,N_9475,N_9327);
nor U14377 (N_14377,N_9945,N_10543);
or U14378 (N_14378,N_9295,N_10465);
and U14379 (N_14379,N_11402,N_10497);
xor U14380 (N_14380,N_9506,N_10284);
nor U14381 (N_14381,N_11151,N_9063);
and U14382 (N_14382,N_9687,N_10172);
nand U14383 (N_14383,N_11957,N_10452);
nor U14384 (N_14384,N_11684,N_10549);
and U14385 (N_14385,N_9726,N_11156);
nor U14386 (N_14386,N_11165,N_11220);
nand U14387 (N_14387,N_10801,N_10976);
xor U14388 (N_14388,N_9778,N_10097);
and U14389 (N_14389,N_9792,N_9676);
or U14390 (N_14390,N_10955,N_10232);
or U14391 (N_14391,N_11310,N_11832);
nor U14392 (N_14392,N_9887,N_9415);
or U14393 (N_14393,N_10151,N_11017);
and U14394 (N_14394,N_9437,N_9156);
xor U14395 (N_14395,N_11246,N_9409);
or U14396 (N_14396,N_11680,N_10461);
xor U14397 (N_14397,N_9510,N_11523);
or U14398 (N_14398,N_11168,N_11176);
xnor U14399 (N_14399,N_9069,N_11583);
xnor U14400 (N_14400,N_9330,N_11480);
xor U14401 (N_14401,N_10336,N_9437);
nand U14402 (N_14402,N_10060,N_9510);
xor U14403 (N_14403,N_9291,N_11186);
xnor U14404 (N_14404,N_9835,N_11357);
or U14405 (N_14405,N_11696,N_10624);
nand U14406 (N_14406,N_11593,N_9168);
xor U14407 (N_14407,N_10626,N_9825);
xnor U14408 (N_14408,N_9801,N_9260);
nor U14409 (N_14409,N_10869,N_11845);
and U14410 (N_14410,N_9273,N_10551);
or U14411 (N_14411,N_11117,N_9146);
nand U14412 (N_14412,N_10961,N_9455);
nand U14413 (N_14413,N_10371,N_9987);
xor U14414 (N_14414,N_9213,N_9263);
and U14415 (N_14415,N_10957,N_11053);
or U14416 (N_14416,N_9789,N_9777);
or U14417 (N_14417,N_9748,N_10004);
or U14418 (N_14418,N_11595,N_9410);
and U14419 (N_14419,N_10249,N_11682);
or U14420 (N_14420,N_9980,N_10826);
or U14421 (N_14421,N_11329,N_11395);
nand U14422 (N_14422,N_10425,N_10383);
or U14423 (N_14423,N_11264,N_11505);
or U14424 (N_14424,N_11720,N_10764);
and U14425 (N_14425,N_11588,N_10816);
nand U14426 (N_14426,N_9244,N_9836);
and U14427 (N_14427,N_10416,N_10290);
and U14428 (N_14428,N_9525,N_11665);
or U14429 (N_14429,N_9011,N_11421);
and U14430 (N_14430,N_10807,N_9035);
nor U14431 (N_14431,N_10972,N_11280);
and U14432 (N_14432,N_11082,N_9876);
nand U14433 (N_14433,N_11180,N_10428);
nor U14434 (N_14434,N_10669,N_9706);
nor U14435 (N_14435,N_10814,N_11529);
nand U14436 (N_14436,N_10441,N_9171);
or U14437 (N_14437,N_9754,N_9743);
nor U14438 (N_14438,N_9627,N_9264);
and U14439 (N_14439,N_11598,N_9718);
and U14440 (N_14440,N_10072,N_10859);
nor U14441 (N_14441,N_9974,N_9348);
nor U14442 (N_14442,N_11988,N_10527);
or U14443 (N_14443,N_9146,N_9434);
nor U14444 (N_14444,N_11502,N_11990);
and U14445 (N_14445,N_9774,N_11620);
nand U14446 (N_14446,N_10941,N_11405);
and U14447 (N_14447,N_10740,N_11088);
or U14448 (N_14448,N_9719,N_11750);
xor U14449 (N_14449,N_11366,N_11394);
xnor U14450 (N_14450,N_11437,N_10158);
nand U14451 (N_14451,N_9886,N_10395);
nor U14452 (N_14452,N_10401,N_10939);
or U14453 (N_14453,N_11772,N_10087);
xor U14454 (N_14454,N_9746,N_10650);
nor U14455 (N_14455,N_11546,N_10571);
nand U14456 (N_14456,N_10326,N_11614);
nor U14457 (N_14457,N_9619,N_11090);
and U14458 (N_14458,N_11605,N_11586);
or U14459 (N_14459,N_10703,N_9391);
nor U14460 (N_14460,N_9608,N_10951);
xor U14461 (N_14461,N_9607,N_10146);
and U14462 (N_14462,N_10401,N_11632);
xor U14463 (N_14463,N_9054,N_9841);
nor U14464 (N_14464,N_11640,N_10931);
nor U14465 (N_14465,N_11197,N_10401);
and U14466 (N_14466,N_10752,N_9904);
or U14467 (N_14467,N_11792,N_10950);
and U14468 (N_14468,N_10010,N_9160);
or U14469 (N_14469,N_11405,N_11489);
nor U14470 (N_14470,N_9931,N_11649);
nor U14471 (N_14471,N_9069,N_10771);
nand U14472 (N_14472,N_11391,N_10135);
and U14473 (N_14473,N_9897,N_11929);
nand U14474 (N_14474,N_11123,N_9820);
nand U14475 (N_14475,N_10948,N_10229);
nor U14476 (N_14476,N_11912,N_9408);
nand U14477 (N_14477,N_11385,N_9743);
nor U14478 (N_14478,N_11587,N_11738);
or U14479 (N_14479,N_9835,N_11818);
nand U14480 (N_14480,N_10990,N_10179);
nor U14481 (N_14481,N_11874,N_11812);
nand U14482 (N_14482,N_9868,N_10270);
nand U14483 (N_14483,N_10888,N_10617);
nor U14484 (N_14484,N_9543,N_10876);
and U14485 (N_14485,N_10543,N_10892);
xnor U14486 (N_14486,N_10644,N_11367);
xor U14487 (N_14487,N_9454,N_10122);
nor U14488 (N_14488,N_11067,N_9511);
or U14489 (N_14489,N_9188,N_11701);
nor U14490 (N_14490,N_9801,N_9455);
xor U14491 (N_14491,N_11133,N_11331);
nor U14492 (N_14492,N_9732,N_9147);
or U14493 (N_14493,N_9381,N_10227);
and U14494 (N_14494,N_10026,N_9846);
nand U14495 (N_14495,N_9270,N_11144);
or U14496 (N_14496,N_11927,N_10627);
nor U14497 (N_14497,N_9977,N_10882);
and U14498 (N_14498,N_9539,N_11123);
or U14499 (N_14499,N_9704,N_11521);
and U14500 (N_14500,N_11777,N_9226);
nand U14501 (N_14501,N_10550,N_11842);
or U14502 (N_14502,N_10712,N_10525);
or U14503 (N_14503,N_10511,N_9619);
xnor U14504 (N_14504,N_9186,N_9325);
or U14505 (N_14505,N_9139,N_11306);
nor U14506 (N_14506,N_9058,N_9414);
xor U14507 (N_14507,N_9277,N_9971);
nand U14508 (N_14508,N_10496,N_10223);
xnor U14509 (N_14509,N_11694,N_9256);
nor U14510 (N_14510,N_9177,N_11015);
nor U14511 (N_14511,N_9840,N_11249);
nor U14512 (N_14512,N_10987,N_10640);
nand U14513 (N_14513,N_11027,N_10882);
or U14514 (N_14514,N_11745,N_10701);
nand U14515 (N_14515,N_10880,N_11542);
and U14516 (N_14516,N_9402,N_10848);
and U14517 (N_14517,N_10665,N_10384);
nor U14518 (N_14518,N_10303,N_9981);
xor U14519 (N_14519,N_11512,N_10986);
or U14520 (N_14520,N_11931,N_11889);
and U14521 (N_14521,N_11932,N_9850);
nand U14522 (N_14522,N_9501,N_11416);
xnor U14523 (N_14523,N_11983,N_11702);
and U14524 (N_14524,N_11261,N_10866);
or U14525 (N_14525,N_9442,N_10107);
or U14526 (N_14526,N_10246,N_10893);
and U14527 (N_14527,N_11505,N_10702);
nand U14528 (N_14528,N_10616,N_11762);
nand U14529 (N_14529,N_11992,N_9954);
nor U14530 (N_14530,N_9625,N_11276);
and U14531 (N_14531,N_11650,N_10213);
nand U14532 (N_14532,N_11182,N_11441);
nor U14533 (N_14533,N_9422,N_10014);
nor U14534 (N_14534,N_11949,N_9866);
and U14535 (N_14535,N_9155,N_9521);
and U14536 (N_14536,N_9404,N_10641);
nor U14537 (N_14537,N_9564,N_10829);
and U14538 (N_14538,N_10047,N_11710);
nor U14539 (N_14539,N_9095,N_9663);
xor U14540 (N_14540,N_9537,N_9528);
or U14541 (N_14541,N_10688,N_11506);
nor U14542 (N_14542,N_10239,N_11492);
and U14543 (N_14543,N_10962,N_10884);
xnor U14544 (N_14544,N_11931,N_11985);
or U14545 (N_14545,N_10130,N_11275);
nor U14546 (N_14546,N_10587,N_10066);
xnor U14547 (N_14547,N_11874,N_9513);
and U14548 (N_14548,N_10334,N_10805);
xnor U14549 (N_14549,N_9341,N_11081);
nand U14550 (N_14550,N_11761,N_10592);
xor U14551 (N_14551,N_11807,N_11279);
nand U14552 (N_14552,N_10007,N_11126);
nor U14553 (N_14553,N_9642,N_9533);
nor U14554 (N_14554,N_10367,N_9597);
nand U14555 (N_14555,N_10588,N_9885);
nand U14556 (N_14556,N_11927,N_9851);
xor U14557 (N_14557,N_9465,N_10672);
and U14558 (N_14558,N_9180,N_9634);
nor U14559 (N_14559,N_9445,N_9367);
or U14560 (N_14560,N_11807,N_11539);
xor U14561 (N_14561,N_11631,N_10879);
nor U14562 (N_14562,N_10174,N_11568);
or U14563 (N_14563,N_10308,N_9912);
or U14564 (N_14564,N_9254,N_10137);
and U14565 (N_14565,N_11802,N_10590);
or U14566 (N_14566,N_9781,N_11584);
xnor U14567 (N_14567,N_9074,N_11310);
nor U14568 (N_14568,N_10017,N_11762);
and U14569 (N_14569,N_9176,N_9053);
nand U14570 (N_14570,N_10019,N_9001);
nand U14571 (N_14571,N_10559,N_9552);
nand U14572 (N_14572,N_11286,N_11067);
or U14573 (N_14573,N_10878,N_10072);
xnor U14574 (N_14574,N_11846,N_11311);
xor U14575 (N_14575,N_10325,N_11290);
nand U14576 (N_14576,N_10967,N_10475);
nand U14577 (N_14577,N_11633,N_9202);
and U14578 (N_14578,N_9179,N_11085);
nor U14579 (N_14579,N_10022,N_10651);
nand U14580 (N_14580,N_10504,N_10312);
and U14581 (N_14581,N_11480,N_9456);
and U14582 (N_14582,N_9108,N_9078);
nand U14583 (N_14583,N_11673,N_9524);
or U14584 (N_14584,N_10158,N_9055);
xor U14585 (N_14585,N_11942,N_10469);
xnor U14586 (N_14586,N_10062,N_9793);
nand U14587 (N_14587,N_10966,N_10729);
nor U14588 (N_14588,N_9890,N_9886);
or U14589 (N_14589,N_9221,N_10457);
xor U14590 (N_14590,N_10195,N_9416);
or U14591 (N_14591,N_9012,N_11390);
nor U14592 (N_14592,N_10159,N_10823);
or U14593 (N_14593,N_10988,N_10372);
or U14594 (N_14594,N_9767,N_11720);
and U14595 (N_14595,N_10114,N_9483);
nor U14596 (N_14596,N_10028,N_11469);
xor U14597 (N_14597,N_9449,N_9839);
and U14598 (N_14598,N_11263,N_11411);
or U14599 (N_14599,N_11313,N_10866);
xnor U14600 (N_14600,N_9710,N_9156);
or U14601 (N_14601,N_9954,N_10764);
xnor U14602 (N_14602,N_9805,N_10503);
nand U14603 (N_14603,N_11032,N_9104);
nor U14604 (N_14604,N_9873,N_10141);
nand U14605 (N_14605,N_10741,N_10830);
and U14606 (N_14606,N_9691,N_9260);
and U14607 (N_14607,N_10597,N_11835);
or U14608 (N_14608,N_10351,N_10089);
or U14609 (N_14609,N_11560,N_10048);
and U14610 (N_14610,N_11256,N_11899);
xor U14611 (N_14611,N_9411,N_10227);
nand U14612 (N_14612,N_9451,N_11161);
xnor U14613 (N_14613,N_9997,N_10322);
nand U14614 (N_14614,N_9478,N_9439);
xnor U14615 (N_14615,N_9123,N_9047);
xor U14616 (N_14616,N_9090,N_10886);
or U14617 (N_14617,N_11357,N_11970);
xnor U14618 (N_14618,N_9311,N_10430);
xor U14619 (N_14619,N_10415,N_10261);
or U14620 (N_14620,N_10434,N_9130);
or U14621 (N_14621,N_9053,N_11456);
nor U14622 (N_14622,N_10338,N_9585);
and U14623 (N_14623,N_10215,N_10572);
or U14624 (N_14624,N_9146,N_9801);
nor U14625 (N_14625,N_10061,N_11156);
xnor U14626 (N_14626,N_10547,N_10588);
nand U14627 (N_14627,N_11414,N_9291);
nand U14628 (N_14628,N_9565,N_9183);
nor U14629 (N_14629,N_9551,N_11099);
nand U14630 (N_14630,N_9864,N_10177);
xnor U14631 (N_14631,N_10241,N_9013);
nand U14632 (N_14632,N_10657,N_11467);
and U14633 (N_14633,N_10745,N_11485);
nand U14634 (N_14634,N_11103,N_10102);
or U14635 (N_14635,N_11590,N_11846);
nand U14636 (N_14636,N_10865,N_9337);
xor U14637 (N_14637,N_11279,N_11549);
xor U14638 (N_14638,N_10834,N_10039);
and U14639 (N_14639,N_9816,N_11693);
nand U14640 (N_14640,N_9196,N_11740);
xnor U14641 (N_14641,N_9233,N_11277);
nand U14642 (N_14642,N_9878,N_10015);
xnor U14643 (N_14643,N_9998,N_11998);
xor U14644 (N_14644,N_10272,N_9553);
nor U14645 (N_14645,N_11716,N_9709);
or U14646 (N_14646,N_11367,N_9381);
nand U14647 (N_14647,N_11117,N_11856);
nand U14648 (N_14648,N_11204,N_11436);
nand U14649 (N_14649,N_11531,N_11161);
nand U14650 (N_14650,N_9381,N_9649);
xor U14651 (N_14651,N_10641,N_11472);
nor U14652 (N_14652,N_9405,N_9787);
or U14653 (N_14653,N_9338,N_9461);
nand U14654 (N_14654,N_11544,N_9764);
or U14655 (N_14655,N_10192,N_11253);
and U14656 (N_14656,N_9236,N_9253);
nand U14657 (N_14657,N_10781,N_11503);
nor U14658 (N_14658,N_11360,N_10184);
or U14659 (N_14659,N_11857,N_11503);
nand U14660 (N_14660,N_11785,N_10085);
nor U14661 (N_14661,N_10151,N_11391);
xnor U14662 (N_14662,N_11763,N_10759);
or U14663 (N_14663,N_9553,N_9172);
nand U14664 (N_14664,N_10795,N_10366);
or U14665 (N_14665,N_9331,N_10535);
or U14666 (N_14666,N_9818,N_10222);
nand U14667 (N_14667,N_9214,N_10005);
nand U14668 (N_14668,N_10997,N_9766);
nand U14669 (N_14669,N_11642,N_9858);
nor U14670 (N_14670,N_9119,N_11180);
and U14671 (N_14671,N_10836,N_10621);
and U14672 (N_14672,N_11118,N_10986);
or U14673 (N_14673,N_11481,N_9226);
or U14674 (N_14674,N_10275,N_9653);
and U14675 (N_14675,N_11102,N_10264);
xnor U14676 (N_14676,N_9148,N_10082);
xor U14677 (N_14677,N_9605,N_10859);
nand U14678 (N_14678,N_10384,N_11729);
or U14679 (N_14679,N_11531,N_11484);
nor U14680 (N_14680,N_9764,N_10604);
nand U14681 (N_14681,N_9435,N_10503);
xnor U14682 (N_14682,N_9338,N_11648);
xor U14683 (N_14683,N_10049,N_11461);
xnor U14684 (N_14684,N_9706,N_9259);
nor U14685 (N_14685,N_11678,N_10020);
nand U14686 (N_14686,N_10667,N_9198);
or U14687 (N_14687,N_11091,N_9850);
nor U14688 (N_14688,N_9375,N_10360);
and U14689 (N_14689,N_9118,N_11623);
nand U14690 (N_14690,N_11222,N_9860);
nand U14691 (N_14691,N_10732,N_10992);
or U14692 (N_14692,N_11198,N_9346);
nand U14693 (N_14693,N_9848,N_9348);
nand U14694 (N_14694,N_10429,N_11569);
or U14695 (N_14695,N_11341,N_10625);
nor U14696 (N_14696,N_11188,N_11192);
or U14697 (N_14697,N_9093,N_9529);
nor U14698 (N_14698,N_9578,N_9126);
xnor U14699 (N_14699,N_10764,N_9460);
and U14700 (N_14700,N_9993,N_9896);
nor U14701 (N_14701,N_9113,N_10192);
nand U14702 (N_14702,N_10889,N_11514);
or U14703 (N_14703,N_9546,N_11011);
nand U14704 (N_14704,N_9891,N_10813);
or U14705 (N_14705,N_10400,N_10192);
and U14706 (N_14706,N_10665,N_10188);
xnor U14707 (N_14707,N_11076,N_9364);
or U14708 (N_14708,N_11889,N_11145);
and U14709 (N_14709,N_10076,N_9755);
and U14710 (N_14710,N_9993,N_9337);
or U14711 (N_14711,N_11912,N_11692);
and U14712 (N_14712,N_9785,N_11953);
or U14713 (N_14713,N_9189,N_11667);
and U14714 (N_14714,N_9971,N_10958);
and U14715 (N_14715,N_9069,N_10618);
and U14716 (N_14716,N_9134,N_10858);
xnor U14717 (N_14717,N_10670,N_11920);
nand U14718 (N_14718,N_10642,N_11304);
and U14719 (N_14719,N_10975,N_11081);
or U14720 (N_14720,N_10993,N_11771);
nor U14721 (N_14721,N_9781,N_9690);
or U14722 (N_14722,N_11673,N_11593);
nand U14723 (N_14723,N_9819,N_10885);
nand U14724 (N_14724,N_10510,N_11030);
nand U14725 (N_14725,N_10313,N_10327);
xnor U14726 (N_14726,N_10295,N_9891);
nor U14727 (N_14727,N_10885,N_11990);
xnor U14728 (N_14728,N_10718,N_9963);
xor U14729 (N_14729,N_10074,N_9163);
and U14730 (N_14730,N_11226,N_11535);
and U14731 (N_14731,N_10952,N_10909);
or U14732 (N_14732,N_11357,N_9792);
or U14733 (N_14733,N_11247,N_10025);
nor U14734 (N_14734,N_9385,N_11836);
or U14735 (N_14735,N_9808,N_11188);
xnor U14736 (N_14736,N_9131,N_10474);
nand U14737 (N_14737,N_9374,N_11436);
xor U14738 (N_14738,N_9448,N_9591);
or U14739 (N_14739,N_10575,N_10988);
nor U14740 (N_14740,N_10835,N_9995);
nor U14741 (N_14741,N_9225,N_9202);
nor U14742 (N_14742,N_10364,N_9032);
nand U14743 (N_14743,N_10671,N_9969);
nor U14744 (N_14744,N_9241,N_9158);
nand U14745 (N_14745,N_9907,N_9035);
and U14746 (N_14746,N_9775,N_10286);
and U14747 (N_14747,N_11925,N_11906);
or U14748 (N_14748,N_11290,N_10056);
xor U14749 (N_14749,N_10849,N_10578);
and U14750 (N_14750,N_9720,N_11493);
and U14751 (N_14751,N_11378,N_11088);
nand U14752 (N_14752,N_11200,N_9315);
xnor U14753 (N_14753,N_11127,N_10160);
xnor U14754 (N_14754,N_11284,N_9420);
or U14755 (N_14755,N_10590,N_11344);
xnor U14756 (N_14756,N_10441,N_11063);
nand U14757 (N_14757,N_10111,N_10766);
nor U14758 (N_14758,N_9229,N_9676);
or U14759 (N_14759,N_11887,N_11368);
and U14760 (N_14760,N_11314,N_11633);
or U14761 (N_14761,N_11917,N_9952);
nand U14762 (N_14762,N_11001,N_11921);
nor U14763 (N_14763,N_10671,N_10442);
nor U14764 (N_14764,N_11473,N_9802);
and U14765 (N_14765,N_9404,N_9519);
xor U14766 (N_14766,N_11531,N_11481);
and U14767 (N_14767,N_9206,N_10136);
nand U14768 (N_14768,N_9377,N_9554);
nor U14769 (N_14769,N_10321,N_10275);
nor U14770 (N_14770,N_11508,N_9041);
or U14771 (N_14771,N_10866,N_10108);
nor U14772 (N_14772,N_11147,N_10067);
nor U14773 (N_14773,N_9996,N_10500);
nand U14774 (N_14774,N_9744,N_11891);
or U14775 (N_14775,N_11081,N_11870);
xor U14776 (N_14776,N_11750,N_9507);
and U14777 (N_14777,N_9825,N_10829);
or U14778 (N_14778,N_10684,N_11450);
xnor U14779 (N_14779,N_11009,N_10575);
nand U14780 (N_14780,N_9048,N_10304);
nor U14781 (N_14781,N_9099,N_10400);
and U14782 (N_14782,N_9719,N_10078);
nor U14783 (N_14783,N_11085,N_10875);
and U14784 (N_14784,N_9755,N_9427);
nor U14785 (N_14785,N_11867,N_9449);
nand U14786 (N_14786,N_9423,N_10161);
nor U14787 (N_14787,N_9731,N_11706);
nor U14788 (N_14788,N_9130,N_11026);
or U14789 (N_14789,N_9848,N_10759);
or U14790 (N_14790,N_11633,N_11351);
and U14791 (N_14791,N_11847,N_10625);
xor U14792 (N_14792,N_11968,N_11330);
xnor U14793 (N_14793,N_11710,N_10839);
nand U14794 (N_14794,N_11509,N_9763);
or U14795 (N_14795,N_11039,N_10686);
xor U14796 (N_14796,N_9342,N_10666);
and U14797 (N_14797,N_11697,N_11148);
and U14798 (N_14798,N_9677,N_10052);
xnor U14799 (N_14799,N_11783,N_9750);
nand U14800 (N_14800,N_11464,N_10847);
xnor U14801 (N_14801,N_11980,N_10661);
or U14802 (N_14802,N_11048,N_11533);
nand U14803 (N_14803,N_10417,N_9389);
xnor U14804 (N_14804,N_11418,N_11586);
and U14805 (N_14805,N_9609,N_11391);
and U14806 (N_14806,N_9520,N_9174);
xor U14807 (N_14807,N_11168,N_10330);
nand U14808 (N_14808,N_9230,N_10902);
nand U14809 (N_14809,N_11772,N_10786);
nand U14810 (N_14810,N_10405,N_10403);
xor U14811 (N_14811,N_9473,N_10185);
nand U14812 (N_14812,N_10648,N_11337);
xor U14813 (N_14813,N_11965,N_11259);
nand U14814 (N_14814,N_11949,N_10845);
and U14815 (N_14815,N_11690,N_10839);
nand U14816 (N_14816,N_11039,N_9771);
nand U14817 (N_14817,N_9638,N_10504);
nor U14818 (N_14818,N_11417,N_9148);
nor U14819 (N_14819,N_10901,N_9482);
nand U14820 (N_14820,N_9451,N_11199);
and U14821 (N_14821,N_11120,N_11515);
and U14822 (N_14822,N_11140,N_11046);
and U14823 (N_14823,N_10073,N_10728);
nand U14824 (N_14824,N_11021,N_11259);
or U14825 (N_14825,N_11286,N_11908);
and U14826 (N_14826,N_11806,N_11116);
nor U14827 (N_14827,N_9842,N_10025);
xnor U14828 (N_14828,N_10149,N_10746);
nand U14829 (N_14829,N_11264,N_11318);
nand U14830 (N_14830,N_9290,N_10662);
nand U14831 (N_14831,N_10211,N_9895);
nor U14832 (N_14832,N_9435,N_9694);
xor U14833 (N_14833,N_11802,N_10924);
nand U14834 (N_14834,N_11711,N_9573);
nand U14835 (N_14835,N_11612,N_10326);
and U14836 (N_14836,N_10801,N_9422);
or U14837 (N_14837,N_10163,N_9428);
nor U14838 (N_14838,N_11706,N_11769);
or U14839 (N_14839,N_10252,N_11536);
and U14840 (N_14840,N_9858,N_9058);
nand U14841 (N_14841,N_9581,N_11627);
nor U14842 (N_14842,N_11224,N_10170);
nor U14843 (N_14843,N_10191,N_10775);
or U14844 (N_14844,N_11307,N_11252);
or U14845 (N_14845,N_9053,N_9788);
xnor U14846 (N_14846,N_11195,N_10937);
or U14847 (N_14847,N_9831,N_10424);
nor U14848 (N_14848,N_10616,N_10458);
xor U14849 (N_14849,N_9306,N_9414);
and U14850 (N_14850,N_10041,N_10984);
nand U14851 (N_14851,N_9384,N_9638);
nor U14852 (N_14852,N_10238,N_11990);
nor U14853 (N_14853,N_11470,N_10528);
nand U14854 (N_14854,N_9291,N_9207);
nand U14855 (N_14855,N_10742,N_10854);
and U14856 (N_14856,N_10639,N_9069);
nand U14857 (N_14857,N_9706,N_9688);
nor U14858 (N_14858,N_10869,N_11807);
nor U14859 (N_14859,N_9753,N_9412);
and U14860 (N_14860,N_11379,N_10781);
and U14861 (N_14861,N_10885,N_11649);
nand U14862 (N_14862,N_10817,N_11023);
and U14863 (N_14863,N_10495,N_10440);
nor U14864 (N_14864,N_11701,N_11662);
nand U14865 (N_14865,N_10296,N_10707);
and U14866 (N_14866,N_10455,N_11121);
nor U14867 (N_14867,N_11070,N_9892);
nor U14868 (N_14868,N_10287,N_9524);
nand U14869 (N_14869,N_9696,N_10785);
or U14870 (N_14870,N_11012,N_11963);
nor U14871 (N_14871,N_9966,N_10784);
xnor U14872 (N_14872,N_9829,N_10908);
xnor U14873 (N_14873,N_9840,N_9142);
nand U14874 (N_14874,N_11842,N_9596);
nor U14875 (N_14875,N_9492,N_9569);
and U14876 (N_14876,N_10838,N_11789);
and U14877 (N_14877,N_11486,N_11858);
nor U14878 (N_14878,N_9221,N_10384);
xnor U14879 (N_14879,N_10848,N_10139);
nor U14880 (N_14880,N_10426,N_10918);
nand U14881 (N_14881,N_11986,N_11716);
and U14882 (N_14882,N_9564,N_10544);
xor U14883 (N_14883,N_10154,N_11146);
nor U14884 (N_14884,N_9715,N_9815);
nor U14885 (N_14885,N_11837,N_11029);
nor U14886 (N_14886,N_11028,N_9791);
and U14887 (N_14887,N_10688,N_11128);
nand U14888 (N_14888,N_10959,N_11673);
xnor U14889 (N_14889,N_11434,N_10187);
nand U14890 (N_14890,N_11538,N_11279);
nand U14891 (N_14891,N_10762,N_9984);
nor U14892 (N_14892,N_10043,N_9621);
nand U14893 (N_14893,N_9517,N_10926);
nor U14894 (N_14894,N_9255,N_11261);
nor U14895 (N_14895,N_10241,N_9670);
xnor U14896 (N_14896,N_9775,N_10284);
nand U14897 (N_14897,N_11240,N_9695);
and U14898 (N_14898,N_11753,N_9029);
or U14899 (N_14899,N_10000,N_10608);
or U14900 (N_14900,N_9960,N_10528);
nand U14901 (N_14901,N_10414,N_10884);
or U14902 (N_14902,N_11850,N_10321);
xor U14903 (N_14903,N_9900,N_10446);
xor U14904 (N_14904,N_9999,N_10104);
nor U14905 (N_14905,N_11436,N_9361);
xnor U14906 (N_14906,N_11876,N_10360);
xnor U14907 (N_14907,N_9693,N_9394);
nor U14908 (N_14908,N_10037,N_10802);
and U14909 (N_14909,N_11892,N_11899);
or U14910 (N_14910,N_10107,N_10831);
nor U14911 (N_14911,N_10662,N_10285);
nor U14912 (N_14912,N_11595,N_9247);
nand U14913 (N_14913,N_9847,N_9027);
and U14914 (N_14914,N_10822,N_11744);
nor U14915 (N_14915,N_9393,N_11983);
or U14916 (N_14916,N_11699,N_9030);
xor U14917 (N_14917,N_11602,N_9177);
nor U14918 (N_14918,N_10497,N_10323);
and U14919 (N_14919,N_9953,N_11907);
and U14920 (N_14920,N_9686,N_11932);
or U14921 (N_14921,N_9490,N_11462);
xnor U14922 (N_14922,N_11677,N_10515);
or U14923 (N_14923,N_11842,N_10972);
xor U14924 (N_14924,N_10494,N_10673);
and U14925 (N_14925,N_9809,N_10184);
and U14926 (N_14926,N_10706,N_11135);
or U14927 (N_14927,N_10658,N_9396);
nor U14928 (N_14928,N_9511,N_9268);
or U14929 (N_14929,N_10784,N_11394);
nor U14930 (N_14930,N_10376,N_10544);
and U14931 (N_14931,N_11839,N_9522);
or U14932 (N_14932,N_9978,N_10700);
and U14933 (N_14933,N_10187,N_11207);
and U14934 (N_14934,N_11950,N_11990);
nand U14935 (N_14935,N_11165,N_9148);
nor U14936 (N_14936,N_10759,N_11329);
and U14937 (N_14937,N_9121,N_10060);
xor U14938 (N_14938,N_11763,N_9224);
nand U14939 (N_14939,N_10080,N_9916);
nor U14940 (N_14940,N_10205,N_9912);
xor U14941 (N_14941,N_10235,N_11088);
nor U14942 (N_14942,N_10956,N_9701);
and U14943 (N_14943,N_10373,N_10225);
nand U14944 (N_14944,N_11384,N_10325);
or U14945 (N_14945,N_10961,N_9245);
xor U14946 (N_14946,N_11045,N_10700);
xnor U14947 (N_14947,N_9163,N_9045);
nor U14948 (N_14948,N_10757,N_10338);
and U14949 (N_14949,N_11079,N_11168);
and U14950 (N_14950,N_11434,N_11351);
xnor U14951 (N_14951,N_11303,N_11928);
xnor U14952 (N_14952,N_9032,N_11930);
or U14953 (N_14953,N_9492,N_9371);
xnor U14954 (N_14954,N_9014,N_11075);
and U14955 (N_14955,N_10047,N_10336);
nor U14956 (N_14956,N_10407,N_9596);
nand U14957 (N_14957,N_10596,N_9519);
or U14958 (N_14958,N_10633,N_10077);
and U14959 (N_14959,N_10664,N_11366);
nand U14960 (N_14960,N_10601,N_11035);
and U14961 (N_14961,N_11521,N_9654);
xor U14962 (N_14962,N_10687,N_9656);
and U14963 (N_14963,N_11592,N_11850);
and U14964 (N_14964,N_9397,N_9860);
or U14965 (N_14965,N_10820,N_11532);
and U14966 (N_14966,N_9540,N_11449);
nand U14967 (N_14967,N_9610,N_9248);
or U14968 (N_14968,N_11652,N_10623);
or U14969 (N_14969,N_10687,N_11376);
xor U14970 (N_14970,N_11975,N_11370);
or U14971 (N_14971,N_9753,N_9326);
or U14972 (N_14972,N_10494,N_10028);
and U14973 (N_14973,N_9979,N_9414);
and U14974 (N_14974,N_11934,N_9854);
or U14975 (N_14975,N_10977,N_10888);
or U14976 (N_14976,N_11060,N_11949);
nor U14977 (N_14977,N_9186,N_9020);
and U14978 (N_14978,N_10756,N_11026);
nor U14979 (N_14979,N_10852,N_9726);
xnor U14980 (N_14980,N_10693,N_9551);
nor U14981 (N_14981,N_10624,N_10002);
nand U14982 (N_14982,N_9047,N_10404);
or U14983 (N_14983,N_11919,N_9524);
nor U14984 (N_14984,N_9036,N_11264);
and U14985 (N_14985,N_10083,N_11695);
xnor U14986 (N_14986,N_10621,N_9942);
nor U14987 (N_14987,N_9289,N_10309);
xnor U14988 (N_14988,N_11021,N_11909);
or U14989 (N_14989,N_10471,N_10945);
or U14990 (N_14990,N_9879,N_11702);
and U14991 (N_14991,N_11489,N_11459);
nor U14992 (N_14992,N_10455,N_11058);
or U14993 (N_14993,N_9360,N_10298);
xor U14994 (N_14994,N_11667,N_9330);
nor U14995 (N_14995,N_10561,N_9730);
or U14996 (N_14996,N_9276,N_10930);
nor U14997 (N_14997,N_10529,N_9842);
xnor U14998 (N_14998,N_11044,N_10150);
nor U14999 (N_14999,N_9327,N_10381);
or UO_0 (O_0,N_12904,N_12127);
nand UO_1 (O_1,N_13515,N_12625);
or UO_2 (O_2,N_13319,N_13477);
xor UO_3 (O_3,N_13247,N_13103);
or UO_4 (O_4,N_12209,N_14098);
nand UO_5 (O_5,N_14305,N_13169);
nand UO_6 (O_6,N_14085,N_13969);
nor UO_7 (O_7,N_12293,N_12007);
xor UO_8 (O_8,N_12800,N_13026);
nand UO_9 (O_9,N_13012,N_14042);
or UO_10 (O_10,N_12238,N_13532);
xnor UO_11 (O_11,N_14809,N_13170);
xnor UO_12 (O_12,N_13375,N_13866);
and UO_13 (O_13,N_12867,N_14655);
or UO_14 (O_14,N_12469,N_14377);
xor UO_15 (O_15,N_12754,N_14977);
or UO_16 (O_16,N_12567,N_13140);
xor UO_17 (O_17,N_14472,N_14631);
and UO_18 (O_18,N_12268,N_12724);
or UO_19 (O_19,N_14213,N_13071);
xnor UO_20 (O_20,N_14758,N_13489);
and UO_21 (O_21,N_13225,N_13983);
or UO_22 (O_22,N_13855,N_12711);
nor UO_23 (O_23,N_12964,N_14505);
xor UO_24 (O_24,N_14450,N_13014);
or UO_25 (O_25,N_13464,N_14818);
xnor UO_26 (O_26,N_13807,N_12126);
nor UO_27 (O_27,N_12504,N_12161);
or UO_28 (O_28,N_14076,N_14964);
and UO_29 (O_29,N_14700,N_12100);
nor UO_30 (O_30,N_14326,N_14715);
or UO_31 (O_31,N_14183,N_12651);
xnor UO_32 (O_32,N_14403,N_14469);
nor UO_33 (O_33,N_13896,N_13781);
or UO_34 (O_34,N_12124,N_13978);
and UO_35 (O_35,N_14981,N_13461);
and UO_36 (O_36,N_14506,N_12187);
xor UO_37 (O_37,N_12873,N_12328);
or UO_38 (O_38,N_14238,N_13186);
nand UO_39 (O_39,N_13571,N_13282);
and UO_40 (O_40,N_13151,N_12888);
or UO_41 (O_41,N_14214,N_13490);
and UO_42 (O_42,N_12384,N_14125);
or UO_43 (O_43,N_12700,N_12967);
xor UO_44 (O_44,N_12212,N_13079);
nor UO_45 (O_45,N_13775,N_13637);
nor UO_46 (O_46,N_12620,N_14392);
and UO_47 (O_47,N_14270,N_13408);
nand UO_48 (O_48,N_12676,N_13200);
xor UO_49 (O_49,N_13799,N_14934);
xnor UO_50 (O_50,N_14870,N_13626);
nand UO_51 (O_51,N_13344,N_14113);
xor UO_52 (O_52,N_12222,N_13924);
nand UO_53 (O_53,N_13195,N_14847);
nand UO_54 (O_54,N_13697,N_12242);
nor UO_55 (O_55,N_14976,N_12540);
nor UO_56 (O_56,N_14857,N_12405);
nand UO_57 (O_57,N_12198,N_14293);
nand UO_58 (O_58,N_12740,N_13792);
or UO_59 (O_59,N_13309,N_12284);
and UO_60 (O_60,N_14661,N_13046);
nor UO_61 (O_61,N_13573,N_14146);
nor UO_62 (O_62,N_12677,N_12588);
xnor UO_63 (O_63,N_12152,N_12653);
nor UO_64 (O_64,N_12235,N_13446);
nor UO_65 (O_65,N_12020,N_12704);
and UO_66 (O_66,N_13033,N_12257);
nor UO_67 (O_67,N_14866,N_12546);
nor UO_68 (O_68,N_12299,N_12699);
and UO_69 (O_69,N_13996,N_14625);
or UO_70 (O_70,N_12478,N_13849);
and UO_71 (O_71,N_13735,N_13350);
nand UO_72 (O_72,N_12038,N_14956);
nor UO_73 (O_73,N_13640,N_14320);
nand UO_74 (O_74,N_14583,N_12997);
nor UO_75 (O_75,N_14304,N_14424);
nand UO_76 (O_76,N_13055,N_12370);
nor UO_77 (O_77,N_12428,N_12648);
and UO_78 (O_78,N_12880,N_13514);
nor UO_79 (O_79,N_12534,N_12414);
nand UO_80 (O_80,N_13859,N_14840);
or UO_81 (O_81,N_14679,N_13847);
and UO_82 (O_82,N_13154,N_13812);
nand UO_83 (O_83,N_14779,N_12218);
xnor UO_84 (O_84,N_13441,N_12556);
and UO_85 (O_85,N_14371,N_12348);
or UO_86 (O_86,N_14845,N_14792);
or UO_87 (O_87,N_14582,N_14228);
nand UO_88 (O_88,N_12241,N_13031);
nand UO_89 (O_89,N_13094,N_14930);
or UO_90 (O_90,N_14397,N_14775);
nand UO_91 (O_91,N_14528,N_14493);
nor UO_92 (O_92,N_12833,N_14375);
nand UO_93 (O_93,N_12454,N_13006);
and UO_94 (O_94,N_13434,N_14459);
nand UO_95 (O_95,N_12542,N_13471);
xnor UO_96 (O_96,N_14102,N_13992);
or UO_97 (O_97,N_12615,N_12785);
nor UO_98 (O_98,N_14491,N_14249);
nand UO_99 (O_99,N_13345,N_13882);
nor UO_100 (O_100,N_12176,N_13892);
xor UO_101 (O_101,N_13168,N_13073);
nor UO_102 (O_102,N_13376,N_12025);
or UO_103 (O_103,N_12617,N_13625);
nor UO_104 (O_104,N_12563,N_13361);
nand UO_105 (O_105,N_14226,N_14704);
nor UO_106 (O_106,N_14157,N_14209);
nand UO_107 (O_107,N_13234,N_13582);
nor UO_108 (O_108,N_12995,N_14701);
or UO_109 (O_109,N_14826,N_13653);
and UO_110 (O_110,N_12940,N_14292);
and UO_111 (O_111,N_12452,N_14003);
nand UO_112 (O_112,N_13479,N_12360);
or UO_113 (O_113,N_13262,N_14350);
and UO_114 (O_114,N_13687,N_13960);
and UO_115 (O_115,N_14947,N_14210);
xnor UO_116 (O_116,N_12051,N_12467);
or UO_117 (O_117,N_14634,N_14240);
or UO_118 (O_118,N_13290,N_14475);
and UO_119 (O_119,N_14652,N_13463);
nor UO_120 (O_120,N_12852,N_12426);
xnor UO_121 (O_121,N_12816,N_12164);
xor UO_122 (O_122,N_14605,N_13485);
nor UO_123 (O_123,N_13893,N_14205);
and UO_124 (O_124,N_14300,N_12498);
nor UO_125 (O_125,N_12906,N_14184);
nor UO_126 (O_126,N_13136,N_14974);
nor UO_127 (O_127,N_12443,N_13386);
nor UO_128 (O_128,N_13105,N_13391);
or UO_129 (O_129,N_14055,N_14440);
nor UO_130 (O_130,N_14707,N_13438);
and UO_131 (O_131,N_13809,N_14702);
or UO_132 (O_132,N_12446,N_13482);
nand UO_133 (O_133,N_14781,N_13134);
nand UO_134 (O_134,N_12632,N_13180);
nand UO_135 (O_135,N_12543,N_12207);
or UO_136 (O_136,N_14285,N_12703);
or UO_137 (O_137,N_14031,N_12357);
and UO_138 (O_138,N_12154,N_12600);
nand UO_139 (O_139,N_12231,N_12386);
xnor UO_140 (O_140,N_14991,N_12132);
nand UO_141 (O_141,N_14289,N_13576);
and UO_142 (O_142,N_14369,N_13908);
and UO_143 (O_143,N_14002,N_13585);
or UO_144 (O_144,N_14959,N_13481);
or UO_145 (O_145,N_14393,N_14541);
nor UO_146 (O_146,N_13873,N_14684);
xnor UO_147 (O_147,N_14021,N_14112);
or UO_148 (O_148,N_12914,N_13598);
or UO_149 (O_149,N_12566,N_13927);
xnor UO_150 (O_150,N_13836,N_14729);
nor UO_151 (O_151,N_14982,N_13433);
and UO_152 (O_152,N_12407,N_12297);
nand UO_153 (O_153,N_12728,N_13512);
or UO_154 (O_154,N_12643,N_14429);
or UO_155 (O_155,N_14572,N_13129);
and UO_156 (O_156,N_12385,N_12654);
nor UO_157 (O_157,N_14717,N_12591);
and UO_158 (O_158,N_13374,N_14025);
or UO_159 (O_159,N_14803,N_13534);
or UO_160 (O_160,N_12944,N_12398);
or UO_161 (O_161,N_12850,N_13752);
and UO_162 (O_162,N_14907,N_14576);
nand UO_163 (O_163,N_14137,N_14639);
nor UO_164 (O_164,N_13476,N_12892);
and UO_165 (O_165,N_13586,N_14063);
or UO_166 (O_166,N_14748,N_12551);
nand UO_167 (O_167,N_14175,N_13674);
nor UO_168 (O_168,N_13911,N_14149);
and UO_169 (O_169,N_13043,N_13284);
and UO_170 (O_170,N_13497,N_14227);
or UO_171 (O_171,N_12966,N_12039);
and UO_172 (O_172,N_12349,N_13469);
or UO_173 (O_173,N_14989,N_14136);
nor UO_174 (O_174,N_13861,N_12688);
or UO_175 (O_175,N_12712,N_12952);
xnor UO_176 (O_176,N_13793,N_12974);
xor UO_177 (O_177,N_12623,N_12579);
and UO_178 (O_178,N_12517,N_13891);
nor UO_179 (O_179,N_14372,N_13182);
xnor UO_180 (O_180,N_14396,N_14299);
xnor UO_181 (O_181,N_12658,N_12741);
xnor UO_182 (O_182,N_14246,N_14574);
nand UO_183 (O_183,N_12520,N_13721);
or UO_184 (O_184,N_13047,N_14916);
and UO_185 (O_185,N_12010,N_12810);
and UO_186 (O_186,N_12069,N_14551);
and UO_187 (O_187,N_12784,N_14278);
or UO_188 (O_188,N_12705,N_13985);
nand UO_189 (O_189,N_14894,N_12341);
or UO_190 (O_190,N_13961,N_13541);
nand UO_191 (O_191,N_13679,N_12781);
and UO_192 (O_192,N_12383,N_12709);
or UO_193 (O_193,N_14519,N_12505);
nand UO_194 (O_194,N_13786,N_13106);
and UO_195 (O_195,N_12689,N_12934);
or UO_196 (O_196,N_12539,N_14897);
nand UO_197 (O_197,N_12495,N_14448);
and UO_198 (O_198,N_13691,N_13835);
and UO_199 (O_199,N_13716,N_13628);
or UO_200 (O_200,N_12091,N_12048);
or UO_201 (O_201,N_14562,N_14789);
nand UO_202 (O_202,N_14455,N_14362);
nor UO_203 (O_203,N_14948,N_13652);
nand UO_204 (O_204,N_14570,N_14736);
nand UO_205 (O_205,N_13456,N_14105);
xnor UO_206 (O_206,N_12763,N_13508);
xor UO_207 (O_207,N_13147,N_12645);
nor UO_208 (O_208,N_13377,N_14993);
xnor UO_209 (O_209,N_12497,N_13370);
or UO_210 (O_210,N_13209,N_14494);
and UO_211 (O_211,N_14919,N_13495);
nand UO_212 (O_212,N_12114,N_13233);
nor UO_213 (O_213,N_12919,N_12691);
xnor UO_214 (O_214,N_12076,N_13493);
and UO_215 (O_215,N_14130,N_13132);
xnor UO_216 (O_216,N_12224,N_14263);
and UO_217 (O_217,N_12101,N_14568);
and UO_218 (O_218,N_12544,N_12080);
nand UO_219 (O_219,N_13226,N_13492);
nand UO_220 (O_220,N_12547,N_12589);
xnor UO_221 (O_221,N_12327,N_12747);
xnor UO_222 (O_222,N_13126,N_12861);
xor UO_223 (O_223,N_12968,N_12847);
or UO_224 (O_224,N_12537,N_13700);
nor UO_225 (O_225,N_12418,N_12463);
and UO_226 (O_226,N_14722,N_14622);
xor UO_227 (O_227,N_13300,N_13592);
nand UO_228 (O_228,N_12570,N_14851);
nor UO_229 (O_229,N_14873,N_12851);
or UO_230 (O_230,N_13114,N_13651);
nand UO_231 (O_231,N_14347,N_14407);
xnor UO_232 (O_232,N_12420,N_12029);
and UO_233 (O_233,N_14339,N_12994);
or UO_234 (O_234,N_14973,N_14928);
nand UO_235 (O_235,N_14875,N_13056);
nor UO_236 (O_236,N_12649,N_12969);
and UO_237 (O_237,N_14337,N_12484);
nand UO_238 (O_238,N_13712,N_12722);
nor UO_239 (O_239,N_12376,N_14859);
nor UO_240 (O_240,N_12337,N_12147);
xor UO_241 (O_241,N_14998,N_12373);
xor UO_242 (O_242,N_14705,N_14280);
nand UO_243 (O_243,N_12144,N_13451);
and UO_244 (O_244,N_12917,N_13159);
nand UO_245 (O_245,N_13806,N_14026);
xnor UO_246 (O_246,N_13028,N_13805);
or UO_247 (O_247,N_12380,N_13384);
and UO_248 (O_248,N_13920,N_14417);
and UO_249 (O_249,N_14121,N_12447);
or UO_250 (O_250,N_13342,N_13137);
nor UO_251 (O_251,N_13810,N_12464);
nand UO_252 (O_252,N_12901,N_14747);
nand UO_253 (O_253,N_12434,N_14259);
xnor UO_254 (O_254,N_14617,N_12808);
or UO_255 (O_255,N_12815,N_12775);
or UO_256 (O_256,N_13241,N_13709);
nand UO_257 (O_257,N_13141,N_12437);
or UO_258 (O_258,N_12767,N_13678);
xnor UO_259 (O_259,N_14423,N_13577);
xnor UO_260 (O_260,N_13513,N_13516);
or UO_261 (O_261,N_13813,N_13884);
and UO_262 (O_262,N_12353,N_13946);
nor UO_263 (O_263,N_12422,N_12225);
nand UO_264 (O_264,N_13327,N_13693);
nor UO_265 (O_265,N_12282,N_14905);
nand UO_266 (O_266,N_14378,N_12335);
xor UO_267 (O_267,N_14800,N_14122);
nand UO_268 (O_268,N_13118,N_13449);
xnor UO_269 (O_269,N_14331,N_12638);
or UO_270 (O_270,N_14181,N_13142);
and UO_271 (O_271,N_13102,N_14309);
and UO_272 (O_272,N_12825,N_13853);
or UO_273 (O_273,N_13979,N_13174);
or UO_274 (O_274,N_13395,N_14391);
and UO_275 (O_275,N_13183,N_13278);
nor UO_276 (O_276,N_12339,N_12772);
nand UO_277 (O_277,N_14969,N_14813);
or UO_278 (O_278,N_12028,N_12683);
nor UO_279 (O_279,N_14173,N_12323);
and UO_280 (O_280,N_13509,N_12482);
or UO_281 (O_281,N_12564,N_12204);
nand UO_282 (O_282,N_14155,N_14850);
and UO_283 (O_283,N_13879,N_14496);
xor UO_284 (O_284,N_14757,N_14148);
nor UO_285 (O_285,N_12948,N_13216);
nand UO_286 (O_286,N_13351,N_14476);
xor UO_287 (O_287,N_14784,N_12840);
nor UO_288 (O_288,N_14699,N_14557);
or UO_289 (O_289,N_14560,N_12807);
and UO_290 (O_290,N_12494,N_13846);
or UO_291 (O_291,N_12590,N_13682);
nand UO_292 (O_292,N_12347,N_12510);
nor UO_293 (O_293,N_12098,N_14812);
nor UO_294 (O_294,N_12644,N_13037);
nor UO_295 (O_295,N_14158,N_14303);
nand UO_296 (O_296,N_14338,N_12898);
xor UO_297 (O_297,N_12254,N_13669);
nor UO_298 (O_298,N_12983,N_12957);
or UO_299 (O_299,N_12762,N_12011);
or UO_300 (O_300,N_14336,N_14487);
xnor UO_301 (O_301,N_14946,N_12227);
nor UO_302 (O_302,N_13007,N_12755);
and UO_303 (O_303,N_14683,N_12287);
or UO_304 (O_304,N_12945,N_12338);
nor UO_305 (O_305,N_12460,N_13967);
xor UO_306 (O_306,N_13860,N_12153);
nor UO_307 (O_307,N_13372,N_13423);
and UO_308 (O_308,N_12083,N_13714);
or UO_309 (O_309,N_14222,N_12167);
or UO_310 (O_310,N_14438,N_12938);
and UO_311 (O_311,N_13773,N_14832);
nand UO_312 (O_312,N_12402,N_13688);
nand UO_313 (O_313,N_13845,N_12766);
or UO_314 (O_314,N_13346,N_13308);
xor UO_315 (O_315,N_14006,N_14162);
nor UO_316 (O_316,N_12052,N_14301);
and UO_317 (O_317,N_12263,N_13095);
xnor UO_318 (O_318,N_14888,N_13178);
or UO_319 (O_319,N_13984,N_14647);
nand UO_320 (O_320,N_12726,N_12723);
xor UO_321 (O_321,N_14997,N_12826);
and UO_322 (O_322,N_12260,N_12435);
nor UO_323 (O_323,N_13522,N_12552);
nand UO_324 (O_324,N_12886,N_14376);
or UO_325 (O_325,N_13165,N_12999);
xnor UO_326 (O_326,N_13191,N_14348);
nand UO_327 (O_327,N_13093,N_13591);
nand UO_328 (O_328,N_12839,N_14477);
and UO_329 (O_329,N_13850,N_13176);
and UO_330 (O_330,N_14234,N_12532);
nor UO_331 (O_331,N_13757,N_12596);
xnor UO_332 (O_332,N_13316,N_13112);
and UO_333 (O_333,N_14189,N_12856);
nand UO_334 (O_334,N_13325,N_12047);
or UO_335 (O_335,N_13890,N_13569);
and UO_336 (O_336,N_12560,N_12985);
xor UO_337 (O_337,N_14614,N_14751);
or UO_338 (O_338,N_14057,N_12923);
and UO_339 (O_339,N_12671,N_13197);
and UO_340 (O_340,N_12594,N_14590);
xnor UO_341 (O_341,N_12910,N_12916);
or UO_342 (O_342,N_14323,N_14269);
nor UO_343 (O_343,N_14449,N_13296);
and UO_344 (O_344,N_12681,N_13705);
nand UO_345 (O_345,N_13416,N_12765);
nand UO_346 (O_346,N_14180,N_13915);
xnor UO_347 (O_347,N_12611,N_14474);
nand UO_348 (O_348,N_13430,N_12330);
and UO_349 (O_349,N_12479,N_13644);
and UO_350 (O_350,N_12064,N_12234);
nor UO_351 (O_351,N_12641,N_12354);
and UO_352 (O_352,N_13221,N_12812);
xor UO_353 (O_353,N_12058,N_14525);
nor UO_354 (O_354,N_12441,N_14322);
nor UO_355 (O_355,N_12525,N_14467);
nand UO_356 (O_356,N_14204,N_14743);
nor UO_357 (O_357,N_14490,N_12310);
nand UO_358 (O_358,N_13326,N_14093);
xor UO_359 (O_359,N_12773,N_13264);
xor UO_360 (O_360,N_14624,N_13298);
nor UO_361 (O_361,N_13388,N_14852);
or UO_362 (O_362,N_13362,N_14685);
xnor UO_363 (O_363,N_14062,N_13196);
or UO_364 (O_364,N_12145,N_14837);
nor UO_365 (O_365,N_12618,N_13239);
and UO_366 (O_366,N_14400,N_13702);
or UO_367 (O_367,N_14900,N_14435);
and UO_368 (O_368,N_13562,N_12377);
or UO_369 (O_369,N_14485,N_12637);
or UO_370 (O_370,N_14092,N_12827);
xnor UO_371 (O_371,N_12308,N_12461);
nor UO_372 (O_372,N_14554,N_14343);
or UO_373 (O_373,N_12859,N_12776);
nand UO_374 (O_374,N_14547,N_12729);
xor UO_375 (O_375,N_13425,N_14906);
nand UO_376 (O_376,N_14019,N_13964);
xnor UO_377 (O_377,N_12318,N_12770);
or UO_378 (O_378,N_12838,N_13612);
nand UO_379 (O_379,N_12920,N_12211);
nand UO_380 (O_380,N_12250,N_13401);
or UO_381 (O_381,N_14730,N_12610);
and UO_382 (O_382,N_14697,N_14915);
nor UO_383 (O_383,N_14172,N_12118);
nand UO_384 (O_384,N_13641,N_13567);
nand UO_385 (O_385,N_14575,N_14524);
and UO_386 (O_386,N_12698,N_12890);
or UO_387 (O_387,N_12245,N_12499);
xnor UO_388 (O_388,N_13215,N_12120);
nand UO_389 (O_389,N_13815,N_14830);
and UO_390 (O_390,N_13686,N_13973);
nor UO_391 (O_391,N_14515,N_12274);
or UO_392 (O_392,N_14692,N_14073);
and UO_393 (O_393,N_13801,N_14698);
or UO_394 (O_394,N_12882,N_12096);
nand UO_395 (O_395,N_14637,N_12030);
xnor UO_396 (O_396,N_13287,N_12431);
nor UO_397 (O_397,N_13312,N_13645);
xnor UO_398 (O_398,N_13783,N_14497);
and UO_399 (O_399,N_13426,N_13096);
xnor UO_400 (O_400,N_13692,N_12468);
nand UO_401 (O_401,N_12270,N_14241);
or UO_402 (O_402,N_12971,N_13161);
and UO_403 (O_403,N_13066,N_14546);
nor UO_404 (O_404,N_12415,N_12958);
and UO_405 (O_405,N_12909,N_13756);
or UO_406 (O_406,N_13177,N_13092);
or UO_407 (O_407,N_13791,N_14365);
or UO_408 (O_408,N_12140,N_13696);
nand UO_409 (O_409,N_14566,N_14077);
xnor UO_410 (O_410,N_13348,N_12180);
nand UO_411 (O_411,N_12669,N_13870);
and UO_412 (O_412,N_14434,N_14714);
nand UO_413 (O_413,N_13555,N_13382);
or UO_414 (O_414,N_14910,N_13009);
nand UO_415 (O_415,N_13905,N_13694);
or UO_416 (O_416,N_14436,N_12921);
or UO_417 (O_417,N_12046,N_12023);
or UO_418 (O_418,N_14636,N_12021);
and UO_419 (O_419,N_14095,N_12244);
and UO_420 (O_420,N_12977,N_13610);
nor UO_421 (O_421,N_14719,N_12408);
and UO_422 (O_422,N_14385,N_13402);
xnor UO_423 (O_423,N_14752,N_14677);
or UO_424 (O_424,N_12078,N_12223);
and UO_425 (O_425,N_12757,N_13494);
or UO_426 (O_426,N_12561,N_13754);
and UO_427 (O_427,N_13088,N_13748);
and UO_428 (O_428,N_14972,N_14680);
nand UO_429 (O_429,N_13248,N_13635);
xnor UO_430 (O_430,N_14893,N_14366);
xor UO_431 (O_431,N_14861,N_12199);
nand UO_432 (O_432,N_13910,N_13989);
xor UO_433 (O_433,N_13938,N_12758);
nand UO_434 (O_434,N_14353,N_14819);
xor UO_435 (O_435,N_13280,N_13881);
or UO_436 (O_436,N_12586,N_13899);
xor UO_437 (O_437,N_12674,N_13643);
xnor UO_438 (O_438,N_12014,N_14089);
nor UO_439 (O_439,N_13914,N_14821);
xor UO_440 (O_440,N_12150,N_12060);
nand UO_441 (O_441,N_14018,N_12291);
xnor UO_442 (O_442,N_14877,N_12387);
and UO_443 (O_443,N_14167,N_14272);
and UO_444 (O_444,N_14544,N_13778);
xor UO_445 (O_445,N_12631,N_13286);
and UO_446 (O_446,N_12549,N_14509);
nor UO_447 (O_447,N_12178,N_14931);
nand UO_448 (O_448,N_12003,N_14653);
xor UO_449 (O_449,N_12364,N_14886);
xor UO_450 (O_450,N_12417,N_12887);
xnor UO_451 (O_451,N_13214,N_14820);
nand UO_452 (O_452,N_13085,N_13854);
xnor UO_453 (O_453,N_14643,N_13042);
nand UO_454 (O_454,N_12922,N_14675);
or UO_455 (O_455,N_12451,N_12043);
nand UO_456 (O_456,N_12019,N_13788);
and UO_457 (O_457,N_12587,N_14522);
nand UO_458 (O_458,N_13942,N_13468);
or UO_459 (O_459,N_12093,N_12992);
and UO_460 (O_460,N_13857,N_14790);
and UO_461 (O_461,N_13759,N_14398);
or UO_462 (O_462,N_12197,N_13663);
xor UO_463 (O_463,N_12137,N_14777);
or UO_464 (O_464,N_13774,N_14580);
nand UO_465 (O_465,N_12599,N_13201);
nor UO_466 (O_466,N_14668,N_14160);
xor UO_467 (O_467,N_13422,N_13213);
xor UO_468 (O_468,N_13704,N_12169);
xor UO_469 (O_469,N_13901,N_14903);
and UO_470 (O_470,N_13466,N_14329);
nor UO_471 (O_471,N_13962,N_12951);
and UO_472 (O_472,N_14333,N_14945);
nand UO_473 (O_473,N_13655,N_13257);
and UO_474 (O_474,N_12913,N_14594);
nor UO_475 (O_475,N_14732,N_13117);
or UO_476 (O_476,N_14111,N_13083);
or UO_477 (O_477,N_14060,N_13507);
or UO_478 (O_478,N_13930,N_12759);
xor UO_479 (O_479,N_12665,N_12811);
nand UO_480 (O_480,N_13725,N_13755);
nor UO_481 (O_481,N_12237,N_14716);
nor UO_482 (O_482,N_14480,N_14404);
nand UO_483 (O_483,N_12527,N_12979);
and UO_484 (O_484,N_14843,N_12267);
nand UO_485 (O_485,N_13087,N_14884);
and UO_486 (O_486,N_12508,N_12174);
nor UO_487 (O_487,N_14927,N_13480);
nor UO_488 (O_488,N_14070,N_13381);
or UO_489 (O_489,N_14510,N_14785);
xnor UO_490 (O_490,N_13412,N_12733);
or UO_491 (O_491,N_14444,N_13738);
and UO_492 (O_492,N_12210,N_12796);
nand UO_493 (O_493,N_13283,N_14726);
and UO_494 (O_494,N_14232,N_13061);
or UO_495 (O_495,N_12819,N_12301);
nor UO_496 (O_496,N_13305,N_13608);
and UO_497 (O_497,N_12926,N_13187);
and UO_498 (O_498,N_12954,N_13599);
nand UO_499 (O_499,N_13909,N_12433);
and UO_500 (O_500,N_14912,N_13768);
xnor UO_501 (O_501,N_13670,N_14874);
xor UO_502 (O_502,N_12107,N_13649);
and UO_503 (O_503,N_14761,N_14581);
and UO_504 (O_504,N_13546,N_12406);
xnor UO_505 (O_505,N_14841,N_13077);
or UO_506 (O_506,N_12392,N_13366);
nand UO_507 (O_507,N_14678,N_12369);
and UO_508 (O_508,N_13518,N_13208);
xor UO_509 (O_509,N_13837,N_14923);
or UO_510 (O_510,N_14538,N_12113);
nor UO_511 (O_511,N_13259,N_12253);
xor UO_512 (O_512,N_12395,N_13131);
nor UO_513 (O_513,N_13075,N_12305);
nand UO_514 (O_514,N_14769,N_14161);
and UO_515 (O_515,N_14169,N_12061);
xnor UO_516 (O_516,N_12798,N_14489);
nand UO_517 (O_517,N_13051,N_14159);
nand UO_518 (O_518,N_14221,N_13820);
or UO_519 (O_519,N_13542,N_14010);
xor UO_520 (O_520,N_12929,N_14271);
xnor UO_521 (O_521,N_12598,N_13951);
or UO_522 (O_522,N_13601,N_14252);
nor UO_523 (O_523,N_12822,N_13204);
nor UO_524 (O_524,N_12663,N_14988);
nand UO_525 (O_525,N_12727,N_14523);
nor UO_526 (O_526,N_13076,N_14426);
and UO_527 (O_527,N_12123,N_14527);
nor UO_528 (O_528,N_14782,N_13572);
nor UO_529 (O_529,N_13138,N_14577);
and UO_530 (O_530,N_13564,N_13976);
and UO_531 (O_531,N_14120,N_12526);
or UO_532 (O_532,N_12202,N_14356);
and UO_533 (O_533,N_13419,N_12442);
xnor UO_534 (O_534,N_12953,N_12646);
or UO_535 (O_535,N_14855,N_12089);
and UO_536 (O_536,N_12229,N_14153);
or UO_537 (O_537,N_14737,N_13355);
or UO_538 (O_538,N_14374,N_13109);
and UO_539 (O_539,N_14170,N_14265);
nor UO_540 (O_540,N_12325,N_12166);
xor UO_541 (O_541,N_13963,N_12515);
nor UO_542 (O_542,N_12311,N_14542);
and UO_543 (O_543,N_14926,N_12378);
xnor UO_544 (O_544,N_12790,N_14735);
or UO_545 (O_545,N_14609,N_12465);
nand UO_546 (O_546,N_14144,N_14176);
and UO_547 (O_547,N_12304,N_13701);
and UO_548 (O_548,N_14957,N_14831);
nand UO_549 (O_549,N_13038,N_13365);
or UO_550 (O_550,N_13580,N_14386);
nor UO_551 (O_551,N_12062,N_14539);
nand UO_552 (O_552,N_14119,N_14607);
nor UO_553 (O_553,N_12000,N_14033);
xor UO_554 (O_554,N_14618,N_13741);
nand UO_555 (O_555,N_13583,N_14216);
xnor UO_556 (O_556,N_13166,N_13135);
nand UO_557 (O_557,N_14443,N_13916);
nand UO_558 (O_558,N_14050,N_13399);
nand UO_559 (O_559,N_13724,N_13273);
and UO_560 (O_560,N_14082,N_13329);
xor UO_561 (O_561,N_12281,N_12670);
xnor UO_562 (O_562,N_14041,N_13662);
or UO_563 (O_563,N_14413,N_12425);
nand UO_564 (O_564,N_13212,N_14862);
nor UO_565 (O_565,N_12506,N_14567);
nor UO_566 (O_566,N_13929,N_14584);
xnor UO_567 (O_567,N_13110,N_13198);
xnor UO_568 (O_568,N_13907,N_12622);
xnor UO_569 (O_569,N_14412,N_14445);
nand UO_570 (O_570,N_12191,N_13199);
xor UO_571 (O_571,N_13023,N_14207);
xor UO_572 (O_572,N_13611,N_13747);
xor UO_573 (O_573,N_13880,N_14882);
nand UO_574 (O_574,N_12389,N_13897);
nor UO_575 (O_575,N_12018,N_12962);
nor UO_576 (O_576,N_14656,N_12131);
nand UO_577 (O_577,N_13185,N_14034);
or UO_578 (O_578,N_12528,N_13703);
and UO_579 (O_579,N_12165,N_12184);
xor UO_580 (O_580,N_14481,N_12739);
and UO_581 (O_581,N_14532,N_14835);
nand UO_582 (O_582,N_13537,N_13931);
and UO_583 (O_583,N_12725,N_14370);
or UO_584 (O_584,N_12055,N_12372);
nand UO_585 (O_585,N_12889,N_14457);
nor UO_586 (O_586,N_14858,N_14279);
xnor UO_587 (O_587,N_14810,N_13369);
or UO_588 (O_588,N_12491,N_13770);
and UO_589 (O_589,N_14471,N_12970);
nand UO_590 (O_590,N_13314,N_12915);
xnor UO_591 (O_591,N_14197,N_14453);
or UO_592 (O_592,N_12088,N_14264);
or UO_593 (O_593,N_13749,N_12130);
xor UO_594 (O_594,N_13323,N_12661);
or UO_595 (O_595,N_14447,N_13044);
and UO_596 (O_596,N_12634,N_12714);
or UO_597 (O_597,N_13743,N_12821);
nor UO_598 (O_598,N_12361,N_12908);
xor UO_599 (O_599,N_14571,N_13173);
nand UO_600 (O_600,N_12445,N_13953);
or UO_601 (O_601,N_14885,N_14166);
xnor UO_602 (O_602,N_14463,N_14029);
or UO_603 (O_603,N_14150,N_13804);
and UO_604 (O_604,N_12288,N_12151);
or UO_605 (O_605,N_13823,N_12743);
xor UO_606 (O_606,N_13478,N_14569);
and UO_607 (O_607,N_12273,N_12424);
and UO_608 (O_608,N_12272,N_14012);
or UO_609 (O_609,N_13207,N_14788);
nor UO_610 (O_610,N_13266,N_12667);
xnor UO_611 (O_611,N_13631,N_12697);
nor UO_612 (O_612,N_14721,N_12215);
nor UO_613 (O_613,N_14415,N_12846);
xor UO_614 (O_614,N_14838,N_13181);
nand UO_615 (O_615,N_12448,N_14297);
nor UO_616 (O_616,N_12403,N_12717);
and UO_617 (O_617,N_13711,N_12117);
xor UO_618 (O_618,N_14774,N_14816);
nor UO_619 (O_619,N_13097,N_14099);
nor UO_620 (O_620,N_12991,N_12230);
nor UO_621 (O_621,N_13274,N_14441);
nand UO_622 (O_622,N_13380,N_14899);
or UO_623 (O_623,N_12500,N_13359);
xnor UO_624 (O_624,N_14996,N_13874);
xnor UO_625 (O_625,N_13941,N_12057);
or UO_626 (O_626,N_13833,N_12232);
and UO_627 (O_627,N_12022,N_13206);
and UO_628 (O_628,N_13642,N_14013);
nand UO_629 (O_629,N_12652,N_12592);
xor UO_630 (O_630,N_14286,N_13943);
nor UO_631 (O_631,N_13977,N_14724);
nor UO_632 (O_632,N_14291,N_14203);
or UO_633 (O_633,N_13227,N_12624);
or UO_634 (O_634,N_12314,N_13552);
nor UO_635 (O_635,N_12135,N_14937);
nand UO_636 (O_636,N_14828,N_14596);
or UO_637 (O_637,N_14925,N_14140);
or UO_638 (O_638,N_13604,N_13503);
or UO_639 (O_639,N_14939,N_12320);
nor UO_640 (O_640,N_13010,N_13831);
xnor UO_641 (O_641,N_12657,N_13887);
nor UO_642 (O_642,N_13392,N_13722);
and UO_643 (O_643,N_14044,N_14254);
xnor UO_644 (O_644,N_14896,N_14104);
xor UO_645 (O_645,N_14387,N_12139);
or UO_646 (O_646,N_12365,N_13289);
nor UO_647 (O_647,N_13364,N_12458);
xor UO_648 (O_648,N_14552,N_12261);
nor UO_649 (O_649,N_14037,N_13766);
and UO_650 (O_650,N_14533,N_12580);
xor UO_651 (O_651,N_12196,N_13230);
and UO_652 (O_652,N_14865,N_13172);
xor UO_653 (O_653,N_13935,N_12419);
or UO_654 (O_654,N_13068,N_13627);
nand UO_655 (O_655,N_13324,N_12302);
nand UO_656 (O_656,N_13647,N_13971);
nor UO_657 (O_657,N_13713,N_12903);
nor UO_658 (O_658,N_14648,N_12475);
xor UO_659 (O_659,N_14045,N_14518);
or UO_660 (O_660,N_12629,N_12097);
nor UO_661 (O_661,N_14890,N_14014);
nand UO_662 (O_662,N_13529,N_12686);
xnor UO_663 (O_663,N_14548,N_14768);
and UO_664 (O_664,N_13228,N_14142);
and UO_665 (O_665,N_13378,N_13554);
nor UO_666 (O_666,N_14940,N_14849);
or UO_667 (O_667,N_14913,N_14219);
xnor UO_668 (O_668,N_12483,N_13616);
xnor UO_669 (O_669,N_14421,N_12855);
and UO_670 (O_670,N_13800,N_12959);
xor UO_671 (O_671,N_14236,N_14174);
nor UO_672 (O_672,N_14399,N_12079);
or UO_673 (O_673,N_14307,N_14151);
xor UO_674 (O_674,N_13527,N_12413);
xnor UO_675 (O_675,N_12837,N_13660);
xnor UO_676 (O_676,N_12771,N_13510);
xor UO_677 (O_677,N_13018,N_13834);
or UO_678 (O_678,N_13246,N_13251);
nor UO_679 (O_679,N_14420,N_13057);
xor UO_680 (O_680,N_14983,N_14979);
or UO_681 (O_681,N_12960,N_13544);
and UO_682 (O_682,N_12163,N_13205);
nand UO_683 (O_683,N_13997,N_12283);
xnor UO_684 (O_684,N_13780,N_13184);
and UO_685 (O_685,N_12899,N_12397);
xor UO_686 (O_686,N_14712,N_13561);
and UO_687 (O_687,N_14578,N_12266);
xnor UO_688 (O_688,N_12466,N_13668);
nor UO_689 (O_689,N_12764,N_13538);
xnor UO_690 (O_690,N_14058,N_12243);
nor UO_691 (O_691,N_14586,N_13718);
nor UO_692 (O_692,N_13966,N_13622);
or UO_693 (O_693,N_12834,N_14091);
or UO_694 (O_694,N_12626,N_13436);
nand UO_695 (O_695,N_14990,N_14047);
and UO_696 (O_696,N_12344,N_12858);
or UO_697 (O_697,N_13148,N_14295);
and UO_698 (O_698,N_12780,N_12603);
nand UO_699 (O_699,N_14638,N_14938);
xnor UO_700 (O_700,N_13340,N_14612);
nor UO_701 (O_701,N_13027,N_14009);
nand UO_702 (O_702,N_13158,N_13525);
nor UO_703 (O_703,N_13666,N_14132);
nand UO_704 (O_704,N_14880,N_14723);
nand UO_705 (O_705,N_14096,N_14495);
nor UO_706 (O_706,N_13020,N_13925);
and UO_707 (O_707,N_13275,N_13084);
nand UO_708 (O_708,N_13435,N_14950);
or UO_709 (O_709,N_12794,N_12706);
and UO_710 (O_710,N_14559,N_14842);
or UO_711 (O_711,N_13863,N_14688);
nand UO_712 (O_712,N_13830,N_13506);
and UO_713 (O_713,N_14134,N_14177);
xor UO_714 (O_714,N_12156,N_13584);
xor UO_715 (O_715,N_14411,N_13240);
nor UO_716 (O_716,N_13021,N_13022);
nand UO_717 (O_717,N_14442,N_14749);
or UO_718 (O_718,N_14315,N_14962);
xnor UO_719 (O_719,N_14258,N_14776);
and UO_720 (O_720,N_14654,N_14330);
xor UO_721 (O_721,N_14537,N_13429);
or UO_722 (O_722,N_12660,N_14917);
or UO_723 (O_723,N_14186,N_14185);
xor UO_724 (O_724,N_13974,N_13279);
nor UO_725 (O_725,N_14658,N_14573);
nand UO_726 (O_726,N_13472,N_14281);
xnor UO_727 (O_727,N_14650,N_14592);
or UO_728 (O_728,N_13517,N_14230);
xor UO_729 (O_729,N_14564,N_14054);
nand UO_730 (O_730,N_14536,N_13950);
or UO_731 (O_731,N_13818,N_13041);
nor UO_732 (O_732,N_14056,N_13383);
or UO_733 (O_733,N_13035,N_14454);
and UO_734 (O_734,N_12558,N_13271);
nor UO_735 (O_735,N_12956,N_12536);
and UO_736 (O_736,N_12400,N_12359);
nand UO_737 (O_737,N_12568,N_12555);
nand UO_738 (O_738,N_13785,N_13218);
and UO_739 (O_739,N_12262,N_12015);
nand UO_740 (O_740,N_12947,N_12744);
xor UO_741 (O_741,N_14296,N_13970);
or UO_742 (O_742,N_14711,N_14966);
and UO_743 (O_743,N_12666,N_13826);
or UO_744 (O_744,N_13306,N_13450);
xor UO_745 (O_745,N_12894,N_14277);
and UO_746 (O_746,N_14878,N_13437);
xor UO_747 (O_747,N_14124,N_14114);
nor UO_748 (O_748,N_12049,N_12731);
xnor UO_749 (O_749,N_14335,N_12835);
or UO_750 (O_750,N_12316,N_13121);
nor UO_751 (O_751,N_14008,N_14895);
and UO_752 (O_752,N_14742,N_14666);
xnor UO_753 (O_753,N_14825,N_14223);
nor UO_754 (O_754,N_12514,N_12912);
or UO_755 (O_755,N_13462,N_13107);
and UO_756 (O_756,N_12613,N_14390);
nor UO_757 (O_757,N_14727,N_13867);
xnor UO_758 (O_758,N_13267,N_14516);
xnor UO_759 (O_759,N_13814,N_13630);
and UO_760 (O_760,N_13453,N_14935);
xor UO_761 (O_761,N_12809,N_14106);
nor UO_762 (O_762,N_13394,N_12041);
nor UO_763 (O_763,N_12607,N_14345);
nand UO_764 (O_764,N_12640,N_12574);
xnor UO_765 (O_765,N_13913,N_13779);
nor UO_766 (O_766,N_13428,N_12285);
nand UO_767 (O_767,N_14090,N_12192);
nor UO_768 (O_768,N_12814,N_14953);
or UO_769 (O_769,N_14908,N_14233);
nand UO_770 (O_770,N_14951,N_13727);
nor UO_771 (O_771,N_12803,N_13261);
and UO_772 (O_772,N_14640,N_13171);
xnor UO_773 (O_773,N_13856,N_13049);
nor UO_774 (O_774,N_12309,N_14229);
and UO_775 (O_775,N_12981,N_13069);
and UO_776 (O_776,N_12462,N_13223);
or UO_777 (O_777,N_13104,N_12628);
and UO_778 (O_778,N_14190,N_12375);
and UO_779 (O_779,N_13356,N_12436);
or UO_780 (O_780,N_13162,N_14817);
or UO_781 (O_781,N_13557,N_13519);
nor UO_782 (O_782,N_14135,N_14341);
xnor UO_783 (O_783,N_12769,N_12975);
or UO_784 (O_784,N_12219,N_13396);
or UO_785 (O_785,N_14256,N_14970);
or UO_786 (O_786,N_12577,N_13934);
nand UO_787 (O_787,N_12829,N_12173);
nand UO_788 (O_788,N_14778,N_12099);
nor UO_789 (O_789,N_12553,N_12358);
nand UO_790 (O_790,N_12409,N_12978);
and UO_791 (O_791,N_12830,N_13921);
and UO_792 (O_792,N_14046,N_13556);
or UO_793 (O_793,N_14960,N_13858);
xor UO_794 (O_794,N_13589,N_13675);
nand UO_795 (O_795,N_14225,N_12279);
nor UO_796 (O_796,N_13763,N_13417);
or UO_797 (O_797,N_14904,N_12621);
or UO_798 (O_798,N_13811,N_14242);
and UO_799 (O_799,N_14623,N_13618);
or UO_800 (O_800,N_13335,N_13771);
xor UO_801 (O_801,N_14015,N_14553);
xnor UO_802 (O_802,N_13232,N_13116);
and UO_803 (O_803,N_14344,N_12842);
xnor UO_804 (O_804,N_12987,N_13883);
nand UO_805 (O_805,N_12675,N_13098);
nand UO_806 (O_806,N_12845,N_14629);
xor UO_807 (O_807,N_14043,N_14967);
nand UO_808 (O_808,N_12548,N_13533);
and UO_809 (O_809,N_13081,N_14363);
nand UO_810 (O_810,N_13875,N_13839);
nor UO_811 (O_811,N_12033,N_12993);
and UO_812 (O_812,N_12655,N_14382);
xor UO_813 (O_813,N_13091,N_14670);
and UO_814 (O_814,N_12133,N_13219);
nor UO_815 (O_815,N_14806,N_13194);
xnor UO_816 (O_816,N_13540,N_14791);
xnor UO_817 (O_817,N_13500,N_12955);
nand UO_818 (O_818,N_13690,N_14720);
xor UO_819 (O_819,N_14500,N_12965);
or UO_820 (O_820,N_12486,N_13334);
nand UO_821 (O_821,N_13578,N_12129);
and UO_822 (O_822,N_13609,N_14478);
or UO_823 (O_823,N_13764,N_12844);
and UO_824 (O_824,N_14048,N_12932);
or UO_825 (O_825,N_14083,N_13190);
nor UO_826 (O_826,N_13052,N_14540);
or UO_827 (O_827,N_12393,N_12559);
and UO_828 (O_828,N_14432,N_12251);
nor UO_829 (O_829,N_14253,N_14016);
nor UO_830 (O_830,N_14649,N_12027);
or UO_831 (O_831,N_13543,N_13301);
xnor UO_832 (O_832,N_12067,N_14995);
nor UO_833 (O_833,N_13203,N_13443);
or UO_834 (O_834,N_13149,N_14762);
and UO_835 (O_835,N_13231,N_14084);
nor UO_836 (O_836,N_13475,N_12489);
xnor UO_837 (O_837,N_13189,N_12220);
xor UO_838 (O_838,N_13520,N_13496);
or UO_839 (O_839,N_13803,N_13065);
xor UO_840 (O_840,N_12942,N_12158);
or UO_841 (O_841,N_13596,N_12692);
nand UO_842 (O_842,N_12925,N_12181);
nand UO_843 (O_843,N_13153,N_12802);
and UO_844 (O_844,N_12550,N_12512);
nor UO_845 (O_845,N_14416,N_13371);
xor UO_846 (O_846,N_14744,N_12258);
xnor UO_847 (O_847,N_14632,N_12476);
nand UO_848 (O_848,N_12684,N_14734);
nand UO_849 (O_849,N_12980,N_13133);
xor UO_850 (O_850,N_14689,N_14275);
xor UO_851 (O_851,N_13353,N_13015);
xor UO_852 (O_852,N_13621,N_14359);
nand UO_853 (O_853,N_13698,N_12017);
nor UO_854 (O_854,N_14049,N_12849);
or UO_855 (O_855,N_12715,N_14141);
nand UO_856 (O_856,N_13124,N_14868);
or UO_857 (O_857,N_14133,N_13072);
xor UO_858 (O_858,N_14587,N_13790);
nand UO_859 (O_859,N_12719,N_14691);
xor UO_860 (O_860,N_13017,N_12429);
and UO_861 (O_861,N_14239,N_14827);
nand UO_862 (O_862,N_13320,N_13318);
nand UO_863 (O_863,N_13277,N_13511);
or UO_864 (O_864,N_13844,N_14787);
and UO_865 (O_865,N_13036,N_14388);
xor UO_866 (O_866,N_13745,N_14911);
and UO_867 (O_867,N_13994,N_13829);
nand UO_868 (O_868,N_14844,N_14793);
nand UO_869 (O_869,N_13202,N_12680);
or UO_870 (O_870,N_12831,N_12190);
or UO_871 (O_871,N_13600,N_14389);
nor UO_872 (O_872,N_13936,N_14708);
and UO_873 (O_873,N_13728,N_13832);
nand UO_874 (O_874,N_14218,N_14965);
xnor UO_875 (O_875,N_13723,N_14284);
and UO_876 (O_876,N_14922,N_14795);
xor UO_877 (O_877,N_13265,N_13864);
and UO_878 (O_878,N_13403,N_14152);
xor UO_879 (O_879,N_12248,N_14921);
or UO_880 (O_880,N_13291,N_12737);
xnor UO_881 (O_881,N_13090,N_12366);
nor UO_882 (O_882,N_14310,N_14549);
nand UO_883 (O_883,N_12742,N_14520);
xnor UO_884 (O_884,N_12633,N_14354);
or UO_885 (O_885,N_13322,N_14914);
xnor UO_886 (O_886,N_12294,N_14503);
nand UO_887 (O_887,N_13968,N_12122);
nand UO_888 (O_888,N_14512,N_12008);
nor UO_889 (O_889,N_14131,N_13357);
nor UO_890 (O_890,N_12650,N_12050);
nand UO_891 (O_891,N_12247,N_12300);
and UO_892 (O_892,N_12854,N_12928);
or UO_893 (O_893,N_12095,N_13945);
xnor UO_894 (O_894,N_12531,N_12259);
nand UO_895 (O_895,N_13575,N_12860);
nor UO_896 (O_896,N_14262,N_14860);
nand UO_897 (O_897,N_12584,N_12298);
or UO_898 (O_898,N_13898,N_14342);
xor UO_899 (O_899,N_13235,N_13794);
and UO_900 (O_900,N_14555,N_14188);
xor UO_901 (O_901,N_12134,N_12042);
or UO_902 (O_902,N_13784,N_13294);
nor UO_903 (O_903,N_12350,N_13560);
or UO_904 (O_904,N_14848,N_13986);
or UO_905 (O_905,N_13684,N_14273);
nand UO_906 (O_906,N_13144,N_12472);
nand UO_907 (O_907,N_13156,N_12216);
nor UO_908 (O_908,N_14030,N_14201);
nand UO_909 (O_909,N_13633,N_14401);
and UO_910 (O_910,N_14839,N_14000);
nor UO_911 (O_911,N_12943,N_14876);
nor UO_912 (O_912,N_14488,N_13058);
nand UO_913 (O_913,N_14287,N_13455);
nor UO_914 (O_914,N_14325,N_13796);
xor UO_915 (O_915,N_13445,N_14804);
nor UO_916 (O_916,N_12941,N_12306);
nor UO_917 (O_917,N_13648,N_13904);
and UO_918 (O_918,N_12585,N_14941);
nand UO_919 (O_919,N_14695,N_14115);
nor UO_920 (O_920,N_12183,N_12582);
nor UO_921 (O_921,N_12866,N_13415);
or UO_922 (O_922,N_14143,N_14486);
nand UO_923 (O_923,N_12931,N_12687);
nand UO_924 (O_924,N_14462,N_13397);
nor UO_925 (O_925,N_12949,N_14199);
xor UO_926 (O_926,N_14534,N_14439);
or UO_927 (O_927,N_12189,N_12416);
xnor UO_928 (O_928,N_12946,N_13646);
xnor UO_929 (O_929,N_13368,N_13276);
nor UO_930 (O_930,N_12545,N_13730);
nand UO_931 (O_931,N_12054,N_13067);
xor UO_932 (O_932,N_13029,N_12459);
nand UO_933 (O_933,N_12427,N_12756);
and UO_934 (O_934,N_14088,N_14406);
nand UO_935 (O_935,N_12111,N_13602);
nand UO_936 (O_936,N_13667,N_13535);
xor UO_937 (O_937,N_14834,N_13551);
or UO_938 (O_938,N_13016,N_13563);
xor UO_939 (O_939,N_13470,N_12871);
xor UO_940 (O_940,N_14943,N_13523);
nand UO_941 (O_941,N_13328,N_12608);
nand UO_942 (O_942,N_13536,N_13848);
nand UO_943 (O_943,N_13949,N_14846);
or UO_944 (O_944,N_13473,N_12214);
xnor UO_945 (O_945,N_14713,N_13816);
nor UO_946 (O_946,N_13762,N_14068);
nand UO_947 (O_947,N_13179,N_12084);
and UO_948 (O_948,N_12355,N_12109);
xnor UO_949 (O_949,N_14094,N_12106);
nand UO_950 (O_950,N_14430,N_14606);
and UO_951 (O_951,N_12672,N_12843);
and UO_952 (O_952,N_14765,N_14007);
nor UO_953 (O_953,N_13064,N_13317);
nor UO_954 (O_954,N_12296,N_14394);
xor UO_955 (O_955,N_12604,N_14268);
nor UO_956 (O_956,N_14833,N_12004);
nor UO_957 (O_957,N_12695,N_13452);
nand UO_958 (O_958,N_14733,N_12321);
xnor UO_959 (O_959,N_14616,N_14645);
and UO_960 (O_960,N_14081,N_14610);
xnor UO_961 (O_961,N_13566,N_13139);
nand UO_962 (O_962,N_14479,N_13164);
xor UO_963 (O_963,N_13797,N_14419);
and UO_964 (O_964,N_12148,N_14492);
xnor UO_965 (O_965,N_14410,N_14687);
and UO_966 (O_966,N_12168,N_12511);
nor UO_967 (O_967,N_12315,N_12290);
and UO_968 (O_968,N_13975,N_14011);
nor UO_969 (O_969,N_12063,N_12787);
and UO_970 (O_970,N_13547,N_12455);
or UO_971 (O_971,N_12034,N_14052);
nand UO_972 (O_972,N_13448,N_14414);
or UO_973 (O_973,N_12457,N_12324);
and UO_974 (O_974,N_13409,N_13163);
and UO_975 (O_975,N_13530,N_13146);
xor UO_976 (O_976,N_12410,N_13192);
xnor UO_977 (O_977,N_12449,N_13130);
xnor UO_978 (O_978,N_14460,N_14072);
nor UO_979 (O_979,N_12075,N_12753);
and UO_980 (O_980,N_12477,N_13385);
xor UO_981 (O_981,N_14766,N_14739);
nor UO_982 (O_982,N_13005,N_14508);
nor UO_983 (O_983,N_14869,N_13272);
nand UO_984 (O_984,N_12973,N_13777);
nor UO_985 (O_985,N_14327,N_12509);
and UO_986 (O_986,N_12155,N_13360);
xor UO_987 (O_987,N_14340,N_12523);
and UO_988 (O_988,N_12748,N_14604);
nand UO_989 (O_989,N_13260,N_14165);
nor UO_990 (O_990,N_12368,N_14984);
or UO_991 (O_991,N_13876,N_13155);
and UO_992 (O_992,N_14276,N_14064);
nand UO_993 (O_993,N_14282,N_14987);
xor UO_994 (O_994,N_12864,N_13677);
xnor UO_995 (O_995,N_13825,N_14763);
and UO_996 (O_996,N_12313,N_13944);
and UO_997 (O_997,N_14328,N_14118);
xnor UO_998 (O_998,N_12768,N_12110);
and UO_999 (O_999,N_14191,N_12388);
xnor UO_1000 (O_1000,N_13354,N_13053);
xor UO_1001 (O_1001,N_14808,N_14944);
nor UO_1002 (O_1002,N_12252,N_12885);
and UO_1003 (O_1003,N_14901,N_12918);
xor UO_1004 (O_1004,N_12783,N_14040);
and UO_1005 (O_1005,N_12721,N_12732);
xor UO_1006 (O_1006,N_14644,N_13258);
nand UO_1007 (O_1007,N_14889,N_13268);
nand UO_1008 (O_1008,N_13358,N_12094);
xor UO_1009 (O_1009,N_14673,N_14061);
nor UO_1010 (O_1010,N_12752,N_12186);
nand UO_1011 (O_1011,N_12059,N_13410);
and UO_1012 (O_1012,N_14428,N_12832);
or UO_1013 (O_1013,N_12751,N_13750);
nor UO_1014 (O_1014,N_12857,N_14770);
nand UO_1015 (O_1015,N_13243,N_14949);
and UO_1016 (O_1016,N_14452,N_12006);
and UO_1017 (O_1017,N_12356,N_12044);
xnor UO_1018 (O_1018,N_13990,N_14822);
nor UO_1019 (O_1019,N_14163,N_12193);
or UO_1020 (O_1020,N_13011,N_14892);
nand UO_1021 (O_1021,N_14243,N_13993);
nand UO_1022 (O_1022,N_12884,N_12569);
and UO_1023 (O_1023,N_13623,N_14306);
or UO_1024 (O_1024,N_13379,N_12045);
nor UO_1025 (O_1025,N_12233,N_12379);
nand UO_1026 (O_1026,N_13304,N_13001);
or UO_1027 (O_1027,N_14069,N_14498);
or UO_1028 (O_1028,N_12138,N_14468);
nand UO_1029 (O_1029,N_14994,N_14642);
or UO_1030 (O_1030,N_12332,N_12501);
nand UO_1031 (O_1031,N_12639,N_14290);
xor UO_1032 (O_1032,N_13504,N_12085);
or UO_1033 (O_1033,N_12121,N_14932);
and UO_1034 (O_1034,N_13054,N_14302);
xor UO_1035 (O_1035,N_12430,N_13998);
or UO_1036 (O_1036,N_13101,N_14728);
xor UO_1037 (O_1037,N_13581,N_13111);
xor UO_1038 (O_1038,N_12972,N_14871);
nand UO_1039 (O_1039,N_14690,N_13614);
and UO_1040 (O_1040,N_12317,N_14550);
nand UO_1041 (O_1041,N_12933,N_13991);
nand UO_1042 (O_1042,N_14200,N_14108);
and UO_1043 (O_1043,N_12503,N_12362);
nand UO_1044 (O_1044,N_13315,N_13868);
nor UO_1045 (O_1045,N_14379,N_13707);
or UO_1046 (O_1046,N_14215,N_12792);
nand UO_1047 (O_1047,N_14220,N_14179);
nand UO_1048 (O_1048,N_14360,N_14872);
xor UO_1049 (O_1049,N_14796,N_13352);
xnor UO_1050 (O_1050,N_14318,N_12642);
nor UO_1051 (O_1051,N_12848,N_14332);
xnor UO_1052 (O_1052,N_12172,N_13400);
nor UO_1053 (O_1053,N_13013,N_14355);
nand UO_1054 (O_1054,N_12513,N_12450);
nor UO_1055 (O_1055,N_14772,N_13224);
and UO_1056 (O_1056,N_12401,N_13442);
nand UO_1057 (O_1057,N_12730,N_12881);
nor UO_1058 (O_1058,N_14261,N_12679);
or UO_1059 (O_1059,N_12071,N_12185);
or UO_1060 (O_1060,N_12179,N_12382);
xnor UO_1061 (O_1061,N_12205,N_14381);
xor UO_1062 (O_1062,N_13579,N_13746);
and UO_1063 (O_1063,N_14126,N_12636);
xnor UO_1064 (O_1064,N_14663,N_13157);
or UO_1065 (O_1065,N_13842,N_13789);
or UO_1066 (O_1066,N_14156,N_14352);
xnor UO_1067 (O_1067,N_12656,N_12777);
nor UO_1068 (O_1068,N_12541,N_14671);
and UO_1069 (O_1069,N_13336,N_12616);
nand UO_1070 (O_1070,N_14615,N_14667);
nand UO_1071 (O_1071,N_12562,N_13889);
or UO_1072 (O_1072,N_13720,N_14676);
and UO_1073 (O_1073,N_13654,N_12102);
nand UO_1074 (O_1074,N_13488,N_14038);
nor UO_1075 (O_1075,N_12982,N_12108);
nand UO_1076 (O_1076,N_12673,N_12249);
nor UO_1077 (O_1077,N_13404,N_12009);
nand UO_1078 (O_1078,N_14257,N_12893);
and UO_1079 (O_1079,N_12601,N_12269);
nor UO_1080 (O_1080,N_14696,N_14591);
or UO_1081 (O_1081,N_14718,N_13821);
xor UO_1082 (O_1082,N_14531,N_13739);
and UO_1083 (O_1083,N_12820,N_12718);
or UO_1084 (O_1084,N_13828,N_13937);
nand UO_1085 (O_1085,N_13238,N_14109);
xor UO_1086 (O_1086,N_14071,N_14395);
nand UO_1087 (O_1087,N_14458,N_14517);
or UO_1088 (O_1088,N_12391,N_12493);
and UO_1089 (O_1089,N_13605,N_12895);
or UO_1090 (O_1090,N_12896,N_12786);
nor UO_1091 (O_1091,N_12905,N_12791);
and UO_1092 (O_1092,N_14373,N_13565);
and UO_1093 (O_1093,N_14672,N_12708);
and UO_1094 (O_1094,N_14473,N_13719);
or UO_1095 (O_1095,N_12659,N_14319);
and UO_1096 (O_1096,N_13080,N_13003);
nor UO_1097 (O_1097,N_13245,N_14357);
or UO_1098 (O_1098,N_13699,N_12171);
or UO_1099 (O_1099,N_12813,N_12105);
and UO_1100 (O_1100,N_12824,N_12453);
nand UO_1101 (O_1101,N_14526,N_13742);
nor UO_1102 (O_1102,N_13871,N_14080);
nand UO_1103 (O_1103,N_14384,N_13708);
and UO_1104 (O_1104,N_12240,N_13431);
or UO_1105 (O_1105,N_13389,N_13956);
or UO_1106 (O_1106,N_12065,N_14929);
or UO_1107 (O_1107,N_14248,N_12103);
nand UO_1108 (O_1108,N_14409,N_13840);
or UO_1109 (O_1109,N_12217,N_14097);
xnor UO_1110 (O_1110,N_14465,N_14565);
and UO_1111 (O_1111,N_13025,N_13550);
nand UO_1112 (O_1112,N_14863,N_13119);
nor UO_1113 (O_1113,N_14854,N_13465);
xnor UO_1114 (O_1114,N_14975,N_12779);
xor UO_1115 (O_1115,N_14035,N_13888);
nor UO_1116 (O_1116,N_13253,N_12583);
nor UO_1117 (O_1117,N_14154,N_13769);
nor UO_1118 (O_1118,N_14267,N_12440);
xor UO_1119 (O_1119,N_13958,N_12116);
xnor UO_1120 (O_1120,N_14641,N_13593);
xor UO_1121 (O_1121,N_13270,N_12841);
xor UO_1122 (O_1122,N_12986,N_12005);
and UO_1123 (O_1123,N_14978,N_14051);
or UO_1124 (O_1124,N_12818,N_12989);
and UO_1125 (O_1125,N_14317,N_12438);
and UO_1126 (O_1126,N_13957,N_13367);
nor UO_1127 (O_1127,N_12115,N_14556);
xor UO_1128 (O_1128,N_14980,N_13034);
nor UO_1129 (O_1129,N_14368,N_13638);
or UO_1130 (O_1130,N_12322,N_14499);
nand UO_1131 (O_1131,N_13740,N_13965);
and UO_1132 (O_1132,N_12874,N_14316);
nor UO_1133 (O_1133,N_13753,N_12883);
nand UO_1134 (O_1134,N_14783,N_12907);
nand UO_1135 (O_1135,N_12998,N_12012);
nand UO_1136 (O_1136,N_14313,N_13980);
xor UO_1137 (O_1137,N_14502,N_12984);
or UO_1138 (O_1138,N_12265,N_12471);
nand UO_1139 (O_1139,N_12481,N_13869);
xor UO_1140 (O_1140,N_13959,N_13363);
and UO_1141 (O_1141,N_12292,N_13432);
nor UO_1142 (O_1142,N_13751,N_13440);
or UO_1143 (O_1143,N_13587,N_13460);
nor UO_1144 (O_1144,N_14260,N_12862);
xnor UO_1145 (O_1145,N_14662,N_14881);
nor UO_1146 (O_1146,N_13074,N_14773);
or UO_1147 (O_1147,N_14545,N_14182);
nor UO_1148 (O_1148,N_14294,N_14750);
and UO_1149 (O_1149,N_12690,N_12891);
nand UO_1150 (O_1150,N_12935,N_14805);
xnor UO_1151 (O_1151,N_13903,N_13115);
nand UO_1152 (O_1152,N_14351,N_12412);
nand UO_1153 (O_1153,N_14933,N_13928);
and UO_1154 (O_1154,N_14380,N_14608);
or UO_1155 (O_1155,N_12789,N_13413);
nand UO_1156 (O_1156,N_14563,N_13999);
xnor UO_1157 (O_1157,N_13872,N_13715);
or UO_1158 (O_1158,N_13843,N_13082);
and UO_1159 (O_1159,N_13817,N_14710);
nand UO_1160 (O_1160,N_14244,N_14589);
xnor UO_1161 (O_1161,N_13000,N_14138);
xor UO_1162 (O_1162,N_14665,N_14483);
or UO_1163 (O_1163,N_12485,N_14952);
and UO_1164 (O_1164,N_14504,N_12228);
nor UO_1165 (O_1165,N_13886,N_12806);
and UO_1166 (O_1166,N_12612,N_14065);
or UO_1167 (O_1167,N_13767,N_12206);
xor UO_1168 (O_1168,N_12072,N_13695);
xor UO_1169 (O_1169,N_13862,N_13414);
nand UO_1170 (O_1170,N_13613,N_14660);
nand UO_1171 (O_1171,N_13424,N_12399);
and UO_1172 (O_1172,N_14621,N_14543);
or UO_1173 (O_1173,N_13737,N_12521);
or UO_1174 (O_1174,N_12170,N_14484);
or UO_1175 (O_1175,N_14759,N_14603);
and UO_1176 (O_1176,N_12801,N_13483);
xor UO_1177 (O_1177,N_12939,N_12319);
xor UO_1178 (O_1178,N_12352,N_12664);
xnor UO_1179 (O_1179,N_13673,N_13427);
xor UO_1180 (O_1180,N_14027,N_12963);
nand UO_1181 (O_1181,N_12710,N_12037);
or UO_1182 (O_1182,N_13313,N_14251);
nand UO_1183 (O_1183,N_12203,N_14746);
nand UO_1184 (O_1184,N_13347,N_14836);
xor UO_1185 (O_1185,N_12694,N_13220);
or UO_1186 (O_1186,N_12439,N_14422);
and UO_1187 (O_1187,N_13467,N_12761);
and UO_1188 (O_1188,N_13160,N_12593);
xnor UO_1189 (O_1189,N_13393,N_12001);
nand UO_1190 (O_1190,N_13255,N_14703);
and UO_1191 (O_1191,N_14482,N_14992);
nor UO_1192 (O_1192,N_13900,N_13917);
nand UO_1193 (O_1193,N_13539,N_13981);
or UO_1194 (O_1194,N_12456,N_13545);
and UO_1195 (O_1195,N_12828,N_13444);
and UO_1196 (O_1196,N_12647,N_12609);
xnor UO_1197 (O_1197,N_14231,N_13659);
nor UO_1198 (O_1198,N_12996,N_13229);
nand UO_1199 (O_1199,N_13032,N_13787);
nor UO_1200 (O_1200,N_12575,N_12053);
and UO_1201 (O_1201,N_14958,N_13152);
and UO_1202 (O_1202,N_14464,N_14139);
nand UO_1203 (O_1203,N_13281,N_13923);
nor UO_1204 (O_1204,N_12516,N_13955);
nand UO_1205 (O_1205,N_12035,N_14867);
and UO_1206 (O_1206,N_12578,N_12538);
nor UO_1207 (O_1207,N_12423,N_12868);
xnor UO_1208 (O_1208,N_14198,N_12255);
and UO_1209 (O_1209,N_12875,N_14694);
nor UO_1210 (O_1210,N_12619,N_12507);
nor UO_1211 (O_1211,N_12602,N_14224);
xnor UO_1212 (O_1212,N_14128,N_14036);
and UO_1213 (O_1213,N_13636,N_12863);
xnor UO_1214 (O_1214,N_13250,N_13841);
nor UO_1215 (O_1215,N_14529,N_13827);
and UO_1216 (O_1216,N_12490,N_13406);
xor UO_1217 (O_1217,N_12351,N_13498);
and UO_1218 (O_1218,N_12805,N_13499);
nand UO_1219 (O_1219,N_12502,N_14602);
xnor UO_1220 (O_1220,N_14633,N_14446);
and UO_1221 (O_1221,N_14588,N_14613);
nand UO_1222 (O_1222,N_13632,N_14619);
nand UO_1223 (O_1223,N_14461,N_12087);
nor UO_1224 (O_1224,N_13744,N_13302);
and UO_1225 (O_1225,N_13039,N_14823);
and UO_1226 (O_1226,N_12678,N_13331);
nand UO_1227 (O_1227,N_12200,N_14693);
nand UO_1228 (O_1228,N_13939,N_13919);
xor UO_1229 (O_1229,N_13059,N_13947);
or UO_1230 (O_1230,N_12930,N_12597);
and UO_1231 (O_1231,N_14164,N_12635);
nand UO_1232 (O_1232,N_13252,N_12421);
nand UO_1233 (O_1233,N_14274,N_13885);
xnor UO_1234 (O_1234,N_14079,N_12474);
or UO_1235 (O_1235,N_14521,N_14887);
or UO_1236 (O_1236,N_13060,N_12782);
or UO_1237 (O_1237,N_13045,N_12162);
nand UO_1238 (O_1238,N_14405,N_14725);
nor UO_1239 (O_1239,N_14985,N_12092);
and UO_1240 (O_1240,N_14954,N_14601);
and UO_1241 (O_1241,N_13620,N_14620);
and UO_1242 (O_1242,N_14212,N_14936);
nand UO_1243 (O_1243,N_14288,N_14075);
nor UO_1244 (O_1244,N_12572,N_12275);
and UO_1245 (O_1245,N_12295,N_12760);
nand UO_1246 (O_1246,N_14771,N_12016);
or UO_1247 (O_1247,N_14147,N_14308);
xor UO_1248 (O_1248,N_12177,N_14067);
or UO_1249 (O_1249,N_14074,N_13524);
and UO_1250 (O_1250,N_14202,N_13030);
and UO_1251 (O_1251,N_13619,N_13671);
nor UO_1252 (O_1252,N_13050,N_13122);
xnor UO_1253 (O_1253,N_12605,N_13933);
nor UO_1254 (O_1254,N_13553,N_12125);
nand UO_1255 (O_1255,N_13263,N_12702);
and UO_1256 (O_1256,N_13782,N_12326);
nor UO_1257 (O_1257,N_13078,N_13595);
nand UO_1258 (O_1258,N_12990,N_13310);
or UO_1259 (O_1259,N_12788,N_13484);
or UO_1260 (O_1260,N_13952,N_12797);
nand UO_1261 (O_1261,N_12736,N_12286);
nor UO_1262 (O_1262,N_13531,N_14206);
and UO_1263 (O_1263,N_12278,N_12363);
or UO_1264 (O_1264,N_12066,N_13597);
and UO_1265 (O_1265,N_12031,N_14918);
xor UO_1266 (O_1266,N_13123,N_14283);
or UO_1267 (O_1267,N_12799,N_13339);
nand UO_1268 (O_1268,N_14611,N_12068);
and UO_1269 (O_1269,N_12529,N_12394);
or UO_1270 (O_1270,N_12937,N_14123);
or UO_1271 (O_1271,N_12090,N_14250);
and UO_1272 (O_1272,N_13650,N_14312);
nor UO_1273 (O_1273,N_12713,N_14686);
nand UO_1274 (O_1274,N_12195,N_12221);
or UO_1275 (O_1275,N_13948,N_12872);
xnor UO_1276 (O_1276,N_13603,N_14814);
and UO_1277 (O_1277,N_14682,N_13411);
and UO_1278 (O_1278,N_14324,N_14909);
nor UO_1279 (O_1279,N_14194,N_13297);
xnor UO_1280 (O_1280,N_14192,N_12519);
nand UO_1281 (O_1281,N_14364,N_12208);
nand UO_1282 (O_1282,N_14709,N_14195);
xnor UO_1283 (O_1283,N_14630,N_13311);
and UO_1284 (O_1284,N_13439,N_13558);
nand UO_1285 (O_1285,N_13995,N_13617);
or UO_1286 (O_1286,N_14598,N_13972);
or UO_1287 (O_1287,N_13024,N_12876);
xor UO_1288 (O_1288,N_13062,N_13988);
nor UO_1289 (O_1289,N_13902,N_14883);
and UO_1290 (O_1290,N_13293,N_13285);
nor UO_1291 (O_1291,N_12988,N_14208);
nand UO_1292 (O_1292,N_14942,N_13526);
nor UO_1293 (O_1293,N_13337,N_13590);
nand UO_1294 (O_1294,N_13236,N_14311);
xor UO_1295 (O_1295,N_13940,N_13681);
and UO_1296 (O_1296,N_14740,N_12159);
nor UO_1297 (O_1297,N_12836,N_13795);
xor UO_1298 (O_1298,N_12289,N_12902);
nand UO_1299 (O_1299,N_13217,N_13672);
nand UO_1300 (O_1300,N_12213,N_13776);
nand UO_1301 (O_1301,N_13568,N_13125);
nor UO_1302 (O_1302,N_13676,N_14628);
nand UO_1303 (O_1303,N_12738,N_12976);
nor UO_1304 (O_1304,N_13254,N_14657);
nand UO_1305 (O_1305,N_14217,N_14425);
nor UO_1306 (O_1306,N_12795,N_12056);
or UO_1307 (O_1307,N_13706,N_13877);
nor UO_1308 (O_1308,N_14266,N_12390);
nor UO_1309 (O_1309,N_12236,N_13726);
and UO_1310 (O_1310,N_14627,N_14780);
xor UO_1311 (O_1311,N_14145,N_13405);
and UO_1312 (O_1312,N_14367,N_13528);
xnor UO_1313 (O_1313,N_13918,N_14753);
and UO_1314 (O_1314,N_12936,N_14402);
xnor UO_1315 (O_1315,N_12522,N_13459);
nor UO_1316 (O_1316,N_13143,N_12804);
nand UO_1317 (O_1317,N_12013,N_12911);
nor UO_1318 (O_1318,N_14431,N_14920);
nand UO_1319 (O_1319,N_14129,N_14127);
nor UO_1320 (O_1320,N_12432,N_14807);
nor UO_1321 (O_1321,N_14235,N_14087);
nand UO_1322 (O_1322,N_13656,N_13019);
or UO_1323 (O_1323,N_13926,N_12246);
or UO_1324 (O_1324,N_14334,N_13865);
nor UO_1325 (O_1325,N_12961,N_14891);
xor UO_1326 (O_1326,N_14856,N_12480);
nor UO_1327 (O_1327,N_14456,N_14756);
nor UO_1328 (O_1328,N_14110,N_13559);
and UO_1329 (O_1329,N_13491,N_12188);
or UO_1330 (O_1330,N_12573,N_13851);
nand UO_1331 (O_1331,N_12682,N_13269);
xnor UO_1332 (O_1332,N_14053,N_14530);
and UO_1333 (O_1333,N_14674,N_12026);
and UO_1334 (O_1334,N_12182,N_12226);
nor UO_1335 (O_1335,N_12239,N_13321);
xnor UO_1336 (O_1336,N_13607,N_12565);
nand UO_1337 (O_1337,N_14986,N_14902);
xor UO_1338 (O_1338,N_13332,N_14864);
and UO_1339 (O_1339,N_13487,N_12336);
and UO_1340 (O_1340,N_13120,N_12024);
xor UO_1341 (O_1341,N_12685,N_13244);
xnor UO_1342 (O_1342,N_12334,N_14593);
or UO_1343 (O_1343,N_14101,N_14245);
xor UO_1344 (O_1344,N_13822,N_13731);
xnor UO_1345 (O_1345,N_13588,N_12036);
xnor UO_1346 (O_1346,N_13188,N_12662);
nand UO_1347 (O_1347,N_14924,N_12877);
or UO_1348 (O_1348,N_14117,N_14349);
nor UO_1349 (O_1349,N_13634,N_13150);
nand UO_1350 (O_1350,N_12518,N_13210);
nor UO_1351 (O_1351,N_14561,N_13894);
nor UO_1352 (O_1352,N_13100,N_14824);
nor UO_1353 (O_1353,N_14408,N_14196);
xor UO_1354 (O_1354,N_13502,N_12576);
nand UO_1355 (O_1355,N_14600,N_12256);
nor UO_1356 (O_1356,N_12823,N_13549);
xor UO_1357 (O_1357,N_12201,N_14059);
nor UO_1358 (O_1358,N_13665,N_12340);
xor UO_1359 (O_1359,N_13760,N_14361);
or UO_1360 (O_1360,N_12870,N_13729);
nor UO_1361 (O_1361,N_14741,N_12329);
nor UO_1362 (O_1362,N_12086,N_13689);
and UO_1363 (O_1363,N_14193,N_13407);
xor UO_1364 (O_1364,N_14786,N_14626);
nand UO_1365 (O_1365,N_12143,N_13680);
xnor UO_1366 (O_1366,N_13717,N_12746);
xor UO_1367 (O_1367,N_12927,N_12119);
and UO_1368 (O_1368,N_14168,N_14511);
or UO_1369 (O_1369,N_13501,N_13505);
nand UO_1370 (O_1370,N_12897,N_12082);
nand UO_1371 (O_1371,N_12774,N_12002);
or UO_1372 (O_1372,N_13167,N_12749);
or UO_1373 (O_1373,N_14738,N_14418);
nand UO_1374 (O_1374,N_12488,N_13099);
nand UO_1375 (O_1375,N_12701,N_14004);
or UO_1376 (O_1376,N_12411,N_12141);
or UO_1377 (O_1377,N_13685,N_14107);
xnor UO_1378 (O_1378,N_14513,N_13338);
nor UO_1379 (O_1379,N_12950,N_14171);
or UO_1380 (O_1380,N_12146,N_14955);
nor UO_1381 (O_1381,N_13606,N_13288);
nand UO_1382 (O_1382,N_13454,N_14879);
and UO_1383 (O_1383,N_13710,N_13639);
nor UO_1384 (O_1384,N_12878,N_14020);
or UO_1385 (O_1385,N_12040,N_13798);
nor UO_1386 (O_1386,N_13398,N_13128);
nand UO_1387 (O_1387,N_12073,N_12778);
and UO_1388 (O_1388,N_14797,N_13145);
xor UO_1389 (O_1389,N_12693,N_14066);
xnor UO_1390 (O_1390,N_12668,N_14802);
or UO_1391 (O_1391,N_13954,N_13852);
xnor UO_1392 (O_1392,N_12396,N_14799);
and UO_1393 (O_1393,N_13594,N_12307);
and UO_1394 (O_1394,N_12371,N_14314);
nand UO_1395 (O_1395,N_14028,N_14681);
nor UO_1396 (O_1396,N_14032,N_14963);
or UO_1397 (O_1397,N_13002,N_14086);
or UO_1398 (O_1398,N_12571,N_14595);
and UO_1399 (O_1399,N_13390,N_13734);
nand UO_1400 (O_1400,N_13040,N_13664);
and UO_1401 (O_1401,N_12444,N_13838);
and UO_1402 (O_1402,N_14187,N_14507);
xor UO_1403 (O_1403,N_13222,N_12853);
nand UO_1404 (O_1404,N_14745,N_12750);
and UO_1405 (O_1405,N_14754,N_14017);
nand UO_1406 (O_1406,N_14585,N_12533);
nor UO_1407 (O_1407,N_14501,N_12869);
or UO_1408 (O_1408,N_13295,N_12032);
xnor UO_1409 (O_1409,N_13772,N_14764);
or UO_1410 (O_1410,N_12194,N_14853);
nor UO_1411 (O_1411,N_14659,N_13683);
xnor UO_1412 (O_1412,N_14470,N_12492);
nor UO_1413 (O_1413,N_14599,N_12745);
nand UO_1414 (O_1414,N_12535,N_13307);
and UO_1415 (O_1415,N_14466,N_13574);
and UO_1416 (O_1416,N_14669,N_13548);
and UO_1417 (O_1417,N_14798,N_13193);
or UO_1418 (O_1418,N_12381,N_14829);
or UO_1419 (O_1419,N_14961,N_14755);
or UO_1420 (O_1420,N_12346,N_14579);
nand UO_1421 (O_1421,N_13237,N_14433);
nor UO_1422 (O_1422,N_12104,N_14651);
nor UO_1423 (O_1423,N_12557,N_14971);
or UO_1424 (O_1424,N_12077,N_13657);
and UO_1425 (O_1425,N_13819,N_12735);
and UO_1426 (O_1426,N_13629,N_14437);
xnor UO_1427 (O_1427,N_13765,N_14794);
nand UO_1428 (O_1428,N_14255,N_12924);
nand UO_1429 (O_1429,N_13175,N_12345);
or UO_1430 (O_1430,N_13089,N_13418);
nor UO_1431 (O_1431,N_12716,N_13242);
nor UO_1432 (O_1432,N_13758,N_13008);
and UO_1433 (O_1433,N_12793,N_12074);
and UO_1434 (O_1434,N_14635,N_13486);
xnor UO_1435 (O_1435,N_14358,N_14451);
xor UO_1436 (O_1436,N_12081,N_12524);
xor UO_1437 (O_1437,N_14022,N_12136);
nor UO_1438 (O_1438,N_12333,N_14706);
and UO_1439 (O_1439,N_12160,N_14514);
nand UO_1440 (O_1440,N_13256,N_12554);
xor UO_1441 (O_1441,N_12343,N_12367);
or UO_1442 (O_1442,N_14078,N_12606);
nor UO_1443 (O_1443,N_14815,N_14321);
and UO_1444 (O_1444,N_13658,N_14024);
or UO_1445 (O_1445,N_13932,N_12342);
nor UO_1446 (O_1446,N_14039,N_13211);
nor UO_1447 (O_1447,N_14103,N_12581);
nor UO_1448 (O_1448,N_14383,N_13303);
nand UO_1449 (O_1449,N_13458,N_13333);
nand UO_1450 (O_1450,N_12470,N_12627);
and UO_1451 (O_1451,N_14298,N_12070);
or UO_1452 (O_1452,N_14731,N_12149);
or UO_1453 (O_1453,N_14116,N_12734);
nand UO_1454 (O_1454,N_13341,N_13127);
nand UO_1455 (O_1455,N_13878,N_14005);
nor UO_1456 (O_1456,N_14100,N_14999);
xnor UO_1457 (O_1457,N_12614,N_14767);
xor UO_1458 (O_1458,N_13421,N_12303);
or UO_1459 (O_1459,N_13987,N_13802);
and UO_1460 (O_1460,N_12271,N_14023);
or UO_1461 (O_1461,N_13906,N_13299);
or UO_1462 (O_1462,N_12276,N_12277);
or UO_1463 (O_1463,N_13349,N_13048);
and UO_1464 (O_1464,N_14178,N_12112);
and UO_1465 (O_1465,N_13615,N_14427);
and UO_1466 (O_1466,N_14247,N_12530);
nand UO_1467 (O_1467,N_12487,N_12865);
nand UO_1468 (O_1468,N_12264,N_13447);
and UO_1469 (O_1469,N_14968,N_13474);
nand UO_1470 (O_1470,N_12331,N_12496);
nand UO_1471 (O_1471,N_12404,N_13292);
xor UO_1472 (O_1472,N_14558,N_13070);
xor UO_1473 (O_1473,N_14664,N_12696);
nor UO_1474 (O_1474,N_14211,N_12157);
or UO_1475 (O_1475,N_12142,N_13343);
xor UO_1476 (O_1476,N_12879,N_12720);
xor UO_1477 (O_1477,N_13521,N_13570);
or UO_1478 (O_1478,N_13373,N_13982);
nor UO_1479 (O_1479,N_13736,N_13063);
nor UO_1480 (O_1480,N_13912,N_13895);
xor UO_1481 (O_1481,N_14898,N_14597);
and UO_1482 (O_1482,N_14646,N_14760);
nand UO_1483 (O_1483,N_13108,N_14535);
and UO_1484 (O_1484,N_13086,N_13661);
xnor UO_1485 (O_1485,N_13733,N_12630);
or UO_1486 (O_1486,N_13113,N_12900);
and UO_1487 (O_1487,N_12707,N_13387);
nor UO_1488 (O_1488,N_12817,N_13004);
and UO_1489 (O_1489,N_14801,N_13761);
and UO_1490 (O_1490,N_13808,N_12175);
xnor UO_1491 (O_1491,N_13824,N_13922);
and UO_1492 (O_1492,N_14346,N_13330);
or UO_1493 (O_1493,N_13457,N_13732);
nand UO_1494 (O_1494,N_14811,N_12312);
xnor UO_1495 (O_1495,N_13420,N_14237);
or UO_1496 (O_1496,N_12473,N_12595);
or UO_1497 (O_1497,N_12374,N_13624);
nand UO_1498 (O_1498,N_12128,N_14001);
and UO_1499 (O_1499,N_12280,N_13249);
or UO_1500 (O_1500,N_12534,N_14404);
nand UO_1501 (O_1501,N_12277,N_14635);
nand UO_1502 (O_1502,N_12907,N_13875);
nand UO_1503 (O_1503,N_12890,N_12837);
xor UO_1504 (O_1504,N_14067,N_12463);
nand UO_1505 (O_1505,N_13505,N_12408);
nor UO_1506 (O_1506,N_14854,N_14992);
nand UO_1507 (O_1507,N_12126,N_12310);
and UO_1508 (O_1508,N_13618,N_13295);
nand UO_1509 (O_1509,N_14437,N_12658);
nand UO_1510 (O_1510,N_12827,N_13300);
xnor UO_1511 (O_1511,N_12088,N_12212);
and UO_1512 (O_1512,N_12099,N_13495);
or UO_1513 (O_1513,N_14782,N_12552);
nand UO_1514 (O_1514,N_12966,N_14398);
and UO_1515 (O_1515,N_12298,N_13434);
nand UO_1516 (O_1516,N_12385,N_14554);
nor UO_1517 (O_1517,N_14564,N_14740);
and UO_1518 (O_1518,N_12774,N_13786);
nor UO_1519 (O_1519,N_14903,N_14123);
nand UO_1520 (O_1520,N_12189,N_14750);
xor UO_1521 (O_1521,N_14049,N_14287);
nor UO_1522 (O_1522,N_12850,N_12481);
and UO_1523 (O_1523,N_14893,N_13729);
nor UO_1524 (O_1524,N_12903,N_12219);
xnor UO_1525 (O_1525,N_12047,N_14474);
nand UO_1526 (O_1526,N_13805,N_14170);
and UO_1527 (O_1527,N_13164,N_13910);
nor UO_1528 (O_1528,N_13915,N_14297);
and UO_1529 (O_1529,N_14993,N_14118);
nand UO_1530 (O_1530,N_13698,N_14797);
and UO_1531 (O_1531,N_12910,N_13356);
and UO_1532 (O_1532,N_13148,N_13152);
nor UO_1533 (O_1533,N_12863,N_13780);
xnor UO_1534 (O_1534,N_13905,N_12126);
and UO_1535 (O_1535,N_14484,N_12895);
nor UO_1536 (O_1536,N_12730,N_12800);
nand UO_1537 (O_1537,N_14988,N_12565);
or UO_1538 (O_1538,N_13521,N_12204);
xor UO_1539 (O_1539,N_12052,N_12445);
nand UO_1540 (O_1540,N_13364,N_13864);
xor UO_1541 (O_1541,N_12849,N_14670);
nor UO_1542 (O_1542,N_13194,N_14398);
or UO_1543 (O_1543,N_12723,N_14610);
nor UO_1544 (O_1544,N_13006,N_12684);
nor UO_1545 (O_1545,N_14616,N_13252);
xor UO_1546 (O_1546,N_13426,N_13476);
xnor UO_1547 (O_1547,N_12498,N_12178);
xnor UO_1548 (O_1548,N_14156,N_12939);
xnor UO_1549 (O_1549,N_14789,N_12895);
and UO_1550 (O_1550,N_14812,N_14932);
nor UO_1551 (O_1551,N_12433,N_14085);
and UO_1552 (O_1552,N_12282,N_12851);
xor UO_1553 (O_1553,N_13738,N_14808);
and UO_1554 (O_1554,N_14771,N_12931);
and UO_1555 (O_1555,N_12346,N_14768);
or UO_1556 (O_1556,N_12275,N_12957);
or UO_1557 (O_1557,N_12476,N_14848);
nor UO_1558 (O_1558,N_13346,N_14467);
nor UO_1559 (O_1559,N_13437,N_12246);
nand UO_1560 (O_1560,N_12222,N_13347);
xor UO_1561 (O_1561,N_13191,N_12735);
and UO_1562 (O_1562,N_12902,N_13924);
nand UO_1563 (O_1563,N_12463,N_14426);
or UO_1564 (O_1564,N_14335,N_12534);
nand UO_1565 (O_1565,N_14669,N_14605);
and UO_1566 (O_1566,N_14621,N_14167);
and UO_1567 (O_1567,N_12670,N_12087);
nand UO_1568 (O_1568,N_13718,N_13410);
xnor UO_1569 (O_1569,N_13000,N_12018);
nor UO_1570 (O_1570,N_12597,N_12153);
or UO_1571 (O_1571,N_13785,N_14467);
and UO_1572 (O_1572,N_12108,N_12964);
and UO_1573 (O_1573,N_13785,N_13125);
nand UO_1574 (O_1574,N_13366,N_14299);
and UO_1575 (O_1575,N_13957,N_14991);
nand UO_1576 (O_1576,N_12149,N_12036);
nand UO_1577 (O_1577,N_14308,N_13247);
nand UO_1578 (O_1578,N_12356,N_12161);
nor UO_1579 (O_1579,N_12515,N_13195);
nor UO_1580 (O_1580,N_12064,N_14343);
xnor UO_1581 (O_1581,N_13918,N_12335);
and UO_1582 (O_1582,N_14387,N_13322);
nand UO_1583 (O_1583,N_14986,N_13661);
nand UO_1584 (O_1584,N_14031,N_13117);
xnor UO_1585 (O_1585,N_12705,N_12702);
and UO_1586 (O_1586,N_14564,N_12603);
nor UO_1587 (O_1587,N_12213,N_14538);
or UO_1588 (O_1588,N_13853,N_14765);
or UO_1589 (O_1589,N_12120,N_13188);
or UO_1590 (O_1590,N_12401,N_13314);
and UO_1591 (O_1591,N_13725,N_13440);
xnor UO_1592 (O_1592,N_14972,N_13967);
xnor UO_1593 (O_1593,N_14127,N_13691);
nand UO_1594 (O_1594,N_13537,N_13482);
and UO_1595 (O_1595,N_14279,N_14585);
and UO_1596 (O_1596,N_14301,N_13727);
nand UO_1597 (O_1597,N_14754,N_14250);
and UO_1598 (O_1598,N_12794,N_14620);
or UO_1599 (O_1599,N_14162,N_12582);
nor UO_1600 (O_1600,N_13081,N_12658);
nand UO_1601 (O_1601,N_14405,N_13339);
and UO_1602 (O_1602,N_13714,N_12084);
nand UO_1603 (O_1603,N_14905,N_14153);
nand UO_1604 (O_1604,N_13243,N_14235);
or UO_1605 (O_1605,N_14729,N_14114);
xor UO_1606 (O_1606,N_14078,N_14677);
xor UO_1607 (O_1607,N_14755,N_13179);
nor UO_1608 (O_1608,N_13252,N_14056);
nand UO_1609 (O_1609,N_12930,N_12665);
or UO_1610 (O_1610,N_12813,N_13636);
xnor UO_1611 (O_1611,N_13536,N_13812);
xnor UO_1612 (O_1612,N_12369,N_12117);
nand UO_1613 (O_1613,N_12193,N_13749);
nor UO_1614 (O_1614,N_12634,N_13585);
or UO_1615 (O_1615,N_13503,N_13779);
nand UO_1616 (O_1616,N_13629,N_14517);
and UO_1617 (O_1617,N_14060,N_13589);
nor UO_1618 (O_1618,N_13471,N_12779);
nand UO_1619 (O_1619,N_14556,N_14119);
or UO_1620 (O_1620,N_14881,N_14537);
or UO_1621 (O_1621,N_12401,N_14086);
or UO_1622 (O_1622,N_14499,N_13386);
nor UO_1623 (O_1623,N_12224,N_12512);
xor UO_1624 (O_1624,N_12961,N_12750);
or UO_1625 (O_1625,N_14068,N_12706);
nor UO_1626 (O_1626,N_12512,N_13282);
nor UO_1627 (O_1627,N_12795,N_12745);
and UO_1628 (O_1628,N_13484,N_13286);
nand UO_1629 (O_1629,N_12392,N_12104);
nor UO_1630 (O_1630,N_12005,N_13815);
or UO_1631 (O_1631,N_14413,N_14156);
nand UO_1632 (O_1632,N_13979,N_12675);
xor UO_1633 (O_1633,N_13078,N_12821);
and UO_1634 (O_1634,N_13857,N_14778);
nand UO_1635 (O_1635,N_14440,N_14383);
xor UO_1636 (O_1636,N_14338,N_14450);
nand UO_1637 (O_1637,N_12551,N_13119);
or UO_1638 (O_1638,N_13063,N_14485);
and UO_1639 (O_1639,N_14204,N_14425);
nand UO_1640 (O_1640,N_12908,N_14617);
or UO_1641 (O_1641,N_13650,N_12107);
nand UO_1642 (O_1642,N_13951,N_14739);
xnor UO_1643 (O_1643,N_14995,N_13034);
nand UO_1644 (O_1644,N_12750,N_12615);
nand UO_1645 (O_1645,N_13031,N_12752);
nor UO_1646 (O_1646,N_14114,N_13882);
xnor UO_1647 (O_1647,N_12120,N_14670);
or UO_1648 (O_1648,N_12551,N_13223);
xnor UO_1649 (O_1649,N_12567,N_12007);
or UO_1650 (O_1650,N_13972,N_12643);
nor UO_1651 (O_1651,N_12210,N_14820);
nor UO_1652 (O_1652,N_12226,N_14465);
nor UO_1653 (O_1653,N_14940,N_14413);
nand UO_1654 (O_1654,N_13872,N_13831);
nand UO_1655 (O_1655,N_13995,N_12614);
nor UO_1656 (O_1656,N_14602,N_12419);
nand UO_1657 (O_1657,N_13201,N_12865);
xor UO_1658 (O_1658,N_12589,N_14710);
nor UO_1659 (O_1659,N_14196,N_14437);
nand UO_1660 (O_1660,N_12274,N_14169);
nor UO_1661 (O_1661,N_13537,N_14824);
or UO_1662 (O_1662,N_14917,N_14628);
nor UO_1663 (O_1663,N_13281,N_13948);
and UO_1664 (O_1664,N_12037,N_13907);
or UO_1665 (O_1665,N_14456,N_14722);
and UO_1666 (O_1666,N_12310,N_14778);
xnor UO_1667 (O_1667,N_13155,N_13270);
and UO_1668 (O_1668,N_12970,N_14723);
and UO_1669 (O_1669,N_12530,N_12833);
nor UO_1670 (O_1670,N_14963,N_12844);
nand UO_1671 (O_1671,N_12336,N_14909);
nand UO_1672 (O_1672,N_12576,N_14613);
or UO_1673 (O_1673,N_13484,N_14115);
nand UO_1674 (O_1674,N_13268,N_13181);
or UO_1675 (O_1675,N_14358,N_14398);
nand UO_1676 (O_1676,N_13565,N_12498);
xor UO_1677 (O_1677,N_12615,N_13754);
xor UO_1678 (O_1678,N_12872,N_14357);
nor UO_1679 (O_1679,N_14274,N_13864);
and UO_1680 (O_1680,N_12483,N_13157);
and UO_1681 (O_1681,N_12797,N_14287);
and UO_1682 (O_1682,N_12242,N_12434);
or UO_1683 (O_1683,N_12518,N_13798);
and UO_1684 (O_1684,N_12669,N_13997);
and UO_1685 (O_1685,N_12456,N_14611);
nor UO_1686 (O_1686,N_12689,N_13794);
nand UO_1687 (O_1687,N_14410,N_12757);
or UO_1688 (O_1688,N_14848,N_14914);
and UO_1689 (O_1689,N_12822,N_13949);
or UO_1690 (O_1690,N_13606,N_12417);
nor UO_1691 (O_1691,N_12197,N_13014);
nand UO_1692 (O_1692,N_12031,N_12904);
nor UO_1693 (O_1693,N_12448,N_12719);
nor UO_1694 (O_1694,N_14130,N_13947);
xnor UO_1695 (O_1695,N_13647,N_12423);
nor UO_1696 (O_1696,N_14643,N_14973);
nand UO_1697 (O_1697,N_14180,N_13528);
or UO_1698 (O_1698,N_12155,N_14763);
or UO_1699 (O_1699,N_12596,N_14618);
nor UO_1700 (O_1700,N_12519,N_12841);
nand UO_1701 (O_1701,N_13147,N_14529);
nor UO_1702 (O_1702,N_13154,N_12176);
and UO_1703 (O_1703,N_12095,N_14179);
nand UO_1704 (O_1704,N_13046,N_12339);
xnor UO_1705 (O_1705,N_13710,N_14345);
and UO_1706 (O_1706,N_14599,N_13140);
nand UO_1707 (O_1707,N_14742,N_13843);
xor UO_1708 (O_1708,N_14103,N_14079);
xnor UO_1709 (O_1709,N_12562,N_12600);
nor UO_1710 (O_1710,N_14583,N_12712);
and UO_1711 (O_1711,N_14188,N_13858);
and UO_1712 (O_1712,N_13541,N_14340);
xnor UO_1713 (O_1713,N_12013,N_13063);
and UO_1714 (O_1714,N_14545,N_13814);
and UO_1715 (O_1715,N_12800,N_14278);
or UO_1716 (O_1716,N_14784,N_14631);
nor UO_1717 (O_1717,N_14121,N_12807);
or UO_1718 (O_1718,N_13489,N_13911);
and UO_1719 (O_1719,N_13156,N_12103);
nand UO_1720 (O_1720,N_12480,N_14832);
nor UO_1721 (O_1721,N_14970,N_13601);
or UO_1722 (O_1722,N_13533,N_14703);
nor UO_1723 (O_1723,N_14543,N_14052);
nor UO_1724 (O_1724,N_12406,N_14632);
nor UO_1725 (O_1725,N_12692,N_13812);
xnor UO_1726 (O_1726,N_13905,N_12403);
and UO_1727 (O_1727,N_13201,N_13691);
nor UO_1728 (O_1728,N_13179,N_13164);
nand UO_1729 (O_1729,N_14114,N_12397);
or UO_1730 (O_1730,N_13311,N_12158);
xor UO_1731 (O_1731,N_12536,N_12119);
and UO_1732 (O_1732,N_13897,N_12794);
and UO_1733 (O_1733,N_12553,N_13475);
or UO_1734 (O_1734,N_12235,N_12568);
xor UO_1735 (O_1735,N_12176,N_14126);
nand UO_1736 (O_1736,N_13209,N_13067);
nor UO_1737 (O_1737,N_13722,N_13547);
nand UO_1738 (O_1738,N_12834,N_12447);
or UO_1739 (O_1739,N_12956,N_12944);
nor UO_1740 (O_1740,N_12365,N_13458);
nand UO_1741 (O_1741,N_13058,N_13017);
or UO_1742 (O_1742,N_14454,N_14203);
and UO_1743 (O_1743,N_13990,N_13952);
nor UO_1744 (O_1744,N_14859,N_14158);
nor UO_1745 (O_1745,N_13484,N_13806);
or UO_1746 (O_1746,N_13104,N_14070);
xor UO_1747 (O_1747,N_13451,N_12325);
and UO_1748 (O_1748,N_14477,N_12032);
nand UO_1749 (O_1749,N_12637,N_14968);
or UO_1750 (O_1750,N_13691,N_14994);
nor UO_1751 (O_1751,N_13820,N_13315);
or UO_1752 (O_1752,N_14878,N_13020);
nor UO_1753 (O_1753,N_13577,N_14921);
or UO_1754 (O_1754,N_12976,N_12900);
xor UO_1755 (O_1755,N_13196,N_13969);
nand UO_1756 (O_1756,N_14988,N_14564);
nor UO_1757 (O_1757,N_13664,N_13186);
nor UO_1758 (O_1758,N_12400,N_13771);
nand UO_1759 (O_1759,N_13217,N_12097);
and UO_1760 (O_1760,N_14167,N_13507);
nor UO_1761 (O_1761,N_14154,N_12482);
xnor UO_1762 (O_1762,N_13634,N_14672);
nand UO_1763 (O_1763,N_12350,N_14759);
and UO_1764 (O_1764,N_14895,N_14445);
nor UO_1765 (O_1765,N_12968,N_14207);
xnor UO_1766 (O_1766,N_12549,N_14442);
and UO_1767 (O_1767,N_14111,N_14681);
xor UO_1768 (O_1768,N_13245,N_14242);
and UO_1769 (O_1769,N_13750,N_14429);
xor UO_1770 (O_1770,N_13585,N_13688);
nand UO_1771 (O_1771,N_14978,N_13683);
and UO_1772 (O_1772,N_12263,N_13475);
nand UO_1773 (O_1773,N_12142,N_12103);
and UO_1774 (O_1774,N_13294,N_14750);
and UO_1775 (O_1775,N_12569,N_14251);
or UO_1776 (O_1776,N_14222,N_13849);
nand UO_1777 (O_1777,N_12660,N_14374);
nand UO_1778 (O_1778,N_14410,N_12392);
nand UO_1779 (O_1779,N_12619,N_12477);
nor UO_1780 (O_1780,N_14362,N_12943);
nand UO_1781 (O_1781,N_14926,N_14495);
nor UO_1782 (O_1782,N_12312,N_13349);
xnor UO_1783 (O_1783,N_13676,N_13899);
nor UO_1784 (O_1784,N_14169,N_13835);
nor UO_1785 (O_1785,N_14110,N_14051);
nand UO_1786 (O_1786,N_12298,N_13726);
or UO_1787 (O_1787,N_12298,N_13714);
nor UO_1788 (O_1788,N_14450,N_14052);
or UO_1789 (O_1789,N_14263,N_12197);
xnor UO_1790 (O_1790,N_14807,N_14234);
nor UO_1791 (O_1791,N_12789,N_14257);
or UO_1792 (O_1792,N_13189,N_14132);
nor UO_1793 (O_1793,N_12534,N_12684);
xnor UO_1794 (O_1794,N_14415,N_13814);
nand UO_1795 (O_1795,N_14921,N_14716);
or UO_1796 (O_1796,N_12668,N_13925);
nor UO_1797 (O_1797,N_14314,N_14890);
or UO_1798 (O_1798,N_14170,N_14535);
or UO_1799 (O_1799,N_14149,N_13475);
nor UO_1800 (O_1800,N_14500,N_14589);
and UO_1801 (O_1801,N_12896,N_12581);
and UO_1802 (O_1802,N_14252,N_14808);
nand UO_1803 (O_1803,N_13172,N_14014);
nor UO_1804 (O_1804,N_14287,N_14592);
or UO_1805 (O_1805,N_13745,N_13238);
nor UO_1806 (O_1806,N_13152,N_12032);
or UO_1807 (O_1807,N_14910,N_12719);
nand UO_1808 (O_1808,N_14680,N_14532);
xnor UO_1809 (O_1809,N_13149,N_14673);
or UO_1810 (O_1810,N_13948,N_12859);
or UO_1811 (O_1811,N_12479,N_14145);
or UO_1812 (O_1812,N_13835,N_13218);
or UO_1813 (O_1813,N_13655,N_13621);
xnor UO_1814 (O_1814,N_13084,N_13877);
and UO_1815 (O_1815,N_13350,N_13118);
xnor UO_1816 (O_1816,N_12221,N_14614);
xor UO_1817 (O_1817,N_14676,N_12442);
nand UO_1818 (O_1818,N_14336,N_14581);
or UO_1819 (O_1819,N_12751,N_14037);
or UO_1820 (O_1820,N_12286,N_12429);
and UO_1821 (O_1821,N_12340,N_12429);
and UO_1822 (O_1822,N_12654,N_12554);
xnor UO_1823 (O_1823,N_14727,N_12724);
xnor UO_1824 (O_1824,N_12881,N_14784);
xor UO_1825 (O_1825,N_14538,N_14728);
and UO_1826 (O_1826,N_12556,N_14997);
nor UO_1827 (O_1827,N_14586,N_13162);
xnor UO_1828 (O_1828,N_14919,N_14125);
nand UO_1829 (O_1829,N_13022,N_14695);
nand UO_1830 (O_1830,N_12711,N_13322);
and UO_1831 (O_1831,N_13249,N_13017);
xor UO_1832 (O_1832,N_12877,N_14740);
nor UO_1833 (O_1833,N_14321,N_12001);
or UO_1834 (O_1834,N_12212,N_12107);
nor UO_1835 (O_1835,N_12607,N_14051);
nor UO_1836 (O_1836,N_12148,N_14601);
or UO_1837 (O_1837,N_12373,N_13400);
nand UO_1838 (O_1838,N_12397,N_13124);
nor UO_1839 (O_1839,N_12428,N_12788);
nand UO_1840 (O_1840,N_13282,N_13934);
nand UO_1841 (O_1841,N_14508,N_14298);
xor UO_1842 (O_1842,N_13283,N_13906);
or UO_1843 (O_1843,N_12856,N_12958);
nor UO_1844 (O_1844,N_14995,N_13713);
nand UO_1845 (O_1845,N_14555,N_12584);
nand UO_1846 (O_1846,N_12959,N_13520);
and UO_1847 (O_1847,N_13686,N_13111);
and UO_1848 (O_1848,N_12995,N_13775);
or UO_1849 (O_1849,N_13558,N_13268);
and UO_1850 (O_1850,N_13339,N_14303);
and UO_1851 (O_1851,N_14728,N_14112);
nand UO_1852 (O_1852,N_14670,N_14923);
xnor UO_1853 (O_1853,N_13605,N_12308);
and UO_1854 (O_1854,N_14562,N_12814);
nand UO_1855 (O_1855,N_14693,N_13229);
and UO_1856 (O_1856,N_12971,N_14787);
nor UO_1857 (O_1857,N_13880,N_14601);
nor UO_1858 (O_1858,N_14457,N_14578);
xor UO_1859 (O_1859,N_14213,N_14353);
nand UO_1860 (O_1860,N_13584,N_13788);
and UO_1861 (O_1861,N_13627,N_13964);
and UO_1862 (O_1862,N_13623,N_12409);
or UO_1863 (O_1863,N_14147,N_12454);
and UO_1864 (O_1864,N_14678,N_12986);
nor UO_1865 (O_1865,N_14112,N_13106);
and UO_1866 (O_1866,N_13385,N_13854);
nand UO_1867 (O_1867,N_14188,N_13770);
or UO_1868 (O_1868,N_12015,N_12974);
or UO_1869 (O_1869,N_13822,N_13479);
nand UO_1870 (O_1870,N_14282,N_13768);
xor UO_1871 (O_1871,N_14853,N_12099);
xnor UO_1872 (O_1872,N_12513,N_12093);
or UO_1873 (O_1873,N_12608,N_14823);
nand UO_1874 (O_1874,N_12479,N_14858);
nand UO_1875 (O_1875,N_13010,N_12598);
or UO_1876 (O_1876,N_12000,N_12646);
and UO_1877 (O_1877,N_13289,N_14190);
nand UO_1878 (O_1878,N_13300,N_12482);
nor UO_1879 (O_1879,N_14504,N_12879);
xnor UO_1880 (O_1880,N_14130,N_13495);
and UO_1881 (O_1881,N_12906,N_14586);
nor UO_1882 (O_1882,N_13770,N_12823);
xor UO_1883 (O_1883,N_13271,N_12608);
or UO_1884 (O_1884,N_14824,N_13629);
nand UO_1885 (O_1885,N_12499,N_14212);
xor UO_1886 (O_1886,N_14928,N_13666);
or UO_1887 (O_1887,N_14051,N_14357);
and UO_1888 (O_1888,N_12618,N_12464);
nand UO_1889 (O_1889,N_13243,N_14358);
or UO_1890 (O_1890,N_12946,N_12091);
nand UO_1891 (O_1891,N_12622,N_14721);
or UO_1892 (O_1892,N_14819,N_14881);
nand UO_1893 (O_1893,N_14916,N_14667);
or UO_1894 (O_1894,N_14520,N_12498);
and UO_1895 (O_1895,N_12860,N_14084);
nor UO_1896 (O_1896,N_13768,N_13441);
and UO_1897 (O_1897,N_13868,N_13405);
nor UO_1898 (O_1898,N_14061,N_12086);
xor UO_1899 (O_1899,N_13052,N_13390);
nand UO_1900 (O_1900,N_12075,N_13008);
xor UO_1901 (O_1901,N_13448,N_14868);
xor UO_1902 (O_1902,N_12463,N_14869);
or UO_1903 (O_1903,N_12648,N_14498);
nor UO_1904 (O_1904,N_13179,N_12742);
xnor UO_1905 (O_1905,N_13188,N_13355);
and UO_1906 (O_1906,N_14092,N_14549);
nand UO_1907 (O_1907,N_14989,N_14367);
nor UO_1908 (O_1908,N_13673,N_13699);
and UO_1909 (O_1909,N_13130,N_12532);
xor UO_1910 (O_1910,N_12991,N_13871);
nand UO_1911 (O_1911,N_13021,N_14638);
nand UO_1912 (O_1912,N_14706,N_14508);
nor UO_1913 (O_1913,N_13213,N_12746);
xnor UO_1914 (O_1914,N_12385,N_12500);
and UO_1915 (O_1915,N_12003,N_14373);
or UO_1916 (O_1916,N_12796,N_13690);
or UO_1917 (O_1917,N_13665,N_12611);
or UO_1918 (O_1918,N_13224,N_12022);
and UO_1919 (O_1919,N_13222,N_12843);
nor UO_1920 (O_1920,N_12598,N_12420);
nor UO_1921 (O_1921,N_12963,N_13444);
nor UO_1922 (O_1922,N_13541,N_12081);
nand UO_1923 (O_1923,N_12182,N_14632);
nor UO_1924 (O_1924,N_13918,N_12229);
xnor UO_1925 (O_1925,N_14340,N_12302);
xor UO_1926 (O_1926,N_12539,N_13366);
nor UO_1927 (O_1927,N_12631,N_12061);
or UO_1928 (O_1928,N_14079,N_13972);
nor UO_1929 (O_1929,N_13822,N_13991);
nand UO_1930 (O_1930,N_12896,N_12546);
nand UO_1931 (O_1931,N_13661,N_12227);
nor UO_1932 (O_1932,N_12054,N_12156);
or UO_1933 (O_1933,N_13283,N_14814);
and UO_1934 (O_1934,N_12425,N_14280);
or UO_1935 (O_1935,N_12947,N_12337);
or UO_1936 (O_1936,N_12257,N_14500);
and UO_1937 (O_1937,N_12240,N_13026);
nand UO_1938 (O_1938,N_12314,N_13385);
and UO_1939 (O_1939,N_14077,N_13125);
and UO_1940 (O_1940,N_14567,N_14539);
or UO_1941 (O_1941,N_14670,N_13641);
nand UO_1942 (O_1942,N_12766,N_13627);
nand UO_1943 (O_1943,N_12715,N_13362);
nor UO_1944 (O_1944,N_13300,N_14593);
nand UO_1945 (O_1945,N_12261,N_14953);
nand UO_1946 (O_1946,N_13668,N_14662);
xor UO_1947 (O_1947,N_14657,N_14728);
nand UO_1948 (O_1948,N_12386,N_14772);
or UO_1949 (O_1949,N_12193,N_14736);
and UO_1950 (O_1950,N_12251,N_14415);
and UO_1951 (O_1951,N_12718,N_12213);
nand UO_1952 (O_1952,N_14052,N_12664);
nand UO_1953 (O_1953,N_12492,N_13913);
and UO_1954 (O_1954,N_13098,N_14560);
and UO_1955 (O_1955,N_14351,N_13935);
nor UO_1956 (O_1956,N_14108,N_14477);
and UO_1957 (O_1957,N_12788,N_12134);
xnor UO_1958 (O_1958,N_14237,N_14024);
nand UO_1959 (O_1959,N_12148,N_12167);
nor UO_1960 (O_1960,N_14802,N_12220);
xnor UO_1961 (O_1961,N_13857,N_13822);
nand UO_1962 (O_1962,N_13826,N_14330);
or UO_1963 (O_1963,N_12269,N_12355);
nor UO_1964 (O_1964,N_13518,N_14833);
or UO_1965 (O_1965,N_12721,N_14569);
or UO_1966 (O_1966,N_13440,N_13577);
nand UO_1967 (O_1967,N_14136,N_14917);
nand UO_1968 (O_1968,N_12101,N_13362);
nand UO_1969 (O_1969,N_12488,N_12490);
xor UO_1970 (O_1970,N_12120,N_13784);
nand UO_1971 (O_1971,N_13763,N_12511);
and UO_1972 (O_1972,N_12474,N_13768);
nor UO_1973 (O_1973,N_13031,N_14062);
nand UO_1974 (O_1974,N_13921,N_12479);
and UO_1975 (O_1975,N_12045,N_14821);
and UO_1976 (O_1976,N_12146,N_14900);
xor UO_1977 (O_1977,N_12821,N_12247);
nand UO_1978 (O_1978,N_12845,N_12979);
xnor UO_1979 (O_1979,N_12901,N_12310);
xnor UO_1980 (O_1980,N_12051,N_12203);
or UO_1981 (O_1981,N_13969,N_12055);
or UO_1982 (O_1982,N_13610,N_14120);
nor UO_1983 (O_1983,N_12487,N_12670);
nor UO_1984 (O_1984,N_14191,N_14568);
and UO_1985 (O_1985,N_13692,N_12612);
and UO_1986 (O_1986,N_13370,N_14713);
and UO_1987 (O_1987,N_12893,N_12915);
or UO_1988 (O_1988,N_12019,N_14927);
and UO_1989 (O_1989,N_12532,N_12484);
or UO_1990 (O_1990,N_13705,N_12137);
nand UO_1991 (O_1991,N_12213,N_13454);
xnor UO_1992 (O_1992,N_12756,N_14580);
nand UO_1993 (O_1993,N_13330,N_14849);
or UO_1994 (O_1994,N_13603,N_13442);
xor UO_1995 (O_1995,N_14343,N_12866);
xnor UO_1996 (O_1996,N_14442,N_12539);
nor UO_1997 (O_1997,N_13908,N_13789);
xor UO_1998 (O_1998,N_14723,N_14849);
nor UO_1999 (O_1999,N_12164,N_14464);
endmodule