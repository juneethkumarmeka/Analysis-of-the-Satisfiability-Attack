module basic_750_5000_1000_2_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2520,N_2522,N_2525,N_2526,N_2527,N_2529,N_2530,N_2531,N_2532,N_2534,N_2535,N_2536,N_2537,N_2539,N_2540,N_2541,N_2542,N_2543,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2552,N_2553,N_2555,N_2556,N_2557,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2585,N_2587,N_2588,N_2589,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2607,N_2608,N_2609,N_2610,N_2611,N_2613,N_2614,N_2617,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2626,N_2628,N_2630,N_2631,N_2634,N_2635,N_2636,N_2637,N_2638,N_2640,N_2641,N_2642,N_2644,N_2645,N_2648,N_2649,N_2650,N_2651,N_2653,N_2654,N_2655,N_2656,N_2658,N_2659,N_2660,N_2662,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2673,N_2674,N_2677,N_2678,N_2679,N_2682,N_2684,N_2685,N_2686,N_2687,N_2689,N_2690,N_2691,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2705,N_2706,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2730,N_2731,N_2732,N_2733,N_2734,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2748,N_2749,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2779,N_2781,N_2782,N_2783,N_2784,N_2785,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2806,N_2807,N_2809,N_2810,N_2811,N_2812,N_2813,N_2815,N_2818,N_2819,N_2820,N_2823,N_2824,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2833,N_2834,N_2835,N_2836,N_2837,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2852,N_2853,N_2855,N_2856,N_2858,N_2859,N_2860,N_2863,N_2864,N_2865,N_2867,N_2868,N_2870,N_2871,N_2872,N_2873,N_2874,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2884,N_2885,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2894,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2906,N_2907,N_2908,N_2909,N_2912,N_2913,N_2917,N_2918,N_2919,N_2921,N_2922,N_2924,N_2925,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2987,N_2988,N_2989,N_2990,N_2991,N_2993,N_2994,N_2995,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3052,N_3053,N_3055,N_3056,N_3058,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3073,N_3074,N_3075,N_3076,N_3078,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3092,N_3093,N_3094,N_3095,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3108,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3117,N_3118,N_3119,N_3120,N_3121,N_3124,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3146,N_3147,N_3148,N_3149,N_3151,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3163,N_3165,N_3166,N_3167,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3179,N_3181,N_3182,N_3185,N_3186,N_3189,N_3190,N_3191,N_3192,N_3193,N_3195,N_3196,N_3197,N_3200,N_3201,N_3202,N_3204,N_3207,N_3208,N_3210,N_3211,N_3212,N_3213,N_3215,N_3216,N_3217,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3231,N_3232,N_3233,N_3234,N_3236,N_3238,N_3239,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3249,N_3250,N_3252,N_3253,N_3254,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3276,N_3277,N_3279,N_3280,N_3282,N_3283,N_3284,N_3285,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3310,N_3311,N_3312,N_3313,N_3314,N_3316,N_3319,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3334,N_3335,N_3336,N_3337,N_3338,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3350,N_3351,N_3355,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3374,N_3375,N_3376,N_3378,N_3381,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3391,N_3392,N_3393,N_3394,N_3395,N_3397,N_3398,N_3400,N_3401,N_3403,N_3405,N_3406,N_3408,N_3409,N_3410,N_3411,N_3413,N_3414,N_3416,N_3417,N_3418,N_3419,N_3420,N_3423,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3438,N_3439,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3452,N_3453,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3477,N_3479,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3493,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3504,N_3505,N_3506,N_3508,N_3509,N_3510,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3527,N_3528,N_3529,N_3531,N_3532,N_3533,N_3535,N_3536,N_3537,N_3539,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3557,N_3560,N_3562,N_3564,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3579,N_3580,N_3581,N_3583,N_3584,N_3585,N_3588,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3677,N_3678,N_3679,N_3682,N_3683,N_3685,N_3686,N_3688,N_3689,N_3690,N_3691,N_3693,N_3694,N_3695,N_3696,N_3697,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3711,N_3712,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3742,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3769,N_3770,N_3771,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3781,N_3782,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3791,N_3792,N_3793,N_3794,N_3796,N_3797,N_3799,N_3800,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3823,N_3824,N_3825,N_3827,N_3828,N_3830,N_3832,N_3833,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3846,N_3848,N_3849,N_3850,N_3853,N_3855,N_3856,N_3857,N_3858,N_3859,N_3861,N_3862,N_3863,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3873,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3892,N_3893,N_3894,N_3895,N_3897,N_3899,N_3900,N_3902,N_3904,N_3908,N_3909,N_3910,N_3911,N_3912,N_3914,N_3915,N_3916,N_3918,N_3920,N_3921,N_3922,N_3923,N_3924,N_3926,N_3927,N_3928,N_3929,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3943,N_3944,N_3945,N_3946,N_3948,N_3949,N_3950,N_3952,N_3953,N_3954,N_3956,N_3958,N_3959,N_3960,N_3963,N_3965,N_3966,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3977,N_3978,N_3979,N_3980,N_3982,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3991,N_3992,N_3993,N_3994,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4005,N_4006,N_4007,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4027,N_4028,N_4030,N_4032,N_4033,N_4035,N_4036,N_4038,N_4039,N_4040,N_4042,N_4043,N_4044,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4053,N_4054,N_4055,N_4056,N_4057,N_4059,N_4060,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4076,N_4077,N_4078,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4097,N_4099,N_4100,N_4101,N_4103,N_4104,N_4105,N_4107,N_4109,N_4110,N_4111,N_4112,N_4113,N_4115,N_4116,N_4118,N_4119,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4134,N_4135,N_4136,N_4137,N_4139,N_4140,N_4141,N_4142,N_4143,N_4145,N_4148,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4160,N_4161,N_4162,N_4163,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4196,N_4198,N_4199,N_4201,N_4202,N_4203,N_4204,N_4205,N_4207,N_4208,N_4210,N_4211,N_4212,N_4215,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4227,N_4228,N_4229,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4267,N_4268,N_4269,N_4270,N_4272,N_4273,N_4274,N_4276,N_4277,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4287,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4298,N_4301,N_4303,N_4304,N_4305,N_4307,N_4308,N_4309,N_4311,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4332,N_4333,N_4334,N_4336,N_4337,N_4338,N_4339,N_4342,N_4344,N_4345,N_4346,N_4348,N_4350,N_4351,N_4352,N_4353,N_4355,N_4356,N_4358,N_4359,N_4360,N_4362,N_4363,N_4365,N_4366,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4383,N_4384,N_4385,N_4386,N_4389,N_4390,N_4391,N_4392,N_4393,N_4395,N_4397,N_4398,N_4400,N_4401,N_4402,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4414,N_4415,N_4416,N_4418,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4447,N_4448,N_4449,N_4450,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4460,N_4461,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4470,N_4471,N_4472,N_4473,N_4475,N_4477,N_4478,N_4479,N_4480,N_4482,N_4483,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4496,N_4498,N_4499,N_4501,N_4502,N_4503,N_4505,N_4506,N_4507,N_4509,N_4510,N_4511,N_4512,N_4516,N_4517,N_4518,N_4520,N_4522,N_4523,N_4524,N_4525,N_4526,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4548,N_4549,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4572,N_4574,N_4575,N_4576,N_4577,N_4578,N_4580,N_4581,N_4583,N_4584,N_4585,N_4586,N_4588,N_4590,N_4592,N_4593,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4605,N_4606,N_4607,N_4608,N_4610,N_4611,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4636,N_4638,N_4639,N_4640,N_4641,N_4642,N_4644,N_4647,N_4648,N_4650,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4661,N_4662,N_4664,N_4666,N_4667,N_4668,N_4672,N_4673,N_4674,N_4675,N_4676,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4692,N_4693,N_4694,N_4696,N_4697,N_4699,N_4700,N_4701,N_4702,N_4704,N_4705,N_4706,N_4707,N_4709,N_4711,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4743,N_4744,N_4745,N_4746,N_4748,N_4749,N_4750,N_4752,N_4753,N_4754,N_4755,N_4758,N_4759,N_4760,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4779,N_4780,N_4781,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4808,N_4809,N_4811,N_4812,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4822,N_4823,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4834,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4864,N_4866,N_4867,N_4868,N_4869,N_4870,N_4872,N_4873,N_4875,N_4876,N_4878,N_4879,N_4881,N_4882,N_4883,N_4884,N_4885,N_4887,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4898,N_4899,N_4900,N_4901,N_4902,N_4904,N_4905,N_4907,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4935,N_4936,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4968,N_4969,N_4972,N_4973,N_4974,N_4976,N_4977,N_4978,N_4982,N_4983,N_4984,N_4985,N_4987,N_4988,N_4989,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_378,In_386);
and U1 (N_1,In_690,In_650);
nand U2 (N_2,In_583,In_248);
or U3 (N_3,In_548,In_568);
or U4 (N_4,In_192,In_246);
xnor U5 (N_5,In_534,In_12);
nand U6 (N_6,In_405,In_197);
and U7 (N_7,In_418,In_586);
nand U8 (N_8,In_183,In_210);
or U9 (N_9,In_116,In_440);
nand U10 (N_10,In_654,In_622);
xor U11 (N_11,In_279,In_656);
xor U12 (N_12,In_642,In_708);
nand U13 (N_13,In_265,In_610);
and U14 (N_14,In_659,In_446);
nor U15 (N_15,In_312,In_663);
or U16 (N_16,In_571,In_67);
xor U17 (N_17,In_83,In_53);
xor U18 (N_18,In_219,In_303);
nor U19 (N_19,In_614,In_481);
xnor U20 (N_20,In_124,In_19);
and U21 (N_21,In_304,In_676);
and U22 (N_22,In_422,In_531);
nor U23 (N_23,In_218,In_747);
xnor U24 (N_24,In_383,In_213);
xnor U25 (N_25,In_742,In_193);
nand U26 (N_26,In_289,In_229);
or U27 (N_27,In_287,In_117);
nor U28 (N_28,In_703,In_662);
or U29 (N_29,In_370,In_371);
and U30 (N_30,In_221,In_484);
and U31 (N_31,In_477,In_189);
and U32 (N_32,In_11,In_724);
and U33 (N_33,In_273,In_665);
or U34 (N_34,In_206,In_627);
xnor U35 (N_35,In_329,In_224);
nand U36 (N_36,In_630,In_558);
nor U37 (N_37,In_466,In_731);
or U38 (N_38,In_14,In_403);
xor U39 (N_39,In_98,In_309);
nand U40 (N_40,In_290,In_156);
and U41 (N_41,In_328,In_138);
nand U42 (N_42,In_150,In_260);
nand U43 (N_43,In_283,In_575);
and U44 (N_44,In_305,In_331);
nand U45 (N_45,In_672,In_175);
or U46 (N_46,In_31,In_400);
or U47 (N_47,In_508,In_23);
nor U48 (N_48,In_443,In_174);
and U49 (N_49,In_85,In_164);
xor U50 (N_50,In_638,In_486);
and U51 (N_51,In_306,In_651);
nor U52 (N_52,In_130,In_566);
or U53 (N_53,In_66,In_626);
and U54 (N_54,In_748,In_122);
xnor U55 (N_55,In_38,In_373);
or U56 (N_56,In_216,In_295);
xor U57 (N_57,In_608,In_467);
nor U58 (N_58,In_511,In_611);
xor U59 (N_59,In_255,In_345);
xnor U60 (N_60,In_453,In_40);
nand U61 (N_61,In_41,In_4);
xor U62 (N_62,In_700,In_445);
nand U63 (N_63,In_101,In_570);
nor U64 (N_64,In_252,In_71);
nor U65 (N_65,In_518,In_18);
and U66 (N_66,In_177,In_103);
or U67 (N_67,In_93,In_44);
and U68 (N_68,In_264,In_152);
nor U69 (N_69,In_498,In_173);
or U70 (N_70,In_390,In_408);
and U71 (N_71,In_320,In_491);
and U72 (N_72,In_186,In_104);
or U73 (N_73,In_687,In_431);
nor U74 (N_74,In_8,In_119);
nor U75 (N_75,In_313,In_109);
xnor U76 (N_76,In_182,In_27);
and U77 (N_77,In_494,In_121);
and U78 (N_78,In_190,In_576);
nand U79 (N_79,In_314,In_726);
xor U80 (N_80,In_348,In_513);
and U81 (N_81,In_679,In_427);
xnor U82 (N_82,In_298,In_161);
nand U83 (N_83,In_459,In_17);
and U84 (N_84,In_384,In_195);
nor U85 (N_85,In_238,In_424);
nand U86 (N_86,In_244,In_222);
or U87 (N_87,In_358,In_392);
nand U88 (N_88,In_205,In_158);
xor U89 (N_89,In_135,In_52);
or U90 (N_90,In_520,In_455);
or U91 (N_91,In_664,In_737);
nand U92 (N_92,In_73,In_151);
or U93 (N_93,In_556,In_354);
nor U94 (N_94,In_202,In_507);
nor U95 (N_95,In_465,In_214);
nand U96 (N_96,In_68,In_670);
or U97 (N_97,In_648,In_375);
and U98 (N_98,In_167,In_426);
xor U99 (N_99,In_74,In_624);
xor U100 (N_100,In_585,In_30);
xor U101 (N_101,In_569,In_634);
and U102 (N_102,In_263,In_284);
and U103 (N_103,In_510,In_154);
nor U104 (N_104,In_474,In_419);
or U105 (N_105,In_269,In_363);
and U106 (N_106,In_613,In_712);
nand U107 (N_107,In_734,In_172);
xor U108 (N_108,In_646,In_729);
nor U109 (N_109,In_685,In_645);
nand U110 (N_110,In_538,In_357);
and U111 (N_111,In_521,In_155);
and U112 (N_112,In_318,In_744);
nor U113 (N_113,In_524,In_6);
xor U114 (N_114,In_594,In_48);
nand U115 (N_115,In_230,In_153);
or U116 (N_116,In_452,In_26);
xor U117 (N_117,In_24,In_165);
xor U118 (N_118,In_675,In_87);
nand U119 (N_119,In_159,In_526);
nor U120 (N_120,In_573,In_515);
or U121 (N_121,In_63,In_547);
and U122 (N_122,In_69,In_535);
nand U123 (N_123,In_251,In_361);
and U124 (N_124,In_90,In_62);
or U125 (N_125,In_188,In_274);
nor U126 (N_126,In_652,In_128);
and U127 (N_127,In_557,In_201);
or U128 (N_128,In_315,In_641);
xor U129 (N_129,In_564,In_36);
nand U130 (N_130,In_442,In_285);
nor U131 (N_131,In_721,In_533);
xnor U132 (N_132,In_550,In_198);
xor U133 (N_133,In_497,In_559);
xnor U134 (N_134,In_15,In_432);
nor U135 (N_135,In_34,In_522);
nor U136 (N_136,In_364,In_257);
and U137 (N_137,In_606,In_407);
xnor U138 (N_138,In_79,In_503);
xor U139 (N_139,In_458,In_242);
nand U140 (N_140,In_730,In_292);
nor U141 (N_141,In_187,In_323);
or U142 (N_142,In_65,In_447);
or U143 (N_143,In_61,In_324);
and U144 (N_144,In_243,In_462);
and U145 (N_145,In_204,In_341);
xor U146 (N_146,In_72,In_359);
or U147 (N_147,In_655,In_728);
nand U148 (N_148,In_369,In_59);
and U149 (N_149,In_625,In_636);
xor U150 (N_150,In_338,In_600);
nand U151 (N_151,In_719,In_232);
nor U152 (N_152,In_411,In_179);
nand U153 (N_153,In_683,In_668);
nand U154 (N_154,In_249,In_723);
xor U155 (N_155,In_565,In_438);
nand U156 (N_156,In_226,In_60);
and U157 (N_157,In_166,In_220);
and U158 (N_158,In_108,In_247);
xor U159 (N_159,In_605,In_615);
or U160 (N_160,In_170,In_391);
xor U161 (N_161,In_28,In_302);
nand U162 (N_162,In_563,In_333);
nand U163 (N_163,In_32,In_346);
nand U164 (N_164,In_591,In_393);
or U165 (N_165,In_653,In_335);
nand U166 (N_166,In_114,In_682);
or U167 (N_167,In_476,In_94);
nor U168 (N_168,In_696,In_560);
nor U169 (N_169,In_82,In_437);
xnor U170 (N_170,In_543,In_29);
nor U171 (N_171,In_529,In_326);
and U172 (N_172,In_102,In_643);
xor U173 (N_173,In_80,In_25);
xor U174 (N_174,In_480,In_372);
nand U175 (N_175,In_532,In_711);
xor U176 (N_176,In_123,In_640);
xor U177 (N_177,In_301,In_196);
nand U178 (N_178,In_612,In_350);
or U179 (N_179,In_381,In_322);
xnor U180 (N_180,In_0,In_506);
and U181 (N_181,In_496,In_250);
or U182 (N_182,In_537,In_512);
and U183 (N_183,In_546,In_554);
or U184 (N_184,In_635,In_176);
or U185 (N_185,In_46,In_293);
nand U186 (N_186,In_578,In_344);
nor U187 (N_187,In_110,In_592);
nor U188 (N_188,In_401,In_549);
nor U189 (N_189,In_347,In_96);
nor U190 (N_190,In_297,In_42);
or U191 (N_191,In_542,In_144);
and U192 (N_192,In_516,In_727);
or U193 (N_193,In_572,In_581);
or U194 (N_194,In_689,In_236);
nor U195 (N_195,In_146,In_310);
nand U196 (N_196,In_275,In_291);
nand U197 (N_197,In_50,In_413);
nand U198 (N_198,In_436,In_749);
nor U199 (N_199,In_541,In_16);
xnor U200 (N_200,In_715,In_261);
nand U201 (N_201,In_81,In_178);
xnor U202 (N_202,In_136,In_409);
and U203 (N_203,In_268,In_10);
xnor U204 (N_204,In_661,In_701);
nand U205 (N_205,In_502,In_430);
xor U206 (N_206,In_389,In_368);
nor U207 (N_207,In_688,In_595);
nor U208 (N_208,In_330,In_589);
nand U209 (N_209,In_92,In_417);
nand U210 (N_210,In_362,In_351);
nand U211 (N_211,In_332,In_396);
or U212 (N_212,In_253,In_134);
nor U213 (N_213,In_735,In_658);
and U214 (N_214,In_262,In_519);
nor U215 (N_215,In_716,In_468);
nor U216 (N_216,In_91,In_399);
nand U217 (N_217,In_514,In_698);
and U218 (N_218,In_428,In_105);
xnor U219 (N_219,In_20,In_551);
nand U220 (N_220,In_470,In_340);
nor U221 (N_221,In_717,In_609);
and U222 (N_222,In_596,In_464);
nor U223 (N_223,In_709,In_601);
and U224 (N_224,In_603,In_131);
or U225 (N_225,In_695,In_483);
and U226 (N_226,In_147,In_412);
nor U227 (N_227,In_281,In_523);
or U228 (N_228,In_597,In_686);
xnor U229 (N_229,In_233,In_528);
nor U230 (N_230,In_37,In_671);
nand U231 (N_231,In_200,In_713);
and U232 (N_232,In_540,In_317);
xor U233 (N_233,In_78,In_120);
or U234 (N_234,In_492,In_420);
nand U235 (N_235,In_75,In_544);
xnor U236 (N_236,In_142,In_241);
nand U237 (N_237,In_379,In_223);
and U238 (N_238,In_89,In_617);
or U239 (N_239,In_501,In_725);
and U240 (N_240,In_272,In_194);
nor U241 (N_241,In_618,In_423);
nand U242 (N_242,In_527,In_148);
or U243 (N_243,In_582,In_3);
or U244 (N_244,In_574,In_334);
nand U245 (N_245,In_212,In_580);
nor U246 (N_246,In_111,In_509);
xnor U247 (N_247,In_681,In_140);
and U248 (N_248,In_308,In_479);
nand U249 (N_249,In_504,In_235);
xnor U250 (N_250,In_33,In_282);
and U251 (N_251,In_217,In_180);
nand U252 (N_252,In_337,In_215);
or U253 (N_253,In_705,In_660);
nand U254 (N_254,In_402,In_95);
nor U255 (N_255,In_450,In_694);
and U256 (N_256,In_410,In_145);
or U257 (N_257,In_499,In_181);
xnor U258 (N_258,In_739,In_118);
nor U259 (N_259,In_21,In_552);
nand U260 (N_260,In_394,In_395);
or U261 (N_261,In_536,In_86);
xor U262 (N_262,In_133,In_444);
nand U263 (N_263,In_633,In_84);
xnor U264 (N_264,In_632,In_457);
and U265 (N_265,In_674,In_49);
nor U266 (N_266,In_398,In_441);
xnor U267 (N_267,In_129,In_307);
nor U268 (N_268,In_294,In_456);
xor U269 (N_269,In_628,In_157);
xnor U270 (N_270,In_245,In_397);
xor U271 (N_271,In_266,In_143);
or U272 (N_272,In_404,In_746);
nand U273 (N_273,In_277,In_460);
or U274 (N_274,In_590,In_316);
and U275 (N_275,In_382,In_487);
nand U276 (N_276,In_692,In_355);
xnor U277 (N_277,In_593,In_475);
nor U278 (N_278,In_619,In_22);
nor U279 (N_279,In_228,In_599);
or U280 (N_280,In_488,In_184);
or U281 (N_281,In_714,In_691);
or U282 (N_282,In_132,In_607);
or U283 (N_283,In_677,In_139);
xor U284 (N_284,In_718,In_288);
nand U285 (N_285,In_525,In_360);
nand U286 (N_286,In_448,In_299);
or U287 (N_287,In_1,In_207);
nand U288 (N_288,In_141,In_163);
and U289 (N_289,In_325,In_352);
or U290 (N_290,In_342,In_740);
and U291 (N_291,In_616,In_58);
nand U292 (N_292,In_168,In_254);
xor U293 (N_293,In_657,In_267);
nor U294 (N_294,In_620,In_738);
nor U295 (N_295,In_39,In_602);
nor U296 (N_296,In_587,In_493);
and U297 (N_297,In_225,In_505);
and U298 (N_298,In_271,In_545);
and U299 (N_299,In_227,In_300);
and U300 (N_300,In_639,In_473);
or U301 (N_301,In_259,In_349);
xor U302 (N_302,In_421,In_45);
nand U303 (N_303,In_644,In_97);
nand U304 (N_304,In_647,In_100);
nand U305 (N_305,In_743,In_490);
xor U306 (N_306,In_240,In_598);
nand U307 (N_307,In_365,In_380);
nand U308 (N_308,In_171,In_678);
or U309 (N_309,In_667,In_489);
nor U310 (N_310,In_673,In_35);
nor U311 (N_311,In_234,In_669);
or U312 (N_312,In_706,In_9);
xnor U313 (N_313,In_343,In_339);
nor U314 (N_314,In_736,In_629);
and U315 (N_315,In_693,In_149);
nand U316 (N_316,In_461,In_54);
nand U317 (N_317,In_454,In_366);
nor U318 (N_318,In_435,In_374);
xnor U319 (N_319,In_621,In_732);
xnor U320 (N_320,In_680,In_463);
or U321 (N_321,In_43,In_433);
or U322 (N_322,In_162,In_115);
nor U323 (N_323,In_126,In_296);
xor U324 (N_324,In_562,In_406);
or U325 (N_325,In_745,In_185);
nand U326 (N_326,In_127,In_649);
nand U327 (N_327,In_485,In_137);
or U328 (N_328,In_449,In_414);
nand U329 (N_329,In_702,In_107);
nand U330 (N_330,In_631,In_57);
nor U331 (N_331,In_704,In_353);
nand U332 (N_332,In_697,In_482);
nor U333 (N_333,In_707,In_434);
nor U334 (N_334,In_203,In_385);
xor U335 (N_335,In_319,In_553);
or U336 (N_336,In_555,In_106);
xor U337 (N_337,In_577,In_64);
and U338 (N_338,In_720,In_425);
xor U339 (N_339,In_211,In_256);
nor U340 (N_340,In_567,In_270);
nand U341 (N_341,In_561,In_377);
or U342 (N_342,In_336,In_416);
xor U343 (N_343,In_7,In_699);
xor U344 (N_344,In_112,In_70);
xnor U345 (N_345,In_579,In_286);
nor U346 (N_346,In_666,In_231);
xor U347 (N_347,In_47,In_51);
nor U348 (N_348,In_77,In_495);
nand U349 (N_349,In_710,In_280);
nor U350 (N_350,In_517,In_623);
nand U351 (N_351,In_88,In_327);
xnor U352 (N_352,In_539,In_13);
xnor U353 (N_353,In_471,In_478);
nor U354 (N_354,In_169,In_604);
xnor U355 (N_355,In_278,In_208);
xnor U356 (N_356,In_191,In_2);
xnor U357 (N_357,In_367,In_55);
nor U358 (N_358,In_500,In_469);
nor U359 (N_359,In_741,In_588);
nor U360 (N_360,In_113,In_388);
nand U361 (N_361,In_733,In_722);
nand U362 (N_362,In_584,In_56);
nor U363 (N_363,In_276,In_209);
nor U364 (N_364,In_637,In_199);
nand U365 (N_365,In_451,In_684);
and U366 (N_366,In_356,In_387);
and U367 (N_367,In_76,In_99);
xor U368 (N_368,In_530,In_376);
nor U369 (N_369,In_239,In_439);
nand U370 (N_370,In_429,In_321);
nor U371 (N_371,In_160,In_472);
nor U372 (N_372,In_5,In_258);
or U373 (N_373,In_415,In_125);
and U374 (N_374,In_237,In_311);
nor U375 (N_375,In_20,In_268);
and U376 (N_376,In_585,In_522);
xor U377 (N_377,In_512,In_547);
nand U378 (N_378,In_624,In_725);
nor U379 (N_379,In_343,In_84);
nor U380 (N_380,In_504,In_392);
xor U381 (N_381,In_543,In_747);
xor U382 (N_382,In_272,In_371);
and U383 (N_383,In_95,In_236);
xor U384 (N_384,In_449,In_532);
nor U385 (N_385,In_457,In_728);
or U386 (N_386,In_501,In_318);
nand U387 (N_387,In_456,In_749);
or U388 (N_388,In_541,In_147);
and U389 (N_389,In_652,In_430);
or U390 (N_390,In_140,In_304);
nor U391 (N_391,In_538,In_580);
and U392 (N_392,In_527,In_302);
or U393 (N_393,In_320,In_522);
xnor U394 (N_394,In_616,In_370);
nand U395 (N_395,In_253,In_672);
nor U396 (N_396,In_186,In_744);
nand U397 (N_397,In_732,In_642);
nand U398 (N_398,In_740,In_429);
nor U399 (N_399,In_700,In_486);
nor U400 (N_400,In_607,In_328);
nor U401 (N_401,In_239,In_690);
xnor U402 (N_402,In_414,In_318);
and U403 (N_403,In_299,In_469);
or U404 (N_404,In_3,In_259);
xor U405 (N_405,In_571,In_736);
and U406 (N_406,In_565,In_687);
and U407 (N_407,In_502,In_714);
or U408 (N_408,In_747,In_345);
xnor U409 (N_409,In_80,In_370);
and U410 (N_410,In_101,In_704);
or U411 (N_411,In_672,In_294);
nand U412 (N_412,In_640,In_369);
nand U413 (N_413,In_279,In_672);
nor U414 (N_414,In_539,In_497);
nor U415 (N_415,In_549,In_370);
or U416 (N_416,In_253,In_426);
or U417 (N_417,In_363,In_672);
nand U418 (N_418,In_441,In_492);
xor U419 (N_419,In_19,In_449);
and U420 (N_420,In_483,In_318);
xnor U421 (N_421,In_186,In_383);
or U422 (N_422,In_525,In_60);
nor U423 (N_423,In_352,In_249);
nor U424 (N_424,In_51,In_423);
xnor U425 (N_425,In_596,In_409);
and U426 (N_426,In_485,In_128);
or U427 (N_427,In_301,In_572);
nor U428 (N_428,In_297,In_664);
and U429 (N_429,In_715,In_7);
nand U430 (N_430,In_302,In_741);
and U431 (N_431,In_659,In_301);
or U432 (N_432,In_749,In_435);
xor U433 (N_433,In_441,In_256);
and U434 (N_434,In_544,In_557);
nor U435 (N_435,In_461,In_706);
or U436 (N_436,In_36,In_701);
xor U437 (N_437,In_476,In_722);
nand U438 (N_438,In_136,In_168);
or U439 (N_439,In_262,In_528);
nor U440 (N_440,In_421,In_117);
nand U441 (N_441,In_403,In_296);
and U442 (N_442,In_175,In_111);
xnor U443 (N_443,In_616,In_354);
or U444 (N_444,In_336,In_671);
nand U445 (N_445,In_561,In_727);
or U446 (N_446,In_522,In_747);
and U447 (N_447,In_296,In_568);
nand U448 (N_448,In_47,In_471);
xnor U449 (N_449,In_236,In_429);
nand U450 (N_450,In_556,In_183);
nor U451 (N_451,In_163,In_50);
and U452 (N_452,In_146,In_84);
xnor U453 (N_453,In_490,In_485);
xor U454 (N_454,In_503,In_681);
and U455 (N_455,In_235,In_516);
xnor U456 (N_456,In_698,In_593);
nor U457 (N_457,In_253,In_24);
nand U458 (N_458,In_627,In_260);
and U459 (N_459,In_113,In_468);
nand U460 (N_460,In_111,In_118);
nor U461 (N_461,In_238,In_42);
nor U462 (N_462,In_334,In_729);
or U463 (N_463,In_73,In_686);
and U464 (N_464,In_661,In_50);
xor U465 (N_465,In_636,In_148);
nand U466 (N_466,In_288,In_245);
nor U467 (N_467,In_499,In_594);
xnor U468 (N_468,In_218,In_182);
nor U469 (N_469,In_77,In_633);
xnor U470 (N_470,In_697,In_743);
nor U471 (N_471,In_20,In_27);
xor U472 (N_472,In_33,In_167);
nand U473 (N_473,In_641,In_316);
nor U474 (N_474,In_749,In_413);
nand U475 (N_475,In_732,In_23);
nand U476 (N_476,In_632,In_323);
nor U477 (N_477,In_435,In_282);
nor U478 (N_478,In_219,In_430);
nand U479 (N_479,In_361,In_569);
nor U480 (N_480,In_389,In_220);
and U481 (N_481,In_169,In_480);
xnor U482 (N_482,In_350,In_435);
or U483 (N_483,In_688,In_623);
or U484 (N_484,In_321,In_436);
xor U485 (N_485,In_274,In_548);
nor U486 (N_486,In_511,In_346);
or U487 (N_487,In_581,In_303);
or U488 (N_488,In_216,In_102);
xor U489 (N_489,In_48,In_443);
nand U490 (N_490,In_314,In_165);
nand U491 (N_491,In_478,In_399);
nand U492 (N_492,In_186,In_6);
and U493 (N_493,In_339,In_467);
nor U494 (N_494,In_211,In_363);
xor U495 (N_495,In_397,In_267);
and U496 (N_496,In_482,In_8);
nand U497 (N_497,In_536,In_207);
nor U498 (N_498,In_359,In_545);
nor U499 (N_499,In_220,In_652);
or U500 (N_500,In_698,In_236);
xor U501 (N_501,In_487,In_194);
nand U502 (N_502,In_468,In_9);
and U503 (N_503,In_134,In_739);
xor U504 (N_504,In_401,In_159);
nor U505 (N_505,In_545,In_396);
or U506 (N_506,In_265,In_173);
nand U507 (N_507,In_194,In_421);
nand U508 (N_508,In_51,In_266);
or U509 (N_509,In_650,In_408);
xnor U510 (N_510,In_139,In_28);
and U511 (N_511,In_166,In_639);
and U512 (N_512,In_292,In_344);
nor U513 (N_513,In_631,In_695);
nand U514 (N_514,In_725,In_651);
and U515 (N_515,In_703,In_191);
or U516 (N_516,In_120,In_369);
nand U517 (N_517,In_164,In_105);
nand U518 (N_518,In_445,In_143);
xor U519 (N_519,In_682,In_239);
nor U520 (N_520,In_486,In_22);
xnor U521 (N_521,In_255,In_644);
nor U522 (N_522,In_632,In_262);
xor U523 (N_523,In_310,In_205);
and U524 (N_524,In_391,In_142);
or U525 (N_525,In_70,In_134);
nor U526 (N_526,In_135,In_144);
or U527 (N_527,In_461,In_197);
xnor U528 (N_528,In_561,In_652);
or U529 (N_529,In_634,In_428);
nand U530 (N_530,In_261,In_431);
xnor U531 (N_531,In_151,In_300);
nand U532 (N_532,In_373,In_184);
and U533 (N_533,In_285,In_227);
and U534 (N_534,In_362,In_479);
nand U535 (N_535,In_536,In_444);
or U536 (N_536,In_166,In_129);
nand U537 (N_537,In_469,In_636);
nor U538 (N_538,In_140,In_172);
or U539 (N_539,In_489,In_110);
xor U540 (N_540,In_258,In_280);
nor U541 (N_541,In_360,In_182);
nor U542 (N_542,In_674,In_203);
nand U543 (N_543,In_477,In_632);
nor U544 (N_544,In_463,In_230);
or U545 (N_545,In_217,In_659);
or U546 (N_546,In_0,In_638);
xnor U547 (N_547,In_564,In_709);
xnor U548 (N_548,In_656,In_496);
nor U549 (N_549,In_228,In_524);
or U550 (N_550,In_373,In_421);
nor U551 (N_551,In_719,In_54);
and U552 (N_552,In_306,In_388);
and U553 (N_553,In_3,In_728);
nor U554 (N_554,In_475,In_284);
and U555 (N_555,In_478,In_404);
or U556 (N_556,In_637,In_388);
or U557 (N_557,In_423,In_692);
nand U558 (N_558,In_77,In_284);
nor U559 (N_559,In_403,In_116);
nand U560 (N_560,In_1,In_619);
or U561 (N_561,In_694,In_170);
or U562 (N_562,In_632,In_235);
and U563 (N_563,In_263,In_613);
nand U564 (N_564,In_645,In_600);
nand U565 (N_565,In_485,In_311);
and U566 (N_566,In_40,In_237);
xnor U567 (N_567,In_489,In_681);
nor U568 (N_568,In_356,In_509);
nand U569 (N_569,In_710,In_602);
nor U570 (N_570,In_725,In_460);
or U571 (N_571,In_713,In_202);
xnor U572 (N_572,In_608,In_133);
nand U573 (N_573,In_163,In_78);
or U574 (N_574,In_208,In_72);
and U575 (N_575,In_40,In_48);
or U576 (N_576,In_558,In_258);
xnor U577 (N_577,In_658,In_288);
nor U578 (N_578,In_335,In_25);
nand U579 (N_579,In_408,In_81);
and U580 (N_580,In_206,In_253);
nor U581 (N_581,In_579,In_298);
and U582 (N_582,In_502,In_519);
nor U583 (N_583,In_123,In_214);
or U584 (N_584,In_112,In_368);
and U585 (N_585,In_97,In_655);
or U586 (N_586,In_312,In_193);
nand U587 (N_587,In_317,In_223);
xor U588 (N_588,In_249,In_501);
xnor U589 (N_589,In_380,In_361);
nand U590 (N_590,In_561,In_317);
nand U591 (N_591,In_454,In_75);
or U592 (N_592,In_122,In_169);
xnor U593 (N_593,In_354,In_396);
nor U594 (N_594,In_21,In_166);
nor U595 (N_595,In_409,In_168);
or U596 (N_596,In_589,In_93);
or U597 (N_597,In_174,In_215);
nand U598 (N_598,In_643,In_274);
nor U599 (N_599,In_262,In_53);
nor U600 (N_600,In_547,In_721);
and U601 (N_601,In_412,In_365);
nor U602 (N_602,In_701,In_529);
nor U603 (N_603,In_641,In_538);
xor U604 (N_604,In_2,In_655);
and U605 (N_605,In_18,In_702);
nor U606 (N_606,In_254,In_385);
or U607 (N_607,In_656,In_415);
and U608 (N_608,In_247,In_460);
or U609 (N_609,In_431,In_622);
and U610 (N_610,In_172,In_700);
nand U611 (N_611,In_76,In_467);
or U612 (N_612,In_594,In_361);
and U613 (N_613,In_454,In_284);
nor U614 (N_614,In_124,In_167);
and U615 (N_615,In_488,In_569);
nor U616 (N_616,In_565,In_614);
and U617 (N_617,In_362,In_466);
nand U618 (N_618,In_726,In_213);
nand U619 (N_619,In_76,In_390);
nand U620 (N_620,In_222,In_558);
xor U621 (N_621,In_0,In_361);
and U622 (N_622,In_111,In_440);
xnor U623 (N_623,In_706,In_394);
and U624 (N_624,In_291,In_492);
and U625 (N_625,In_664,In_550);
nor U626 (N_626,In_140,In_377);
and U627 (N_627,In_164,In_631);
and U628 (N_628,In_706,In_730);
or U629 (N_629,In_372,In_404);
nand U630 (N_630,In_352,In_652);
xnor U631 (N_631,In_743,In_646);
nor U632 (N_632,In_125,In_127);
nor U633 (N_633,In_528,In_556);
xnor U634 (N_634,In_507,In_301);
xnor U635 (N_635,In_439,In_175);
and U636 (N_636,In_471,In_247);
xnor U637 (N_637,In_394,In_608);
or U638 (N_638,In_740,In_205);
nand U639 (N_639,In_237,In_737);
xor U640 (N_640,In_492,In_499);
or U641 (N_641,In_605,In_353);
xnor U642 (N_642,In_172,In_563);
nor U643 (N_643,In_544,In_257);
and U644 (N_644,In_488,In_652);
nor U645 (N_645,In_323,In_263);
nor U646 (N_646,In_222,In_90);
and U647 (N_647,In_23,In_140);
or U648 (N_648,In_737,In_595);
nor U649 (N_649,In_111,In_115);
or U650 (N_650,In_101,In_432);
xnor U651 (N_651,In_732,In_434);
xnor U652 (N_652,In_369,In_525);
or U653 (N_653,In_534,In_556);
and U654 (N_654,In_313,In_28);
nand U655 (N_655,In_586,In_407);
or U656 (N_656,In_369,In_58);
nor U657 (N_657,In_638,In_181);
and U658 (N_658,In_580,In_202);
xnor U659 (N_659,In_22,In_623);
xnor U660 (N_660,In_280,In_261);
nand U661 (N_661,In_230,In_73);
and U662 (N_662,In_3,In_714);
or U663 (N_663,In_121,In_260);
nand U664 (N_664,In_581,In_69);
or U665 (N_665,In_461,In_739);
nor U666 (N_666,In_108,In_277);
nor U667 (N_667,In_354,In_517);
nor U668 (N_668,In_230,In_7);
or U669 (N_669,In_484,In_178);
nand U670 (N_670,In_520,In_115);
nor U671 (N_671,In_274,In_25);
xnor U672 (N_672,In_743,In_621);
or U673 (N_673,In_181,In_451);
nor U674 (N_674,In_418,In_475);
nor U675 (N_675,In_700,In_640);
nor U676 (N_676,In_582,In_27);
and U677 (N_677,In_488,In_381);
and U678 (N_678,In_687,In_66);
or U679 (N_679,In_431,In_442);
and U680 (N_680,In_38,In_544);
or U681 (N_681,In_639,In_449);
xor U682 (N_682,In_266,In_440);
nor U683 (N_683,In_742,In_520);
nand U684 (N_684,In_213,In_162);
nand U685 (N_685,In_504,In_140);
or U686 (N_686,In_153,In_450);
xnor U687 (N_687,In_579,In_546);
nand U688 (N_688,In_460,In_374);
or U689 (N_689,In_220,In_423);
xnor U690 (N_690,In_118,In_140);
nand U691 (N_691,In_474,In_362);
and U692 (N_692,In_451,In_605);
and U693 (N_693,In_730,In_641);
nor U694 (N_694,In_121,In_487);
xor U695 (N_695,In_100,In_132);
xnor U696 (N_696,In_325,In_658);
xnor U697 (N_697,In_24,In_296);
and U698 (N_698,In_708,In_280);
xnor U699 (N_699,In_178,In_503);
nand U700 (N_700,In_614,In_407);
nand U701 (N_701,In_486,In_2);
and U702 (N_702,In_133,In_227);
and U703 (N_703,In_128,In_733);
nand U704 (N_704,In_615,In_84);
nand U705 (N_705,In_620,In_208);
and U706 (N_706,In_727,In_370);
nor U707 (N_707,In_274,In_662);
xor U708 (N_708,In_262,In_333);
nand U709 (N_709,In_360,In_667);
or U710 (N_710,In_511,In_26);
xor U711 (N_711,In_683,In_605);
nor U712 (N_712,In_718,In_249);
and U713 (N_713,In_17,In_342);
and U714 (N_714,In_242,In_564);
nand U715 (N_715,In_569,In_574);
xnor U716 (N_716,In_394,In_619);
xnor U717 (N_717,In_202,In_611);
or U718 (N_718,In_517,In_667);
nor U719 (N_719,In_427,In_27);
nand U720 (N_720,In_187,In_510);
xnor U721 (N_721,In_222,In_546);
nand U722 (N_722,In_552,In_642);
or U723 (N_723,In_715,In_147);
or U724 (N_724,In_398,In_163);
or U725 (N_725,In_215,In_463);
nand U726 (N_726,In_122,In_518);
and U727 (N_727,In_342,In_217);
or U728 (N_728,In_390,In_138);
and U729 (N_729,In_572,In_13);
nor U730 (N_730,In_136,In_650);
xnor U731 (N_731,In_736,In_500);
xnor U732 (N_732,In_663,In_137);
or U733 (N_733,In_583,In_182);
nand U734 (N_734,In_407,In_218);
nor U735 (N_735,In_97,In_346);
and U736 (N_736,In_31,In_453);
or U737 (N_737,In_446,In_33);
nor U738 (N_738,In_612,In_29);
nand U739 (N_739,In_333,In_717);
nor U740 (N_740,In_344,In_477);
nand U741 (N_741,In_117,In_484);
nand U742 (N_742,In_138,In_610);
or U743 (N_743,In_69,In_582);
and U744 (N_744,In_706,In_16);
and U745 (N_745,In_394,In_632);
and U746 (N_746,In_545,In_745);
or U747 (N_747,In_703,In_269);
and U748 (N_748,In_334,In_717);
nand U749 (N_749,In_481,In_234);
and U750 (N_750,In_396,In_331);
nand U751 (N_751,In_155,In_91);
xor U752 (N_752,In_150,In_572);
xor U753 (N_753,In_457,In_358);
and U754 (N_754,In_334,In_133);
nand U755 (N_755,In_186,In_131);
xnor U756 (N_756,In_288,In_438);
nor U757 (N_757,In_467,In_704);
and U758 (N_758,In_248,In_278);
nand U759 (N_759,In_457,In_257);
xor U760 (N_760,In_330,In_421);
and U761 (N_761,In_375,In_475);
nor U762 (N_762,In_247,In_41);
and U763 (N_763,In_369,In_206);
and U764 (N_764,In_402,In_334);
and U765 (N_765,In_54,In_228);
nor U766 (N_766,In_250,In_495);
xnor U767 (N_767,In_724,In_35);
and U768 (N_768,In_469,In_197);
nand U769 (N_769,In_431,In_10);
and U770 (N_770,In_160,In_669);
nor U771 (N_771,In_245,In_548);
nor U772 (N_772,In_708,In_40);
or U773 (N_773,In_715,In_67);
xnor U774 (N_774,In_49,In_511);
and U775 (N_775,In_429,In_507);
nand U776 (N_776,In_71,In_369);
or U777 (N_777,In_579,In_573);
nand U778 (N_778,In_729,In_503);
xnor U779 (N_779,In_709,In_662);
nand U780 (N_780,In_550,In_419);
nand U781 (N_781,In_195,In_74);
or U782 (N_782,In_239,In_191);
or U783 (N_783,In_743,In_512);
xor U784 (N_784,In_724,In_215);
nand U785 (N_785,In_458,In_351);
and U786 (N_786,In_600,In_436);
xnor U787 (N_787,In_399,In_248);
nand U788 (N_788,In_33,In_674);
xnor U789 (N_789,In_38,In_719);
nor U790 (N_790,In_736,In_558);
nor U791 (N_791,In_656,In_404);
nor U792 (N_792,In_122,In_553);
xor U793 (N_793,In_272,In_164);
xnor U794 (N_794,In_210,In_327);
or U795 (N_795,In_28,In_446);
nand U796 (N_796,In_452,In_616);
nand U797 (N_797,In_606,In_388);
xnor U798 (N_798,In_239,In_444);
and U799 (N_799,In_169,In_485);
xor U800 (N_800,In_360,In_226);
xnor U801 (N_801,In_448,In_1);
xor U802 (N_802,In_257,In_105);
xnor U803 (N_803,In_517,In_572);
or U804 (N_804,In_595,In_83);
nor U805 (N_805,In_267,In_621);
nor U806 (N_806,In_285,In_338);
xnor U807 (N_807,In_475,In_297);
nand U808 (N_808,In_168,In_633);
xor U809 (N_809,In_114,In_662);
or U810 (N_810,In_205,In_26);
xnor U811 (N_811,In_119,In_332);
nand U812 (N_812,In_466,In_391);
nand U813 (N_813,In_397,In_537);
xnor U814 (N_814,In_56,In_562);
and U815 (N_815,In_466,In_577);
nand U816 (N_816,In_255,In_635);
or U817 (N_817,In_570,In_679);
and U818 (N_818,In_580,In_699);
xnor U819 (N_819,In_327,In_208);
nor U820 (N_820,In_499,In_724);
and U821 (N_821,In_194,In_448);
and U822 (N_822,In_666,In_317);
xor U823 (N_823,In_344,In_25);
or U824 (N_824,In_3,In_458);
nand U825 (N_825,In_477,In_517);
xnor U826 (N_826,In_63,In_116);
or U827 (N_827,In_22,In_663);
xnor U828 (N_828,In_454,In_648);
or U829 (N_829,In_136,In_443);
or U830 (N_830,In_633,In_746);
nor U831 (N_831,In_735,In_498);
and U832 (N_832,In_594,In_53);
xor U833 (N_833,In_628,In_745);
nor U834 (N_834,In_411,In_307);
or U835 (N_835,In_217,In_257);
nand U836 (N_836,In_294,In_268);
and U837 (N_837,In_485,In_585);
and U838 (N_838,In_430,In_3);
or U839 (N_839,In_660,In_615);
or U840 (N_840,In_272,In_712);
and U841 (N_841,In_746,In_35);
and U842 (N_842,In_349,In_649);
nand U843 (N_843,In_394,In_276);
nand U844 (N_844,In_273,In_711);
nand U845 (N_845,In_567,In_493);
and U846 (N_846,In_98,In_577);
xnor U847 (N_847,In_499,In_368);
and U848 (N_848,In_39,In_337);
xor U849 (N_849,In_59,In_457);
xnor U850 (N_850,In_73,In_688);
nor U851 (N_851,In_187,In_56);
and U852 (N_852,In_156,In_540);
xnor U853 (N_853,In_273,In_485);
or U854 (N_854,In_473,In_288);
and U855 (N_855,In_605,In_619);
xor U856 (N_856,In_217,In_412);
xnor U857 (N_857,In_15,In_59);
nor U858 (N_858,In_478,In_181);
and U859 (N_859,In_478,In_711);
nand U860 (N_860,In_319,In_119);
nand U861 (N_861,In_291,In_671);
nor U862 (N_862,In_146,In_177);
nor U863 (N_863,In_702,In_440);
nand U864 (N_864,In_699,In_95);
nand U865 (N_865,In_349,In_402);
nor U866 (N_866,In_441,In_677);
or U867 (N_867,In_692,In_685);
nand U868 (N_868,In_63,In_391);
or U869 (N_869,In_553,In_609);
xor U870 (N_870,In_101,In_513);
nor U871 (N_871,In_561,In_232);
nor U872 (N_872,In_141,In_80);
xor U873 (N_873,In_167,In_326);
and U874 (N_874,In_8,In_334);
nor U875 (N_875,In_359,In_99);
and U876 (N_876,In_226,In_216);
nor U877 (N_877,In_68,In_345);
nor U878 (N_878,In_195,In_9);
or U879 (N_879,In_357,In_199);
xnor U880 (N_880,In_238,In_643);
nor U881 (N_881,In_587,In_592);
and U882 (N_882,In_73,In_387);
and U883 (N_883,In_16,In_185);
xor U884 (N_884,In_456,In_203);
nor U885 (N_885,In_697,In_479);
or U886 (N_886,In_504,In_701);
xnor U887 (N_887,In_591,In_120);
xor U888 (N_888,In_439,In_248);
nor U889 (N_889,In_79,In_173);
nand U890 (N_890,In_490,In_114);
or U891 (N_891,In_439,In_120);
xnor U892 (N_892,In_101,In_206);
nor U893 (N_893,In_355,In_232);
nand U894 (N_894,In_49,In_110);
and U895 (N_895,In_540,In_109);
or U896 (N_896,In_704,In_391);
nor U897 (N_897,In_352,In_369);
and U898 (N_898,In_180,In_94);
nor U899 (N_899,In_213,In_178);
xor U900 (N_900,In_215,In_189);
nor U901 (N_901,In_392,In_16);
xor U902 (N_902,In_340,In_408);
nor U903 (N_903,In_659,In_328);
and U904 (N_904,In_134,In_742);
or U905 (N_905,In_681,In_688);
xnor U906 (N_906,In_481,In_326);
or U907 (N_907,In_201,In_647);
xnor U908 (N_908,In_291,In_591);
xor U909 (N_909,In_746,In_301);
nand U910 (N_910,In_309,In_540);
nor U911 (N_911,In_327,In_676);
nor U912 (N_912,In_611,In_664);
xor U913 (N_913,In_512,In_181);
nor U914 (N_914,In_725,In_653);
and U915 (N_915,In_94,In_667);
nand U916 (N_916,In_379,In_54);
nand U917 (N_917,In_429,In_679);
nand U918 (N_918,In_392,In_620);
nor U919 (N_919,In_555,In_305);
nor U920 (N_920,In_554,In_26);
xnor U921 (N_921,In_553,In_361);
nand U922 (N_922,In_511,In_696);
nand U923 (N_923,In_259,In_222);
or U924 (N_924,In_273,In_44);
and U925 (N_925,In_684,In_673);
nand U926 (N_926,In_148,In_63);
xor U927 (N_927,In_391,In_314);
or U928 (N_928,In_277,In_556);
nor U929 (N_929,In_73,In_367);
or U930 (N_930,In_666,In_648);
nor U931 (N_931,In_273,In_264);
or U932 (N_932,In_110,In_19);
xor U933 (N_933,In_727,In_155);
nor U934 (N_934,In_426,In_302);
nor U935 (N_935,In_630,In_567);
xor U936 (N_936,In_490,In_55);
or U937 (N_937,In_523,In_240);
nand U938 (N_938,In_739,In_174);
and U939 (N_939,In_457,In_695);
or U940 (N_940,In_718,In_553);
nor U941 (N_941,In_662,In_74);
and U942 (N_942,In_517,In_299);
and U943 (N_943,In_672,In_81);
and U944 (N_944,In_429,In_522);
and U945 (N_945,In_222,In_4);
nand U946 (N_946,In_242,In_317);
or U947 (N_947,In_508,In_488);
and U948 (N_948,In_544,In_168);
or U949 (N_949,In_642,In_316);
or U950 (N_950,In_386,In_114);
and U951 (N_951,In_462,In_743);
xor U952 (N_952,In_467,In_432);
xnor U953 (N_953,In_329,In_89);
nand U954 (N_954,In_138,In_499);
or U955 (N_955,In_637,In_358);
or U956 (N_956,In_186,In_250);
nor U957 (N_957,In_436,In_196);
nand U958 (N_958,In_18,In_215);
or U959 (N_959,In_340,In_642);
xor U960 (N_960,In_603,In_667);
and U961 (N_961,In_469,In_450);
xnor U962 (N_962,In_352,In_425);
and U963 (N_963,In_711,In_148);
xor U964 (N_964,In_331,In_346);
nand U965 (N_965,In_223,In_439);
xnor U966 (N_966,In_162,In_148);
nand U967 (N_967,In_49,In_630);
and U968 (N_968,In_514,In_175);
nor U969 (N_969,In_444,In_582);
xnor U970 (N_970,In_744,In_407);
and U971 (N_971,In_495,In_371);
xnor U972 (N_972,In_260,In_601);
xnor U973 (N_973,In_213,In_537);
xor U974 (N_974,In_328,In_593);
nor U975 (N_975,In_423,In_401);
and U976 (N_976,In_573,In_430);
nor U977 (N_977,In_111,In_394);
nor U978 (N_978,In_295,In_396);
nor U979 (N_979,In_666,In_160);
xor U980 (N_980,In_257,In_621);
or U981 (N_981,In_84,In_23);
nor U982 (N_982,In_250,In_54);
or U983 (N_983,In_164,In_72);
or U984 (N_984,In_50,In_124);
and U985 (N_985,In_196,In_240);
nor U986 (N_986,In_544,In_371);
or U987 (N_987,In_570,In_478);
or U988 (N_988,In_295,In_461);
and U989 (N_989,In_674,In_745);
xnor U990 (N_990,In_11,In_3);
or U991 (N_991,In_353,In_230);
and U992 (N_992,In_542,In_501);
nand U993 (N_993,In_591,In_154);
or U994 (N_994,In_650,In_127);
nor U995 (N_995,In_159,In_35);
and U996 (N_996,In_42,In_311);
or U997 (N_997,In_364,In_743);
xor U998 (N_998,In_523,In_267);
xor U999 (N_999,In_226,In_395);
or U1000 (N_1000,In_736,In_303);
and U1001 (N_1001,In_286,In_34);
xor U1002 (N_1002,In_221,In_227);
nand U1003 (N_1003,In_521,In_329);
xnor U1004 (N_1004,In_509,In_714);
nor U1005 (N_1005,In_33,In_213);
and U1006 (N_1006,In_400,In_592);
nand U1007 (N_1007,In_181,In_423);
and U1008 (N_1008,In_392,In_740);
xor U1009 (N_1009,In_134,In_117);
or U1010 (N_1010,In_273,In_667);
or U1011 (N_1011,In_724,In_734);
and U1012 (N_1012,In_404,In_108);
xor U1013 (N_1013,In_538,In_257);
nor U1014 (N_1014,In_120,In_438);
and U1015 (N_1015,In_297,In_129);
nand U1016 (N_1016,In_588,In_4);
and U1017 (N_1017,In_415,In_193);
nor U1018 (N_1018,In_543,In_0);
nand U1019 (N_1019,In_732,In_584);
nand U1020 (N_1020,In_289,In_536);
or U1021 (N_1021,In_525,In_284);
or U1022 (N_1022,In_117,In_601);
nand U1023 (N_1023,In_434,In_711);
nor U1024 (N_1024,In_292,In_200);
nand U1025 (N_1025,In_197,In_185);
or U1026 (N_1026,In_207,In_489);
nor U1027 (N_1027,In_27,In_596);
nor U1028 (N_1028,In_607,In_7);
or U1029 (N_1029,In_532,In_94);
xor U1030 (N_1030,In_47,In_453);
nor U1031 (N_1031,In_308,In_682);
nor U1032 (N_1032,In_49,In_705);
nor U1033 (N_1033,In_204,In_458);
nand U1034 (N_1034,In_105,In_434);
xor U1035 (N_1035,In_613,In_582);
nor U1036 (N_1036,In_746,In_474);
nand U1037 (N_1037,In_615,In_42);
nor U1038 (N_1038,In_446,In_440);
nor U1039 (N_1039,In_607,In_590);
or U1040 (N_1040,In_70,In_325);
nor U1041 (N_1041,In_389,In_27);
xnor U1042 (N_1042,In_744,In_160);
or U1043 (N_1043,In_409,In_744);
nand U1044 (N_1044,In_429,In_31);
xor U1045 (N_1045,In_103,In_747);
xor U1046 (N_1046,In_673,In_131);
nand U1047 (N_1047,In_287,In_575);
nand U1048 (N_1048,In_140,In_619);
or U1049 (N_1049,In_458,In_410);
nor U1050 (N_1050,In_252,In_722);
or U1051 (N_1051,In_49,In_374);
nor U1052 (N_1052,In_587,In_523);
or U1053 (N_1053,In_519,In_229);
xor U1054 (N_1054,In_241,In_694);
nor U1055 (N_1055,In_396,In_713);
nor U1056 (N_1056,In_480,In_641);
nand U1057 (N_1057,In_591,In_644);
and U1058 (N_1058,In_130,In_107);
and U1059 (N_1059,In_574,In_232);
nand U1060 (N_1060,In_589,In_66);
nand U1061 (N_1061,In_745,In_181);
nor U1062 (N_1062,In_288,In_521);
xnor U1063 (N_1063,In_453,In_76);
nor U1064 (N_1064,In_482,In_40);
and U1065 (N_1065,In_693,In_699);
nor U1066 (N_1066,In_707,In_70);
or U1067 (N_1067,In_627,In_603);
or U1068 (N_1068,In_735,In_539);
or U1069 (N_1069,In_738,In_474);
or U1070 (N_1070,In_571,In_548);
nor U1071 (N_1071,In_571,In_703);
or U1072 (N_1072,In_358,In_207);
xnor U1073 (N_1073,In_8,In_691);
nand U1074 (N_1074,In_41,In_531);
nor U1075 (N_1075,In_665,In_477);
xor U1076 (N_1076,In_499,In_207);
and U1077 (N_1077,In_148,In_224);
nand U1078 (N_1078,In_341,In_274);
and U1079 (N_1079,In_381,In_210);
nand U1080 (N_1080,In_486,In_74);
or U1081 (N_1081,In_524,In_187);
and U1082 (N_1082,In_289,In_730);
or U1083 (N_1083,In_246,In_662);
or U1084 (N_1084,In_268,In_235);
xnor U1085 (N_1085,In_466,In_236);
and U1086 (N_1086,In_532,In_531);
nor U1087 (N_1087,In_347,In_540);
or U1088 (N_1088,In_489,In_42);
or U1089 (N_1089,In_317,In_84);
nand U1090 (N_1090,In_80,In_306);
nor U1091 (N_1091,In_694,In_630);
and U1092 (N_1092,In_477,In_96);
or U1093 (N_1093,In_491,In_354);
or U1094 (N_1094,In_397,In_279);
xnor U1095 (N_1095,In_705,In_48);
and U1096 (N_1096,In_156,In_136);
xor U1097 (N_1097,In_585,In_110);
nand U1098 (N_1098,In_135,In_699);
or U1099 (N_1099,In_148,In_413);
xnor U1100 (N_1100,In_380,In_201);
nand U1101 (N_1101,In_151,In_585);
nor U1102 (N_1102,In_647,In_178);
nor U1103 (N_1103,In_346,In_739);
nand U1104 (N_1104,In_725,In_38);
and U1105 (N_1105,In_697,In_52);
xor U1106 (N_1106,In_578,In_198);
xnor U1107 (N_1107,In_507,In_393);
or U1108 (N_1108,In_578,In_328);
and U1109 (N_1109,In_627,In_593);
nand U1110 (N_1110,In_440,In_448);
and U1111 (N_1111,In_304,In_101);
xnor U1112 (N_1112,In_142,In_687);
or U1113 (N_1113,In_148,In_27);
or U1114 (N_1114,In_42,In_290);
xnor U1115 (N_1115,In_284,In_656);
or U1116 (N_1116,In_247,In_396);
and U1117 (N_1117,In_57,In_454);
or U1118 (N_1118,In_61,In_448);
and U1119 (N_1119,In_320,In_111);
nor U1120 (N_1120,In_534,In_37);
nor U1121 (N_1121,In_669,In_333);
nor U1122 (N_1122,In_620,In_700);
and U1123 (N_1123,In_303,In_160);
nand U1124 (N_1124,In_294,In_617);
and U1125 (N_1125,In_193,In_91);
nor U1126 (N_1126,In_727,In_197);
xor U1127 (N_1127,In_10,In_22);
xnor U1128 (N_1128,In_118,In_666);
xnor U1129 (N_1129,In_415,In_10);
and U1130 (N_1130,In_67,In_714);
nand U1131 (N_1131,In_197,In_497);
nor U1132 (N_1132,In_621,In_62);
xnor U1133 (N_1133,In_501,In_612);
xor U1134 (N_1134,In_705,In_233);
nand U1135 (N_1135,In_534,In_742);
nand U1136 (N_1136,In_365,In_604);
nor U1137 (N_1137,In_457,In_313);
nand U1138 (N_1138,In_495,In_608);
xnor U1139 (N_1139,In_677,In_29);
nor U1140 (N_1140,In_263,In_650);
and U1141 (N_1141,In_437,In_603);
nand U1142 (N_1142,In_46,In_649);
nand U1143 (N_1143,In_493,In_53);
and U1144 (N_1144,In_498,In_481);
nor U1145 (N_1145,In_564,In_174);
or U1146 (N_1146,In_69,In_652);
nor U1147 (N_1147,In_367,In_438);
or U1148 (N_1148,In_516,In_420);
xor U1149 (N_1149,In_465,In_630);
and U1150 (N_1150,In_99,In_48);
and U1151 (N_1151,In_615,In_567);
nor U1152 (N_1152,In_511,In_467);
and U1153 (N_1153,In_167,In_408);
nand U1154 (N_1154,In_484,In_309);
nor U1155 (N_1155,In_139,In_89);
or U1156 (N_1156,In_28,In_234);
nor U1157 (N_1157,In_552,In_317);
and U1158 (N_1158,In_580,In_247);
xnor U1159 (N_1159,In_718,In_356);
and U1160 (N_1160,In_163,In_339);
and U1161 (N_1161,In_110,In_233);
nand U1162 (N_1162,In_590,In_422);
nand U1163 (N_1163,In_153,In_552);
nor U1164 (N_1164,In_507,In_560);
and U1165 (N_1165,In_246,In_274);
and U1166 (N_1166,In_64,In_658);
xnor U1167 (N_1167,In_664,In_426);
nand U1168 (N_1168,In_721,In_87);
nor U1169 (N_1169,In_186,In_312);
nand U1170 (N_1170,In_74,In_393);
or U1171 (N_1171,In_721,In_579);
nand U1172 (N_1172,In_214,In_81);
nor U1173 (N_1173,In_570,In_536);
nor U1174 (N_1174,In_392,In_102);
nand U1175 (N_1175,In_175,In_311);
and U1176 (N_1176,In_13,In_607);
or U1177 (N_1177,In_342,In_216);
nand U1178 (N_1178,In_431,In_246);
and U1179 (N_1179,In_714,In_233);
or U1180 (N_1180,In_255,In_49);
nor U1181 (N_1181,In_147,In_431);
xor U1182 (N_1182,In_132,In_401);
and U1183 (N_1183,In_523,In_691);
nand U1184 (N_1184,In_686,In_510);
and U1185 (N_1185,In_133,In_179);
nor U1186 (N_1186,In_266,In_132);
or U1187 (N_1187,In_307,In_201);
nor U1188 (N_1188,In_375,In_425);
nand U1189 (N_1189,In_563,In_730);
or U1190 (N_1190,In_636,In_80);
nand U1191 (N_1191,In_586,In_625);
xor U1192 (N_1192,In_391,In_100);
or U1193 (N_1193,In_98,In_295);
or U1194 (N_1194,In_439,In_133);
nand U1195 (N_1195,In_8,In_463);
nor U1196 (N_1196,In_374,In_660);
nand U1197 (N_1197,In_374,In_509);
xor U1198 (N_1198,In_193,In_614);
or U1199 (N_1199,In_655,In_609);
nand U1200 (N_1200,In_587,In_374);
xnor U1201 (N_1201,In_720,In_293);
nor U1202 (N_1202,In_33,In_692);
and U1203 (N_1203,In_260,In_245);
nand U1204 (N_1204,In_724,In_296);
xnor U1205 (N_1205,In_97,In_569);
xor U1206 (N_1206,In_87,In_207);
or U1207 (N_1207,In_619,In_112);
nor U1208 (N_1208,In_701,In_340);
and U1209 (N_1209,In_630,In_725);
and U1210 (N_1210,In_441,In_229);
xor U1211 (N_1211,In_489,In_83);
and U1212 (N_1212,In_359,In_644);
and U1213 (N_1213,In_118,In_37);
nor U1214 (N_1214,In_80,In_711);
nor U1215 (N_1215,In_362,In_520);
or U1216 (N_1216,In_267,In_599);
and U1217 (N_1217,In_585,In_375);
nor U1218 (N_1218,In_180,In_41);
xor U1219 (N_1219,In_521,In_43);
or U1220 (N_1220,In_722,In_417);
xor U1221 (N_1221,In_204,In_309);
or U1222 (N_1222,In_479,In_707);
nor U1223 (N_1223,In_746,In_535);
nor U1224 (N_1224,In_444,In_2);
and U1225 (N_1225,In_411,In_73);
nand U1226 (N_1226,In_524,In_350);
or U1227 (N_1227,In_289,In_73);
nand U1228 (N_1228,In_234,In_534);
nor U1229 (N_1229,In_432,In_593);
nor U1230 (N_1230,In_488,In_225);
or U1231 (N_1231,In_474,In_223);
xor U1232 (N_1232,In_591,In_255);
and U1233 (N_1233,In_487,In_241);
and U1234 (N_1234,In_359,In_604);
xnor U1235 (N_1235,In_433,In_94);
nor U1236 (N_1236,In_437,In_92);
and U1237 (N_1237,In_722,In_98);
xor U1238 (N_1238,In_601,In_233);
nand U1239 (N_1239,In_402,In_88);
or U1240 (N_1240,In_664,In_84);
and U1241 (N_1241,In_519,In_593);
or U1242 (N_1242,In_630,In_472);
xnor U1243 (N_1243,In_387,In_357);
nor U1244 (N_1244,In_528,In_522);
nor U1245 (N_1245,In_60,In_313);
and U1246 (N_1246,In_630,In_166);
xor U1247 (N_1247,In_424,In_7);
nor U1248 (N_1248,In_219,In_12);
nand U1249 (N_1249,In_709,In_92);
nor U1250 (N_1250,In_33,In_386);
nand U1251 (N_1251,In_185,In_222);
nand U1252 (N_1252,In_401,In_704);
xnor U1253 (N_1253,In_193,In_258);
or U1254 (N_1254,In_193,In_539);
and U1255 (N_1255,In_745,In_22);
and U1256 (N_1256,In_10,In_737);
or U1257 (N_1257,In_541,In_662);
nor U1258 (N_1258,In_613,In_73);
xor U1259 (N_1259,In_401,In_686);
and U1260 (N_1260,In_100,In_304);
xnor U1261 (N_1261,In_574,In_659);
nor U1262 (N_1262,In_202,In_517);
and U1263 (N_1263,In_589,In_345);
and U1264 (N_1264,In_359,In_737);
nor U1265 (N_1265,In_41,In_205);
nand U1266 (N_1266,In_416,In_570);
and U1267 (N_1267,In_673,In_477);
nand U1268 (N_1268,In_330,In_572);
xnor U1269 (N_1269,In_80,In_538);
nand U1270 (N_1270,In_51,In_716);
and U1271 (N_1271,In_208,In_261);
nand U1272 (N_1272,In_680,In_319);
and U1273 (N_1273,In_336,In_461);
xnor U1274 (N_1274,In_278,In_413);
nand U1275 (N_1275,In_379,In_664);
or U1276 (N_1276,In_527,In_136);
nor U1277 (N_1277,In_88,In_468);
xor U1278 (N_1278,In_538,In_668);
nor U1279 (N_1279,In_74,In_337);
or U1280 (N_1280,In_532,In_442);
or U1281 (N_1281,In_219,In_726);
nand U1282 (N_1282,In_28,In_623);
and U1283 (N_1283,In_402,In_600);
xor U1284 (N_1284,In_627,In_577);
nand U1285 (N_1285,In_155,In_136);
nand U1286 (N_1286,In_343,In_130);
nor U1287 (N_1287,In_676,In_610);
xnor U1288 (N_1288,In_688,In_613);
nor U1289 (N_1289,In_103,In_473);
or U1290 (N_1290,In_91,In_243);
xor U1291 (N_1291,In_739,In_184);
or U1292 (N_1292,In_743,In_668);
nor U1293 (N_1293,In_340,In_347);
nor U1294 (N_1294,In_539,In_364);
xnor U1295 (N_1295,In_607,In_594);
and U1296 (N_1296,In_491,In_702);
and U1297 (N_1297,In_332,In_625);
and U1298 (N_1298,In_276,In_426);
nand U1299 (N_1299,In_336,In_323);
nor U1300 (N_1300,In_451,In_406);
xor U1301 (N_1301,In_415,In_99);
xor U1302 (N_1302,In_464,In_274);
and U1303 (N_1303,In_276,In_572);
or U1304 (N_1304,In_16,In_704);
nand U1305 (N_1305,In_427,In_255);
xnor U1306 (N_1306,In_438,In_736);
xnor U1307 (N_1307,In_35,In_458);
or U1308 (N_1308,In_284,In_628);
nand U1309 (N_1309,In_11,In_37);
xor U1310 (N_1310,In_525,In_48);
nand U1311 (N_1311,In_67,In_698);
or U1312 (N_1312,In_358,In_174);
nand U1313 (N_1313,In_440,In_707);
nand U1314 (N_1314,In_599,In_352);
xnor U1315 (N_1315,In_603,In_20);
nor U1316 (N_1316,In_492,In_565);
nand U1317 (N_1317,In_468,In_269);
nand U1318 (N_1318,In_387,In_478);
nor U1319 (N_1319,In_516,In_457);
or U1320 (N_1320,In_112,In_248);
xor U1321 (N_1321,In_645,In_625);
nor U1322 (N_1322,In_589,In_596);
nand U1323 (N_1323,In_314,In_184);
nor U1324 (N_1324,In_665,In_595);
and U1325 (N_1325,In_440,In_268);
xor U1326 (N_1326,In_624,In_430);
and U1327 (N_1327,In_308,In_3);
and U1328 (N_1328,In_588,In_154);
nand U1329 (N_1329,In_111,In_392);
or U1330 (N_1330,In_174,In_514);
xor U1331 (N_1331,In_445,In_682);
or U1332 (N_1332,In_662,In_686);
nor U1333 (N_1333,In_175,In_330);
or U1334 (N_1334,In_553,In_31);
xor U1335 (N_1335,In_699,In_2);
nor U1336 (N_1336,In_183,In_731);
or U1337 (N_1337,In_85,In_235);
or U1338 (N_1338,In_730,In_453);
or U1339 (N_1339,In_656,In_178);
nor U1340 (N_1340,In_119,In_38);
xnor U1341 (N_1341,In_467,In_0);
and U1342 (N_1342,In_592,In_658);
nor U1343 (N_1343,In_539,In_372);
nand U1344 (N_1344,In_107,In_498);
or U1345 (N_1345,In_21,In_630);
nor U1346 (N_1346,In_477,In_677);
nand U1347 (N_1347,In_53,In_742);
nor U1348 (N_1348,In_624,In_516);
xor U1349 (N_1349,In_506,In_72);
and U1350 (N_1350,In_700,In_419);
or U1351 (N_1351,In_215,In_664);
xnor U1352 (N_1352,In_222,In_469);
xnor U1353 (N_1353,In_145,In_154);
or U1354 (N_1354,In_446,In_498);
or U1355 (N_1355,In_229,In_13);
nand U1356 (N_1356,In_697,In_466);
or U1357 (N_1357,In_603,In_73);
or U1358 (N_1358,In_623,In_523);
or U1359 (N_1359,In_602,In_633);
nand U1360 (N_1360,In_328,In_747);
nor U1361 (N_1361,In_267,In_390);
or U1362 (N_1362,In_197,In_297);
nand U1363 (N_1363,In_533,In_462);
nand U1364 (N_1364,In_438,In_291);
xor U1365 (N_1365,In_184,In_253);
nand U1366 (N_1366,In_298,In_584);
nand U1367 (N_1367,In_594,In_59);
xor U1368 (N_1368,In_749,In_629);
nor U1369 (N_1369,In_697,In_638);
or U1370 (N_1370,In_8,In_662);
or U1371 (N_1371,In_413,In_424);
xnor U1372 (N_1372,In_260,In_243);
nand U1373 (N_1373,In_116,In_199);
or U1374 (N_1374,In_33,In_80);
nand U1375 (N_1375,In_74,In_234);
nor U1376 (N_1376,In_127,In_218);
and U1377 (N_1377,In_445,In_710);
nand U1378 (N_1378,In_32,In_113);
xor U1379 (N_1379,In_515,In_160);
or U1380 (N_1380,In_268,In_389);
or U1381 (N_1381,In_511,In_682);
and U1382 (N_1382,In_134,In_460);
or U1383 (N_1383,In_452,In_725);
and U1384 (N_1384,In_626,In_419);
or U1385 (N_1385,In_456,In_535);
or U1386 (N_1386,In_542,In_147);
nor U1387 (N_1387,In_284,In_511);
and U1388 (N_1388,In_514,In_253);
nor U1389 (N_1389,In_344,In_162);
xor U1390 (N_1390,In_108,In_554);
nor U1391 (N_1391,In_28,In_575);
xor U1392 (N_1392,In_154,In_463);
or U1393 (N_1393,In_524,In_216);
or U1394 (N_1394,In_363,In_74);
and U1395 (N_1395,In_150,In_472);
nor U1396 (N_1396,In_120,In_500);
nor U1397 (N_1397,In_651,In_515);
and U1398 (N_1398,In_728,In_725);
or U1399 (N_1399,In_201,In_293);
or U1400 (N_1400,In_426,In_748);
xor U1401 (N_1401,In_670,In_405);
or U1402 (N_1402,In_99,In_190);
or U1403 (N_1403,In_293,In_321);
or U1404 (N_1404,In_734,In_250);
or U1405 (N_1405,In_411,In_178);
xor U1406 (N_1406,In_349,In_385);
xnor U1407 (N_1407,In_724,In_223);
or U1408 (N_1408,In_591,In_563);
and U1409 (N_1409,In_520,In_655);
xor U1410 (N_1410,In_33,In_16);
xor U1411 (N_1411,In_542,In_432);
nor U1412 (N_1412,In_626,In_85);
nand U1413 (N_1413,In_721,In_558);
xnor U1414 (N_1414,In_136,In_530);
or U1415 (N_1415,In_513,In_392);
nand U1416 (N_1416,In_60,In_386);
nor U1417 (N_1417,In_685,In_105);
xnor U1418 (N_1418,In_659,In_565);
xor U1419 (N_1419,In_688,In_274);
xor U1420 (N_1420,In_459,In_604);
or U1421 (N_1421,In_641,In_308);
nor U1422 (N_1422,In_228,In_659);
nand U1423 (N_1423,In_210,In_137);
xnor U1424 (N_1424,In_446,In_735);
nor U1425 (N_1425,In_422,In_503);
xnor U1426 (N_1426,In_650,In_70);
and U1427 (N_1427,In_661,In_113);
and U1428 (N_1428,In_377,In_614);
or U1429 (N_1429,In_602,In_130);
nor U1430 (N_1430,In_546,In_532);
nand U1431 (N_1431,In_487,In_654);
and U1432 (N_1432,In_429,In_44);
xor U1433 (N_1433,In_683,In_247);
nor U1434 (N_1434,In_331,In_711);
nor U1435 (N_1435,In_182,In_345);
nor U1436 (N_1436,In_10,In_652);
nand U1437 (N_1437,In_138,In_482);
or U1438 (N_1438,In_432,In_664);
or U1439 (N_1439,In_607,In_314);
nand U1440 (N_1440,In_748,In_3);
and U1441 (N_1441,In_370,In_494);
nand U1442 (N_1442,In_196,In_676);
nand U1443 (N_1443,In_387,In_376);
or U1444 (N_1444,In_325,In_733);
nor U1445 (N_1445,In_432,In_226);
nor U1446 (N_1446,In_229,In_0);
xnor U1447 (N_1447,In_528,In_253);
nand U1448 (N_1448,In_556,In_251);
nand U1449 (N_1449,In_81,In_130);
nand U1450 (N_1450,In_477,In_425);
or U1451 (N_1451,In_299,In_668);
or U1452 (N_1452,In_646,In_37);
nor U1453 (N_1453,In_136,In_718);
and U1454 (N_1454,In_584,In_55);
xor U1455 (N_1455,In_615,In_512);
and U1456 (N_1456,In_247,In_65);
and U1457 (N_1457,In_170,In_280);
or U1458 (N_1458,In_549,In_17);
and U1459 (N_1459,In_742,In_126);
xnor U1460 (N_1460,In_283,In_638);
nand U1461 (N_1461,In_633,In_647);
xnor U1462 (N_1462,In_42,In_271);
and U1463 (N_1463,In_295,In_441);
xor U1464 (N_1464,In_486,In_277);
nand U1465 (N_1465,In_151,In_739);
nand U1466 (N_1466,In_353,In_455);
nor U1467 (N_1467,In_52,In_424);
and U1468 (N_1468,In_189,In_234);
and U1469 (N_1469,In_565,In_673);
and U1470 (N_1470,In_187,In_151);
nor U1471 (N_1471,In_83,In_80);
and U1472 (N_1472,In_571,In_439);
nand U1473 (N_1473,In_194,In_114);
nor U1474 (N_1474,In_108,In_678);
and U1475 (N_1475,In_58,In_724);
nand U1476 (N_1476,In_385,In_636);
nor U1477 (N_1477,In_708,In_251);
or U1478 (N_1478,In_174,In_722);
xor U1479 (N_1479,In_677,In_651);
nor U1480 (N_1480,In_533,In_662);
xor U1481 (N_1481,In_135,In_432);
or U1482 (N_1482,In_121,In_645);
nand U1483 (N_1483,In_569,In_243);
nor U1484 (N_1484,In_414,In_392);
xnor U1485 (N_1485,In_203,In_274);
nor U1486 (N_1486,In_92,In_273);
xnor U1487 (N_1487,In_443,In_444);
and U1488 (N_1488,In_421,In_285);
nand U1489 (N_1489,In_526,In_210);
xor U1490 (N_1490,In_636,In_527);
nor U1491 (N_1491,In_196,In_481);
or U1492 (N_1492,In_416,In_744);
xor U1493 (N_1493,In_148,In_251);
nor U1494 (N_1494,In_695,In_726);
nand U1495 (N_1495,In_246,In_411);
nand U1496 (N_1496,In_627,In_221);
or U1497 (N_1497,In_313,In_370);
and U1498 (N_1498,In_647,In_141);
or U1499 (N_1499,In_307,In_377);
or U1500 (N_1500,In_88,In_346);
and U1501 (N_1501,In_689,In_598);
or U1502 (N_1502,In_193,In_532);
nor U1503 (N_1503,In_656,In_485);
nor U1504 (N_1504,In_32,In_559);
or U1505 (N_1505,In_176,In_168);
xor U1506 (N_1506,In_276,In_96);
nand U1507 (N_1507,In_252,In_96);
nand U1508 (N_1508,In_668,In_304);
and U1509 (N_1509,In_75,In_321);
and U1510 (N_1510,In_419,In_385);
and U1511 (N_1511,In_733,In_639);
nand U1512 (N_1512,In_507,In_158);
and U1513 (N_1513,In_497,In_465);
or U1514 (N_1514,In_143,In_88);
xnor U1515 (N_1515,In_344,In_280);
nand U1516 (N_1516,In_286,In_44);
xnor U1517 (N_1517,In_302,In_681);
and U1518 (N_1518,In_385,In_506);
and U1519 (N_1519,In_127,In_300);
nand U1520 (N_1520,In_387,In_445);
or U1521 (N_1521,In_145,In_19);
nor U1522 (N_1522,In_715,In_438);
xnor U1523 (N_1523,In_63,In_207);
or U1524 (N_1524,In_197,In_655);
and U1525 (N_1525,In_575,In_3);
nand U1526 (N_1526,In_177,In_218);
and U1527 (N_1527,In_212,In_657);
or U1528 (N_1528,In_699,In_466);
nand U1529 (N_1529,In_386,In_362);
nor U1530 (N_1530,In_120,In_130);
nand U1531 (N_1531,In_365,In_460);
or U1532 (N_1532,In_14,In_564);
or U1533 (N_1533,In_405,In_695);
xor U1534 (N_1534,In_103,In_537);
nor U1535 (N_1535,In_115,In_182);
or U1536 (N_1536,In_70,In_235);
nor U1537 (N_1537,In_53,In_348);
or U1538 (N_1538,In_354,In_669);
nor U1539 (N_1539,In_530,In_129);
and U1540 (N_1540,In_204,In_107);
nor U1541 (N_1541,In_127,In_258);
nor U1542 (N_1542,In_47,In_495);
nor U1543 (N_1543,In_678,In_246);
nand U1544 (N_1544,In_273,In_483);
xnor U1545 (N_1545,In_469,In_600);
nand U1546 (N_1546,In_498,In_179);
xor U1547 (N_1547,In_312,In_604);
and U1548 (N_1548,In_133,In_743);
or U1549 (N_1549,In_328,In_646);
nor U1550 (N_1550,In_396,In_167);
nand U1551 (N_1551,In_698,In_293);
and U1552 (N_1552,In_710,In_590);
or U1553 (N_1553,In_211,In_507);
or U1554 (N_1554,In_408,In_324);
and U1555 (N_1555,In_416,In_138);
xor U1556 (N_1556,In_111,In_209);
nor U1557 (N_1557,In_518,In_538);
xor U1558 (N_1558,In_164,In_405);
and U1559 (N_1559,In_276,In_347);
xnor U1560 (N_1560,In_672,In_180);
nand U1561 (N_1561,In_437,In_588);
and U1562 (N_1562,In_435,In_644);
or U1563 (N_1563,In_389,In_667);
or U1564 (N_1564,In_359,In_207);
nor U1565 (N_1565,In_141,In_184);
or U1566 (N_1566,In_635,In_716);
and U1567 (N_1567,In_68,In_691);
or U1568 (N_1568,In_460,In_147);
xnor U1569 (N_1569,In_96,In_367);
and U1570 (N_1570,In_177,In_206);
and U1571 (N_1571,In_221,In_687);
xnor U1572 (N_1572,In_162,In_97);
nand U1573 (N_1573,In_350,In_701);
xor U1574 (N_1574,In_168,In_214);
xnor U1575 (N_1575,In_170,In_87);
xnor U1576 (N_1576,In_303,In_605);
and U1577 (N_1577,In_571,In_633);
nand U1578 (N_1578,In_644,In_59);
xnor U1579 (N_1579,In_336,In_150);
or U1580 (N_1580,In_11,In_270);
nand U1581 (N_1581,In_218,In_455);
nand U1582 (N_1582,In_9,In_733);
xor U1583 (N_1583,In_245,In_225);
xor U1584 (N_1584,In_483,In_216);
nor U1585 (N_1585,In_123,In_396);
nand U1586 (N_1586,In_661,In_15);
and U1587 (N_1587,In_468,In_301);
nor U1588 (N_1588,In_3,In_94);
xor U1589 (N_1589,In_30,In_487);
nor U1590 (N_1590,In_177,In_135);
and U1591 (N_1591,In_372,In_615);
nor U1592 (N_1592,In_587,In_113);
and U1593 (N_1593,In_606,In_305);
nor U1594 (N_1594,In_116,In_621);
nor U1595 (N_1595,In_143,In_357);
or U1596 (N_1596,In_180,In_593);
nor U1597 (N_1597,In_136,In_198);
nor U1598 (N_1598,In_597,In_122);
nand U1599 (N_1599,In_542,In_224);
or U1600 (N_1600,In_397,In_579);
nor U1601 (N_1601,In_96,In_468);
or U1602 (N_1602,In_655,In_187);
and U1603 (N_1603,In_447,In_563);
nand U1604 (N_1604,In_455,In_319);
nor U1605 (N_1605,In_300,In_193);
and U1606 (N_1606,In_27,In_521);
and U1607 (N_1607,In_160,In_354);
nand U1608 (N_1608,In_368,In_277);
or U1609 (N_1609,In_657,In_345);
or U1610 (N_1610,In_391,In_420);
xnor U1611 (N_1611,In_675,In_618);
or U1612 (N_1612,In_367,In_642);
xor U1613 (N_1613,In_585,In_321);
xnor U1614 (N_1614,In_190,In_392);
xnor U1615 (N_1615,In_71,In_24);
nor U1616 (N_1616,In_231,In_429);
nor U1617 (N_1617,In_375,In_647);
nand U1618 (N_1618,In_91,In_644);
or U1619 (N_1619,In_212,In_497);
nor U1620 (N_1620,In_244,In_62);
nand U1621 (N_1621,In_660,In_356);
and U1622 (N_1622,In_741,In_173);
nor U1623 (N_1623,In_529,In_689);
xnor U1624 (N_1624,In_102,In_193);
nand U1625 (N_1625,In_354,In_580);
and U1626 (N_1626,In_360,In_110);
or U1627 (N_1627,In_673,In_418);
and U1628 (N_1628,In_388,In_480);
nand U1629 (N_1629,In_715,In_165);
xnor U1630 (N_1630,In_500,In_238);
or U1631 (N_1631,In_459,In_287);
nor U1632 (N_1632,In_625,In_305);
nor U1633 (N_1633,In_515,In_438);
nor U1634 (N_1634,In_551,In_694);
and U1635 (N_1635,In_89,In_170);
or U1636 (N_1636,In_338,In_574);
xor U1637 (N_1637,In_132,In_649);
nor U1638 (N_1638,In_671,In_369);
xnor U1639 (N_1639,In_419,In_606);
xor U1640 (N_1640,In_554,In_249);
or U1641 (N_1641,In_641,In_655);
nor U1642 (N_1642,In_6,In_615);
or U1643 (N_1643,In_670,In_305);
and U1644 (N_1644,In_721,In_521);
xnor U1645 (N_1645,In_71,In_525);
nand U1646 (N_1646,In_711,In_47);
xnor U1647 (N_1647,In_18,In_533);
nor U1648 (N_1648,In_541,In_292);
and U1649 (N_1649,In_512,In_689);
xor U1650 (N_1650,In_721,In_276);
or U1651 (N_1651,In_165,In_173);
nor U1652 (N_1652,In_181,In_395);
nand U1653 (N_1653,In_564,In_76);
or U1654 (N_1654,In_336,In_7);
and U1655 (N_1655,In_449,In_692);
and U1656 (N_1656,In_513,In_148);
nor U1657 (N_1657,In_8,In_397);
nor U1658 (N_1658,In_101,In_596);
nor U1659 (N_1659,In_34,In_547);
nor U1660 (N_1660,In_275,In_580);
nand U1661 (N_1661,In_212,In_495);
nand U1662 (N_1662,In_306,In_116);
nand U1663 (N_1663,In_217,In_70);
nor U1664 (N_1664,In_187,In_324);
xor U1665 (N_1665,In_370,In_694);
xnor U1666 (N_1666,In_297,In_363);
or U1667 (N_1667,In_732,In_664);
xor U1668 (N_1668,In_250,In_210);
nor U1669 (N_1669,In_416,In_158);
or U1670 (N_1670,In_583,In_71);
and U1671 (N_1671,In_733,In_358);
or U1672 (N_1672,In_472,In_344);
xor U1673 (N_1673,In_589,In_554);
xnor U1674 (N_1674,In_290,In_634);
nor U1675 (N_1675,In_634,In_321);
or U1676 (N_1676,In_297,In_182);
and U1677 (N_1677,In_652,In_642);
xnor U1678 (N_1678,In_464,In_181);
nand U1679 (N_1679,In_649,In_17);
nand U1680 (N_1680,In_145,In_593);
nor U1681 (N_1681,In_706,In_683);
nand U1682 (N_1682,In_151,In_75);
xor U1683 (N_1683,In_537,In_307);
or U1684 (N_1684,In_234,In_216);
nand U1685 (N_1685,In_691,In_522);
or U1686 (N_1686,In_720,In_212);
and U1687 (N_1687,In_331,In_185);
nor U1688 (N_1688,In_413,In_314);
nand U1689 (N_1689,In_293,In_289);
or U1690 (N_1690,In_79,In_12);
nand U1691 (N_1691,In_720,In_288);
and U1692 (N_1692,In_584,In_637);
xor U1693 (N_1693,In_35,In_486);
nand U1694 (N_1694,In_472,In_132);
xor U1695 (N_1695,In_553,In_615);
xnor U1696 (N_1696,In_84,In_383);
xnor U1697 (N_1697,In_728,In_628);
xnor U1698 (N_1698,In_701,In_122);
or U1699 (N_1699,In_609,In_516);
or U1700 (N_1700,In_551,In_241);
nor U1701 (N_1701,In_464,In_470);
or U1702 (N_1702,In_7,In_471);
xor U1703 (N_1703,In_307,In_572);
nor U1704 (N_1704,In_120,In_278);
nor U1705 (N_1705,In_588,In_68);
nor U1706 (N_1706,In_62,In_290);
nor U1707 (N_1707,In_475,In_121);
or U1708 (N_1708,In_685,In_635);
nand U1709 (N_1709,In_642,In_355);
xor U1710 (N_1710,In_617,In_444);
nor U1711 (N_1711,In_697,In_289);
nand U1712 (N_1712,In_414,In_8);
and U1713 (N_1713,In_639,In_186);
nor U1714 (N_1714,In_205,In_634);
xnor U1715 (N_1715,In_301,In_665);
nand U1716 (N_1716,In_68,In_298);
or U1717 (N_1717,In_111,In_47);
nor U1718 (N_1718,In_349,In_62);
nor U1719 (N_1719,In_117,In_139);
nand U1720 (N_1720,In_397,In_667);
and U1721 (N_1721,In_284,In_430);
nand U1722 (N_1722,In_442,In_568);
and U1723 (N_1723,In_84,In_450);
nor U1724 (N_1724,In_73,In_742);
or U1725 (N_1725,In_446,In_593);
nand U1726 (N_1726,In_70,In_5);
nand U1727 (N_1727,In_126,In_161);
or U1728 (N_1728,In_75,In_559);
and U1729 (N_1729,In_732,In_543);
and U1730 (N_1730,In_609,In_374);
nor U1731 (N_1731,In_373,In_365);
xor U1732 (N_1732,In_76,In_617);
nor U1733 (N_1733,In_263,In_164);
nor U1734 (N_1734,In_731,In_328);
and U1735 (N_1735,In_653,In_643);
nand U1736 (N_1736,In_180,In_470);
and U1737 (N_1737,In_136,In_14);
or U1738 (N_1738,In_745,In_533);
or U1739 (N_1739,In_391,In_532);
xor U1740 (N_1740,In_427,In_324);
xnor U1741 (N_1741,In_220,In_141);
nand U1742 (N_1742,In_15,In_419);
nand U1743 (N_1743,In_67,In_429);
nor U1744 (N_1744,In_206,In_338);
nor U1745 (N_1745,In_659,In_112);
nand U1746 (N_1746,In_227,In_416);
or U1747 (N_1747,In_41,In_571);
nor U1748 (N_1748,In_362,In_487);
nor U1749 (N_1749,In_484,In_311);
and U1750 (N_1750,In_725,In_532);
xnor U1751 (N_1751,In_392,In_562);
nor U1752 (N_1752,In_134,In_55);
nor U1753 (N_1753,In_79,In_481);
or U1754 (N_1754,In_96,In_666);
nand U1755 (N_1755,In_36,In_220);
nand U1756 (N_1756,In_519,In_410);
xnor U1757 (N_1757,In_317,In_287);
or U1758 (N_1758,In_30,In_734);
xor U1759 (N_1759,In_401,In_612);
and U1760 (N_1760,In_641,In_583);
nor U1761 (N_1761,In_74,In_445);
nand U1762 (N_1762,In_669,In_315);
or U1763 (N_1763,In_205,In_111);
nor U1764 (N_1764,In_153,In_681);
nand U1765 (N_1765,In_742,In_30);
and U1766 (N_1766,In_637,In_744);
nor U1767 (N_1767,In_108,In_365);
xor U1768 (N_1768,In_116,In_574);
and U1769 (N_1769,In_237,In_92);
nand U1770 (N_1770,In_460,In_252);
and U1771 (N_1771,In_267,In_241);
xnor U1772 (N_1772,In_25,In_528);
and U1773 (N_1773,In_126,In_69);
nor U1774 (N_1774,In_317,In_712);
xnor U1775 (N_1775,In_646,In_749);
nand U1776 (N_1776,In_251,In_285);
or U1777 (N_1777,In_397,In_262);
nand U1778 (N_1778,In_350,In_159);
or U1779 (N_1779,In_236,In_11);
nand U1780 (N_1780,In_560,In_673);
or U1781 (N_1781,In_184,In_680);
or U1782 (N_1782,In_355,In_395);
or U1783 (N_1783,In_191,In_124);
or U1784 (N_1784,In_195,In_485);
xor U1785 (N_1785,In_128,In_257);
or U1786 (N_1786,In_227,In_741);
or U1787 (N_1787,In_47,In_421);
nand U1788 (N_1788,In_506,In_699);
nand U1789 (N_1789,In_2,In_214);
or U1790 (N_1790,In_567,In_440);
or U1791 (N_1791,In_290,In_38);
xor U1792 (N_1792,In_742,In_714);
xor U1793 (N_1793,In_329,In_272);
nand U1794 (N_1794,In_205,In_335);
xnor U1795 (N_1795,In_447,In_428);
nand U1796 (N_1796,In_328,In_69);
nand U1797 (N_1797,In_259,In_421);
or U1798 (N_1798,In_115,In_438);
nand U1799 (N_1799,In_532,In_466);
nor U1800 (N_1800,In_10,In_1);
nor U1801 (N_1801,In_67,In_410);
xnor U1802 (N_1802,In_694,In_287);
nand U1803 (N_1803,In_600,In_714);
nand U1804 (N_1804,In_228,In_239);
xor U1805 (N_1805,In_150,In_479);
xor U1806 (N_1806,In_380,In_743);
or U1807 (N_1807,In_238,In_14);
nor U1808 (N_1808,In_287,In_196);
xor U1809 (N_1809,In_515,In_212);
nand U1810 (N_1810,In_588,In_125);
nor U1811 (N_1811,In_624,In_362);
nand U1812 (N_1812,In_120,In_653);
nor U1813 (N_1813,In_313,In_293);
nand U1814 (N_1814,In_29,In_84);
nand U1815 (N_1815,In_463,In_72);
xnor U1816 (N_1816,In_475,In_237);
nand U1817 (N_1817,In_87,In_643);
or U1818 (N_1818,In_653,In_210);
or U1819 (N_1819,In_264,In_669);
nand U1820 (N_1820,In_494,In_394);
nor U1821 (N_1821,In_185,In_223);
or U1822 (N_1822,In_640,In_261);
and U1823 (N_1823,In_508,In_576);
nand U1824 (N_1824,In_561,In_549);
nor U1825 (N_1825,In_742,In_725);
nor U1826 (N_1826,In_545,In_650);
or U1827 (N_1827,In_529,In_268);
and U1828 (N_1828,In_731,In_285);
and U1829 (N_1829,In_715,In_520);
and U1830 (N_1830,In_280,In_745);
xor U1831 (N_1831,In_412,In_474);
nand U1832 (N_1832,In_203,In_22);
xnor U1833 (N_1833,In_275,In_176);
nand U1834 (N_1834,In_247,In_689);
or U1835 (N_1835,In_242,In_83);
or U1836 (N_1836,In_279,In_372);
nor U1837 (N_1837,In_128,In_222);
nand U1838 (N_1838,In_398,In_224);
nor U1839 (N_1839,In_90,In_441);
or U1840 (N_1840,In_29,In_188);
xor U1841 (N_1841,In_97,In_109);
xor U1842 (N_1842,In_280,In_357);
nor U1843 (N_1843,In_377,In_583);
or U1844 (N_1844,In_738,In_575);
and U1845 (N_1845,In_120,In_572);
nand U1846 (N_1846,In_380,In_551);
and U1847 (N_1847,In_634,In_264);
or U1848 (N_1848,In_245,In_298);
or U1849 (N_1849,In_46,In_16);
and U1850 (N_1850,In_209,In_156);
and U1851 (N_1851,In_691,In_518);
nor U1852 (N_1852,In_731,In_170);
nand U1853 (N_1853,In_719,In_217);
nor U1854 (N_1854,In_338,In_115);
xnor U1855 (N_1855,In_189,In_634);
nor U1856 (N_1856,In_619,In_329);
and U1857 (N_1857,In_685,In_476);
xor U1858 (N_1858,In_539,In_399);
nand U1859 (N_1859,In_164,In_420);
or U1860 (N_1860,In_335,In_527);
xor U1861 (N_1861,In_500,In_611);
xor U1862 (N_1862,In_516,In_86);
nor U1863 (N_1863,In_687,In_56);
nor U1864 (N_1864,In_100,In_505);
or U1865 (N_1865,In_532,In_395);
xor U1866 (N_1866,In_503,In_38);
nor U1867 (N_1867,In_124,In_182);
or U1868 (N_1868,In_190,In_222);
and U1869 (N_1869,In_291,In_117);
and U1870 (N_1870,In_546,In_512);
and U1871 (N_1871,In_305,In_251);
nor U1872 (N_1872,In_522,In_488);
nor U1873 (N_1873,In_664,In_656);
nand U1874 (N_1874,In_686,In_610);
or U1875 (N_1875,In_23,In_742);
nand U1876 (N_1876,In_372,In_312);
nand U1877 (N_1877,In_725,In_94);
nor U1878 (N_1878,In_48,In_224);
xor U1879 (N_1879,In_744,In_594);
nor U1880 (N_1880,In_393,In_531);
or U1881 (N_1881,In_376,In_720);
xor U1882 (N_1882,In_583,In_102);
or U1883 (N_1883,In_666,In_95);
xor U1884 (N_1884,In_458,In_150);
and U1885 (N_1885,In_230,In_542);
and U1886 (N_1886,In_342,In_351);
or U1887 (N_1887,In_216,In_703);
and U1888 (N_1888,In_573,In_679);
nor U1889 (N_1889,In_291,In_185);
xnor U1890 (N_1890,In_395,In_412);
or U1891 (N_1891,In_604,In_31);
nand U1892 (N_1892,In_133,In_452);
xor U1893 (N_1893,In_75,In_275);
and U1894 (N_1894,In_467,In_427);
nor U1895 (N_1895,In_37,In_193);
nand U1896 (N_1896,In_170,In_685);
nor U1897 (N_1897,In_401,In_286);
nor U1898 (N_1898,In_567,In_457);
and U1899 (N_1899,In_327,In_260);
nand U1900 (N_1900,In_548,In_492);
xnor U1901 (N_1901,In_484,In_520);
nor U1902 (N_1902,In_285,In_64);
or U1903 (N_1903,In_712,In_140);
or U1904 (N_1904,In_727,In_655);
xor U1905 (N_1905,In_536,In_302);
nand U1906 (N_1906,In_579,In_24);
nand U1907 (N_1907,In_170,In_668);
xnor U1908 (N_1908,In_95,In_605);
nand U1909 (N_1909,In_439,In_446);
and U1910 (N_1910,In_474,In_66);
xnor U1911 (N_1911,In_634,In_433);
nand U1912 (N_1912,In_285,In_351);
xor U1913 (N_1913,In_440,In_379);
and U1914 (N_1914,In_52,In_404);
xnor U1915 (N_1915,In_135,In_669);
nor U1916 (N_1916,In_650,In_281);
or U1917 (N_1917,In_285,In_223);
and U1918 (N_1918,In_720,In_702);
xor U1919 (N_1919,In_436,In_30);
nand U1920 (N_1920,In_359,In_126);
nor U1921 (N_1921,In_57,In_284);
nand U1922 (N_1922,In_689,In_1);
nor U1923 (N_1923,In_1,In_342);
or U1924 (N_1924,In_544,In_511);
or U1925 (N_1925,In_47,In_596);
xnor U1926 (N_1926,In_696,In_678);
xnor U1927 (N_1927,In_681,In_106);
or U1928 (N_1928,In_30,In_704);
nor U1929 (N_1929,In_366,In_732);
xnor U1930 (N_1930,In_230,In_166);
and U1931 (N_1931,In_42,In_697);
or U1932 (N_1932,In_649,In_670);
and U1933 (N_1933,In_80,In_6);
nor U1934 (N_1934,In_220,In_227);
or U1935 (N_1935,In_417,In_226);
nand U1936 (N_1936,In_590,In_565);
nand U1937 (N_1937,In_131,In_341);
xnor U1938 (N_1938,In_555,In_243);
and U1939 (N_1939,In_526,In_79);
xnor U1940 (N_1940,In_644,In_115);
nor U1941 (N_1941,In_194,In_728);
nor U1942 (N_1942,In_315,In_250);
xnor U1943 (N_1943,In_400,In_179);
or U1944 (N_1944,In_612,In_520);
xor U1945 (N_1945,In_76,In_505);
or U1946 (N_1946,In_337,In_209);
and U1947 (N_1947,In_53,In_311);
xor U1948 (N_1948,In_491,In_503);
xnor U1949 (N_1949,In_428,In_131);
xor U1950 (N_1950,In_532,In_401);
or U1951 (N_1951,In_361,In_353);
or U1952 (N_1952,In_565,In_515);
nand U1953 (N_1953,In_236,In_387);
nand U1954 (N_1954,In_220,In_603);
nor U1955 (N_1955,In_516,In_278);
and U1956 (N_1956,In_643,In_167);
and U1957 (N_1957,In_527,In_515);
or U1958 (N_1958,In_562,In_81);
nor U1959 (N_1959,In_255,In_25);
and U1960 (N_1960,In_108,In_478);
and U1961 (N_1961,In_73,In_628);
nor U1962 (N_1962,In_304,In_552);
nor U1963 (N_1963,In_531,In_284);
nor U1964 (N_1964,In_691,In_22);
nand U1965 (N_1965,In_277,In_527);
xnor U1966 (N_1966,In_570,In_360);
xor U1967 (N_1967,In_19,In_171);
nor U1968 (N_1968,In_205,In_660);
and U1969 (N_1969,In_594,In_37);
xnor U1970 (N_1970,In_660,In_305);
or U1971 (N_1971,In_153,In_316);
and U1972 (N_1972,In_649,In_399);
or U1973 (N_1973,In_186,In_30);
and U1974 (N_1974,In_392,In_613);
or U1975 (N_1975,In_374,In_31);
nand U1976 (N_1976,In_35,In_93);
xnor U1977 (N_1977,In_130,In_53);
and U1978 (N_1978,In_611,In_221);
nor U1979 (N_1979,In_579,In_445);
nand U1980 (N_1980,In_219,In_400);
nand U1981 (N_1981,In_224,In_574);
xnor U1982 (N_1982,In_290,In_431);
or U1983 (N_1983,In_694,In_73);
nand U1984 (N_1984,In_328,In_355);
nor U1985 (N_1985,In_383,In_136);
or U1986 (N_1986,In_195,In_331);
nor U1987 (N_1987,In_142,In_339);
or U1988 (N_1988,In_657,In_119);
xnor U1989 (N_1989,In_407,In_351);
nor U1990 (N_1990,In_20,In_1);
or U1991 (N_1991,In_351,In_723);
xnor U1992 (N_1992,In_127,In_416);
and U1993 (N_1993,In_96,In_553);
or U1994 (N_1994,In_163,In_682);
and U1995 (N_1995,In_29,In_141);
nor U1996 (N_1996,In_620,In_334);
and U1997 (N_1997,In_451,In_353);
and U1998 (N_1998,In_349,In_130);
xor U1999 (N_1999,In_510,In_598);
or U2000 (N_2000,In_105,In_24);
nand U2001 (N_2001,In_530,In_397);
xor U2002 (N_2002,In_673,In_678);
and U2003 (N_2003,In_415,In_384);
xor U2004 (N_2004,In_608,In_709);
nor U2005 (N_2005,In_362,In_149);
or U2006 (N_2006,In_509,In_343);
or U2007 (N_2007,In_609,In_700);
nand U2008 (N_2008,In_103,In_559);
xor U2009 (N_2009,In_370,In_189);
or U2010 (N_2010,In_249,In_312);
and U2011 (N_2011,In_198,In_55);
xnor U2012 (N_2012,In_589,In_246);
nand U2013 (N_2013,In_93,In_573);
or U2014 (N_2014,In_323,In_725);
nor U2015 (N_2015,In_371,In_466);
nand U2016 (N_2016,In_138,In_422);
or U2017 (N_2017,In_603,In_577);
nand U2018 (N_2018,In_621,In_417);
xnor U2019 (N_2019,In_623,In_404);
nor U2020 (N_2020,In_267,In_276);
xor U2021 (N_2021,In_496,In_377);
and U2022 (N_2022,In_223,In_49);
xnor U2023 (N_2023,In_594,In_408);
xnor U2024 (N_2024,In_592,In_76);
xnor U2025 (N_2025,In_506,In_548);
nand U2026 (N_2026,In_722,In_310);
nand U2027 (N_2027,In_251,In_311);
nand U2028 (N_2028,In_390,In_205);
and U2029 (N_2029,In_703,In_207);
nor U2030 (N_2030,In_573,In_358);
nor U2031 (N_2031,In_315,In_497);
nor U2032 (N_2032,In_63,In_352);
nand U2033 (N_2033,In_639,In_349);
xnor U2034 (N_2034,In_359,In_409);
nor U2035 (N_2035,In_725,In_89);
and U2036 (N_2036,In_702,In_190);
xnor U2037 (N_2037,In_411,In_36);
and U2038 (N_2038,In_65,In_388);
and U2039 (N_2039,In_206,In_449);
nand U2040 (N_2040,In_273,In_627);
nand U2041 (N_2041,In_176,In_30);
nand U2042 (N_2042,In_567,In_586);
nand U2043 (N_2043,In_509,In_643);
or U2044 (N_2044,In_624,In_383);
and U2045 (N_2045,In_312,In_131);
and U2046 (N_2046,In_159,In_112);
and U2047 (N_2047,In_537,In_162);
and U2048 (N_2048,In_223,In_409);
or U2049 (N_2049,In_534,In_498);
nand U2050 (N_2050,In_691,In_311);
nor U2051 (N_2051,In_422,In_415);
nand U2052 (N_2052,In_369,In_119);
or U2053 (N_2053,In_340,In_453);
and U2054 (N_2054,In_349,In_41);
xor U2055 (N_2055,In_596,In_725);
nand U2056 (N_2056,In_371,In_444);
xnor U2057 (N_2057,In_635,In_293);
nor U2058 (N_2058,In_278,In_19);
nor U2059 (N_2059,In_142,In_70);
nand U2060 (N_2060,In_401,In_257);
nor U2061 (N_2061,In_609,In_697);
nor U2062 (N_2062,In_117,In_622);
nor U2063 (N_2063,In_652,In_5);
xnor U2064 (N_2064,In_188,In_401);
and U2065 (N_2065,In_523,In_487);
or U2066 (N_2066,In_493,In_488);
and U2067 (N_2067,In_726,In_596);
xnor U2068 (N_2068,In_291,In_426);
nand U2069 (N_2069,In_110,In_156);
nor U2070 (N_2070,In_239,In_568);
or U2071 (N_2071,In_114,In_684);
xor U2072 (N_2072,In_420,In_212);
nand U2073 (N_2073,In_65,In_739);
nor U2074 (N_2074,In_511,In_685);
xor U2075 (N_2075,In_655,In_650);
nor U2076 (N_2076,In_532,In_289);
or U2077 (N_2077,In_224,In_556);
and U2078 (N_2078,In_403,In_317);
xor U2079 (N_2079,In_32,In_645);
nand U2080 (N_2080,In_251,In_254);
xor U2081 (N_2081,In_242,In_186);
xor U2082 (N_2082,In_117,In_318);
nand U2083 (N_2083,In_232,In_188);
or U2084 (N_2084,In_721,In_123);
xnor U2085 (N_2085,In_710,In_730);
and U2086 (N_2086,In_102,In_556);
and U2087 (N_2087,In_711,In_272);
and U2088 (N_2088,In_121,In_585);
xor U2089 (N_2089,In_503,In_47);
nand U2090 (N_2090,In_242,In_499);
xnor U2091 (N_2091,In_239,In_580);
and U2092 (N_2092,In_21,In_667);
nor U2093 (N_2093,In_57,In_249);
xor U2094 (N_2094,In_253,In_660);
nand U2095 (N_2095,In_100,In_671);
xnor U2096 (N_2096,In_87,In_122);
and U2097 (N_2097,In_604,In_731);
or U2098 (N_2098,In_727,In_244);
or U2099 (N_2099,In_10,In_441);
nand U2100 (N_2100,In_613,In_705);
xnor U2101 (N_2101,In_629,In_624);
nand U2102 (N_2102,In_172,In_559);
nand U2103 (N_2103,In_223,In_80);
nor U2104 (N_2104,In_127,In_319);
or U2105 (N_2105,In_296,In_150);
and U2106 (N_2106,In_122,In_744);
nor U2107 (N_2107,In_75,In_241);
nor U2108 (N_2108,In_577,In_163);
or U2109 (N_2109,In_7,In_268);
xor U2110 (N_2110,In_520,In_326);
xnor U2111 (N_2111,In_174,In_597);
nand U2112 (N_2112,In_514,In_221);
and U2113 (N_2113,In_671,In_10);
nor U2114 (N_2114,In_65,In_632);
xnor U2115 (N_2115,In_28,In_459);
nand U2116 (N_2116,In_145,In_391);
nand U2117 (N_2117,In_411,In_585);
or U2118 (N_2118,In_209,In_302);
or U2119 (N_2119,In_430,In_296);
nor U2120 (N_2120,In_472,In_332);
xor U2121 (N_2121,In_167,In_719);
nand U2122 (N_2122,In_118,In_683);
and U2123 (N_2123,In_417,In_334);
nand U2124 (N_2124,In_381,In_172);
and U2125 (N_2125,In_212,In_728);
xnor U2126 (N_2126,In_376,In_49);
or U2127 (N_2127,In_19,In_254);
xor U2128 (N_2128,In_562,In_243);
and U2129 (N_2129,In_562,In_276);
nor U2130 (N_2130,In_463,In_140);
or U2131 (N_2131,In_478,In_577);
xor U2132 (N_2132,In_21,In_643);
xnor U2133 (N_2133,In_509,In_693);
or U2134 (N_2134,In_170,In_249);
or U2135 (N_2135,In_14,In_83);
or U2136 (N_2136,In_470,In_729);
nand U2137 (N_2137,In_306,In_500);
and U2138 (N_2138,In_317,In_393);
nor U2139 (N_2139,In_30,In_146);
xnor U2140 (N_2140,In_345,In_650);
and U2141 (N_2141,In_677,In_600);
and U2142 (N_2142,In_17,In_197);
nor U2143 (N_2143,In_100,In_346);
and U2144 (N_2144,In_428,In_617);
or U2145 (N_2145,In_570,In_477);
xor U2146 (N_2146,In_420,In_649);
and U2147 (N_2147,In_214,In_178);
or U2148 (N_2148,In_311,In_257);
nor U2149 (N_2149,In_33,In_191);
nor U2150 (N_2150,In_642,In_263);
nand U2151 (N_2151,In_671,In_550);
and U2152 (N_2152,In_527,In_235);
nand U2153 (N_2153,In_460,In_543);
and U2154 (N_2154,In_469,In_34);
nor U2155 (N_2155,In_322,In_527);
nor U2156 (N_2156,In_330,In_355);
and U2157 (N_2157,In_502,In_351);
nor U2158 (N_2158,In_132,In_572);
or U2159 (N_2159,In_179,In_584);
nand U2160 (N_2160,In_162,In_497);
xor U2161 (N_2161,In_189,In_226);
or U2162 (N_2162,In_690,In_463);
xnor U2163 (N_2163,In_356,In_104);
and U2164 (N_2164,In_149,In_269);
or U2165 (N_2165,In_300,In_697);
or U2166 (N_2166,In_475,In_224);
nand U2167 (N_2167,In_671,In_728);
and U2168 (N_2168,In_749,In_743);
xor U2169 (N_2169,In_623,In_349);
xor U2170 (N_2170,In_464,In_629);
and U2171 (N_2171,In_198,In_42);
and U2172 (N_2172,In_431,In_210);
and U2173 (N_2173,In_545,In_47);
and U2174 (N_2174,In_366,In_456);
or U2175 (N_2175,In_308,In_221);
or U2176 (N_2176,In_132,In_618);
nor U2177 (N_2177,In_46,In_705);
or U2178 (N_2178,In_619,In_494);
xor U2179 (N_2179,In_367,In_623);
xnor U2180 (N_2180,In_209,In_705);
or U2181 (N_2181,In_505,In_343);
nand U2182 (N_2182,In_98,In_24);
nor U2183 (N_2183,In_517,In_600);
nor U2184 (N_2184,In_434,In_28);
xor U2185 (N_2185,In_426,In_573);
or U2186 (N_2186,In_336,In_75);
and U2187 (N_2187,In_420,In_205);
and U2188 (N_2188,In_151,In_618);
and U2189 (N_2189,In_137,In_560);
nor U2190 (N_2190,In_635,In_524);
or U2191 (N_2191,In_269,In_132);
xnor U2192 (N_2192,In_454,In_396);
xnor U2193 (N_2193,In_218,In_159);
nand U2194 (N_2194,In_369,In_6);
or U2195 (N_2195,In_529,In_707);
or U2196 (N_2196,In_510,In_511);
nor U2197 (N_2197,In_366,In_275);
and U2198 (N_2198,In_726,In_745);
xnor U2199 (N_2199,In_626,In_678);
xor U2200 (N_2200,In_354,In_245);
nand U2201 (N_2201,In_741,In_7);
and U2202 (N_2202,In_419,In_410);
or U2203 (N_2203,In_462,In_188);
nand U2204 (N_2204,In_77,In_345);
xnor U2205 (N_2205,In_348,In_585);
and U2206 (N_2206,In_736,In_703);
xor U2207 (N_2207,In_461,In_57);
and U2208 (N_2208,In_103,In_396);
nand U2209 (N_2209,In_37,In_135);
nor U2210 (N_2210,In_6,In_193);
nor U2211 (N_2211,In_66,In_546);
xnor U2212 (N_2212,In_637,In_317);
nor U2213 (N_2213,In_269,In_382);
nor U2214 (N_2214,In_126,In_141);
or U2215 (N_2215,In_497,In_483);
xnor U2216 (N_2216,In_547,In_116);
nor U2217 (N_2217,In_327,In_35);
nand U2218 (N_2218,In_421,In_619);
xnor U2219 (N_2219,In_620,In_200);
and U2220 (N_2220,In_241,In_32);
or U2221 (N_2221,In_15,In_546);
nand U2222 (N_2222,In_496,In_44);
xor U2223 (N_2223,In_177,In_189);
nand U2224 (N_2224,In_518,In_331);
nand U2225 (N_2225,In_327,In_489);
or U2226 (N_2226,In_101,In_2);
xor U2227 (N_2227,In_382,In_603);
xor U2228 (N_2228,In_617,In_352);
nand U2229 (N_2229,In_401,In_713);
xor U2230 (N_2230,In_337,In_43);
and U2231 (N_2231,In_629,In_438);
nand U2232 (N_2232,In_61,In_146);
nor U2233 (N_2233,In_79,In_134);
xor U2234 (N_2234,In_26,In_636);
xnor U2235 (N_2235,In_695,In_524);
or U2236 (N_2236,In_222,In_72);
xnor U2237 (N_2237,In_542,In_645);
nand U2238 (N_2238,In_388,In_336);
xnor U2239 (N_2239,In_504,In_420);
or U2240 (N_2240,In_626,In_742);
nor U2241 (N_2241,In_12,In_631);
nand U2242 (N_2242,In_113,In_53);
nand U2243 (N_2243,In_229,In_90);
nor U2244 (N_2244,In_517,In_136);
nor U2245 (N_2245,In_340,In_710);
nor U2246 (N_2246,In_605,In_712);
nor U2247 (N_2247,In_690,In_692);
xnor U2248 (N_2248,In_703,In_436);
nor U2249 (N_2249,In_138,In_84);
xnor U2250 (N_2250,In_137,In_256);
nor U2251 (N_2251,In_14,In_163);
xnor U2252 (N_2252,In_106,In_452);
or U2253 (N_2253,In_578,In_130);
nand U2254 (N_2254,In_617,In_333);
nand U2255 (N_2255,In_48,In_741);
or U2256 (N_2256,In_544,In_114);
nand U2257 (N_2257,In_237,In_626);
or U2258 (N_2258,In_306,In_0);
xnor U2259 (N_2259,In_547,In_444);
xnor U2260 (N_2260,In_430,In_232);
or U2261 (N_2261,In_494,In_518);
or U2262 (N_2262,In_709,In_345);
nand U2263 (N_2263,In_728,In_582);
nand U2264 (N_2264,In_119,In_490);
and U2265 (N_2265,In_482,In_11);
nand U2266 (N_2266,In_175,In_573);
nor U2267 (N_2267,In_649,In_634);
and U2268 (N_2268,In_556,In_554);
or U2269 (N_2269,In_620,In_231);
or U2270 (N_2270,In_656,In_525);
and U2271 (N_2271,In_662,In_478);
nand U2272 (N_2272,In_469,In_95);
nor U2273 (N_2273,In_735,In_588);
nor U2274 (N_2274,In_19,In_271);
and U2275 (N_2275,In_112,In_178);
xnor U2276 (N_2276,In_618,In_269);
nor U2277 (N_2277,In_179,In_349);
nand U2278 (N_2278,In_645,In_91);
or U2279 (N_2279,In_231,In_63);
or U2280 (N_2280,In_395,In_90);
nand U2281 (N_2281,In_324,In_241);
xnor U2282 (N_2282,In_334,In_469);
nand U2283 (N_2283,In_459,In_674);
nor U2284 (N_2284,In_228,In_6);
xor U2285 (N_2285,In_176,In_466);
xnor U2286 (N_2286,In_698,In_455);
nand U2287 (N_2287,In_218,In_82);
xor U2288 (N_2288,In_56,In_184);
nand U2289 (N_2289,In_628,In_626);
nand U2290 (N_2290,In_601,In_450);
nor U2291 (N_2291,In_536,In_509);
nand U2292 (N_2292,In_222,In_570);
nor U2293 (N_2293,In_254,In_640);
and U2294 (N_2294,In_591,In_605);
nand U2295 (N_2295,In_95,In_225);
nand U2296 (N_2296,In_463,In_112);
nor U2297 (N_2297,In_483,In_171);
nor U2298 (N_2298,In_367,In_739);
or U2299 (N_2299,In_563,In_142);
or U2300 (N_2300,In_610,In_229);
nand U2301 (N_2301,In_523,In_197);
and U2302 (N_2302,In_299,In_438);
xor U2303 (N_2303,In_722,In_459);
xnor U2304 (N_2304,In_463,In_663);
nand U2305 (N_2305,In_185,In_141);
and U2306 (N_2306,In_477,In_698);
and U2307 (N_2307,In_285,In_305);
or U2308 (N_2308,In_520,In_460);
nand U2309 (N_2309,In_520,In_270);
and U2310 (N_2310,In_341,In_466);
and U2311 (N_2311,In_575,In_43);
and U2312 (N_2312,In_232,In_601);
nor U2313 (N_2313,In_728,In_718);
or U2314 (N_2314,In_592,In_78);
and U2315 (N_2315,In_583,In_318);
nor U2316 (N_2316,In_425,In_190);
xnor U2317 (N_2317,In_697,In_237);
nor U2318 (N_2318,In_480,In_241);
and U2319 (N_2319,In_360,In_592);
nand U2320 (N_2320,In_470,In_132);
nand U2321 (N_2321,In_615,In_97);
nand U2322 (N_2322,In_272,In_546);
nand U2323 (N_2323,In_731,In_391);
nor U2324 (N_2324,In_395,In_1);
nand U2325 (N_2325,In_581,In_294);
nor U2326 (N_2326,In_607,In_209);
nor U2327 (N_2327,In_145,In_526);
and U2328 (N_2328,In_724,In_628);
nand U2329 (N_2329,In_411,In_182);
or U2330 (N_2330,In_286,In_500);
or U2331 (N_2331,In_369,In_628);
or U2332 (N_2332,In_706,In_559);
or U2333 (N_2333,In_279,In_552);
and U2334 (N_2334,In_492,In_672);
xnor U2335 (N_2335,In_487,In_173);
and U2336 (N_2336,In_218,In_186);
xnor U2337 (N_2337,In_43,In_480);
xnor U2338 (N_2338,In_385,In_367);
xnor U2339 (N_2339,In_309,In_609);
xnor U2340 (N_2340,In_72,In_238);
or U2341 (N_2341,In_104,In_541);
nor U2342 (N_2342,In_428,In_629);
nor U2343 (N_2343,In_363,In_203);
and U2344 (N_2344,In_604,In_207);
or U2345 (N_2345,In_630,In_708);
nand U2346 (N_2346,In_572,In_563);
or U2347 (N_2347,In_675,In_3);
nand U2348 (N_2348,In_302,In_14);
nand U2349 (N_2349,In_180,In_361);
and U2350 (N_2350,In_237,In_214);
nand U2351 (N_2351,In_299,In_174);
xnor U2352 (N_2352,In_616,In_83);
and U2353 (N_2353,In_64,In_680);
nand U2354 (N_2354,In_637,In_377);
xor U2355 (N_2355,In_512,In_83);
nand U2356 (N_2356,In_312,In_644);
or U2357 (N_2357,In_217,In_311);
or U2358 (N_2358,In_464,In_637);
nand U2359 (N_2359,In_151,In_224);
xnor U2360 (N_2360,In_94,In_388);
and U2361 (N_2361,In_744,In_54);
xor U2362 (N_2362,In_285,In_168);
xor U2363 (N_2363,In_445,In_708);
xor U2364 (N_2364,In_39,In_412);
nor U2365 (N_2365,In_553,In_398);
or U2366 (N_2366,In_174,In_678);
and U2367 (N_2367,In_644,In_128);
or U2368 (N_2368,In_240,In_405);
nor U2369 (N_2369,In_284,In_715);
nand U2370 (N_2370,In_645,In_35);
or U2371 (N_2371,In_306,In_285);
nand U2372 (N_2372,In_312,In_53);
or U2373 (N_2373,In_37,In_382);
xor U2374 (N_2374,In_528,In_357);
or U2375 (N_2375,In_82,In_160);
and U2376 (N_2376,In_61,In_226);
and U2377 (N_2377,In_662,In_542);
nand U2378 (N_2378,In_43,In_22);
xor U2379 (N_2379,In_392,In_288);
xor U2380 (N_2380,In_282,In_6);
and U2381 (N_2381,In_395,In_473);
and U2382 (N_2382,In_513,In_560);
nor U2383 (N_2383,In_262,In_106);
or U2384 (N_2384,In_506,In_280);
and U2385 (N_2385,In_401,In_144);
nand U2386 (N_2386,In_743,In_671);
and U2387 (N_2387,In_117,In_505);
nand U2388 (N_2388,In_636,In_73);
and U2389 (N_2389,In_586,In_9);
or U2390 (N_2390,In_196,In_669);
nand U2391 (N_2391,In_75,In_338);
nand U2392 (N_2392,In_644,In_650);
nor U2393 (N_2393,In_700,In_284);
and U2394 (N_2394,In_58,In_218);
and U2395 (N_2395,In_560,In_29);
nand U2396 (N_2396,In_142,In_602);
and U2397 (N_2397,In_328,In_488);
and U2398 (N_2398,In_524,In_142);
nor U2399 (N_2399,In_74,In_355);
or U2400 (N_2400,In_384,In_193);
xor U2401 (N_2401,In_238,In_558);
nand U2402 (N_2402,In_248,In_67);
or U2403 (N_2403,In_554,In_235);
or U2404 (N_2404,In_225,In_130);
or U2405 (N_2405,In_98,In_645);
nor U2406 (N_2406,In_361,In_575);
and U2407 (N_2407,In_281,In_412);
xnor U2408 (N_2408,In_631,In_142);
nor U2409 (N_2409,In_204,In_116);
and U2410 (N_2410,In_415,In_599);
nand U2411 (N_2411,In_392,In_522);
and U2412 (N_2412,In_558,In_549);
and U2413 (N_2413,In_40,In_207);
or U2414 (N_2414,In_161,In_121);
nor U2415 (N_2415,In_725,In_194);
xnor U2416 (N_2416,In_327,In_8);
and U2417 (N_2417,In_547,In_602);
and U2418 (N_2418,In_460,In_559);
nand U2419 (N_2419,In_285,In_116);
nand U2420 (N_2420,In_99,In_84);
xor U2421 (N_2421,In_314,In_442);
nand U2422 (N_2422,In_497,In_680);
and U2423 (N_2423,In_688,In_114);
nand U2424 (N_2424,In_727,In_503);
nor U2425 (N_2425,In_159,In_431);
nand U2426 (N_2426,In_10,In_304);
nor U2427 (N_2427,In_121,In_264);
nand U2428 (N_2428,In_369,In_740);
nor U2429 (N_2429,In_433,In_747);
and U2430 (N_2430,In_303,In_708);
nor U2431 (N_2431,In_386,In_141);
nand U2432 (N_2432,In_471,In_403);
and U2433 (N_2433,In_161,In_283);
xor U2434 (N_2434,In_187,In_83);
nor U2435 (N_2435,In_157,In_159);
or U2436 (N_2436,In_319,In_314);
nand U2437 (N_2437,In_101,In_163);
nor U2438 (N_2438,In_344,In_630);
nand U2439 (N_2439,In_684,In_369);
nand U2440 (N_2440,In_419,In_452);
nand U2441 (N_2441,In_342,In_194);
xnor U2442 (N_2442,In_80,In_525);
or U2443 (N_2443,In_246,In_115);
and U2444 (N_2444,In_673,In_702);
nand U2445 (N_2445,In_220,In_562);
nor U2446 (N_2446,In_20,In_285);
or U2447 (N_2447,In_53,In_361);
nor U2448 (N_2448,In_659,In_40);
and U2449 (N_2449,In_558,In_345);
or U2450 (N_2450,In_189,In_347);
nand U2451 (N_2451,In_465,In_691);
xor U2452 (N_2452,In_662,In_401);
nand U2453 (N_2453,In_431,In_309);
xnor U2454 (N_2454,In_124,In_556);
and U2455 (N_2455,In_87,In_683);
xnor U2456 (N_2456,In_701,In_35);
xor U2457 (N_2457,In_163,In_238);
or U2458 (N_2458,In_437,In_577);
xor U2459 (N_2459,In_582,In_605);
or U2460 (N_2460,In_86,In_628);
xor U2461 (N_2461,In_332,In_609);
xor U2462 (N_2462,In_244,In_86);
nand U2463 (N_2463,In_353,In_513);
and U2464 (N_2464,In_36,In_305);
nor U2465 (N_2465,In_210,In_505);
nor U2466 (N_2466,In_204,In_135);
nand U2467 (N_2467,In_90,In_560);
or U2468 (N_2468,In_200,In_275);
nand U2469 (N_2469,In_199,In_489);
and U2470 (N_2470,In_372,In_590);
nor U2471 (N_2471,In_348,In_260);
nor U2472 (N_2472,In_295,In_533);
and U2473 (N_2473,In_607,In_721);
and U2474 (N_2474,In_232,In_642);
xnor U2475 (N_2475,In_464,In_54);
or U2476 (N_2476,In_25,In_271);
and U2477 (N_2477,In_333,In_340);
and U2478 (N_2478,In_69,In_82);
nor U2479 (N_2479,In_17,In_144);
xnor U2480 (N_2480,In_495,In_64);
or U2481 (N_2481,In_503,In_164);
nand U2482 (N_2482,In_560,In_81);
or U2483 (N_2483,In_123,In_346);
nand U2484 (N_2484,In_72,In_156);
xor U2485 (N_2485,In_542,In_20);
xor U2486 (N_2486,In_420,In_295);
nand U2487 (N_2487,In_713,In_726);
xnor U2488 (N_2488,In_28,In_24);
nand U2489 (N_2489,In_543,In_220);
and U2490 (N_2490,In_317,In_30);
nor U2491 (N_2491,In_682,In_311);
nand U2492 (N_2492,In_228,In_265);
nor U2493 (N_2493,In_737,In_471);
xnor U2494 (N_2494,In_567,In_75);
xor U2495 (N_2495,In_658,In_161);
nand U2496 (N_2496,In_28,In_155);
xor U2497 (N_2497,In_291,In_723);
nand U2498 (N_2498,In_6,In_3);
nor U2499 (N_2499,In_724,In_696);
nand U2500 (N_2500,N_944,N_973);
nand U2501 (N_2501,N_118,N_2398);
nand U2502 (N_2502,N_524,N_1405);
and U2503 (N_2503,N_1533,N_375);
or U2504 (N_2504,N_2056,N_999);
nor U2505 (N_2505,N_1613,N_1300);
nand U2506 (N_2506,N_1386,N_2345);
nand U2507 (N_2507,N_691,N_1628);
or U2508 (N_2508,N_2144,N_1189);
nor U2509 (N_2509,N_210,N_2491);
or U2510 (N_2510,N_702,N_78);
xnor U2511 (N_2511,N_2153,N_1426);
xor U2512 (N_2512,N_211,N_2011);
or U2513 (N_2513,N_615,N_892);
or U2514 (N_2514,N_161,N_1511);
nand U2515 (N_2515,N_618,N_522);
xor U2516 (N_2516,N_247,N_1507);
nand U2517 (N_2517,N_2361,N_1281);
and U2518 (N_2518,N_1732,N_1453);
nor U2519 (N_2519,N_2162,N_1124);
xor U2520 (N_2520,N_435,N_1761);
xnor U2521 (N_2521,N_170,N_769);
nor U2522 (N_2522,N_2040,N_826);
or U2523 (N_2523,N_560,N_1471);
xor U2524 (N_2524,N_955,N_1152);
xor U2525 (N_2525,N_1747,N_1530);
xor U2526 (N_2526,N_214,N_1457);
nor U2527 (N_2527,N_2081,N_94);
nor U2528 (N_2528,N_485,N_122);
or U2529 (N_2529,N_796,N_624);
and U2530 (N_2530,N_539,N_2044);
xor U2531 (N_2531,N_449,N_2132);
or U2532 (N_2532,N_302,N_1657);
nand U2533 (N_2533,N_2383,N_917);
and U2534 (N_2534,N_1009,N_1602);
nand U2535 (N_2535,N_801,N_90);
xnor U2536 (N_2536,N_1772,N_984);
nand U2537 (N_2537,N_272,N_1329);
nor U2538 (N_2538,N_767,N_577);
or U2539 (N_2539,N_57,N_1996);
nand U2540 (N_2540,N_376,N_844);
or U2541 (N_2541,N_395,N_709);
or U2542 (N_2542,N_1295,N_2419);
nand U2543 (N_2543,N_15,N_2313);
xnor U2544 (N_2544,N_1210,N_986);
nand U2545 (N_2545,N_1010,N_1722);
nor U2546 (N_2546,N_2113,N_1040);
nand U2547 (N_2547,N_2292,N_2171);
and U2548 (N_2548,N_1696,N_924);
nand U2549 (N_2549,N_1516,N_1836);
and U2550 (N_2550,N_699,N_1114);
or U2551 (N_2551,N_2079,N_1249);
and U2552 (N_2552,N_322,N_453);
nand U2553 (N_2553,N_199,N_109);
nor U2554 (N_2554,N_1684,N_2413);
or U2555 (N_2555,N_1894,N_858);
nor U2556 (N_2556,N_1018,N_922);
nor U2557 (N_2557,N_295,N_935);
or U2558 (N_2558,N_2229,N_897);
nand U2559 (N_2559,N_953,N_2082);
nand U2560 (N_2560,N_415,N_870);
nor U2561 (N_2561,N_903,N_827);
xor U2562 (N_2562,N_2001,N_1011);
nand U2563 (N_2563,N_213,N_1096);
or U2564 (N_2564,N_311,N_1918);
and U2565 (N_2565,N_253,N_723);
or U2566 (N_2566,N_2017,N_2076);
nor U2567 (N_2567,N_1265,N_1335);
and U2568 (N_2568,N_197,N_2067);
and U2569 (N_2569,N_1239,N_245);
xnor U2570 (N_2570,N_1687,N_291);
or U2571 (N_2571,N_1640,N_1539);
or U2572 (N_2572,N_753,N_259);
and U2573 (N_2573,N_2069,N_1926);
xnor U2574 (N_2574,N_2386,N_2377);
and U2575 (N_2575,N_2471,N_541);
nand U2576 (N_2576,N_2042,N_2484);
or U2577 (N_2577,N_987,N_2299);
nand U2578 (N_2578,N_1446,N_419);
nand U2579 (N_2579,N_1321,N_1056);
nor U2580 (N_2580,N_1244,N_1846);
and U2581 (N_2581,N_713,N_694);
or U2582 (N_2582,N_800,N_1535);
nand U2583 (N_2583,N_312,N_2031);
xor U2584 (N_2584,N_394,N_1729);
or U2585 (N_2585,N_1266,N_1987);
and U2586 (N_2586,N_1596,N_2094);
nor U2587 (N_2587,N_1938,N_2370);
and U2588 (N_2588,N_848,N_1370);
nand U2589 (N_2589,N_467,N_1514);
nor U2590 (N_2590,N_1254,N_1315);
and U2591 (N_2591,N_379,N_487);
xnor U2592 (N_2592,N_640,N_1434);
and U2593 (N_2593,N_1225,N_719);
xnor U2594 (N_2594,N_1805,N_1155);
and U2595 (N_2595,N_7,N_1898);
nor U2596 (N_2596,N_2028,N_531);
and U2597 (N_2597,N_2208,N_1624);
nor U2598 (N_2598,N_910,N_1175);
nor U2599 (N_2599,N_1889,N_1544);
or U2600 (N_2600,N_1956,N_1402);
nand U2601 (N_2601,N_403,N_654);
nor U2602 (N_2602,N_770,N_1665);
xnor U2603 (N_2603,N_356,N_2092);
xnor U2604 (N_2604,N_318,N_167);
nand U2605 (N_2605,N_1866,N_1140);
nor U2606 (N_2606,N_0,N_147);
and U2607 (N_2607,N_1397,N_2124);
xor U2608 (N_2608,N_1332,N_2248);
and U2609 (N_2609,N_519,N_2116);
nand U2610 (N_2610,N_962,N_1737);
and U2611 (N_2611,N_1029,N_85);
xnor U2612 (N_2612,N_932,N_2478);
nand U2613 (N_2613,N_1769,N_1653);
xor U2614 (N_2614,N_875,N_120);
or U2615 (N_2615,N_2135,N_483);
nor U2616 (N_2616,N_1981,N_2454);
xnor U2617 (N_2617,N_2328,N_286);
and U2618 (N_2618,N_331,N_59);
or U2619 (N_2619,N_184,N_423);
nor U2620 (N_2620,N_856,N_1553);
or U2621 (N_2621,N_1631,N_546);
xor U2622 (N_2622,N_2397,N_1765);
nor U2623 (N_2623,N_86,N_2086);
nor U2624 (N_2624,N_111,N_2257);
nor U2625 (N_2625,N_1051,N_270);
and U2626 (N_2626,N_1026,N_1803);
or U2627 (N_2627,N_226,N_528);
or U2628 (N_2628,N_2101,N_592);
or U2629 (N_2629,N_1792,N_2360);
nor U2630 (N_2630,N_2331,N_1752);
and U2631 (N_2631,N_559,N_682);
xor U2632 (N_2632,N_387,N_24);
and U2633 (N_2633,N_879,N_507);
nor U2634 (N_2634,N_1773,N_390);
or U2635 (N_2635,N_157,N_2442);
nand U2636 (N_2636,N_533,N_2145);
or U2637 (N_2637,N_1555,N_202);
nor U2638 (N_2638,N_764,N_1787);
nand U2639 (N_2639,N_16,N_1727);
nor U2640 (N_2640,N_461,N_906);
xor U2641 (N_2641,N_1042,N_1581);
or U2642 (N_2642,N_1537,N_1969);
or U2643 (N_2643,N_717,N_1481);
nand U2644 (N_2644,N_2307,N_1670);
nand U2645 (N_2645,N_622,N_1261);
and U2646 (N_2646,N_1437,N_1549);
xnor U2647 (N_2647,N_2007,N_2203);
nor U2648 (N_2648,N_1991,N_243);
and U2649 (N_2649,N_396,N_29);
xnor U2650 (N_2650,N_1919,N_833);
nor U2651 (N_2651,N_159,N_681);
nor U2652 (N_2652,N_1608,N_1288);
nand U2653 (N_2653,N_2142,N_225);
xor U2654 (N_2654,N_136,N_365);
nor U2655 (N_2655,N_97,N_1320);
nand U2656 (N_2656,N_84,N_1185);
xnor U2657 (N_2657,N_363,N_1387);
xor U2658 (N_2658,N_1510,N_162);
xnor U2659 (N_2659,N_2433,N_738);
or U2660 (N_2660,N_484,N_1799);
nand U2661 (N_2661,N_781,N_860);
and U2662 (N_2662,N_2420,N_822);
and U2663 (N_2663,N_1348,N_328);
or U2664 (N_2664,N_1313,N_1234);
nor U2665 (N_2665,N_612,N_278);
nor U2666 (N_2666,N_2010,N_1188);
and U2667 (N_2667,N_1049,N_1691);
xor U2668 (N_2668,N_1391,N_446);
or U2669 (N_2669,N_1672,N_1468);
xor U2670 (N_2670,N_1063,N_762);
or U2671 (N_2671,N_1986,N_676);
xnor U2672 (N_2672,N_251,N_2108);
nor U2673 (N_2673,N_125,N_840);
nand U2674 (N_2674,N_1186,N_2078);
nor U2675 (N_2675,N_510,N_2220);
nand U2676 (N_2676,N_207,N_1933);
and U2677 (N_2677,N_1193,N_1911);
nand U2678 (N_2678,N_1551,N_273);
xor U2679 (N_2679,N_2279,N_1654);
or U2680 (N_2680,N_544,N_1366);
nor U2681 (N_2681,N_1078,N_1499);
xor U2682 (N_2682,N_1614,N_1780);
nand U2683 (N_2683,N_2295,N_536);
xor U2684 (N_2684,N_2430,N_916);
nor U2685 (N_2685,N_911,N_2194);
nand U2686 (N_2686,N_1506,N_634);
xnor U2687 (N_2687,N_530,N_422);
or U2688 (N_2688,N_1885,N_1381);
nor U2689 (N_2689,N_750,N_1872);
and U2690 (N_2690,N_1497,N_165);
nor U2691 (N_2691,N_2255,N_308);
xor U2692 (N_2692,N_2016,N_1813);
nand U2693 (N_2693,N_409,N_630);
or U2694 (N_2694,N_1572,N_1854);
nor U2695 (N_2695,N_2315,N_2384);
or U2696 (N_2696,N_1117,N_1401);
nand U2697 (N_2697,N_2106,N_1062);
nand U2698 (N_2698,N_1382,N_1970);
nand U2699 (N_2699,N_149,N_2320);
nor U2700 (N_2700,N_1954,N_2466);
nand U2701 (N_2701,N_1768,N_664);
xor U2702 (N_2702,N_1131,N_1831);
nand U2703 (N_2703,N_1992,N_2000);
xor U2704 (N_2704,N_1943,N_785);
nand U2705 (N_2705,N_2390,N_2446);
nand U2706 (N_2706,N_1388,N_1941);
and U2707 (N_2707,N_565,N_1130);
or U2708 (N_2708,N_594,N_2140);
nor U2709 (N_2709,N_1662,N_581);
or U2710 (N_2710,N_873,N_2278);
nor U2711 (N_2711,N_2364,N_2274);
and U2712 (N_2712,N_2335,N_1174);
and U2713 (N_2713,N_141,N_1467);
and U2714 (N_2714,N_320,N_1998);
nor U2715 (N_2715,N_1482,N_1441);
xor U2716 (N_2716,N_2321,N_1709);
or U2717 (N_2717,N_1036,N_1743);
and U2718 (N_2718,N_183,N_988);
nor U2719 (N_2719,N_1913,N_1909);
and U2720 (N_2720,N_2084,N_1564);
nor U2721 (N_2721,N_1203,N_760);
nand U2722 (N_2722,N_2114,N_580);
and U2723 (N_2723,N_1173,N_1766);
or U2724 (N_2724,N_1790,N_1022);
xor U2725 (N_2725,N_166,N_334);
and U2726 (N_2726,N_735,N_454);
or U2727 (N_2727,N_69,N_2136);
nand U2728 (N_2728,N_739,N_439);
or U2729 (N_2729,N_1604,N_337);
or U2730 (N_2730,N_521,N_1050);
xnor U2731 (N_2731,N_1949,N_443);
nor U2732 (N_2732,N_607,N_1304);
nor U2733 (N_2733,N_558,N_2048);
or U2734 (N_2734,N_1749,N_817);
nor U2735 (N_2735,N_786,N_1597);
nor U2736 (N_2736,N_151,N_2090);
or U2737 (N_2737,N_502,N_2176);
nor U2738 (N_2738,N_472,N_244);
and U2739 (N_2739,N_679,N_1069);
xor U2740 (N_2740,N_1995,N_2441);
nor U2741 (N_2741,N_2272,N_391);
nor U2742 (N_2742,N_2151,N_300);
nor U2743 (N_2743,N_1923,N_1420);
nand U2744 (N_2744,N_1110,N_269);
xor U2745 (N_2745,N_918,N_1303);
and U2746 (N_2746,N_1905,N_372);
or U2747 (N_2747,N_1912,N_677);
and U2748 (N_2748,N_1024,N_1679);
and U2749 (N_2749,N_1519,N_2421);
nor U2750 (N_2750,N_495,N_359);
or U2751 (N_2751,N_1751,N_36);
xor U2752 (N_2752,N_1668,N_1294);
nand U2753 (N_2753,N_1406,N_816);
nor U2754 (N_2754,N_881,N_447);
xor U2755 (N_2755,N_1385,N_437);
nand U2756 (N_2756,N_1637,N_2165);
nor U2757 (N_2757,N_382,N_2318);
or U2758 (N_2758,N_142,N_1159);
or U2759 (N_2759,N_1946,N_132);
or U2760 (N_2760,N_1044,N_515);
nor U2761 (N_2761,N_1617,N_1168);
xnor U2762 (N_2762,N_1522,N_23);
or U2763 (N_2763,N_1763,N_1047);
or U2764 (N_2764,N_2236,N_731);
nor U2765 (N_2765,N_1312,N_148);
nand U2766 (N_2766,N_143,N_2030);
nand U2767 (N_2767,N_2179,N_212);
or U2768 (N_2768,N_959,N_774);
nand U2769 (N_2769,N_2283,N_428);
nor U2770 (N_2770,N_799,N_1529);
nand U2771 (N_2771,N_620,N_1973);
xor U2772 (N_2772,N_1361,N_19);
nand U2773 (N_2773,N_1620,N_1444);
and U2774 (N_2774,N_1292,N_1480);
nor U2775 (N_2775,N_51,N_2180);
or U2776 (N_2776,N_145,N_1735);
xnor U2777 (N_2777,N_357,N_757);
nand U2778 (N_2778,N_1139,N_692);
xor U2779 (N_2779,N_1455,N_1652);
nor U2780 (N_2780,N_1744,N_48);
and U2781 (N_2781,N_909,N_2183);
or U2782 (N_2782,N_705,N_1494);
and U2783 (N_2783,N_246,N_205);
nand U2784 (N_2784,N_832,N_146);
or U2785 (N_2785,N_2493,N_1326);
and U2786 (N_2786,N_2399,N_1198);
xor U2787 (N_2787,N_2095,N_2459);
nor U2788 (N_2788,N_2359,N_2188);
and U2789 (N_2789,N_1934,N_610);
nand U2790 (N_2790,N_2439,N_1043);
nand U2791 (N_2791,N_1804,N_1196);
nor U2792 (N_2792,N_513,N_1486);
or U2793 (N_2793,N_2200,N_196);
xnor U2794 (N_2794,N_35,N_627);
xnor U2795 (N_2795,N_1068,N_586);
and U2796 (N_2796,N_1259,N_11);
and U2797 (N_2797,N_1490,N_2083);
nor U2798 (N_2798,N_2436,N_1694);
or U2799 (N_2799,N_1648,N_47);
nor U2800 (N_2800,N_633,N_2099);
or U2801 (N_2801,N_2468,N_693);
xnor U2802 (N_2802,N_283,N_1861);
nand U2803 (N_2803,N_882,N_758);
nand U2804 (N_2804,N_2411,N_53);
and U2805 (N_2805,N_591,N_1738);
xor U2806 (N_2806,N_964,N_1028);
and U2807 (N_2807,N_1690,N_890);
or U2808 (N_2808,N_2358,N_1342);
and U2809 (N_2809,N_298,N_2227);
xnor U2810 (N_2810,N_1376,N_1367);
or U2811 (N_2811,N_2449,N_787);
nand U2812 (N_2812,N_119,N_1534);
xnor U2813 (N_2813,N_740,N_2382);
nor U2814 (N_2814,N_672,N_1364);
xnor U2815 (N_2815,N_836,N_2087);
or U2816 (N_2816,N_1052,N_333);
and U2817 (N_2817,N_2038,N_1681);
nand U2818 (N_2818,N_1673,N_1758);
xor U2819 (N_2819,N_2221,N_2489);
nor U2820 (N_2820,N_1856,N_2309);
nor U2821 (N_2821,N_1160,N_1205);
nor U2822 (N_2822,N_1095,N_1711);
xnor U2823 (N_2823,N_2340,N_1310);
nor U2824 (N_2824,N_2102,N_771);
and U2825 (N_2825,N_1966,N_2029);
xor U2826 (N_2826,N_1742,N_2074);
or U2827 (N_2827,N_2275,N_730);
or U2828 (N_2828,N_72,N_863);
and U2829 (N_2829,N_229,N_724);
nor U2830 (N_2830,N_1255,N_1422);
and U2831 (N_2831,N_1726,N_1791);
and U2832 (N_2832,N_1398,N_2350);
xor U2833 (N_2833,N_1611,N_1427);
nor U2834 (N_2834,N_2476,N_1659);
nor U2835 (N_2835,N_1194,N_2117);
or U2836 (N_2836,N_660,N_1623);
or U2837 (N_2837,N_1983,N_330);
or U2838 (N_2838,N_1561,N_1890);
xor U2839 (N_2839,N_1524,N_1282);
and U2840 (N_2840,N_498,N_604);
nor U2841 (N_2841,N_56,N_1513);
or U2842 (N_2842,N_1085,N_2267);
or U2843 (N_2843,N_919,N_73);
nor U2844 (N_2844,N_1646,N_2302);
nand U2845 (N_2845,N_1045,N_354);
and U2846 (N_2846,N_1906,N_2496);
or U2847 (N_2847,N_1939,N_928);
nor U2848 (N_2848,N_1375,N_1932);
xor U2849 (N_2849,N_497,N_288);
or U2850 (N_2850,N_641,N_1599);
xor U2851 (N_2851,N_1407,N_179);
and U2852 (N_2852,N_1263,N_745);
or U2853 (N_2853,N_1048,N_1287);
and U2854 (N_2854,N_1087,N_1167);
nand U2855 (N_2855,N_71,N_941);
and U2856 (N_2856,N_1466,N_1746);
or U2857 (N_2857,N_1546,N_950);
or U2858 (N_2858,N_350,N_1323);
nand U2859 (N_2859,N_1324,N_2189);
and U2860 (N_2860,N_2034,N_1756);
nor U2861 (N_2861,N_1638,N_88);
and U2862 (N_2862,N_1750,N_908);
nand U2863 (N_2863,N_1788,N_1863);
and U2864 (N_2864,N_2282,N_233);
nor U2865 (N_2865,N_2043,N_80);
nand U2866 (N_2866,N_765,N_402);
or U2867 (N_2867,N_1945,N_869);
and U2868 (N_2868,N_1814,N_611);
and U2869 (N_2869,N_942,N_2064);
xor U2870 (N_2870,N_304,N_2210);
or U2871 (N_2871,N_2423,N_1908);
or U2872 (N_2872,N_405,N_1014);
xor U2873 (N_2873,N_242,N_279);
nor U2874 (N_2874,N_1097,N_407);
xnor U2875 (N_2875,N_386,N_728);
or U2876 (N_2876,N_63,N_1019);
or U2877 (N_2877,N_2298,N_54);
nand U2878 (N_2878,N_1178,N_2105);
or U2879 (N_2879,N_749,N_652);
nand U2880 (N_2880,N_1264,N_1182);
and U2881 (N_2881,N_1824,N_451);
or U2882 (N_2882,N_2089,N_1416);
nand U2883 (N_2883,N_2393,N_2365);
and U2884 (N_2884,N_1200,N_2431);
xor U2885 (N_2885,N_504,N_32);
and U2886 (N_2886,N_2418,N_1658);
and U2887 (N_2887,N_1171,N_20);
nand U2888 (N_2888,N_703,N_34);
nor U2889 (N_2889,N_271,N_1536);
nand U2890 (N_2890,N_946,N_401);
nand U2891 (N_2891,N_1666,N_2149);
and U2892 (N_2892,N_1412,N_2344);
and U2893 (N_2893,N_1118,N_1710);
nor U2894 (N_2894,N_1218,N_222);
or U2895 (N_2895,N_1410,N_27);
or U2896 (N_2896,N_1308,N_1394);
nor U2897 (N_2897,N_2241,N_1251);
or U2898 (N_2898,N_940,N_277);
xnor U2899 (N_2899,N_2058,N_1475);
nor U2900 (N_2900,N_1689,N_2260);
nor U2901 (N_2901,N_1578,N_2415);
nor U2902 (N_2902,N_680,N_232);
and U2903 (N_2903,N_1917,N_104);
nor U2904 (N_2904,N_2450,N_673);
xor U2905 (N_2905,N_562,N_175);
nand U2906 (N_2906,N_1635,N_163);
xnor U2907 (N_2907,N_543,N_127);
xor U2908 (N_2908,N_1584,N_2329);
nand U2909 (N_2909,N_2374,N_31);
nor U2910 (N_2910,N_2125,N_1020);
or U2911 (N_2911,N_1418,N_974);
and U2912 (N_2912,N_1123,N_10);
and U2913 (N_2913,N_2262,N_50);
xnor U2914 (N_2914,N_429,N_642);
or U2915 (N_2915,N_2300,N_789);
nor U2916 (N_2916,N_2404,N_378);
nor U2917 (N_2917,N_1834,N_33);
and U2918 (N_2918,N_1301,N_1760);
or U2919 (N_2919,N_2264,N_1296);
xnor U2920 (N_2920,N_2258,N_1120);
xnor U2921 (N_2921,N_1504,N_835);
nor U2922 (N_2922,N_306,N_1650);
nor U2923 (N_2923,N_715,N_1027);
and U2924 (N_2924,N_563,N_1115);
nor U2925 (N_2925,N_1518,N_2222);
nor U2926 (N_2926,N_1465,N_2405);
nand U2927 (N_2927,N_1899,N_2230);
and U2928 (N_2928,N_1074,N_1811);
xor U2929 (N_2929,N_1080,N_1840);
nor U2930 (N_2930,N_2205,N_2324);
or U2931 (N_2931,N_496,N_436);
nor U2932 (N_2932,N_79,N_1462);
xnor U2933 (N_2933,N_725,N_203);
and U2934 (N_2934,N_1794,N_1065);
nand U2935 (N_2935,N_667,N_1012);
and U2936 (N_2936,N_2080,N_2379);
nand U2937 (N_2937,N_1858,N_527);
nor U2938 (N_2938,N_1195,N_2035);
nor U2939 (N_2939,N_1793,N_1072);
or U2940 (N_2940,N_360,N_1930);
xnor U2941 (N_2941,N_2005,N_995);
nand U2942 (N_2942,N_1428,N_1165);
and U2943 (N_2943,N_284,N_914);
nor U2944 (N_2944,N_1461,N_182);
nor U2945 (N_2945,N_2052,N_2472);
nor U2946 (N_2946,N_169,N_107);
nor U2947 (N_2947,N_2167,N_638);
or U2948 (N_2948,N_2479,N_239);
or U2949 (N_2949,N_1344,N_1247);
and U2950 (N_2950,N_1897,N_1779);
nor U2951 (N_2951,N_1515,N_1474);
nand U2952 (N_2952,N_711,N_2243);
or U2953 (N_2953,N_2098,N_1390);
nor U2954 (N_2954,N_1651,N_2057);
or U2955 (N_2955,N_980,N_1431);
and U2956 (N_2956,N_458,N_1700);
xnor U2957 (N_2957,N_1354,N_158);
xnor U2958 (N_2958,N_688,N_1839);
and U2959 (N_2959,N_2212,N_1357);
nor U2960 (N_2960,N_1695,N_150);
nor U2961 (N_2961,N_416,N_6);
xor U2962 (N_2962,N_818,N_123);
nor U2963 (N_2963,N_1180,N_2311);
nor U2964 (N_2964,N_784,N_223);
and U2965 (N_2965,N_520,N_961);
nor U2966 (N_2966,N_1980,N_847);
nor U2967 (N_2967,N_658,N_1377);
and U2968 (N_2968,N_798,N_208);
xor U2969 (N_2969,N_1825,N_275);
and U2970 (N_2970,N_91,N_412);
or U2971 (N_2971,N_2215,N_550);
or U2972 (N_2972,N_2452,N_2334);
and U2973 (N_2973,N_1976,N_904);
or U2974 (N_2974,N_1920,N_2066);
nand U2975 (N_2975,N_1977,N_1770);
nor U2976 (N_2976,N_266,N_1092);
or U2977 (N_2977,N_761,N_1565);
and U2978 (N_2978,N_1338,N_1360);
nor U2979 (N_2979,N_662,N_281);
xor U2980 (N_2980,N_138,N_368);
nor U2981 (N_2981,N_2326,N_1902);
or U2982 (N_2982,N_2163,N_1447);
or U2983 (N_2983,N_2234,N_1176);
or U2984 (N_2984,N_1339,N_128);
nand U2985 (N_2985,N_1086,N_1242);
nor U2986 (N_2986,N_893,N_1419);
or U2987 (N_2987,N_297,N_1273);
or U2988 (N_2988,N_2182,N_476);
nor U2989 (N_2989,N_1699,N_716);
and U2990 (N_2990,N_1707,N_1240);
or U2991 (N_2991,N_1669,N_2191);
nand U2992 (N_2992,N_1712,N_2143);
and U2993 (N_2993,N_305,N_2438);
and U2994 (N_2994,N_545,N_2025);
nor U2995 (N_2995,N_975,N_1843);
nor U2996 (N_2996,N_1199,N_583);
xor U2997 (N_2997,N_2103,N_1560);
and U2998 (N_2998,N_256,N_1521);
nor U2999 (N_2999,N_663,N_1606);
nor U3000 (N_3000,N_89,N_853);
nor U3001 (N_3001,N_2457,N_2198);
or U3002 (N_3002,N_564,N_2138);
or U3003 (N_3003,N_1107,N_377);
or U3004 (N_3004,N_712,N_1774);
nor U3005 (N_3005,N_1503,N_1297);
nand U3006 (N_3006,N_871,N_82);
nor U3007 (N_3007,N_990,N_17);
nand U3008 (N_3008,N_1319,N_2062);
or U3009 (N_3009,N_2408,N_1104);
xor U3010 (N_3010,N_597,N_155);
and U3011 (N_3011,N_2297,N_532);
and U3012 (N_3012,N_2172,N_907);
nand U3013 (N_3013,N_1172,N_1731);
xor U3014 (N_3014,N_413,N_1879);
nand U3015 (N_3015,N_76,N_1099);
nand U3016 (N_3016,N_2263,N_1484);
or U3017 (N_3017,N_224,N_2410);
xnor U3018 (N_3018,N_1383,N_737);
nand U3019 (N_3019,N_1125,N_201);
and U3020 (N_3020,N_626,N_2376);
xor U3021 (N_3021,N_2181,N_579);
or U3022 (N_3022,N_152,N_2199);
nor U3023 (N_3023,N_2231,N_1088);
or U3024 (N_3024,N_810,N_335);
and U3025 (N_3025,N_1046,N_1238);
or U3026 (N_3026,N_1579,N_655);
xnor U3027 (N_3027,N_803,N_2495);
xor U3028 (N_3028,N_478,N_262);
and U3029 (N_3029,N_978,N_287);
nand U3030 (N_3030,N_2281,N_1371);
nor U3031 (N_3031,N_2285,N_2333);
and U3032 (N_3032,N_1346,N_1676);
xnor U3033 (N_3033,N_280,N_1368);
or U3034 (N_3034,N_1119,N_825);
nand U3035 (N_3035,N_1157,N_1001);
and U3036 (N_3036,N_351,N_629);
or U3037 (N_3037,N_1291,N_570);
and U3038 (N_3038,N_28,N_948);
nor U3039 (N_3039,N_252,N_1111);
nand U3040 (N_3040,N_1716,N_1055);
and U3041 (N_3041,N_135,N_631);
and U3042 (N_3042,N_2266,N_2127);
xnor U3043 (N_3043,N_1910,N_866);
and U3044 (N_3044,N_96,N_465);
xor U3045 (N_3045,N_2091,N_3);
xnor U3046 (N_3046,N_2371,N_1972);
nand U3047 (N_3047,N_1821,N_915);
or U3048 (N_3048,N_2417,N_2341);
nand U3049 (N_3049,N_1962,N_1789);
nand U3050 (N_3050,N_1083,N_2259);
xnor U3051 (N_3051,N_886,N_1267);
nand U3052 (N_3052,N_77,N_1639);
or U3053 (N_3053,N_1587,N_81);
and U3054 (N_3054,N_1122,N_1845);
or U3055 (N_3055,N_913,N_285);
and U3056 (N_3056,N_2435,N_795);
nor U3057 (N_3057,N_734,N_1656);
and U3058 (N_3058,N_95,N_2032);
and U3059 (N_3059,N_1891,N_1285);
nor U3060 (N_3060,N_1706,N_1206);
and U3061 (N_3061,N_381,N_1243);
nand U3062 (N_3062,N_1632,N_977);
xnor U3063 (N_3063,N_1823,N_1215);
nand U3064 (N_3064,N_555,N_993);
nand U3065 (N_3065,N_837,N_1307);
or U3066 (N_3066,N_1526,N_2235);
nand U3067 (N_3067,N_1450,N_296);
xnor U3068 (N_3068,N_574,N_1595);
or U3069 (N_3069,N_1132,N_2173);
or U3070 (N_3070,N_1870,N_380);
and U3071 (N_3071,N_659,N_1904);
or U3072 (N_3072,N_831,N_889);
xnor U3073 (N_3073,N_503,N_1302);
and U3074 (N_3074,N_600,N_1438);
xor U3075 (N_3075,N_1571,N_40);
xor U3076 (N_3076,N_1903,N_2407);
and U3077 (N_3077,N_1143,N_1984);
nor U3078 (N_3078,N_1502,N_1947);
nor U3079 (N_3079,N_2289,N_1877);
xnor U3080 (N_3080,N_931,N_790);
and U3081 (N_3081,N_1137,N_1717);
xnor U3082 (N_3082,N_773,N_1305);
nor U3083 (N_3083,N_174,N_783);
or U3084 (N_3084,N_1720,N_1950);
nor U3085 (N_3085,N_2369,N_1968);
or U3086 (N_3086,N_2050,N_1181);
and U3087 (N_3087,N_1795,N_2487);
and U3088 (N_3088,N_464,N_2387);
or U3089 (N_3089,N_824,N_951);
xnor U3090 (N_3090,N_1322,N_2458);
xor U3091 (N_3091,N_121,N_1728);
nand U3092 (N_3092,N_1975,N_1600);
or U3093 (N_3093,N_87,N_1718);
or U3094 (N_3094,N_1098,N_1016);
or U3095 (N_3095,N_1257,N_2332);
nor U3096 (N_3096,N_1289,N_1369);
nand U3097 (N_3097,N_905,N_1349);
nand U3098 (N_3098,N_133,N_1358);
nand U3099 (N_3099,N_1776,N_1921);
and U3100 (N_3100,N_1064,N_2046);
nand U3101 (N_3101,N_900,N_839);
and U3102 (N_3102,N_1272,N_2239);
nor U3103 (N_3103,N_254,N_240);
and U3104 (N_3104,N_685,N_294);
nand U3105 (N_3105,N_1594,N_1822);
xnor U3106 (N_3106,N_991,N_1054);
nand U3107 (N_3107,N_60,N_399);
nand U3108 (N_3108,N_1232,N_1686);
and U3109 (N_3109,N_2395,N_804);
xor U3110 (N_3110,N_1443,N_2244);
or U3111 (N_3111,N_2460,N_1211);
and U3112 (N_3112,N_1871,N_237);
or U3113 (N_3113,N_2107,N_1878);
and U3114 (N_3114,N_326,N_452);
nand U3115 (N_3115,N_267,N_92);
and U3116 (N_3116,N_1100,N_2277);
xnor U3117 (N_3117,N_1757,N_1489);
nand U3118 (N_3118,N_1641,N_2440);
nor U3119 (N_3119,N_516,N_336);
nor U3120 (N_3120,N_584,N_921);
nand U3121 (N_3121,N_2185,N_2023);
xnor U3122 (N_3122,N_1008,N_2119);
and U3123 (N_3123,N_1838,N_511);
or U3124 (N_3124,N_1771,N_1830);
or U3125 (N_3125,N_1299,N_1655);
nand U3126 (N_3126,N_61,N_2347);
nor U3127 (N_3127,N_2049,N_623);
xor U3128 (N_3128,N_1963,N_2403);
or U3129 (N_3129,N_362,N_2070);
and U3130 (N_3130,N_707,N_2228);
nor U3131 (N_3131,N_1135,N_553);
or U3132 (N_3132,N_896,N_1187);
nand U3133 (N_3133,N_52,N_1059);
nor U3134 (N_3134,N_231,N_883);
nand U3135 (N_3135,N_1231,N_1586);
nor U3136 (N_3136,N_1477,N_2271);
nand U3137 (N_3137,N_1618,N_744);
nand U3138 (N_3138,N_2224,N_115);
nand U3139 (N_3139,N_139,N_571);
nand U3140 (N_3140,N_2314,N_561);
nor U3141 (N_3141,N_1463,N_2490);
nand U3142 (N_3142,N_1558,N_420);
and U3143 (N_3143,N_1929,N_265);
nand U3144 (N_3144,N_2045,N_1030);
nor U3145 (N_3145,N_101,N_1309);
nand U3146 (N_3146,N_18,N_639);
nor U3147 (N_3147,N_2317,N_1914);
or U3148 (N_3148,N_2322,N_1129);
or U3149 (N_3149,N_2485,N_217);
and U3150 (N_3150,N_1424,N_2319);
or U3151 (N_3151,N_648,N_49);
nor U3152 (N_3152,N_313,N_117);
and U3153 (N_3153,N_859,N_105);
or U3154 (N_3154,N_2465,N_1076);
nand U3155 (N_3155,N_392,N_898);
nand U3156 (N_3156,N_367,N_752);
and U3157 (N_3157,N_834,N_1311);
and U3158 (N_3158,N_2093,N_1985);
nand U3159 (N_3159,N_1415,N_2150);
and U3160 (N_3160,N_1868,N_164);
nor U3161 (N_3161,N_2131,N_2186);
or U3162 (N_3162,N_998,N_1867);
xnor U3163 (N_3163,N_481,N_1031);
or U3164 (N_3164,N_621,N_970);
and U3165 (N_3165,N_2428,N_608);
xnor U3166 (N_3166,N_657,N_2473);
xnor U3167 (N_3167,N_1456,N_2367);
nor U3168 (N_3168,N_292,N_1873);
and U3169 (N_3169,N_2156,N_1645);
xor U3170 (N_3170,N_2021,N_967);
nor U3171 (N_3171,N_2327,N_2217);
nand U3172 (N_3172,N_1248,N_972);
nor U3173 (N_3173,N_780,N_746);
or U3174 (N_3174,N_66,N_2346);
or U3175 (N_3175,N_456,N_156);
or U3176 (N_3176,N_1671,N_2422);
xor U3177 (N_3177,N_1343,N_849);
xnor U3178 (N_3178,N_1767,N_1246);
xnor U3179 (N_3179,N_819,N_1552);
nor U3180 (N_3180,N_714,N_1708);
or U3181 (N_3181,N_846,N_989);
xnor U3182 (N_3182,N_878,N_2184);
and U3183 (N_3183,N_2424,N_1812);
nand U3184 (N_3184,N_1142,N_727);
or U3185 (N_3185,N_2022,N_2161);
and U3186 (N_3186,N_1621,N_2197);
and U3187 (N_3187,N_2343,N_2024);
and U3188 (N_3188,N_1826,N_1547);
nand U3189 (N_3189,N_1622,N_671);
nor U3190 (N_3190,N_1960,N_114);
xor U3191 (N_3191,N_2388,N_1961);
nand U3192 (N_3192,N_2475,N_1061);
xnor U3193 (N_3193,N_2443,N_1566);
nor U3194 (N_3194,N_2096,N_751);
nor U3195 (N_3195,N_768,N_4);
and U3196 (N_3196,N_383,N_857);
nor U3197 (N_3197,N_1778,N_1959);
xnor U3198 (N_3198,N_340,N_364);
nor U3199 (N_3199,N_569,N_2306);
nor U3200 (N_3200,N_43,N_1892);
nand U3201 (N_3201,N_83,N_1148);
and U3202 (N_3202,N_2133,N_2392);
or U3203 (N_3203,N_1883,N_316);
xnor U3204 (N_3204,N_2463,N_1619);
xnor U3205 (N_3205,N_1893,N_289);
or U3206 (N_3206,N_488,N_1372);
xor U3207 (N_3207,N_1164,N_1278);
xor U3208 (N_3208,N_181,N_1634);
or U3209 (N_3209,N_1875,N_341);
or U3210 (N_3210,N_1071,N_408);
or U3211 (N_3211,N_2448,N_418);
nand U3212 (N_3212,N_1833,N_1340);
and U3213 (N_3213,N_171,N_2254);
xnor U3214 (N_3214,N_249,N_1347);
and U3215 (N_3215,N_2111,N_2118);
xor U3216 (N_3216,N_1520,N_1379);
xor U3217 (N_3217,N_344,N_1041);
nor U3218 (N_3218,N_1126,N_1191);
or U3219 (N_3219,N_1352,N_2462);
nor U3220 (N_3220,N_1409,N_1154);
or U3221 (N_3221,N_2253,N_178);
xor U3222 (N_3222,N_2206,N_1698);
xor U3223 (N_3223,N_1527,N_1224);
and U3224 (N_3224,N_1213,N_2303);
nor U3225 (N_3225,N_276,N_1819);
nand U3226 (N_3226,N_960,N_301);
xor U3227 (N_3227,N_2152,N_1577);
or U3228 (N_3228,N_2071,N_1820);
nand U3229 (N_3229,N_1882,N_1556);
and U3230 (N_3230,N_872,N_2391);
nand U3231 (N_3231,N_732,N_1219);
or U3232 (N_3232,N_299,N_1660);
or U3233 (N_3233,N_2480,N_741);
nor U3234 (N_3234,N_426,N_777);
xnor U3235 (N_3235,N_2494,N_1633);
or U3236 (N_3236,N_899,N_1940);
xnor U3237 (N_3237,N_2469,N_1032);
nand U3238 (N_3238,N_968,N_1505);
nand U3239 (N_3239,N_1314,N_339);
and U3240 (N_3240,N_1417,N_1538);
or U3241 (N_3241,N_490,N_1517);
nand U3242 (N_3242,N_2169,N_599);
nand U3243 (N_3243,N_191,N_41);
or U3244 (N_3244,N_925,N_1928);
nor U3245 (N_3245,N_2196,N_678);
xor U3246 (N_3246,N_593,N_2363);
nand U3247 (N_3247,N_255,N_1179);
nor U3248 (N_3248,N_25,N_1680);
and U3249 (N_3249,N_13,N_424);
xor U3250 (N_3250,N_1724,N_459);
and U3251 (N_3251,N_1719,N_1039);
or U3252 (N_3252,N_567,N_1937);
or U3253 (N_3253,N_865,N_1333);
xnor U3254 (N_3254,N_2416,N_1378);
and U3255 (N_3255,N_1967,N_971);
nor U3256 (N_3256,N_176,N_1341);
xor U3257 (N_3257,N_1924,N_352);
xor U3258 (N_3258,N_1105,N_772);
xor U3259 (N_3259,N_651,N_369);
nand U3260 (N_3260,N_901,N_1276);
nand U3261 (N_3261,N_384,N_1274);
xnor U3262 (N_3262,N_1807,N_802);
xnor U3263 (N_3263,N_523,N_2357);
nor U3264 (N_3264,N_1576,N_1161);
or U3265 (N_3265,N_462,N_329);
and U3266 (N_3266,N_1554,N_548);
or U3267 (N_3267,N_877,N_1134);
nand U3268 (N_3268,N_1440,N_706);
nor U3269 (N_3269,N_2486,N_2325);
nor U3270 (N_3270,N_1077,N_1759);
nor U3271 (N_3271,N_1753,N_1647);
nand U3272 (N_3272,N_1978,N_547);
nor U3273 (N_3273,N_1153,N_64);
nor U3274 (N_3274,N_1237,N_404);
nand U3275 (N_3275,N_1850,N_2120);
xor U3276 (N_3276,N_1569,N_241);
nor U3277 (N_3277,N_62,N_1084);
xor U3278 (N_3278,N_1745,N_665);
or U3279 (N_3279,N_1488,N_2204);
or U3280 (N_3280,N_137,N_718);
nand U3281 (N_3281,N_1589,N_596);
nand U3282 (N_3282,N_894,N_1330);
and U3283 (N_3283,N_1715,N_1331);
xor U3284 (N_3284,N_1403,N_656);
nor U3285 (N_3285,N_1345,N_108);
and U3286 (N_3286,N_1636,N_1853);
nor U3287 (N_3287,N_862,N_2245);
or U3288 (N_3288,N_1013,N_2409);
nand U3289 (N_3289,N_1423,N_806);
or U3290 (N_3290,N_67,N_216);
xor U3291 (N_3291,N_1796,N_1433);
nor U3292 (N_3292,N_1034,N_2178);
and U3293 (N_3293,N_371,N_1138);
xnor U3294 (N_3294,N_1075,N_131);
nor U3295 (N_3295,N_410,N_590);
xnor U3296 (N_3296,N_75,N_2276);
or U3297 (N_3297,N_976,N_2225);
or U3298 (N_3298,N_1038,N_2051);
and U3299 (N_3299,N_2240,N_68);
and U3300 (N_3300,N_1365,N_852);
and U3301 (N_3301,N_1989,N_1663);
nor U3302 (N_3302,N_2033,N_1800);
and U3303 (N_3303,N_1809,N_1886);
or U3304 (N_3304,N_766,N_1693);
nand U3305 (N_3305,N_116,N_2251);
or U3306 (N_3306,N_1740,N_1979);
xnor U3307 (N_3307,N_1208,N_1350);
and U3308 (N_3308,N_26,N_319);
nor U3309 (N_3309,N_1942,N_864);
xor U3310 (N_3310,N_1221,N_1837);
nand U3311 (N_3311,N_1844,N_2444);
xor U3312 (N_3312,N_421,N_126);
nand U3313 (N_3313,N_2159,N_2130);
nand U3314 (N_3314,N_637,N_2211);
nand U3315 (N_3315,N_1133,N_1005);
nand U3316 (N_3316,N_1101,N_2014);
nor U3317 (N_3317,N_30,N_1067);
nand U3318 (N_3318,N_2366,N_1733);
nand U3319 (N_3319,N_1927,N_1944);
or U3320 (N_3320,N_669,N_100);
xnor U3321 (N_3321,N_2432,N_448);
xnor U3322 (N_3322,N_470,N_1207);
nor U3323 (N_3323,N_1649,N_2004);
nor U3324 (N_3324,N_2214,N_982);
or U3325 (N_3325,N_686,N_1607);
xnor U3326 (N_3326,N_2308,N_45);
xnor U3327 (N_3327,N_2470,N_549);
nor U3328 (N_3328,N_963,N_1583);
nand U3329 (N_3329,N_1449,N_185);
nor U3330 (N_3330,N_460,N_2218);
nor U3331 (N_3331,N_1201,N_1815);
nand U3332 (N_3332,N_792,N_2400);
nor U3333 (N_3333,N_1730,N_2112);
and U3334 (N_3334,N_1306,N_2003);
and U3335 (N_3335,N_500,N_2414);
and U3336 (N_3336,N_1493,N_605);
nand U3337 (N_3337,N_1786,N_1204);
and U3338 (N_3338,N_1952,N_1058);
and U3339 (N_3339,N_361,N_2055);
or U3340 (N_3340,N_811,N_813);
or U3341 (N_3341,N_1675,N_2269);
nand U3342 (N_3342,N_1540,N_884);
nand U3343 (N_3343,N_1835,N_230);
and U3344 (N_3344,N_1542,N_506);
xnor U3345 (N_3345,N_1082,N_1430);
and U3346 (N_3346,N_645,N_1253);
nor U3347 (N_3347,N_1592,N_829);
and U3348 (N_3348,N_2337,N_1396);
nor U3349 (N_3349,N_160,N_2190);
and U3350 (N_3350,N_965,N_701);
xnor U3351 (N_3351,N_957,N_1714);
xor U3352 (N_3352,N_708,N_1334);
and U3353 (N_3353,N_442,N_1762);
and U3354 (N_3354,N_512,N_891);
or U3355 (N_3355,N_635,N_260);
nand U3356 (N_3356,N_1721,N_575);
and U3357 (N_3357,N_981,N_1070);
nor U3358 (N_3358,N_1500,N_2498);
and U3359 (N_3359,N_168,N_850);
or U3360 (N_3360,N_1318,N_743);
nand U3361 (N_3361,N_1245,N_1217);
and U3362 (N_3362,N_1852,N_1881);
nor U3363 (N_3363,N_2467,N_324);
nand U3364 (N_3364,N_140,N_2237);
nor U3365 (N_3365,N_1550,N_888);
nor U3366 (N_3366,N_509,N_2026);
nor U3367 (N_3367,N_1121,N_2287);
xor U3368 (N_3368,N_2141,N_2013);
nor U3369 (N_3369,N_2039,N_325);
and U3370 (N_3370,N_2073,N_353);
and U3371 (N_3371,N_1476,N_556);
nand U3372 (N_3372,N_2310,N_1775);
nor U3373 (N_3373,N_366,N_1990);
and U3374 (N_3374,N_38,N_812);
and U3375 (N_3375,N_1452,N_2437);
nand U3376 (N_3376,N_228,N_1573);
and U3377 (N_3377,N_93,N_1563);
or U3378 (N_3378,N_992,N_938);
nand U3379 (N_3379,N_1832,N_1588);
or U3380 (N_3380,N_2488,N_1901);
nand U3381 (N_3381,N_2193,N_1151);
or U3382 (N_3382,N_1209,N_1150);
nor U3383 (N_3383,N_235,N_1971);
nor U3384 (N_3384,N_349,N_1270);
and U3385 (N_3385,N_1739,N_742);
nand U3386 (N_3386,N_2061,N_1806);
nor U3387 (N_3387,N_9,N_1864);
or U3388 (N_3388,N_1235,N_2213);
nor U3389 (N_3389,N_1532,N_1141);
xnor U3390 (N_3390,N_1701,N_668);
or U3391 (N_3391,N_2246,N_566);
or U3392 (N_3392,N_2195,N_2097);
nor U3393 (N_3393,N_1228,N_601);
nor U3394 (N_3394,N_1575,N_134);
and U3395 (N_3395,N_200,N_1400);
or U3396 (N_3396,N_188,N_1582);
and U3397 (N_3397,N_841,N_1828);
and U3398 (N_3398,N_153,N_1703);
or U3399 (N_3399,N_1158,N_2280);
nor U3400 (N_3400,N_710,N_463);
and U3401 (N_3401,N_1688,N_809);
and U3402 (N_3402,N_1781,N_1256);
xor U3403 (N_3403,N_1764,N_2110);
or U3404 (N_3404,N_1674,N_2294);
nand U3405 (N_3405,N_2170,N_417);
and U3406 (N_3406,N_431,N_1678);
or U3407 (N_3407,N_1713,N_2261);
and U3408 (N_3408,N_1585,N_321);
xnor U3409 (N_3409,N_2284,N_39);
or U3410 (N_3410,N_2242,N_912);
xor U3411 (N_3411,N_616,N_775);
and U3412 (N_3412,N_1874,N_2247);
and U3413 (N_3413,N_609,N_997);
xor U3414 (N_3414,N_1091,N_695);
nand U3415 (N_3415,N_186,N_1362);
xor U3416 (N_3416,N_343,N_1848);
nand U3417 (N_3417,N_2301,N_1353);
nand U3418 (N_3418,N_754,N_1216);
nor U3419 (N_3419,N_814,N_2268);
or U3420 (N_3420,N_1214,N_1953);
nand U3421 (N_3421,N_939,N_112);
xor U3422 (N_3422,N_687,N_323);
and U3423 (N_3423,N_1784,N_1487);
xnor U3424 (N_3424,N_1483,N_1328);
nor U3425 (N_3425,N_797,N_310);
nor U3426 (N_3426,N_2075,N_625);
or U3427 (N_3427,N_398,N_2296);
or U3428 (N_3428,N_845,N_966);
nor U3429 (N_3429,N_263,N_2085);
nor U3430 (N_3430,N_1591,N_1439);
and U3431 (N_3431,N_1895,N_1988);
xor U3432 (N_3432,N_1202,N_902);
or U3433 (N_3433,N_1736,N_1492);
nor U3434 (N_3434,N_1829,N_930);
and U3435 (N_3435,N_885,N_2305);
or U3436 (N_3436,N_952,N_315);
xor U3437 (N_3437,N_499,N_1593);
and U3438 (N_3438,N_1460,N_1629);
or U3439 (N_3439,N_282,N_1545);
nand U3440 (N_3440,N_736,N_2019);
xor U3441 (N_3441,N_1997,N_2155);
nor U3442 (N_3442,N_1808,N_1915);
nand U3443 (N_3443,N_1568,N_1432);
xor U3444 (N_3444,N_189,N_1233);
and U3445 (N_3445,N_2158,N_411);
or U3446 (N_3446,N_1448,N_348);
nor U3447 (N_3447,N_2,N_475);
and U3448 (N_3448,N_374,N_1496);
nor U3449 (N_3449,N_1184,N_2015);
or U3450 (N_3450,N_861,N_1625);
nor U3451 (N_3451,N_2396,N_144);
xnor U3452 (N_3452,N_1798,N_1404);
nand U3453 (N_3453,N_110,N_1269);
nor U3454 (N_3454,N_2373,N_2312);
xnor U3455 (N_3455,N_1197,N_1955);
and U3456 (N_3456,N_1017,N_1037);
nand U3457 (N_3457,N_923,N_1112);
nor U3458 (N_3458,N_598,N_1327);
nand U3459 (N_3459,N_2349,N_195);
nand U3460 (N_3460,N_830,N_450);
and U3461 (N_3461,N_747,N_2427);
nor U3462 (N_3462,N_1442,N_776);
nand U3463 (N_3463,N_2447,N_1057);
nor U3464 (N_3464,N_2216,N_1993);
nand U3465 (N_3465,N_2394,N_650);
nor U3466 (N_3466,N_1958,N_327);
or U3467 (N_3467,N_535,N_2425);
nor U3468 (N_3468,N_2233,N_945);
and U3469 (N_3469,N_220,N_1325);
xnor U3470 (N_3470,N_720,N_956);
or U3471 (N_3471,N_2381,N_1994);
xnor U3472 (N_3472,N_2372,N_514);
nand U3473 (N_3473,N_2041,N_1359);
xor U3474 (N_3474,N_2226,N_1683);
xor U3475 (N_3475,N_1106,N_1236);
nand U3476 (N_3476,N_2219,N_1907);
nor U3477 (N_3477,N_58,N_274);
xor U3478 (N_3478,N_303,N_479);
and U3479 (N_3479,N_763,N_1900);
and U3480 (N_3480,N_2461,N_489);
and U3481 (N_3481,N_1399,N_851);
or U3482 (N_3482,N_823,N_268);
xor U3483 (N_3483,N_209,N_636);
and U3484 (N_3484,N_1512,N_1393);
and U3485 (N_3485,N_1754,N_927);
and U3486 (N_3486,N_2353,N_1644);
nor U3487 (N_3487,N_194,N_1896);
and U3488 (N_3488,N_1590,N_526);
and U3489 (N_3489,N_1337,N_370);
nor U3490 (N_3490,N_1931,N_1275);
nand U3491 (N_3491,N_494,N_2072);
or U3492 (N_3492,N_698,N_1102);
xor U3493 (N_3493,N_37,N_1498);
or U3494 (N_3494,N_2068,N_1280);
nand U3495 (N_3495,N_2291,N_258);
xnor U3496 (N_3496,N_468,N_1170);
xnor U3497 (N_3497,N_700,N_1144);
nand U3498 (N_3498,N_2201,N_1374);
or U3499 (N_3499,N_2037,N_538);
nor U3500 (N_3500,N_1093,N_1562);
xor U3501 (N_3501,N_480,N_1777);
nor U3502 (N_3502,N_1531,N_778);
nand U3503 (N_3503,N_1965,N_177);
xor U3504 (N_3504,N_1286,N_880);
nand U3505 (N_3505,N_1661,N_2474);
nor U3506 (N_3506,N_2354,N_578);
xor U3507 (N_3507,N_1000,N_1869);
and U3508 (N_3508,N_855,N_508);
and U3509 (N_3509,N_293,N_2273);
and U3510 (N_3510,N_1974,N_1007);
or U3511 (N_3511,N_1865,N_949);
nor U3512 (N_3512,N_572,N_1459);
xnor U3513 (N_3513,N_643,N_2012);
nand U3514 (N_3514,N_486,N_1705);
nand U3515 (N_3515,N_2238,N_1612);
and U3516 (N_3516,N_2401,N_1841);
and U3517 (N_3517,N_1643,N_1277);
or U3518 (N_3518,N_748,N_44);
and U3519 (N_3519,N_393,N_1473);
nand U3520 (N_3520,N_455,N_2160);
nand U3521 (N_3521,N_755,N_1847);
and U3522 (N_3522,N_2356,N_22);
or U3523 (N_3523,N_264,N_2088);
nor U3524 (N_3524,N_215,N_1177);
and U3525 (N_3525,N_2109,N_568);
or U3526 (N_3526,N_2139,N_2157);
xnor U3527 (N_3527,N_389,N_1279);
nand U3528 (N_3528,N_1002,N_585);
or U3529 (N_3529,N_603,N_1220);
nor U3530 (N_3530,N_2464,N_876);
nand U3531 (N_3531,N_2348,N_2122);
xor U3532 (N_3532,N_2175,N_1810);
nand U3533 (N_3533,N_534,N_2174);
or U3534 (N_3534,N_469,N_2483);
and U3535 (N_3535,N_2177,N_219);
xor U3536 (N_3536,N_1827,N_1025);
xnor U3537 (N_3537,N_342,N_248);
nand U3538 (N_3538,N_936,N_619);
and U3539 (N_3539,N_2256,N_1156);
nor U3540 (N_3540,N_1936,N_2445);
nand U3541 (N_3541,N_1284,N_1147);
xnor U3542 (N_3542,N_113,N_1702);
nand U3543 (N_3543,N_1015,N_2100);
and U3544 (N_3544,N_355,N_1627);
nor U3545 (N_3545,N_2355,N_505);
xnor U3546 (N_3546,N_704,N_1925);
and U3547 (N_3547,N_55,N_12);
and U3548 (N_3548,N_1509,N_1136);
or U3549 (N_3549,N_867,N_926);
nor U3550 (N_3550,N_1580,N_1094);
nor U3551 (N_3551,N_2368,N_42);
or U3552 (N_3552,N_1356,N_1818);
and U3553 (N_3553,N_1857,N_2290);
nor U3554 (N_3554,N_1293,N_1704);
xor U3555 (N_3555,N_791,N_2065);
or U3556 (N_3556,N_21,N_2123);
xor U3557 (N_3557,N_2252,N_2412);
xor U3558 (N_3558,N_445,N_332);
and U3559 (N_3559,N_103,N_1501);
xor U3560 (N_3560,N_807,N_440);
or U3561 (N_3561,N_187,N_613);
nor U3562 (N_3562,N_2168,N_1922);
or U3563 (N_3563,N_1855,N_2147);
xnor U3564 (N_3564,N_1222,N_2166);
nor U3565 (N_3565,N_1081,N_2380);
or U3566 (N_3566,N_2134,N_1523);
nor U3567 (N_3567,N_958,N_1336);
xor U3568 (N_3568,N_1692,N_441);
nand U3569 (N_3569,N_1411,N_1271);
and U3570 (N_3570,N_696,N_493);
and U3571 (N_3571,N_1,N_874);
nor U3572 (N_3572,N_1317,N_1227);
or U3573 (N_3573,N_1816,N_1478);
and U3574 (N_3574,N_388,N_573);
nor U3575 (N_3575,N_689,N_1862);
and U3576 (N_3576,N_854,N_759);
nor U3577 (N_3577,N_617,N_347);
or U3578 (N_3578,N_929,N_1351);
and U3579 (N_3579,N_821,N_1103);
nor U3580 (N_3580,N_1023,N_198);
and U3581 (N_3581,N_1851,N_1006);
nor U3582 (N_3582,N_646,N_653);
nand U3583 (N_3583,N_587,N_1888);
xnor U3584 (N_3584,N_192,N_2385);
nor U3585 (N_3585,N_1252,N_1021);
xnor U3586 (N_3586,N_2316,N_722);
or U3587 (N_3587,N_1421,N_1212);
and U3588 (N_3588,N_190,N_1108);
xnor U3589 (N_3589,N_346,N_74);
and U3590 (N_3590,N_1603,N_2453);
and U3591 (N_3591,N_947,N_2146);
nor U3592 (N_3592,N_1472,N_582);
xnor U3593 (N_3593,N_557,N_1485);
and U3594 (N_3594,N_425,N_2286);
and U3595 (N_3595,N_1723,N_1260);
xnor U3596 (N_3596,N_1363,N_2137);
and U3597 (N_3597,N_1559,N_2429);
nand U3598 (N_3598,N_2223,N_1250);
nand U3599 (N_3599,N_1435,N_1283);
and U3600 (N_3600,N_2192,N_2009);
and U3601 (N_3601,N_1697,N_943);
nand U3602 (N_3602,N_427,N_1183);
xor U3603 (N_3603,N_2434,N_2121);
nor U3604 (N_3604,N_2104,N_969);
nor U3605 (N_3605,N_733,N_979);
nor U3606 (N_3606,N_1880,N_1642);
nand U3607 (N_3607,N_1884,N_2063);
xor U3608 (N_3608,N_2336,N_1741);
nand U3609 (N_3609,N_1066,N_1429);
and U3610 (N_3610,N_2451,N_430);
nor U3611 (N_3611,N_1782,N_794);
nor U3612 (N_3612,N_218,N_2406);
xnor U3613 (N_3613,N_1162,N_2232);
nand U3614 (N_3614,N_129,N_98);
and U3615 (N_3615,N_649,N_1454);
and U3616 (N_3616,N_2128,N_1859);
nand U3617 (N_3617,N_606,N_1004);
or U3618 (N_3618,N_1469,N_2323);
or U3619 (N_3619,N_1598,N_1033);
and U3620 (N_3620,N_250,N_793);
and U3621 (N_3621,N_434,N_552);
or U3622 (N_3622,N_1414,N_1145);
nand U3623 (N_3623,N_2482,N_1860);
nor U3624 (N_3624,N_1887,N_2375);
xor U3625 (N_3625,N_2187,N_1682);
xnor U3626 (N_3626,N_193,N_102);
and U3627 (N_3627,N_1169,N_1999);
nand U3628 (N_3628,N_2477,N_1229);
nand U3629 (N_3629,N_1630,N_529);
or U3630 (N_3630,N_1685,N_173);
nor U3631 (N_3631,N_808,N_290);
and U3632 (N_3632,N_721,N_540);
or U3633 (N_3633,N_2389,N_124);
and U3634 (N_3634,N_1425,N_1230);
or U3635 (N_3635,N_756,N_994);
or U3636 (N_3636,N_954,N_1003);
nand U3637 (N_3637,N_1223,N_309);
xnor U3638 (N_3638,N_542,N_2209);
nand U3639 (N_3639,N_1610,N_1127);
nand U3640 (N_3640,N_788,N_843);
or U3641 (N_3641,N_2036,N_206);
and U3642 (N_3642,N_2020,N_1801);
or U3643 (N_3643,N_317,N_1957);
nor U3644 (N_3644,N_2154,N_466);
and U3645 (N_3645,N_2330,N_937);
or U3646 (N_3646,N_887,N_805);
or U3647 (N_3647,N_471,N_492);
or U3648 (N_3648,N_257,N_920);
xor U3649 (N_3649,N_820,N_1964);
and U3650 (N_3650,N_684,N_314);
nand U3651 (N_3651,N_934,N_1557);
or U3652 (N_3652,N_1567,N_1035);
nor U3653 (N_3653,N_983,N_517);
or U3654 (N_3654,N_473,N_99);
xor U3655 (N_3655,N_1543,N_537);
nand U3656 (N_3656,N_551,N_2288);
nor U3657 (N_3657,N_1948,N_1876);
nor U3658 (N_3658,N_1667,N_933);
or U3659 (N_3659,N_1073,N_2352);
xnor U3660 (N_3660,N_2077,N_2338);
nand U3661 (N_3661,N_1262,N_1116);
xor U3662 (N_3662,N_1734,N_1384);
nor U3663 (N_3663,N_2018,N_985);
xnor U3664 (N_3664,N_2455,N_815);
nor U3665 (N_3665,N_589,N_1113);
xnor U3666 (N_3666,N_261,N_1491);
nor U3667 (N_3667,N_477,N_576);
nand U3668 (N_3668,N_996,N_895);
nand U3669 (N_3669,N_1605,N_345);
nand U3670 (N_3670,N_1785,N_2351);
nor U3671 (N_3671,N_729,N_130);
nor U3672 (N_3672,N_2027,N_482);
xor U3673 (N_3673,N_2402,N_2378);
nand U3674 (N_3674,N_2492,N_1060);
nor U3675 (N_3675,N_683,N_238);
nand U3676 (N_3676,N_1146,N_1109);
or U3677 (N_3677,N_2202,N_2265);
nand U3678 (N_3678,N_2115,N_1451);
or U3679 (N_3679,N_602,N_1574);
or U3680 (N_3680,N_1783,N_1495);
or U3681 (N_3681,N_70,N_1445);
nand U3682 (N_3682,N_2129,N_221);
nand U3683 (N_3683,N_444,N_2497);
nor U3684 (N_3684,N_2059,N_46);
xnor U3685 (N_3685,N_1389,N_670);
nand U3686 (N_3686,N_1725,N_1609);
and U3687 (N_3687,N_457,N_644);
nand U3688 (N_3688,N_1616,N_2250);
nand U3689 (N_3689,N_1458,N_2047);
xnor U3690 (N_3690,N_525,N_838);
nand U3691 (N_3691,N_2060,N_1149);
nor U3692 (N_3692,N_204,N_1479);
or U3693 (N_3693,N_1664,N_1316);
xor U3694 (N_3694,N_1541,N_2362);
and U3695 (N_3695,N_438,N_2148);
nand U3696 (N_3696,N_406,N_397);
or U3697 (N_3697,N_1163,N_1802);
or U3698 (N_3698,N_1226,N_5);
xor U3699 (N_3699,N_1797,N_106);
nand U3700 (N_3700,N_1849,N_1395);
nand U3701 (N_3701,N_1748,N_1548);
and U3702 (N_3702,N_1053,N_588);
nand U3703 (N_3703,N_2342,N_1470);
xor U3704 (N_3704,N_554,N_338);
xnor U3705 (N_3705,N_65,N_2164);
nor U3706 (N_3706,N_1380,N_385);
or U3707 (N_3707,N_2249,N_2002);
xnor U3708 (N_3708,N_632,N_1090);
nand U3709 (N_3709,N_782,N_1413);
or U3710 (N_3710,N_2339,N_595);
or U3711 (N_3711,N_1464,N_8);
and U3712 (N_3712,N_661,N_180);
and U3713 (N_3713,N_842,N_236);
or U3714 (N_3714,N_1241,N_2426);
nor U3715 (N_3715,N_2006,N_227);
nand U3716 (N_3716,N_1601,N_1166);
nand U3717 (N_3717,N_628,N_2481);
and U3718 (N_3718,N_154,N_1615);
and U3719 (N_3719,N_1528,N_675);
xor U3720 (N_3720,N_779,N_1677);
xnor U3721 (N_3721,N_1392,N_726);
and U3722 (N_3722,N_1982,N_2126);
xnor U3723 (N_3723,N_1916,N_1626);
and U3724 (N_3724,N_614,N_501);
and U3725 (N_3725,N_1525,N_518);
nor U3726 (N_3726,N_2304,N_2456);
or U3727 (N_3727,N_234,N_1298);
or U3728 (N_3728,N_491,N_2270);
or U3729 (N_3729,N_1408,N_358);
or U3730 (N_3730,N_432,N_697);
nand U3731 (N_3731,N_433,N_1508);
or U3732 (N_3732,N_1089,N_1079);
or U3733 (N_3733,N_474,N_647);
and U3734 (N_3734,N_690,N_172);
nor U3735 (N_3735,N_2054,N_1355);
and U3736 (N_3736,N_307,N_2207);
xnor U3737 (N_3737,N_2499,N_2293);
and U3738 (N_3738,N_1290,N_868);
and U3739 (N_3739,N_373,N_1373);
or U3740 (N_3740,N_1268,N_14);
and U3741 (N_3741,N_1755,N_1817);
xor U3742 (N_3742,N_1935,N_1570);
nor U3743 (N_3743,N_1842,N_1128);
and U3744 (N_3744,N_2008,N_2053);
xnor U3745 (N_3745,N_828,N_414);
and U3746 (N_3746,N_1951,N_674);
or U3747 (N_3747,N_1258,N_1436);
nand U3748 (N_3748,N_1192,N_666);
or U3749 (N_3749,N_1190,N_400);
nor U3750 (N_3750,N_1322,N_2352);
or U3751 (N_3751,N_415,N_745);
nor U3752 (N_3752,N_1474,N_1268);
nand U3753 (N_3753,N_1820,N_1435);
nor U3754 (N_3754,N_2441,N_2087);
and U3755 (N_3755,N_320,N_750);
nor U3756 (N_3756,N_712,N_272);
nand U3757 (N_3757,N_131,N_799);
and U3758 (N_3758,N_998,N_1624);
or U3759 (N_3759,N_1618,N_248);
nand U3760 (N_3760,N_144,N_2120);
and U3761 (N_3761,N_1902,N_1765);
nor U3762 (N_3762,N_2278,N_975);
and U3763 (N_3763,N_2477,N_1028);
and U3764 (N_3764,N_698,N_1454);
and U3765 (N_3765,N_1896,N_1963);
nor U3766 (N_3766,N_1171,N_1632);
nand U3767 (N_3767,N_588,N_1223);
xnor U3768 (N_3768,N_949,N_177);
xor U3769 (N_3769,N_432,N_422);
nor U3770 (N_3770,N_308,N_1054);
nor U3771 (N_3771,N_737,N_2320);
and U3772 (N_3772,N_2138,N_1227);
nor U3773 (N_3773,N_985,N_800);
nand U3774 (N_3774,N_16,N_163);
and U3775 (N_3775,N_1401,N_274);
xor U3776 (N_3776,N_781,N_747);
xor U3777 (N_3777,N_2492,N_2390);
and U3778 (N_3778,N_1686,N_1480);
nand U3779 (N_3779,N_213,N_510);
nor U3780 (N_3780,N_2485,N_1836);
nand U3781 (N_3781,N_21,N_1917);
xnor U3782 (N_3782,N_2364,N_1992);
nand U3783 (N_3783,N_2271,N_1958);
xor U3784 (N_3784,N_314,N_200);
nand U3785 (N_3785,N_2376,N_766);
or U3786 (N_3786,N_2269,N_1700);
and U3787 (N_3787,N_560,N_1172);
nor U3788 (N_3788,N_2497,N_2025);
nor U3789 (N_3789,N_1608,N_1984);
and U3790 (N_3790,N_2454,N_1838);
and U3791 (N_3791,N_1989,N_1000);
and U3792 (N_3792,N_2299,N_2117);
nand U3793 (N_3793,N_353,N_1633);
nor U3794 (N_3794,N_789,N_2336);
and U3795 (N_3795,N_2018,N_1736);
xnor U3796 (N_3796,N_1918,N_1682);
xor U3797 (N_3797,N_2010,N_1526);
nor U3798 (N_3798,N_1158,N_790);
xor U3799 (N_3799,N_2455,N_1582);
and U3800 (N_3800,N_1811,N_1318);
and U3801 (N_3801,N_1155,N_1590);
and U3802 (N_3802,N_349,N_1837);
nand U3803 (N_3803,N_369,N_151);
xnor U3804 (N_3804,N_1048,N_1763);
nand U3805 (N_3805,N_2462,N_949);
or U3806 (N_3806,N_552,N_4);
xnor U3807 (N_3807,N_2175,N_846);
and U3808 (N_3808,N_1271,N_1191);
and U3809 (N_3809,N_642,N_1717);
and U3810 (N_3810,N_2249,N_190);
nor U3811 (N_3811,N_1180,N_1588);
xnor U3812 (N_3812,N_1314,N_693);
or U3813 (N_3813,N_1264,N_969);
xor U3814 (N_3814,N_1341,N_394);
xor U3815 (N_3815,N_638,N_858);
xor U3816 (N_3816,N_2394,N_1722);
or U3817 (N_3817,N_1400,N_1421);
xor U3818 (N_3818,N_2215,N_707);
nand U3819 (N_3819,N_1907,N_1333);
xor U3820 (N_3820,N_857,N_958);
and U3821 (N_3821,N_215,N_2412);
or U3822 (N_3822,N_602,N_2052);
and U3823 (N_3823,N_558,N_805);
nor U3824 (N_3824,N_950,N_1237);
or U3825 (N_3825,N_903,N_285);
nand U3826 (N_3826,N_2288,N_2024);
and U3827 (N_3827,N_1314,N_2355);
nand U3828 (N_3828,N_2211,N_1877);
xor U3829 (N_3829,N_1748,N_581);
nand U3830 (N_3830,N_110,N_1782);
xor U3831 (N_3831,N_2002,N_58);
or U3832 (N_3832,N_2292,N_1758);
xnor U3833 (N_3833,N_2348,N_2272);
and U3834 (N_3834,N_1752,N_2297);
or U3835 (N_3835,N_301,N_849);
and U3836 (N_3836,N_752,N_1112);
or U3837 (N_3837,N_1560,N_1744);
nand U3838 (N_3838,N_409,N_63);
and U3839 (N_3839,N_1839,N_1427);
xor U3840 (N_3840,N_133,N_530);
xnor U3841 (N_3841,N_1457,N_2364);
xnor U3842 (N_3842,N_334,N_2341);
nor U3843 (N_3843,N_626,N_1476);
and U3844 (N_3844,N_2483,N_886);
nor U3845 (N_3845,N_2399,N_791);
nand U3846 (N_3846,N_2475,N_1379);
or U3847 (N_3847,N_630,N_146);
or U3848 (N_3848,N_387,N_371);
xnor U3849 (N_3849,N_1332,N_1642);
nor U3850 (N_3850,N_244,N_1551);
xor U3851 (N_3851,N_132,N_1803);
xor U3852 (N_3852,N_982,N_1100);
and U3853 (N_3853,N_2178,N_843);
nand U3854 (N_3854,N_1734,N_380);
or U3855 (N_3855,N_689,N_2022);
nor U3856 (N_3856,N_1856,N_2325);
or U3857 (N_3857,N_992,N_454);
nand U3858 (N_3858,N_382,N_1985);
nor U3859 (N_3859,N_1419,N_764);
or U3860 (N_3860,N_1878,N_2452);
and U3861 (N_3861,N_1841,N_280);
xor U3862 (N_3862,N_231,N_596);
xor U3863 (N_3863,N_1893,N_528);
or U3864 (N_3864,N_272,N_1392);
or U3865 (N_3865,N_1196,N_1486);
xor U3866 (N_3866,N_316,N_956);
nor U3867 (N_3867,N_896,N_2118);
nand U3868 (N_3868,N_567,N_2174);
or U3869 (N_3869,N_355,N_1393);
and U3870 (N_3870,N_2387,N_2288);
xnor U3871 (N_3871,N_1166,N_744);
xor U3872 (N_3872,N_343,N_2007);
nand U3873 (N_3873,N_531,N_781);
nand U3874 (N_3874,N_179,N_1856);
nand U3875 (N_3875,N_501,N_1454);
xnor U3876 (N_3876,N_1481,N_326);
or U3877 (N_3877,N_1728,N_718);
or U3878 (N_3878,N_1935,N_668);
and U3879 (N_3879,N_497,N_759);
xnor U3880 (N_3880,N_1459,N_983);
xor U3881 (N_3881,N_50,N_1261);
and U3882 (N_3882,N_2010,N_44);
nor U3883 (N_3883,N_623,N_2277);
and U3884 (N_3884,N_1867,N_128);
nor U3885 (N_3885,N_576,N_2410);
nand U3886 (N_3886,N_1382,N_1282);
and U3887 (N_3887,N_1817,N_228);
and U3888 (N_3888,N_834,N_1823);
or U3889 (N_3889,N_1771,N_2482);
nor U3890 (N_3890,N_834,N_1959);
and U3891 (N_3891,N_2446,N_781);
nor U3892 (N_3892,N_2256,N_2081);
or U3893 (N_3893,N_192,N_211);
nand U3894 (N_3894,N_658,N_27);
nand U3895 (N_3895,N_303,N_390);
nor U3896 (N_3896,N_826,N_1235);
or U3897 (N_3897,N_1584,N_1974);
and U3898 (N_3898,N_2490,N_474);
nor U3899 (N_3899,N_1881,N_1436);
nor U3900 (N_3900,N_95,N_1272);
and U3901 (N_3901,N_695,N_1316);
and U3902 (N_3902,N_2344,N_2097);
nand U3903 (N_3903,N_2051,N_1690);
nor U3904 (N_3904,N_2120,N_1919);
or U3905 (N_3905,N_148,N_1744);
nand U3906 (N_3906,N_1556,N_890);
nand U3907 (N_3907,N_289,N_146);
or U3908 (N_3908,N_918,N_2222);
nor U3909 (N_3909,N_1329,N_422);
or U3910 (N_3910,N_1327,N_2397);
nor U3911 (N_3911,N_295,N_131);
nand U3912 (N_3912,N_152,N_2264);
or U3913 (N_3913,N_1563,N_1071);
or U3914 (N_3914,N_542,N_1796);
nand U3915 (N_3915,N_1948,N_188);
or U3916 (N_3916,N_859,N_586);
nand U3917 (N_3917,N_661,N_1175);
nor U3918 (N_3918,N_1672,N_1242);
or U3919 (N_3919,N_2012,N_1393);
or U3920 (N_3920,N_1659,N_1687);
or U3921 (N_3921,N_2445,N_994);
nor U3922 (N_3922,N_1151,N_808);
and U3923 (N_3923,N_842,N_1589);
nor U3924 (N_3924,N_1908,N_1153);
nand U3925 (N_3925,N_2049,N_27);
nor U3926 (N_3926,N_1818,N_425);
nor U3927 (N_3927,N_1578,N_1762);
and U3928 (N_3928,N_2232,N_1442);
or U3929 (N_3929,N_2213,N_552);
or U3930 (N_3930,N_1386,N_158);
nand U3931 (N_3931,N_188,N_148);
nor U3932 (N_3932,N_926,N_962);
nor U3933 (N_3933,N_2150,N_2112);
nor U3934 (N_3934,N_379,N_2045);
nor U3935 (N_3935,N_1606,N_1924);
and U3936 (N_3936,N_1723,N_1206);
nand U3937 (N_3937,N_769,N_1570);
xnor U3938 (N_3938,N_1303,N_1107);
or U3939 (N_3939,N_2121,N_600);
nor U3940 (N_3940,N_898,N_86);
and U3941 (N_3941,N_1828,N_2226);
and U3942 (N_3942,N_993,N_1324);
nand U3943 (N_3943,N_1306,N_1651);
nand U3944 (N_3944,N_1011,N_1930);
and U3945 (N_3945,N_1114,N_347);
nand U3946 (N_3946,N_1721,N_2397);
and U3947 (N_3947,N_1307,N_1709);
nor U3948 (N_3948,N_1345,N_542);
xor U3949 (N_3949,N_260,N_2302);
nor U3950 (N_3950,N_1944,N_1415);
nand U3951 (N_3951,N_1369,N_1269);
nor U3952 (N_3952,N_1688,N_184);
and U3953 (N_3953,N_201,N_1933);
and U3954 (N_3954,N_1564,N_427);
or U3955 (N_3955,N_1766,N_1142);
xor U3956 (N_3956,N_1971,N_1287);
and U3957 (N_3957,N_111,N_530);
nor U3958 (N_3958,N_1923,N_1863);
nand U3959 (N_3959,N_2059,N_238);
and U3960 (N_3960,N_931,N_1107);
and U3961 (N_3961,N_876,N_456);
or U3962 (N_3962,N_5,N_1277);
and U3963 (N_3963,N_1014,N_974);
nor U3964 (N_3964,N_2368,N_767);
xor U3965 (N_3965,N_1964,N_296);
nor U3966 (N_3966,N_1949,N_1984);
and U3967 (N_3967,N_2026,N_112);
and U3968 (N_3968,N_1657,N_1500);
nand U3969 (N_3969,N_1549,N_1060);
or U3970 (N_3970,N_107,N_2316);
or U3971 (N_3971,N_993,N_1092);
nor U3972 (N_3972,N_849,N_1052);
and U3973 (N_3973,N_1835,N_1353);
nor U3974 (N_3974,N_325,N_1147);
and U3975 (N_3975,N_182,N_1768);
nor U3976 (N_3976,N_603,N_1652);
and U3977 (N_3977,N_1908,N_1202);
or U3978 (N_3978,N_1416,N_1643);
nand U3979 (N_3979,N_655,N_811);
and U3980 (N_3980,N_2035,N_128);
nand U3981 (N_3981,N_1047,N_1509);
nand U3982 (N_3982,N_283,N_556);
nor U3983 (N_3983,N_701,N_3);
xnor U3984 (N_3984,N_1867,N_536);
nand U3985 (N_3985,N_2165,N_1487);
xor U3986 (N_3986,N_1261,N_611);
or U3987 (N_3987,N_237,N_266);
and U3988 (N_3988,N_1920,N_2465);
and U3989 (N_3989,N_535,N_2155);
nand U3990 (N_3990,N_760,N_2300);
nand U3991 (N_3991,N_1585,N_1072);
nand U3992 (N_3992,N_990,N_2100);
and U3993 (N_3993,N_1898,N_477);
or U3994 (N_3994,N_831,N_602);
and U3995 (N_3995,N_2470,N_1653);
xnor U3996 (N_3996,N_1862,N_28);
xor U3997 (N_3997,N_920,N_1982);
nand U3998 (N_3998,N_1501,N_1395);
and U3999 (N_3999,N_2226,N_1162);
xor U4000 (N_4000,N_1145,N_2496);
nand U4001 (N_4001,N_32,N_775);
nand U4002 (N_4002,N_718,N_1357);
xor U4003 (N_4003,N_206,N_2005);
or U4004 (N_4004,N_1456,N_876);
nand U4005 (N_4005,N_2223,N_1643);
or U4006 (N_4006,N_1110,N_1715);
nand U4007 (N_4007,N_2201,N_1008);
xor U4008 (N_4008,N_638,N_565);
or U4009 (N_4009,N_1518,N_1276);
or U4010 (N_4010,N_82,N_2327);
nand U4011 (N_4011,N_853,N_1001);
nor U4012 (N_4012,N_1137,N_759);
nor U4013 (N_4013,N_2208,N_1130);
and U4014 (N_4014,N_1507,N_973);
nor U4015 (N_4015,N_1144,N_1262);
nor U4016 (N_4016,N_1161,N_2348);
nor U4017 (N_4017,N_605,N_1899);
xnor U4018 (N_4018,N_1099,N_441);
or U4019 (N_4019,N_1374,N_1909);
xor U4020 (N_4020,N_1034,N_836);
xnor U4021 (N_4021,N_762,N_2121);
xnor U4022 (N_4022,N_791,N_338);
nand U4023 (N_4023,N_1788,N_853);
nor U4024 (N_4024,N_2122,N_1765);
nand U4025 (N_4025,N_863,N_2171);
and U4026 (N_4026,N_447,N_1418);
or U4027 (N_4027,N_777,N_647);
xor U4028 (N_4028,N_1358,N_2467);
or U4029 (N_4029,N_1896,N_1441);
nand U4030 (N_4030,N_888,N_2143);
nand U4031 (N_4031,N_803,N_102);
nor U4032 (N_4032,N_1490,N_734);
nand U4033 (N_4033,N_533,N_2155);
nand U4034 (N_4034,N_1154,N_2446);
nand U4035 (N_4035,N_344,N_1126);
and U4036 (N_4036,N_2072,N_777);
xor U4037 (N_4037,N_994,N_242);
xnor U4038 (N_4038,N_1580,N_1566);
nand U4039 (N_4039,N_1526,N_2155);
nand U4040 (N_4040,N_785,N_1344);
or U4041 (N_4041,N_1774,N_412);
and U4042 (N_4042,N_809,N_695);
and U4043 (N_4043,N_2333,N_849);
nand U4044 (N_4044,N_1773,N_1431);
or U4045 (N_4045,N_361,N_1972);
and U4046 (N_4046,N_1598,N_1825);
and U4047 (N_4047,N_2155,N_2283);
or U4048 (N_4048,N_1979,N_768);
and U4049 (N_4049,N_2079,N_881);
nand U4050 (N_4050,N_1981,N_2262);
nor U4051 (N_4051,N_683,N_1715);
nor U4052 (N_4052,N_184,N_448);
nor U4053 (N_4053,N_155,N_760);
nor U4054 (N_4054,N_1026,N_438);
or U4055 (N_4055,N_1576,N_133);
or U4056 (N_4056,N_2188,N_739);
nor U4057 (N_4057,N_817,N_1099);
nand U4058 (N_4058,N_449,N_1707);
or U4059 (N_4059,N_798,N_194);
nor U4060 (N_4060,N_2465,N_405);
or U4061 (N_4061,N_620,N_55);
and U4062 (N_4062,N_1720,N_123);
xor U4063 (N_4063,N_919,N_2054);
and U4064 (N_4064,N_2378,N_1685);
and U4065 (N_4065,N_2003,N_324);
nand U4066 (N_4066,N_1701,N_1127);
nand U4067 (N_4067,N_1168,N_1887);
xor U4068 (N_4068,N_1336,N_1801);
or U4069 (N_4069,N_1894,N_278);
and U4070 (N_4070,N_968,N_416);
xnor U4071 (N_4071,N_763,N_2070);
nor U4072 (N_4072,N_125,N_490);
nor U4073 (N_4073,N_1522,N_687);
and U4074 (N_4074,N_2276,N_1845);
xor U4075 (N_4075,N_724,N_1013);
nor U4076 (N_4076,N_1310,N_2258);
nor U4077 (N_4077,N_1311,N_1891);
nand U4078 (N_4078,N_1445,N_2111);
nor U4079 (N_4079,N_743,N_215);
xor U4080 (N_4080,N_1980,N_1474);
nand U4081 (N_4081,N_1287,N_2248);
and U4082 (N_4082,N_2439,N_1828);
xnor U4083 (N_4083,N_1533,N_1122);
or U4084 (N_4084,N_2273,N_761);
nor U4085 (N_4085,N_178,N_2330);
and U4086 (N_4086,N_699,N_1335);
xnor U4087 (N_4087,N_418,N_79);
nand U4088 (N_4088,N_555,N_1609);
xor U4089 (N_4089,N_1424,N_1384);
nor U4090 (N_4090,N_287,N_2291);
nand U4091 (N_4091,N_2192,N_2227);
xor U4092 (N_4092,N_2378,N_1037);
nand U4093 (N_4093,N_1847,N_2446);
nor U4094 (N_4094,N_2471,N_1886);
and U4095 (N_4095,N_476,N_1073);
nand U4096 (N_4096,N_315,N_1303);
xor U4097 (N_4097,N_649,N_1048);
or U4098 (N_4098,N_1210,N_1709);
or U4099 (N_4099,N_55,N_2307);
or U4100 (N_4100,N_690,N_2166);
nand U4101 (N_4101,N_1789,N_1357);
and U4102 (N_4102,N_2075,N_988);
nor U4103 (N_4103,N_325,N_1841);
nor U4104 (N_4104,N_1772,N_739);
xnor U4105 (N_4105,N_699,N_1682);
nor U4106 (N_4106,N_1305,N_483);
or U4107 (N_4107,N_2229,N_1846);
xor U4108 (N_4108,N_874,N_2326);
xnor U4109 (N_4109,N_19,N_477);
nor U4110 (N_4110,N_754,N_656);
nand U4111 (N_4111,N_1846,N_1580);
nand U4112 (N_4112,N_1459,N_1680);
xnor U4113 (N_4113,N_441,N_2374);
and U4114 (N_4114,N_1266,N_2316);
nand U4115 (N_4115,N_2307,N_1991);
xor U4116 (N_4116,N_1819,N_683);
nand U4117 (N_4117,N_201,N_1897);
nand U4118 (N_4118,N_390,N_111);
or U4119 (N_4119,N_48,N_466);
and U4120 (N_4120,N_2047,N_744);
xnor U4121 (N_4121,N_461,N_1369);
or U4122 (N_4122,N_1672,N_1049);
or U4123 (N_4123,N_1866,N_1513);
xor U4124 (N_4124,N_1028,N_1014);
and U4125 (N_4125,N_1084,N_222);
nand U4126 (N_4126,N_529,N_962);
nand U4127 (N_4127,N_60,N_1028);
or U4128 (N_4128,N_2170,N_1887);
and U4129 (N_4129,N_840,N_1087);
xor U4130 (N_4130,N_28,N_1629);
nor U4131 (N_4131,N_2053,N_2082);
and U4132 (N_4132,N_2009,N_2170);
xnor U4133 (N_4133,N_682,N_286);
nor U4134 (N_4134,N_598,N_869);
nand U4135 (N_4135,N_2212,N_1516);
xor U4136 (N_4136,N_1217,N_683);
or U4137 (N_4137,N_326,N_1020);
and U4138 (N_4138,N_1252,N_2109);
and U4139 (N_4139,N_664,N_1673);
and U4140 (N_4140,N_1259,N_727);
nand U4141 (N_4141,N_1670,N_2214);
nand U4142 (N_4142,N_579,N_1768);
nand U4143 (N_4143,N_1761,N_1580);
and U4144 (N_4144,N_1030,N_1544);
nand U4145 (N_4145,N_1937,N_1941);
xor U4146 (N_4146,N_1479,N_2350);
xnor U4147 (N_4147,N_365,N_1888);
nor U4148 (N_4148,N_1550,N_578);
and U4149 (N_4149,N_2299,N_472);
nor U4150 (N_4150,N_2339,N_1690);
and U4151 (N_4151,N_269,N_2265);
or U4152 (N_4152,N_1855,N_1951);
xor U4153 (N_4153,N_2067,N_567);
nor U4154 (N_4154,N_1426,N_2183);
nand U4155 (N_4155,N_2294,N_474);
or U4156 (N_4156,N_516,N_2197);
nor U4157 (N_4157,N_2050,N_1676);
or U4158 (N_4158,N_274,N_1295);
xnor U4159 (N_4159,N_558,N_950);
and U4160 (N_4160,N_820,N_589);
nand U4161 (N_4161,N_937,N_732);
or U4162 (N_4162,N_2255,N_1502);
and U4163 (N_4163,N_2338,N_2215);
and U4164 (N_4164,N_363,N_2181);
and U4165 (N_4165,N_2184,N_697);
or U4166 (N_4166,N_2267,N_92);
nor U4167 (N_4167,N_201,N_2180);
and U4168 (N_4168,N_362,N_1821);
xnor U4169 (N_4169,N_963,N_37);
and U4170 (N_4170,N_1130,N_1091);
or U4171 (N_4171,N_1193,N_2339);
nor U4172 (N_4172,N_971,N_2358);
xnor U4173 (N_4173,N_1196,N_2287);
nand U4174 (N_4174,N_1897,N_1525);
xnor U4175 (N_4175,N_30,N_279);
nor U4176 (N_4176,N_769,N_634);
and U4177 (N_4177,N_2411,N_698);
xnor U4178 (N_4178,N_46,N_423);
nand U4179 (N_4179,N_1951,N_2002);
or U4180 (N_4180,N_436,N_1053);
nor U4181 (N_4181,N_1983,N_2477);
nand U4182 (N_4182,N_1084,N_1799);
and U4183 (N_4183,N_17,N_1239);
nor U4184 (N_4184,N_2142,N_1854);
nor U4185 (N_4185,N_1412,N_1814);
and U4186 (N_4186,N_2316,N_1797);
or U4187 (N_4187,N_224,N_352);
xor U4188 (N_4188,N_189,N_2115);
nor U4189 (N_4189,N_1873,N_2319);
and U4190 (N_4190,N_931,N_2467);
nand U4191 (N_4191,N_960,N_1610);
nor U4192 (N_4192,N_460,N_2254);
nand U4193 (N_4193,N_930,N_624);
nand U4194 (N_4194,N_1461,N_855);
nor U4195 (N_4195,N_2466,N_1854);
xnor U4196 (N_4196,N_2145,N_1636);
nor U4197 (N_4197,N_629,N_1082);
nand U4198 (N_4198,N_1351,N_2194);
or U4199 (N_4199,N_1681,N_961);
nor U4200 (N_4200,N_281,N_78);
and U4201 (N_4201,N_1919,N_1968);
xor U4202 (N_4202,N_210,N_1366);
or U4203 (N_4203,N_1454,N_569);
xor U4204 (N_4204,N_399,N_211);
nand U4205 (N_4205,N_1044,N_143);
nor U4206 (N_4206,N_1369,N_1592);
nor U4207 (N_4207,N_2266,N_2167);
nor U4208 (N_4208,N_1249,N_1750);
nand U4209 (N_4209,N_1046,N_1715);
nand U4210 (N_4210,N_1445,N_1130);
and U4211 (N_4211,N_2086,N_158);
nand U4212 (N_4212,N_337,N_1028);
and U4213 (N_4213,N_959,N_584);
nand U4214 (N_4214,N_223,N_1333);
and U4215 (N_4215,N_2002,N_1044);
or U4216 (N_4216,N_426,N_1150);
nor U4217 (N_4217,N_2406,N_1882);
and U4218 (N_4218,N_279,N_2359);
nand U4219 (N_4219,N_2208,N_660);
or U4220 (N_4220,N_271,N_2062);
or U4221 (N_4221,N_345,N_130);
and U4222 (N_4222,N_1361,N_2476);
or U4223 (N_4223,N_123,N_421);
or U4224 (N_4224,N_1820,N_1458);
and U4225 (N_4225,N_56,N_1161);
nand U4226 (N_4226,N_1059,N_1898);
nor U4227 (N_4227,N_2008,N_386);
or U4228 (N_4228,N_2131,N_2283);
or U4229 (N_4229,N_69,N_2267);
xor U4230 (N_4230,N_669,N_1257);
xnor U4231 (N_4231,N_1264,N_1296);
xnor U4232 (N_4232,N_237,N_128);
nand U4233 (N_4233,N_1077,N_664);
nor U4234 (N_4234,N_1636,N_1290);
xor U4235 (N_4235,N_632,N_2150);
xnor U4236 (N_4236,N_214,N_247);
or U4237 (N_4237,N_34,N_2493);
or U4238 (N_4238,N_2323,N_1856);
nor U4239 (N_4239,N_249,N_415);
and U4240 (N_4240,N_781,N_1946);
nor U4241 (N_4241,N_1615,N_1695);
nor U4242 (N_4242,N_2235,N_1322);
xor U4243 (N_4243,N_1407,N_2287);
nor U4244 (N_4244,N_223,N_2194);
and U4245 (N_4245,N_2484,N_1125);
nor U4246 (N_4246,N_890,N_1868);
or U4247 (N_4247,N_1687,N_346);
nor U4248 (N_4248,N_1463,N_846);
nor U4249 (N_4249,N_1323,N_355);
xnor U4250 (N_4250,N_1833,N_2446);
xnor U4251 (N_4251,N_442,N_1464);
and U4252 (N_4252,N_1202,N_2487);
nor U4253 (N_4253,N_2404,N_2363);
xor U4254 (N_4254,N_1439,N_1398);
xnor U4255 (N_4255,N_486,N_144);
nor U4256 (N_4256,N_741,N_2087);
nand U4257 (N_4257,N_2123,N_1184);
or U4258 (N_4258,N_1514,N_977);
nand U4259 (N_4259,N_2076,N_2153);
nand U4260 (N_4260,N_1267,N_2355);
nor U4261 (N_4261,N_19,N_375);
and U4262 (N_4262,N_2230,N_1196);
or U4263 (N_4263,N_470,N_2421);
nor U4264 (N_4264,N_2157,N_2219);
or U4265 (N_4265,N_1017,N_1756);
or U4266 (N_4266,N_2096,N_1749);
xor U4267 (N_4267,N_1195,N_677);
nand U4268 (N_4268,N_1658,N_2373);
nand U4269 (N_4269,N_622,N_2047);
and U4270 (N_4270,N_476,N_540);
xnor U4271 (N_4271,N_1702,N_1270);
and U4272 (N_4272,N_19,N_2360);
nor U4273 (N_4273,N_663,N_94);
nand U4274 (N_4274,N_165,N_1986);
nor U4275 (N_4275,N_382,N_478);
xnor U4276 (N_4276,N_840,N_1428);
nand U4277 (N_4277,N_1234,N_2120);
xor U4278 (N_4278,N_890,N_1476);
and U4279 (N_4279,N_1977,N_383);
nand U4280 (N_4280,N_1586,N_806);
nor U4281 (N_4281,N_2021,N_918);
or U4282 (N_4282,N_1368,N_1901);
or U4283 (N_4283,N_868,N_1757);
xor U4284 (N_4284,N_2472,N_668);
nand U4285 (N_4285,N_1911,N_2167);
or U4286 (N_4286,N_1985,N_1275);
nor U4287 (N_4287,N_240,N_1001);
and U4288 (N_4288,N_81,N_506);
xnor U4289 (N_4289,N_155,N_2286);
and U4290 (N_4290,N_1505,N_264);
and U4291 (N_4291,N_270,N_296);
nand U4292 (N_4292,N_2139,N_1436);
and U4293 (N_4293,N_1745,N_1926);
and U4294 (N_4294,N_1301,N_2164);
xnor U4295 (N_4295,N_1904,N_331);
nand U4296 (N_4296,N_1883,N_834);
nor U4297 (N_4297,N_517,N_1291);
nor U4298 (N_4298,N_38,N_2362);
and U4299 (N_4299,N_2462,N_1809);
and U4300 (N_4300,N_550,N_1851);
or U4301 (N_4301,N_510,N_1460);
xor U4302 (N_4302,N_1329,N_15);
nor U4303 (N_4303,N_2374,N_1883);
and U4304 (N_4304,N_1574,N_759);
nor U4305 (N_4305,N_2293,N_390);
nor U4306 (N_4306,N_2134,N_237);
nand U4307 (N_4307,N_745,N_2254);
nor U4308 (N_4308,N_2205,N_50);
and U4309 (N_4309,N_734,N_1213);
and U4310 (N_4310,N_1047,N_408);
and U4311 (N_4311,N_2427,N_838);
or U4312 (N_4312,N_1531,N_1151);
nand U4313 (N_4313,N_1424,N_985);
nand U4314 (N_4314,N_134,N_39);
or U4315 (N_4315,N_195,N_1426);
xnor U4316 (N_4316,N_2314,N_256);
nand U4317 (N_4317,N_35,N_810);
xor U4318 (N_4318,N_842,N_697);
or U4319 (N_4319,N_1203,N_404);
xor U4320 (N_4320,N_519,N_1949);
nor U4321 (N_4321,N_1245,N_327);
nand U4322 (N_4322,N_1289,N_676);
or U4323 (N_4323,N_2304,N_1325);
and U4324 (N_4324,N_895,N_1919);
xor U4325 (N_4325,N_451,N_1815);
nand U4326 (N_4326,N_221,N_2137);
nand U4327 (N_4327,N_2406,N_1146);
and U4328 (N_4328,N_3,N_487);
xnor U4329 (N_4329,N_1409,N_282);
or U4330 (N_4330,N_2112,N_1920);
xnor U4331 (N_4331,N_612,N_1642);
or U4332 (N_4332,N_1366,N_1048);
or U4333 (N_4333,N_1950,N_489);
nand U4334 (N_4334,N_998,N_1232);
and U4335 (N_4335,N_2079,N_581);
nor U4336 (N_4336,N_1535,N_1610);
xnor U4337 (N_4337,N_227,N_1204);
or U4338 (N_4338,N_2326,N_2122);
or U4339 (N_4339,N_389,N_2473);
nor U4340 (N_4340,N_43,N_867);
and U4341 (N_4341,N_1350,N_2036);
xor U4342 (N_4342,N_1737,N_1893);
nor U4343 (N_4343,N_1031,N_2146);
xor U4344 (N_4344,N_2122,N_80);
xor U4345 (N_4345,N_1566,N_1783);
nor U4346 (N_4346,N_362,N_2209);
xor U4347 (N_4347,N_1034,N_628);
or U4348 (N_4348,N_1360,N_46);
or U4349 (N_4349,N_522,N_2187);
nand U4350 (N_4350,N_2324,N_1995);
nor U4351 (N_4351,N_1214,N_2104);
and U4352 (N_4352,N_2166,N_306);
nand U4353 (N_4353,N_1015,N_1771);
nor U4354 (N_4354,N_1534,N_34);
and U4355 (N_4355,N_1558,N_1547);
nand U4356 (N_4356,N_1382,N_374);
nand U4357 (N_4357,N_727,N_874);
xor U4358 (N_4358,N_2343,N_1632);
or U4359 (N_4359,N_1782,N_800);
nand U4360 (N_4360,N_1144,N_28);
or U4361 (N_4361,N_82,N_2408);
or U4362 (N_4362,N_50,N_810);
nand U4363 (N_4363,N_2171,N_574);
xor U4364 (N_4364,N_157,N_2483);
xnor U4365 (N_4365,N_2487,N_1062);
nor U4366 (N_4366,N_2294,N_58);
or U4367 (N_4367,N_837,N_2368);
or U4368 (N_4368,N_706,N_2209);
nor U4369 (N_4369,N_1013,N_1968);
nand U4370 (N_4370,N_311,N_440);
or U4371 (N_4371,N_817,N_2072);
xor U4372 (N_4372,N_1828,N_1463);
or U4373 (N_4373,N_485,N_295);
and U4374 (N_4374,N_1621,N_2160);
xnor U4375 (N_4375,N_2177,N_129);
and U4376 (N_4376,N_1433,N_1353);
or U4377 (N_4377,N_783,N_362);
nor U4378 (N_4378,N_1003,N_1502);
nor U4379 (N_4379,N_462,N_1712);
or U4380 (N_4380,N_1991,N_1560);
or U4381 (N_4381,N_993,N_1154);
nand U4382 (N_4382,N_1757,N_2382);
nand U4383 (N_4383,N_571,N_731);
or U4384 (N_4384,N_2120,N_802);
and U4385 (N_4385,N_1832,N_1290);
nor U4386 (N_4386,N_1600,N_786);
and U4387 (N_4387,N_2166,N_1537);
xor U4388 (N_4388,N_14,N_397);
xnor U4389 (N_4389,N_1071,N_1376);
xnor U4390 (N_4390,N_2003,N_1865);
or U4391 (N_4391,N_941,N_204);
and U4392 (N_4392,N_1088,N_959);
xnor U4393 (N_4393,N_621,N_1613);
nor U4394 (N_4394,N_2043,N_2205);
nor U4395 (N_4395,N_1032,N_387);
or U4396 (N_4396,N_514,N_1451);
nand U4397 (N_4397,N_649,N_453);
nor U4398 (N_4398,N_2210,N_789);
or U4399 (N_4399,N_2080,N_1617);
xor U4400 (N_4400,N_359,N_166);
or U4401 (N_4401,N_408,N_891);
nor U4402 (N_4402,N_2136,N_2042);
xnor U4403 (N_4403,N_614,N_1768);
nor U4404 (N_4404,N_2205,N_997);
or U4405 (N_4405,N_2251,N_232);
and U4406 (N_4406,N_1002,N_2198);
or U4407 (N_4407,N_864,N_2393);
xnor U4408 (N_4408,N_1806,N_2152);
nand U4409 (N_4409,N_1083,N_1308);
or U4410 (N_4410,N_1063,N_579);
nor U4411 (N_4411,N_1275,N_850);
nand U4412 (N_4412,N_240,N_1433);
xnor U4413 (N_4413,N_1820,N_2002);
and U4414 (N_4414,N_492,N_359);
nand U4415 (N_4415,N_2190,N_1206);
nand U4416 (N_4416,N_2016,N_1420);
xnor U4417 (N_4417,N_2256,N_689);
xor U4418 (N_4418,N_434,N_1087);
nand U4419 (N_4419,N_1091,N_2123);
or U4420 (N_4420,N_1445,N_1356);
nand U4421 (N_4421,N_1339,N_1292);
nand U4422 (N_4422,N_2094,N_1897);
or U4423 (N_4423,N_480,N_437);
nor U4424 (N_4424,N_986,N_938);
and U4425 (N_4425,N_1893,N_2422);
nand U4426 (N_4426,N_1119,N_1318);
and U4427 (N_4427,N_1996,N_2178);
and U4428 (N_4428,N_1203,N_1184);
xnor U4429 (N_4429,N_1505,N_1070);
and U4430 (N_4430,N_1808,N_1751);
xor U4431 (N_4431,N_549,N_278);
xnor U4432 (N_4432,N_1068,N_1220);
xnor U4433 (N_4433,N_446,N_59);
nor U4434 (N_4434,N_960,N_2268);
xor U4435 (N_4435,N_6,N_2164);
or U4436 (N_4436,N_1107,N_2147);
or U4437 (N_4437,N_1088,N_906);
or U4438 (N_4438,N_1803,N_53);
nand U4439 (N_4439,N_942,N_1890);
nand U4440 (N_4440,N_171,N_1811);
or U4441 (N_4441,N_1092,N_446);
or U4442 (N_4442,N_203,N_223);
nand U4443 (N_4443,N_2253,N_1277);
or U4444 (N_4444,N_990,N_2087);
and U4445 (N_4445,N_1442,N_1424);
xor U4446 (N_4446,N_2449,N_187);
or U4447 (N_4447,N_2451,N_2348);
and U4448 (N_4448,N_193,N_732);
and U4449 (N_4449,N_96,N_115);
nor U4450 (N_4450,N_1407,N_493);
xnor U4451 (N_4451,N_207,N_2184);
nor U4452 (N_4452,N_262,N_754);
nand U4453 (N_4453,N_1891,N_1885);
nor U4454 (N_4454,N_916,N_664);
xnor U4455 (N_4455,N_1826,N_1623);
and U4456 (N_4456,N_436,N_419);
and U4457 (N_4457,N_925,N_74);
nor U4458 (N_4458,N_722,N_233);
xor U4459 (N_4459,N_139,N_1667);
or U4460 (N_4460,N_726,N_2439);
nand U4461 (N_4461,N_1832,N_1748);
or U4462 (N_4462,N_1296,N_2391);
and U4463 (N_4463,N_1195,N_2478);
and U4464 (N_4464,N_1031,N_1708);
nand U4465 (N_4465,N_338,N_2331);
nand U4466 (N_4466,N_2166,N_1487);
nor U4467 (N_4467,N_619,N_1024);
and U4468 (N_4468,N_891,N_1932);
or U4469 (N_4469,N_2048,N_1440);
xor U4470 (N_4470,N_1143,N_517);
or U4471 (N_4471,N_1513,N_1161);
or U4472 (N_4472,N_200,N_2494);
or U4473 (N_4473,N_1041,N_2152);
nand U4474 (N_4474,N_1142,N_1144);
nor U4475 (N_4475,N_2376,N_89);
nor U4476 (N_4476,N_2407,N_2143);
and U4477 (N_4477,N_1570,N_264);
nand U4478 (N_4478,N_254,N_1286);
xor U4479 (N_4479,N_2099,N_621);
or U4480 (N_4480,N_2332,N_1303);
nor U4481 (N_4481,N_1602,N_708);
xor U4482 (N_4482,N_1292,N_703);
xnor U4483 (N_4483,N_1951,N_1498);
or U4484 (N_4484,N_2207,N_1512);
or U4485 (N_4485,N_1957,N_363);
or U4486 (N_4486,N_2391,N_956);
nand U4487 (N_4487,N_156,N_277);
nor U4488 (N_4488,N_975,N_483);
nor U4489 (N_4489,N_2480,N_1772);
nand U4490 (N_4490,N_2148,N_1784);
nand U4491 (N_4491,N_372,N_1087);
and U4492 (N_4492,N_594,N_1606);
nand U4493 (N_4493,N_1462,N_1125);
or U4494 (N_4494,N_1426,N_180);
nand U4495 (N_4495,N_1920,N_1154);
nor U4496 (N_4496,N_2354,N_1294);
nand U4497 (N_4497,N_2312,N_585);
or U4498 (N_4498,N_2395,N_502);
or U4499 (N_4499,N_2050,N_142);
or U4500 (N_4500,N_492,N_558);
or U4501 (N_4501,N_406,N_1373);
nand U4502 (N_4502,N_1962,N_2145);
and U4503 (N_4503,N_198,N_507);
nand U4504 (N_4504,N_32,N_1504);
and U4505 (N_4505,N_2364,N_2472);
and U4506 (N_4506,N_456,N_979);
and U4507 (N_4507,N_1114,N_99);
xnor U4508 (N_4508,N_514,N_1738);
or U4509 (N_4509,N_995,N_2328);
nor U4510 (N_4510,N_2135,N_1791);
xor U4511 (N_4511,N_831,N_1404);
or U4512 (N_4512,N_1983,N_2367);
xor U4513 (N_4513,N_1849,N_1117);
or U4514 (N_4514,N_29,N_2390);
nor U4515 (N_4515,N_27,N_1126);
nor U4516 (N_4516,N_1477,N_1050);
nor U4517 (N_4517,N_2403,N_2394);
nor U4518 (N_4518,N_795,N_1841);
nor U4519 (N_4519,N_1593,N_1206);
nor U4520 (N_4520,N_462,N_1411);
xnor U4521 (N_4521,N_1932,N_1210);
xor U4522 (N_4522,N_701,N_60);
nand U4523 (N_4523,N_236,N_2360);
xor U4524 (N_4524,N_1112,N_915);
and U4525 (N_4525,N_420,N_303);
or U4526 (N_4526,N_484,N_2107);
xnor U4527 (N_4527,N_2466,N_231);
xnor U4528 (N_4528,N_1576,N_381);
and U4529 (N_4529,N_2287,N_1132);
xnor U4530 (N_4530,N_477,N_1152);
xor U4531 (N_4531,N_2256,N_248);
nor U4532 (N_4532,N_2161,N_1768);
xnor U4533 (N_4533,N_2036,N_2192);
xor U4534 (N_4534,N_1842,N_1633);
or U4535 (N_4535,N_1863,N_1361);
and U4536 (N_4536,N_1641,N_704);
or U4537 (N_4537,N_897,N_1736);
nor U4538 (N_4538,N_718,N_143);
nand U4539 (N_4539,N_2346,N_527);
nor U4540 (N_4540,N_1013,N_1800);
and U4541 (N_4541,N_2447,N_2116);
xor U4542 (N_4542,N_2018,N_2024);
nand U4543 (N_4543,N_1024,N_955);
nand U4544 (N_4544,N_1034,N_314);
xor U4545 (N_4545,N_1121,N_2176);
xor U4546 (N_4546,N_809,N_950);
and U4547 (N_4547,N_580,N_704);
nor U4548 (N_4548,N_2257,N_1765);
nor U4549 (N_4549,N_1460,N_2038);
xnor U4550 (N_4550,N_1841,N_1282);
or U4551 (N_4551,N_1830,N_1133);
nand U4552 (N_4552,N_1935,N_836);
or U4553 (N_4553,N_140,N_443);
xor U4554 (N_4554,N_47,N_1369);
or U4555 (N_4555,N_1198,N_223);
nor U4556 (N_4556,N_316,N_1199);
or U4557 (N_4557,N_1967,N_1679);
and U4558 (N_4558,N_2289,N_74);
nor U4559 (N_4559,N_2350,N_2067);
and U4560 (N_4560,N_2013,N_2130);
nand U4561 (N_4561,N_1236,N_2205);
or U4562 (N_4562,N_187,N_1802);
nor U4563 (N_4563,N_974,N_264);
nand U4564 (N_4564,N_752,N_115);
nand U4565 (N_4565,N_1899,N_1072);
and U4566 (N_4566,N_266,N_318);
and U4567 (N_4567,N_863,N_390);
xor U4568 (N_4568,N_2116,N_542);
or U4569 (N_4569,N_619,N_278);
nand U4570 (N_4570,N_1640,N_315);
and U4571 (N_4571,N_441,N_815);
and U4572 (N_4572,N_2198,N_397);
nand U4573 (N_4573,N_1857,N_2123);
xor U4574 (N_4574,N_1243,N_1236);
nand U4575 (N_4575,N_1347,N_1927);
or U4576 (N_4576,N_1458,N_1922);
and U4577 (N_4577,N_2476,N_1539);
or U4578 (N_4578,N_1439,N_754);
xor U4579 (N_4579,N_209,N_153);
xor U4580 (N_4580,N_2235,N_681);
and U4581 (N_4581,N_446,N_2071);
nor U4582 (N_4582,N_2180,N_844);
xor U4583 (N_4583,N_811,N_2485);
xnor U4584 (N_4584,N_826,N_69);
xnor U4585 (N_4585,N_959,N_2264);
xnor U4586 (N_4586,N_97,N_1562);
xor U4587 (N_4587,N_1216,N_1090);
nand U4588 (N_4588,N_340,N_1096);
or U4589 (N_4589,N_652,N_102);
nand U4590 (N_4590,N_435,N_1425);
nand U4591 (N_4591,N_60,N_859);
nand U4592 (N_4592,N_2205,N_307);
nand U4593 (N_4593,N_1130,N_597);
xnor U4594 (N_4594,N_1572,N_180);
nor U4595 (N_4595,N_587,N_2065);
nand U4596 (N_4596,N_1457,N_415);
nand U4597 (N_4597,N_2250,N_681);
nand U4598 (N_4598,N_1759,N_51);
and U4599 (N_4599,N_774,N_1130);
nor U4600 (N_4600,N_1468,N_2384);
or U4601 (N_4601,N_727,N_69);
xor U4602 (N_4602,N_1187,N_947);
or U4603 (N_4603,N_200,N_692);
xor U4604 (N_4604,N_568,N_144);
nor U4605 (N_4605,N_466,N_2352);
nand U4606 (N_4606,N_1660,N_13);
nor U4607 (N_4607,N_789,N_299);
or U4608 (N_4608,N_995,N_430);
nor U4609 (N_4609,N_1284,N_2119);
or U4610 (N_4610,N_601,N_1493);
or U4611 (N_4611,N_284,N_2160);
xnor U4612 (N_4612,N_2499,N_510);
or U4613 (N_4613,N_802,N_1084);
nand U4614 (N_4614,N_2152,N_859);
nor U4615 (N_4615,N_1961,N_1672);
and U4616 (N_4616,N_860,N_285);
or U4617 (N_4617,N_647,N_738);
xnor U4618 (N_4618,N_1012,N_1532);
or U4619 (N_4619,N_871,N_1067);
nor U4620 (N_4620,N_1877,N_1955);
or U4621 (N_4621,N_182,N_2302);
xor U4622 (N_4622,N_1306,N_2041);
and U4623 (N_4623,N_1774,N_1728);
or U4624 (N_4624,N_1168,N_1709);
and U4625 (N_4625,N_2379,N_1764);
and U4626 (N_4626,N_1193,N_1262);
xor U4627 (N_4627,N_2353,N_2171);
or U4628 (N_4628,N_1250,N_2042);
or U4629 (N_4629,N_1281,N_1572);
nor U4630 (N_4630,N_164,N_1301);
or U4631 (N_4631,N_279,N_1738);
nor U4632 (N_4632,N_1313,N_893);
xnor U4633 (N_4633,N_1744,N_169);
nor U4634 (N_4634,N_507,N_1853);
nand U4635 (N_4635,N_1240,N_1151);
nor U4636 (N_4636,N_2028,N_1851);
xnor U4637 (N_4637,N_1075,N_1238);
nor U4638 (N_4638,N_830,N_2347);
xor U4639 (N_4639,N_927,N_1102);
nor U4640 (N_4640,N_1857,N_987);
nand U4641 (N_4641,N_855,N_1441);
or U4642 (N_4642,N_1614,N_1914);
and U4643 (N_4643,N_757,N_643);
nor U4644 (N_4644,N_2373,N_1198);
nand U4645 (N_4645,N_2378,N_2247);
xnor U4646 (N_4646,N_424,N_1915);
and U4647 (N_4647,N_364,N_2231);
nor U4648 (N_4648,N_925,N_1481);
nor U4649 (N_4649,N_1080,N_1177);
nand U4650 (N_4650,N_1759,N_523);
xor U4651 (N_4651,N_1757,N_1822);
nor U4652 (N_4652,N_512,N_33);
xnor U4653 (N_4653,N_1155,N_259);
nor U4654 (N_4654,N_1002,N_1166);
or U4655 (N_4655,N_1037,N_49);
and U4656 (N_4656,N_632,N_1042);
or U4657 (N_4657,N_1744,N_1432);
nand U4658 (N_4658,N_2499,N_1572);
nor U4659 (N_4659,N_410,N_739);
or U4660 (N_4660,N_630,N_2195);
or U4661 (N_4661,N_2373,N_1768);
nor U4662 (N_4662,N_2494,N_1730);
and U4663 (N_4663,N_366,N_293);
nor U4664 (N_4664,N_1720,N_582);
or U4665 (N_4665,N_1588,N_855);
xnor U4666 (N_4666,N_2004,N_1818);
or U4667 (N_4667,N_1435,N_1862);
and U4668 (N_4668,N_2292,N_1371);
or U4669 (N_4669,N_1984,N_83);
nand U4670 (N_4670,N_2239,N_569);
nand U4671 (N_4671,N_1817,N_756);
or U4672 (N_4672,N_209,N_2264);
or U4673 (N_4673,N_844,N_2097);
nor U4674 (N_4674,N_578,N_50);
xor U4675 (N_4675,N_386,N_840);
nand U4676 (N_4676,N_1839,N_1716);
nand U4677 (N_4677,N_1708,N_1645);
or U4678 (N_4678,N_1291,N_1223);
nor U4679 (N_4679,N_1704,N_869);
xnor U4680 (N_4680,N_288,N_1596);
or U4681 (N_4681,N_543,N_596);
and U4682 (N_4682,N_295,N_1606);
nor U4683 (N_4683,N_1998,N_877);
nand U4684 (N_4684,N_156,N_2486);
and U4685 (N_4685,N_1927,N_50);
nand U4686 (N_4686,N_498,N_1821);
nand U4687 (N_4687,N_594,N_2061);
or U4688 (N_4688,N_1871,N_126);
nand U4689 (N_4689,N_2103,N_2120);
xnor U4690 (N_4690,N_71,N_1340);
or U4691 (N_4691,N_131,N_568);
nand U4692 (N_4692,N_2313,N_391);
and U4693 (N_4693,N_628,N_1373);
nand U4694 (N_4694,N_1342,N_1039);
xor U4695 (N_4695,N_1539,N_551);
xnor U4696 (N_4696,N_1002,N_1615);
or U4697 (N_4697,N_1909,N_1044);
nand U4698 (N_4698,N_1042,N_877);
nand U4699 (N_4699,N_1838,N_2146);
xnor U4700 (N_4700,N_1569,N_316);
or U4701 (N_4701,N_587,N_1392);
nor U4702 (N_4702,N_416,N_1881);
and U4703 (N_4703,N_2455,N_2220);
and U4704 (N_4704,N_2239,N_220);
xnor U4705 (N_4705,N_1843,N_1574);
xor U4706 (N_4706,N_671,N_336);
nor U4707 (N_4707,N_213,N_1924);
or U4708 (N_4708,N_1051,N_1454);
xnor U4709 (N_4709,N_355,N_1132);
and U4710 (N_4710,N_1810,N_1041);
and U4711 (N_4711,N_2092,N_32);
nand U4712 (N_4712,N_1082,N_1012);
and U4713 (N_4713,N_1921,N_101);
and U4714 (N_4714,N_706,N_680);
nand U4715 (N_4715,N_305,N_770);
nor U4716 (N_4716,N_1525,N_1822);
nand U4717 (N_4717,N_1030,N_402);
or U4718 (N_4718,N_1190,N_1953);
xor U4719 (N_4719,N_977,N_390);
or U4720 (N_4720,N_162,N_861);
or U4721 (N_4721,N_1298,N_480);
xnor U4722 (N_4722,N_1487,N_1364);
nand U4723 (N_4723,N_707,N_2281);
xnor U4724 (N_4724,N_1926,N_1811);
or U4725 (N_4725,N_2220,N_1987);
nand U4726 (N_4726,N_1998,N_1585);
nand U4727 (N_4727,N_1758,N_236);
nor U4728 (N_4728,N_1924,N_1670);
nand U4729 (N_4729,N_318,N_2130);
and U4730 (N_4730,N_1228,N_2421);
nand U4731 (N_4731,N_1816,N_93);
and U4732 (N_4732,N_810,N_2489);
xnor U4733 (N_4733,N_1554,N_348);
and U4734 (N_4734,N_466,N_1995);
nor U4735 (N_4735,N_1639,N_117);
xnor U4736 (N_4736,N_1132,N_1926);
nand U4737 (N_4737,N_918,N_1435);
nor U4738 (N_4738,N_1380,N_200);
nand U4739 (N_4739,N_2379,N_1674);
nand U4740 (N_4740,N_608,N_1201);
nor U4741 (N_4741,N_178,N_1694);
xnor U4742 (N_4742,N_82,N_358);
xnor U4743 (N_4743,N_1563,N_415);
and U4744 (N_4744,N_1260,N_1831);
or U4745 (N_4745,N_430,N_1745);
xor U4746 (N_4746,N_1660,N_1581);
xor U4747 (N_4747,N_2142,N_2311);
nor U4748 (N_4748,N_661,N_2457);
nor U4749 (N_4749,N_398,N_2426);
or U4750 (N_4750,N_1137,N_857);
nor U4751 (N_4751,N_222,N_924);
or U4752 (N_4752,N_841,N_1038);
and U4753 (N_4753,N_1442,N_370);
and U4754 (N_4754,N_1761,N_121);
and U4755 (N_4755,N_892,N_2361);
and U4756 (N_4756,N_737,N_58);
xor U4757 (N_4757,N_715,N_726);
nand U4758 (N_4758,N_1330,N_1329);
and U4759 (N_4759,N_2067,N_1339);
nor U4760 (N_4760,N_533,N_936);
and U4761 (N_4761,N_2449,N_1602);
and U4762 (N_4762,N_1309,N_1518);
xor U4763 (N_4763,N_20,N_1024);
or U4764 (N_4764,N_1186,N_49);
or U4765 (N_4765,N_1984,N_544);
nor U4766 (N_4766,N_174,N_725);
and U4767 (N_4767,N_2058,N_1025);
nand U4768 (N_4768,N_1912,N_623);
nor U4769 (N_4769,N_1753,N_2319);
nand U4770 (N_4770,N_609,N_2003);
xnor U4771 (N_4771,N_103,N_146);
nand U4772 (N_4772,N_240,N_1690);
nor U4773 (N_4773,N_2057,N_1038);
nand U4774 (N_4774,N_1440,N_1784);
nor U4775 (N_4775,N_2125,N_485);
xnor U4776 (N_4776,N_2189,N_2294);
xor U4777 (N_4777,N_1381,N_931);
nand U4778 (N_4778,N_2399,N_209);
or U4779 (N_4779,N_440,N_2334);
nor U4780 (N_4780,N_1892,N_239);
nand U4781 (N_4781,N_1899,N_1792);
nand U4782 (N_4782,N_1615,N_578);
or U4783 (N_4783,N_561,N_1120);
nand U4784 (N_4784,N_1219,N_1757);
nor U4785 (N_4785,N_0,N_986);
nor U4786 (N_4786,N_117,N_1930);
and U4787 (N_4787,N_2158,N_1200);
and U4788 (N_4788,N_2450,N_973);
xor U4789 (N_4789,N_1917,N_1498);
and U4790 (N_4790,N_639,N_160);
xnor U4791 (N_4791,N_2488,N_2276);
xnor U4792 (N_4792,N_1928,N_1401);
nand U4793 (N_4793,N_2001,N_1666);
xor U4794 (N_4794,N_1390,N_2265);
and U4795 (N_4795,N_159,N_1175);
xnor U4796 (N_4796,N_2163,N_1700);
nand U4797 (N_4797,N_191,N_46);
nor U4798 (N_4798,N_655,N_1973);
nand U4799 (N_4799,N_1435,N_162);
and U4800 (N_4800,N_2089,N_2302);
and U4801 (N_4801,N_2188,N_560);
and U4802 (N_4802,N_2184,N_1355);
and U4803 (N_4803,N_2224,N_1233);
xor U4804 (N_4804,N_703,N_1145);
or U4805 (N_4805,N_35,N_225);
and U4806 (N_4806,N_1034,N_944);
or U4807 (N_4807,N_2034,N_514);
xnor U4808 (N_4808,N_1504,N_704);
nor U4809 (N_4809,N_2163,N_2351);
xor U4810 (N_4810,N_2347,N_854);
or U4811 (N_4811,N_900,N_1648);
and U4812 (N_4812,N_346,N_1053);
xnor U4813 (N_4813,N_557,N_188);
xnor U4814 (N_4814,N_2094,N_680);
xnor U4815 (N_4815,N_1157,N_2420);
nor U4816 (N_4816,N_856,N_509);
nand U4817 (N_4817,N_1582,N_1332);
nand U4818 (N_4818,N_601,N_1409);
xor U4819 (N_4819,N_528,N_870);
nand U4820 (N_4820,N_2402,N_2318);
nand U4821 (N_4821,N_1868,N_1029);
or U4822 (N_4822,N_129,N_1730);
and U4823 (N_4823,N_2181,N_1902);
or U4824 (N_4824,N_2038,N_973);
or U4825 (N_4825,N_844,N_391);
or U4826 (N_4826,N_976,N_1781);
or U4827 (N_4827,N_2070,N_1407);
and U4828 (N_4828,N_1727,N_167);
nor U4829 (N_4829,N_2428,N_124);
nor U4830 (N_4830,N_422,N_2478);
xnor U4831 (N_4831,N_770,N_2274);
or U4832 (N_4832,N_852,N_346);
or U4833 (N_4833,N_2343,N_300);
or U4834 (N_4834,N_156,N_2096);
xor U4835 (N_4835,N_1267,N_1458);
nor U4836 (N_4836,N_491,N_830);
nor U4837 (N_4837,N_1185,N_645);
xnor U4838 (N_4838,N_2304,N_924);
nor U4839 (N_4839,N_692,N_263);
xor U4840 (N_4840,N_1477,N_263);
xnor U4841 (N_4841,N_1133,N_1230);
or U4842 (N_4842,N_814,N_1393);
nand U4843 (N_4843,N_347,N_144);
xnor U4844 (N_4844,N_147,N_607);
nor U4845 (N_4845,N_270,N_1175);
or U4846 (N_4846,N_274,N_2483);
or U4847 (N_4847,N_2111,N_820);
nand U4848 (N_4848,N_838,N_1357);
nand U4849 (N_4849,N_367,N_1425);
xnor U4850 (N_4850,N_1934,N_13);
xnor U4851 (N_4851,N_1488,N_1120);
nand U4852 (N_4852,N_1054,N_244);
nor U4853 (N_4853,N_1847,N_1487);
nor U4854 (N_4854,N_1369,N_2260);
xnor U4855 (N_4855,N_1594,N_1017);
and U4856 (N_4856,N_1698,N_1313);
nand U4857 (N_4857,N_1167,N_1716);
or U4858 (N_4858,N_1030,N_1617);
or U4859 (N_4859,N_2461,N_206);
or U4860 (N_4860,N_821,N_2037);
nand U4861 (N_4861,N_1244,N_1935);
and U4862 (N_4862,N_1198,N_2159);
nor U4863 (N_4863,N_318,N_730);
and U4864 (N_4864,N_2268,N_453);
nor U4865 (N_4865,N_2370,N_827);
and U4866 (N_4866,N_542,N_954);
or U4867 (N_4867,N_1027,N_2318);
xnor U4868 (N_4868,N_382,N_195);
nor U4869 (N_4869,N_1617,N_893);
or U4870 (N_4870,N_268,N_508);
or U4871 (N_4871,N_2156,N_2089);
xor U4872 (N_4872,N_1974,N_583);
nor U4873 (N_4873,N_2421,N_20);
and U4874 (N_4874,N_1681,N_1762);
or U4875 (N_4875,N_952,N_476);
or U4876 (N_4876,N_2475,N_1555);
nor U4877 (N_4877,N_735,N_945);
or U4878 (N_4878,N_1460,N_637);
nand U4879 (N_4879,N_2120,N_2138);
or U4880 (N_4880,N_2095,N_1366);
and U4881 (N_4881,N_1241,N_1199);
xnor U4882 (N_4882,N_518,N_1028);
nor U4883 (N_4883,N_1615,N_2226);
nand U4884 (N_4884,N_1545,N_536);
nor U4885 (N_4885,N_1212,N_803);
and U4886 (N_4886,N_1921,N_2029);
and U4887 (N_4887,N_1377,N_1128);
nand U4888 (N_4888,N_2319,N_2215);
nor U4889 (N_4889,N_1836,N_627);
nand U4890 (N_4890,N_608,N_1705);
xnor U4891 (N_4891,N_346,N_710);
xnor U4892 (N_4892,N_1308,N_1482);
or U4893 (N_4893,N_2111,N_348);
or U4894 (N_4894,N_1906,N_2099);
or U4895 (N_4895,N_2066,N_2369);
nand U4896 (N_4896,N_876,N_1818);
and U4897 (N_4897,N_1180,N_295);
xnor U4898 (N_4898,N_2468,N_2124);
xor U4899 (N_4899,N_1300,N_1700);
nand U4900 (N_4900,N_1322,N_924);
nand U4901 (N_4901,N_1815,N_1167);
or U4902 (N_4902,N_2326,N_2);
nand U4903 (N_4903,N_1489,N_2377);
and U4904 (N_4904,N_323,N_1156);
xnor U4905 (N_4905,N_35,N_1802);
or U4906 (N_4906,N_1764,N_1748);
nor U4907 (N_4907,N_1188,N_1518);
and U4908 (N_4908,N_1707,N_819);
and U4909 (N_4909,N_64,N_2198);
nor U4910 (N_4910,N_1116,N_1848);
xnor U4911 (N_4911,N_1186,N_2006);
nand U4912 (N_4912,N_97,N_2404);
and U4913 (N_4913,N_2106,N_238);
nand U4914 (N_4914,N_884,N_1663);
or U4915 (N_4915,N_2320,N_1108);
and U4916 (N_4916,N_1981,N_1160);
or U4917 (N_4917,N_455,N_2100);
xnor U4918 (N_4918,N_1923,N_2003);
nand U4919 (N_4919,N_2110,N_2162);
nor U4920 (N_4920,N_1230,N_1480);
and U4921 (N_4921,N_2387,N_630);
nor U4922 (N_4922,N_802,N_2368);
nand U4923 (N_4923,N_42,N_2090);
nand U4924 (N_4924,N_407,N_2261);
nor U4925 (N_4925,N_2214,N_2132);
nor U4926 (N_4926,N_303,N_1567);
xor U4927 (N_4927,N_2436,N_1906);
nor U4928 (N_4928,N_1206,N_2248);
or U4929 (N_4929,N_1996,N_1794);
xnor U4930 (N_4930,N_1409,N_969);
nor U4931 (N_4931,N_1843,N_1822);
nor U4932 (N_4932,N_1325,N_399);
or U4933 (N_4933,N_1807,N_645);
xor U4934 (N_4934,N_663,N_1865);
and U4935 (N_4935,N_1968,N_720);
nor U4936 (N_4936,N_1090,N_1365);
or U4937 (N_4937,N_1445,N_566);
nor U4938 (N_4938,N_2169,N_827);
xnor U4939 (N_4939,N_1009,N_2063);
and U4940 (N_4940,N_194,N_2141);
or U4941 (N_4941,N_562,N_488);
nand U4942 (N_4942,N_1761,N_266);
nand U4943 (N_4943,N_295,N_217);
and U4944 (N_4944,N_1767,N_1817);
nor U4945 (N_4945,N_509,N_295);
and U4946 (N_4946,N_153,N_967);
nor U4947 (N_4947,N_562,N_1732);
nand U4948 (N_4948,N_2390,N_2368);
or U4949 (N_4949,N_2419,N_2177);
and U4950 (N_4950,N_354,N_792);
xor U4951 (N_4951,N_1905,N_657);
nand U4952 (N_4952,N_135,N_698);
nor U4953 (N_4953,N_1339,N_2044);
xor U4954 (N_4954,N_389,N_2065);
nand U4955 (N_4955,N_1264,N_2495);
xor U4956 (N_4956,N_494,N_2262);
xnor U4957 (N_4957,N_1446,N_705);
and U4958 (N_4958,N_635,N_407);
or U4959 (N_4959,N_1953,N_2120);
nor U4960 (N_4960,N_1211,N_2016);
nand U4961 (N_4961,N_2104,N_2258);
and U4962 (N_4962,N_2358,N_205);
nand U4963 (N_4963,N_1647,N_1245);
and U4964 (N_4964,N_2233,N_56);
nor U4965 (N_4965,N_1255,N_1458);
nor U4966 (N_4966,N_2310,N_2196);
nand U4967 (N_4967,N_2039,N_469);
nand U4968 (N_4968,N_2408,N_319);
nor U4969 (N_4969,N_890,N_701);
nand U4970 (N_4970,N_173,N_380);
and U4971 (N_4971,N_1560,N_7);
or U4972 (N_4972,N_1073,N_505);
or U4973 (N_4973,N_2115,N_1225);
xor U4974 (N_4974,N_1755,N_260);
nand U4975 (N_4975,N_978,N_1195);
and U4976 (N_4976,N_1117,N_1536);
xnor U4977 (N_4977,N_1206,N_966);
nand U4978 (N_4978,N_466,N_2329);
or U4979 (N_4979,N_1450,N_1995);
nor U4980 (N_4980,N_693,N_819);
nand U4981 (N_4981,N_374,N_1384);
nor U4982 (N_4982,N_1448,N_2139);
nand U4983 (N_4983,N_2276,N_55);
and U4984 (N_4984,N_131,N_1117);
xnor U4985 (N_4985,N_2119,N_1802);
and U4986 (N_4986,N_737,N_869);
nor U4987 (N_4987,N_1811,N_1402);
nor U4988 (N_4988,N_2499,N_1669);
or U4989 (N_4989,N_1887,N_2119);
or U4990 (N_4990,N_2134,N_665);
and U4991 (N_4991,N_664,N_2327);
nand U4992 (N_4992,N_315,N_2086);
nor U4993 (N_4993,N_552,N_998);
xnor U4994 (N_4994,N_1459,N_1601);
nor U4995 (N_4995,N_643,N_1973);
xor U4996 (N_4996,N_1210,N_1319);
and U4997 (N_4997,N_486,N_422);
nand U4998 (N_4998,N_488,N_1729);
nor U4999 (N_4999,N_86,N_1989);
nor UO_0 (O_0,N_4994,N_4304);
xor UO_1 (O_1,N_3813,N_4452);
nand UO_2 (O_2,N_3617,N_4855);
nand UO_3 (O_3,N_3794,N_3954);
nor UO_4 (O_4,N_3938,N_4661);
and UO_5 (O_5,N_2511,N_3978);
xor UO_6 (O_6,N_4430,N_4130);
nor UO_7 (O_7,N_2953,N_3588);
and UO_8 (O_8,N_2743,N_2865);
nor UO_9 (O_9,N_4822,N_3920);
nand UO_10 (O_10,N_4815,N_4962);
xor UO_11 (O_11,N_3304,N_4140);
and UO_12 (O_12,N_4239,N_2972);
and UO_13 (O_13,N_4720,N_2947);
or UO_14 (O_14,N_4235,N_3838);
nand UO_15 (O_15,N_4112,N_3550);
xor UO_16 (O_16,N_3715,N_4639);
or UO_17 (O_17,N_4001,N_2885);
nand UO_18 (O_18,N_3496,N_3258);
xor UO_19 (O_19,N_2775,N_3773);
or UO_20 (O_20,N_4447,N_3171);
nand UO_21 (O_21,N_2712,N_2505);
nand UO_22 (O_22,N_2561,N_2662);
or UO_23 (O_23,N_2679,N_2813);
nand UO_24 (O_24,N_4148,N_4467);
xor UO_25 (O_25,N_2855,N_4921);
nor UO_26 (O_26,N_4719,N_3118);
xor UO_27 (O_27,N_2532,N_2526);
and UO_28 (O_28,N_3030,N_3193);
nand UO_29 (O_29,N_4552,N_3102);
nor UO_30 (O_30,N_3014,N_2769);
nand UO_31 (O_31,N_3517,N_4224);
nand UO_32 (O_32,N_2710,N_4081);
and UO_33 (O_33,N_4648,N_4972);
nand UO_34 (O_34,N_2605,N_3015);
and UO_35 (O_35,N_2849,N_3600);
and UO_36 (O_36,N_3971,N_3204);
xor UO_37 (O_37,N_4849,N_4656);
xnor UO_38 (O_38,N_4966,N_2755);
or UO_39 (O_39,N_2727,N_3417);
nand UO_40 (O_40,N_3634,N_2623);
xor UO_41 (O_41,N_3261,N_3993);
nand UO_42 (O_42,N_2581,N_3828);
nor UO_43 (O_43,N_3620,N_2576);
xnor UO_44 (O_44,N_2758,N_4135);
and UO_45 (O_45,N_2669,N_4716);
or UO_46 (O_46,N_4958,N_4366);
or UO_47 (O_47,N_3393,N_3104);
nand UO_48 (O_48,N_2541,N_3155);
xnor UO_49 (O_49,N_3016,N_4423);
xor UO_50 (O_50,N_2837,N_3101);
and UO_51 (O_51,N_2725,N_3282);
nor UO_52 (O_52,N_3005,N_3175);
nor UO_53 (O_53,N_4441,N_4047);
and UO_54 (O_54,N_3312,N_4395);
nand UO_55 (O_55,N_3464,N_4957);
xnor UO_56 (O_56,N_4787,N_4125);
nor UO_57 (O_57,N_4085,N_2995);
xor UO_58 (O_58,N_2931,N_4477);
or UO_59 (O_59,N_3737,N_2859);
nor UO_60 (O_60,N_4955,N_4836);
and UO_61 (O_61,N_3513,N_2513);
xnor UO_62 (O_62,N_4898,N_3927);
xnor UO_63 (O_63,N_3348,N_4666);
nor UO_64 (O_64,N_3113,N_3568);
or UO_65 (O_65,N_2694,N_3824);
nor UO_66 (O_66,N_2984,N_2603);
xnor UO_67 (O_67,N_3560,N_3749);
nor UO_68 (O_68,N_4878,N_2839);
or UO_69 (O_69,N_3409,N_4056);
xor UO_70 (O_70,N_3472,N_4654);
nor UO_71 (O_71,N_4290,N_3112);
nor UO_72 (O_72,N_3148,N_4548);
nor UO_73 (O_73,N_4371,N_4884);
xnor UO_74 (O_74,N_3557,N_4843);
or UO_75 (O_75,N_3637,N_4383);
nand UO_76 (O_76,N_3952,N_3992);
and UO_77 (O_77,N_4759,N_4949);
or UO_78 (O_78,N_4786,N_4317);
nor UO_79 (O_79,N_4509,N_2858);
xnor UO_80 (O_80,N_2740,N_3013);
or UO_81 (O_81,N_4812,N_4160);
xor UO_82 (O_82,N_4920,N_4458);
and UO_83 (O_83,N_3621,N_4252);
xnor UO_84 (O_84,N_2934,N_4418);
nor UO_85 (O_85,N_3270,N_3453);
nand UO_86 (O_86,N_4192,N_4892);
or UO_87 (O_87,N_3514,N_3173);
xnor UO_88 (O_88,N_4109,N_3615);
xnor UO_89 (O_89,N_3049,N_3073);
or UO_90 (O_90,N_2973,N_4816);
or UO_91 (O_91,N_3524,N_2748);
nand UO_92 (O_92,N_2506,N_3987);
or UO_93 (O_93,N_4205,N_3571);
xor UO_94 (O_94,N_3010,N_3279);
xor UO_95 (O_95,N_2570,N_3144);
or UO_96 (O_96,N_2556,N_2990);
nor UO_97 (O_97,N_4705,N_4040);
or UO_98 (O_98,N_2978,N_3050);
or UO_99 (O_99,N_3252,N_4963);
and UO_100 (O_100,N_3475,N_3832);
nor UO_101 (O_101,N_2803,N_3149);
or UO_102 (O_102,N_4583,N_4473);
and UO_103 (O_103,N_4905,N_4498);
and UO_104 (O_104,N_4675,N_3969);
xor UO_105 (O_105,N_3973,N_3400);
or UO_106 (O_106,N_2763,N_4210);
or UO_107 (O_107,N_3291,N_2881);
nor UO_108 (O_108,N_3853,N_3157);
and UO_109 (O_109,N_4536,N_2687);
xor UO_110 (O_110,N_4731,N_3280);
and UO_111 (O_111,N_4243,N_2771);
nand UO_112 (O_112,N_4922,N_3242);
and UO_113 (O_113,N_4015,N_4723);
nor UO_114 (O_114,N_4690,N_4895);
and UO_115 (O_115,N_2644,N_2820);
and UO_116 (O_116,N_4273,N_4261);
nand UO_117 (O_117,N_3369,N_2912);
nor UO_118 (O_118,N_4439,N_3146);
nand UO_119 (O_119,N_4483,N_4960);
nand UO_120 (O_120,N_3061,N_3167);
xnor UO_121 (O_121,N_3081,N_4770);
or UO_122 (O_122,N_3551,N_3895);
nand UO_123 (O_123,N_4686,N_2982);
nand UO_124 (O_124,N_4060,N_3166);
or UO_125 (O_125,N_4861,N_2515);
or UO_126 (O_126,N_4944,N_4097);
nor UO_127 (O_127,N_4581,N_3616);
or UO_128 (O_128,N_4121,N_3484);
nor UO_129 (O_129,N_3124,N_3186);
nor UO_130 (O_130,N_4607,N_3974);
nor UO_131 (O_131,N_4104,N_3923);
or UO_132 (O_132,N_3355,N_2974);
xor UO_133 (O_133,N_3911,N_3998);
nand UO_134 (O_134,N_4755,N_2921);
and UO_135 (O_135,N_4840,N_3950);
nand UO_136 (O_136,N_4881,N_3088);
nand UO_137 (O_137,N_3758,N_3098);
nor UO_138 (O_138,N_3858,N_3461);
nor UO_139 (O_139,N_2557,N_4127);
or UO_140 (O_140,N_4292,N_3351);
nand UO_141 (O_141,N_4242,N_4739);
nor UO_142 (O_142,N_4709,N_4351);
nor UO_143 (O_143,N_2760,N_3667);
or UO_144 (O_144,N_4942,N_4071);
nor UO_145 (O_145,N_4198,N_2943);
and UO_146 (O_146,N_3189,N_3001);
xor UO_147 (O_147,N_3532,N_4456);
nor UO_148 (O_148,N_3859,N_4562);
nand UO_149 (O_149,N_4334,N_4584);
xor UO_150 (O_150,N_2502,N_3784);
or UO_151 (O_151,N_3276,N_4976);
nor UO_152 (O_152,N_3678,N_3890);
and UO_153 (O_153,N_3985,N_4543);
nand UO_154 (O_154,N_3856,N_2764);
xnor UO_155 (O_155,N_3506,N_4505);
nand UO_156 (O_156,N_2503,N_3546);
or UO_157 (O_157,N_3966,N_3537);
nor UO_158 (O_158,N_4801,N_2626);
nor UO_159 (O_159,N_3185,N_3746);
or UO_160 (O_160,N_2717,N_4478);
and UO_161 (O_161,N_2542,N_3357);
xor UO_162 (O_162,N_4064,N_4194);
xnor UO_163 (O_163,N_2949,N_2574);
nand UO_164 (O_164,N_2660,N_3446);
nand UO_165 (O_165,N_3863,N_4480);
nand UO_166 (O_166,N_3306,N_4529);
and UO_167 (O_167,N_3130,N_4689);
nor UO_168 (O_168,N_4379,N_4876);
and UO_169 (O_169,N_2566,N_3239);
xor UO_170 (O_170,N_4868,N_3988);
or UO_171 (O_171,N_3322,N_3121);
xnor UO_172 (O_172,N_4841,N_4636);
nor UO_173 (O_173,N_3378,N_2983);
xnor UO_174 (O_174,N_3728,N_4974);
and UO_175 (O_175,N_4819,N_3143);
xor UO_176 (O_176,N_3986,N_3395);
nor UO_177 (O_177,N_4400,N_4680);
nand UO_178 (O_178,N_2935,N_4390);
nand UO_179 (O_179,N_4618,N_3575);
xor UO_180 (O_180,N_2737,N_4487);
nand UO_181 (O_181,N_3533,N_4434);
and UO_182 (O_182,N_3724,N_2834);
xnor UO_183 (O_183,N_2980,N_2564);
or UO_184 (O_184,N_4901,N_2565);
or UO_185 (O_185,N_3751,N_4391);
or UO_186 (O_186,N_3222,N_4282);
nand UO_187 (O_187,N_2728,N_4714);
and UO_188 (O_188,N_2696,N_3714);
nor UO_189 (O_189,N_4363,N_3495);
xor UO_190 (O_190,N_4613,N_3117);
or UO_191 (O_191,N_2835,N_3661);
nand UO_192 (O_192,N_4332,N_4186);
nand UO_193 (O_193,N_2939,N_2703);
or UO_194 (O_194,N_4416,N_4511);
and UO_195 (O_195,N_4577,N_4322);
xnor UO_196 (O_196,N_4154,N_2531);
and UO_197 (O_197,N_4540,N_4392);
nand UO_198 (O_198,N_2779,N_3577);
nor UO_199 (O_199,N_2537,N_3094);
and UO_200 (O_200,N_4526,N_3596);
nand UO_201 (O_201,N_4927,N_3518);
nand UO_202 (O_202,N_2613,N_3755);
nand UO_203 (O_203,N_2938,N_4095);
xnor UO_204 (O_204,N_3300,N_4212);
and UO_205 (O_205,N_2945,N_4555);
xor UO_206 (O_206,N_3690,N_2827);
and UO_207 (O_207,N_3093,N_3350);
nor UO_208 (O_208,N_3640,N_3169);
and UO_209 (O_209,N_3008,N_4805);
and UO_210 (O_210,N_2645,N_3114);
xor UO_211 (O_211,N_4522,N_4157);
or UO_212 (O_212,N_3426,N_3949);
or UO_213 (O_213,N_3980,N_3319);
or UO_214 (O_214,N_4472,N_3877);
xor UO_215 (O_215,N_2894,N_3862);
nand UO_216 (O_216,N_2967,N_3745);
nand UO_217 (O_217,N_4621,N_2846);
nor UO_218 (O_218,N_2977,N_3221);
and UO_219 (O_219,N_3731,N_3067);
and UO_220 (O_220,N_3959,N_3111);
nor UO_221 (O_221,N_4496,N_3935);
or UO_222 (O_222,N_3501,N_3074);
nand UO_223 (O_223,N_2724,N_4236);
xnor UO_224 (O_224,N_4204,N_3766);
nand UO_225 (O_225,N_4729,N_2545);
nor UO_226 (O_226,N_2655,N_3960);
nand UO_227 (O_227,N_4406,N_3630);
nand UO_228 (O_228,N_4435,N_3254);
nand UO_229 (O_229,N_4455,N_4077);
nand UO_230 (O_230,N_3344,N_3761);
nor UO_231 (O_231,N_4409,N_2514);
and UO_232 (O_232,N_3359,N_4655);
nand UO_233 (O_233,N_4411,N_3583);
and UO_234 (O_234,N_3500,N_3597);
nor UO_235 (O_235,N_2954,N_2516);
or UO_236 (O_236,N_3585,N_4486);
or UO_237 (O_237,N_4059,N_4580);
or UO_238 (O_238,N_3796,N_2691);
and UO_239 (O_239,N_4407,N_3153);
xor UO_240 (O_240,N_2787,N_2897);
and UO_241 (O_241,N_3841,N_2530);
and UO_242 (O_242,N_2709,N_2994);
xor UO_243 (O_243,N_2930,N_4785);
or UO_244 (O_244,N_2936,N_4325);
xnor UO_245 (O_245,N_4168,N_3701);
and UO_246 (O_246,N_3991,N_2772);
or UO_247 (O_247,N_4365,N_4838);
nand UO_248 (O_248,N_3411,N_4067);
and UO_249 (O_249,N_3570,N_4510);
or UO_250 (O_250,N_3769,N_4679);
nand UO_251 (O_251,N_2925,N_3914);
or UO_252 (O_252,N_2731,N_4030);
nand UO_253 (O_253,N_4432,N_2720);
or UO_254 (O_254,N_3401,N_2843);
nor UO_255 (O_255,N_2852,N_4339);
nor UO_256 (O_256,N_4802,N_3817);
or UO_257 (O_257,N_3848,N_3662);
nor UO_258 (O_258,N_4142,N_2909);
or UO_259 (O_259,N_3671,N_3463);
and UO_260 (O_260,N_3882,N_4065);
nor UO_261 (O_261,N_3201,N_4667);
nand UO_262 (O_262,N_3739,N_3347);
or UO_263 (O_263,N_4996,N_3139);
xnor UO_264 (O_264,N_3246,N_3628);
or UO_265 (O_265,N_3483,N_4576);
nand UO_266 (O_266,N_4867,N_4269);
nand UO_267 (O_267,N_4875,N_2879);
xor UO_268 (O_268,N_2906,N_2826);
and UO_269 (O_269,N_3843,N_2601);
xor UO_270 (O_270,N_2955,N_3024);
or UO_271 (O_271,N_3984,N_3133);
nor UO_272 (O_272,N_3445,N_4171);
nand UO_273 (O_273,N_2598,N_4634);
xor UO_274 (O_274,N_4203,N_2887);
nor UO_275 (O_275,N_4305,N_4683);
nand UO_276 (O_276,N_3574,N_3044);
nor UO_277 (O_277,N_4389,N_3754);
nor UO_278 (O_278,N_4935,N_4315);
or UO_279 (O_279,N_4567,N_2810);
nor UO_280 (O_280,N_3591,N_3011);
and UO_281 (O_281,N_3336,N_4845);
nand UO_282 (O_282,N_2525,N_4162);
nand UO_283 (O_283,N_3786,N_3934);
xor UO_284 (O_284,N_2988,N_4992);
nand UO_285 (O_285,N_3815,N_2933);
nor UO_286 (O_286,N_3314,N_2721);
nand UO_287 (O_287,N_4596,N_3612);
or UO_288 (O_288,N_3177,N_4402);
nor UO_289 (O_289,N_2884,N_4479);
or UO_290 (O_290,N_4023,N_2577);
nor UO_291 (O_291,N_2559,N_3244);
nand UO_292 (O_292,N_4002,N_3569);
or UO_293 (O_293,N_3217,N_4831);
or UO_294 (O_294,N_3165,N_4330);
xor UO_295 (O_295,N_3002,N_4344);
nand UO_296 (O_296,N_3084,N_2856);
nand UO_297 (O_297,N_3553,N_3631);
nor UO_298 (O_298,N_3607,N_4068);
xnor UO_299 (O_299,N_3190,N_4775);
or UO_300 (O_300,N_2784,N_3384);
nand UO_301 (O_301,N_2579,N_4941);
and UO_302 (O_302,N_4232,N_4123);
nand UO_303 (O_303,N_4143,N_3414);
or UO_304 (O_304,N_3200,N_2742);
nor UO_305 (O_305,N_3224,N_4764);
or UO_306 (O_306,N_4961,N_4249);
xor UO_307 (O_307,N_3147,N_3581);
or UO_308 (O_308,N_2658,N_4381);
and UO_309 (O_309,N_3519,N_3599);
nor UO_310 (O_310,N_4553,N_2653);
and UO_311 (O_311,N_4166,N_4124);
and UO_312 (O_312,N_4426,N_4488);
or UO_313 (O_313,N_4532,N_2848);
nor UO_314 (O_314,N_4279,N_2635);
or UO_315 (O_315,N_2636,N_2588);
and UO_316 (O_316,N_4076,N_2971);
or UO_317 (O_317,N_4404,N_2845);
and UO_318 (O_318,N_4700,N_3869);
xor UO_319 (O_319,N_2918,N_2951);
and UO_320 (O_320,N_2993,N_2882);
or UO_321 (O_321,N_2761,N_2965);
nor UO_322 (O_322,N_4018,N_4664);
nand UO_323 (O_323,N_3850,N_3844);
nand UO_324 (O_324,N_4453,N_4748);
xor UO_325 (O_325,N_4285,N_4189);
nor UO_326 (O_326,N_4632,N_2788);
nor UO_327 (O_327,N_2888,N_3435);
or UO_328 (O_328,N_4470,N_2901);
and UO_329 (O_329,N_2500,N_4699);
nand UO_330 (O_330,N_4169,N_2591);
and UO_331 (O_331,N_3213,N_4028);
or UO_332 (O_332,N_4973,N_4464);
xnor UO_333 (O_333,N_3902,N_2975);
nand UO_334 (O_334,N_4115,N_4153);
and UO_335 (O_335,N_2738,N_4804);
and UO_336 (O_336,N_4009,N_4570);
and UO_337 (O_337,N_3305,N_3590);
and UO_338 (O_338,N_2668,N_4846);
or UO_339 (O_339,N_4909,N_4046);
nand UO_340 (O_340,N_3712,N_3362);
or UO_341 (O_341,N_4750,N_4616);
and UO_342 (O_342,N_3156,N_4244);
xnor UO_343 (O_343,N_3682,N_4155);
or UO_344 (O_344,N_3394,N_4156);
or UO_345 (O_345,N_2981,N_4779);
and UO_346 (O_346,N_4531,N_3127);
and UO_347 (O_347,N_4987,N_2783);
or UO_348 (O_348,N_3290,N_2842);
nand UO_349 (O_349,N_4674,N_4427);
xnor UO_350 (O_350,N_4482,N_2942);
nand UO_351 (O_351,N_3215,N_2656);
xor UO_352 (O_352,N_4638,N_2549);
and UO_353 (O_353,N_4415,N_2819);
and UO_354 (O_354,N_4223,N_4721);
nor UO_355 (O_355,N_3818,N_3835);
and UO_356 (O_356,N_4926,N_3564);
xor UO_357 (O_357,N_4743,N_4329);
nand UO_358 (O_358,N_4858,N_4676);
or UO_359 (O_359,N_3037,N_2908);
and UO_360 (O_360,N_3642,N_3083);
nand UO_361 (O_361,N_3708,N_4247);
nor UO_362 (O_362,N_4545,N_2723);
nor UO_363 (O_363,N_4995,N_3075);
nand UO_364 (O_364,N_4631,N_3372);
nand UO_365 (O_365,N_4007,N_3479);
nor UO_366 (O_366,N_3499,N_4066);
and UO_367 (O_367,N_4137,N_3736);
xnor UO_368 (O_368,N_2527,N_3163);
and UO_369 (O_369,N_3220,N_2754);
or UO_370 (O_370,N_3626,N_4762);
xnor UO_371 (O_371,N_3100,N_3757);
nand UO_372 (O_372,N_4736,N_4600);
xor UO_373 (O_373,N_3181,N_4735);
xor UO_374 (O_374,N_2631,N_2841);
or UO_375 (O_375,N_3875,N_4408);
or UO_376 (O_376,N_3376,N_3137);
xnor UO_377 (O_377,N_4188,N_4180);
xor UO_378 (O_378,N_3006,N_4597);
nor UO_379 (O_379,N_2714,N_4219);
nor UO_380 (O_380,N_4611,N_3272);
and UO_381 (O_381,N_3465,N_4113);
and UO_382 (O_382,N_4501,N_3691);
nor UO_383 (O_383,N_2781,N_3331);
xnor UO_384 (O_384,N_3756,N_4930);
nand UO_385 (O_385,N_4346,N_3498);
and UO_386 (O_386,N_2562,N_3543);
nand UO_387 (O_387,N_3752,N_3374);
and UO_388 (O_388,N_2929,N_4701);
xnor UO_389 (O_389,N_2666,N_2773);
xor UO_390 (O_390,N_3129,N_3965);
and UO_391 (O_391,N_4145,N_4283);
nor UO_392 (O_392,N_3764,N_3115);
and UO_393 (O_393,N_4533,N_3438);
and UO_394 (O_394,N_2850,N_3197);
and UO_395 (O_395,N_2800,N_3063);
and UO_396 (O_396,N_3549,N_4763);
nor UO_397 (O_397,N_3142,N_2550);
nor UO_398 (O_398,N_3026,N_3644);
and UO_399 (O_399,N_4733,N_4889);
and UO_400 (O_400,N_3576,N_4376);
nand UO_401 (O_401,N_3211,N_4254);
nand UO_402 (O_402,N_2637,N_4181);
and UO_403 (O_403,N_2958,N_4959);
and UO_404 (O_404,N_4516,N_4842);
or UO_405 (O_405,N_4818,N_4038);
nor UO_406 (O_406,N_3939,N_2711);
nor UO_407 (O_407,N_3562,N_3179);
nor UO_408 (O_408,N_3338,N_4817);
xnor UO_409 (O_409,N_4590,N_4673);
nor UO_410 (O_410,N_2927,N_4575);
or UO_411 (O_411,N_4605,N_4658);
or UO_412 (O_412,N_2560,N_3141);
xnor UO_413 (O_413,N_4998,N_2739);
nor UO_414 (O_414,N_2670,N_4378);
and UO_415 (O_415,N_2815,N_3779);
nand UO_416 (O_416,N_3799,N_3436);
nand UO_417 (O_417,N_4270,N_4375);
nor UO_418 (O_418,N_4176,N_2890);
nor UO_419 (O_419,N_4592,N_2649);
and UO_420 (O_420,N_4692,N_2534);
nor UO_421 (O_421,N_4754,N_3065);
nor UO_422 (O_422,N_4820,N_4678);
nor UO_423 (O_423,N_4360,N_4051);
nand UO_424 (O_424,N_3509,N_3485);
or UO_425 (O_425,N_3656,N_3434);
nor UO_426 (O_426,N_2708,N_3140);
nor UO_427 (O_427,N_3210,N_3316);
or UO_428 (O_428,N_3289,N_4425);
nand UO_429 (O_429,N_3808,N_4221);
or UO_430 (O_430,N_3932,N_3629);
and UO_431 (O_431,N_3018,N_3154);
nor UO_432 (O_432,N_2790,N_2540);
xnor UO_433 (O_433,N_2699,N_3921);
and UO_434 (O_434,N_3486,N_3516);
nand UO_435 (O_435,N_4094,N_4758);
xor UO_436 (O_436,N_3313,N_4852);
and UO_437 (O_437,N_3759,N_2940);
xor UO_438 (O_438,N_4010,N_2998);
or UO_439 (O_439,N_4267,N_2677);
and UO_440 (O_440,N_3929,N_4257);
nor UO_441 (O_441,N_3493,N_3223);
nor UO_442 (O_442,N_3652,N_3572);
or UO_443 (O_443,N_3420,N_2966);
nor UO_444 (O_444,N_3323,N_4620);
nand UO_445 (O_445,N_4560,N_2634);
xor UO_446 (O_446,N_4525,N_3800);
nand UO_447 (O_447,N_4373,N_2844);
and UO_448 (O_448,N_3337,N_3439);
or UO_449 (O_449,N_3721,N_4837);
and UO_450 (O_450,N_3849,N_4713);
nand UO_451 (O_451,N_3593,N_2611);
nor UO_452 (O_452,N_4238,N_3311);
or UO_453 (O_453,N_4049,N_4608);
nor UO_454 (O_454,N_3457,N_4016);
or UO_455 (O_455,N_3447,N_3602);
and UO_456 (O_456,N_4965,N_3025);
or UO_457 (O_457,N_3688,N_4551);
xnor UO_458 (O_458,N_4380,N_2609);
nand UO_459 (O_459,N_2767,N_3734);
and UO_460 (O_460,N_3529,N_3366);
xor UO_461 (O_461,N_4940,N_2624);
nand UO_462 (O_462,N_4256,N_3090);
or UO_463 (O_463,N_2950,N_2555);
xor UO_464 (O_464,N_2917,N_3326);
or UO_465 (O_465,N_2745,N_3277);
nor UO_466 (O_466,N_3041,N_4208);
xor UO_467 (O_467,N_3912,N_3055);
nand UO_468 (O_468,N_4165,N_3078);
nor UO_469 (O_469,N_3310,N_3383);
nor UO_470 (O_470,N_3332,N_3885);
xor UO_471 (O_471,N_3528,N_4101);
and UO_472 (O_472,N_3870,N_4564);
nand UO_473 (O_473,N_3466,N_2547);
or UO_474 (O_474,N_3043,N_3716);
nor UO_475 (O_475,N_2682,N_3029);
or UO_476 (O_476,N_2878,N_4687);
xor UO_477 (O_477,N_4882,N_4945);
or UO_478 (O_478,N_4179,N_4436);
nand UO_479 (O_479,N_2896,N_4336);
nor UO_480 (O_480,N_2713,N_2785);
nor UO_481 (O_481,N_4727,N_4088);
or UO_482 (O_482,N_2757,N_3131);
nand UO_483 (O_483,N_2695,N_3294);
nor UO_484 (O_484,N_3012,N_2774);
and UO_485 (O_485,N_4215,N_4000);
nand UO_486 (O_486,N_3095,N_3653);
and UO_487 (O_487,N_4640,N_2684);
xnor UO_488 (O_488,N_2831,N_3723);
nor UO_489 (O_489,N_3535,N_4997);
xor UO_490 (O_490,N_3389,N_3975);
xnor UO_491 (O_491,N_4653,N_3789);
nor UO_492 (O_492,N_4309,N_4444);
nand UO_493 (O_493,N_4494,N_3624);
and UO_494 (O_494,N_4158,N_4445);
and UO_495 (O_495,N_4414,N_3227);
or UO_496 (O_496,N_3982,N_4627);
nor UO_497 (O_497,N_3738,N_4092);
nand UO_498 (O_498,N_4303,N_4193);
and UO_499 (O_499,N_3618,N_2868);
nor UO_500 (O_500,N_4796,N_2512);
and UO_501 (O_501,N_4784,N_4977);
or UO_502 (O_502,N_3742,N_3397);
or UO_503 (O_503,N_3391,N_4428);
nor UO_504 (O_504,N_4610,N_3473);
nor UO_505 (O_505,N_4724,N_4118);
nand UO_506 (O_506,N_3944,N_4844);
xnor UO_507 (O_507,N_4136,N_4569);
xnor UO_508 (O_508,N_4806,N_4103);
xnor UO_509 (O_509,N_4187,N_3398);
nand UO_510 (O_510,N_3997,N_4268);
and UO_511 (O_511,N_2964,N_3260);
nand UO_512 (O_512,N_4912,N_3253);
nand UO_513 (O_513,N_3767,N_4745);
xor UO_514 (O_514,N_4246,N_2572);
xor UO_515 (O_515,N_2715,N_3170);
and UO_516 (O_516,N_4832,N_4311);
or UO_517 (O_517,N_3510,N_4730);
xor UO_518 (O_518,N_4021,N_4662);
nor UO_519 (O_519,N_3508,N_4100);
and UO_520 (O_520,N_2812,N_4915);
or UO_521 (O_521,N_3660,N_2768);
or UO_522 (O_522,N_4020,N_3491);
or UO_523 (O_523,N_4043,N_4749);
and UO_524 (O_524,N_3867,N_4936);
and UO_525 (O_525,N_4307,N_4466);
or UO_526 (O_526,N_3782,N_2628);
or UO_527 (O_527,N_4220,N_4042);
and UO_528 (O_528,N_4925,N_2698);
nand UO_529 (O_529,N_4598,N_3884);
nor UO_530 (O_530,N_2928,N_4826);
xnor UO_531 (O_531,N_3428,N_3456);
and UO_532 (O_532,N_3654,N_3899);
xor UO_533 (O_533,N_2678,N_2674);
nand UO_534 (O_534,N_2829,N_4800);
xor UO_535 (O_535,N_3274,N_3448);
and UO_536 (O_536,N_2697,N_3733);
nand UO_537 (O_537,N_3547,N_3881);
and UO_538 (O_538,N_2833,N_3196);
xnor UO_539 (O_539,N_3873,N_2919);
nor UO_540 (O_540,N_2640,N_3017);
or UO_541 (O_541,N_3138,N_3490);
xnor UO_542 (O_542,N_3257,N_3342);
xnor UO_543 (O_543,N_3299,N_4542);
nand UO_544 (O_544,N_4984,N_4013);
nand UO_545 (O_545,N_4358,N_3830);
nand UO_546 (O_546,N_3056,N_3622);
nand UO_547 (O_547,N_3636,N_4629);
and UO_548 (O_548,N_4211,N_4233);
or UO_549 (O_549,N_2932,N_3649);
or UO_550 (O_550,N_3579,N_3926);
nor UO_551 (O_551,N_4546,N_4893);
nor UO_552 (O_552,N_2867,N_3989);
or UO_553 (O_553,N_3249,N_4834);
nand UO_554 (O_554,N_4790,N_3718);
nor UO_555 (O_555,N_2880,N_3686);
and UO_556 (O_556,N_4711,N_3031);
nor UO_557 (O_557,N_4601,N_3022);
and UO_558 (O_558,N_2801,N_3288);
xor UO_559 (O_559,N_2863,N_3776);
or UO_560 (O_560,N_3937,N_2573);
nand UO_561 (O_561,N_4116,N_4641);
nand UO_562 (O_562,N_4350,N_3837);
nand UO_563 (O_563,N_3488,N_3216);
nand UO_564 (O_564,N_3505,N_4728);
nand UO_565 (O_565,N_4110,N_3416);
and UO_566 (O_566,N_4659,N_3470);
or UO_567 (O_567,N_3788,N_4253);
or UO_568 (O_568,N_4900,N_3335);
or UO_569 (O_569,N_4767,N_4359);
nor UO_570 (O_570,N_3064,N_3857);
nor UO_571 (O_571,N_3028,N_3385);
nand UO_572 (O_572,N_4122,N_2922);
xnor UO_573 (O_573,N_4776,N_3936);
and UO_574 (O_574,N_4696,N_3777);
xor UO_575 (O_575,N_4693,N_3241);
nand UO_576 (O_576,N_4207,N_4947);
or UO_577 (O_577,N_2582,N_3471);
xor UO_578 (O_578,N_3459,N_4294);
and UO_579 (O_579,N_4566,N_2600);
and UO_580 (O_580,N_4386,N_4005);
xnor UO_581 (O_581,N_2730,N_3105);
nand UO_582 (O_582,N_3632,N_2741);
xnor UO_583 (O_583,N_2807,N_3027);
xnor UO_584 (O_584,N_3979,N_4603);
xor UO_585 (O_585,N_4265,N_3668);
xor UO_586 (O_586,N_2756,N_2766);
xor UO_587 (O_587,N_4864,N_2509);
nor UO_588 (O_588,N_4668,N_4139);
or UO_589 (O_589,N_4163,N_4412);
and UO_590 (O_590,N_3702,N_3038);
and UO_591 (O_591,N_4704,N_4929);
nor UO_592 (O_592,N_3172,N_4277);
and UO_593 (O_593,N_3387,N_2948);
and UO_594 (O_594,N_3047,N_3020);
xor UO_595 (O_595,N_4794,N_3555);
nand UO_596 (O_596,N_3497,N_2587);
nand UO_597 (O_597,N_3605,N_3807);
nor UO_598 (O_598,N_3176,N_4321);
and UO_599 (O_599,N_2693,N_2508);
xor UO_600 (O_600,N_4829,N_3245);
nor UO_601 (O_601,N_4493,N_4465);
xor UO_602 (O_602,N_4287,N_3639);
nand UO_603 (O_603,N_2999,N_4196);
nand UO_604 (O_604,N_3968,N_4369);
nor UO_605 (O_605,N_4384,N_3135);
and UO_606 (O_606,N_4554,N_3487);
nand UO_607 (O_607,N_4856,N_3208);
xor UO_608 (O_608,N_4272,N_3108);
nand UO_609 (O_609,N_4174,N_3840);
nand UO_610 (O_610,N_4541,N_3092);
and UO_611 (O_611,N_4968,N_4823);
nand UO_612 (O_612,N_4964,N_4619);
xnor UO_613 (O_613,N_3693,N_4070);
or UO_614 (O_614,N_4565,N_3119);
or UO_615 (O_615,N_4771,N_4732);
xor UO_616 (O_616,N_4086,N_2510);
or UO_617 (O_617,N_3298,N_3089);
and UO_618 (O_618,N_4141,N_4792);
or UO_619 (O_619,N_3151,N_4150);
and UO_620 (O_620,N_4222,N_4185);
and UO_621 (O_621,N_2604,N_3233);
xor UO_622 (O_622,N_4032,N_4506);
nor UO_623 (O_623,N_3765,N_3036);
and UO_624 (O_624,N_4885,N_3334);
xnor UO_625 (O_625,N_4345,N_2796);
nor UO_626 (O_626,N_4326,N_2673);
or UO_627 (O_627,N_3343,N_2782);
nor UO_628 (O_628,N_3259,N_3823);
nand UO_629 (O_629,N_2568,N_2593);
nor UO_630 (O_630,N_3821,N_2642);
nor UO_631 (O_631,N_2571,N_3068);
nor UO_632 (O_632,N_3803,N_2809);
nor UO_633 (O_633,N_2719,N_3806);
or UO_634 (O_634,N_3234,N_4420);
or UO_635 (O_635,N_3449,N_3771);
and UO_636 (O_636,N_4578,N_3243);
and UO_637 (O_637,N_3191,N_3705);
xor UO_638 (O_638,N_4460,N_4083);
nand UO_639 (O_639,N_3595,N_3696);
or UO_640 (O_640,N_3916,N_4951);
or UO_641 (O_641,N_3946,N_3819);
or UO_642 (O_642,N_2961,N_2970);
nor UO_643 (O_643,N_4450,N_3103);
nor UO_644 (O_644,N_3611,N_2686);
xor UO_645 (O_645,N_3918,N_4172);
or UO_646 (O_646,N_4873,N_3633);
nor UO_647 (O_647,N_4923,N_4938);
and UO_648 (O_648,N_3042,N_4499);
xnor UO_649 (O_649,N_3330,N_4685);
or UO_650 (O_650,N_4293,N_3900);
xor UO_651 (O_651,N_2794,N_3933);
nor UO_652 (O_652,N_3598,N_4825);
and UO_653 (O_653,N_3046,N_2539);
xor UO_654 (O_654,N_4523,N_3392);
nor UO_655 (O_655,N_3674,N_2962);
and UO_656 (O_656,N_4799,N_4328);
nor UO_657 (O_657,N_3866,N_3536);
and UO_658 (O_658,N_4320,N_4862);
and UO_659 (O_659,N_4475,N_2553);
and UO_660 (O_660,N_4626,N_3943);
nor UO_661 (O_661,N_3023,N_3080);
and UO_662 (O_662,N_4617,N_2517);
nand UO_663 (O_663,N_3956,N_4512);
nor UO_664 (O_664,N_4585,N_3880);
or UO_665 (O_665,N_3897,N_3909);
nor UO_666 (O_666,N_4370,N_4872);
or UO_667 (O_667,N_2959,N_4119);
or UO_668 (O_668,N_2722,N_3106);
nand UO_669 (O_669,N_4006,N_4348);
xor UO_670 (O_670,N_3825,N_4218);
nand UO_671 (O_671,N_4913,N_2596);
nand UO_672 (O_672,N_3886,N_3273);
nor UO_673 (O_673,N_4549,N_4946);
and UO_674 (O_674,N_3325,N_3264);
or UO_675 (O_675,N_4352,N_4538);
or UO_676 (O_676,N_4887,N_3212);
nor UO_677 (O_677,N_2543,N_3232);
nand UO_678 (O_678,N_2651,N_3539);
xnor UO_679 (O_679,N_3876,N_3531);
xnor UO_680 (O_680,N_3474,N_3542);
nor UO_681 (O_681,N_3683,N_3515);
nor UO_682 (O_682,N_3820,N_4401);
or UO_683 (O_683,N_4789,N_4890);
nor UO_684 (O_684,N_4191,N_4574);
or UO_685 (O_685,N_4982,N_4202);
or UO_686 (O_686,N_2617,N_2536);
nor UO_687 (O_687,N_4393,N_2913);
nor UO_688 (O_688,N_2899,N_4783);
nand UO_689 (O_689,N_2900,N_4250);
nor UO_690 (O_690,N_3658,N_2903);
xnor UO_691 (O_691,N_3052,N_2734);
or UO_692 (O_692,N_4780,N_4572);
nand UO_693 (O_693,N_2706,N_3839);
or UO_694 (O_694,N_2602,N_3427);
or UO_695 (O_695,N_4082,N_2770);
xnor UO_696 (O_696,N_2607,N_4593);
and UO_697 (O_697,N_3285,N_2641);
and UO_698 (O_698,N_4022,N_3887);
and UO_699 (O_699,N_4053,N_3452);
xnor UO_700 (O_700,N_4866,N_3827);
xor UO_701 (O_701,N_3722,N_3889);
nand UO_702 (O_702,N_3669,N_4746);
xnor UO_703 (O_703,N_4883,N_3619);
or UO_704 (O_704,N_3469,N_4518);
and UO_705 (O_705,N_3677,N_4251);
xor UO_706 (O_706,N_3623,N_2968);
nor UO_707 (O_707,N_3520,N_2529);
or UO_708 (O_708,N_2690,N_3704);
nor UO_709 (O_709,N_4991,N_4904);
and UO_710 (O_710,N_3371,N_3878);
and UO_711 (O_711,N_3158,N_3861);
xnor UO_712 (O_712,N_3904,N_4828);
and UO_713 (O_713,N_3999,N_3816);
or UO_714 (O_714,N_4175,N_4943);
xnor UO_715 (O_715,N_2749,N_2753);
xnor UO_716 (O_716,N_4760,N_2797);
and UO_717 (O_717,N_4642,N_3033);
xnor UO_718 (O_718,N_3226,N_3879);
xor UO_719 (O_719,N_3729,N_3610);
nor UO_720 (O_720,N_3888,N_4308);
nor UO_721 (O_721,N_3265,N_4437);
nor UO_722 (O_722,N_4356,N_4027);
nand UO_723 (O_723,N_4534,N_3747);
nand UO_724 (O_724,N_4461,N_2718);
and UO_725 (O_725,N_4491,N_2762);
or UO_726 (O_726,N_3225,N_3792);
xnor UO_727 (O_727,N_4777,N_3522);
xnor UO_728 (O_728,N_3648,N_3341);
or UO_729 (O_729,N_4170,N_3267);
or UO_730 (O_730,N_3908,N_4422);
nor UO_731 (O_731,N_2776,N_2798);
nand UO_732 (O_732,N_4993,N_2580);
nor UO_733 (O_733,N_4410,N_4044);
nand UO_734 (O_734,N_3297,N_4517);
nor UO_735 (O_735,N_3871,N_4107);
or UO_736 (O_736,N_4338,N_3707);
nor UO_737 (O_737,N_3120,N_4902);
nand UO_738 (O_738,N_2614,N_2599);
or UO_739 (O_739,N_4072,N_4752);
and UO_740 (O_740,N_3231,N_3019);
xor UO_741 (O_741,N_4182,N_4602);
nand UO_742 (O_742,N_4228,N_2799);
nand UO_743 (O_743,N_3793,N_3365);
nor UO_744 (O_744,N_4245,N_4024);
and UO_745 (O_745,N_4078,N_4442);
nand UO_746 (O_746,N_3697,N_2585);
xnor UO_747 (O_747,N_4561,N_4342);
xor UO_748 (O_748,N_2594,N_3296);
xnor UO_749 (O_749,N_3604,N_4795);
or UO_750 (O_750,N_4443,N_3527);
and UO_751 (O_751,N_3039,N_3641);
nor UO_752 (O_752,N_3521,N_4468);
nor UO_753 (O_753,N_4928,N_4258);
nand UO_754 (O_754,N_4259,N_2665);
nand UO_755 (O_755,N_4050,N_4152);
nor UO_756 (O_756,N_4781,N_2563);
xnor UO_757 (O_757,N_3429,N_4948);
xor UO_758 (O_758,N_3573,N_2840);
or UO_759 (O_759,N_2732,N_4327);
and UO_760 (O_760,N_4353,N_4622);
nand UO_761 (O_761,N_2716,N_4847);
and UO_762 (O_762,N_4939,N_4039);
and UO_763 (O_763,N_3774,N_3045);
nand UO_764 (O_764,N_4774,N_4405);
xnor UO_765 (O_765,N_3327,N_3360);
nand UO_766 (O_766,N_3048,N_3948);
or UO_767 (O_767,N_3229,N_2567);
nor UO_768 (O_768,N_3679,N_2907);
or UO_769 (O_769,N_3086,N_4301);
xnor UO_770 (O_770,N_3651,N_3410);
nor UO_771 (O_771,N_2504,N_3160);
and UO_772 (O_772,N_4431,N_3703);
xnor UO_773 (O_773,N_4894,N_4503);
or UO_774 (O_774,N_3580,N_3963);
xor UO_775 (O_775,N_3763,N_2806);
nand UO_776 (O_776,N_3953,N_3544);
and UO_777 (O_777,N_3431,N_4036);
nor UO_778 (O_778,N_4151,N_3732);
nor UO_779 (O_779,N_3159,N_3003);
or UO_780 (O_780,N_3804,N_4524);
nor UO_781 (O_781,N_4697,N_2610);
nand UO_782 (O_782,N_3787,N_2620);
nor UO_783 (O_783,N_4859,N_2736);
and UO_784 (O_784,N_4463,N_3207);
xor UO_785 (O_785,N_2864,N_4355);
and UO_786 (O_786,N_4803,N_3000);
xnor UO_787 (O_787,N_3502,N_4931);
and UO_788 (O_788,N_3670,N_4563);
or UO_789 (O_789,N_2650,N_2937);
xnor UO_790 (O_790,N_4237,N_3760);
and UO_791 (O_791,N_4190,N_4424);
and UO_792 (O_792,N_4091,N_3603);
nand UO_793 (O_793,N_3664,N_3287);
and UO_794 (O_794,N_4398,N_4385);
and UO_795 (O_795,N_4853,N_3346);
xor UO_796 (O_796,N_3802,N_3405);
or UO_797 (O_797,N_3945,N_2860);
nor UO_798 (O_798,N_3442,N_4454);
xor UO_799 (O_799,N_3666,N_3770);
xor UO_800 (O_800,N_4911,N_2700);
or UO_801 (O_801,N_3489,N_4291);
and UO_802 (O_802,N_4048,N_2622);
or UO_803 (O_803,N_3053,N_3364);
or UO_804 (O_804,N_4681,N_2667);
nand UO_805 (O_805,N_4848,N_4615);
xor UO_806 (O_806,N_3386,N_3262);
xor UO_807 (O_807,N_4628,N_3504);
nor UO_808 (O_808,N_3552,N_3627);
nor UO_809 (O_809,N_4033,N_3592);
or UO_810 (O_810,N_3638,N_4744);
xor UO_811 (O_811,N_2830,N_3202);
or UO_812 (O_812,N_2985,N_3894);
nor UO_813 (O_813,N_3432,N_3087);
nor UO_814 (O_814,N_4229,N_4262);
and UO_815 (O_815,N_3657,N_3717);
nand UO_816 (O_816,N_4316,N_4054);
xnor UO_817 (O_817,N_3345,N_3284);
or UO_818 (O_818,N_3740,N_2823);
nand UO_819 (O_819,N_4014,N_4850);
or UO_820 (O_820,N_2619,N_3381);
or UO_821 (O_821,N_4544,N_3762);
and UO_822 (O_822,N_4568,N_4625);
xor UO_823 (O_823,N_4167,N_4672);
xnor UO_824 (O_824,N_4089,N_4827);
or UO_825 (O_825,N_3419,N_3477);
or UO_826 (O_826,N_2871,N_4988);
nand UO_827 (O_827,N_2960,N_3846);
or UO_828 (O_828,N_3865,N_4740);
and UO_829 (O_829,N_3922,N_4688);
or UO_830 (O_830,N_4539,N_2979);
and UO_831 (O_831,N_4492,N_2733);
or UO_832 (O_832,N_4814,N_4019);
nand UO_833 (O_833,N_3744,N_4791);
and UO_834 (O_834,N_4644,N_4924);
nand UO_835 (O_835,N_4557,N_4323);
or UO_836 (O_836,N_4372,N_3748);
xor UO_837 (O_837,N_4099,N_4234);
xor UO_838 (O_838,N_4313,N_3625);
or UO_839 (O_839,N_2789,N_4722);
or UO_840 (O_840,N_2891,N_2791);
nand UO_841 (O_841,N_3996,N_2991);
or UO_842 (O_842,N_4199,N_3730);
nor UO_843 (O_843,N_3594,N_3238);
nor UO_844 (O_844,N_3958,N_3814);
and UO_845 (O_845,N_3753,N_2575);
and UO_846 (O_846,N_2546,N_4765);
xor UO_847 (O_847,N_4530,N_2824);
and UO_848 (O_848,N_4080,N_2726);
nand UO_849 (O_849,N_3977,N_2946);
xnor UO_850 (O_850,N_3097,N_2792);
nor UO_851 (O_851,N_4055,N_3467);
nor UO_852 (O_852,N_4717,N_3842);
or UO_853 (O_853,N_4969,N_4956);
xor UO_854 (O_854,N_3940,N_2987);
or UO_855 (O_855,N_2595,N_2989);
and UO_856 (O_856,N_4035,N_2630);
or UO_857 (O_857,N_4857,N_4854);
and UO_858 (O_858,N_2702,N_3655);
or UO_859 (O_859,N_3301,N_3303);
xnor UO_860 (O_860,N_4161,N_4914);
xor UO_861 (O_861,N_4177,N_4012);
and UO_862 (O_862,N_4647,N_4295);
xnor UO_863 (O_863,N_3247,N_3082);
nand UO_864 (O_864,N_4178,N_4738);
nor UO_865 (O_865,N_2853,N_4264);
and UO_866 (O_866,N_3941,N_2746);
and UO_867 (O_867,N_3785,N_2874);
or UO_868 (O_868,N_4797,N_4073);
nand UO_869 (O_869,N_4440,N_3647);
nand UO_870 (O_870,N_4105,N_3085);
nand UO_871 (O_871,N_4281,N_3719);
xor UO_872 (O_872,N_4011,N_4368);
nor UO_873 (O_873,N_3302,N_4983);
nand UO_874 (O_874,N_3195,N_4891);
nand UO_875 (O_875,N_2941,N_3271);
nand UO_876 (O_876,N_3468,N_3328);
nor UO_877 (O_877,N_4830,N_4274);
nor UO_878 (O_878,N_4694,N_3423);
xor UO_879 (O_879,N_4706,N_2765);
nor UO_880 (O_880,N_2904,N_2520);
and UO_881 (O_881,N_2589,N_3236);
or UO_882 (O_882,N_4421,N_4173);
nor UO_883 (O_883,N_3910,N_3735);
xnor UO_884 (O_884,N_4606,N_4377);
and UO_885 (O_885,N_4773,N_3481);
or UO_886 (O_886,N_3126,N_3709);
nor UO_887 (O_887,N_3994,N_3368);
or UO_888 (O_888,N_3673,N_3388);
xnor UO_889 (O_889,N_4707,N_4111);
xnor UO_890 (O_890,N_4599,N_4556);
xnor UO_891 (O_891,N_3418,N_3805);
nor UO_892 (O_892,N_3672,N_4624);
and UO_893 (O_893,N_3523,N_3358);
nor UO_894 (O_894,N_4870,N_3250);
xnor UO_895 (O_895,N_3893,N_2701);
xnor UO_896 (O_896,N_4449,N_4989);
and UO_897 (O_897,N_3868,N_4284);
or UO_898 (O_898,N_3443,N_2828);
or UO_899 (O_899,N_3110,N_2638);
nand UO_900 (O_900,N_3413,N_3924);
and UO_901 (O_901,N_3694,N_3069);
or UO_902 (O_902,N_3646,N_3781);
xor UO_903 (O_903,N_3430,N_4090);
nand UO_904 (O_904,N_4633,N_3128);
or UO_905 (O_905,N_3408,N_3584);
nand UO_906 (O_906,N_4839,N_2548);
xor UO_907 (O_907,N_4718,N_3425);
xor UO_908 (O_908,N_4950,N_4134);
nor UO_909 (O_909,N_3972,N_4457);
xnor UO_910 (O_910,N_2898,N_3367);
nand UO_911 (O_911,N_4588,N_4657);
nand UO_912 (O_912,N_2892,N_2752);
nor UO_913 (O_913,N_4471,N_3268);
nand UO_914 (O_914,N_4084,N_3855);
or UO_915 (O_915,N_4280,N_3833);
xnor UO_916 (O_916,N_3444,N_3458);
and UO_917 (O_917,N_4684,N_3608);
or UO_918 (O_918,N_4333,N_2877);
nor UO_919 (O_919,N_3812,N_4811);
or UO_920 (O_920,N_3554,N_4808);
or UO_921 (O_921,N_4231,N_3136);
nand UO_922 (O_922,N_4558,N_2963);
xnor UO_923 (O_923,N_3403,N_2654);
xor UO_924 (O_924,N_4184,N_3797);
and UO_925 (O_925,N_2952,N_4314);
nor UO_926 (O_926,N_4586,N_2811);
nand UO_927 (O_927,N_4650,N_3460);
xor UO_928 (O_928,N_2804,N_2944);
xnor UO_929 (O_929,N_3970,N_4227);
and UO_930 (O_930,N_4490,N_2648);
or UO_931 (O_931,N_3066,N_3228);
xor UO_932 (O_932,N_3182,N_4276);
and UO_933 (O_933,N_2847,N_2744);
nand UO_934 (O_934,N_3062,N_4318);
xor UO_935 (O_935,N_4614,N_2793);
xnor UO_936 (O_936,N_4260,N_4630);
nand UO_937 (O_937,N_4535,N_3406);
or UO_938 (O_938,N_4899,N_2705);
nand UO_939 (O_939,N_3725,N_3329);
nand UO_940 (O_940,N_2870,N_3375);
xnor UO_941 (O_941,N_4809,N_4741);
nor UO_942 (O_942,N_4429,N_3040);
nor UO_943 (O_943,N_4507,N_3883);
and UO_944 (O_944,N_3665,N_3643);
xnor UO_945 (O_945,N_4753,N_3836);
xor UO_946 (O_946,N_2535,N_2569);
xor UO_947 (O_947,N_3892,N_3433);
and UO_948 (O_948,N_4263,N_4017);
xnor UO_949 (O_949,N_3791,N_2873);
and UO_950 (O_950,N_4298,N_2578);
and UO_951 (O_951,N_4715,N_3928);
nor UO_952 (O_952,N_4798,N_4362);
nand UO_953 (O_953,N_3689,N_4978);
and UO_954 (O_954,N_2872,N_2689);
nand UO_955 (O_955,N_2552,N_4985);
xor UO_956 (O_956,N_4999,N_3545);
or UO_957 (O_957,N_4682,N_3035);
xor UO_958 (O_958,N_2836,N_2818);
xnor UO_959 (O_959,N_3269,N_3711);
and UO_960 (O_960,N_3750,N_3266);
and UO_961 (O_961,N_3076,N_4520);
and UO_962 (O_962,N_3606,N_2997);
and UO_963 (O_963,N_4448,N_2685);
or UO_964 (O_964,N_4201,N_4766);
nand UO_965 (O_965,N_3455,N_3809);
or UO_966 (O_966,N_3292,N_4772);
and UO_967 (O_967,N_4241,N_2802);
and UO_968 (O_968,N_3695,N_4702);
nand UO_969 (O_969,N_2507,N_3613);
and UO_970 (O_970,N_3283,N_3324);
nand UO_971 (O_971,N_3361,N_3726);
xnor UO_972 (O_972,N_3099,N_3007);
nor UO_973 (O_973,N_3293,N_4502);
nand UO_974 (O_974,N_4337,N_2621);
nand UO_975 (O_975,N_4128,N_4240);
nor UO_976 (O_976,N_4397,N_3070);
or UO_977 (O_977,N_3685,N_4129);
xnor UO_978 (O_978,N_3058,N_4057);
nand UO_979 (O_979,N_4489,N_3775);
xnor UO_980 (O_980,N_3192,N_3915);
and UO_981 (O_981,N_3706,N_4869);
and UO_982 (O_982,N_3307,N_2522);
nor UO_983 (O_983,N_4074,N_2759);
nor UO_984 (O_984,N_3659,N_4737);
and UO_985 (O_985,N_2777,N_3321);
or UO_986 (O_986,N_2902,N_3609);
or UO_987 (O_987,N_2924,N_4217);
nor UO_988 (O_988,N_4126,N_3004);
nor UO_989 (O_989,N_3032,N_3778);
and UO_990 (O_990,N_4768,N_4069);
and UO_991 (O_991,N_4788,N_4879);
and UO_992 (O_992,N_4324,N_2659);
and UO_993 (O_993,N_3650,N_2592);
xnor UO_994 (O_994,N_4860,N_4093);
and UO_995 (O_995,N_3482,N_3174);
xnor UO_996 (O_996,N_4559,N_4433);
or UO_997 (O_997,N_3134,N_3370);
or UO_998 (O_998,N_4907,N_2608);
and UO_999 (O_999,N_4910,N_2889);
endmodule