module basic_1000_10000_1500_10_levels_1xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_293,In_617);
and U1 (N_1,In_867,In_553);
or U2 (N_2,In_728,In_564);
or U3 (N_3,In_840,In_118);
or U4 (N_4,In_628,In_649);
nor U5 (N_5,In_490,In_813);
and U6 (N_6,In_53,In_644);
or U7 (N_7,In_292,In_541);
nor U8 (N_8,In_909,In_522);
nor U9 (N_9,In_47,In_52);
nor U10 (N_10,In_991,In_414);
and U11 (N_11,In_876,In_161);
nor U12 (N_12,In_401,In_784);
and U13 (N_13,In_800,In_589);
nor U14 (N_14,In_865,In_86);
nor U15 (N_15,In_45,In_312);
and U16 (N_16,In_910,In_382);
nand U17 (N_17,In_677,In_939);
nand U18 (N_18,In_925,In_374);
or U19 (N_19,In_466,In_605);
or U20 (N_20,In_378,In_363);
nor U21 (N_21,In_210,In_237);
or U22 (N_22,In_282,In_569);
and U23 (N_23,In_445,In_127);
and U24 (N_24,In_64,In_600);
or U25 (N_25,In_744,In_970);
nor U26 (N_26,In_60,In_413);
nand U27 (N_27,In_188,In_333);
and U28 (N_28,In_460,In_380);
or U29 (N_29,In_701,In_219);
or U30 (N_30,In_325,In_354);
and U31 (N_31,In_515,In_969);
nor U32 (N_32,In_906,In_448);
nand U33 (N_33,In_789,In_355);
and U34 (N_34,In_83,In_781);
and U35 (N_35,In_443,In_560);
nand U36 (N_36,In_27,In_262);
nor U37 (N_37,In_539,In_832);
and U38 (N_38,In_25,In_624);
xnor U39 (N_39,In_533,In_598);
nor U40 (N_40,In_159,In_62);
nand U41 (N_41,In_544,In_16);
or U42 (N_42,In_635,In_756);
or U43 (N_43,In_696,In_556);
and U44 (N_44,In_698,In_362);
nor U45 (N_45,In_69,In_441);
and U46 (N_46,In_552,In_904);
and U47 (N_47,In_493,In_622);
nand U48 (N_48,In_810,In_695);
nor U49 (N_49,In_654,In_120);
nor U50 (N_50,In_152,In_202);
nand U51 (N_51,In_599,In_97);
or U52 (N_52,In_452,In_594);
and U53 (N_53,In_924,In_46);
nor U54 (N_54,In_176,In_956);
nor U55 (N_55,In_863,In_754);
or U56 (N_56,In_128,In_835);
nor U57 (N_57,In_763,In_423);
or U58 (N_58,In_418,In_108);
nor U59 (N_59,In_146,In_839);
and U60 (N_60,In_726,In_997);
xnor U61 (N_61,In_618,In_36);
nor U62 (N_62,In_203,In_211);
or U63 (N_63,In_171,In_933);
nor U64 (N_64,In_962,In_399);
nor U65 (N_65,In_735,In_430);
nand U66 (N_66,In_106,In_667);
nand U67 (N_67,In_186,In_115);
and U68 (N_68,In_940,In_65);
nand U69 (N_69,In_982,In_191);
or U70 (N_70,In_602,In_737);
nor U71 (N_71,In_929,In_75);
and U72 (N_72,In_145,In_234);
or U73 (N_73,In_243,In_782);
nand U74 (N_74,In_139,In_995);
nor U75 (N_75,In_137,In_240);
nor U76 (N_76,In_93,In_897);
nor U77 (N_77,In_946,In_3);
and U78 (N_78,In_314,In_932);
and U79 (N_79,In_10,In_536);
and U80 (N_80,In_623,In_576);
and U81 (N_81,In_257,In_558);
and U82 (N_82,In_117,In_831);
and U83 (N_83,In_548,In_579);
nand U84 (N_84,In_542,In_738);
nor U85 (N_85,In_793,In_361);
and U86 (N_86,In_266,In_410);
and U87 (N_87,In_678,In_196);
or U88 (N_88,In_141,In_583);
and U89 (N_89,In_439,In_705);
nand U90 (N_90,In_389,In_388);
nand U91 (N_91,In_534,In_577);
xnor U92 (N_92,In_893,In_258);
nor U93 (N_93,In_862,In_421);
or U94 (N_94,In_952,In_947);
or U95 (N_95,In_37,In_222);
and U96 (N_96,In_755,In_487);
or U97 (N_97,In_442,In_926);
nand U98 (N_98,In_658,In_456);
or U99 (N_99,In_309,In_360);
or U100 (N_100,In_974,In_177);
nor U101 (N_101,In_61,In_422);
nor U102 (N_102,In_149,In_209);
nand U103 (N_103,In_261,In_565);
and U104 (N_104,In_610,In_281);
or U105 (N_105,In_400,In_291);
nand U106 (N_106,In_223,In_693);
nor U107 (N_107,In_778,In_464);
and U108 (N_108,In_918,In_406);
nor U109 (N_109,In_265,In_129);
or U110 (N_110,In_836,In_160);
nand U111 (N_111,In_285,In_734);
nand U112 (N_112,In_31,In_263);
nand U113 (N_113,In_514,In_878);
nor U114 (N_114,In_516,In_773);
nand U115 (N_115,In_271,In_408);
nor U116 (N_116,In_71,In_531);
nand U117 (N_117,In_59,In_471);
and U118 (N_118,In_297,In_339);
or U119 (N_119,In_168,In_777);
nor U120 (N_120,In_32,In_581);
nor U121 (N_121,In_767,In_409);
nand U122 (N_122,In_669,In_978);
and U123 (N_123,In_283,In_627);
or U124 (N_124,In_397,In_747);
nor U125 (N_125,In_686,In_395);
or U126 (N_126,In_608,In_670);
nor U127 (N_127,In_84,In_461);
nor U128 (N_128,In_869,In_329);
nand U129 (N_129,In_807,In_509);
nand U130 (N_130,In_647,In_819);
nor U131 (N_131,In_379,In_742);
or U132 (N_132,In_157,In_603);
or U133 (N_133,In_462,In_525);
xor U134 (N_134,In_614,In_943);
nand U135 (N_135,In_275,In_692);
nor U136 (N_136,In_711,In_844);
and U137 (N_137,In_934,In_167);
and U138 (N_138,In_340,In_561);
nor U139 (N_139,In_975,In_759);
nand U140 (N_140,In_967,In_130);
and U141 (N_141,In_226,In_923);
and U142 (N_142,In_444,In_426);
or U143 (N_143,In_214,In_690);
nor U144 (N_144,In_620,In_402);
or U145 (N_145,In_597,In_290);
or U146 (N_146,In_529,In_310);
or U147 (N_147,In_775,In_392);
nor U148 (N_148,In_963,In_135);
and U149 (N_149,In_357,In_0);
and U150 (N_150,In_125,In_899);
and U151 (N_151,In_621,In_829);
nor U152 (N_152,In_197,In_304);
nor U153 (N_153,In_50,In_900);
and U154 (N_154,In_609,In_142);
nor U155 (N_155,In_945,In_676);
and U156 (N_156,In_748,In_496);
or U157 (N_157,In_364,In_371);
nor U158 (N_158,In_668,In_110);
and U159 (N_159,In_791,In_732);
and U160 (N_160,In_858,In_51);
nor U161 (N_161,In_871,In_868);
nand U162 (N_162,In_350,In_313);
nand U163 (N_163,In_903,In_804);
and U164 (N_164,In_733,In_834);
nor U165 (N_165,In_109,In_156);
and U166 (N_166,In_198,In_774);
nand U167 (N_167,In_592,In_163);
or U168 (N_168,In_739,In_985);
or U169 (N_169,In_316,In_227);
or U170 (N_170,In_495,In_301);
nor U171 (N_171,In_342,In_42);
or U172 (N_172,In_207,In_749);
nor U173 (N_173,In_625,In_450);
or U174 (N_174,In_231,In_429);
or U175 (N_175,In_102,In_555);
or U176 (N_176,In_540,In_331);
and U177 (N_177,In_381,In_545);
or U178 (N_178,In_612,In_817);
nor U179 (N_179,In_914,In_386);
nor U180 (N_180,In_626,In_74);
nand U181 (N_181,In_870,In_845);
nor U182 (N_182,In_478,In_849);
nor U183 (N_183,In_15,In_131);
nand U184 (N_184,In_475,In_172);
nand U185 (N_185,In_930,In_937);
and U186 (N_186,In_76,In_327);
nor U187 (N_187,In_730,In_228);
nor U188 (N_188,In_242,In_277);
nor U189 (N_189,In_48,In_886);
or U190 (N_190,In_827,In_498);
nand U191 (N_191,In_124,In_526);
or U192 (N_192,In_185,In_528);
nor U193 (N_193,In_861,In_595);
or U194 (N_194,In_665,In_562);
or U195 (N_195,In_935,In_916);
or U196 (N_196,In_494,In_786);
or U197 (N_197,In_499,In_586);
or U198 (N_198,In_416,In_335);
nor U199 (N_199,In_57,In_814);
and U200 (N_200,In_484,In_472);
or U201 (N_201,In_806,In_317);
nor U202 (N_202,In_492,In_994);
nand U203 (N_203,In_305,In_680);
and U204 (N_204,In_879,In_745);
or U205 (N_205,In_613,In_255);
nor U206 (N_206,In_259,In_403);
nand U207 (N_207,In_353,In_717);
nor U208 (N_208,In_640,In_768);
or U209 (N_209,In_706,In_104);
and U210 (N_210,In_841,In_384);
and U211 (N_211,In_999,In_979);
and U212 (N_212,In_532,In_746);
nor U213 (N_213,In_769,In_44);
nand U214 (N_214,In_811,In_891);
and U215 (N_215,In_855,In_770);
xnor U216 (N_216,In_713,In_289);
and U217 (N_217,In_675,In_238);
nand U218 (N_218,In_771,In_85);
nor U219 (N_219,In_828,In_17);
nor U220 (N_220,In_981,In_761);
nand U221 (N_221,In_465,In_480);
and U222 (N_222,In_479,In_885);
or U223 (N_223,In_467,In_998);
or U224 (N_224,In_303,In_294);
xnor U225 (N_225,In_311,In_977);
nand U226 (N_226,In_474,In_296);
nor U227 (N_227,In_537,In_356);
nor U228 (N_228,In_966,In_77);
nand U229 (N_229,In_323,In_92);
nand U230 (N_230,In_366,In_941);
nor U231 (N_231,In_107,In_567);
nor U232 (N_232,In_319,In_425);
nor U233 (N_233,In_741,In_679);
and U234 (N_234,In_375,In_489);
nor U235 (N_235,In_919,In_182);
or U236 (N_236,In_368,In_708);
nand U237 (N_237,In_349,In_136);
nor U238 (N_238,In_189,In_992);
nor U239 (N_239,In_477,In_411);
nand U240 (N_240,In_387,In_35);
or U241 (N_241,In_961,In_760);
or U242 (N_242,In_41,In_417);
and U243 (N_243,In_229,In_587);
nor U244 (N_244,In_87,In_795);
or U245 (N_245,In_954,In_121);
or U246 (N_246,In_653,In_779);
nand U247 (N_247,In_434,In_950);
nor U248 (N_248,In_43,In_500);
and U249 (N_249,In_113,In_199);
nand U250 (N_250,In_476,In_220);
nand U251 (N_251,In_549,In_905);
nand U252 (N_252,In_269,In_601);
xnor U253 (N_253,In_812,In_272);
and U254 (N_254,In_527,In_816);
nor U255 (N_255,In_607,In_138);
and U256 (N_256,In_968,In_568);
nand U257 (N_257,In_896,In_436);
nand U258 (N_258,In_24,In_922);
nor U259 (N_259,In_632,In_112);
or U260 (N_260,In_345,In_184);
or U261 (N_261,In_236,In_547);
nor U262 (N_262,In_169,In_641);
nand U263 (N_263,In_502,In_661);
and U264 (N_264,In_78,In_405);
nand U265 (N_265,In_765,In_433);
nand U266 (N_266,In_630,In_302);
nand U267 (N_267,In_100,In_799);
nand U268 (N_268,In_797,In_338);
and U269 (N_269,In_902,In_508);
or U270 (N_270,In_344,In_246);
or U271 (N_271,In_13,In_287);
nor U272 (N_272,In_268,In_758);
or U273 (N_273,In_235,In_481);
nand U274 (N_274,In_6,In_221);
and U275 (N_275,In_723,In_88);
or U276 (N_276,In_279,In_650);
and U277 (N_277,In_151,In_873);
or U278 (N_278,In_582,In_501);
nor U279 (N_279,In_491,In_79);
nor U280 (N_280,In_611,In_521);
nor U281 (N_281,In_651,In_63);
and U282 (N_282,In_288,In_833);
or U283 (N_283,In_91,In_751);
and U284 (N_284,In_419,In_306);
nand U285 (N_285,In_672,In_574);
nand U286 (N_286,In_38,In_396);
and U287 (N_287,In_762,In_857);
nand U288 (N_288,In_173,In_822);
and U289 (N_289,In_449,In_123);
nand U290 (N_290,In_4,In_116);
nor U291 (N_291,In_206,In_95);
nor U292 (N_292,In_81,In_883);
and U293 (N_293,In_18,In_82);
or U294 (N_294,In_11,In_394);
nor U295 (N_295,In_854,In_359);
or U296 (N_296,In_267,In_575);
nor U297 (N_297,In_321,In_105);
nor U298 (N_298,In_927,In_133);
nand U299 (N_299,In_913,In_504);
nand U300 (N_300,In_615,In_720);
nand U301 (N_301,In_792,In_270);
or U302 (N_302,In_468,In_944);
and U303 (N_303,In_94,In_119);
or U304 (N_304,In_964,In_34);
nor U305 (N_305,In_393,In_346);
nor U306 (N_306,In_390,In_908);
and U307 (N_307,In_566,In_239);
or U308 (N_308,In_90,In_593);
nand U309 (N_309,In_699,In_253);
xnor U310 (N_310,In_830,In_874);
and U311 (N_311,In_218,In_358);
nor U312 (N_312,In_629,In_546);
nand U313 (N_313,In_54,In_164);
nand U314 (N_314,In_636,In_326);
nand U315 (N_315,In_457,In_158);
or U316 (N_316,In_300,In_570);
nand U317 (N_317,In_482,In_217);
or U318 (N_318,In_451,In_681);
nand U319 (N_319,In_40,In_469);
nor U320 (N_320,In_510,In_590);
nand U321 (N_321,In_483,In_215);
or U322 (N_322,In_702,In_420);
and U323 (N_323,In_73,In_39);
and U324 (N_324,In_122,In_685);
nor U325 (N_325,In_972,In_192);
and U326 (N_326,In_634,In_488);
and U327 (N_327,In_459,In_264);
xnor U328 (N_328,In_783,In_30);
nor U329 (N_329,In_260,In_704);
nor U330 (N_330,In_703,In_497);
nor U331 (N_331,In_660,In_148);
nor U332 (N_332,In_5,In_183);
xnor U333 (N_333,In_66,In_14);
nand U334 (N_334,In_274,In_524);
nor U335 (N_335,In_225,In_803);
or U336 (N_336,In_233,In_67);
xnor U337 (N_337,In_820,In_864);
nand U338 (N_338,In_398,In_664);
and U339 (N_339,In_330,In_557);
nor U340 (N_340,In_385,In_463);
nor U341 (N_341,In_616,In_788);
or U342 (N_342,In_241,In_951);
nor U343 (N_343,In_458,In_798);
and U344 (N_344,In_373,In_376);
nand U345 (N_345,In_26,In_689);
nand U346 (N_346,In_752,In_193);
nand U347 (N_347,In_980,In_538);
nand U348 (N_348,In_727,In_805);
nor U349 (N_349,In_716,In_996);
or U350 (N_350,In_147,In_881);
or U351 (N_351,In_697,In_837);
or U352 (N_352,In_101,In_989);
and U353 (N_353,In_165,In_652);
nand U354 (N_354,In_959,In_446);
and U355 (N_355,In_518,In_9);
nor U356 (N_356,In_986,In_72);
nor U357 (N_357,In_308,In_729);
or U358 (N_358,In_983,In_298);
nor U359 (N_359,In_20,In_520);
and U360 (N_360,In_990,In_875);
or U361 (N_361,In_580,In_440);
or U362 (N_362,In_8,In_573);
nand U363 (N_363,In_7,In_852);
or U364 (N_364,In_725,In_843);
nand U365 (N_365,In_960,In_334);
and U366 (N_366,In_470,In_993);
nor U367 (N_367,In_190,In_688);
nand U368 (N_368,In_780,In_889);
nand U369 (N_369,In_332,In_80);
nor U370 (N_370,In_322,In_432);
nand U371 (N_371,In_656,In_796);
nor U372 (N_372,In_352,In_888);
or U373 (N_373,In_642,In_847);
nand U374 (N_374,In_776,In_68);
or U375 (N_375,In_764,In_958);
nand U376 (N_376,In_588,In_682);
or U377 (N_377,In_415,In_49);
nand U378 (N_378,In_825,In_412);
or U379 (N_379,In_637,In_866);
nor U380 (N_380,In_507,In_787);
or U381 (N_381,In_216,In_766);
and U382 (N_382,In_424,In_872);
or U383 (N_383,In_324,In_153);
or U384 (N_384,In_683,In_709);
and U385 (N_385,In_743,In_427);
or U386 (N_386,In_802,In_377);
or U387 (N_387,In_824,In_250);
and U388 (N_388,In_638,In_585);
nand U389 (N_389,In_848,In_180);
and U390 (N_390,In_920,In_99);
nor U391 (N_391,In_860,In_794);
nand U392 (N_392,In_150,In_56);
and U393 (N_393,In_691,In_643);
nand U394 (N_394,In_284,In_174);
or U395 (N_395,In_687,In_965);
and U396 (N_396,In_299,In_140);
nor U397 (N_397,In_208,In_256);
or U398 (N_398,In_367,In_821);
or U399 (N_399,In_971,In_563);
and U400 (N_400,In_645,In_513);
nor U401 (N_401,In_204,In_249);
nor U402 (N_402,In_245,In_984);
nand U403 (N_403,In_921,In_273);
nor U404 (N_404,In_365,In_280);
nand U405 (N_405,In_278,In_659);
nor U406 (N_406,In_205,In_372);
nand U407 (N_407,In_949,In_486);
or U408 (N_408,In_200,In_724);
nand U409 (N_409,In_276,In_604);
and U410 (N_410,In_631,In_2);
and U411 (N_411,In_347,In_503);
and U412 (N_412,In_719,In_596);
nand U413 (N_413,In_315,In_407);
nor U414 (N_414,In_619,In_251);
nor U415 (N_415,In_58,In_166);
and U416 (N_416,In_838,In_431);
and U417 (N_417,In_815,In_254);
nand U418 (N_418,In_987,In_114);
or U419 (N_419,In_790,In_224);
nor U420 (N_420,In_884,In_715);
and U421 (N_421,In_428,In_955);
and U422 (N_422,In_391,In_320);
and U423 (N_423,In_912,In_181);
nor U424 (N_424,In_383,In_21);
and U425 (N_425,In_1,In_170);
nor U426 (N_426,In_447,In_195);
nor U427 (N_427,In_646,In_530);
or U428 (N_428,In_307,In_559);
and U429 (N_429,In_895,In_132);
nor U430 (N_430,In_712,In_936);
and U431 (N_431,In_19,In_907);
nor U432 (N_432,In_808,In_584);
and U433 (N_433,In_571,In_673);
nand U434 (N_434,In_230,In_694);
or U435 (N_435,In_882,In_212);
or U436 (N_436,In_370,In_684);
nor U437 (N_437,In_901,In_785);
nor U438 (N_438,In_674,In_12);
or U439 (N_439,In_853,In_578);
and U440 (N_440,In_519,In_942);
and U441 (N_441,In_714,In_194);
and U442 (N_442,In_33,In_155);
nor U443 (N_443,In_337,In_823);
and U444 (N_444,In_55,In_454);
and U445 (N_445,In_740,In_973);
nor U446 (N_446,In_328,In_455);
and U447 (N_447,In_134,In_655);
nor U448 (N_448,In_898,In_473);
and U449 (N_449,In_517,In_554);
and U450 (N_450,In_666,In_976);
nor U451 (N_451,In_736,In_178);
nand U452 (N_452,In_126,In_809);
nor U453 (N_453,In_437,In_505);
nor U454 (N_454,In_369,In_22);
nor U455 (N_455,In_232,In_850);
nor U456 (N_456,In_404,In_957);
nor U457 (N_457,In_928,In_890);
or U458 (N_458,In_931,In_948);
or U459 (N_459,In_144,In_648);
nor U460 (N_460,In_591,In_248);
nor U461 (N_461,In_818,In_154);
or U462 (N_462,In_856,In_721);
nand U463 (N_463,In_606,In_103);
nor U464 (N_464,In_213,In_318);
nand U465 (N_465,In_911,In_523);
nor U466 (N_466,In_718,In_750);
nor U467 (N_467,In_143,In_295);
or U468 (N_468,In_753,In_826);
xor U469 (N_469,In_535,In_252);
nor U470 (N_470,In_663,In_187);
or U471 (N_471,In_700,In_550);
or U472 (N_472,In_96,In_731);
nor U473 (N_473,In_453,In_572);
and U474 (N_474,In_772,In_70);
or U475 (N_475,In_201,In_162);
and U476 (N_476,In_551,In_89);
nand U477 (N_477,In_707,In_543);
nor U478 (N_478,In_842,In_846);
xnor U479 (N_479,In_28,In_722);
nor U480 (N_480,In_657,In_343);
nor U481 (N_481,In_894,In_988);
nand U482 (N_482,In_179,In_348);
and U483 (N_483,In_98,In_953);
and U484 (N_484,In_351,In_633);
nand U485 (N_485,In_286,In_880);
nor U486 (N_486,In_801,In_917);
nand U487 (N_487,In_757,In_851);
nand U488 (N_488,In_671,In_938);
and U489 (N_489,In_662,In_438);
and U490 (N_490,In_244,In_710);
or U491 (N_491,In_341,In_336);
and U492 (N_492,In_512,In_506);
and U493 (N_493,In_511,In_915);
nor U494 (N_494,In_887,In_435);
nand U495 (N_495,In_859,In_892);
nand U496 (N_496,In_111,In_29);
and U497 (N_497,In_639,In_247);
and U498 (N_498,In_877,In_175);
nand U499 (N_499,In_23,In_485);
nand U500 (N_500,In_168,In_317);
and U501 (N_501,In_455,In_547);
or U502 (N_502,In_610,In_379);
nand U503 (N_503,In_393,In_484);
and U504 (N_504,In_398,In_38);
and U505 (N_505,In_886,In_993);
nor U506 (N_506,In_759,In_797);
nand U507 (N_507,In_395,In_155);
nand U508 (N_508,In_806,In_613);
nand U509 (N_509,In_374,In_157);
nor U510 (N_510,In_888,In_96);
nor U511 (N_511,In_115,In_654);
nand U512 (N_512,In_126,In_949);
nor U513 (N_513,In_839,In_811);
nand U514 (N_514,In_360,In_688);
and U515 (N_515,In_406,In_168);
and U516 (N_516,In_366,In_49);
and U517 (N_517,In_771,In_351);
nand U518 (N_518,In_252,In_606);
or U519 (N_519,In_381,In_674);
and U520 (N_520,In_659,In_384);
nor U521 (N_521,In_899,In_748);
and U522 (N_522,In_836,In_497);
nor U523 (N_523,In_834,In_340);
or U524 (N_524,In_773,In_892);
and U525 (N_525,In_627,In_180);
and U526 (N_526,In_848,In_348);
or U527 (N_527,In_330,In_649);
and U528 (N_528,In_451,In_148);
and U529 (N_529,In_202,In_642);
or U530 (N_530,In_279,In_589);
nor U531 (N_531,In_785,In_386);
nor U532 (N_532,In_996,In_984);
nor U533 (N_533,In_926,In_418);
nor U534 (N_534,In_431,In_432);
or U535 (N_535,In_886,In_252);
nor U536 (N_536,In_835,In_700);
or U537 (N_537,In_835,In_247);
or U538 (N_538,In_333,In_626);
nor U539 (N_539,In_704,In_130);
nor U540 (N_540,In_997,In_812);
or U541 (N_541,In_687,In_372);
nand U542 (N_542,In_684,In_310);
or U543 (N_543,In_601,In_772);
nand U544 (N_544,In_551,In_930);
nand U545 (N_545,In_333,In_273);
and U546 (N_546,In_894,In_475);
and U547 (N_547,In_567,In_677);
nand U548 (N_548,In_621,In_38);
and U549 (N_549,In_536,In_914);
nand U550 (N_550,In_987,In_118);
nor U551 (N_551,In_177,In_87);
and U552 (N_552,In_344,In_219);
nor U553 (N_553,In_292,In_670);
nand U554 (N_554,In_338,In_763);
nand U555 (N_555,In_300,In_295);
and U556 (N_556,In_292,In_901);
nand U557 (N_557,In_449,In_953);
and U558 (N_558,In_703,In_485);
nand U559 (N_559,In_961,In_954);
and U560 (N_560,In_622,In_149);
and U561 (N_561,In_936,In_952);
or U562 (N_562,In_442,In_846);
nor U563 (N_563,In_332,In_692);
and U564 (N_564,In_600,In_537);
or U565 (N_565,In_58,In_168);
nand U566 (N_566,In_529,In_85);
nor U567 (N_567,In_519,In_135);
and U568 (N_568,In_322,In_529);
nand U569 (N_569,In_278,In_218);
nor U570 (N_570,In_718,In_228);
or U571 (N_571,In_376,In_515);
or U572 (N_572,In_289,In_909);
nand U573 (N_573,In_322,In_487);
and U574 (N_574,In_524,In_112);
nand U575 (N_575,In_737,In_575);
or U576 (N_576,In_681,In_118);
or U577 (N_577,In_129,In_555);
or U578 (N_578,In_615,In_246);
and U579 (N_579,In_700,In_825);
or U580 (N_580,In_213,In_803);
nor U581 (N_581,In_430,In_531);
nand U582 (N_582,In_781,In_775);
nand U583 (N_583,In_478,In_247);
and U584 (N_584,In_606,In_759);
and U585 (N_585,In_728,In_744);
nand U586 (N_586,In_856,In_243);
nand U587 (N_587,In_38,In_980);
nand U588 (N_588,In_681,In_265);
nand U589 (N_589,In_740,In_918);
and U590 (N_590,In_836,In_257);
or U591 (N_591,In_946,In_580);
nand U592 (N_592,In_264,In_652);
and U593 (N_593,In_66,In_201);
xnor U594 (N_594,In_305,In_942);
nand U595 (N_595,In_359,In_677);
nand U596 (N_596,In_881,In_830);
nor U597 (N_597,In_156,In_206);
nand U598 (N_598,In_82,In_785);
nand U599 (N_599,In_568,In_297);
nor U600 (N_600,In_959,In_60);
and U601 (N_601,In_794,In_658);
or U602 (N_602,In_720,In_11);
nand U603 (N_603,In_866,In_652);
nand U604 (N_604,In_113,In_798);
nand U605 (N_605,In_793,In_348);
nand U606 (N_606,In_444,In_772);
and U607 (N_607,In_249,In_172);
nand U608 (N_608,In_715,In_50);
and U609 (N_609,In_680,In_426);
and U610 (N_610,In_98,In_289);
nor U611 (N_611,In_23,In_136);
nor U612 (N_612,In_271,In_546);
nor U613 (N_613,In_589,In_372);
or U614 (N_614,In_699,In_364);
and U615 (N_615,In_479,In_803);
and U616 (N_616,In_335,In_178);
or U617 (N_617,In_489,In_920);
nand U618 (N_618,In_152,In_963);
nor U619 (N_619,In_604,In_51);
nand U620 (N_620,In_308,In_447);
nand U621 (N_621,In_553,In_552);
and U622 (N_622,In_382,In_889);
or U623 (N_623,In_575,In_783);
and U624 (N_624,In_99,In_973);
nor U625 (N_625,In_916,In_366);
or U626 (N_626,In_745,In_83);
nor U627 (N_627,In_723,In_439);
and U628 (N_628,In_839,In_85);
or U629 (N_629,In_981,In_341);
and U630 (N_630,In_60,In_675);
nor U631 (N_631,In_706,In_586);
or U632 (N_632,In_575,In_858);
nand U633 (N_633,In_820,In_263);
and U634 (N_634,In_291,In_585);
nor U635 (N_635,In_154,In_712);
nor U636 (N_636,In_41,In_309);
nor U637 (N_637,In_710,In_679);
or U638 (N_638,In_229,In_92);
and U639 (N_639,In_543,In_388);
or U640 (N_640,In_505,In_438);
or U641 (N_641,In_777,In_514);
or U642 (N_642,In_506,In_20);
and U643 (N_643,In_735,In_608);
or U644 (N_644,In_506,In_827);
nor U645 (N_645,In_505,In_119);
nor U646 (N_646,In_555,In_261);
nor U647 (N_647,In_782,In_661);
and U648 (N_648,In_780,In_397);
and U649 (N_649,In_826,In_77);
or U650 (N_650,In_283,In_976);
or U651 (N_651,In_500,In_834);
nor U652 (N_652,In_242,In_337);
nor U653 (N_653,In_850,In_805);
or U654 (N_654,In_976,In_129);
nor U655 (N_655,In_368,In_179);
or U656 (N_656,In_150,In_927);
and U657 (N_657,In_506,In_184);
or U658 (N_658,In_315,In_311);
and U659 (N_659,In_546,In_568);
nand U660 (N_660,In_709,In_729);
and U661 (N_661,In_321,In_630);
and U662 (N_662,In_73,In_704);
or U663 (N_663,In_395,In_674);
or U664 (N_664,In_106,In_531);
nor U665 (N_665,In_289,In_646);
and U666 (N_666,In_361,In_722);
and U667 (N_667,In_351,In_399);
nand U668 (N_668,In_312,In_831);
or U669 (N_669,In_652,In_198);
nand U670 (N_670,In_273,In_764);
nand U671 (N_671,In_143,In_316);
and U672 (N_672,In_631,In_466);
xor U673 (N_673,In_773,In_814);
or U674 (N_674,In_567,In_933);
or U675 (N_675,In_293,In_452);
and U676 (N_676,In_568,In_435);
nor U677 (N_677,In_276,In_315);
nor U678 (N_678,In_514,In_281);
nand U679 (N_679,In_704,In_682);
or U680 (N_680,In_294,In_364);
and U681 (N_681,In_209,In_376);
and U682 (N_682,In_547,In_38);
nand U683 (N_683,In_634,In_394);
and U684 (N_684,In_633,In_941);
nand U685 (N_685,In_438,In_761);
nand U686 (N_686,In_660,In_879);
or U687 (N_687,In_969,In_718);
nor U688 (N_688,In_293,In_201);
or U689 (N_689,In_787,In_570);
nand U690 (N_690,In_205,In_364);
or U691 (N_691,In_325,In_65);
nor U692 (N_692,In_19,In_815);
nor U693 (N_693,In_602,In_520);
nand U694 (N_694,In_989,In_62);
and U695 (N_695,In_14,In_786);
nor U696 (N_696,In_345,In_486);
nand U697 (N_697,In_590,In_68);
and U698 (N_698,In_240,In_668);
or U699 (N_699,In_232,In_604);
and U700 (N_700,In_89,In_843);
nor U701 (N_701,In_288,In_920);
or U702 (N_702,In_461,In_35);
or U703 (N_703,In_645,In_581);
nand U704 (N_704,In_535,In_207);
or U705 (N_705,In_278,In_104);
nand U706 (N_706,In_521,In_158);
and U707 (N_707,In_291,In_340);
nand U708 (N_708,In_477,In_909);
and U709 (N_709,In_280,In_217);
nor U710 (N_710,In_169,In_15);
nor U711 (N_711,In_672,In_962);
or U712 (N_712,In_526,In_385);
and U713 (N_713,In_775,In_433);
and U714 (N_714,In_822,In_615);
nand U715 (N_715,In_398,In_679);
nor U716 (N_716,In_277,In_843);
nor U717 (N_717,In_594,In_660);
or U718 (N_718,In_453,In_219);
or U719 (N_719,In_544,In_405);
or U720 (N_720,In_57,In_886);
or U721 (N_721,In_429,In_261);
xnor U722 (N_722,In_745,In_154);
or U723 (N_723,In_733,In_445);
or U724 (N_724,In_398,In_553);
or U725 (N_725,In_810,In_149);
and U726 (N_726,In_533,In_321);
or U727 (N_727,In_513,In_966);
nor U728 (N_728,In_535,In_331);
nand U729 (N_729,In_567,In_533);
or U730 (N_730,In_244,In_800);
and U731 (N_731,In_207,In_772);
nand U732 (N_732,In_216,In_783);
and U733 (N_733,In_473,In_278);
nor U734 (N_734,In_134,In_604);
nor U735 (N_735,In_991,In_721);
nand U736 (N_736,In_884,In_382);
or U737 (N_737,In_408,In_213);
nor U738 (N_738,In_709,In_635);
or U739 (N_739,In_189,In_286);
nor U740 (N_740,In_93,In_793);
nand U741 (N_741,In_964,In_450);
or U742 (N_742,In_769,In_575);
nor U743 (N_743,In_483,In_916);
nor U744 (N_744,In_385,In_414);
nand U745 (N_745,In_132,In_896);
or U746 (N_746,In_183,In_679);
nand U747 (N_747,In_272,In_24);
or U748 (N_748,In_622,In_872);
nand U749 (N_749,In_127,In_75);
or U750 (N_750,In_195,In_18);
nor U751 (N_751,In_814,In_11);
or U752 (N_752,In_100,In_106);
or U753 (N_753,In_705,In_185);
or U754 (N_754,In_134,In_728);
and U755 (N_755,In_512,In_754);
or U756 (N_756,In_551,In_482);
nand U757 (N_757,In_129,In_859);
and U758 (N_758,In_564,In_50);
and U759 (N_759,In_337,In_878);
or U760 (N_760,In_725,In_652);
nor U761 (N_761,In_686,In_578);
nor U762 (N_762,In_660,In_33);
or U763 (N_763,In_278,In_612);
xor U764 (N_764,In_767,In_106);
and U765 (N_765,In_97,In_548);
nand U766 (N_766,In_420,In_717);
nand U767 (N_767,In_438,In_829);
nor U768 (N_768,In_80,In_319);
nor U769 (N_769,In_73,In_88);
and U770 (N_770,In_718,In_126);
or U771 (N_771,In_237,In_689);
nand U772 (N_772,In_781,In_664);
nor U773 (N_773,In_675,In_713);
or U774 (N_774,In_519,In_522);
nand U775 (N_775,In_458,In_993);
nand U776 (N_776,In_308,In_942);
or U777 (N_777,In_429,In_921);
nor U778 (N_778,In_546,In_138);
nor U779 (N_779,In_446,In_175);
nand U780 (N_780,In_826,In_911);
and U781 (N_781,In_765,In_955);
nand U782 (N_782,In_457,In_19);
nor U783 (N_783,In_958,In_718);
or U784 (N_784,In_648,In_689);
or U785 (N_785,In_295,In_348);
and U786 (N_786,In_959,In_549);
nor U787 (N_787,In_863,In_109);
nand U788 (N_788,In_802,In_964);
or U789 (N_789,In_340,In_819);
or U790 (N_790,In_647,In_856);
or U791 (N_791,In_408,In_737);
nor U792 (N_792,In_128,In_175);
nor U793 (N_793,In_592,In_111);
or U794 (N_794,In_96,In_225);
and U795 (N_795,In_493,In_198);
nor U796 (N_796,In_418,In_750);
nor U797 (N_797,In_893,In_937);
or U798 (N_798,In_956,In_509);
and U799 (N_799,In_815,In_140);
nor U800 (N_800,In_143,In_869);
and U801 (N_801,In_78,In_970);
and U802 (N_802,In_412,In_918);
nand U803 (N_803,In_699,In_105);
nand U804 (N_804,In_523,In_378);
or U805 (N_805,In_8,In_884);
or U806 (N_806,In_110,In_447);
nand U807 (N_807,In_639,In_600);
and U808 (N_808,In_131,In_463);
and U809 (N_809,In_132,In_621);
nor U810 (N_810,In_600,In_946);
and U811 (N_811,In_578,In_690);
and U812 (N_812,In_496,In_596);
or U813 (N_813,In_315,In_549);
and U814 (N_814,In_437,In_504);
nand U815 (N_815,In_618,In_823);
nand U816 (N_816,In_117,In_756);
or U817 (N_817,In_125,In_265);
and U818 (N_818,In_160,In_78);
xor U819 (N_819,In_875,In_223);
nor U820 (N_820,In_950,In_16);
and U821 (N_821,In_701,In_691);
nand U822 (N_822,In_107,In_720);
nor U823 (N_823,In_103,In_449);
and U824 (N_824,In_827,In_781);
or U825 (N_825,In_109,In_796);
and U826 (N_826,In_954,In_586);
and U827 (N_827,In_407,In_825);
nand U828 (N_828,In_48,In_207);
nor U829 (N_829,In_808,In_439);
or U830 (N_830,In_291,In_542);
nor U831 (N_831,In_695,In_489);
nor U832 (N_832,In_142,In_109);
nor U833 (N_833,In_171,In_268);
and U834 (N_834,In_503,In_829);
nand U835 (N_835,In_325,In_977);
and U836 (N_836,In_321,In_683);
xor U837 (N_837,In_674,In_978);
and U838 (N_838,In_456,In_685);
nor U839 (N_839,In_372,In_748);
or U840 (N_840,In_528,In_331);
nor U841 (N_841,In_911,In_434);
or U842 (N_842,In_924,In_355);
or U843 (N_843,In_321,In_402);
and U844 (N_844,In_731,In_784);
or U845 (N_845,In_546,In_133);
nand U846 (N_846,In_613,In_751);
nor U847 (N_847,In_380,In_354);
nor U848 (N_848,In_174,In_608);
or U849 (N_849,In_35,In_931);
nor U850 (N_850,In_570,In_963);
nand U851 (N_851,In_264,In_918);
or U852 (N_852,In_782,In_238);
nand U853 (N_853,In_553,In_451);
nor U854 (N_854,In_284,In_848);
or U855 (N_855,In_571,In_406);
and U856 (N_856,In_766,In_877);
nor U857 (N_857,In_343,In_901);
and U858 (N_858,In_231,In_446);
nor U859 (N_859,In_191,In_844);
nor U860 (N_860,In_33,In_644);
and U861 (N_861,In_399,In_322);
or U862 (N_862,In_228,In_538);
nor U863 (N_863,In_591,In_161);
nand U864 (N_864,In_224,In_418);
and U865 (N_865,In_263,In_235);
nand U866 (N_866,In_479,In_899);
or U867 (N_867,In_452,In_627);
nor U868 (N_868,In_685,In_683);
or U869 (N_869,In_110,In_656);
or U870 (N_870,In_493,In_162);
nand U871 (N_871,In_290,In_415);
nor U872 (N_872,In_516,In_581);
or U873 (N_873,In_508,In_850);
and U874 (N_874,In_532,In_122);
and U875 (N_875,In_297,In_138);
nand U876 (N_876,In_211,In_135);
nor U877 (N_877,In_820,In_476);
or U878 (N_878,In_302,In_530);
and U879 (N_879,In_246,In_116);
nand U880 (N_880,In_317,In_709);
nor U881 (N_881,In_927,In_328);
or U882 (N_882,In_16,In_639);
nand U883 (N_883,In_176,In_191);
or U884 (N_884,In_124,In_240);
nor U885 (N_885,In_554,In_843);
nor U886 (N_886,In_310,In_668);
or U887 (N_887,In_698,In_883);
nand U888 (N_888,In_973,In_421);
and U889 (N_889,In_348,In_720);
nor U890 (N_890,In_956,In_305);
or U891 (N_891,In_311,In_336);
nor U892 (N_892,In_142,In_981);
nor U893 (N_893,In_331,In_868);
or U894 (N_894,In_239,In_217);
and U895 (N_895,In_560,In_118);
or U896 (N_896,In_555,In_862);
and U897 (N_897,In_868,In_971);
or U898 (N_898,In_91,In_146);
nand U899 (N_899,In_392,In_305);
or U900 (N_900,In_33,In_82);
nand U901 (N_901,In_489,In_445);
or U902 (N_902,In_237,In_272);
nor U903 (N_903,In_327,In_152);
or U904 (N_904,In_40,In_28);
nor U905 (N_905,In_242,In_775);
or U906 (N_906,In_53,In_404);
nand U907 (N_907,In_217,In_633);
nor U908 (N_908,In_467,In_564);
nor U909 (N_909,In_192,In_907);
and U910 (N_910,In_782,In_929);
nor U911 (N_911,In_81,In_431);
nor U912 (N_912,In_273,In_860);
or U913 (N_913,In_645,In_783);
and U914 (N_914,In_27,In_942);
or U915 (N_915,In_92,In_449);
or U916 (N_916,In_988,In_964);
nor U917 (N_917,In_676,In_555);
nand U918 (N_918,In_955,In_756);
nor U919 (N_919,In_166,In_113);
nor U920 (N_920,In_881,In_618);
nand U921 (N_921,In_345,In_928);
or U922 (N_922,In_837,In_99);
or U923 (N_923,In_472,In_596);
or U924 (N_924,In_785,In_638);
and U925 (N_925,In_690,In_549);
or U926 (N_926,In_56,In_277);
or U927 (N_927,In_782,In_993);
or U928 (N_928,In_487,In_493);
or U929 (N_929,In_776,In_648);
and U930 (N_930,In_741,In_968);
or U931 (N_931,In_841,In_716);
and U932 (N_932,In_96,In_512);
and U933 (N_933,In_511,In_671);
nand U934 (N_934,In_821,In_416);
nor U935 (N_935,In_209,In_880);
or U936 (N_936,In_954,In_839);
nand U937 (N_937,In_173,In_838);
nor U938 (N_938,In_157,In_137);
nand U939 (N_939,In_582,In_85);
and U940 (N_940,In_438,In_300);
nor U941 (N_941,In_452,In_78);
and U942 (N_942,In_446,In_377);
nor U943 (N_943,In_220,In_475);
nor U944 (N_944,In_78,In_750);
or U945 (N_945,In_195,In_773);
or U946 (N_946,In_783,In_320);
nor U947 (N_947,In_852,In_229);
nor U948 (N_948,In_663,In_118);
and U949 (N_949,In_909,In_149);
nor U950 (N_950,In_371,In_902);
and U951 (N_951,In_211,In_687);
or U952 (N_952,In_865,In_575);
nand U953 (N_953,In_292,In_233);
nand U954 (N_954,In_340,In_385);
xor U955 (N_955,In_646,In_768);
nand U956 (N_956,In_786,In_813);
nor U957 (N_957,In_826,In_91);
nand U958 (N_958,In_180,In_658);
or U959 (N_959,In_938,In_894);
nand U960 (N_960,In_884,In_128);
nor U961 (N_961,In_430,In_82);
or U962 (N_962,In_680,In_225);
nand U963 (N_963,In_908,In_325);
nand U964 (N_964,In_739,In_557);
and U965 (N_965,In_889,In_972);
nand U966 (N_966,In_98,In_50);
nand U967 (N_967,In_695,In_791);
or U968 (N_968,In_613,In_637);
nor U969 (N_969,In_4,In_18);
nand U970 (N_970,In_306,In_558);
nand U971 (N_971,In_263,In_0);
or U972 (N_972,In_601,In_767);
or U973 (N_973,In_88,In_111);
or U974 (N_974,In_944,In_640);
or U975 (N_975,In_211,In_948);
nand U976 (N_976,In_570,In_293);
and U977 (N_977,In_783,In_105);
and U978 (N_978,In_637,In_544);
nor U979 (N_979,In_919,In_539);
nor U980 (N_980,In_618,In_450);
and U981 (N_981,In_513,In_639);
or U982 (N_982,In_571,In_52);
or U983 (N_983,In_760,In_248);
or U984 (N_984,In_231,In_308);
and U985 (N_985,In_23,In_689);
and U986 (N_986,In_101,In_557);
and U987 (N_987,In_442,In_741);
nor U988 (N_988,In_375,In_635);
nand U989 (N_989,In_99,In_329);
and U990 (N_990,In_379,In_772);
nand U991 (N_991,In_119,In_271);
nor U992 (N_992,In_142,In_260);
nand U993 (N_993,In_97,In_511);
xnor U994 (N_994,In_81,In_720);
nand U995 (N_995,In_695,In_780);
nor U996 (N_996,In_644,In_361);
nand U997 (N_997,In_237,In_297);
nand U998 (N_998,In_554,In_438);
nand U999 (N_999,In_673,In_728);
nor U1000 (N_1000,N_6,N_949);
or U1001 (N_1001,N_987,N_384);
or U1002 (N_1002,N_293,N_883);
nand U1003 (N_1003,N_918,N_508);
nor U1004 (N_1004,N_386,N_421);
or U1005 (N_1005,N_194,N_604);
nor U1006 (N_1006,N_335,N_104);
nand U1007 (N_1007,N_704,N_866);
nor U1008 (N_1008,N_734,N_171);
and U1009 (N_1009,N_702,N_84);
or U1010 (N_1010,N_499,N_433);
or U1011 (N_1011,N_338,N_698);
nor U1012 (N_1012,N_462,N_321);
and U1013 (N_1013,N_515,N_929);
or U1014 (N_1014,N_332,N_182);
and U1015 (N_1015,N_145,N_583);
nor U1016 (N_1016,N_270,N_616);
or U1017 (N_1017,N_306,N_831);
and U1018 (N_1018,N_134,N_699);
and U1019 (N_1019,N_888,N_633);
or U1020 (N_1020,N_302,N_18);
or U1021 (N_1021,N_453,N_994);
nor U1022 (N_1022,N_512,N_853);
nand U1023 (N_1023,N_377,N_798);
and U1024 (N_1024,N_86,N_920);
nor U1025 (N_1025,N_37,N_347);
or U1026 (N_1026,N_303,N_305);
nor U1027 (N_1027,N_580,N_196);
and U1028 (N_1028,N_792,N_658);
and U1029 (N_1029,N_596,N_96);
or U1030 (N_1030,N_353,N_467);
nand U1031 (N_1031,N_264,N_575);
nand U1032 (N_1032,N_198,N_985);
or U1033 (N_1033,N_183,N_706);
and U1034 (N_1034,N_805,N_563);
nor U1035 (N_1035,N_739,N_214);
nand U1036 (N_1036,N_149,N_869);
nor U1037 (N_1037,N_552,N_279);
or U1038 (N_1038,N_861,N_581);
nand U1039 (N_1039,N_252,N_199);
nor U1040 (N_1040,N_285,N_585);
and U1041 (N_1041,N_218,N_977);
nand U1042 (N_1042,N_594,N_161);
nand U1043 (N_1043,N_954,N_615);
or U1044 (N_1044,N_942,N_814);
nand U1045 (N_1045,N_811,N_259);
and U1046 (N_1046,N_97,N_3);
nand U1047 (N_1047,N_824,N_40);
nand U1048 (N_1048,N_849,N_317);
nand U1049 (N_1049,N_930,N_513);
or U1050 (N_1050,N_634,N_968);
or U1051 (N_1051,N_309,N_554);
nand U1052 (N_1052,N_291,N_101);
and U1053 (N_1053,N_555,N_464);
nor U1054 (N_1054,N_736,N_156);
nand U1055 (N_1055,N_403,N_835);
nand U1056 (N_1056,N_622,N_586);
nand U1057 (N_1057,N_844,N_778);
nor U1058 (N_1058,N_848,N_1);
nand U1059 (N_1059,N_732,N_95);
or U1060 (N_1060,N_116,N_981);
nor U1061 (N_1061,N_751,N_990);
nor U1062 (N_1062,N_846,N_478);
nor U1063 (N_1063,N_39,N_928);
and U1064 (N_1064,N_414,N_221);
nand U1065 (N_1065,N_55,N_26);
and U1066 (N_1066,N_388,N_53);
nand U1067 (N_1067,N_442,N_412);
nor U1068 (N_1068,N_102,N_503);
nor U1069 (N_1069,N_986,N_187);
and U1070 (N_1070,N_885,N_185);
nand U1071 (N_1071,N_470,N_640);
and U1072 (N_1072,N_263,N_868);
nor U1073 (N_1073,N_812,N_471);
or U1074 (N_1074,N_77,N_659);
nor U1075 (N_1075,N_253,N_864);
and U1076 (N_1076,N_799,N_678);
and U1077 (N_1077,N_663,N_110);
or U1078 (N_1078,N_341,N_953);
or U1079 (N_1079,N_204,N_376);
nand U1080 (N_1080,N_489,N_813);
or U1081 (N_1081,N_289,N_141);
nor U1082 (N_1082,N_613,N_358);
and U1083 (N_1083,N_645,N_135);
nand U1084 (N_1084,N_408,N_463);
or U1085 (N_1085,N_67,N_315);
nand U1086 (N_1086,N_261,N_999);
nor U1087 (N_1087,N_184,N_875);
or U1088 (N_1088,N_806,N_748);
nand U1089 (N_1089,N_859,N_984);
and U1090 (N_1090,N_36,N_559);
and U1091 (N_1091,N_298,N_20);
nor U1092 (N_1092,N_560,N_741);
or U1093 (N_1093,N_569,N_164);
nor U1094 (N_1094,N_224,N_605);
or U1095 (N_1095,N_79,N_670);
nand U1096 (N_1096,N_617,N_44);
or U1097 (N_1097,N_111,N_874);
nor U1098 (N_1098,N_38,N_689);
nor U1099 (N_1099,N_712,N_176);
nand U1100 (N_1100,N_380,N_891);
nor U1101 (N_1101,N_480,N_206);
and U1102 (N_1102,N_11,N_200);
or U1103 (N_1103,N_375,N_250);
nor U1104 (N_1104,N_541,N_127);
nor U1105 (N_1105,N_56,N_72);
nor U1106 (N_1106,N_331,N_667);
nand U1107 (N_1107,N_34,N_351);
nor U1108 (N_1108,N_547,N_719);
nand U1109 (N_1109,N_902,N_316);
or U1110 (N_1110,N_180,N_795);
nor U1111 (N_1111,N_531,N_349);
nor U1112 (N_1112,N_644,N_657);
nor U1113 (N_1113,N_266,N_409);
and U1114 (N_1114,N_459,N_383);
nor U1115 (N_1115,N_995,N_972);
and U1116 (N_1116,N_635,N_277);
nor U1117 (N_1117,N_256,N_418);
or U1118 (N_1118,N_286,N_829);
and U1119 (N_1119,N_147,N_693);
and U1120 (N_1120,N_631,N_858);
or U1121 (N_1121,N_340,N_401);
nor U1122 (N_1122,N_235,N_679);
or U1123 (N_1123,N_788,N_852);
nor U1124 (N_1124,N_240,N_257);
nand U1125 (N_1125,N_979,N_422);
nand U1126 (N_1126,N_385,N_879);
or U1127 (N_1127,N_174,N_917);
or U1128 (N_1128,N_744,N_465);
or U1129 (N_1129,N_653,N_915);
nor U1130 (N_1130,N_241,N_405);
nor U1131 (N_1131,N_881,N_638);
or U1132 (N_1132,N_964,N_57);
or U1133 (N_1133,N_757,N_228);
nor U1134 (N_1134,N_24,N_609);
or U1135 (N_1135,N_714,N_607);
nand U1136 (N_1136,N_434,N_551);
nor U1137 (N_1137,N_121,N_25);
and U1138 (N_1138,N_724,N_664);
nand U1139 (N_1139,N_483,N_673);
nor U1140 (N_1140,N_445,N_624);
or U1141 (N_1141,N_170,N_661);
and U1142 (N_1142,N_701,N_239);
nand U1143 (N_1143,N_790,N_460);
and U1144 (N_1144,N_152,N_65);
nand U1145 (N_1145,N_991,N_826);
nor U1146 (N_1146,N_82,N_504);
or U1147 (N_1147,N_727,N_320);
or U1148 (N_1148,N_713,N_961);
or U1149 (N_1149,N_535,N_676);
and U1150 (N_1150,N_600,N_46);
nor U1151 (N_1151,N_629,N_17);
nor U1152 (N_1152,N_166,N_572);
nand U1153 (N_1153,N_735,N_907);
nand U1154 (N_1154,N_295,N_362);
nand U1155 (N_1155,N_426,N_246);
and U1156 (N_1156,N_425,N_947);
and U1157 (N_1157,N_567,N_743);
or U1158 (N_1158,N_630,N_30);
and U1159 (N_1159,N_162,N_606);
and U1160 (N_1160,N_420,N_593);
and U1161 (N_1161,N_215,N_172);
nor U1162 (N_1162,N_21,N_410);
and U1163 (N_1163,N_119,N_366);
and U1164 (N_1164,N_956,N_357);
nor U1165 (N_1165,N_820,N_530);
nor U1166 (N_1166,N_822,N_35);
nand U1167 (N_1167,N_998,N_601);
nor U1168 (N_1168,N_177,N_599);
and U1169 (N_1169,N_280,N_863);
and U1170 (N_1170,N_804,N_59);
nand U1171 (N_1171,N_900,N_330);
nand U1172 (N_1172,N_536,N_22);
nand U1173 (N_1173,N_391,N_73);
nand U1174 (N_1174,N_0,N_733);
and U1175 (N_1175,N_217,N_777);
and U1176 (N_1176,N_83,N_143);
or U1177 (N_1177,N_13,N_430);
nor U1178 (N_1178,N_534,N_131);
and U1179 (N_1179,N_4,N_784);
nor U1180 (N_1180,N_721,N_636);
nand U1181 (N_1181,N_595,N_506);
and U1182 (N_1182,N_989,N_982);
or U1183 (N_1183,N_823,N_108);
xnor U1184 (N_1184,N_85,N_202);
nor U1185 (N_1185,N_66,N_731);
or U1186 (N_1186,N_927,N_244);
nor U1187 (N_1187,N_345,N_872);
and U1188 (N_1188,N_650,N_314);
and U1189 (N_1189,N_910,N_509);
nand U1190 (N_1190,N_931,N_685);
or U1191 (N_1191,N_262,N_138);
and U1192 (N_1192,N_816,N_921);
nand U1193 (N_1193,N_120,N_943);
nand U1194 (N_1194,N_756,N_238);
or U1195 (N_1195,N_452,N_197);
nand U1196 (N_1196,N_461,N_457);
nand U1197 (N_1197,N_919,N_662);
or U1198 (N_1198,N_697,N_890);
nor U1199 (N_1199,N_807,N_873);
nor U1200 (N_1200,N_114,N_254);
nor U1201 (N_1201,N_587,N_803);
and U1202 (N_1202,N_548,N_140);
and U1203 (N_1203,N_404,N_539);
nor U1204 (N_1204,N_973,N_146);
nand U1205 (N_1205,N_287,N_359);
nor U1206 (N_1206,N_500,N_550);
and U1207 (N_1207,N_192,N_821);
or U1208 (N_1208,N_68,N_354);
or U1209 (N_1209,N_516,N_273);
nor U1210 (N_1210,N_451,N_759);
or U1211 (N_1211,N_723,N_878);
and U1212 (N_1212,N_776,N_817);
or U1213 (N_1213,N_479,N_269);
and U1214 (N_1214,N_836,N_494);
nand U1215 (N_1215,N_27,N_668);
nor U1216 (N_1216,N_571,N_641);
nor U1217 (N_1217,N_274,N_540);
and U1218 (N_1218,N_708,N_771);
and U1219 (N_1219,N_490,N_237);
nor U1220 (N_1220,N_230,N_877);
nor U1221 (N_1221,N_181,N_473);
and U1222 (N_1222,N_628,N_70);
and U1223 (N_1223,N_976,N_974);
and U1224 (N_1224,N_468,N_178);
and U1225 (N_1225,N_851,N_518);
nand U1226 (N_1226,N_389,N_847);
and U1227 (N_1227,N_325,N_382);
nor U1228 (N_1228,N_924,N_369);
and U1229 (N_1229,N_243,N_137);
nor U1230 (N_1230,N_755,N_313);
and U1231 (N_1231,N_381,N_647);
nor U1232 (N_1232,N_148,N_155);
or U1233 (N_1233,N_810,N_307);
nand U1234 (N_1234,N_406,N_481);
nand U1235 (N_1235,N_42,N_106);
or U1236 (N_1236,N_971,N_466);
nor U1237 (N_1237,N_157,N_169);
nor U1238 (N_1238,N_603,N_672);
nor U1239 (N_1239,N_703,N_220);
or U1240 (N_1240,N_781,N_87);
or U1241 (N_1241,N_850,N_533);
nand U1242 (N_1242,N_233,N_576);
nand U1243 (N_1243,N_524,N_343);
or U1244 (N_1244,N_677,N_819);
and U1245 (N_1245,N_213,N_399);
nor U1246 (N_1246,N_154,N_772);
nor U1247 (N_1247,N_520,N_591);
or U1248 (N_1248,N_397,N_128);
nand U1249 (N_1249,N_941,N_705);
nand U1250 (N_1250,N_916,N_521);
nand U1251 (N_1251,N_290,N_226);
or U1252 (N_1252,N_561,N_742);
and U1253 (N_1253,N_683,N_914);
nor U1254 (N_1254,N_249,N_808);
and U1255 (N_1255,N_894,N_654);
nor U1256 (N_1256,N_136,N_660);
nand U1257 (N_1257,N_845,N_651);
nor U1258 (N_1258,N_909,N_52);
nand U1259 (N_1259,N_933,N_416);
or U1260 (N_1260,N_492,N_589);
nand U1261 (N_1261,N_818,N_411);
nor U1262 (N_1262,N_901,N_783);
nor U1263 (N_1263,N_722,N_525);
and U1264 (N_1264,N_179,N_758);
and U1265 (N_1265,N_529,N_281);
and U1266 (N_1266,N_502,N_598);
nor U1267 (N_1267,N_276,N_711);
and U1268 (N_1268,N_203,N_940);
nor U1269 (N_1269,N_553,N_28);
or U1270 (N_1270,N_681,N_472);
nand U1271 (N_1271,N_669,N_564);
nand U1272 (N_1272,N_671,N_590);
or U1273 (N_1273,N_336,N_532);
or U1274 (N_1274,N_770,N_123);
nor U1275 (N_1275,N_895,N_173);
nand U1276 (N_1276,N_841,N_730);
and U1277 (N_1277,N_620,N_160);
nand U1278 (N_1278,N_9,N_800);
nand U1279 (N_1279,N_398,N_746);
nor U1280 (N_1280,N_912,N_7);
and U1281 (N_1281,N_584,N_328);
nor U1282 (N_1282,N_725,N_275);
nand U1283 (N_1283,N_691,N_687);
nor U1284 (N_1284,N_477,N_402);
nand U1285 (N_1285,N_579,N_519);
nand U1286 (N_1286,N_260,N_71);
nand U1287 (N_1287,N_573,N_311);
nand U1288 (N_1288,N_210,N_793);
or U1289 (N_1289,N_454,N_151);
xor U1290 (N_1290,N_505,N_392);
and U1291 (N_1291,N_74,N_892);
or U1292 (N_1292,N_674,N_545);
nand U1293 (N_1293,N_886,N_939);
and U1294 (N_1294,N_718,N_248);
nand U1295 (N_1295,N_150,N_365);
nor U1296 (N_1296,N_549,N_132);
or U1297 (N_1297,N_62,N_117);
or U1298 (N_1298,N_245,N_191);
nand U1299 (N_1299,N_193,N_165);
nand U1300 (N_1300,N_642,N_766);
nand U1301 (N_1301,N_448,N_692);
nor U1302 (N_1302,N_337,N_458);
nand U1303 (N_1303,N_301,N_159);
nand U1304 (N_1304,N_913,N_326);
nand U1305 (N_1305,N_163,N_501);
or U1306 (N_1306,N_544,N_537);
nand U1307 (N_1307,N_429,N_809);
nor U1308 (N_1308,N_396,N_843);
nand U1309 (N_1309,N_577,N_566);
nor U1310 (N_1310,N_334,N_686);
nand U1311 (N_1311,N_839,N_431);
nand U1312 (N_1312,N_574,N_267);
or U1313 (N_1313,N_94,N_107);
and U1314 (N_1314,N_284,N_729);
nor U1315 (N_1315,N_690,N_133);
and U1316 (N_1316,N_887,N_542);
and U1317 (N_1317,N_374,N_675);
nor U1318 (N_1318,N_455,N_578);
and U1319 (N_1319,N_632,N_379);
nor U1320 (N_1320,N_967,N_614);
nand U1321 (N_1321,N_830,N_324);
and U1322 (N_1322,N_911,N_763);
and U1323 (N_1323,N_996,N_882);
and U1324 (N_1324,N_762,N_205);
nor U1325 (N_1325,N_89,N_978);
or U1326 (N_1326,N_970,N_854);
or U1327 (N_1327,N_960,N_282);
or U1328 (N_1328,N_342,N_61);
and U1329 (N_1329,N_76,N_568);
nor U1330 (N_1330,N_372,N_597);
or U1331 (N_1331,N_292,N_760);
or U1332 (N_1332,N_112,N_526);
nor U1333 (N_1333,N_618,N_47);
nor U1334 (N_1334,N_415,N_925);
nor U1335 (N_1335,N_258,N_906);
and U1336 (N_1336,N_958,N_219);
or U1337 (N_1337,N_236,N_125);
nand U1338 (N_1338,N_265,N_364);
and U1339 (N_1339,N_728,N_842);
and U1340 (N_1340,N_435,N_153);
and U1341 (N_1341,N_754,N_427);
nor U1342 (N_1342,N_951,N_90);
or U1343 (N_1343,N_955,N_498);
and U1344 (N_1344,N_761,N_139);
or U1345 (N_1345,N_207,N_283);
and U1346 (N_1346,N_333,N_223);
or U1347 (N_1347,N_495,N_41);
nor U1348 (N_1348,N_707,N_216);
nand U1349 (N_1349,N_440,N_255);
nand U1350 (N_1350,N_78,N_740);
nand U1351 (N_1351,N_833,N_959);
nor U1352 (N_1352,N_827,N_656);
nand U1353 (N_1353,N_898,N_558);
nor U1354 (N_1354,N_31,N_60);
and U1355 (N_1355,N_749,N_680);
nand U1356 (N_1356,N_363,N_105);
and U1357 (N_1357,N_825,N_15);
and U1358 (N_1358,N_118,N_130);
and U1359 (N_1359,N_511,N_393);
or U1360 (N_1360,N_665,N_528);
and U1361 (N_1361,N_45,N_5);
and U1362 (N_1362,N_952,N_700);
nand U1363 (N_1363,N_14,N_937);
nand U1364 (N_1364,N_715,N_58);
nand U1365 (N_1365,N_945,N_493);
nor U1366 (N_1366,N_175,N_838);
or U1367 (N_1367,N_889,N_791);
nor U1368 (N_1368,N_815,N_753);
or U1369 (N_1369,N_684,N_122);
or U1370 (N_1370,N_562,N_626);
nor U1371 (N_1371,N_497,N_507);
nand U1372 (N_1372,N_908,N_946);
and U1373 (N_1373,N_441,N_229);
nor U1374 (N_1374,N_49,N_247);
nor U1375 (N_1375,N_787,N_720);
or U1376 (N_1376,N_510,N_447);
nor U1377 (N_1377,N_201,N_208);
xor U1378 (N_1378,N_950,N_648);
and U1379 (N_1379,N_2,N_546);
or U1380 (N_1380,N_75,N_438);
nand U1381 (N_1381,N_491,N_966);
nor U1382 (N_1382,N_789,N_649);
or U1383 (N_1383,N_474,N_752);
and U1384 (N_1384,N_69,N_329);
nor U1385 (N_1385,N_469,N_80);
nor U1386 (N_1386,N_352,N_965);
and U1387 (N_1387,N_834,N_932);
nand U1388 (N_1388,N_304,N_768);
and U1389 (N_1389,N_738,N_802);
and U1390 (N_1390,N_33,N_299);
and U1391 (N_1391,N_637,N_419);
nor U1392 (N_1392,N_319,N_840);
nor U1393 (N_1393,N_227,N_860);
and U1394 (N_1394,N_983,N_610);
nor U1395 (N_1395,N_934,N_767);
or U1396 (N_1396,N_23,N_407);
and U1397 (N_1397,N_450,N_242);
nand U1398 (N_1398,N_167,N_710);
nand U1399 (N_1399,N_129,N_485);
nor U1400 (N_1400,N_837,N_8);
or U1401 (N_1401,N_627,N_764);
nand U1402 (N_1402,N_32,N_969);
and U1403 (N_1403,N_271,N_186);
xnor U1404 (N_1404,N_619,N_300);
or U1405 (N_1405,N_88,N_871);
and U1406 (N_1406,N_592,N_361);
and U1407 (N_1407,N_896,N_444);
and U1408 (N_1408,N_993,N_437);
nor U1409 (N_1409,N_211,N_523);
and U1410 (N_1410,N_666,N_439);
nor U1411 (N_1411,N_99,N_115);
and U1412 (N_1412,N_655,N_527);
and U1413 (N_1413,N_50,N_312);
nand U1414 (N_1414,N_588,N_310);
nand U1415 (N_1415,N_517,N_63);
nand U1416 (N_1416,N_988,N_904);
or U1417 (N_1417,N_785,N_98);
or U1418 (N_1418,N_16,N_142);
nor U1419 (N_1419,N_225,N_144);
nor U1420 (N_1420,N_64,N_963);
nor U1421 (N_1421,N_602,N_297);
nor U1422 (N_1422,N_621,N_780);
nor U1423 (N_1423,N_944,N_387);
and U1424 (N_1424,N_476,N_926);
nor U1425 (N_1425,N_371,N_694);
or U1426 (N_1426,N_980,N_456);
and U1427 (N_1427,N_54,N_124);
or U1428 (N_1428,N_899,N_514);
or U1429 (N_1429,N_884,N_696);
or U1430 (N_1430,N_737,N_828);
and U1431 (N_1431,N_765,N_623);
nor U1432 (N_1432,N_350,N_796);
nor U1433 (N_1433,N_272,N_346);
or U1434 (N_1434,N_323,N_475);
nand U1435 (N_1435,N_126,N_368);
nand U1436 (N_1436,N_234,N_231);
or U1437 (N_1437,N_488,N_19);
nand U1438 (N_1438,N_832,N_557);
or U1439 (N_1439,N_268,N_413);
nand U1440 (N_1440,N_10,N_93);
and U1441 (N_1441,N_893,N_936);
nor U1442 (N_1442,N_327,N_774);
nor U1443 (N_1443,N_100,N_482);
nor U1444 (N_1444,N_356,N_782);
nand U1445 (N_1445,N_29,N_611);
and U1446 (N_1446,N_773,N_652);
nor U1447 (N_1447,N_903,N_709);
and U1448 (N_1448,N_188,N_582);
nand U1449 (N_1449,N_367,N_390);
nand U1450 (N_1450,N_747,N_432);
nand U1451 (N_1451,N_318,N_189);
and U1452 (N_1452,N_113,N_570);
or U1453 (N_1453,N_103,N_543);
nand U1454 (N_1454,N_688,N_639);
nand U1455 (N_1455,N_797,N_308);
nor U1456 (N_1456,N_209,N_905);
xnor U1457 (N_1457,N_296,N_643);
or U1458 (N_1458,N_922,N_158);
or U1459 (N_1459,N_794,N_190);
nor U1460 (N_1460,N_565,N_923);
nor U1461 (N_1461,N_12,N_195);
nand U1462 (N_1462,N_935,N_355);
or U1463 (N_1463,N_51,N_436);
and U1464 (N_1464,N_556,N_443);
and U1465 (N_1465,N_339,N_92);
xor U1466 (N_1466,N_344,N_880);
nor U1467 (N_1467,N_484,N_486);
or U1468 (N_1468,N_109,N_938);
nor U1469 (N_1469,N_856,N_538);
or U1470 (N_1470,N_865,N_682);
and U1471 (N_1471,N_717,N_378);
nand U1472 (N_1472,N_855,N_769);
or U1473 (N_1473,N_294,N_948);
or U1474 (N_1474,N_322,N_348);
nand U1475 (N_1475,N_222,N_962);
nor U1476 (N_1476,N_625,N_360);
and U1477 (N_1477,N_801,N_775);
nand U1478 (N_1478,N_779,N_695);
or U1479 (N_1479,N_750,N_997);
nand U1480 (N_1480,N_394,N_424);
or U1481 (N_1481,N_370,N_212);
nand U1482 (N_1482,N_168,N_876);
nand U1483 (N_1483,N_251,N_957);
or U1484 (N_1484,N_43,N_608);
and U1485 (N_1485,N_857,N_867);
nor U1486 (N_1486,N_975,N_395);
or U1487 (N_1487,N_522,N_400);
nand U1488 (N_1488,N_446,N_726);
or U1489 (N_1489,N_646,N_81);
and U1490 (N_1490,N_496,N_278);
or U1491 (N_1491,N_288,N_91);
nor U1492 (N_1492,N_870,N_423);
and U1493 (N_1493,N_612,N_487);
nand U1494 (N_1494,N_373,N_417);
nand U1495 (N_1495,N_992,N_449);
or U1496 (N_1496,N_745,N_862);
and U1497 (N_1497,N_897,N_786);
xor U1498 (N_1498,N_716,N_48);
nor U1499 (N_1499,N_428,N_232);
xor U1500 (N_1500,N_743,N_403);
and U1501 (N_1501,N_869,N_133);
and U1502 (N_1502,N_121,N_199);
nand U1503 (N_1503,N_614,N_409);
nor U1504 (N_1504,N_214,N_787);
and U1505 (N_1505,N_381,N_273);
nor U1506 (N_1506,N_932,N_219);
or U1507 (N_1507,N_277,N_983);
nor U1508 (N_1508,N_679,N_312);
nor U1509 (N_1509,N_786,N_787);
nor U1510 (N_1510,N_642,N_545);
and U1511 (N_1511,N_69,N_85);
and U1512 (N_1512,N_594,N_646);
nand U1513 (N_1513,N_602,N_511);
or U1514 (N_1514,N_108,N_681);
and U1515 (N_1515,N_966,N_232);
or U1516 (N_1516,N_45,N_934);
nand U1517 (N_1517,N_144,N_143);
and U1518 (N_1518,N_380,N_767);
nor U1519 (N_1519,N_88,N_547);
or U1520 (N_1520,N_191,N_242);
and U1521 (N_1521,N_547,N_865);
nand U1522 (N_1522,N_890,N_669);
or U1523 (N_1523,N_250,N_918);
or U1524 (N_1524,N_807,N_886);
and U1525 (N_1525,N_961,N_418);
or U1526 (N_1526,N_44,N_796);
nor U1527 (N_1527,N_924,N_824);
or U1528 (N_1528,N_129,N_251);
nand U1529 (N_1529,N_639,N_768);
nor U1530 (N_1530,N_562,N_69);
or U1531 (N_1531,N_902,N_113);
and U1532 (N_1532,N_699,N_264);
and U1533 (N_1533,N_659,N_366);
nand U1534 (N_1534,N_858,N_108);
nand U1535 (N_1535,N_266,N_325);
nand U1536 (N_1536,N_800,N_807);
and U1537 (N_1537,N_582,N_740);
nor U1538 (N_1538,N_209,N_774);
nand U1539 (N_1539,N_658,N_345);
and U1540 (N_1540,N_666,N_914);
and U1541 (N_1541,N_346,N_779);
nand U1542 (N_1542,N_709,N_620);
nand U1543 (N_1543,N_545,N_287);
and U1544 (N_1544,N_969,N_805);
or U1545 (N_1545,N_795,N_617);
nand U1546 (N_1546,N_478,N_439);
nor U1547 (N_1547,N_99,N_197);
nor U1548 (N_1548,N_361,N_573);
and U1549 (N_1549,N_750,N_18);
nand U1550 (N_1550,N_21,N_670);
nand U1551 (N_1551,N_396,N_360);
nand U1552 (N_1552,N_823,N_728);
and U1553 (N_1553,N_793,N_329);
nand U1554 (N_1554,N_367,N_546);
nor U1555 (N_1555,N_732,N_173);
nand U1556 (N_1556,N_152,N_863);
nand U1557 (N_1557,N_160,N_578);
nand U1558 (N_1558,N_672,N_69);
and U1559 (N_1559,N_710,N_815);
and U1560 (N_1560,N_850,N_642);
and U1561 (N_1561,N_282,N_287);
nand U1562 (N_1562,N_50,N_859);
and U1563 (N_1563,N_755,N_971);
and U1564 (N_1564,N_641,N_862);
or U1565 (N_1565,N_258,N_419);
nand U1566 (N_1566,N_274,N_485);
or U1567 (N_1567,N_918,N_895);
or U1568 (N_1568,N_966,N_386);
nand U1569 (N_1569,N_908,N_360);
or U1570 (N_1570,N_148,N_75);
or U1571 (N_1571,N_932,N_916);
nor U1572 (N_1572,N_470,N_925);
and U1573 (N_1573,N_665,N_436);
nor U1574 (N_1574,N_293,N_643);
nand U1575 (N_1575,N_661,N_292);
or U1576 (N_1576,N_811,N_649);
nand U1577 (N_1577,N_726,N_508);
or U1578 (N_1578,N_262,N_492);
nor U1579 (N_1579,N_303,N_259);
nor U1580 (N_1580,N_390,N_522);
or U1581 (N_1581,N_228,N_497);
nor U1582 (N_1582,N_253,N_714);
or U1583 (N_1583,N_498,N_809);
and U1584 (N_1584,N_364,N_585);
xnor U1585 (N_1585,N_95,N_773);
nor U1586 (N_1586,N_416,N_378);
nand U1587 (N_1587,N_990,N_97);
and U1588 (N_1588,N_870,N_680);
and U1589 (N_1589,N_353,N_564);
nand U1590 (N_1590,N_28,N_502);
and U1591 (N_1591,N_849,N_35);
nand U1592 (N_1592,N_443,N_536);
or U1593 (N_1593,N_658,N_597);
nor U1594 (N_1594,N_138,N_539);
xor U1595 (N_1595,N_345,N_705);
and U1596 (N_1596,N_3,N_222);
nand U1597 (N_1597,N_988,N_181);
nand U1598 (N_1598,N_824,N_467);
or U1599 (N_1599,N_785,N_25);
nand U1600 (N_1600,N_713,N_202);
or U1601 (N_1601,N_68,N_595);
nand U1602 (N_1602,N_851,N_947);
and U1603 (N_1603,N_211,N_253);
and U1604 (N_1604,N_619,N_784);
nor U1605 (N_1605,N_624,N_995);
nor U1606 (N_1606,N_436,N_240);
nand U1607 (N_1607,N_802,N_403);
nand U1608 (N_1608,N_74,N_489);
nand U1609 (N_1609,N_993,N_495);
nor U1610 (N_1610,N_481,N_468);
and U1611 (N_1611,N_344,N_404);
or U1612 (N_1612,N_923,N_23);
nor U1613 (N_1613,N_157,N_861);
and U1614 (N_1614,N_580,N_471);
or U1615 (N_1615,N_716,N_644);
nor U1616 (N_1616,N_678,N_341);
nor U1617 (N_1617,N_276,N_95);
nand U1618 (N_1618,N_486,N_889);
nor U1619 (N_1619,N_673,N_595);
nor U1620 (N_1620,N_594,N_525);
nand U1621 (N_1621,N_524,N_919);
nor U1622 (N_1622,N_981,N_854);
nor U1623 (N_1623,N_824,N_113);
nand U1624 (N_1624,N_178,N_511);
or U1625 (N_1625,N_881,N_462);
and U1626 (N_1626,N_293,N_31);
xnor U1627 (N_1627,N_159,N_780);
nand U1628 (N_1628,N_28,N_195);
nand U1629 (N_1629,N_27,N_327);
and U1630 (N_1630,N_653,N_78);
nor U1631 (N_1631,N_476,N_254);
and U1632 (N_1632,N_850,N_161);
and U1633 (N_1633,N_351,N_318);
nand U1634 (N_1634,N_539,N_895);
nand U1635 (N_1635,N_249,N_661);
nand U1636 (N_1636,N_626,N_475);
and U1637 (N_1637,N_769,N_531);
nand U1638 (N_1638,N_699,N_490);
nand U1639 (N_1639,N_551,N_158);
and U1640 (N_1640,N_338,N_827);
nor U1641 (N_1641,N_291,N_626);
and U1642 (N_1642,N_909,N_768);
nand U1643 (N_1643,N_795,N_335);
or U1644 (N_1644,N_962,N_63);
nor U1645 (N_1645,N_253,N_565);
nand U1646 (N_1646,N_368,N_364);
and U1647 (N_1647,N_252,N_470);
and U1648 (N_1648,N_935,N_839);
or U1649 (N_1649,N_937,N_50);
and U1650 (N_1650,N_3,N_521);
nand U1651 (N_1651,N_6,N_703);
nand U1652 (N_1652,N_892,N_213);
nor U1653 (N_1653,N_327,N_271);
nor U1654 (N_1654,N_574,N_22);
and U1655 (N_1655,N_428,N_583);
nor U1656 (N_1656,N_990,N_101);
and U1657 (N_1657,N_220,N_345);
nand U1658 (N_1658,N_578,N_613);
nor U1659 (N_1659,N_42,N_435);
or U1660 (N_1660,N_102,N_850);
or U1661 (N_1661,N_115,N_566);
and U1662 (N_1662,N_800,N_945);
nand U1663 (N_1663,N_762,N_738);
or U1664 (N_1664,N_38,N_925);
and U1665 (N_1665,N_97,N_967);
and U1666 (N_1666,N_731,N_558);
or U1667 (N_1667,N_686,N_931);
or U1668 (N_1668,N_136,N_446);
nor U1669 (N_1669,N_596,N_514);
nand U1670 (N_1670,N_842,N_654);
nor U1671 (N_1671,N_365,N_80);
nand U1672 (N_1672,N_945,N_351);
and U1673 (N_1673,N_337,N_154);
nor U1674 (N_1674,N_385,N_201);
nand U1675 (N_1675,N_857,N_375);
nor U1676 (N_1676,N_305,N_92);
nor U1677 (N_1677,N_648,N_614);
nor U1678 (N_1678,N_3,N_596);
or U1679 (N_1679,N_598,N_21);
nor U1680 (N_1680,N_738,N_308);
nand U1681 (N_1681,N_567,N_8);
nand U1682 (N_1682,N_472,N_680);
and U1683 (N_1683,N_101,N_106);
or U1684 (N_1684,N_958,N_424);
nand U1685 (N_1685,N_921,N_234);
nand U1686 (N_1686,N_626,N_526);
or U1687 (N_1687,N_922,N_250);
or U1688 (N_1688,N_755,N_298);
nor U1689 (N_1689,N_291,N_240);
nand U1690 (N_1690,N_859,N_903);
xnor U1691 (N_1691,N_529,N_770);
nor U1692 (N_1692,N_334,N_368);
and U1693 (N_1693,N_415,N_945);
nor U1694 (N_1694,N_470,N_805);
or U1695 (N_1695,N_828,N_968);
nor U1696 (N_1696,N_488,N_964);
and U1697 (N_1697,N_622,N_382);
and U1698 (N_1698,N_225,N_286);
nand U1699 (N_1699,N_336,N_214);
and U1700 (N_1700,N_399,N_531);
or U1701 (N_1701,N_462,N_661);
nand U1702 (N_1702,N_767,N_929);
and U1703 (N_1703,N_868,N_792);
and U1704 (N_1704,N_484,N_885);
and U1705 (N_1705,N_160,N_883);
nand U1706 (N_1706,N_870,N_158);
nor U1707 (N_1707,N_748,N_965);
and U1708 (N_1708,N_19,N_39);
nand U1709 (N_1709,N_981,N_156);
or U1710 (N_1710,N_719,N_33);
and U1711 (N_1711,N_650,N_588);
or U1712 (N_1712,N_557,N_14);
or U1713 (N_1713,N_813,N_35);
xnor U1714 (N_1714,N_375,N_89);
or U1715 (N_1715,N_333,N_920);
nor U1716 (N_1716,N_489,N_278);
or U1717 (N_1717,N_827,N_783);
and U1718 (N_1718,N_459,N_455);
nor U1719 (N_1719,N_635,N_848);
and U1720 (N_1720,N_902,N_694);
and U1721 (N_1721,N_802,N_858);
and U1722 (N_1722,N_796,N_535);
nor U1723 (N_1723,N_398,N_829);
nor U1724 (N_1724,N_703,N_379);
or U1725 (N_1725,N_729,N_260);
nand U1726 (N_1726,N_452,N_63);
nor U1727 (N_1727,N_776,N_246);
nor U1728 (N_1728,N_9,N_484);
and U1729 (N_1729,N_689,N_299);
nand U1730 (N_1730,N_300,N_851);
nand U1731 (N_1731,N_350,N_102);
and U1732 (N_1732,N_165,N_461);
and U1733 (N_1733,N_904,N_175);
nand U1734 (N_1734,N_437,N_915);
nand U1735 (N_1735,N_259,N_851);
nand U1736 (N_1736,N_102,N_388);
or U1737 (N_1737,N_929,N_865);
nor U1738 (N_1738,N_322,N_729);
and U1739 (N_1739,N_341,N_76);
or U1740 (N_1740,N_1,N_407);
xnor U1741 (N_1741,N_131,N_63);
nor U1742 (N_1742,N_263,N_711);
or U1743 (N_1743,N_999,N_73);
nand U1744 (N_1744,N_911,N_312);
and U1745 (N_1745,N_389,N_58);
nand U1746 (N_1746,N_503,N_28);
nor U1747 (N_1747,N_417,N_687);
and U1748 (N_1748,N_310,N_355);
xnor U1749 (N_1749,N_36,N_13);
nor U1750 (N_1750,N_399,N_763);
or U1751 (N_1751,N_707,N_571);
or U1752 (N_1752,N_131,N_828);
nand U1753 (N_1753,N_677,N_359);
and U1754 (N_1754,N_213,N_905);
nor U1755 (N_1755,N_640,N_292);
and U1756 (N_1756,N_840,N_184);
and U1757 (N_1757,N_856,N_991);
nand U1758 (N_1758,N_712,N_394);
and U1759 (N_1759,N_502,N_277);
nor U1760 (N_1760,N_502,N_599);
or U1761 (N_1761,N_773,N_134);
nor U1762 (N_1762,N_390,N_627);
nor U1763 (N_1763,N_369,N_26);
and U1764 (N_1764,N_523,N_779);
and U1765 (N_1765,N_720,N_698);
and U1766 (N_1766,N_707,N_662);
or U1767 (N_1767,N_755,N_34);
or U1768 (N_1768,N_701,N_346);
nand U1769 (N_1769,N_999,N_182);
nand U1770 (N_1770,N_436,N_352);
nand U1771 (N_1771,N_648,N_754);
xor U1772 (N_1772,N_724,N_288);
or U1773 (N_1773,N_998,N_630);
or U1774 (N_1774,N_846,N_381);
nand U1775 (N_1775,N_660,N_509);
or U1776 (N_1776,N_320,N_526);
or U1777 (N_1777,N_791,N_630);
nand U1778 (N_1778,N_593,N_623);
nand U1779 (N_1779,N_277,N_431);
nand U1780 (N_1780,N_3,N_144);
nor U1781 (N_1781,N_655,N_773);
or U1782 (N_1782,N_215,N_26);
or U1783 (N_1783,N_987,N_753);
and U1784 (N_1784,N_371,N_609);
xnor U1785 (N_1785,N_666,N_565);
nand U1786 (N_1786,N_699,N_528);
nand U1787 (N_1787,N_487,N_827);
or U1788 (N_1788,N_105,N_360);
or U1789 (N_1789,N_517,N_515);
and U1790 (N_1790,N_973,N_592);
and U1791 (N_1791,N_230,N_998);
nand U1792 (N_1792,N_92,N_683);
nand U1793 (N_1793,N_455,N_972);
or U1794 (N_1794,N_491,N_28);
and U1795 (N_1795,N_719,N_842);
nand U1796 (N_1796,N_149,N_366);
nor U1797 (N_1797,N_750,N_966);
nor U1798 (N_1798,N_328,N_233);
and U1799 (N_1799,N_13,N_104);
or U1800 (N_1800,N_925,N_118);
and U1801 (N_1801,N_883,N_52);
nor U1802 (N_1802,N_668,N_926);
nor U1803 (N_1803,N_87,N_4);
or U1804 (N_1804,N_91,N_531);
nand U1805 (N_1805,N_996,N_787);
and U1806 (N_1806,N_348,N_375);
nand U1807 (N_1807,N_243,N_136);
nor U1808 (N_1808,N_859,N_597);
or U1809 (N_1809,N_4,N_892);
or U1810 (N_1810,N_337,N_949);
nor U1811 (N_1811,N_560,N_0);
or U1812 (N_1812,N_71,N_841);
nand U1813 (N_1813,N_303,N_906);
nor U1814 (N_1814,N_807,N_901);
nand U1815 (N_1815,N_659,N_507);
nor U1816 (N_1816,N_780,N_71);
and U1817 (N_1817,N_702,N_666);
nor U1818 (N_1818,N_550,N_964);
nor U1819 (N_1819,N_305,N_658);
nand U1820 (N_1820,N_531,N_449);
or U1821 (N_1821,N_843,N_376);
nand U1822 (N_1822,N_991,N_394);
and U1823 (N_1823,N_370,N_166);
nand U1824 (N_1824,N_352,N_530);
or U1825 (N_1825,N_834,N_251);
or U1826 (N_1826,N_84,N_186);
nand U1827 (N_1827,N_8,N_322);
or U1828 (N_1828,N_374,N_822);
nor U1829 (N_1829,N_385,N_36);
nand U1830 (N_1830,N_823,N_196);
nand U1831 (N_1831,N_848,N_517);
and U1832 (N_1832,N_146,N_267);
nand U1833 (N_1833,N_163,N_187);
and U1834 (N_1834,N_106,N_287);
nand U1835 (N_1835,N_756,N_327);
nand U1836 (N_1836,N_40,N_768);
and U1837 (N_1837,N_990,N_193);
nand U1838 (N_1838,N_45,N_344);
or U1839 (N_1839,N_456,N_322);
and U1840 (N_1840,N_165,N_115);
nor U1841 (N_1841,N_392,N_230);
and U1842 (N_1842,N_385,N_111);
nor U1843 (N_1843,N_856,N_979);
nor U1844 (N_1844,N_810,N_284);
nand U1845 (N_1845,N_532,N_338);
or U1846 (N_1846,N_130,N_35);
and U1847 (N_1847,N_615,N_676);
nand U1848 (N_1848,N_65,N_565);
nand U1849 (N_1849,N_898,N_856);
nor U1850 (N_1850,N_578,N_571);
nand U1851 (N_1851,N_792,N_959);
or U1852 (N_1852,N_318,N_719);
or U1853 (N_1853,N_670,N_582);
nand U1854 (N_1854,N_540,N_248);
nand U1855 (N_1855,N_290,N_898);
or U1856 (N_1856,N_20,N_403);
and U1857 (N_1857,N_176,N_462);
nor U1858 (N_1858,N_167,N_991);
nor U1859 (N_1859,N_778,N_369);
and U1860 (N_1860,N_402,N_259);
or U1861 (N_1861,N_201,N_140);
nand U1862 (N_1862,N_466,N_821);
nor U1863 (N_1863,N_21,N_860);
nor U1864 (N_1864,N_77,N_920);
nand U1865 (N_1865,N_145,N_849);
nor U1866 (N_1866,N_206,N_827);
nand U1867 (N_1867,N_315,N_6);
or U1868 (N_1868,N_976,N_317);
nand U1869 (N_1869,N_156,N_388);
nand U1870 (N_1870,N_466,N_120);
or U1871 (N_1871,N_61,N_586);
and U1872 (N_1872,N_467,N_775);
nor U1873 (N_1873,N_922,N_479);
nor U1874 (N_1874,N_601,N_82);
and U1875 (N_1875,N_977,N_403);
nand U1876 (N_1876,N_375,N_792);
nand U1877 (N_1877,N_962,N_902);
nand U1878 (N_1878,N_442,N_671);
nand U1879 (N_1879,N_820,N_232);
nand U1880 (N_1880,N_631,N_728);
nor U1881 (N_1881,N_592,N_142);
nand U1882 (N_1882,N_372,N_342);
nand U1883 (N_1883,N_851,N_175);
nand U1884 (N_1884,N_169,N_900);
nor U1885 (N_1885,N_515,N_966);
nand U1886 (N_1886,N_745,N_578);
and U1887 (N_1887,N_456,N_631);
nor U1888 (N_1888,N_718,N_918);
and U1889 (N_1889,N_852,N_903);
nor U1890 (N_1890,N_164,N_765);
or U1891 (N_1891,N_423,N_90);
nand U1892 (N_1892,N_663,N_67);
and U1893 (N_1893,N_661,N_493);
nand U1894 (N_1894,N_729,N_746);
and U1895 (N_1895,N_107,N_239);
or U1896 (N_1896,N_519,N_15);
and U1897 (N_1897,N_198,N_266);
nor U1898 (N_1898,N_50,N_788);
and U1899 (N_1899,N_228,N_513);
nor U1900 (N_1900,N_424,N_100);
nand U1901 (N_1901,N_619,N_138);
or U1902 (N_1902,N_854,N_380);
nor U1903 (N_1903,N_757,N_78);
and U1904 (N_1904,N_423,N_573);
nor U1905 (N_1905,N_70,N_858);
nor U1906 (N_1906,N_502,N_527);
nand U1907 (N_1907,N_594,N_937);
and U1908 (N_1908,N_239,N_225);
and U1909 (N_1909,N_918,N_638);
and U1910 (N_1910,N_112,N_821);
nor U1911 (N_1911,N_221,N_92);
and U1912 (N_1912,N_633,N_119);
and U1913 (N_1913,N_357,N_496);
nand U1914 (N_1914,N_245,N_153);
nand U1915 (N_1915,N_572,N_577);
and U1916 (N_1916,N_85,N_451);
and U1917 (N_1917,N_745,N_968);
nor U1918 (N_1918,N_143,N_796);
or U1919 (N_1919,N_872,N_30);
or U1920 (N_1920,N_686,N_270);
nand U1921 (N_1921,N_82,N_42);
and U1922 (N_1922,N_847,N_995);
nor U1923 (N_1923,N_807,N_727);
and U1924 (N_1924,N_500,N_666);
and U1925 (N_1925,N_370,N_986);
nand U1926 (N_1926,N_305,N_864);
nor U1927 (N_1927,N_966,N_764);
and U1928 (N_1928,N_357,N_220);
nor U1929 (N_1929,N_363,N_770);
nand U1930 (N_1930,N_395,N_819);
nand U1931 (N_1931,N_555,N_888);
and U1932 (N_1932,N_622,N_215);
or U1933 (N_1933,N_929,N_863);
and U1934 (N_1934,N_142,N_753);
nand U1935 (N_1935,N_424,N_867);
or U1936 (N_1936,N_706,N_199);
and U1937 (N_1937,N_24,N_141);
or U1938 (N_1938,N_748,N_459);
nor U1939 (N_1939,N_697,N_884);
nor U1940 (N_1940,N_111,N_223);
and U1941 (N_1941,N_860,N_410);
xor U1942 (N_1942,N_183,N_302);
or U1943 (N_1943,N_732,N_214);
nand U1944 (N_1944,N_27,N_735);
xor U1945 (N_1945,N_411,N_227);
or U1946 (N_1946,N_626,N_61);
or U1947 (N_1947,N_997,N_682);
nor U1948 (N_1948,N_711,N_406);
nand U1949 (N_1949,N_454,N_331);
and U1950 (N_1950,N_125,N_963);
and U1951 (N_1951,N_231,N_726);
or U1952 (N_1952,N_718,N_514);
nand U1953 (N_1953,N_562,N_512);
and U1954 (N_1954,N_896,N_491);
or U1955 (N_1955,N_144,N_541);
nor U1956 (N_1956,N_754,N_418);
nor U1957 (N_1957,N_588,N_982);
or U1958 (N_1958,N_490,N_133);
nor U1959 (N_1959,N_46,N_877);
and U1960 (N_1960,N_472,N_56);
or U1961 (N_1961,N_898,N_121);
or U1962 (N_1962,N_485,N_334);
nor U1963 (N_1963,N_17,N_223);
and U1964 (N_1964,N_319,N_992);
nand U1965 (N_1965,N_151,N_996);
nor U1966 (N_1966,N_976,N_943);
and U1967 (N_1967,N_226,N_376);
and U1968 (N_1968,N_493,N_279);
nand U1969 (N_1969,N_510,N_76);
nor U1970 (N_1970,N_325,N_632);
or U1971 (N_1971,N_513,N_245);
nor U1972 (N_1972,N_616,N_767);
nand U1973 (N_1973,N_84,N_666);
or U1974 (N_1974,N_138,N_463);
nand U1975 (N_1975,N_908,N_650);
and U1976 (N_1976,N_164,N_445);
nand U1977 (N_1977,N_321,N_635);
or U1978 (N_1978,N_736,N_342);
or U1979 (N_1979,N_124,N_240);
and U1980 (N_1980,N_824,N_831);
nor U1981 (N_1981,N_78,N_775);
and U1982 (N_1982,N_428,N_225);
nor U1983 (N_1983,N_346,N_429);
nand U1984 (N_1984,N_566,N_392);
xnor U1985 (N_1985,N_910,N_566);
nor U1986 (N_1986,N_496,N_133);
nand U1987 (N_1987,N_176,N_818);
or U1988 (N_1988,N_356,N_978);
and U1989 (N_1989,N_839,N_895);
or U1990 (N_1990,N_81,N_709);
or U1991 (N_1991,N_483,N_83);
nor U1992 (N_1992,N_338,N_363);
nand U1993 (N_1993,N_867,N_210);
and U1994 (N_1994,N_408,N_262);
nand U1995 (N_1995,N_597,N_234);
nand U1996 (N_1996,N_201,N_547);
and U1997 (N_1997,N_812,N_4);
nor U1998 (N_1998,N_91,N_496);
nand U1999 (N_1999,N_740,N_20);
and U2000 (N_2000,N_1863,N_1989);
or U2001 (N_2001,N_1488,N_1802);
xor U2002 (N_2002,N_1729,N_1569);
or U2003 (N_2003,N_1107,N_1462);
nand U2004 (N_2004,N_1810,N_1111);
nor U2005 (N_2005,N_1927,N_1380);
nor U2006 (N_2006,N_1419,N_1495);
nor U2007 (N_2007,N_1946,N_1526);
and U2008 (N_2008,N_1990,N_1058);
and U2009 (N_2009,N_1013,N_1698);
or U2010 (N_2010,N_1327,N_1391);
nand U2011 (N_2011,N_1922,N_1967);
and U2012 (N_2012,N_1828,N_1935);
nor U2013 (N_2013,N_1708,N_1601);
and U2014 (N_2014,N_1904,N_1038);
and U2015 (N_2015,N_1814,N_1332);
and U2016 (N_2016,N_1934,N_1352);
nand U2017 (N_2017,N_1424,N_1580);
nor U2018 (N_2018,N_1079,N_1021);
nor U2019 (N_2019,N_1543,N_1545);
nand U2020 (N_2020,N_1217,N_1684);
nor U2021 (N_2021,N_1808,N_1242);
and U2022 (N_2022,N_1821,N_1225);
or U2023 (N_2023,N_1534,N_1407);
nand U2024 (N_2024,N_1344,N_1224);
or U2025 (N_2025,N_1266,N_1248);
and U2026 (N_2026,N_1194,N_1265);
or U2027 (N_2027,N_1109,N_1435);
nand U2028 (N_2028,N_1535,N_1650);
nor U2029 (N_2029,N_1176,N_1649);
or U2030 (N_2030,N_1900,N_1908);
nand U2031 (N_2031,N_1532,N_1511);
nand U2032 (N_2032,N_1491,N_1556);
nand U2033 (N_2033,N_1337,N_1733);
and U2034 (N_2034,N_1849,N_1606);
nand U2035 (N_2035,N_1884,N_1370);
nand U2036 (N_2036,N_1146,N_1104);
and U2037 (N_2037,N_1529,N_1644);
or U2038 (N_2038,N_1091,N_1151);
and U2039 (N_2039,N_1402,N_1240);
nor U2040 (N_2040,N_1972,N_1894);
and U2041 (N_2041,N_1289,N_1539);
or U2042 (N_2042,N_1164,N_1952);
or U2043 (N_2043,N_1641,N_1899);
and U2044 (N_2044,N_1768,N_1173);
or U2045 (N_2045,N_1062,N_1185);
or U2046 (N_2046,N_1498,N_1076);
and U2047 (N_2047,N_1216,N_1983);
nor U2048 (N_2048,N_1541,N_1027);
nand U2049 (N_2049,N_1203,N_1788);
nor U2050 (N_2050,N_1367,N_1865);
nor U2051 (N_2051,N_1519,N_1279);
nand U2052 (N_2052,N_1818,N_1537);
nand U2053 (N_2053,N_1234,N_1709);
nor U2054 (N_2054,N_1453,N_1060);
nand U2055 (N_2055,N_1065,N_1917);
and U2056 (N_2056,N_1041,N_1964);
nor U2057 (N_2057,N_1014,N_1283);
and U2058 (N_2058,N_1315,N_1158);
and U2059 (N_2059,N_1017,N_1906);
and U2060 (N_2060,N_1575,N_1735);
nand U2061 (N_2061,N_1571,N_1809);
and U2062 (N_2062,N_1770,N_1582);
nor U2063 (N_2063,N_1813,N_1343);
or U2064 (N_2064,N_1039,N_1138);
nand U2065 (N_2065,N_1492,N_1730);
or U2066 (N_2066,N_1516,N_1154);
nand U2067 (N_2067,N_1219,N_1475);
nand U2068 (N_2068,N_1574,N_1879);
nand U2069 (N_2069,N_1531,N_1565);
nor U2070 (N_2070,N_1004,N_1755);
nor U2071 (N_2071,N_1218,N_1783);
nor U2072 (N_2072,N_1763,N_1386);
nand U2073 (N_2073,N_1795,N_1699);
and U2074 (N_2074,N_1888,N_1136);
or U2075 (N_2075,N_1237,N_1794);
and U2076 (N_2076,N_1336,N_1489);
nor U2077 (N_2077,N_1263,N_1406);
nand U2078 (N_2078,N_1920,N_1375);
or U2079 (N_2079,N_1259,N_1165);
nor U2080 (N_2080,N_1521,N_1055);
nor U2081 (N_2081,N_1069,N_1561);
or U2082 (N_2082,N_1328,N_1673);
or U2083 (N_2083,N_1648,N_1550);
and U2084 (N_2084,N_1985,N_1803);
or U2085 (N_2085,N_1468,N_1448);
and U2086 (N_2086,N_1595,N_1287);
or U2087 (N_2087,N_1000,N_1705);
nor U2088 (N_2088,N_1348,N_1782);
or U2089 (N_2089,N_1500,N_1001);
nor U2090 (N_2090,N_1999,N_1536);
nor U2091 (N_2091,N_1241,N_1126);
or U2092 (N_2092,N_1396,N_1321);
or U2093 (N_2093,N_1702,N_1078);
and U2094 (N_2094,N_1867,N_1118);
and U2095 (N_2095,N_1411,N_1602);
or U2096 (N_2096,N_1307,N_1861);
or U2097 (N_2097,N_1198,N_1269);
nand U2098 (N_2098,N_1678,N_1008);
and U2099 (N_2099,N_1859,N_1638);
nor U2100 (N_2100,N_1098,N_1421);
or U2101 (N_2101,N_1450,N_1410);
or U2102 (N_2102,N_1817,N_1681);
or U2103 (N_2103,N_1778,N_1262);
and U2104 (N_2104,N_1258,N_1767);
nor U2105 (N_2105,N_1553,N_1851);
nand U2106 (N_2106,N_1656,N_1969);
nor U2107 (N_2107,N_1799,N_1339);
or U2108 (N_2108,N_1083,N_1680);
nand U2109 (N_2109,N_1953,N_1340);
and U2110 (N_2110,N_1011,N_1664);
or U2111 (N_2111,N_1622,N_1246);
or U2112 (N_2112,N_1806,N_1135);
or U2113 (N_2113,N_1432,N_1551);
or U2114 (N_2114,N_1254,N_1499);
and U2115 (N_2115,N_1272,N_1436);
nor U2116 (N_2116,N_1088,N_1192);
and U2117 (N_2117,N_1632,N_1179);
nor U2118 (N_2118,N_1189,N_1830);
nand U2119 (N_2119,N_1002,N_1071);
nand U2120 (N_2120,N_1092,N_1652);
or U2121 (N_2121,N_1190,N_1115);
and U2122 (N_2122,N_1170,N_1161);
or U2123 (N_2123,N_1626,N_1555);
and U2124 (N_2124,N_1019,N_1593);
or U2125 (N_2125,N_1048,N_1360);
and U2126 (N_2126,N_1764,N_1881);
nor U2127 (N_2127,N_1400,N_1522);
nor U2128 (N_2128,N_1777,N_1449);
and U2129 (N_2129,N_1268,N_1568);
and U2130 (N_2130,N_1987,N_1210);
nor U2131 (N_2131,N_1059,N_1581);
and U2132 (N_2132,N_1538,N_1501);
and U2133 (N_2133,N_1563,N_1931);
nand U2134 (N_2134,N_1653,N_1113);
nor U2135 (N_2135,N_1996,N_1253);
nor U2136 (N_2136,N_1719,N_1883);
or U2137 (N_2137,N_1527,N_1966);
nor U2138 (N_2138,N_1979,N_1822);
and U2139 (N_2139,N_1721,N_1372);
and U2140 (N_2140,N_1609,N_1611);
or U2141 (N_2141,N_1962,N_1137);
nor U2142 (N_2142,N_1308,N_1508);
nand U2143 (N_2143,N_1358,N_1270);
and U2144 (N_2144,N_1542,N_1383);
or U2145 (N_2145,N_1560,N_1666);
and U2146 (N_2146,N_1914,N_1096);
nand U2147 (N_2147,N_1081,N_1378);
and U2148 (N_2148,N_1629,N_1162);
nor U2149 (N_2149,N_1007,N_1064);
and U2150 (N_2150,N_1594,N_1376);
nand U2151 (N_2151,N_1752,N_1873);
or U2152 (N_2152,N_1141,N_1408);
and U2153 (N_2153,N_1322,N_1397);
or U2154 (N_2154,N_1211,N_1297);
and U2155 (N_2155,N_1919,N_1018);
or U2156 (N_2156,N_1477,N_1466);
and U2157 (N_2157,N_1356,N_1995);
and U2158 (N_2158,N_1988,N_1944);
and U2159 (N_2159,N_1936,N_1950);
nor U2160 (N_2160,N_1122,N_1195);
nand U2161 (N_2161,N_1621,N_1087);
and U2162 (N_2162,N_1547,N_1633);
nand U2163 (N_2163,N_1986,N_1613);
nand U2164 (N_2164,N_1033,N_1831);
or U2165 (N_2165,N_1452,N_1155);
and U2166 (N_2166,N_1331,N_1267);
nand U2167 (N_2167,N_1319,N_1774);
or U2168 (N_2168,N_1790,N_1746);
or U2169 (N_2169,N_1362,N_1816);
or U2170 (N_2170,N_1490,N_1020);
and U2171 (N_2171,N_1896,N_1024);
nor U2172 (N_2172,N_1932,N_1226);
nor U2173 (N_2173,N_1204,N_1695);
and U2174 (N_2174,N_1704,N_1393);
and U2175 (N_2175,N_1443,N_1685);
nor U2176 (N_2176,N_1618,N_1469);
nor U2177 (N_2177,N_1530,N_1892);
or U2178 (N_2178,N_1607,N_1583);
nand U2179 (N_2179,N_1288,N_1954);
nor U2180 (N_2180,N_1334,N_1876);
nor U2181 (N_2181,N_1635,N_1924);
nor U2182 (N_2182,N_1642,N_1025);
nand U2183 (N_2183,N_1026,N_1981);
or U2184 (N_2184,N_1423,N_1197);
nand U2185 (N_2185,N_1505,N_1199);
nor U2186 (N_2186,N_1674,N_1961);
and U2187 (N_2187,N_1409,N_1659);
nand U2188 (N_2188,N_1015,N_1303);
nand U2189 (N_2189,N_1619,N_1665);
nor U2190 (N_2190,N_1054,N_1751);
and U2191 (N_2191,N_1824,N_1416);
and U2192 (N_2192,N_1510,N_1335);
or U2193 (N_2193,N_1341,N_1683);
nand U2194 (N_2194,N_1460,N_1139);
nand U2195 (N_2195,N_1196,N_1067);
nand U2196 (N_2196,N_1291,N_1549);
or U2197 (N_2197,N_1320,N_1734);
and U2198 (N_2198,N_1057,N_1231);
nor U2199 (N_2199,N_1509,N_1933);
nand U2200 (N_2200,N_1903,N_1564);
nor U2201 (N_2201,N_1294,N_1446);
xnor U2202 (N_2202,N_1119,N_1840);
or U2203 (N_2203,N_1412,N_1201);
and U2204 (N_2204,N_1731,N_1589);
nor U2205 (N_2205,N_1779,N_1086);
and U2206 (N_2206,N_1784,N_1902);
and U2207 (N_2207,N_1689,N_1235);
nand U2208 (N_2208,N_1608,N_1796);
and U2209 (N_2209,N_1804,N_1174);
nand U2210 (N_2210,N_1703,N_1675);
nand U2211 (N_2211,N_1243,N_1117);
nor U2212 (N_2212,N_1373,N_1006);
or U2213 (N_2213,N_1839,N_1780);
nand U2214 (N_2214,N_1732,N_1129);
or U2215 (N_2215,N_1982,N_1425);
nor U2216 (N_2216,N_1364,N_1725);
nor U2217 (N_2217,N_1692,N_1302);
nand U2218 (N_2218,N_1942,N_1044);
nor U2219 (N_2219,N_1515,N_1728);
or U2220 (N_2220,N_1377,N_1760);
nand U2221 (N_2221,N_1434,N_1891);
nand U2222 (N_2222,N_1325,N_1132);
nand U2223 (N_2223,N_1750,N_1353);
and U2224 (N_2224,N_1853,N_1528);
or U2225 (N_2225,N_1395,N_1120);
or U2226 (N_2226,N_1739,N_1414);
nor U2227 (N_2227,N_1366,N_1191);
and U2228 (N_2228,N_1820,N_1326);
or U2229 (N_2229,N_1562,N_1646);
nand U2230 (N_2230,N_1010,N_1514);
nor U2231 (N_2231,N_1843,N_1206);
and U2232 (N_2232,N_1965,N_1623);
nand U2233 (N_2233,N_1103,N_1212);
nand U2234 (N_2234,N_1286,N_1984);
and U2235 (N_2235,N_1754,N_1456);
nand U2236 (N_2236,N_1833,N_1168);
xnor U2237 (N_2237,N_1229,N_1832);
nand U2238 (N_2238,N_1016,N_1451);
and U2239 (N_2239,N_1744,N_1005);
nor U2240 (N_2240,N_1504,N_1338);
nand U2241 (N_2241,N_1072,N_1304);
nor U2242 (N_2242,N_1558,N_1052);
nand U2243 (N_2243,N_1874,N_1455);
nand U2244 (N_2244,N_1357,N_1945);
or U2245 (N_2245,N_1186,N_1647);
nor U2246 (N_2246,N_1958,N_1716);
nand U2247 (N_2247,N_1478,N_1506);
or U2248 (N_2248,N_1715,N_1856);
or U2249 (N_2249,N_1368,N_1256);
or U2250 (N_2250,N_1871,N_1483);
or U2251 (N_2251,N_1815,N_1085);
nand U2252 (N_2252,N_1690,N_1973);
or U2253 (N_2253,N_1793,N_1880);
nand U2254 (N_2254,N_1890,N_1187);
or U2255 (N_2255,N_1740,N_1925);
nand U2256 (N_2256,N_1612,N_1857);
and U2257 (N_2257,N_1912,N_1003);
and U2258 (N_2258,N_1707,N_1390);
xor U2259 (N_2259,N_1940,N_1379);
nor U2260 (N_2260,N_1930,N_1476);
or U2261 (N_2261,N_1605,N_1157);
or U2262 (N_2262,N_1756,N_1587);
and U2263 (N_2263,N_1472,N_1762);
or U2264 (N_2264,N_1603,N_1741);
nor U2265 (N_2265,N_1918,N_1236);
nand U2266 (N_2266,N_1614,N_1854);
nand U2267 (N_2267,N_1722,N_1928);
or U2268 (N_2268,N_1080,N_1503);
and U2269 (N_2269,N_1239,N_1963);
nor U2270 (N_2270,N_1670,N_1260);
nand U2271 (N_2271,N_1032,N_1047);
nand U2272 (N_2272,N_1461,N_1300);
or U2273 (N_2273,N_1130,N_1893);
nand U2274 (N_2274,N_1948,N_1342);
and U2275 (N_2275,N_1482,N_1977);
nand U2276 (N_2276,N_1693,N_1566);
nor U2277 (N_2277,N_1180,N_1588);
and U2278 (N_2278,N_1655,N_1222);
nand U2279 (N_2279,N_1420,N_1970);
or U2280 (N_2280,N_1617,N_1207);
nand U2281 (N_2281,N_1089,N_1264);
or U2282 (N_2282,N_1306,N_1860);
or U2283 (N_2283,N_1616,N_1238);
and U2284 (N_2284,N_1457,N_1147);
and U2285 (N_2285,N_1745,N_1040);
or U2286 (N_2286,N_1374,N_1428);
and U2287 (N_2287,N_1208,N_1398);
nor U2288 (N_2288,N_1776,N_1748);
nor U2289 (N_2289,N_1862,N_1567);
nand U2290 (N_2290,N_1227,N_1710);
nor U2291 (N_2291,N_1724,N_1333);
or U2292 (N_2292,N_1166,N_1718);
nand U2293 (N_2293,N_1034,N_1634);
or U2294 (N_2294,N_1706,N_1167);
nand U2295 (N_2295,N_1929,N_1389);
nor U2296 (N_2296,N_1172,N_1672);
nor U2297 (N_2297,N_1765,N_1388);
nand U2298 (N_2298,N_1074,N_1579);
nor U2299 (N_2299,N_1669,N_1687);
nor U2300 (N_2300,N_1313,N_1882);
nor U2301 (N_2301,N_1145,N_1769);
or U2302 (N_2302,N_1415,N_1175);
nor U2303 (N_2303,N_1597,N_1941);
nor U2304 (N_2304,N_1916,N_1467);
or U2305 (N_2305,N_1781,N_1417);
or U2306 (N_2306,N_1697,N_1772);
nor U2307 (N_2307,N_1823,N_1548);
nand U2308 (N_2308,N_1960,N_1838);
or U2309 (N_2309,N_1178,N_1329);
and U2310 (N_2310,N_1599,N_1310);
or U2311 (N_2311,N_1035,N_1056);
and U2312 (N_2312,N_1975,N_1330);
or U2313 (N_2313,N_1992,N_1834);
or U2314 (N_2314,N_1394,N_1068);
nor U2315 (N_2315,N_1430,N_1586);
and U2316 (N_2316,N_1022,N_1598);
nor U2317 (N_2317,N_1223,N_1789);
and U2318 (N_2318,N_1361,N_1825);
nand U2319 (N_2319,N_1093,N_1512);
nor U2320 (N_2320,N_1464,N_1480);
nand U2321 (N_2321,N_1029,N_1872);
and U2322 (N_2322,N_1524,N_1181);
nand U2323 (N_2323,N_1540,N_1387);
and U2324 (N_2324,N_1371,N_1819);
nor U2325 (N_2325,N_1807,N_1976);
nor U2326 (N_2326,N_1791,N_1949);
nor U2327 (N_2327,N_1637,N_1228);
nor U2328 (N_2328,N_1845,N_1887);
or U2329 (N_2329,N_1926,N_1148);
and U2330 (N_2330,N_1422,N_1713);
nand U2331 (N_2331,N_1484,N_1131);
or U2332 (N_2332,N_1101,N_1518);
and U2333 (N_2333,N_1921,N_1077);
or U2334 (N_2334,N_1444,N_1473);
nor U2335 (N_2335,N_1114,N_1786);
nor U2336 (N_2336,N_1281,N_1668);
or U2337 (N_2337,N_1864,N_1938);
nand U2338 (N_2338,N_1533,N_1787);
nand U2339 (N_2339,N_1075,N_1761);
and U2340 (N_2340,N_1110,N_1736);
and U2341 (N_2341,N_1513,N_1826);
nand U2342 (N_2342,N_1991,N_1610);
and U2343 (N_2343,N_1458,N_1413);
nand U2344 (N_2344,N_1280,N_1905);
nor U2345 (N_2345,N_1030,N_1213);
nand U2346 (N_2346,N_1317,N_1978);
or U2347 (N_2347,N_1250,N_1663);
or U2348 (N_2348,N_1233,N_1577);
or U2349 (N_2349,N_1143,N_1723);
nand U2350 (N_2350,N_1277,N_1720);
nor U2351 (N_2351,N_1994,N_1028);
nor U2352 (N_2352,N_1691,N_1800);
nor U2353 (N_2353,N_1214,N_1046);
or U2354 (N_2354,N_1053,N_1645);
nor U2355 (N_2355,N_1700,N_1576);
or U2356 (N_2356,N_1878,N_1701);
nand U2357 (N_2357,N_1842,N_1318);
nor U2358 (N_2358,N_1600,N_1276);
and U2359 (N_2359,N_1403,N_1205);
nor U2360 (N_2360,N_1230,N_1998);
nor U2361 (N_2361,N_1497,N_1662);
and U2362 (N_2362,N_1439,N_1116);
and U2363 (N_2363,N_1347,N_1712);
nand U2364 (N_2364,N_1743,N_1679);
nand U2365 (N_2365,N_1349,N_1292);
nand U2366 (N_2366,N_1023,N_1628);
or U2367 (N_2367,N_1625,N_1285);
nand U2368 (N_2368,N_1660,N_1084);
nor U2369 (N_2369,N_1596,N_1636);
nor U2370 (N_2370,N_1177,N_1045);
nor U2371 (N_2371,N_1278,N_1445);
nand U2372 (N_2372,N_1271,N_1974);
and U2373 (N_2373,N_1061,N_1951);
and U2374 (N_2374,N_1099,N_1573);
nand U2375 (N_2375,N_1688,N_1247);
nand U2376 (N_2376,N_1639,N_1037);
nand U2377 (N_2377,N_1726,N_1667);
or U2378 (N_2378,N_1171,N_1711);
and U2379 (N_2379,N_1036,N_1812);
xor U2380 (N_2380,N_1836,N_1886);
nand U2381 (N_2381,N_1133,N_1156);
nor U2382 (N_2382,N_1121,N_1897);
or U2383 (N_2383,N_1252,N_1870);
or U2384 (N_2384,N_1980,N_1293);
nand U2385 (N_2385,N_1947,N_1907);
or U2386 (N_2386,N_1163,N_1682);
nor U2387 (N_2387,N_1442,N_1971);
nor U2388 (N_2388,N_1792,N_1844);
nand U2389 (N_2389,N_1221,N_1249);
nand U2390 (N_2390,N_1671,N_1959);
nor U2391 (N_2391,N_1183,N_1624);
xor U2392 (N_2392,N_1801,N_1943);
xnor U2393 (N_2393,N_1100,N_1798);
nand U2394 (N_2394,N_1654,N_1848);
nand U2395 (N_2395,N_1677,N_1841);
xor U2396 (N_2396,N_1128,N_1365);
nand U2397 (N_2397,N_1479,N_1431);
or U2398 (N_2398,N_1717,N_1570);
or U2399 (N_2399,N_1354,N_1852);
nor U2400 (N_2400,N_1070,N_1351);
or U2401 (N_2401,N_1094,N_1050);
nor U2402 (N_2402,N_1591,N_1363);
nor U2403 (N_2403,N_1661,N_1160);
or U2404 (N_2404,N_1875,N_1866);
or U2405 (N_2405,N_1251,N_1284);
nand U2406 (N_2406,N_1232,N_1592);
nand U2407 (N_2407,N_1359,N_1507);
and U2408 (N_2408,N_1889,N_1805);
and U2409 (N_2409,N_1405,N_1152);
nand U2410 (N_2410,N_1309,N_1485);
xor U2411 (N_2411,N_1384,N_1274);
nand U2412 (N_2412,N_1620,N_1073);
and U2413 (N_2413,N_1493,N_1847);
nand U2414 (N_2414,N_1440,N_1993);
nand U2415 (N_2415,N_1727,N_1631);
and U2416 (N_2416,N_1345,N_1911);
and U2417 (N_2417,N_1766,N_1049);
or U2418 (N_2418,N_1520,N_1324);
or U2419 (N_2419,N_1031,N_1149);
nand U2420 (N_2420,N_1494,N_1209);
nor U2421 (N_2421,N_1350,N_1296);
or U2422 (N_2422,N_1290,N_1282);
or U2423 (N_2423,N_1124,N_1082);
nor U2424 (N_2424,N_1441,N_1827);
nand U2425 (N_2425,N_1955,N_1846);
nand U2426 (N_2426,N_1640,N_1470);
or U2427 (N_2427,N_1261,N_1523);
or U2428 (N_2428,N_1202,N_1855);
nor U2429 (N_2429,N_1255,N_1454);
and U2430 (N_2430,N_1696,N_1355);
and U2431 (N_2431,N_1956,N_1502);
or U2432 (N_2432,N_1749,N_1418);
nand U2433 (N_2433,N_1051,N_1433);
nand U2434 (N_2434,N_1651,N_1627);
nand U2435 (N_2435,N_1630,N_1694);
and U2436 (N_2436,N_1142,N_1295);
or U2437 (N_2437,N_1182,N_1298);
nand U2438 (N_2438,N_1471,N_1275);
nand U2439 (N_2439,N_1399,N_1102);
nand U2440 (N_2440,N_1811,N_1898);
nor U2441 (N_2441,N_1200,N_1299);
and U2442 (N_2442,N_1369,N_1557);
or U2443 (N_2443,N_1381,N_1910);
or U2444 (N_2444,N_1244,N_1043);
nand U2445 (N_2445,N_1868,N_1753);
nand U2446 (N_2446,N_1643,N_1063);
nand U2447 (N_2447,N_1486,N_1447);
or U2448 (N_2448,N_1829,N_1106);
and U2449 (N_2449,N_1496,N_1042);
and U2450 (N_2450,N_1775,N_1346);
nor U2451 (N_2451,N_1937,N_1314);
and U2452 (N_2452,N_1184,N_1108);
nor U2453 (N_2453,N_1153,N_1127);
and U2454 (N_2454,N_1112,N_1915);
or U2455 (N_2455,N_1257,N_1487);
xnor U2456 (N_2456,N_1474,N_1968);
and U2457 (N_2457,N_1159,N_1150);
nor U2458 (N_2458,N_1615,N_1554);
nand U2459 (N_2459,N_1758,N_1438);
nand U2460 (N_2460,N_1997,N_1738);
nor U2461 (N_2461,N_1957,N_1714);
and U2462 (N_2462,N_1517,N_1797);
and U2463 (N_2463,N_1066,N_1188);
nand U2464 (N_2464,N_1559,N_1572);
nor U2465 (N_2465,N_1658,N_1125);
nor U2466 (N_2466,N_1095,N_1459);
or U2467 (N_2467,N_1463,N_1427);
and U2468 (N_2468,N_1546,N_1385);
and U2469 (N_2469,N_1437,N_1525);
or U2470 (N_2470,N_1305,N_1392);
or U2471 (N_2471,N_1465,N_1578);
nor U2472 (N_2472,N_1858,N_1301);
or U2473 (N_2473,N_1169,N_1747);
nor U2474 (N_2474,N_1771,N_1869);
nor U2475 (N_2475,N_1404,N_1757);
nor U2476 (N_2476,N_1123,N_1737);
or U2477 (N_2477,N_1676,N_1481);
or U2478 (N_2478,N_1316,N_1901);
nand U2479 (N_2479,N_1604,N_1837);
and U2480 (N_2480,N_1657,N_1913);
and U2481 (N_2481,N_1850,N_1090);
nor U2482 (N_2482,N_1590,N_1009);
nor U2483 (N_2483,N_1909,N_1877);
nand U2484 (N_2484,N_1785,N_1835);
nor U2485 (N_2485,N_1552,N_1895);
or U2486 (N_2486,N_1401,N_1585);
nor U2487 (N_2487,N_1885,N_1012);
or U2488 (N_2488,N_1245,N_1323);
nor U2489 (N_2489,N_1686,N_1429);
or U2490 (N_2490,N_1939,N_1144);
and U2491 (N_2491,N_1773,N_1193);
or U2492 (N_2492,N_1105,N_1220);
nor U2493 (N_2493,N_1273,N_1134);
and U2494 (N_2494,N_1544,N_1382);
nor U2495 (N_2495,N_1923,N_1742);
or U2496 (N_2496,N_1759,N_1215);
nor U2497 (N_2497,N_1426,N_1097);
nor U2498 (N_2498,N_1140,N_1311);
nand U2499 (N_2499,N_1312,N_1584);
nor U2500 (N_2500,N_1216,N_1601);
and U2501 (N_2501,N_1294,N_1988);
and U2502 (N_2502,N_1386,N_1903);
nand U2503 (N_2503,N_1696,N_1357);
and U2504 (N_2504,N_1017,N_1773);
nand U2505 (N_2505,N_1737,N_1686);
or U2506 (N_2506,N_1066,N_1200);
or U2507 (N_2507,N_1994,N_1562);
and U2508 (N_2508,N_1566,N_1766);
xor U2509 (N_2509,N_1099,N_1095);
or U2510 (N_2510,N_1414,N_1736);
nor U2511 (N_2511,N_1789,N_1388);
and U2512 (N_2512,N_1585,N_1539);
and U2513 (N_2513,N_1811,N_1275);
and U2514 (N_2514,N_1145,N_1328);
nand U2515 (N_2515,N_1402,N_1374);
nor U2516 (N_2516,N_1443,N_1491);
or U2517 (N_2517,N_1883,N_1746);
nand U2518 (N_2518,N_1876,N_1102);
nor U2519 (N_2519,N_1472,N_1428);
nand U2520 (N_2520,N_1339,N_1546);
and U2521 (N_2521,N_1113,N_1802);
nand U2522 (N_2522,N_1963,N_1613);
or U2523 (N_2523,N_1209,N_1568);
and U2524 (N_2524,N_1913,N_1378);
and U2525 (N_2525,N_1648,N_1615);
or U2526 (N_2526,N_1547,N_1081);
nor U2527 (N_2527,N_1466,N_1903);
nand U2528 (N_2528,N_1176,N_1545);
or U2529 (N_2529,N_1857,N_1714);
and U2530 (N_2530,N_1811,N_1810);
nor U2531 (N_2531,N_1734,N_1375);
nor U2532 (N_2532,N_1375,N_1788);
and U2533 (N_2533,N_1753,N_1785);
nand U2534 (N_2534,N_1786,N_1270);
or U2535 (N_2535,N_1075,N_1746);
nand U2536 (N_2536,N_1756,N_1422);
and U2537 (N_2537,N_1693,N_1885);
and U2538 (N_2538,N_1654,N_1629);
and U2539 (N_2539,N_1985,N_1756);
or U2540 (N_2540,N_1272,N_1038);
nand U2541 (N_2541,N_1303,N_1431);
nor U2542 (N_2542,N_1761,N_1134);
nand U2543 (N_2543,N_1973,N_1943);
and U2544 (N_2544,N_1050,N_1121);
or U2545 (N_2545,N_1488,N_1110);
and U2546 (N_2546,N_1106,N_1224);
or U2547 (N_2547,N_1392,N_1787);
or U2548 (N_2548,N_1159,N_1931);
nor U2549 (N_2549,N_1265,N_1599);
nor U2550 (N_2550,N_1331,N_1682);
nor U2551 (N_2551,N_1926,N_1853);
and U2552 (N_2552,N_1504,N_1866);
nand U2553 (N_2553,N_1956,N_1429);
nor U2554 (N_2554,N_1348,N_1005);
nand U2555 (N_2555,N_1572,N_1323);
or U2556 (N_2556,N_1273,N_1710);
or U2557 (N_2557,N_1496,N_1565);
nand U2558 (N_2558,N_1565,N_1144);
or U2559 (N_2559,N_1644,N_1258);
or U2560 (N_2560,N_1523,N_1075);
and U2561 (N_2561,N_1676,N_1764);
or U2562 (N_2562,N_1101,N_1644);
nor U2563 (N_2563,N_1753,N_1847);
and U2564 (N_2564,N_1275,N_1263);
nand U2565 (N_2565,N_1798,N_1394);
nand U2566 (N_2566,N_1477,N_1790);
and U2567 (N_2567,N_1917,N_1899);
nor U2568 (N_2568,N_1386,N_1981);
nor U2569 (N_2569,N_1864,N_1155);
or U2570 (N_2570,N_1885,N_1830);
and U2571 (N_2571,N_1286,N_1066);
and U2572 (N_2572,N_1746,N_1318);
or U2573 (N_2573,N_1272,N_1711);
or U2574 (N_2574,N_1019,N_1135);
and U2575 (N_2575,N_1800,N_1861);
and U2576 (N_2576,N_1922,N_1416);
nand U2577 (N_2577,N_1285,N_1295);
and U2578 (N_2578,N_1814,N_1378);
and U2579 (N_2579,N_1196,N_1303);
or U2580 (N_2580,N_1304,N_1919);
or U2581 (N_2581,N_1909,N_1840);
or U2582 (N_2582,N_1737,N_1033);
nand U2583 (N_2583,N_1400,N_1095);
or U2584 (N_2584,N_1019,N_1182);
nand U2585 (N_2585,N_1515,N_1859);
or U2586 (N_2586,N_1154,N_1893);
and U2587 (N_2587,N_1936,N_1998);
nand U2588 (N_2588,N_1486,N_1949);
and U2589 (N_2589,N_1529,N_1025);
nor U2590 (N_2590,N_1948,N_1156);
or U2591 (N_2591,N_1475,N_1098);
or U2592 (N_2592,N_1975,N_1752);
or U2593 (N_2593,N_1279,N_1362);
and U2594 (N_2594,N_1662,N_1706);
or U2595 (N_2595,N_1720,N_1545);
nor U2596 (N_2596,N_1727,N_1217);
or U2597 (N_2597,N_1166,N_1334);
or U2598 (N_2598,N_1074,N_1278);
or U2599 (N_2599,N_1088,N_1437);
nand U2600 (N_2600,N_1120,N_1668);
or U2601 (N_2601,N_1381,N_1925);
or U2602 (N_2602,N_1703,N_1779);
and U2603 (N_2603,N_1576,N_1346);
and U2604 (N_2604,N_1295,N_1181);
nor U2605 (N_2605,N_1339,N_1911);
nor U2606 (N_2606,N_1713,N_1753);
nor U2607 (N_2607,N_1096,N_1137);
xnor U2608 (N_2608,N_1057,N_1175);
nor U2609 (N_2609,N_1893,N_1737);
and U2610 (N_2610,N_1876,N_1054);
and U2611 (N_2611,N_1297,N_1183);
nand U2612 (N_2612,N_1739,N_1442);
nor U2613 (N_2613,N_1177,N_1779);
or U2614 (N_2614,N_1610,N_1770);
or U2615 (N_2615,N_1810,N_1073);
nor U2616 (N_2616,N_1373,N_1859);
nor U2617 (N_2617,N_1856,N_1435);
nand U2618 (N_2618,N_1410,N_1721);
or U2619 (N_2619,N_1503,N_1604);
and U2620 (N_2620,N_1985,N_1032);
or U2621 (N_2621,N_1267,N_1099);
nor U2622 (N_2622,N_1292,N_1282);
and U2623 (N_2623,N_1803,N_1834);
nor U2624 (N_2624,N_1248,N_1419);
or U2625 (N_2625,N_1170,N_1515);
xor U2626 (N_2626,N_1255,N_1844);
nand U2627 (N_2627,N_1954,N_1232);
and U2628 (N_2628,N_1244,N_1458);
and U2629 (N_2629,N_1901,N_1143);
or U2630 (N_2630,N_1557,N_1317);
nand U2631 (N_2631,N_1493,N_1383);
and U2632 (N_2632,N_1787,N_1068);
and U2633 (N_2633,N_1687,N_1064);
and U2634 (N_2634,N_1946,N_1007);
nand U2635 (N_2635,N_1478,N_1955);
or U2636 (N_2636,N_1740,N_1703);
nand U2637 (N_2637,N_1831,N_1447);
or U2638 (N_2638,N_1895,N_1340);
and U2639 (N_2639,N_1296,N_1061);
nand U2640 (N_2640,N_1066,N_1765);
nor U2641 (N_2641,N_1056,N_1091);
or U2642 (N_2642,N_1019,N_1860);
nor U2643 (N_2643,N_1277,N_1991);
and U2644 (N_2644,N_1832,N_1180);
nor U2645 (N_2645,N_1365,N_1966);
and U2646 (N_2646,N_1310,N_1894);
and U2647 (N_2647,N_1761,N_1250);
nor U2648 (N_2648,N_1683,N_1372);
nand U2649 (N_2649,N_1909,N_1815);
nor U2650 (N_2650,N_1505,N_1511);
nor U2651 (N_2651,N_1402,N_1406);
nand U2652 (N_2652,N_1138,N_1282);
nand U2653 (N_2653,N_1270,N_1770);
or U2654 (N_2654,N_1487,N_1701);
nand U2655 (N_2655,N_1538,N_1181);
and U2656 (N_2656,N_1481,N_1082);
and U2657 (N_2657,N_1374,N_1743);
or U2658 (N_2658,N_1512,N_1635);
and U2659 (N_2659,N_1616,N_1683);
or U2660 (N_2660,N_1896,N_1370);
or U2661 (N_2661,N_1039,N_1803);
and U2662 (N_2662,N_1170,N_1273);
or U2663 (N_2663,N_1806,N_1604);
or U2664 (N_2664,N_1699,N_1638);
xor U2665 (N_2665,N_1309,N_1211);
nand U2666 (N_2666,N_1017,N_1320);
nor U2667 (N_2667,N_1706,N_1542);
or U2668 (N_2668,N_1452,N_1658);
or U2669 (N_2669,N_1459,N_1975);
or U2670 (N_2670,N_1034,N_1383);
nor U2671 (N_2671,N_1274,N_1927);
nand U2672 (N_2672,N_1990,N_1137);
or U2673 (N_2673,N_1141,N_1136);
and U2674 (N_2674,N_1792,N_1319);
and U2675 (N_2675,N_1011,N_1305);
and U2676 (N_2676,N_1962,N_1690);
and U2677 (N_2677,N_1940,N_1777);
nor U2678 (N_2678,N_1453,N_1096);
nor U2679 (N_2679,N_1545,N_1171);
nor U2680 (N_2680,N_1235,N_1546);
nor U2681 (N_2681,N_1451,N_1773);
or U2682 (N_2682,N_1671,N_1313);
or U2683 (N_2683,N_1157,N_1060);
or U2684 (N_2684,N_1944,N_1723);
and U2685 (N_2685,N_1171,N_1457);
or U2686 (N_2686,N_1355,N_1051);
and U2687 (N_2687,N_1520,N_1767);
nand U2688 (N_2688,N_1514,N_1500);
nand U2689 (N_2689,N_1183,N_1134);
and U2690 (N_2690,N_1955,N_1395);
or U2691 (N_2691,N_1548,N_1568);
nand U2692 (N_2692,N_1872,N_1374);
and U2693 (N_2693,N_1408,N_1325);
nand U2694 (N_2694,N_1175,N_1216);
or U2695 (N_2695,N_1544,N_1380);
nand U2696 (N_2696,N_1112,N_1888);
and U2697 (N_2697,N_1272,N_1213);
nor U2698 (N_2698,N_1224,N_1937);
and U2699 (N_2699,N_1310,N_1517);
and U2700 (N_2700,N_1190,N_1019);
and U2701 (N_2701,N_1070,N_1920);
and U2702 (N_2702,N_1143,N_1951);
nor U2703 (N_2703,N_1530,N_1876);
and U2704 (N_2704,N_1644,N_1462);
and U2705 (N_2705,N_1216,N_1669);
nand U2706 (N_2706,N_1621,N_1752);
nor U2707 (N_2707,N_1970,N_1818);
nand U2708 (N_2708,N_1101,N_1080);
nand U2709 (N_2709,N_1914,N_1544);
nand U2710 (N_2710,N_1400,N_1809);
nand U2711 (N_2711,N_1387,N_1613);
nand U2712 (N_2712,N_1242,N_1150);
or U2713 (N_2713,N_1000,N_1028);
or U2714 (N_2714,N_1406,N_1637);
nor U2715 (N_2715,N_1075,N_1481);
or U2716 (N_2716,N_1550,N_1024);
and U2717 (N_2717,N_1306,N_1321);
nand U2718 (N_2718,N_1581,N_1318);
and U2719 (N_2719,N_1407,N_1848);
nor U2720 (N_2720,N_1488,N_1316);
and U2721 (N_2721,N_1322,N_1551);
and U2722 (N_2722,N_1438,N_1647);
or U2723 (N_2723,N_1239,N_1428);
nand U2724 (N_2724,N_1628,N_1125);
and U2725 (N_2725,N_1194,N_1202);
nand U2726 (N_2726,N_1650,N_1669);
nor U2727 (N_2727,N_1490,N_1118);
or U2728 (N_2728,N_1980,N_1273);
nand U2729 (N_2729,N_1629,N_1754);
or U2730 (N_2730,N_1124,N_1698);
xnor U2731 (N_2731,N_1233,N_1602);
or U2732 (N_2732,N_1604,N_1489);
or U2733 (N_2733,N_1381,N_1267);
nand U2734 (N_2734,N_1856,N_1908);
or U2735 (N_2735,N_1363,N_1092);
nor U2736 (N_2736,N_1454,N_1527);
and U2737 (N_2737,N_1158,N_1894);
nor U2738 (N_2738,N_1113,N_1722);
nor U2739 (N_2739,N_1773,N_1599);
nand U2740 (N_2740,N_1059,N_1265);
xnor U2741 (N_2741,N_1200,N_1844);
and U2742 (N_2742,N_1719,N_1862);
or U2743 (N_2743,N_1838,N_1191);
nor U2744 (N_2744,N_1589,N_1452);
or U2745 (N_2745,N_1618,N_1620);
and U2746 (N_2746,N_1996,N_1274);
nand U2747 (N_2747,N_1783,N_1315);
nor U2748 (N_2748,N_1395,N_1223);
or U2749 (N_2749,N_1789,N_1042);
nand U2750 (N_2750,N_1025,N_1360);
or U2751 (N_2751,N_1794,N_1713);
nand U2752 (N_2752,N_1723,N_1774);
and U2753 (N_2753,N_1117,N_1823);
nand U2754 (N_2754,N_1566,N_1234);
nor U2755 (N_2755,N_1031,N_1187);
and U2756 (N_2756,N_1556,N_1625);
and U2757 (N_2757,N_1982,N_1693);
or U2758 (N_2758,N_1716,N_1808);
or U2759 (N_2759,N_1867,N_1295);
nand U2760 (N_2760,N_1086,N_1650);
and U2761 (N_2761,N_1597,N_1332);
nor U2762 (N_2762,N_1857,N_1828);
or U2763 (N_2763,N_1908,N_1969);
or U2764 (N_2764,N_1022,N_1724);
or U2765 (N_2765,N_1917,N_1155);
or U2766 (N_2766,N_1414,N_1726);
or U2767 (N_2767,N_1761,N_1366);
or U2768 (N_2768,N_1815,N_1798);
nor U2769 (N_2769,N_1601,N_1812);
nor U2770 (N_2770,N_1134,N_1330);
nor U2771 (N_2771,N_1087,N_1514);
nand U2772 (N_2772,N_1780,N_1649);
nand U2773 (N_2773,N_1462,N_1976);
and U2774 (N_2774,N_1152,N_1679);
or U2775 (N_2775,N_1894,N_1741);
nand U2776 (N_2776,N_1479,N_1460);
or U2777 (N_2777,N_1618,N_1772);
and U2778 (N_2778,N_1824,N_1751);
nand U2779 (N_2779,N_1818,N_1586);
nor U2780 (N_2780,N_1330,N_1970);
or U2781 (N_2781,N_1027,N_1515);
nand U2782 (N_2782,N_1454,N_1091);
nand U2783 (N_2783,N_1192,N_1969);
and U2784 (N_2784,N_1561,N_1711);
and U2785 (N_2785,N_1901,N_1831);
nand U2786 (N_2786,N_1571,N_1993);
nor U2787 (N_2787,N_1048,N_1470);
nand U2788 (N_2788,N_1405,N_1814);
nand U2789 (N_2789,N_1433,N_1104);
nor U2790 (N_2790,N_1595,N_1704);
nor U2791 (N_2791,N_1486,N_1851);
or U2792 (N_2792,N_1378,N_1237);
nand U2793 (N_2793,N_1594,N_1911);
nor U2794 (N_2794,N_1225,N_1444);
and U2795 (N_2795,N_1268,N_1813);
and U2796 (N_2796,N_1150,N_1037);
nor U2797 (N_2797,N_1541,N_1841);
or U2798 (N_2798,N_1918,N_1050);
nor U2799 (N_2799,N_1802,N_1447);
nand U2800 (N_2800,N_1441,N_1471);
nor U2801 (N_2801,N_1119,N_1633);
and U2802 (N_2802,N_1313,N_1990);
and U2803 (N_2803,N_1328,N_1131);
nor U2804 (N_2804,N_1342,N_1182);
or U2805 (N_2805,N_1205,N_1457);
and U2806 (N_2806,N_1044,N_1273);
or U2807 (N_2807,N_1499,N_1986);
or U2808 (N_2808,N_1001,N_1975);
and U2809 (N_2809,N_1669,N_1330);
nand U2810 (N_2810,N_1992,N_1959);
and U2811 (N_2811,N_1286,N_1192);
nor U2812 (N_2812,N_1752,N_1206);
nor U2813 (N_2813,N_1415,N_1347);
and U2814 (N_2814,N_1020,N_1441);
or U2815 (N_2815,N_1318,N_1120);
nor U2816 (N_2816,N_1973,N_1675);
and U2817 (N_2817,N_1349,N_1253);
and U2818 (N_2818,N_1611,N_1709);
and U2819 (N_2819,N_1558,N_1829);
and U2820 (N_2820,N_1348,N_1199);
nand U2821 (N_2821,N_1197,N_1230);
and U2822 (N_2822,N_1206,N_1647);
nand U2823 (N_2823,N_1406,N_1960);
or U2824 (N_2824,N_1915,N_1903);
or U2825 (N_2825,N_1084,N_1671);
or U2826 (N_2826,N_1413,N_1921);
and U2827 (N_2827,N_1745,N_1825);
nand U2828 (N_2828,N_1871,N_1649);
xnor U2829 (N_2829,N_1237,N_1627);
nand U2830 (N_2830,N_1061,N_1568);
nand U2831 (N_2831,N_1335,N_1731);
nand U2832 (N_2832,N_1552,N_1897);
or U2833 (N_2833,N_1390,N_1210);
and U2834 (N_2834,N_1211,N_1129);
and U2835 (N_2835,N_1666,N_1011);
nor U2836 (N_2836,N_1712,N_1572);
nor U2837 (N_2837,N_1550,N_1685);
nand U2838 (N_2838,N_1714,N_1683);
nor U2839 (N_2839,N_1221,N_1412);
and U2840 (N_2840,N_1088,N_1073);
nor U2841 (N_2841,N_1847,N_1499);
and U2842 (N_2842,N_1904,N_1208);
nor U2843 (N_2843,N_1842,N_1711);
nor U2844 (N_2844,N_1294,N_1310);
nor U2845 (N_2845,N_1765,N_1842);
or U2846 (N_2846,N_1764,N_1040);
xor U2847 (N_2847,N_1088,N_1567);
or U2848 (N_2848,N_1073,N_1522);
and U2849 (N_2849,N_1519,N_1494);
or U2850 (N_2850,N_1074,N_1559);
nor U2851 (N_2851,N_1807,N_1006);
or U2852 (N_2852,N_1291,N_1203);
nand U2853 (N_2853,N_1387,N_1398);
or U2854 (N_2854,N_1261,N_1195);
and U2855 (N_2855,N_1603,N_1248);
or U2856 (N_2856,N_1094,N_1430);
and U2857 (N_2857,N_1481,N_1900);
xnor U2858 (N_2858,N_1019,N_1319);
or U2859 (N_2859,N_1069,N_1189);
or U2860 (N_2860,N_1477,N_1386);
nand U2861 (N_2861,N_1652,N_1788);
nor U2862 (N_2862,N_1652,N_1920);
nor U2863 (N_2863,N_1577,N_1952);
nor U2864 (N_2864,N_1725,N_1474);
or U2865 (N_2865,N_1786,N_1759);
nor U2866 (N_2866,N_1267,N_1272);
nor U2867 (N_2867,N_1091,N_1217);
or U2868 (N_2868,N_1117,N_1472);
nand U2869 (N_2869,N_1380,N_1027);
nor U2870 (N_2870,N_1594,N_1506);
or U2871 (N_2871,N_1169,N_1591);
nand U2872 (N_2872,N_1903,N_1262);
nand U2873 (N_2873,N_1171,N_1432);
or U2874 (N_2874,N_1747,N_1194);
nand U2875 (N_2875,N_1244,N_1191);
nand U2876 (N_2876,N_1078,N_1534);
nor U2877 (N_2877,N_1381,N_1764);
nand U2878 (N_2878,N_1908,N_1160);
and U2879 (N_2879,N_1452,N_1960);
or U2880 (N_2880,N_1388,N_1306);
nand U2881 (N_2881,N_1382,N_1360);
nor U2882 (N_2882,N_1964,N_1228);
nand U2883 (N_2883,N_1857,N_1663);
or U2884 (N_2884,N_1785,N_1406);
nor U2885 (N_2885,N_1249,N_1706);
or U2886 (N_2886,N_1387,N_1976);
or U2887 (N_2887,N_1814,N_1168);
nand U2888 (N_2888,N_1636,N_1571);
nor U2889 (N_2889,N_1226,N_1428);
nor U2890 (N_2890,N_1673,N_1966);
or U2891 (N_2891,N_1186,N_1811);
nor U2892 (N_2892,N_1098,N_1389);
and U2893 (N_2893,N_1565,N_1131);
nor U2894 (N_2894,N_1105,N_1168);
and U2895 (N_2895,N_1257,N_1761);
nand U2896 (N_2896,N_1000,N_1844);
or U2897 (N_2897,N_1583,N_1351);
or U2898 (N_2898,N_1254,N_1872);
or U2899 (N_2899,N_1734,N_1152);
or U2900 (N_2900,N_1530,N_1363);
nor U2901 (N_2901,N_1972,N_1354);
nor U2902 (N_2902,N_1607,N_1300);
or U2903 (N_2903,N_1050,N_1105);
nand U2904 (N_2904,N_1634,N_1635);
nand U2905 (N_2905,N_1526,N_1152);
and U2906 (N_2906,N_1758,N_1188);
nor U2907 (N_2907,N_1130,N_1561);
or U2908 (N_2908,N_1500,N_1288);
nor U2909 (N_2909,N_1699,N_1458);
or U2910 (N_2910,N_1420,N_1027);
nor U2911 (N_2911,N_1173,N_1887);
and U2912 (N_2912,N_1441,N_1327);
and U2913 (N_2913,N_1858,N_1669);
nor U2914 (N_2914,N_1079,N_1711);
and U2915 (N_2915,N_1652,N_1080);
and U2916 (N_2916,N_1970,N_1669);
nand U2917 (N_2917,N_1899,N_1324);
nor U2918 (N_2918,N_1672,N_1862);
nand U2919 (N_2919,N_1573,N_1044);
or U2920 (N_2920,N_1122,N_1762);
or U2921 (N_2921,N_1772,N_1456);
nand U2922 (N_2922,N_1392,N_1149);
nor U2923 (N_2923,N_1289,N_1861);
nand U2924 (N_2924,N_1858,N_1727);
or U2925 (N_2925,N_1303,N_1276);
and U2926 (N_2926,N_1343,N_1171);
or U2927 (N_2927,N_1481,N_1390);
nand U2928 (N_2928,N_1210,N_1627);
and U2929 (N_2929,N_1210,N_1906);
and U2930 (N_2930,N_1231,N_1172);
nor U2931 (N_2931,N_1437,N_1158);
or U2932 (N_2932,N_1095,N_1944);
nor U2933 (N_2933,N_1811,N_1857);
nand U2934 (N_2934,N_1585,N_1056);
and U2935 (N_2935,N_1654,N_1235);
nand U2936 (N_2936,N_1251,N_1569);
nor U2937 (N_2937,N_1530,N_1525);
or U2938 (N_2938,N_1227,N_1758);
and U2939 (N_2939,N_1469,N_1555);
nand U2940 (N_2940,N_1665,N_1703);
nor U2941 (N_2941,N_1380,N_1715);
and U2942 (N_2942,N_1200,N_1531);
nor U2943 (N_2943,N_1455,N_1206);
or U2944 (N_2944,N_1925,N_1889);
nor U2945 (N_2945,N_1485,N_1020);
or U2946 (N_2946,N_1099,N_1373);
and U2947 (N_2947,N_1385,N_1611);
and U2948 (N_2948,N_1862,N_1471);
or U2949 (N_2949,N_1115,N_1194);
or U2950 (N_2950,N_1791,N_1100);
nand U2951 (N_2951,N_1625,N_1003);
nor U2952 (N_2952,N_1713,N_1379);
nand U2953 (N_2953,N_1281,N_1554);
and U2954 (N_2954,N_1182,N_1786);
and U2955 (N_2955,N_1381,N_1213);
nor U2956 (N_2956,N_1431,N_1632);
nand U2957 (N_2957,N_1390,N_1884);
nand U2958 (N_2958,N_1475,N_1136);
and U2959 (N_2959,N_1461,N_1953);
nand U2960 (N_2960,N_1671,N_1394);
or U2961 (N_2961,N_1096,N_1960);
and U2962 (N_2962,N_1060,N_1747);
nand U2963 (N_2963,N_1786,N_1375);
nand U2964 (N_2964,N_1450,N_1387);
and U2965 (N_2965,N_1635,N_1879);
and U2966 (N_2966,N_1004,N_1402);
nand U2967 (N_2967,N_1358,N_1432);
or U2968 (N_2968,N_1509,N_1958);
nand U2969 (N_2969,N_1464,N_1877);
nor U2970 (N_2970,N_1705,N_1756);
nand U2971 (N_2971,N_1959,N_1891);
nor U2972 (N_2972,N_1062,N_1134);
nor U2973 (N_2973,N_1756,N_1665);
nor U2974 (N_2974,N_1953,N_1892);
nand U2975 (N_2975,N_1774,N_1268);
and U2976 (N_2976,N_1895,N_1050);
or U2977 (N_2977,N_1792,N_1819);
nor U2978 (N_2978,N_1595,N_1855);
and U2979 (N_2979,N_1505,N_1392);
and U2980 (N_2980,N_1274,N_1956);
nor U2981 (N_2981,N_1296,N_1628);
or U2982 (N_2982,N_1745,N_1882);
and U2983 (N_2983,N_1772,N_1463);
and U2984 (N_2984,N_1510,N_1143);
or U2985 (N_2985,N_1755,N_1109);
and U2986 (N_2986,N_1061,N_1256);
nor U2987 (N_2987,N_1345,N_1567);
and U2988 (N_2988,N_1667,N_1453);
nor U2989 (N_2989,N_1078,N_1797);
and U2990 (N_2990,N_1481,N_1422);
nand U2991 (N_2991,N_1624,N_1217);
nor U2992 (N_2992,N_1023,N_1310);
nand U2993 (N_2993,N_1663,N_1087);
nor U2994 (N_2994,N_1080,N_1069);
or U2995 (N_2995,N_1849,N_1827);
and U2996 (N_2996,N_1673,N_1148);
and U2997 (N_2997,N_1033,N_1340);
and U2998 (N_2998,N_1858,N_1905);
or U2999 (N_2999,N_1964,N_1968);
or U3000 (N_3000,N_2820,N_2491);
or U3001 (N_3001,N_2988,N_2031);
nand U3002 (N_3002,N_2384,N_2624);
nor U3003 (N_3003,N_2387,N_2652);
and U3004 (N_3004,N_2185,N_2457);
and U3005 (N_3005,N_2621,N_2873);
nand U3006 (N_3006,N_2656,N_2774);
nand U3007 (N_3007,N_2461,N_2413);
and U3008 (N_3008,N_2120,N_2095);
and U3009 (N_3009,N_2287,N_2973);
or U3010 (N_3010,N_2051,N_2240);
nor U3011 (N_3011,N_2816,N_2422);
or U3012 (N_3012,N_2212,N_2133);
or U3013 (N_3013,N_2136,N_2008);
and U3014 (N_3014,N_2714,N_2448);
and U3015 (N_3015,N_2719,N_2628);
nor U3016 (N_3016,N_2586,N_2552);
and U3017 (N_3017,N_2900,N_2896);
or U3018 (N_3018,N_2489,N_2919);
or U3019 (N_3019,N_2573,N_2319);
or U3020 (N_3020,N_2084,N_2821);
and U3021 (N_3021,N_2112,N_2864);
or U3022 (N_3022,N_2933,N_2672);
nor U3023 (N_3023,N_2655,N_2829);
and U3024 (N_3024,N_2455,N_2712);
or U3025 (N_3025,N_2951,N_2600);
or U3026 (N_3026,N_2889,N_2412);
and U3027 (N_3027,N_2685,N_2307);
or U3028 (N_3028,N_2151,N_2760);
nand U3029 (N_3029,N_2863,N_2576);
or U3030 (N_3030,N_2474,N_2568);
or U3031 (N_3031,N_2466,N_2983);
nor U3032 (N_3032,N_2056,N_2311);
nand U3033 (N_3033,N_2179,N_2267);
or U3034 (N_3034,N_2742,N_2824);
nand U3035 (N_3035,N_2323,N_2665);
and U3036 (N_3036,N_2555,N_2178);
and U3037 (N_3037,N_2511,N_2172);
nand U3038 (N_3038,N_2407,N_2059);
and U3039 (N_3039,N_2823,N_2246);
or U3040 (N_3040,N_2956,N_2321);
or U3041 (N_3041,N_2334,N_2295);
or U3042 (N_3042,N_2107,N_2764);
or U3043 (N_3043,N_2427,N_2129);
nand U3044 (N_3044,N_2072,N_2625);
nor U3045 (N_3045,N_2339,N_2755);
nor U3046 (N_3046,N_2683,N_2618);
nor U3047 (N_3047,N_2473,N_2849);
and U3048 (N_3048,N_2190,N_2698);
or U3049 (N_3049,N_2214,N_2277);
or U3050 (N_3050,N_2741,N_2164);
and U3051 (N_3051,N_2459,N_2364);
and U3052 (N_3052,N_2541,N_2047);
and U3053 (N_3053,N_2077,N_2961);
or U3054 (N_3054,N_2508,N_2682);
nand U3055 (N_3055,N_2987,N_2464);
and U3056 (N_3056,N_2022,N_2910);
or U3057 (N_3057,N_2397,N_2761);
or U3058 (N_3058,N_2981,N_2963);
nand U3059 (N_3059,N_2377,N_2720);
or U3060 (N_3060,N_2001,N_2302);
nor U3061 (N_3061,N_2724,N_2435);
nand U3062 (N_3062,N_2637,N_2867);
and U3063 (N_3063,N_2644,N_2219);
nand U3064 (N_3064,N_2525,N_2937);
nor U3065 (N_3065,N_2594,N_2275);
nand U3066 (N_3066,N_2395,N_2882);
and U3067 (N_3067,N_2374,N_2404);
nand U3068 (N_3068,N_2335,N_2602);
nor U3069 (N_3069,N_2232,N_2163);
and U3070 (N_3070,N_2106,N_2220);
nand U3071 (N_3071,N_2345,N_2233);
nor U3072 (N_3072,N_2601,N_2936);
nand U3073 (N_3073,N_2043,N_2091);
nand U3074 (N_3074,N_2554,N_2924);
nor U3075 (N_3075,N_2386,N_2265);
or U3076 (N_3076,N_2101,N_2639);
nand U3077 (N_3077,N_2748,N_2708);
nand U3078 (N_3078,N_2128,N_2082);
nand U3079 (N_3079,N_2763,N_2293);
or U3080 (N_3080,N_2213,N_2745);
or U3081 (N_3081,N_2901,N_2279);
nor U3082 (N_3082,N_2790,N_2482);
nand U3083 (N_3083,N_2689,N_2123);
nand U3084 (N_3084,N_2296,N_2607);
and U3085 (N_3085,N_2691,N_2857);
nand U3086 (N_3086,N_2899,N_2142);
and U3087 (N_3087,N_2498,N_2423);
and U3088 (N_3088,N_2958,N_2366);
and U3089 (N_3089,N_2271,N_2440);
or U3090 (N_3090,N_2417,N_2888);
nand U3091 (N_3091,N_2690,N_2484);
nand U3092 (N_3092,N_2941,N_2197);
and U3093 (N_3093,N_2065,N_2913);
nor U3094 (N_3094,N_2674,N_2911);
nand U3095 (N_3095,N_2575,N_2029);
or U3096 (N_3096,N_2881,N_2141);
nor U3097 (N_3097,N_2817,N_2336);
nand U3098 (N_3098,N_2634,N_2673);
nand U3099 (N_3099,N_2752,N_2312);
nor U3100 (N_3100,N_2675,N_2874);
and U3101 (N_3101,N_2587,N_2426);
or U3102 (N_3102,N_2801,N_2795);
nor U3103 (N_3103,N_2458,N_2915);
or U3104 (N_3104,N_2053,N_2415);
or U3105 (N_3105,N_2947,N_2659);
nor U3106 (N_3106,N_2174,N_2728);
or U3107 (N_3107,N_2772,N_2878);
or U3108 (N_3108,N_2476,N_2747);
or U3109 (N_3109,N_2081,N_2750);
and U3110 (N_3110,N_2799,N_2950);
nor U3111 (N_3111,N_2773,N_2049);
nor U3112 (N_3112,N_2884,N_2203);
or U3113 (N_3113,N_2754,N_2006);
or U3114 (N_3114,N_2372,N_2202);
nor U3115 (N_3115,N_2405,N_2356);
nor U3116 (N_3116,N_2429,N_2074);
nor U3117 (N_3117,N_2026,N_2617);
and U3118 (N_3118,N_2650,N_2327);
nor U3119 (N_3119,N_2291,N_2481);
and U3120 (N_3120,N_2431,N_2256);
and U3121 (N_3121,N_2975,N_2488);
nand U3122 (N_3122,N_2547,N_2033);
or U3123 (N_3123,N_2478,N_2124);
nor U3124 (N_3124,N_2117,N_2589);
nand U3125 (N_3125,N_2697,N_2999);
and U3126 (N_3126,N_2768,N_2869);
or U3127 (N_3127,N_2737,N_2616);
or U3128 (N_3128,N_2463,N_2414);
and U3129 (N_3129,N_2753,N_2865);
nor U3130 (N_3130,N_2264,N_2068);
and U3131 (N_3131,N_2964,N_2749);
or U3132 (N_3132,N_2251,N_2798);
or U3133 (N_3133,N_2822,N_2276);
or U3134 (N_3134,N_2574,N_2926);
nand U3135 (N_3135,N_2449,N_2286);
nor U3136 (N_3136,N_2371,N_2177);
and U3137 (N_3137,N_2550,N_2347);
nand U3138 (N_3138,N_2153,N_2005);
nor U3139 (N_3139,N_2322,N_2505);
and U3140 (N_3140,N_2211,N_2711);
and U3141 (N_3141,N_2389,N_2702);
or U3142 (N_3142,N_2931,N_2363);
nor U3143 (N_3143,N_2717,N_2416);
nor U3144 (N_3144,N_2565,N_2272);
nor U3145 (N_3145,N_2832,N_2806);
and U3146 (N_3146,N_2859,N_2846);
or U3147 (N_3147,N_2089,N_2492);
and U3148 (N_3148,N_2024,N_2333);
nor U3149 (N_3149,N_2419,N_2470);
nand U3150 (N_3150,N_2401,N_2793);
or U3151 (N_3151,N_2099,N_2441);
and U3152 (N_3152,N_2180,N_2487);
and U3153 (N_3153,N_2181,N_2553);
and U3154 (N_3154,N_2980,N_2205);
and U3155 (N_3155,N_2224,N_2664);
and U3156 (N_3156,N_2432,N_2680);
and U3157 (N_3157,N_2952,N_2306);
nand U3158 (N_3158,N_2111,N_2192);
and U3159 (N_3159,N_2252,N_2135);
or U3160 (N_3160,N_2653,N_2154);
or U3161 (N_3161,N_2860,N_2222);
or U3162 (N_3162,N_2035,N_2445);
nand U3163 (N_3163,N_2209,N_2703);
or U3164 (N_3164,N_2167,N_2827);
and U3165 (N_3165,N_2434,N_2318);
and U3166 (N_3166,N_2144,N_2007);
nor U3167 (N_3167,N_2626,N_2666);
and U3168 (N_3168,N_2572,N_2578);
or U3169 (N_3169,N_2018,N_2842);
nor U3170 (N_3170,N_2393,N_2088);
and U3171 (N_3171,N_2805,N_2803);
and U3172 (N_3172,N_2942,N_2254);
nand U3173 (N_3173,N_2235,N_2844);
and U3174 (N_3174,N_2733,N_2861);
and U3175 (N_3175,N_2346,N_2613);
and U3176 (N_3176,N_2226,N_2403);
or U3177 (N_3177,N_2160,N_2841);
and U3178 (N_3178,N_2765,N_2198);
nor U3179 (N_3179,N_2273,N_2769);
nor U3180 (N_3180,N_2796,N_2695);
nand U3181 (N_3181,N_2905,N_2012);
nand U3182 (N_3182,N_2974,N_2520);
or U3183 (N_3183,N_2157,N_2965);
or U3184 (N_3184,N_2678,N_2704);
or U3185 (N_3185,N_2169,N_2352);
or U3186 (N_3186,N_2684,N_2620);
nor U3187 (N_3187,N_2766,N_2807);
nor U3188 (N_3188,N_2984,N_2040);
and U3189 (N_3189,N_2996,N_2903);
or U3190 (N_3190,N_2969,N_2204);
nor U3191 (N_3191,N_2571,N_2989);
nor U3192 (N_3192,N_2850,N_2917);
and U3193 (N_3193,N_2130,N_2662);
and U3194 (N_3194,N_2923,N_2789);
nor U3195 (N_3195,N_2243,N_2227);
or U3196 (N_3196,N_2585,N_2623);
and U3197 (N_3197,N_2818,N_2320);
and U3198 (N_3198,N_2109,N_2087);
and U3199 (N_3199,N_2075,N_2062);
or U3200 (N_3200,N_2677,N_2839);
or U3201 (N_3201,N_2730,N_2119);
or U3202 (N_3202,N_2028,N_2097);
nand U3203 (N_3203,N_2593,N_2731);
and U3204 (N_3204,N_2070,N_2184);
and U3205 (N_3205,N_2930,N_2149);
and U3206 (N_3206,N_2260,N_2938);
and U3207 (N_3207,N_2443,N_2004);
nor U3208 (N_3208,N_2994,N_2330);
nand U3209 (N_3209,N_2173,N_2979);
xnor U3210 (N_3210,N_2725,N_2343);
nand U3211 (N_3211,N_2556,N_2436);
nand U3212 (N_3212,N_2701,N_2332);
and U3213 (N_3213,N_2721,N_2244);
nor U3214 (N_3214,N_2094,N_2036);
xor U3215 (N_3215,N_2494,N_2944);
nor U3216 (N_3216,N_2837,N_2073);
or U3217 (N_3217,N_2902,N_2301);
or U3218 (N_3218,N_2229,N_2052);
nor U3219 (N_3219,N_2064,N_2085);
nor U3220 (N_3220,N_2840,N_2230);
nor U3221 (N_3221,N_2398,N_2543);
nor U3222 (N_3222,N_2875,N_2558);
and U3223 (N_3223,N_2048,N_2943);
or U3224 (N_3224,N_2269,N_2446);
nor U3225 (N_3225,N_2636,N_2400);
nand U3226 (N_3226,N_2394,N_2115);
nand U3227 (N_3227,N_2581,N_2206);
or U3228 (N_3228,N_2014,N_2583);
and U3229 (N_3229,N_2971,N_2658);
nand U3230 (N_3230,N_2324,N_2615);
and U3231 (N_3231,N_2557,N_2612);
nor U3232 (N_3232,N_2281,N_2605);
and U3233 (N_3233,N_2299,N_2447);
nor U3234 (N_3234,N_2898,N_2609);
or U3235 (N_3235,N_2978,N_2396);
nor U3236 (N_3236,N_2316,N_2582);
or U3237 (N_3237,N_2158,N_2872);
or U3238 (N_3238,N_2736,N_2468);
or U3239 (N_3239,N_2288,N_2542);
or U3240 (N_3240,N_2392,N_2490);
or U3241 (N_3241,N_2707,N_2800);
or U3242 (N_3242,N_2249,N_2137);
and U3243 (N_3243,N_2757,N_2810);
or U3244 (N_3244,N_2236,N_2966);
or U3245 (N_3245,N_2635,N_2519);
nor U3246 (N_3246,N_2044,N_2102);
nor U3247 (N_3247,N_2080,N_2732);
nor U3248 (N_3248,N_2694,N_2580);
nand U3249 (N_3249,N_2166,N_2200);
nor U3250 (N_3250,N_2485,N_2537);
nor U3251 (N_3251,N_2409,N_2071);
nor U3252 (N_3252,N_2630,N_2223);
or U3253 (N_3253,N_2709,N_2096);
nand U3254 (N_3254,N_2970,N_2960);
or U3255 (N_3255,N_2310,N_2746);
nor U3256 (N_3256,N_2852,N_2165);
nor U3257 (N_3257,N_2686,N_2783);
nand U3258 (N_3258,N_2156,N_2460);
nor U3259 (N_3259,N_2237,N_2125);
and U3260 (N_3260,N_2885,N_2228);
and U3261 (N_3261,N_2002,N_2399);
nor U3262 (N_3262,N_2632,N_2502);
and U3263 (N_3263,N_2912,N_2496);
nand U3264 (N_3264,N_2013,N_2274);
and U3265 (N_3265,N_2886,N_2338);
nor U3266 (N_3266,N_2360,N_2104);
nor U3267 (N_3267,N_2247,N_2268);
nor U3268 (N_3268,N_2738,N_2023);
nor U3269 (N_3269,N_2168,N_2908);
or U3270 (N_3270,N_2292,N_2939);
and U3271 (N_3271,N_2162,N_2055);
nand U3272 (N_3272,N_2530,N_2993);
nand U3273 (N_3273,N_2215,N_2139);
nor U3274 (N_3274,N_2495,N_2559);
or U3275 (N_3275,N_2986,N_2241);
nand U3276 (N_3276,N_2500,N_2300);
nand U3277 (N_3277,N_2182,N_2187);
and U3278 (N_3278,N_2877,N_2497);
and U3279 (N_3279,N_2925,N_2922);
and U3280 (N_3280,N_2619,N_2146);
nand U3281 (N_3281,N_2067,N_2242);
nand U3282 (N_3282,N_2041,N_2315);
or U3283 (N_3283,N_2313,N_2880);
and U3284 (N_3284,N_2606,N_2171);
nand U3285 (N_3285,N_2348,N_2210);
nor U3286 (N_3286,N_2000,N_2114);
or U3287 (N_3287,N_2548,N_2949);
nand U3288 (N_3288,N_2700,N_2991);
or U3289 (N_3289,N_2439,N_2083);
nor U3290 (N_3290,N_2289,N_2437);
or U3291 (N_3291,N_2118,N_2365);
or U3292 (N_3292,N_2479,N_2098);
nand U3293 (N_3293,N_2934,N_2921);
nand U3294 (N_3294,N_2518,N_2452);
and U3295 (N_3295,N_2514,N_2444);
or U3296 (N_3296,N_2003,N_2569);
nor U3297 (N_3297,N_2670,N_2828);
nand U3298 (N_3298,N_2050,N_2929);
and U3299 (N_3299,N_2326,N_2294);
and U3300 (N_3300,N_2853,N_2866);
nand U3301 (N_3301,N_2968,N_2016);
nor U3302 (N_3302,N_2560,N_2862);
or U3303 (N_3303,N_2263,N_2019);
nand U3304 (N_3304,N_2779,N_2245);
or U3305 (N_3305,N_2510,N_2017);
and U3306 (N_3306,N_2608,N_2977);
nand U3307 (N_3307,N_2020,N_2876);
and U3308 (N_3308,N_2826,N_2353);
nand U3309 (N_3309,N_2651,N_2015);
nor U3310 (N_3310,N_2871,N_2471);
and U3311 (N_3311,N_2935,N_2643);
or U3312 (N_3312,N_2596,N_2143);
nor U3313 (N_3313,N_2524,N_2967);
nor U3314 (N_3314,N_2676,N_2152);
nand U3315 (N_3315,N_2113,N_2512);
or U3316 (N_3316,N_2797,N_2893);
and U3317 (N_3317,N_2567,N_2390);
and U3318 (N_3318,N_2134,N_2808);
nand U3319 (N_3319,N_2894,N_2868);
or U3320 (N_3320,N_2904,N_2188);
nor U3321 (N_3321,N_2148,N_2475);
nor U3322 (N_3322,N_2945,N_2713);
xor U3323 (N_3323,N_2592,N_2388);
nor U3324 (N_3324,N_2570,N_2551);
nor U3325 (N_3325,N_2599,N_2283);
nand U3326 (N_3326,N_2349,N_2380);
and U3327 (N_3327,N_2025,N_2428);
nand U3328 (N_3328,N_2325,N_2928);
nor U3329 (N_3329,N_2221,N_2718);
nand U3330 (N_3330,N_2743,N_2406);
or U3331 (N_3331,N_2261,N_2838);
and U3332 (N_3332,N_2830,N_2058);
nand U3333 (N_3333,N_2453,N_2054);
nor U3334 (N_3334,N_2776,N_2465);
and U3335 (N_3335,N_2217,N_2649);
nor U3336 (N_3336,N_2813,N_2507);
nor U3337 (N_3337,N_2706,N_2739);
nand U3338 (N_3338,N_2442,N_2234);
nor U3339 (N_3339,N_2533,N_2410);
nor U3340 (N_3340,N_2314,N_2782);
nor U3341 (N_3341,N_2155,N_2648);
nor U3342 (N_3342,N_2544,N_2784);
nand U3343 (N_3343,N_2430,N_2564);
nand U3344 (N_3344,N_2159,N_2170);
nor U3345 (N_3345,N_2402,N_2424);
and U3346 (N_3346,N_2127,N_2671);
nor U3347 (N_3347,N_2255,N_2657);
or U3348 (N_3348,N_2948,N_2186);
nor U3349 (N_3349,N_2833,N_2549);
nor U3350 (N_3350,N_2278,N_2914);
and U3351 (N_3351,N_2357,N_2751);
and U3352 (N_3352,N_2340,N_2940);
nand U3353 (N_3353,N_2408,N_2317);
nand U3354 (N_3354,N_2831,N_2802);
nor U3355 (N_3355,N_2727,N_2845);
and U3356 (N_3356,N_2982,N_2610);
nor U3357 (N_3357,N_2561,N_2734);
or U3358 (N_3358,N_2391,N_2962);
nand U3359 (N_3359,N_2577,N_2425);
nor U3360 (N_3360,N_2614,N_2641);
and U3361 (N_3361,N_2629,N_2039);
nand U3362 (N_3362,N_2038,N_2250);
and U3363 (N_3363,N_2715,N_2257);
nor U3364 (N_3364,N_2562,N_2042);
nor U3365 (N_3365,N_2383,N_2858);
and U3366 (N_3366,N_2526,N_2010);
and U3367 (N_3367,N_2138,N_2814);
nor U3368 (N_3368,N_2598,N_2385);
nor U3369 (N_3369,N_2262,N_2909);
nand U3370 (N_3370,N_2927,N_2661);
nand U3371 (N_3371,N_2916,N_2955);
nor U3372 (N_3372,N_2093,N_2090);
and U3373 (N_3373,N_2595,N_2775);
and U3374 (N_3374,N_2998,N_2045);
nor U3375 (N_3375,N_2270,N_2483);
or U3376 (N_3376,N_2906,N_2532);
nor U3377 (N_3377,N_2531,N_2344);
nor U3378 (N_3378,N_2195,N_2699);
or U3379 (N_3379,N_2705,N_2856);
nand U3380 (N_3380,N_2959,N_2027);
and U3381 (N_3381,N_2778,N_2780);
nor U3382 (N_3382,N_2835,N_2078);
nor U3383 (N_3383,N_2812,N_2588);
and U3384 (N_3384,N_2451,N_2358);
or U3385 (N_3385,N_2579,N_2216);
or U3386 (N_3386,N_2540,N_2342);
nor U3387 (N_3387,N_2298,N_2034);
nor U3388 (N_3388,N_2480,N_2063);
nor U3389 (N_3389,N_2669,N_2645);
nand U3390 (N_3390,N_2450,N_2030);
and U3391 (N_3391,N_2920,N_2469);
or U3392 (N_3392,N_2193,N_2337);
nand U3393 (N_3393,N_2499,N_2297);
and U3394 (N_3394,N_2726,N_2369);
and U3395 (N_3395,N_2515,N_2069);
and U3396 (N_3396,N_2781,N_2883);
nor U3397 (N_3397,N_2517,N_2819);
or U3398 (N_3398,N_2815,N_2176);
nor U3399 (N_3399,N_2597,N_2723);
nor U3400 (N_3400,N_2590,N_2066);
nor U3401 (N_3401,N_2284,N_2667);
and U3402 (N_3402,N_2785,N_2341);
or U3403 (N_3403,N_2199,N_2021);
nand U3404 (N_3404,N_2032,N_2546);
nor U3405 (N_3405,N_2116,N_2767);
and U3406 (N_3406,N_2642,N_2836);
and U3407 (N_3407,N_2660,N_2654);
nand U3408 (N_3408,N_2362,N_2759);
nor U3409 (N_3409,N_2486,N_2504);
or U3410 (N_3410,N_2638,N_2462);
nand U3411 (N_3411,N_2848,N_2175);
nor U3412 (N_3412,N_2100,N_2382);
xor U3413 (N_3413,N_2282,N_2538);
nor U3414 (N_3414,N_2954,N_2354);
nor U3415 (N_3415,N_2990,N_2527);
nand U3416 (N_3416,N_2140,N_2918);
or U3417 (N_3417,N_2132,N_2604);
and U3418 (N_3418,N_2368,N_2011);
nand U3419 (N_3419,N_2953,N_2477);
nand U3420 (N_3420,N_2603,N_2329);
or U3421 (N_3421,N_2710,N_2304);
and U3422 (N_3422,N_2421,N_2679);
nand U3423 (N_3423,N_2501,N_2566);
and U3424 (N_3424,N_2009,N_2328);
nand U3425 (N_3425,N_2646,N_2418);
or U3426 (N_3426,N_2108,N_2591);
and U3427 (N_3427,N_2456,N_2529);
or U3428 (N_3428,N_2521,N_2259);
nand U3429 (N_3429,N_2290,N_2892);
nand U3430 (N_3430,N_2756,N_2253);
or U3431 (N_3431,N_2771,N_2231);
nor U3432 (N_3432,N_2985,N_2536);
nor U3433 (N_3433,N_2218,N_2631);
nand U3434 (N_3434,N_2788,N_2787);
and U3435 (N_3435,N_2891,N_2611);
nor U3436 (N_3436,N_2309,N_2351);
and U3437 (N_3437,N_2183,N_2897);
nor U3438 (N_3438,N_2758,N_2992);
nor U3439 (N_3439,N_2622,N_2509);
or U3440 (N_3440,N_2331,N_2668);
and U3441 (N_3441,N_2248,N_2522);
nand U3442 (N_3442,N_2126,N_2729);
nor U3443 (N_3443,N_2528,N_2834);
or U3444 (N_3444,N_2870,N_2189);
and U3445 (N_3445,N_2381,N_2121);
and U3446 (N_3446,N_2266,N_2825);
or U3447 (N_3447,N_2305,N_2308);
nand U3448 (N_3448,N_2640,N_2957);
or U3449 (N_3449,N_2145,N_2285);
and U3450 (N_3450,N_2046,N_2225);
and U3451 (N_3451,N_2370,N_2535);
or U3452 (N_3452,N_2086,N_2791);
and U3453 (N_3453,N_2191,N_2681);
or U3454 (N_3454,N_2687,N_2196);
or U3455 (N_3455,N_2379,N_2037);
and U3456 (N_3456,N_2207,N_2740);
and U3457 (N_3457,N_2851,N_2563);
nor U3458 (N_3458,N_2584,N_2361);
or U3459 (N_3459,N_2688,N_2843);
and U3460 (N_3460,N_2373,N_2735);
and U3461 (N_3461,N_2057,N_2907);
nand U3462 (N_3462,N_2545,N_2411);
and U3463 (N_3463,N_2633,N_2895);
and U3464 (N_3464,N_2493,N_2534);
or U3465 (N_3465,N_2367,N_2854);
and U3466 (N_3466,N_2770,N_2280);
or U3467 (N_3467,N_2744,N_2811);
and U3468 (N_3468,N_2539,N_2433);
nor U3469 (N_3469,N_2809,N_2376);
nand U3470 (N_3470,N_2438,N_2467);
nor U3471 (N_3471,N_2777,N_2794);
and U3472 (N_3472,N_2454,N_2103);
or U3473 (N_3473,N_2105,N_2350);
nor U3474 (N_3474,N_2762,N_2359);
and U3475 (N_3475,N_2355,N_2122);
and U3476 (N_3476,N_2506,N_2513);
and U3477 (N_3477,N_2995,N_2150);
or U3478 (N_3478,N_2239,N_2147);
and U3479 (N_3479,N_2378,N_2092);
and U3480 (N_3480,N_2786,N_2847);
and U3481 (N_3481,N_2110,N_2627);
or U3482 (N_3482,N_2855,N_2804);
nand U3483 (N_3483,N_2722,N_2879);
nor U3484 (N_3484,N_2201,N_2420);
and U3485 (N_3485,N_2693,N_2887);
nor U3486 (N_3486,N_2131,N_2076);
nor U3487 (N_3487,N_2946,N_2997);
and U3488 (N_3488,N_2716,N_2523);
or U3489 (N_3489,N_2696,N_2792);
or U3490 (N_3490,N_2976,N_2516);
nor U3491 (N_3491,N_2208,N_2258);
nor U3492 (N_3492,N_2692,N_2503);
nor U3493 (N_3493,N_2303,N_2375);
nand U3494 (N_3494,N_2238,N_2060);
or U3495 (N_3495,N_2194,N_2079);
or U3496 (N_3496,N_2161,N_2647);
and U3497 (N_3497,N_2932,N_2061);
or U3498 (N_3498,N_2663,N_2890);
or U3499 (N_3499,N_2972,N_2472);
nand U3500 (N_3500,N_2251,N_2857);
and U3501 (N_3501,N_2511,N_2941);
and U3502 (N_3502,N_2444,N_2875);
nor U3503 (N_3503,N_2549,N_2971);
and U3504 (N_3504,N_2800,N_2689);
nand U3505 (N_3505,N_2076,N_2019);
or U3506 (N_3506,N_2880,N_2802);
or U3507 (N_3507,N_2930,N_2179);
nor U3508 (N_3508,N_2850,N_2687);
and U3509 (N_3509,N_2312,N_2444);
or U3510 (N_3510,N_2874,N_2212);
nor U3511 (N_3511,N_2405,N_2909);
and U3512 (N_3512,N_2016,N_2368);
or U3513 (N_3513,N_2131,N_2485);
and U3514 (N_3514,N_2966,N_2412);
nand U3515 (N_3515,N_2638,N_2589);
nand U3516 (N_3516,N_2911,N_2448);
xnor U3517 (N_3517,N_2140,N_2317);
or U3518 (N_3518,N_2694,N_2460);
and U3519 (N_3519,N_2164,N_2722);
and U3520 (N_3520,N_2754,N_2522);
or U3521 (N_3521,N_2103,N_2692);
and U3522 (N_3522,N_2737,N_2571);
nand U3523 (N_3523,N_2303,N_2664);
nor U3524 (N_3524,N_2501,N_2373);
nor U3525 (N_3525,N_2403,N_2641);
and U3526 (N_3526,N_2930,N_2943);
nor U3527 (N_3527,N_2402,N_2380);
or U3528 (N_3528,N_2463,N_2691);
and U3529 (N_3529,N_2055,N_2207);
and U3530 (N_3530,N_2423,N_2369);
nand U3531 (N_3531,N_2098,N_2315);
and U3532 (N_3532,N_2732,N_2532);
nor U3533 (N_3533,N_2135,N_2641);
or U3534 (N_3534,N_2040,N_2710);
and U3535 (N_3535,N_2827,N_2151);
or U3536 (N_3536,N_2180,N_2024);
nand U3537 (N_3537,N_2676,N_2163);
nor U3538 (N_3538,N_2655,N_2982);
and U3539 (N_3539,N_2297,N_2833);
or U3540 (N_3540,N_2411,N_2395);
and U3541 (N_3541,N_2591,N_2819);
or U3542 (N_3542,N_2679,N_2533);
or U3543 (N_3543,N_2494,N_2694);
nor U3544 (N_3544,N_2843,N_2948);
or U3545 (N_3545,N_2446,N_2804);
nand U3546 (N_3546,N_2236,N_2493);
and U3547 (N_3547,N_2522,N_2921);
and U3548 (N_3548,N_2420,N_2411);
and U3549 (N_3549,N_2176,N_2272);
nor U3550 (N_3550,N_2002,N_2278);
or U3551 (N_3551,N_2330,N_2717);
and U3552 (N_3552,N_2760,N_2218);
nor U3553 (N_3553,N_2854,N_2322);
nor U3554 (N_3554,N_2776,N_2955);
xor U3555 (N_3555,N_2011,N_2523);
nor U3556 (N_3556,N_2888,N_2669);
nor U3557 (N_3557,N_2220,N_2385);
nand U3558 (N_3558,N_2300,N_2832);
nand U3559 (N_3559,N_2523,N_2472);
nand U3560 (N_3560,N_2684,N_2592);
xor U3561 (N_3561,N_2588,N_2773);
nand U3562 (N_3562,N_2701,N_2278);
or U3563 (N_3563,N_2831,N_2157);
nor U3564 (N_3564,N_2377,N_2825);
nand U3565 (N_3565,N_2634,N_2798);
or U3566 (N_3566,N_2267,N_2070);
or U3567 (N_3567,N_2781,N_2905);
and U3568 (N_3568,N_2850,N_2356);
and U3569 (N_3569,N_2254,N_2988);
nor U3570 (N_3570,N_2404,N_2147);
nand U3571 (N_3571,N_2417,N_2193);
nand U3572 (N_3572,N_2527,N_2072);
and U3573 (N_3573,N_2103,N_2165);
nor U3574 (N_3574,N_2765,N_2495);
and U3575 (N_3575,N_2897,N_2750);
or U3576 (N_3576,N_2688,N_2933);
or U3577 (N_3577,N_2032,N_2358);
and U3578 (N_3578,N_2483,N_2434);
or U3579 (N_3579,N_2485,N_2455);
nand U3580 (N_3580,N_2036,N_2192);
and U3581 (N_3581,N_2643,N_2067);
and U3582 (N_3582,N_2997,N_2479);
and U3583 (N_3583,N_2045,N_2785);
nor U3584 (N_3584,N_2484,N_2604);
nand U3585 (N_3585,N_2043,N_2584);
or U3586 (N_3586,N_2018,N_2216);
and U3587 (N_3587,N_2168,N_2989);
or U3588 (N_3588,N_2806,N_2328);
nor U3589 (N_3589,N_2615,N_2720);
or U3590 (N_3590,N_2526,N_2878);
nand U3591 (N_3591,N_2053,N_2274);
or U3592 (N_3592,N_2722,N_2967);
or U3593 (N_3593,N_2669,N_2166);
nand U3594 (N_3594,N_2907,N_2467);
nand U3595 (N_3595,N_2065,N_2836);
nand U3596 (N_3596,N_2242,N_2651);
or U3597 (N_3597,N_2669,N_2533);
or U3598 (N_3598,N_2074,N_2908);
nand U3599 (N_3599,N_2847,N_2303);
nand U3600 (N_3600,N_2242,N_2653);
nand U3601 (N_3601,N_2620,N_2275);
nand U3602 (N_3602,N_2267,N_2523);
nand U3603 (N_3603,N_2958,N_2023);
nand U3604 (N_3604,N_2900,N_2304);
nor U3605 (N_3605,N_2806,N_2895);
nor U3606 (N_3606,N_2745,N_2785);
nor U3607 (N_3607,N_2995,N_2341);
nand U3608 (N_3608,N_2513,N_2913);
and U3609 (N_3609,N_2733,N_2490);
or U3610 (N_3610,N_2253,N_2598);
nor U3611 (N_3611,N_2242,N_2124);
or U3612 (N_3612,N_2053,N_2838);
or U3613 (N_3613,N_2786,N_2115);
or U3614 (N_3614,N_2687,N_2942);
nor U3615 (N_3615,N_2603,N_2319);
nand U3616 (N_3616,N_2428,N_2858);
nand U3617 (N_3617,N_2021,N_2627);
nand U3618 (N_3618,N_2077,N_2923);
or U3619 (N_3619,N_2101,N_2035);
nor U3620 (N_3620,N_2616,N_2252);
nand U3621 (N_3621,N_2470,N_2668);
and U3622 (N_3622,N_2417,N_2146);
nor U3623 (N_3623,N_2303,N_2007);
nor U3624 (N_3624,N_2185,N_2237);
nor U3625 (N_3625,N_2956,N_2349);
and U3626 (N_3626,N_2400,N_2960);
nor U3627 (N_3627,N_2557,N_2632);
or U3628 (N_3628,N_2355,N_2439);
or U3629 (N_3629,N_2434,N_2398);
and U3630 (N_3630,N_2181,N_2395);
or U3631 (N_3631,N_2530,N_2204);
and U3632 (N_3632,N_2239,N_2292);
nor U3633 (N_3633,N_2960,N_2112);
or U3634 (N_3634,N_2834,N_2648);
nor U3635 (N_3635,N_2794,N_2357);
and U3636 (N_3636,N_2284,N_2271);
and U3637 (N_3637,N_2550,N_2742);
nor U3638 (N_3638,N_2050,N_2450);
and U3639 (N_3639,N_2039,N_2042);
and U3640 (N_3640,N_2891,N_2945);
or U3641 (N_3641,N_2872,N_2366);
or U3642 (N_3642,N_2516,N_2346);
nor U3643 (N_3643,N_2842,N_2257);
nand U3644 (N_3644,N_2610,N_2255);
or U3645 (N_3645,N_2498,N_2730);
nor U3646 (N_3646,N_2306,N_2656);
or U3647 (N_3647,N_2456,N_2214);
nor U3648 (N_3648,N_2401,N_2299);
and U3649 (N_3649,N_2464,N_2353);
nand U3650 (N_3650,N_2475,N_2334);
or U3651 (N_3651,N_2865,N_2277);
and U3652 (N_3652,N_2901,N_2419);
nand U3653 (N_3653,N_2562,N_2015);
nor U3654 (N_3654,N_2075,N_2170);
or U3655 (N_3655,N_2729,N_2555);
and U3656 (N_3656,N_2112,N_2906);
nand U3657 (N_3657,N_2216,N_2809);
or U3658 (N_3658,N_2461,N_2535);
or U3659 (N_3659,N_2072,N_2958);
or U3660 (N_3660,N_2550,N_2693);
nor U3661 (N_3661,N_2469,N_2389);
nand U3662 (N_3662,N_2787,N_2014);
and U3663 (N_3663,N_2618,N_2472);
nor U3664 (N_3664,N_2842,N_2262);
nor U3665 (N_3665,N_2331,N_2974);
and U3666 (N_3666,N_2502,N_2798);
and U3667 (N_3667,N_2976,N_2833);
or U3668 (N_3668,N_2748,N_2863);
nor U3669 (N_3669,N_2218,N_2246);
and U3670 (N_3670,N_2282,N_2498);
nand U3671 (N_3671,N_2807,N_2646);
nand U3672 (N_3672,N_2732,N_2987);
nor U3673 (N_3673,N_2159,N_2468);
nor U3674 (N_3674,N_2387,N_2920);
xor U3675 (N_3675,N_2059,N_2094);
or U3676 (N_3676,N_2441,N_2581);
nand U3677 (N_3677,N_2071,N_2446);
nand U3678 (N_3678,N_2651,N_2200);
nor U3679 (N_3679,N_2129,N_2975);
or U3680 (N_3680,N_2986,N_2740);
and U3681 (N_3681,N_2626,N_2248);
nor U3682 (N_3682,N_2563,N_2375);
or U3683 (N_3683,N_2897,N_2140);
nand U3684 (N_3684,N_2134,N_2765);
or U3685 (N_3685,N_2337,N_2096);
nor U3686 (N_3686,N_2687,N_2256);
nand U3687 (N_3687,N_2739,N_2398);
nor U3688 (N_3688,N_2972,N_2511);
or U3689 (N_3689,N_2407,N_2295);
nor U3690 (N_3690,N_2034,N_2233);
and U3691 (N_3691,N_2783,N_2148);
nand U3692 (N_3692,N_2430,N_2253);
nor U3693 (N_3693,N_2534,N_2882);
and U3694 (N_3694,N_2456,N_2801);
nand U3695 (N_3695,N_2202,N_2084);
or U3696 (N_3696,N_2443,N_2985);
or U3697 (N_3697,N_2061,N_2482);
or U3698 (N_3698,N_2176,N_2447);
nor U3699 (N_3699,N_2593,N_2646);
nand U3700 (N_3700,N_2076,N_2238);
or U3701 (N_3701,N_2027,N_2263);
and U3702 (N_3702,N_2989,N_2613);
nand U3703 (N_3703,N_2999,N_2396);
nor U3704 (N_3704,N_2637,N_2840);
nor U3705 (N_3705,N_2114,N_2668);
nand U3706 (N_3706,N_2267,N_2034);
nor U3707 (N_3707,N_2620,N_2778);
or U3708 (N_3708,N_2860,N_2361);
and U3709 (N_3709,N_2244,N_2254);
nand U3710 (N_3710,N_2222,N_2679);
or U3711 (N_3711,N_2621,N_2396);
nor U3712 (N_3712,N_2296,N_2312);
or U3713 (N_3713,N_2124,N_2739);
nand U3714 (N_3714,N_2679,N_2905);
and U3715 (N_3715,N_2885,N_2899);
or U3716 (N_3716,N_2003,N_2968);
or U3717 (N_3717,N_2724,N_2583);
or U3718 (N_3718,N_2696,N_2286);
and U3719 (N_3719,N_2533,N_2734);
or U3720 (N_3720,N_2991,N_2964);
nor U3721 (N_3721,N_2523,N_2377);
and U3722 (N_3722,N_2363,N_2229);
xnor U3723 (N_3723,N_2142,N_2891);
nor U3724 (N_3724,N_2592,N_2210);
nor U3725 (N_3725,N_2916,N_2160);
nor U3726 (N_3726,N_2908,N_2317);
nand U3727 (N_3727,N_2116,N_2727);
nor U3728 (N_3728,N_2077,N_2914);
and U3729 (N_3729,N_2897,N_2295);
nor U3730 (N_3730,N_2901,N_2907);
nand U3731 (N_3731,N_2220,N_2403);
nor U3732 (N_3732,N_2154,N_2664);
and U3733 (N_3733,N_2745,N_2101);
nand U3734 (N_3734,N_2274,N_2309);
nor U3735 (N_3735,N_2043,N_2891);
nand U3736 (N_3736,N_2615,N_2809);
and U3737 (N_3737,N_2925,N_2760);
nand U3738 (N_3738,N_2247,N_2683);
nand U3739 (N_3739,N_2559,N_2130);
nor U3740 (N_3740,N_2566,N_2967);
nor U3741 (N_3741,N_2753,N_2409);
or U3742 (N_3742,N_2297,N_2771);
and U3743 (N_3743,N_2190,N_2540);
nor U3744 (N_3744,N_2032,N_2256);
nor U3745 (N_3745,N_2437,N_2568);
or U3746 (N_3746,N_2234,N_2343);
or U3747 (N_3747,N_2329,N_2250);
and U3748 (N_3748,N_2760,N_2936);
xnor U3749 (N_3749,N_2992,N_2166);
nand U3750 (N_3750,N_2347,N_2599);
nor U3751 (N_3751,N_2265,N_2676);
nor U3752 (N_3752,N_2508,N_2524);
nor U3753 (N_3753,N_2791,N_2264);
nor U3754 (N_3754,N_2350,N_2079);
and U3755 (N_3755,N_2940,N_2503);
nor U3756 (N_3756,N_2419,N_2044);
or U3757 (N_3757,N_2350,N_2145);
or U3758 (N_3758,N_2825,N_2525);
or U3759 (N_3759,N_2779,N_2743);
nand U3760 (N_3760,N_2803,N_2680);
nand U3761 (N_3761,N_2361,N_2078);
or U3762 (N_3762,N_2532,N_2859);
and U3763 (N_3763,N_2175,N_2508);
or U3764 (N_3764,N_2482,N_2128);
nor U3765 (N_3765,N_2766,N_2564);
nand U3766 (N_3766,N_2423,N_2743);
nand U3767 (N_3767,N_2047,N_2957);
or U3768 (N_3768,N_2263,N_2273);
nand U3769 (N_3769,N_2547,N_2402);
nor U3770 (N_3770,N_2385,N_2104);
or U3771 (N_3771,N_2852,N_2772);
nor U3772 (N_3772,N_2694,N_2094);
nand U3773 (N_3773,N_2526,N_2408);
and U3774 (N_3774,N_2836,N_2155);
and U3775 (N_3775,N_2308,N_2141);
or U3776 (N_3776,N_2392,N_2398);
or U3777 (N_3777,N_2652,N_2617);
nand U3778 (N_3778,N_2227,N_2154);
or U3779 (N_3779,N_2797,N_2786);
and U3780 (N_3780,N_2005,N_2064);
nand U3781 (N_3781,N_2348,N_2944);
and U3782 (N_3782,N_2723,N_2208);
and U3783 (N_3783,N_2429,N_2740);
or U3784 (N_3784,N_2487,N_2146);
or U3785 (N_3785,N_2432,N_2627);
nor U3786 (N_3786,N_2925,N_2911);
nand U3787 (N_3787,N_2684,N_2599);
or U3788 (N_3788,N_2592,N_2408);
nand U3789 (N_3789,N_2063,N_2602);
or U3790 (N_3790,N_2658,N_2588);
and U3791 (N_3791,N_2862,N_2053);
and U3792 (N_3792,N_2097,N_2073);
nand U3793 (N_3793,N_2947,N_2906);
and U3794 (N_3794,N_2901,N_2927);
nor U3795 (N_3795,N_2789,N_2177);
xor U3796 (N_3796,N_2672,N_2886);
and U3797 (N_3797,N_2448,N_2864);
nand U3798 (N_3798,N_2770,N_2326);
and U3799 (N_3799,N_2010,N_2293);
and U3800 (N_3800,N_2446,N_2946);
and U3801 (N_3801,N_2133,N_2760);
and U3802 (N_3802,N_2636,N_2786);
nor U3803 (N_3803,N_2627,N_2739);
and U3804 (N_3804,N_2302,N_2454);
or U3805 (N_3805,N_2560,N_2374);
and U3806 (N_3806,N_2228,N_2121);
and U3807 (N_3807,N_2924,N_2328);
or U3808 (N_3808,N_2220,N_2277);
or U3809 (N_3809,N_2599,N_2379);
nor U3810 (N_3810,N_2518,N_2793);
or U3811 (N_3811,N_2871,N_2637);
or U3812 (N_3812,N_2311,N_2219);
nor U3813 (N_3813,N_2284,N_2794);
or U3814 (N_3814,N_2668,N_2389);
nor U3815 (N_3815,N_2686,N_2442);
and U3816 (N_3816,N_2456,N_2627);
and U3817 (N_3817,N_2124,N_2141);
nand U3818 (N_3818,N_2083,N_2485);
or U3819 (N_3819,N_2332,N_2786);
and U3820 (N_3820,N_2519,N_2285);
nor U3821 (N_3821,N_2365,N_2499);
nor U3822 (N_3822,N_2678,N_2399);
and U3823 (N_3823,N_2916,N_2950);
and U3824 (N_3824,N_2136,N_2190);
nand U3825 (N_3825,N_2811,N_2027);
and U3826 (N_3826,N_2184,N_2003);
nand U3827 (N_3827,N_2614,N_2316);
or U3828 (N_3828,N_2627,N_2844);
nand U3829 (N_3829,N_2098,N_2535);
nor U3830 (N_3830,N_2203,N_2495);
and U3831 (N_3831,N_2668,N_2971);
nand U3832 (N_3832,N_2655,N_2462);
or U3833 (N_3833,N_2082,N_2037);
nand U3834 (N_3834,N_2035,N_2344);
or U3835 (N_3835,N_2952,N_2946);
nand U3836 (N_3836,N_2548,N_2179);
nor U3837 (N_3837,N_2685,N_2818);
and U3838 (N_3838,N_2130,N_2911);
nor U3839 (N_3839,N_2863,N_2418);
or U3840 (N_3840,N_2861,N_2056);
nor U3841 (N_3841,N_2448,N_2208);
or U3842 (N_3842,N_2016,N_2030);
nor U3843 (N_3843,N_2404,N_2993);
or U3844 (N_3844,N_2662,N_2528);
nand U3845 (N_3845,N_2012,N_2936);
nor U3846 (N_3846,N_2346,N_2830);
xor U3847 (N_3847,N_2573,N_2324);
and U3848 (N_3848,N_2856,N_2634);
nor U3849 (N_3849,N_2502,N_2586);
nor U3850 (N_3850,N_2268,N_2761);
and U3851 (N_3851,N_2327,N_2486);
nand U3852 (N_3852,N_2867,N_2071);
nor U3853 (N_3853,N_2229,N_2712);
or U3854 (N_3854,N_2017,N_2048);
nand U3855 (N_3855,N_2123,N_2252);
nor U3856 (N_3856,N_2852,N_2091);
nand U3857 (N_3857,N_2612,N_2393);
nand U3858 (N_3858,N_2292,N_2546);
nand U3859 (N_3859,N_2579,N_2076);
or U3860 (N_3860,N_2697,N_2433);
nor U3861 (N_3861,N_2424,N_2961);
nand U3862 (N_3862,N_2364,N_2668);
nor U3863 (N_3863,N_2471,N_2191);
nand U3864 (N_3864,N_2909,N_2329);
nand U3865 (N_3865,N_2404,N_2367);
and U3866 (N_3866,N_2144,N_2460);
nand U3867 (N_3867,N_2860,N_2059);
nand U3868 (N_3868,N_2774,N_2294);
and U3869 (N_3869,N_2472,N_2585);
nor U3870 (N_3870,N_2635,N_2981);
or U3871 (N_3871,N_2403,N_2758);
and U3872 (N_3872,N_2800,N_2940);
or U3873 (N_3873,N_2475,N_2402);
and U3874 (N_3874,N_2042,N_2016);
and U3875 (N_3875,N_2743,N_2574);
or U3876 (N_3876,N_2022,N_2235);
or U3877 (N_3877,N_2144,N_2070);
nor U3878 (N_3878,N_2777,N_2100);
and U3879 (N_3879,N_2487,N_2689);
nand U3880 (N_3880,N_2342,N_2859);
nor U3881 (N_3881,N_2296,N_2945);
and U3882 (N_3882,N_2637,N_2338);
or U3883 (N_3883,N_2898,N_2165);
or U3884 (N_3884,N_2178,N_2742);
nand U3885 (N_3885,N_2854,N_2209);
nand U3886 (N_3886,N_2658,N_2832);
nor U3887 (N_3887,N_2486,N_2520);
and U3888 (N_3888,N_2427,N_2753);
nor U3889 (N_3889,N_2905,N_2587);
or U3890 (N_3890,N_2586,N_2496);
nand U3891 (N_3891,N_2275,N_2639);
nand U3892 (N_3892,N_2011,N_2456);
or U3893 (N_3893,N_2062,N_2795);
nand U3894 (N_3894,N_2162,N_2195);
and U3895 (N_3895,N_2117,N_2321);
and U3896 (N_3896,N_2235,N_2122);
or U3897 (N_3897,N_2392,N_2638);
nor U3898 (N_3898,N_2655,N_2811);
nand U3899 (N_3899,N_2993,N_2465);
nor U3900 (N_3900,N_2218,N_2468);
nor U3901 (N_3901,N_2909,N_2263);
or U3902 (N_3902,N_2490,N_2204);
and U3903 (N_3903,N_2846,N_2935);
and U3904 (N_3904,N_2483,N_2932);
or U3905 (N_3905,N_2196,N_2350);
nor U3906 (N_3906,N_2560,N_2681);
and U3907 (N_3907,N_2343,N_2989);
nand U3908 (N_3908,N_2836,N_2987);
and U3909 (N_3909,N_2068,N_2485);
nor U3910 (N_3910,N_2165,N_2389);
or U3911 (N_3911,N_2597,N_2229);
or U3912 (N_3912,N_2339,N_2841);
or U3913 (N_3913,N_2384,N_2324);
and U3914 (N_3914,N_2831,N_2982);
or U3915 (N_3915,N_2903,N_2851);
or U3916 (N_3916,N_2494,N_2415);
or U3917 (N_3917,N_2930,N_2615);
and U3918 (N_3918,N_2271,N_2657);
nand U3919 (N_3919,N_2787,N_2515);
or U3920 (N_3920,N_2126,N_2355);
xnor U3921 (N_3921,N_2365,N_2273);
nand U3922 (N_3922,N_2446,N_2355);
and U3923 (N_3923,N_2223,N_2250);
or U3924 (N_3924,N_2189,N_2298);
or U3925 (N_3925,N_2148,N_2735);
and U3926 (N_3926,N_2294,N_2793);
nor U3927 (N_3927,N_2409,N_2895);
or U3928 (N_3928,N_2741,N_2043);
or U3929 (N_3929,N_2387,N_2483);
or U3930 (N_3930,N_2844,N_2569);
xor U3931 (N_3931,N_2659,N_2257);
nor U3932 (N_3932,N_2465,N_2340);
or U3933 (N_3933,N_2930,N_2670);
nor U3934 (N_3934,N_2308,N_2549);
nand U3935 (N_3935,N_2886,N_2424);
nand U3936 (N_3936,N_2941,N_2036);
nor U3937 (N_3937,N_2893,N_2570);
or U3938 (N_3938,N_2382,N_2548);
and U3939 (N_3939,N_2917,N_2042);
and U3940 (N_3940,N_2165,N_2126);
or U3941 (N_3941,N_2478,N_2238);
and U3942 (N_3942,N_2507,N_2419);
nand U3943 (N_3943,N_2028,N_2986);
nor U3944 (N_3944,N_2170,N_2572);
and U3945 (N_3945,N_2251,N_2396);
and U3946 (N_3946,N_2505,N_2930);
and U3947 (N_3947,N_2703,N_2728);
or U3948 (N_3948,N_2222,N_2503);
xnor U3949 (N_3949,N_2347,N_2539);
and U3950 (N_3950,N_2604,N_2252);
nor U3951 (N_3951,N_2814,N_2697);
nand U3952 (N_3952,N_2067,N_2976);
nor U3953 (N_3953,N_2536,N_2579);
or U3954 (N_3954,N_2236,N_2163);
nand U3955 (N_3955,N_2413,N_2525);
nor U3956 (N_3956,N_2421,N_2591);
or U3957 (N_3957,N_2516,N_2012);
or U3958 (N_3958,N_2836,N_2196);
nor U3959 (N_3959,N_2626,N_2731);
nand U3960 (N_3960,N_2874,N_2281);
nor U3961 (N_3961,N_2514,N_2958);
nor U3962 (N_3962,N_2450,N_2705);
nor U3963 (N_3963,N_2266,N_2769);
nand U3964 (N_3964,N_2270,N_2216);
or U3965 (N_3965,N_2247,N_2900);
and U3966 (N_3966,N_2203,N_2688);
nor U3967 (N_3967,N_2796,N_2645);
nand U3968 (N_3968,N_2309,N_2654);
nor U3969 (N_3969,N_2360,N_2414);
nor U3970 (N_3970,N_2734,N_2604);
nand U3971 (N_3971,N_2111,N_2600);
nand U3972 (N_3972,N_2447,N_2008);
or U3973 (N_3973,N_2912,N_2622);
or U3974 (N_3974,N_2591,N_2887);
nand U3975 (N_3975,N_2584,N_2496);
nand U3976 (N_3976,N_2866,N_2158);
or U3977 (N_3977,N_2589,N_2124);
and U3978 (N_3978,N_2895,N_2973);
nand U3979 (N_3979,N_2538,N_2460);
and U3980 (N_3980,N_2576,N_2250);
nor U3981 (N_3981,N_2426,N_2214);
nand U3982 (N_3982,N_2621,N_2976);
or U3983 (N_3983,N_2597,N_2900);
nor U3984 (N_3984,N_2251,N_2729);
nor U3985 (N_3985,N_2528,N_2612);
nor U3986 (N_3986,N_2782,N_2678);
and U3987 (N_3987,N_2434,N_2354);
nand U3988 (N_3988,N_2158,N_2412);
nor U3989 (N_3989,N_2889,N_2352);
nor U3990 (N_3990,N_2056,N_2120);
or U3991 (N_3991,N_2353,N_2118);
and U3992 (N_3992,N_2573,N_2762);
or U3993 (N_3993,N_2512,N_2952);
and U3994 (N_3994,N_2529,N_2880);
or U3995 (N_3995,N_2486,N_2453);
nor U3996 (N_3996,N_2290,N_2527);
nand U3997 (N_3997,N_2292,N_2591);
and U3998 (N_3998,N_2564,N_2546);
and U3999 (N_3999,N_2603,N_2082);
and U4000 (N_4000,N_3258,N_3146);
and U4001 (N_4001,N_3044,N_3664);
and U4002 (N_4002,N_3016,N_3915);
nor U4003 (N_4003,N_3432,N_3376);
nand U4004 (N_4004,N_3125,N_3031);
or U4005 (N_4005,N_3035,N_3195);
and U4006 (N_4006,N_3795,N_3947);
and U4007 (N_4007,N_3580,N_3072);
nor U4008 (N_4008,N_3205,N_3637);
or U4009 (N_4009,N_3078,N_3056);
or U4010 (N_4010,N_3365,N_3410);
nand U4011 (N_4011,N_3149,N_3477);
xor U4012 (N_4012,N_3046,N_3228);
or U4013 (N_4013,N_3610,N_3685);
nand U4014 (N_4014,N_3969,N_3647);
and U4015 (N_4015,N_3671,N_3257);
or U4016 (N_4016,N_3511,N_3583);
or U4017 (N_4017,N_3444,N_3897);
or U4018 (N_4018,N_3634,N_3812);
nand U4019 (N_4019,N_3802,N_3550);
or U4020 (N_4020,N_3927,N_3360);
nand U4021 (N_4021,N_3877,N_3931);
nor U4022 (N_4022,N_3279,N_3638);
and U4023 (N_4023,N_3079,N_3199);
or U4024 (N_4024,N_3361,N_3683);
nand U4025 (N_4025,N_3201,N_3000);
or U4026 (N_4026,N_3820,N_3278);
or U4027 (N_4027,N_3521,N_3250);
or U4028 (N_4028,N_3935,N_3472);
nand U4029 (N_4029,N_3467,N_3619);
nor U4030 (N_4030,N_3810,N_3911);
or U4031 (N_4031,N_3468,N_3417);
and U4032 (N_4032,N_3510,N_3402);
or U4033 (N_4033,N_3355,N_3083);
nand U4034 (N_4034,N_3617,N_3964);
nor U4035 (N_4035,N_3682,N_3639);
nand U4036 (N_4036,N_3584,N_3241);
or U4037 (N_4037,N_3729,N_3796);
nor U4038 (N_4038,N_3663,N_3595);
nor U4039 (N_4039,N_3174,N_3641);
and U4040 (N_4040,N_3751,N_3872);
nand U4041 (N_4041,N_3144,N_3272);
and U4042 (N_4042,N_3559,N_3596);
and U4043 (N_4043,N_3309,N_3322);
or U4044 (N_4044,N_3515,N_3570);
nor U4045 (N_4045,N_3932,N_3533);
or U4046 (N_4046,N_3473,N_3073);
nand U4047 (N_4047,N_3508,N_3501);
and U4048 (N_4048,N_3203,N_3134);
nand U4049 (N_4049,N_3577,N_3007);
nor U4050 (N_4050,N_3921,N_3719);
and U4051 (N_4051,N_3691,N_3088);
nor U4052 (N_4052,N_3839,N_3500);
nor U4053 (N_4053,N_3819,N_3319);
nor U4054 (N_4054,N_3995,N_3827);
nand U4055 (N_4055,N_3843,N_3298);
and U4056 (N_4056,N_3037,N_3200);
or U4057 (N_4057,N_3657,N_3367);
and U4058 (N_4058,N_3227,N_3042);
nor U4059 (N_4059,N_3918,N_3741);
nor U4060 (N_4060,N_3136,N_3387);
nand U4061 (N_4061,N_3863,N_3153);
and U4062 (N_4062,N_3717,N_3141);
nor U4063 (N_4063,N_3254,N_3235);
nor U4064 (N_4064,N_3700,N_3749);
nand U4065 (N_4065,N_3513,N_3553);
and U4066 (N_4066,N_3383,N_3736);
or U4067 (N_4067,N_3528,N_3480);
nor U4068 (N_4068,N_3019,N_3434);
nor U4069 (N_4069,N_3522,N_3930);
nor U4070 (N_4070,N_3160,N_3389);
or U4071 (N_4071,N_3373,N_3699);
or U4072 (N_4072,N_3412,N_3068);
and U4073 (N_4073,N_3280,N_3696);
nor U4074 (N_4074,N_3784,N_3652);
and U4075 (N_4075,N_3460,N_3039);
nor U4076 (N_4076,N_3613,N_3494);
or U4077 (N_4077,N_3658,N_3880);
nand U4078 (N_4078,N_3374,N_3773);
and U4079 (N_4079,N_3715,N_3359);
nor U4080 (N_4080,N_3192,N_3456);
nand U4081 (N_4081,N_3133,N_3369);
and U4082 (N_4082,N_3744,N_3447);
nor U4083 (N_4083,N_3966,N_3172);
and U4084 (N_4084,N_3033,N_3164);
or U4085 (N_4085,N_3045,N_3774);
xnor U4086 (N_4086,N_3343,N_3642);
nor U4087 (N_4087,N_3558,N_3535);
or U4088 (N_4088,N_3152,N_3594);
nor U4089 (N_4089,N_3603,N_3600);
or U4090 (N_4090,N_3540,N_3177);
or U4091 (N_4091,N_3529,N_3938);
or U4092 (N_4092,N_3209,N_3173);
nor U4093 (N_4093,N_3453,N_3390);
nor U4094 (N_4094,N_3411,N_3304);
or U4095 (N_4095,N_3159,N_3585);
or U4096 (N_4096,N_3408,N_3093);
and U4097 (N_4097,N_3789,N_3129);
nor U4098 (N_4098,N_3328,N_3628);
or U4099 (N_4099,N_3573,N_3437);
nand U4100 (N_4100,N_3676,N_3800);
or U4101 (N_4101,N_3622,N_3266);
or U4102 (N_4102,N_3106,N_3380);
or U4103 (N_4103,N_3150,N_3770);
and U4104 (N_4104,N_3348,N_3532);
and U4105 (N_4105,N_3009,N_3739);
nand U4106 (N_4106,N_3002,N_3986);
or U4107 (N_4107,N_3024,N_3527);
and U4108 (N_4108,N_3486,N_3344);
and U4109 (N_4109,N_3755,N_3181);
or U4110 (N_4110,N_3689,N_3245);
nand U4111 (N_4111,N_3405,N_3643);
nand U4112 (N_4112,N_3184,N_3640);
and U4113 (N_4113,N_3894,N_3409);
or U4114 (N_4114,N_3779,N_3831);
or U4115 (N_4115,N_3607,N_3858);
nand U4116 (N_4116,N_3169,N_3273);
nor U4117 (N_4117,N_3957,N_3725);
nand U4118 (N_4118,N_3517,N_3026);
and U4119 (N_4119,N_3162,N_3829);
and U4120 (N_4120,N_3615,N_3945);
or U4121 (N_4121,N_3029,N_3051);
nor U4122 (N_4122,N_3463,N_3104);
and U4123 (N_4123,N_3962,N_3197);
nor U4124 (N_4124,N_3507,N_3978);
nand U4125 (N_4125,N_3666,N_3673);
nand U4126 (N_4126,N_3581,N_3759);
nand U4127 (N_4127,N_3520,N_3857);
or U4128 (N_4128,N_3381,N_3660);
nor U4129 (N_4129,N_3208,N_3826);
or U4130 (N_4130,N_3869,N_3994);
or U4131 (N_4131,N_3238,N_3214);
nand U4132 (N_4132,N_3502,N_3289);
nor U4133 (N_4133,N_3653,N_3956);
or U4134 (N_4134,N_3188,N_3860);
or U4135 (N_4135,N_3959,N_3440);
nor U4136 (N_4136,N_3457,N_3909);
nand U4137 (N_4137,N_3972,N_3549);
nand U4138 (N_4138,N_3572,N_3754);
or U4139 (N_4139,N_3384,N_3284);
nand U4140 (N_4140,N_3287,N_3296);
and U4141 (N_4141,N_3526,N_3183);
or U4142 (N_4142,N_3461,N_3096);
nand U4143 (N_4143,N_3782,N_3849);
or U4144 (N_4144,N_3058,N_3870);
or U4145 (N_4145,N_3053,N_3006);
nor U4146 (N_4146,N_3898,N_3108);
and U4147 (N_4147,N_3524,N_3781);
nor U4148 (N_4148,N_3207,N_3998);
nand U4149 (N_4149,N_3264,N_3004);
nand U4150 (N_4150,N_3302,N_3011);
xnor U4151 (N_4151,N_3990,N_3276);
or U4152 (N_4152,N_3155,N_3234);
and U4153 (N_4153,N_3531,N_3377);
nor U4154 (N_4154,N_3455,N_3138);
nand U4155 (N_4155,N_3769,N_3219);
or U4156 (N_4156,N_3459,N_3232);
nor U4157 (N_4157,N_3274,N_3261);
or U4158 (N_4158,N_3593,N_3678);
and U4159 (N_4159,N_3103,N_3038);
nand U4160 (N_4160,N_3623,N_3226);
and U4161 (N_4161,N_3854,N_3441);
and U4162 (N_4162,N_3043,N_3397);
and U4163 (N_4163,N_3742,N_3571);
and U4164 (N_4164,N_3439,N_3886);
nor U4165 (N_4165,N_3283,N_3675);
nor U4166 (N_4166,N_3269,N_3980);
nor U4167 (N_4167,N_3488,N_3358);
nand U4168 (N_4168,N_3332,N_3776);
nor U4169 (N_4169,N_3780,N_3845);
nand U4170 (N_4170,N_3028,N_3589);
nor U4171 (N_4171,N_3430,N_3888);
nor U4172 (N_4172,N_3331,N_3334);
nand U4173 (N_4173,N_3062,N_3327);
and U4174 (N_4174,N_3132,N_3356);
and U4175 (N_4175,N_3885,N_3102);
nor U4176 (N_4176,N_3963,N_3394);
and U4177 (N_4177,N_3148,N_3620);
nand U4178 (N_4178,N_3388,N_3724);
or U4179 (N_4179,N_3080,N_3731);
nor U4180 (N_4180,N_3255,N_3094);
nand U4181 (N_4181,N_3060,N_3307);
and U4182 (N_4182,N_3974,N_3474);
and U4183 (N_4183,N_3801,N_3993);
or U4184 (N_4184,N_3903,N_3342);
nand U4185 (N_4185,N_3242,N_3793);
or U4186 (N_4186,N_3669,N_3868);
and U4187 (N_4187,N_3562,N_3667);
and U4188 (N_4188,N_3875,N_3730);
or U4189 (N_4189,N_3973,N_3575);
and U4190 (N_4190,N_3567,N_3578);
and U4191 (N_4191,N_3421,N_3352);
or U4192 (N_4192,N_3075,N_3005);
nand U4193 (N_4193,N_3720,N_3262);
and U4194 (N_4194,N_3618,N_3896);
and U4195 (N_4195,N_3027,N_3351);
or U4196 (N_4196,N_3196,N_3491);
and U4197 (N_4197,N_3222,N_3100);
nand U4198 (N_4198,N_3713,N_3282);
nand U4199 (N_4199,N_3218,N_3293);
nand U4200 (N_4200,N_3732,N_3621);
or U4201 (N_4201,N_3568,N_3496);
nor U4202 (N_4202,N_3514,N_3300);
and U4203 (N_4203,N_3167,N_3913);
or U4204 (N_4204,N_3465,N_3876);
and U4205 (N_4205,N_3047,N_3010);
nand U4206 (N_4206,N_3345,N_3081);
and U4207 (N_4207,N_3175,N_3895);
and U4208 (N_4208,N_3265,N_3791);
and U4209 (N_4209,N_3224,N_3818);
or U4210 (N_4210,N_3492,N_3335);
and U4211 (N_4211,N_3185,N_3756);
and U4212 (N_4212,N_3709,N_3955);
or U4213 (N_4213,N_3525,N_3151);
nor U4214 (N_4214,N_3023,N_3252);
or U4215 (N_4215,N_3866,N_3889);
nor U4216 (N_4216,N_3069,N_3560);
or U4217 (N_4217,N_3117,N_3059);
and U4218 (N_4218,N_3630,N_3139);
and U4219 (N_4219,N_3182,N_3048);
nor U4220 (N_4220,N_3497,N_3861);
and U4221 (N_4221,N_3569,N_3566);
and U4222 (N_4222,N_3523,N_3418);
nand U4223 (N_4223,N_3143,N_3967);
nor U4224 (N_4224,N_3464,N_3943);
and U4225 (N_4225,N_3881,N_3579);
and U4226 (N_4226,N_3799,N_3760);
and U4227 (N_4227,N_3837,N_3601);
nor U4228 (N_4228,N_3958,N_3020);
nor U4229 (N_4229,N_3592,N_3735);
or U4230 (N_4230,N_3306,N_3764);
and U4231 (N_4231,N_3771,N_3217);
nor U4232 (N_4232,N_3036,N_3061);
nor U4233 (N_4233,N_3767,N_3968);
nand U4234 (N_4234,N_3256,N_3251);
and U4235 (N_4235,N_3611,N_3055);
or U4236 (N_4236,N_3495,N_3299);
nand U4237 (N_4237,N_3711,N_3338);
nand U4238 (N_4238,N_3612,N_3606);
nor U4239 (N_4239,N_3981,N_3576);
or U4240 (N_4240,N_3864,N_3887);
nand U4241 (N_4241,N_3471,N_3018);
and U4242 (N_4242,N_3707,N_3798);
or U4243 (N_4243,N_3672,N_3318);
and U4244 (N_4244,N_3116,N_3314);
nand U4245 (N_4245,N_3120,N_3105);
nand U4246 (N_4246,N_3066,N_3220);
or U4247 (N_4247,N_3248,N_3899);
and U4248 (N_4248,N_3321,N_3427);
or U4249 (N_4249,N_3127,N_3851);
nor U4250 (N_4250,N_3268,N_3324);
or U4251 (N_4251,N_3161,N_3277);
nor U4252 (N_4252,N_3030,N_3215);
and U4253 (N_4253,N_3140,N_3371);
nand U4254 (N_4254,N_3950,N_3662);
nand U4255 (N_4255,N_3705,N_3907);
nand U4256 (N_4256,N_3126,N_3323);
and U4257 (N_4257,N_3454,N_3399);
and U4258 (N_4258,N_3450,N_3170);
nand U4259 (N_4259,N_3362,N_3650);
nand U4260 (N_4260,N_3841,N_3428);
nand U4261 (N_4261,N_3971,N_3537);
nor U4262 (N_4262,N_3003,N_3703);
nand U4263 (N_4263,N_3848,N_3270);
nand U4264 (N_4264,N_3702,N_3121);
nor U4265 (N_4265,N_3659,N_3301);
nand U4266 (N_4266,N_3189,N_3976);
nand U4267 (N_4267,N_3815,N_3239);
nor U4268 (N_4268,N_3554,N_3142);
xor U4269 (N_4269,N_3590,N_3908);
nand U4270 (N_4270,N_3370,N_3924);
nor U4271 (N_4271,N_3404,N_3347);
and U4272 (N_4272,N_3398,N_3704);
nor U4273 (N_4273,N_3015,N_3824);
nor U4274 (N_4274,N_3385,N_3204);
or U4275 (N_4275,N_3415,N_3679);
and U4276 (N_4276,N_3878,N_3237);
nor U4277 (N_4277,N_3563,N_3057);
and U4278 (N_4278,N_3591,N_3194);
or U4279 (N_4279,N_3340,N_3458);
nand U4280 (N_4280,N_3336,N_3288);
nor U4281 (N_4281,N_3263,N_3478);
and U4282 (N_4282,N_3419,N_3506);
or U4283 (N_4283,N_3165,N_3225);
nor U4284 (N_4284,N_3313,N_3814);
or U4285 (N_4285,N_3626,N_3884);
nand U4286 (N_4286,N_3745,N_3443);
or U4287 (N_4287,N_3008,N_3803);
nor U4288 (N_4288,N_3210,N_3844);
nand U4289 (N_4289,N_3750,N_3556);
nand U4290 (N_4290,N_3180,N_3737);
nand U4291 (N_4291,N_3728,N_3838);
and U4292 (N_4292,N_3503,N_3001);
nand U4293 (N_4293,N_3922,N_3822);
nor U4294 (N_4294,N_3113,N_3614);
nor U4295 (N_4295,N_3193,N_3842);
and U4296 (N_4296,N_3244,N_3156);
and U4297 (N_4297,N_3063,N_3052);
nor U4298 (N_4298,N_3902,N_3305);
nor U4299 (N_4299,N_3420,N_3693);
and U4300 (N_4300,N_3763,N_3236);
or U4301 (N_4301,N_3997,N_3413);
nand U4302 (N_4302,N_3633,N_3722);
nand U4303 (N_4303,N_3948,N_3230);
and U4304 (N_4304,N_3953,N_3442);
and U4305 (N_4305,N_3087,N_3539);
nor U4306 (N_4306,N_3176,N_3608);
nor U4307 (N_4307,N_3115,N_3065);
nor U4308 (N_4308,N_3825,N_3716);
or U4309 (N_4309,N_3123,N_3681);
or U4310 (N_4310,N_3012,N_3761);
and U4311 (N_4311,N_3542,N_3768);
nand U4312 (N_4312,N_3191,N_3587);
and U4313 (N_4313,N_3303,N_3988);
or U4314 (N_4314,N_3890,N_3926);
or U4315 (N_4315,N_3656,N_3840);
nand U4316 (N_4316,N_3645,N_3586);
or U4317 (N_4317,N_3687,N_3989);
and U4318 (N_4318,N_3949,N_3014);
and U4319 (N_4319,N_3747,N_3661);
nor U4320 (N_4320,N_3213,N_3695);
and U4321 (N_4321,N_3493,N_3325);
xnor U4322 (N_4322,N_3157,N_3565);
nor U4323 (N_4323,N_3708,N_3723);
nor U4324 (N_4324,N_3740,N_3588);
or U4325 (N_4325,N_3423,N_3564);
nand U4326 (N_4326,N_3112,N_3145);
xnor U4327 (N_4327,N_3905,N_3762);
and U4328 (N_4328,N_3828,N_3834);
or U4329 (N_4329,N_3445,N_3797);
nand U4330 (N_4330,N_3379,N_3936);
or U4331 (N_4331,N_3984,N_3130);
and U4332 (N_4332,N_3677,N_3929);
or U4333 (N_4333,N_3109,N_3847);
nor U4334 (N_4334,N_3476,N_3941);
nor U4335 (N_4335,N_3179,N_3547);
nor U4336 (N_4336,N_3198,N_3786);
or U4337 (N_4337,N_3940,N_3882);
and U4338 (N_4338,N_3766,N_3091);
nor U4339 (N_4339,N_3483,N_3470);
nand U4340 (N_4340,N_3879,N_3900);
nor U4341 (N_4341,N_3285,N_3893);
and U4342 (N_4342,N_3243,N_3424);
nor U4343 (N_4343,N_3710,N_3353);
nor U4344 (N_4344,N_3267,N_3688);
nor U4345 (N_4345,N_3698,N_3050);
and U4346 (N_4346,N_3469,N_3481);
and U4347 (N_4347,N_3946,N_3690);
and U4348 (N_4348,N_3071,N_3375);
and U4349 (N_4349,N_3871,N_3777);
and U4350 (N_4350,N_3498,N_3316);
nor U4351 (N_4351,N_3904,N_3475);
and U4352 (N_4352,N_3906,N_3807);
and U4353 (N_4353,N_3519,N_3386);
nor U4354 (N_4354,N_3317,N_3668);
and U4355 (N_4355,N_3867,N_3308);
nor U4356 (N_4356,N_3937,N_3504);
and U4357 (N_4357,N_3686,N_3901);
nand U4358 (N_4358,N_3122,N_3646);
or U4359 (N_4359,N_3363,N_3557);
and U4360 (N_4360,N_3574,N_3378);
nor U4361 (N_4361,N_3999,N_3281);
nand U4362 (N_4362,N_3808,N_3961);
nor U4363 (N_4363,N_3718,N_3407);
and U4364 (N_4364,N_3357,N_3084);
and U4365 (N_4365,N_3541,N_3823);
nor U4366 (N_4366,N_3097,N_3836);
or U4367 (N_4367,N_3811,N_3022);
nor U4368 (N_4368,N_3499,N_3406);
nor U4369 (N_4369,N_3960,N_3632);
and U4370 (N_4370,N_3670,N_3330);
nor U4371 (N_4371,N_3883,N_3382);
and U4372 (N_4372,N_3712,N_3734);
and U4373 (N_4373,N_3320,N_3655);
nand U4374 (N_4374,N_3787,N_3414);
or U4375 (N_4375,N_3354,N_3605);
nor U4376 (N_4376,N_3326,N_3484);
and U4377 (N_4377,N_3211,N_3543);
or U4378 (N_4378,N_3545,N_3163);
nand U4379 (N_4379,N_3602,N_3433);
nand U4380 (N_4380,N_3403,N_3850);
or U4381 (N_4381,N_3555,N_3977);
nand U4382 (N_4382,N_3933,N_3436);
and U4383 (N_4383,N_3131,N_3505);
nor U4384 (N_4384,N_3101,N_3085);
or U4385 (N_4385,N_3229,N_3431);
nand U4386 (N_4386,N_3916,N_3074);
or U4387 (N_4387,N_3259,N_3778);
and U4388 (N_4388,N_3785,N_3147);
and U4389 (N_4389,N_3862,N_3021);
nand U4390 (N_4390,N_3082,N_3942);
nor U4391 (N_4391,N_3833,N_3462);
and U4392 (N_4392,N_3435,N_3425);
and U4393 (N_4393,N_3721,N_3552);
or U4394 (N_4394,N_3368,N_3939);
and U4395 (N_4395,N_3996,N_3925);
and U4396 (N_4396,N_3853,N_3449);
or U4397 (N_4397,N_3291,N_3312);
nor U4398 (N_4398,N_3516,N_3631);
or U4399 (N_4399,N_3438,N_3598);
and U4400 (N_4400,N_3654,N_3372);
nand U4401 (N_4401,N_3292,N_3190);
or U4402 (N_4402,N_3487,N_3859);
or U4403 (N_4403,N_3090,N_3804);
or U4404 (N_4404,N_3448,N_3706);
and U4405 (N_4405,N_3099,N_3846);
nand U4406 (N_4406,N_3975,N_3536);
or U4407 (N_4407,N_3954,N_3616);
and U4408 (N_4408,N_3538,N_3395);
and U4409 (N_4409,N_3240,N_3231);
nand U4410 (N_4410,N_3098,N_3124);
and U4411 (N_4411,N_3392,N_3089);
or U4412 (N_4412,N_3346,N_3366);
and U4413 (N_4413,N_3067,N_3874);
nand U4414 (N_4414,N_3512,N_3333);
nand U4415 (N_4415,N_3648,N_3393);
or U4416 (N_4416,N_3983,N_3701);
nand U4417 (N_4417,N_3290,N_3790);
or U4418 (N_4418,N_3684,N_3260);
nor U4419 (N_4419,N_3070,N_3114);
nor U4420 (N_4420,N_3212,N_3987);
nand U4421 (N_4421,N_3625,N_3910);
nor U4422 (N_4422,N_3337,N_3758);
nand U4423 (N_4423,N_3223,N_3757);
nor U4424 (N_4424,N_3813,N_3809);
nand U4425 (N_4425,N_3350,N_3530);
nor U4426 (N_4426,N_3253,N_3271);
nor U4427 (N_4427,N_3830,N_3992);
or U4428 (N_4428,N_3216,N_3485);
nand U4429 (N_4429,N_3429,N_3168);
and U4430 (N_4430,N_3119,N_3597);
or U4431 (N_4431,N_3917,N_3714);
or U4432 (N_4432,N_3738,N_3923);
or U4433 (N_4433,N_3752,N_3743);
nand U4434 (N_4434,N_3339,N_3341);
xnor U4435 (N_4435,N_3609,N_3297);
or U4436 (N_4436,N_3599,N_3891);
and U4437 (N_4437,N_3482,N_3979);
and U4438 (N_4438,N_3107,N_3206);
and U4439 (N_4439,N_3509,N_3128);
and U4440 (N_4440,N_3233,N_3040);
and U4441 (N_4441,N_3746,N_3865);
nand U4442 (N_4442,N_3158,N_3991);
and U4443 (N_4443,N_3951,N_3928);
and U4444 (N_4444,N_3783,N_3013);
nand U4445 (N_4445,N_3086,N_3171);
or U4446 (N_4446,N_3873,N_3692);
nand U4447 (N_4447,N_3364,N_3794);
nand U4448 (N_4448,N_3805,N_3855);
nand U4449 (N_4449,N_3644,N_3892);
or U4450 (N_4450,N_3118,N_3111);
nor U4451 (N_4451,N_3772,N_3806);
nor U4452 (N_4452,N_3315,N_3154);
or U4453 (N_4453,N_3775,N_3635);
nand U4454 (N_4454,N_3032,N_3534);
and U4455 (N_4455,N_3110,N_3310);
or U4456 (N_4456,N_3726,N_3391);
xor U4457 (N_4457,N_3479,N_3246);
or U4458 (N_4458,N_3649,N_3422);
nand U4459 (N_4459,N_3748,N_3852);
nor U4460 (N_4460,N_3095,N_3680);
nand U4461 (N_4461,N_3137,N_3651);
and U4462 (N_4462,N_3187,N_3604);
and U4463 (N_4463,N_3636,N_3311);
nand U4464 (N_4464,N_3416,N_3166);
nor U4465 (N_4465,N_3466,N_3697);
and U4466 (N_4466,N_3753,N_3912);
nor U4467 (N_4467,N_3982,N_3396);
nand U4468 (N_4468,N_3451,N_3546);
or U4469 (N_4469,N_3490,N_3076);
nand U4470 (N_4470,N_3624,N_3054);
and U4471 (N_4471,N_3446,N_3400);
nor U4472 (N_4472,N_3816,N_3452);
or U4473 (N_4473,N_3295,N_3275);
nand U4474 (N_4474,N_3286,N_3186);
and U4475 (N_4475,N_3629,N_3092);
and U4476 (N_4476,N_3727,N_3856);
nor U4477 (N_4477,N_3249,N_3401);
nand U4478 (N_4478,N_3965,N_3178);
and U4479 (N_4479,N_3920,N_3952);
and U4480 (N_4480,N_3561,N_3788);
or U4481 (N_4481,N_3985,N_3970);
and U4482 (N_4482,N_3551,N_3919);
and U4483 (N_4483,N_3934,N_3518);
nand U4484 (N_4484,N_3914,N_3221);
nor U4485 (N_4485,N_3064,N_3247);
or U4486 (N_4486,N_3202,N_3832);
nor U4487 (N_4487,N_3944,N_3765);
nand U4488 (N_4488,N_3135,N_3077);
and U4489 (N_4489,N_3017,N_3821);
or U4490 (N_4490,N_3426,N_3582);
nor U4491 (N_4491,N_3548,N_3049);
and U4492 (N_4492,N_3817,N_3694);
nand U4493 (N_4493,N_3665,N_3349);
and U4494 (N_4494,N_3294,N_3544);
nand U4495 (N_4495,N_3489,N_3329);
and U4496 (N_4496,N_3034,N_3674);
or U4497 (N_4497,N_3627,N_3025);
nand U4498 (N_4498,N_3835,N_3792);
or U4499 (N_4499,N_3041,N_3733);
nor U4500 (N_4500,N_3500,N_3661);
or U4501 (N_4501,N_3913,N_3868);
nand U4502 (N_4502,N_3812,N_3708);
and U4503 (N_4503,N_3657,N_3091);
nor U4504 (N_4504,N_3161,N_3453);
or U4505 (N_4505,N_3832,N_3170);
nand U4506 (N_4506,N_3067,N_3912);
nand U4507 (N_4507,N_3832,N_3591);
or U4508 (N_4508,N_3671,N_3878);
or U4509 (N_4509,N_3941,N_3498);
nor U4510 (N_4510,N_3358,N_3628);
or U4511 (N_4511,N_3501,N_3662);
xor U4512 (N_4512,N_3452,N_3020);
or U4513 (N_4513,N_3713,N_3665);
nor U4514 (N_4514,N_3152,N_3922);
or U4515 (N_4515,N_3840,N_3279);
nor U4516 (N_4516,N_3278,N_3156);
and U4517 (N_4517,N_3536,N_3406);
and U4518 (N_4518,N_3486,N_3392);
or U4519 (N_4519,N_3444,N_3057);
and U4520 (N_4520,N_3897,N_3286);
nand U4521 (N_4521,N_3628,N_3034);
or U4522 (N_4522,N_3193,N_3560);
nor U4523 (N_4523,N_3188,N_3145);
or U4524 (N_4524,N_3941,N_3634);
and U4525 (N_4525,N_3924,N_3428);
nand U4526 (N_4526,N_3484,N_3427);
and U4527 (N_4527,N_3102,N_3533);
nand U4528 (N_4528,N_3844,N_3120);
nor U4529 (N_4529,N_3614,N_3932);
nand U4530 (N_4530,N_3706,N_3170);
nand U4531 (N_4531,N_3111,N_3242);
and U4532 (N_4532,N_3614,N_3742);
nor U4533 (N_4533,N_3617,N_3250);
and U4534 (N_4534,N_3403,N_3641);
nor U4535 (N_4535,N_3389,N_3211);
and U4536 (N_4536,N_3360,N_3740);
or U4537 (N_4537,N_3055,N_3784);
or U4538 (N_4538,N_3096,N_3479);
nand U4539 (N_4539,N_3892,N_3898);
or U4540 (N_4540,N_3103,N_3905);
or U4541 (N_4541,N_3779,N_3265);
nor U4542 (N_4542,N_3780,N_3766);
nor U4543 (N_4543,N_3602,N_3770);
and U4544 (N_4544,N_3183,N_3894);
nor U4545 (N_4545,N_3942,N_3029);
nor U4546 (N_4546,N_3594,N_3516);
nor U4547 (N_4547,N_3878,N_3641);
nor U4548 (N_4548,N_3422,N_3973);
nor U4549 (N_4549,N_3702,N_3583);
nor U4550 (N_4550,N_3760,N_3514);
nor U4551 (N_4551,N_3545,N_3947);
nor U4552 (N_4552,N_3790,N_3517);
nor U4553 (N_4553,N_3043,N_3317);
nand U4554 (N_4554,N_3350,N_3535);
or U4555 (N_4555,N_3340,N_3040);
nand U4556 (N_4556,N_3483,N_3135);
and U4557 (N_4557,N_3540,N_3750);
or U4558 (N_4558,N_3885,N_3435);
or U4559 (N_4559,N_3732,N_3573);
and U4560 (N_4560,N_3135,N_3602);
nor U4561 (N_4561,N_3055,N_3349);
or U4562 (N_4562,N_3595,N_3674);
nand U4563 (N_4563,N_3426,N_3475);
nor U4564 (N_4564,N_3961,N_3867);
or U4565 (N_4565,N_3272,N_3446);
nor U4566 (N_4566,N_3433,N_3262);
and U4567 (N_4567,N_3298,N_3956);
nor U4568 (N_4568,N_3931,N_3843);
and U4569 (N_4569,N_3355,N_3117);
or U4570 (N_4570,N_3296,N_3355);
or U4571 (N_4571,N_3264,N_3349);
nor U4572 (N_4572,N_3933,N_3738);
or U4573 (N_4573,N_3942,N_3744);
nor U4574 (N_4574,N_3723,N_3515);
and U4575 (N_4575,N_3279,N_3474);
nand U4576 (N_4576,N_3886,N_3384);
and U4577 (N_4577,N_3297,N_3173);
or U4578 (N_4578,N_3987,N_3901);
or U4579 (N_4579,N_3930,N_3743);
nand U4580 (N_4580,N_3489,N_3327);
or U4581 (N_4581,N_3622,N_3274);
nor U4582 (N_4582,N_3915,N_3002);
nor U4583 (N_4583,N_3083,N_3414);
nand U4584 (N_4584,N_3141,N_3844);
nand U4585 (N_4585,N_3928,N_3385);
or U4586 (N_4586,N_3733,N_3528);
xor U4587 (N_4587,N_3793,N_3939);
or U4588 (N_4588,N_3238,N_3628);
nor U4589 (N_4589,N_3509,N_3247);
or U4590 (N_4590,N_3340,N_3779);
nand U4591 (N_4591,N_3081,N_3501);
and U4592 (N_4592,N_3798,N_3408);
or U4593 (N_4593,N_3110,N_3909);
or U4594 (N_4594,N_3272,N_3055);
nand U4595 (N_4595,N_3767,N_3055);
nor U4596 (N_4596,N_3115,N_3045);
nand U4597 (N_4597,N_3628,N_3056);
or U4598 (N_4598,N_3274,N_3435);
or U4599 (N_4599,N_3916,N_3031);
or U4600 (N_4600,N_3340,N_3116);
and U4601 (N_4601,N_3641,N_3137);
and U4602 (N_4602,N_3684,N_3784);
and U4603 (N_4603,N_3246,N_3138);
or U4604 (N_4604,N_3842,N_3013);
nand U4605 (N_4605,N_3045,N_3558);
nor U4606 (N_4606,N_3758,N_3687);
or U4607 (N_4607,N_3484,N_3443);
or U4608 (N_4608,N_3550,N_3661);
and U4609 (N_4609,N_3026,N_3699);
nand U4610 (N_4610,N_3693,N_3827);
and U4611 (N_4611,N_3485,N_3566);
or U4612 (N_4612,N_3477,N_3627);
nand U4613 (N_4613,N_3104,N_3905);
or U4614 (N_4614,N_3575,N_3494);
and U4615 (N_4615,N_3302,N_3599);
or U4616 (N_4616,N_3777,N_3152);
and U4617 (N_4617,N_3869,N_3567);
and U4618 (N_4618,N_3284,N_3676);
or U4619 (N_4619,N_3421,N_3484);
or U4620 (N_4620,N_3042,N_3098);
and U4621 (N_4621,N_3621,N_3759);
nand U4622 (N_4622,N_3776,N_3026);
nand U4623 (N_4623,N_3816,N_3647);
or U4624 (N_4624,N_3357,N_3045);
nand U4625 (N_4625,N_3547,N_3931);
or U4626 (N_4626,N_3606,N_3452);
nor U4627 (N_4627,N_3484,N_3295);
nor U4628 (N_4628,N_3075,N_3655);
nor U4629 (N_4629,N_3625,N_3542);
nor U4630 (N_4630,N_3536,N_3281);
and U4631 (N_4631,N_3852,N_3909);
nor U4632 (N_4632,N_3626,N_3378);
or U4633 (N_4633,N_3505,N_3402);
and U4634 (N_4634,N_3792,N_3922);
and U4635 (N_4635,N_3317,N_3045);
or U4636 (N_4636,N_3271,N_3997);
nor U4637 (N_4637,N_3204,N_3337);
and U4638 (N_4638,N_3409,N_3952);
or U4639 (N_4639,N_3508,N_3399);
and U4640 (N_4640,N_3984,N_3247);
nor U4641 (N_4641,N_3007,N_3055);
nand U4642 (N_4642,N_3039,N_3059);
and U4643 (N_4643,N_3950,N_3192);
or U4644 (N_4644,N_3068,N_3024);
or U4645 (N_4645,N_3899,N_3709);
nand U4646 (N_4646,N_3208,N_3671);
nor U4647 (N_4647,N_3150,N_3642);
nor U4648 (N_4648,N_3955,N_3279);
or U4649 (N_4649,N_3692,N_3069);
and U4650 (N_4650,N_3603,N_3337);
or U4651 (N_4651,N_3051,N_3294);
nor U4652 (N_4652,N_3127,N_3163);
and U4653 (N_4653,N_3471,N_3073);
nand U4654 (N_4654,N_3055,N_3169);
or U4655 (N_4655,N_3065,N_3462);
or U4656 (N_4656,N_3949,N_3243);
nand U4657 (N_4657,N_3329,N_3650);
nand U4658 (N_4658,N_3158,N_3210);
nor U4659 (N_4659,N_3704,N_3991);
and U4660 (N_4660,N_3486,N_3964);
or U4661 (N_4661,N_3137,N_3779);
and U4662 (N_4662,N_3649,N_3423);
nor U4663 (N_4663,N_3225,N_3620);
nor U4664 (N_4664,N_3947,N_3723);
nand U4665 (N_4665,N_3368,N_3473);
or U4666 (N_4666,N_3096,N_3271);
nand U4667 (N_4667,N_3240,N_3423);
and U4668 (N_4668,N_3260,N_3509);
and U4669 (N_4669,N_3182,N_3177);
and U4670 (N_4670,N_3774,N_3031);
nor U4671 (N_4671,N_3624,N_3472);
nor U4672 (N_4672,N_3166,N_3330);
nor U4673 (N_4673,N_3242,N_3812);
or U4674 (N_4674,N_3330,N_3715);
nor U4675 (N_4675,N_3260,N_3418);
or U4676 (N_4676,N_3957,N_3038);
nor U4677 (N_4677,N_3573,N_3417);
nor U4678 (N_4678,N_3451,N_3973);
xor U4679 (N_4679,N_3456,N_3116);
nor U4680 (N_4680,N_3537,N_3591);
nor U4681 (N_4681,N_3645,N_3580);
or U4682 (N_4682,N_3650,N_3150);
nor U4683 (N_4683,N_3242,N_3183);
nor U4684 (N_4684,N_3244,N_3953);
or U4685 (N_4685,N_3442,N_3834);
nand U4686 (N_4686,N_3391,N_3242);
or U4687 (N_4687,N_3264,N_3965);
nor U4688 (N_4688,N_3451,N_3746);
nor U4689 (N_4689,N_3677,N_3302);
nand U4690 (N_4690,N_3764,N_3277);
nand U4691 (N_4691,N_3769,N_3504);
or U4692 (N_4692,N_3181,N_3296);
nor U4693 (N_4693,N_3191,N_3137);
nor U4694 (N_4694,N_3415,N_3663);
nor U4695 (N_4695,N_3856,N_3756);
or U4696 (N_4696,N_3175,N_3074);
and U4697 (N_4697,N_3785,N_3251);
nand U4698 (N_4698,N_3831,N_3855);
or U4699 (N_4699,N_3779,N_3063);
and U4700 (N_4700,N_3890,N_3337);
and U4701 (N_4701,N_3001,N_3669);
or U4702 (N_4702,N_3129,N_3657);
or U4703 (N_4703,N_3155,N_3880);
xnor U4704 (N_4704,N_3347,N_3564);
nor U4705 (N_4705,N_3871,N_3784);
or U4706 (N_4706,N_3711,N_3714);
nor U4707 (N_4707,N_3019,N_3597);
or U4708 (N_4708,N_3557,N_3913);
nor U4709 (N_4709,N_3520,N_3476);
or U4710 (N_4710,N_3174,N_3709);
or U4711 (N_4711,N_3447,N_3036);
and U4712 (N_4712,N_3266,N_3918);
nand U4713 (N_4713,N_3789,N_3786);
nand U4714 (N_4714,N_3624,N_3031);
and U4715 (N_4715,N_3877,N_3571);
or U4716 (N_4716,N_3555,N_3734);
nand U4717 (N_4717,N_3319,N_3067);
nor U4718 (N_4718,N_3852,N_3078);
nand U4719 (N_4719,N_3431,N_3633);
nand U4720 (N_4720,N_3067,N_3244);
nor U4721 (N_4721,N_3617,N_3079);
nor U4722 (N_4722,N_3223,N_3910);
nand U4723 (N_4723,N_3709,N_3009);
nor U4724 (N_4724,N_3603,N_3813);
and U4725 (N_4725,N_3317,N_3026);
or U4726 (N_4726,N_3238,N_3412);
nand U4727 (N_4727,N_3422,N_3124);
or U4728 (N_4728,N_3773,N_3504);
and U4729 (N_4729,N_3816,N_3481);
and U4730 (N_4730,N_3580,N_3708);
nor U4731 (N_4731,N_3692,N_3033);
and U4732 (N_4732,N_3320,N_3843);
and U4733 (N_4733,N_3292,N_3668);
and U4734 (N_4734,N_3064,N_3531);
or U4735 (N_4735,N_3434,N_3003);
and U4736 (N_4736,N_3912,N_3450);
nor U4737 (N_4737,N_3539,N_3936);
or U4738 (N_4738,N_3490,N_3637);
nor U4739 (N_4739,N_3400,N_3402);
or U4740 (N_4740,N_3035,N_3909);
or U4741 (N_4741,N_3104,N_3041);
nor U4742 (N_4742,N_3089,N_3524);
and U4743 (N_4743,N_3422,N_3481);
nor U4744 (N_4744,N_3907,N_3987);
nand U4745 (N_4745,N_3953,N_3502);
nand U4746 (N_4746,N_3686,N_3289);
nand U4747 (N_4747,N_3088,N_3176);
nor U4748 (N_4748,N_3982,N_3787);
nor U4749 (N_4749,N_3564,N_3059);
nand U4750 (N_4750,N_3146,N_3527);
and U4751 (N_4751,N_3378,N_3459);
nor U4752 (N_4752,N_3151,N_3569);
nand U4753 (N_4753,N_3471,N_3833);
and U4754 (N_4754,N_3565,N_3926);
nand U4755 (N_4755,N_3751,N_3072);
and U4756 (N_4756,N_3036,N_3448);
and U4757 (N_4757,N_3457,N_3687);
nand U4758 (N_4758,N_3178,N_3919);
nand U4759 (N_4759,N_3585,N_3189);
nand U4760 (N_4760,N_3648,N_3060);
and U4761 (N_4761,N_3826,N_3069);
or U4762 (N_4762,N_3069,N_3544);
nand U4763 (N_4763,N_3015,N_3370);
nor U4764 (N_4764,N_3072,N_3532);
nand U4765 (N_4765,N_3539,N_3581);
nand U4766 (N_4766,N_3107,N_3818);
nand U4767 (N_4767,N_3491,N_3846);
or U4768 (N_4768,N_3770,N_3870);
or U4769 (N_4769,N_3374,N_3381);
and U4770 (N_4770,N_3268,N_3221);
and U4771 (N_4771,N_3483,N_3194);
and U4772 (N_4772,N_3400,N_3849);
and U4773 (N_4773,N_3479,N_3615);
and U4774 (N_4774,N_3006,N_3068);
and U4775 (N_4775,N_3388,N_3552);
and U4776 (N_4776,N_3642,N_3676);
nand U4777 (N_4777,N_3145,N_3020);
nand U4778 (N_4778,N_3804,N_3581);
nor U4779 (N_4779,N_3633,N_3266);
nor U4780 (N_4780,N_3693,N_3109);
nand U4781 (N_4781,N_3535,N_3449);
and U4782 (N_4782,N_3602,N_3581);
nor U4783 (N_4783,N_3840,N_3930);
nor U4784 (N_4784,N_3187,N_3618);
or U4785 (N_4785,N_3874,N_3687);
nand U4786 (N_4786,N_3589,N_3594);
or U4787 (N_4787,N_3814,N_3509);
or U4788 (N_4788,N_3388,N_3378);
nand U4789 (N_4789,N_3977,N_3784);
nand U4790 (N_4790,N_3359,N_3127);
or U4791 (N_4791,N_3798,N_3862);
and U4792 (N_4792,N_3846,N_3837);
nor U4793 (N_4793,N_3642,N_3909);
nor U4794 (N_4794,N_3588,N_3904);
and U4795 (N_4795,N_3314,N_3597);
nand U4796 (N_4796,N_3262,N_3618);
or U4797 (N_4797,N_3864,N_3177);
nand U4798 (N_4798,N_3364,N_3704);
or U4799 (N_4799,N_3537,N_3281);
nand U4800 (N_4800,N_3832,N_3687);
nand U4801 (N_4801,N_3296,N_3765);
and U4802 (N_4802,N_3611,N_3779);
or U4803 (N_4803,N_3879,N_3988);
and U4804 (N_4804,N_3412,N_3731);
nand U4805 (N_4805,N_3402,N_3706);
or U4806 (N_4806,N_3665,N_3581);
and U4807 (N_4807,N_3541,N_3144);
nor U4808 (N_4808,N_3788,N_3807);
nand U4809 (N_4809,N_3747,N_3856);
nand U4810 (N_4810,N_3969,N_3937);
and U4811 (N_4811,N_3871,N_3655);
or U4812 (N_4812,N_3173,N_3160);
nand U4813 (N_4813,N_3094,N_3967);
or U4814 (N_4814,N_3177,N_3647);
nand U4815 (N_4815,N_3375,N_3602);
or U4816 (N_4816,N_3094,N_3719);
and U4817 (N_4817,N_3167,N_3151);
nor U4818 (N_4818,N_3569,N_3763);
and U4819 (N_4819,N_3556,N_3092);
nor U4820 (N_4820,N_3733,N_3001);
nor U4821 (N_4821,N_3610,N_3126);
nand U4822 (N_4822,N_3617,N_3435);
nand U4823 (N_4823,N_3495,N_3829);
nand U4824 (N_4824,N_3792,N_3073);
nor U4825 (N_4825,N_3863,N_3062);
nor U4826 (N_4826,N_3768,N_3402);
nand U4827 (N_4827,N_3462,N_3572);
nand U4828 (N_4828,N_3676,N_3660);
and U4829 (N_4829,N_3898,N_3400);
and U4830 (N_4830,N_3268,N_3872);
nand U4831 (N_4831,N_3922,N_3990);
or U4832 (N_4832,N_3458,N_3037);
nand U4833 (N_4833,N_3397,N_3446);
and U4834 (N_4834,N_3246,N_3006);
and U4835 (N_4835,N_3864,N_3307);
and U4836 (N_4836,N_3622,N_3911);
and U4837 (N_4837,N_3580,N_3517);
nor U4838 (N_4838,N_3303,N_3861);
nor U4839 (N_4839,N_3566,N_3653);
nand U4840 (N_4840,N_3768,N_3171);
or U4841 (N_4841,N_3805,N_3899);
or U4842 (N_4842,N_3572,N_3206);
or U4843 (N_4843,N_3549,N_3108);
nor U4844 (N_4844,N_3066,N_3098);
nand U4845 (N_4845,N_3074,N_3945);
or U4846 (N_4846,N_3526,N_3976);
and U4847 (N_4847,N_3298,N_3732);
and U4848 (N_4848,N_3871,N_3987);
nand U4849 (N_4849,N_3307,N_3277);
or U4850 (N_4850,N_3840,N_3979);
nand U4851 (N_4851,N_3209,N_3485);
nand U4852 (N_4852,N_3619,N_3959);
nand U4853 (N_4853,N_3263,N_3589);
and U4854 (N_4854,N_3406,N_3953);
and U4855 (N_4855,N_3792,N_3382);
nand U4856 (N_4856,N_3319,N_3414);
nand U4857 (N_4857,N_3662,N_3676);
or U4858 (N_4858,N_3218,N_3024);
and U4859 (N_4859,N_3414,N_3651);
or U4860 (N_4860,N_3772,N_3240);
or U4861 (N_4861,N_3559,N_3439);
nor U4862 (N_4862,N_3554,N_3969);
nand U4863 (N_4863,N_3636,N_3205);
nor U4864 (N_4864,N_3694,N_3112);
and U4865 (N_4865,N_3464,N_3090);
nor U4866 (N_4866,N_3294,N_3591);
and U4867 (N_4867,N_3518,N_3653);
or U4868 (N_4868,N_3642,N_3382);
or U4869 (N_4869,N_3892,N_3895);
nor U4870 (N_4870,N_3487,N_3761);
nor U4871 (N_4871,N_3338,N_3241);
xnor U4872 (N_4872,N_3587,N_3052);
nor U4873 (N_4873,N_3310,N_3361);
and U4874 (N_4874,N_3124,N_3854);
nand U4875 (N_4875,N_3072,N_3628);
and U4876 (N_4876,N_3525,N_3758);
nor U4877 (N_4877,N_3123,N_3805);
xnor U4878 (N_4878,N_3796,N_3301);
nor U4879 (N_4879,N_3350,N_3900);
nand U4880 (N_4880,N_3118,N_3139);
nand U4881 (N_4881,N_3900,N_3401);
and U4882 (N_4882,N_3494,N_3604);
nand U4883 (N_4883,N_3016,N_3665);
or U4884 (N_4884,N_3707,N_3982);
and U4885 (N_4885,N_3166,N_3573);
or U4886 (N_4886,N_3661,N_3871);
and U4887 (N_4887,N_3272,N_3701);
or U4888 (N_4888,N_3508,N_3749);
nor U4889 (N_4889,N_3598,N_3290);
nor U4890 (N_4890,N_3357,N_3281);
and U4891 (N_4891,N_3823,N_3691);
nand U4892 (N_4892,N_3689,N_3158);
and U4893 (N_4893,N_3477,N_3342);
xor U4894 (N_4894,N_3182,N_3849);
nor U4895 (N_4895,N_3666,N_3571);
nand U4896 (N_4896,N_3760,N_3015);
nand U4897 (N_4897,N_3305,N_3942);
and U4898 (N_4898,N_3007,N_3727);
xnor U4899 (N_4899,N_3462,N_3400);
or U4900 (N_4900,N_3141,N_3931);
or U4901 (N_4901,N_3271,N_3329);
or U4902 (N_4902,N_3046,N_3836);
and U4903 (N_4903,N_3173,N_3926);
nor U4904 (N_4904,N_3725,N_3533);
nor U4905 (N_4905,N_3085,N_3488);
xor U4906 (N_4906,N_3778,N_3535);
nand U4907 (N_4907,N_3226,N_3244);
or U4908 (N_4908,N_3563,N_3122);
nor U4909 (N_4909,N_3742,N_3838);
nand U4910 (N_4910,N_3042,N_3794);
nand U4911 (N_4911,N_3166,N_3703);
nand U4912 (N_4912,N_3611,N_3637);
or U4913 (N_4913,N_3391,N_3926);
or U4914 (N_4914,N_3764,N_3386);
and U4915 (N_4915,N_3698,N_3670);
or U4916 (N_4916,N_3708,N_3503);
nand U4917 (N_4917,N_3680,N_3798);
nor U4918 (N_4918,N_3301,N_3162);
nor U4919 (N_4919,N_3410,N_3612);
nor U4920 (N_4920,N_3219,N_3675);
or U4921 (N_4921,N_3788,N_3671);
and U4922 (N_4922,N_3479,N_3599);
and U4923 (N_4923,N_3114,N_3247);
nor U4924 (N_4924,N_3807,N_3516);
nor U4925 (N_4925,N_3177,N_3597);
or U4926 (N_4926,N_3799,N_3552);
or U4927 (N_4927,N_3907,N_3301);
and U4928 (N_4928,N_3154,N_3701);
and U4929 (N_4929,N_3909,N_3467);
nor U4930 (N_4930,N_3431,N_3563);
nand U4931 (N_4931,N_3567,N_3272);
nor U4932 (N_4932,N_3418,N_3774);
nor U4933 (N_4933,N_3092,N_3481);
nand U4934 (N_4934,N_3943,N_3636);
nand U4935 (N_4935,N_3211,N_3997);
nor U4936 (N_4936,N_3266,N_3413);
and U4937 (N_4937,N_3789,N_3046);
or U4938 (N_4938,N_3476,N_3501);
nor U4939 (N_4939,N_3616,N_3758);
nor U4940 (N_4940,N_3006,N_3789);
nor U4941 (N_4941,N_3924,N_3482);
nand U4942 (N_4942,N_3711,N_3624);
xor U4943 (N_4943,N_3059,N_3955);
xnor U4944 (N_4944,N_3204,N_3426);
or U4945 (N_4945,N_3378,N_3259);
nand U4946 (N_4946,N_3974,N_3114);
nor U4947 (N_4947,N_3498,N_3140);
nor U4948 (N_4948,N_3657,N_3936);
nor U4949 (N_4949,N_3902,N_3197);
nand U4950 (N_4950,N_3582,N_3394);
xnor U4951 (N_4951,N_3437,N_3832);
nand U4952 (N_4952,N_3669,N_3569);
or U4953 (N_4953,N_3967,N_3475);
nand U4954 (N_4954,N_3911,N_3875);
nand U4955 (N_4955,N_3876,N_3119);
or U4956 (N_4956,N_3483,N_3932);
nand U4957 (N_4957,N_3132,N_3330);
nand U4958 (N_4958,N_3056,N_3086);
and U4959 (N_4959,N_3442,N_3787);
or U4960 (N_4960,N_3170,N_3820);
nor U4961 (N_4961,N_3153,N_3988);
or U4962 (N_4962,N_3579,N_3591);
and U4963 (N_4963,N_3030,N_3752);
or U4964 (N_4964,N_3160,N_3993);
or U4965 (N_4965,N_3305,N_3966);
nor U4966 (N_4966,N_3957,N_3658);
and U4967 (N_4967,N_3221,N_3359);
or U4968 (N_4968,N_3205,N_3778);
nand U4969 (N_4969,N_3033,N_3693);
nor U4970 (N_4970,N_3658,N_3811);
and U4971 (N_4971,N_3028,N_3977);
or U4972 (N_4972,N_3056,N_3491);
nor U4973 (N_4973,N_3252,N_3409);
and U4974 (N_4974,N_3445,N_3278);
nor U4975 (N_4975,N_3806,N_3948);
nor U4976 (N_4976,N_3797,N_3179);
nand U4977 (N_4977,N_3545,N_3161);
or U4978 (N_4978,N_3014,N_3846);
nor U4979 (N_4979,N_3052,N_3059);
nand U4980 (N_4980,N_3114,N_3078);
nor U4981 (N_4981,N_3060,N_3554);
and U4982 (N_4982,N_3413,N_3031);
nand U4983 (N_4983,N_3321,N_3762);
nand U4984 (N_4984,N_3196,N_3399);
nand U4985 (N_4985,N_3807,N_3471);
nor U4986 (N_4986,N_3857,N_3095);
or U4987 (N_4987,N_3087,N_3959);
or U4988 (N_4988,N_3240,N_3598);
nand U4989 (N_4989,N_3446,N_3769);
or U4990 (N_4990,N_3624,N_3486);
nor U4991 (N_4991,N_3545,N_3423);
nor U4992 (N_4992,N_3169,N_3537);
nor U4993 (N_4993,N_3612,N_3603);
and U4994 (N_4994,N_3134,N_3116);
nand U4995 (N_4995,N_3754,N_3088);
nand U4996 (N_4996,N_3105,N_3318);
or U4997 (N_4997,N_3541,N_3188);
nor U4998 (N_4998,N_3126,N_3601);
or U4999 (N_4999,N_3687,N_3281);
or U5000 (N_5000,N_4322,N_4516);
nand U5001 (N_5001,N_4748,N_4009);
and U5002 (N_5002,N_4915,N_4665);
nor U5003 (N_5003,N_4502,N_4415);
nor U5004 (N_5004,N_4115,N_4882);
and U5005 (N_5005,N_4329,N_4035);
nand U5006 (N_5006,N_4313,N_4282);
and U5007 (N_5007,N_4142,N_4382);
nand U5008 (N_5008,N_4623,N_4640);
nand U5009 (N_5009,N_4067,N_4480);
nor U5010 (N_5010,N_4116,N_4332);
nand U5011 (N_5011,N_4759,N_4397);
or U5012 (N_5012,N_4511,N_4696);
nand U5013 (N_5013,N_4834,N_4504);
nand U5014 (N_5014,N_4580,N_4464);
nand U5015 (N_5015,N_4596,N_4838);
and U5016 (N_5016,N_4992,N_4004);
nand U5017 (N_5017,N_4199,N_4242);
nand U5018 (N_5018,N_4751,N_4721);
or U5019 (N_5019,N_4565,N_4019);
or U5020 (N_5020,N_4837,N_4222);
nand U5021 (N_5021,N_4750,N_4600);
and U5022 (N_5022,N_4508,N_4878);
and U5023 (N_5023,N_4051,N_4978);
or U5024 (N_5024,N_4538,N_4128);
or U5025 (N_5025,N_4096,N_4149);
and U5026 (N_5026,N_4003,N_4324);
or U5027 (N_5027,N_4920,N_4496);
nor U5028 (N_5028,N_4688,N_4797);
nor U5029 (N_5029,N_4798,N_4077);
nand U5030 (N_5030,N_4576,N_4917);
or U5031 (N_5031,N_4219,N_4767);
nand U5032 (N_5032,N_4377,N_4432);
or U5033 (N_5033,N_4740,N_4579);
nor U5034 (N_5034,N_4131,N_4409);
nor U5035 (N_5035,N_4652,N_4501);
nor U5036 (N_5036,N_4715,N_4490);
nor U5037 (N_5037,N_4606,N_4791);
and U5038 (N_5038,N_4065,N_4593);
nor U5039 (N_5039,N_4162,N_4817);
and U5040 (N_5040,N_4050,N_4459);
nand U5041 (N_5041,N_4426,N_4028);
nor U5042 (N_5042,N_4530,N_4154);
nor U5043 (N_5043,N_4279,N_4577);
or U5044 (N_5044,N_4477,N_4705);
or U5045 (N_5045,N_4616,N_4068);
or U5046 (N_5046,N_4520,N_4972);
nand U5047 (N_5047,N_4165,N_4047);
nor U5048 (N_5048,N_4239,N_4746);
and U5049 (N_5049,N_4533,N_4308);
nor U5050 (N_5050,N_4618,N_4930);
nand U5051 (N_5051,N_4012,N_4395);
or U5052 (N_5052,N_4626,N_4996);
nor U5053 (N_5053,N_4095,N_4515);
and U5054 (N_5054,N_4947,N_4301);
nand U5055 (N_5055,N_4120,N_4356);
nand U5056 (N_5056,N_4264,N_4923);
and U5057 (N_5057,N_4657,N_4584);
and U5058 (N_5058,N_4566,N_4543);
nor U5059 (N_5059,N_4697,N_4921);
xnor U5060 (N_5060,N_4729,N_4505);
nand U5061 (N_5061,N_4205,N_4429);
or U5062 (N_5062,N_4857,N_4692);
and U5063 (N_5063,N_4621,N_4663);
and U5064 (N_5064,N_4266,N_4155);
or U5065 (N_5065,N_4870,N_4995);
or U5066 (N_5066,N_4387,N_4331);
or U5067 (N_5067,N_4014,N_4918);
and U5068 (N_5068,N_4603,N_4192);
or U5069 (N_5069,N_4981,N_4320);
or U5070 (N_5070,N_4206,N_4934);
xor U5071 (N_5071,N_4103,N_4368);
nand U5072 (N_5072,N_4380,N_4755);
nand U5073 (N_5073,N_4762,N_4107);
nor U5074 (N_5074,N_4772,N_4583);
or U5075 (N_5075,N_4255,N_4300);
and U5076 (N_5076,N_4777,N_4716);
nor U5077 (N_5077,N_4273,N_4805);
nor U5078 (N_5078,N_4269,N_4246);
or U5079 (N_5079,N_4720,N_4902);
or U5080 (N_5080,N_4234,N_4080);
nor U5081 (N_5081,N_4243,N_4043);
or U5082 (N_5082,N_4061,N_4421);
and U5083 (N_5083,N_4253,N_4754);
nor U5084 (N_5084,N_4653,N_4156);
nand U5085 (N_5085,N_4910,N_4202);
nand U5086 (N_5086,N_4851,N_4275);
or U5087 (N_5087,N_4561,N_4430);
or U5088 (N_5088,N_4178,N_4304);
or U5089 (N_5089,N_4581,N_4690);
or U5090 (N_5090,N_4519,N_4517);
nand U5091 (N_5091,N_4763,N_4675);
xor U5092 (N_5092,N_4334,N_4418);
or U5093 (N_5093,N_4109,N_4526);
nor U5094 (N_5094,N_4633,N_4148);
nand U5095 (N_5095,N_4281,N_4969);
and U5096 (N_5096,N_4431,N_4383);
nor U5097 (N_5097,N_4196,N_4417);
or U5098 (N_5098,N_4053,N_4642);
or U5099 (N_5099,N_4303,N_4032);
nor U5100 (N_5100,N_4424,N_4728);
and U5101 (N_5101,N_4201,N_4742);
or U5102 (N_5102,N_4134,N_4340);
and U5103 (N_5103,N_4815,N_4532);
nor U5104 (N_5104,N_4776,N_4673);
nor U5105 (N_5105,N_4539,N_4385);
nand U5106 (N_5106,N_4174,N_4471);
nand U5107 (N_5107,N_4736,N_4326);
nand U5108 (N_5108,N_4738,N_4252);
and U5109 (N_5109,N_4176,N_4585);
nor U5110 (N_5110,N_4040,N_4250);
nor U5111 (N_5111,N_4546,N_4689);
nand U5112 (N_5112,N_4849,N_4254);
and U5113 (N_5113,N_4291,N_4714);
or U5114 (N_5114,N_4608,N_4975);
nand U5115 (N_5115,N_4048,N_4790);
nor U5116 (N_5116,N_4778,N_4564);
and U5117 (N_5117,N_4428,N_4895);
nand U5118 (N_5118,N_4786,N_4647);
nand U5119 (N_5119,N_4744,N_4407);
nor U5120 (N_5120,N_4027,N_4268);
and U5121 (N_5121,N_4771,N_4413);
nor U5122 (N_5122,N_4510,N_4670);
nand U5123 (N_5123,N_4365,N_4658);
and U5124 (N_5124,N_4563,N_4598);
and U5125 (N_5125,N_4884,N_4886);
or U5126 (N_5126,N_4362,N_4865);
or U5127 (N_5127,N_4933,N_4317);
and U5128 (N_5128,N_4829,N_4587);
nor U5129 (N_5129,N_4509,N_4812);
or U5130 (N_5130,N_4601,N_4062);
or U5131 (N_5131,N_4438,N_4400);
and U5132 (N_5132,N_4044,N_4984);
or U5133 (N_5133,N_4871,N_4534);
nor U5134 (N_5134,N_4737,N_4445);
or U5135 (N_5135,N_4309,N_4687);
nand U5136 (N_5136,N_4147,N_4152);
nor U5137 (N_5137,N_4562,N_4030);
nor U5138 (N_5138,N_4924,N_4756);
nor U5139 (N_5139,N_4366,N_4589);
nor U5140 (N_5140,N_4553,N_4549);
nor U5141 (N_5141,N_4926,N_4821);
nand U5142 (N_5142,N_4186,N_4054);
nor U5143 (N_5143,N_4677,N_4726);
or U5144 (N_5144,N_4348,N_4422);
nor U5145 (N_5145,N_4452,N_4169);
nor U5146 (N_5146,N_4506,N_4336);
nor U5147 (N_5147,N_4231,N_4396);
nand U5148 (N_5148,N_4140,N_4747);
nand U5149 (N_5149,N_4212,N_4935);
nor U5150 (N_5150,N_4312,N_4025);
or U5151 (N_5151,N_4957,N_4868);
and U5152 (N_5152,N_4936,N_4375);
nand U5153 (N_5153,N_4143,N_4599);
and U5154 (N_5154,N_4949,N_4079);
and U5155 (N_5155,N_4129,N_4567);
and U5156 (N_5156,N_4345,N_4325);
or U5157 (N_5157,N_4645,N_4316);
and U5158 (N_5158,N_4021,N_4270);
and U5159 (N_5159,N_4944,N_4235);
nand U5160 (N_5160,N_4099,N_4557);
or U5161 (N_5161,N_4609,N_4175);
and U5162 (N_5162,N_4006,N_4338);
nor U5163 (N_5163,N_4288,N_4086);
nand U5164 (N_5164,N_4315,N_4753);
nand U5165 (N_5165,N_4835,N_4018);
and U5166 (N_5166,N_4594,N_4818);
and U5167 (N_5167,N_4794,N_4374);
nor U5168 (N_5168,N_4339,N_4722);
nand U5169 (N_5169,N_4988,N_4993);
and U5170 (N_5170,N_4998,N_4560);
or U5171 (N_5171,N_4251,N_4968);
nand U5172 (N_5172,N_4770,N_4197);
and U5173 (N_5173,N_4110,N_4093);
and U5174 (N_5174,N_4097,N_4441);
or U5175 (N_5175,N_4188,N_4041);
nand U5176 (N_5176,N_4961,N_4962);
or U5177 (N_5177,N_4026,N_4912);
and U5178 (N_5178,N_4830,N_4127);
nor U5179 (N_5179,N_4624,N_4774);
nand U5180 (N_5180,N_4444,N_4700);
and U5181 (N_5181,N_4056,N_4462);
or U5182 (N_5182,N_4071,N_4964);
or U5183 (N_5183,N_4405,N_4284);
or U5184 (N_5184,N_4055,N_4671);
nor U5185 (N_5185,N_4531,N_4063);
nor U5186 (N_5186,N_4792,N_4588);
xnor U5187 (N_5187,N_4904,N_4241);
nand U5188 (N_5188,N_4733,N_4177);
or U5189 (N_5189,N_4986,N_4100);
or U5190 (N_5190,N_4159,N_4059);
nand U5191 (N_5191,N_4038,N_4853);
nor U5192 (N_5192,N_4359,N_4989);
nor U5193 (N_5193,N_4262,N_4832);
or U5194 (N_5194,N_4344,N_4384);
or U5195 (N_5195,N_4209,N_4017);
or U5196 (N_5196,N_4507,N_4213);
or U5197 (N_5197,N_4551,N_4946);
nor U5198 (N_5198,N_4899,N_4245);
and U5199 (N_5199,N_4856,N_4873);
or U5200 (N_5200,N_4394,N_4141);
nor U5201 (N_5201,N_4081,N_4573);
nor U5202 (N_5202,N_4191,N_4411);
and U5203 (N_5203,N_4267,N_4535);
or U5204 (N_5204,N_4780,N_4189);
and U5205 (N_5205,N_4139,N_4458);
and U5206 (N_5206,N_4999,N_4639);
or U5207 (N_5207,N_4341,N_4157);
or U5208 (N_5208,N_4908,N_4492);
or U5209 (N_5209,N_4179,N_4132);
or U5210 (N_5210,N_4078,N_4228);
xor U5211 (N_5211,N_4541,N_4806);
or U5212 (N_5212,N_4160,N_4389);
or U5213 (N_5213,N_4801,N_4111);
nor U5214 (N_5214,N_4090,N_4704);
nor U5215 (N_5215,N_4523,N_4049);
and U5216 (N_5216,N_4967,N_4124);
nor U5217 (N_5217,N_4977,N_4888);
and U5218 (N_5218,N_4355,N_4512);
and U5219 (N_5219,N_4813,N_4119);
and U5220 (N_5220,N_4330,N_4703);
nand U5221 (N_5221,N_4106,N_4550);
nand U5222 (N_5222,N_4295,N_4808);
nor U5223 (N_5223,N_4346,N_4352);
or U5224 (N_5224,N_4901,N_4630);
or U5225 (N_5225,N_4230,N_4455);
or U5226 (N_5226,N_4015,N_4453);
or U5227 (N_5227,N_4826,N_4943);
and U5228 (N_5228,N_4075,N_4574);
nor U5229 (N_5229,N_4604,N_4425);
and U5230 (N_5230,N_4822,N_4513);
and U5231 (N_5231,N_4484,N_4150);
nor U5232 (N_5232,N_4020,N_4758);
nand U5233 (N_5233,N_4360,N_4953);
nand U5234 (N_5234,N_4734,N_4283);
nor U5235 (N_5235,N_4825,N_4376);
xor U5236 (N_5236,N_4745,N_4997);
or U5237 (N_5237,N_4036,N_4823);
nor U5238 (N_5238,N_4433,N_4391);
nor U5239 (N_5239,N_4153,N_4005);
or U5240 (N_5240,N_4906,N_4060);
nand U5241 (N_5241,N_4709,N_4135);
and U5242 (N_5242,N_4854,N_4769);
and U5243 (N_5243,N_4928,N_4617);
or U5244 (N_5244,N_4979,N_4779);
nand U5245 (N_5245,N_4485,N_4536);
or U5246 (N_5246,N_4217,N_4183);
nand U5247 (N_5247,N_4636,N_4874);
or U5248 (N_5248,N_4556,N_4261);
nor U5249 (N_5249,N_4314,N_4592);
and U5250 (N_5250,N_4224,N_4193);
or U5251 (N_5251,N_4207,N_4730);
nand U5252 (N_5252,N_4586,N_4836);
nor U5253 (N_5253,N_4894,N_4809);
nor U5254 (N_5254,N_4666,N_4443);
xnor U5255 (N_5255,N_4613,N_4001);
nor U5256 (N_5256,N_4927,N_4364);
and U5257 (N_5257,N_4723,N_4372);
nor U5258 (N_5258,N_4782,N_4448);
nor U5259 (N_5259,N_4225,N_4974);
or U5260 (N_5260,N_4789,N_4220);
and U5261 (N_5261,N_4337,N_4263);
nor U5262 (N_5262,N_4983,N_4168);
nand U5263 (N_5263,N_4956,N_4223);
and U5264 (N_5264,N_4470,N_4137);
nor U5265 (N_5265,N_4487,N_4649);
or U5266 (N_5266,N_4170,N_4070);
and U5267 (N_5267,N_4521,N_4803);
or U5268 (N_5268,N_4852,N_4475);
nor U5269 (N_5269,N_4824,N_4037);
nor U5270 (N_5270,N_4237,N_4839);
or U5271 (N_5271,N_4820,N_4612);
nor U5272 (N_5272,N_4440,N_4527);
nor U5273 (N_5273,N_4570,N_4064);
xor U5274 (N_5274,N_4138,N_4112);
or U5275 (N_5275,N_4491,N_4572);
and U5276 (N_5276,N_4693,N_4537);
or U5277 (N_5277,N_4073,N_4941);
nor U5278 (N_5278,N_4861,N_4802);
nor U5279 (N_5279,N_4615,N_4766);
nor U5280 (N_5280,N_4691,N_4610);
or U5281 (N_5281,N_4102,N_4859);
nor U5282 (N_5282,N_4292,N_4204);
nand U5283 (N_5283,N_4232,N_4889);
or U5284 (N_5284,N_4469,N_4354);
nor U5285 (N_5285,N_4554,N_4960);
nand U5286 (N_5286,N_4472,N_4402);
and U5287 (N_5287,N_4864,N_4542);
nor U5288 (N_5288,N_4931,N_4247);
nor U5289 (N_5289,N_4486,N_4022);
nor U5290 (N_5290,N_4660,N_4990);
and U5291 (N_5291,N_4386,N_4000);
and U5292 (N_5292,N_4436,N_4710);
or U5293 (N_5293,N_4435,N_4952);
and U5294 (N_5294,N_4877,N_4190);
nor U5295 (N_5295,N_4855,N_4893);
nor U5296 (N_5296,N_4367,N_4558);
or U5297 (N_5297,N_4662,N_4187);
nand U5298 (N_5298,N_4439,N_4891);
and U5299 (N_5299,N_4914,N_4208);
nand U5300 (N_5300,N_4844,N_4088);
or U5301 (N_5301,N_4712,N_4929);
nor U5302 (N_5302,N_4760,N_4765);
nor U5303 (N_5303,N_4136,N_4545);
nor U5304 (N_5304,N_4793,N_4399);
nor U5305 (N_5305,N_4575,N_4629);
or U5306 (N_5306,N_4991,N_4858);
and U5307 (N_5307,N_4265,N_4126);
nand U5308 (N_5308,N_4285,N_4456);
nand U5309 (N_5309,N_4483,N_4890);
nor U5310 (N_5310,N_4181,N_4311);
and U5311 (N_5311,N_4406,N_4258);
nor U5312 (N_5312,N_4350,N_4370);
or U5313 (N_5313,N_4796,N_4296);
nor U5314 (N_5314,N_4667,N_4881);
and U5315 (N_5315,N_4294,N_4706);
and U5316 (N_5316,N_4764,N_4467);
nand U5317 (N_5317,N_4369,N_4994);
and U5318 (N_5318,N_4167,N_4727);
nor U5319 (N_5319,N_4198,N_4862);
or U5320 (N_5320,N_4194,N_4404);
and U5321 (N_5321,N_4379,N_4161);
and U5322 (N_5322,N_4328,N_4937);
nor U5323 (N_5323,N_4632,N_4876);
nand U5324 (N_5324,N_4272,N_4795);
and U5325 (N_5325,N_4672,N_4655);
nor U5326 (N_5326,N_4357,N_4905);
nand U5327 (N_5327,N_4342,N_4683);
nor U5328 (N_5328,N_4547,N_4860);
nor U5329 (N_5329,N_4503,N_4816);
nand U5330 (N_5330,N_4595,N_4416);
and U5331 (N_5331,N_4711,N_4932);
nand U5332 (N_5332,N_4735,N_4218);
nand U5333 (N_5333,N_4437,N_4942);
or U5334 (N_5334,N_4398,N_4450);
and U5335 (N_5335,N_4963,N_4811);
nor U5336 (N_5336,N_4749,N_4800);
nand U5337 (N_5337,N_4681,N_4358);
or U5338 (N_5338,N_4066,N_4244);
nand U5339 (N_5339,N_4403,N_4804);
nor U5340 (N_5340,N_4427,N_4708);
or U5341 (N_5341,N_4732,N_4498);
and U5342 (N_5342,N_4474,N_4434);
nand U5343 (N_5343,N_4828,N_4644);
nor U5344 (N_5344,N_4731,N_4226);
or U5345 (N_5345,N_4104,N_4916);
or U5346 (N_5346,N_4361,N_4171);
nor U5347 (N_5347,N_4656,N_4052);
nor U5348 (N_5348,N_4785,N_4087);
nor U5349 (N_5349,N_4277,N_4892);
nor U5350 (N_5350,N_4117,N_4500);
xnor U5351 (N_5351,N_4105,N_4948);
and U5352 (N_5352,N_4145,N_4694);
or U5353 (N_5353,N_4698,N_4113);
nor U5354 (N_5354,N_4280,N_4680);
and U5355 (N_5355,N_4900,N_4343);
nor U5356 (N_5356,N_4151,N_4590);
nor U5357 (N_5357,N_4982,N_4863);
nor U5358 (N_5358,N_4033,N_4082);
nand U5359 (N_5359,N_4569,N_4872);
and U5360 (N_5360,N_4757,N_4101);
nand U5361 (N_5361,N_4614,N_4114);
or U5362 (N_5362,N_4465,N_4819);
and U5363 (N_5363,N_4724,N_4922);
and U5364 (N_5364,N_4807,N_4831);
xnor U5365 (N_5365,N_4954,N_4306);
nor U5366 (N_5366,N_4602,N_4559);
nor U5367 (N_5367,N_4410,N_4619);
nor U5368 (N_5368,N_4761,N_4980);
and U5369 (N_5369,N_4323,N_4497);
and U5370 (N_5370,N_4184,N_4091);
nor U5371 (N_5371,N_4144,N_4684);
and U5372 (N_5372,N_4845,N_4023);
nand U5373 (N_5373,N_4966,N_4725);
nand U5374 (N_5374,N_4378,N_4842);
nor U5375 (N_5375,N_4869,N_4686);
nand U5376 (N_5376,N_4654,N_4016);
nand U5377 (N_5377,N_4814,N_4046);
nor U5378 (N_5378,N_4955,N_4850);
nand U5379 (N_5379,N_4939,N_4783);
nand U5380 (N_5380,N_4240,N_4985);
or U5381 (N_5381,N_4414,N_4211);
or U5382 (N_5382,N_4122,N_4318);
nand U5383 (N_5383,N_4130,N_4451);
and U5384 (N_5384,N_4058,N_4489);
nor U5385 (N_5385,N_4002,N_4256);
nand U5386 (N_5386,N_4089,N_4166);
nand U5387 (N_5387,N_4039,N_4286);
or U5388 (N_5388,N_4298,N_4185);
and U5389 (N_5389,N_4473,N_4297);
nand U5390 (N_5390,N_4481,N_4200);
or U5391 (N_5391,N_4125,N_4679);
or U5392 (N_5392,N_4799,N_4287);
nor U5393 (N_5393,N_4118,N_4695);
or U5394 (N_5394,N_4008,N_4552);
or U5395 (N_5395,N_4668,N_4401);
nor U5396 (N_5396,N_4307,N_4607);
or U5397 (N_5397,N_4784,N_4646);
or U5398 (N_5398,N_4074,N_4221);
or U5399 (N_5399,N_4203,N_4525);
nand U5400 (N_5400,N_4634,N_4460);
and U5401 (N_5401,N_4664,N_4482);
and U5402 (N_5402,N_4887,N_4381);
and U5403 (N_5403,N_4911,N_4641);
or U5404 (N_5404,N_4092,N_4123);
and U5405 (N_5405,N_4637,N_4685);
nor U5406 (N_5406,N_4973,N_4781);
or U5407 (N_5407,N_4249,N_4271);
nor U5408 (N_5408,N_4042,N_4880);
nand U5409 (N_5409,N_4739,N_4768);
or U5410 (N_5410,N_4743,N_4840);
nand U5411 (N_5411,N_4987,N_4578);
nor U5412 (N_5412,N_4229,N_4072);
and U5413 (N_5413,N_4959,N_4848);
nand U5414 (N_5414,N_4885,N_4528);
nor U5415 (N_5415,N_4259,N_4461);
and U5416 (N_5416,N_4676,N_4643);
or U5417 (N_5417,N_4479,N_4674);
or U5418 (N_5418,N_4010,N_4907);
and U5419 (N_5419,N_4393,N_4390);
nand U5420 (N_5420,N_4493,N_4260);
nor U5421 (N_5421,N_4164,N_4950);
nor U5422 (N_5422,N_4879,N_4085);
nand U5423 (N_5423,N_4622,N_4029);
and U5424 (N_5424,N_4233,N_4773);
or U5425 (N_5425,N_4833,N_4289);
nand U5426 (N_5426,N_4661,N_4925);
nand U5427 (N_5427,N_4146,N_4083);
or U5428 (N_5428,N_4299,N_4741);
nand U5429 (N_5429,N_4958,N_4866);
nor U5430 (N_5430,N_4423,N_4568);
or U5431 (N_5431,N_4591,N_4495);
nand U5432 (N_5432,N_4548,N_4707);
or U5433 (N_5433,N_4976,N_4173);
nand U5434 (N_5434,N_4896,N_4965);
and U5435 (N_5435,N_4057,N_4847);
nand U5436 (N_5436,N_4447,N_4940);
nand U5437 (N_5437,N_4457,N_4408);
nand U5438 (N_5438,N_4752,N_4108);
nand U5439 (N_5439,N_4180,N_4597);
nor U5440 (N_5440,N_4215,N_4970);
and U5441 (N_5441,N_4158,N_4420);
nor U5442 (N_5442,N_4347,N_4718);
nand U5443 (N_5443,N_4419,N_4788);
nand U5444 (N_5444,N_4701,N_4627);
or U5445 (N_5445,N_4529,N_4236);
nand U5446 (N_5446,N_4293,N_4321);
or U5447 (N_5447,N_4463,N_4333);
or U5448 (N_5448,N_4163,N_4945);
and U5449 (N_5449,N_4628,N_4938);
and U5450 (N_5450,N_4571,N_4214);
nand U5451 (N_5451,N_4007,N_4555);
and U5452 (N_5452,N_4305,N_4363);
or U5453 (N_5453,N_4449,N_4897);
nor U5454 (N_5454,N_4867,N_4631);
or U5455 (N_5455,N_4648,N_4238);
nor U5456 (N_5456,N_4466,N_4392);
nand U5457 (N_5457,N_4084,N_4248);
and U5458 (N_5458,N_4524,N_4274);
nor U5459 (N_5459,N_4182,N_4257);
and U5460 (N_5460,N_4883,N_4605);
or U5461 (N_5461,N_4195,N_4625);
and U5462 (N_5462,N_4713,N_4353);
nor U5463 (N_5463,N_4290,N_4682);
nand U5464 (N_5464,N_4210,N_4843);
and U5465 (N_5465,N_4544,N_4717);
and U5466 (N_5466,N_4611,N_4919);
nand U5467 (N_5467,N_4349,N_4846);
xor U5468 (N_5468,N_4121,N_4898);
nor U5469 (N_5469,N_4651,N_4371);
nor U5470 (N_5470,N_4951,N_4013);
nor U5471 (N_5471,N_4650,N_4319);
nor U5472 (N_5472,N_4582,N_4913);
or U5473 (N_5473,N_4276,N_4678);
or U5474 (N_5474,N_4388,N_4522);
and U5475 (N_5475,N_4094,N_4488);
and U5476 (N_5476,N_4310,N_4635);
and U5477 (N_5477,N_4699,N_4476);
nor U5478 (N_5478,N_4446,N_4468);
or U5479 (N_5479,N_4909,N_4031);
nor U5480 (N_5480,N_4454,N_4076);
nor U5481 (N_5481,N_4442,N_4335);
nand U5482 (N_5482,N_4787,N_4875);
nand U5483 (N_5483,N_4373,N_4659);
nand U5484 (N_5484,N_4702,N_4841);
or U5485 (N_5485,N_4827,N_4810);
nand U5486 (N_5486,N_4216,N_4227);
and U5487 (N_5487,N_4638,N_4412);
and U5488 (N_5488,N_4514,N_4133);
and U5489 (N_5489,N_4278,N_4719);
nor U5490 (N_5490,N_4903,N_4024);
nor U5491 (N_5491,N_4478,N_4669);
and U5492 (N_5492,N_4518,N_4098);
and U5493 (N_5493,N_4327,N_4034);
and U5494 (N_5494,N_4045,N_4172);
nand U5495 (N_5495,N_4069,N_4302);
or U5496 (N_5496,N_4011,N_4494);
or U5497 (N_5497,N_4971,N_4620);
or U5498 (N_5498,N_4775,N_4540);
or U5499 (N_5499,N_4351,N_4499);
or U5500 (N_5500,N_4081,N_4001);
nand U5501 (N_5501,N_4660,N_4750);
nor U5502 (N_5502,N_4979,N_4711);
or U5503 (N_5503,N_4899,N_4019);
or U5504 (N_5504,N_4397,N_4903);
xor U5505 (N_5505,N_4522,N_4230);
and U5506 (N_5506,N_4285,N_4806);
nand U5507 (N_5507,N_4298,N_4944);
nand U5508 (N_5508,N_4120,N_4615);
or U5509 (N_5509,N_4754,N_4025);
nand U5510 (N_5510,N_4801,N_4732);
nand U5511 (N_5511,N_4891,N_4026);
nor U5512 (N_5512,N_4322,N_4617);
or U5513 (N_5513,N_4006,N_4516);
nand U5514 (N_5514,N_4400,N_4258);
nand U5515 (N_5515,N_4684,N_4324);
or U5516 (N_5516,N_4112,N_4300);
nand U5517 (N_5517,N_4056,N_4741);
and U5518 (N_5518,N_4322,N_4160);
nor U5519 (N_5519,N_4296,N_4324);
or U5520 (N_5520,N_4514,N_4989);
nor U5521 (N_5521,N_4341,N_4025);
nor U5522 (N_5522,N_4535,N_4103);
nor U5523 (N_5523,N_4900,N_4804);
nor U5524 (N_5524,N_4935,N_4556);
nand U5525 (N_5525,N_4173,N_4747);
nor U5526 (N_5526,N_4243,N_4540);
and U5527 (N_5527,N_4171,N_4581);
nor U5528 (N_5528,N_4636,N_4016);
nor U5529 (N_5529,N_4723,N_4678);
nor U5530 (N_5530,N_4039,N_4396);
or U5531 (N_5531,N_4257,N_4844);
nor U5532 (N_5532,N_4988,N_4095);
and U5533 (N_5533,N_4383,N_4496);
nand U5534 (N_5534,N_4009,N_4595);
or U5535 (N_5535,N_4028,N_4182);
nor U5536 (N_5536,N_4580,N_4499);
nand U5537 (N_5537,N_4114,N_4795);
nand U5538 (N_5538,N_4312,N_4830);
nor U5539 (N_5539,N_4308,N_4859);
or U5540 (N_5540,N_4608,N_4285);
or U5541 (N_5541,N_4099,N_4152);
and U5542 (N_5542,N_4171,N_4042);
or U5543 (N_5543,N_4401,N_4435);
nor U5544 (N_5544,N_4479,N_4553);
nand U5545 (N_5545,N_4344,N_4301);
nand U5546 (N_5546,N_4153,N_4823);
and U5547 (N_5547,N_4743,N_4348);
nor U5548 (N_5548,N_4102,N_4401);
nor U5549 (N_5549,N_4314,N_4986);
or U5550 (N_5550,N_4439,N_4343);
nor U5551 (N_5551,N_4220,N_4659);
or U5552 (N_5552,N_4160,N_4518);
and U5553 (N_5553,N_4784,N_4676);
nor U5554 (N_5554,N_4562,N_4005);
nand U5555 (N_5555,N_4332,N_4050);
and U5556 (N_5556,N_4869,N_4714);
or U5557 (N_5557,N_4571,N_4058);
nand U5558 (N_5558,N_4417,N_4082);
nand U5559 (N_5559,N_4656,N_4891);
nand U5560 (N_5560,N_4043,N_4452);
nand U5561 (N_5561,N_4894,N_4797);
or U5562 (N_5562,N_4092,N_4916);
and U5563 (N_5563,N_4387,N_4172);
and U5564 (N_5564,N_4660,N_4039);
nand U5565 (N_5565,N_4584,N_4844);
nand U5566 (N_5566,N_4083,N_4371);
or U5567 (N_5567,N_4268,N_4141);
and U5568 (N_5568,N_4553,N_4657);
and U5569 (N_5569,N_4709,N_4371);
nand U5570 (N_5570,N_4479,N_4526);
or U5571 (N_5571,N_4452,N_4743);
nand U5572 (N_5572,N_4535,N_4023);
nand U5573 (N_5573,N_4494,N_4132);
and U5574 (N_5574,N_4162,N_4227);
nand U5575 (N_5575,N_4839,N_4342);
and U5576 (N_5576,N_4717,N_4377);
nor U5577 (N_5577,N_4741,N_4256);
and U5578 (N_5578,N_4971,N_4133);
and U5579 (N_5579,N_4954,N_4704);
or U5580 (N_5580,N_4451,N_4994);
nor U5581 (N_5581,N_4690,N_4437);
nand U5582 (N_5582,N_4060,N_4560);
nor U5583 (N_5583,N_4591,N_4579);
and U5584 (N_5584,N_4497,N_4707);
nand U5585 (N_5585,N_4394,N_4179);
or U5586 (N_5586,N_4337,N_4787);
nand U5587 (N_5587,N_4086,N_4543);
or U5588 (N_5588,N_4840,N_4755);
and U5589 (N_5589,N_4220,N_4108);
or U5590 (N_5590,N_4832,N_4462);
nand U5591 (N_5591,N_4913,N_4260);
nor U5592 (N_5592,N_4978,N_4378);
nor U5593 (N_5593,N_4755,N_4046);
nand U5594 (N_5594,N_4735,N_4837);
nor U5595 (N_5595,N_4272,N_4081);
or U5596 (N_5596,N_4425,N_4965);
or U5597 (N_5597,N_4553,N_4389);
nor U5598 (N_5598,N_4447,N_4266);
nor U5599 (N_5599,N_4348,N_4239);
nor U5600 (N_5600,N_4408,N_4663);
or U5601 (N_5601,N_4167,N_4511);
or U5602 (N_5602,N_4319,N_4522);
and U5603 (N_5603,N_4013,N_4142);
and U5604 (N_5604,N_4925,N_4519);
nor U5605 (N_5605,N_4688,N_4999);
nor U5606 (N_5606,N_4343,N_4052);
or U5607 (N_5607,N_4563,N_4185);
nor U5608 (N_5608,N_4357,N_4234);
or U5609 (N_5609,N_4264,N_4231);
or U5610 (N_5610,N_4535,N_4599);
nor U5611 (N_5611,N_4542,N_4517);
and U5612 (N_5612,N_4552,N_4608);
nand U5613 (N_5613,N_4452,N_4561);
and U5614 (N_5614,N_4580,N_4628);
nor U5615 (N_5615,N_4746,N_4930);
and U5616 (N_5616,N_4423,N_4761);
nand U5617 (N_5617,N_4219,N_4621);
or U5618 (N_5618,N_4535,N_4922);
and U5619 (N_5619,N_4991,N_4891);
nor U5620 (N_5620,N_4404,N_4159);
nand U5621 (N_5621,N_4817,N_4845);
or U5622 (N_5622,N_4206,N_4163);
nor U5623 (N_5623,N_4035,N_4172);
nor U5624 (N_5624,N_4749,N_4121);
and U5625 (N_5625,N_4369,N_4862);
xor U5626 (N_5626,N_4374,N_4540);
nor U5627 (N_5627,N_4963,N_4677);
nand U5628 (N_5628,N_4588,N_4493);
nand U5629 (N_5629,N_4552,N_4378);
and U5630 (N_5630,N_4637,N_4772);
or U5631 (N_5631,N_4294,N_4529);
nand U5632 (N_5632,N_4182,N_4953);
nor U5633 (N_5633,N_4603,N_4989);
nand U5634 (N_5634,N_4433,N_4904);
and U5635 (N_5635,N_4997,N_4284);
nor U5636 (N_5636,N_4208,N_4076);
xnor U5637 (N_5637,N_4685,N_4251);
and U5638 (N_5638,N_4354,N_4822);
and U5639 (N_5639,N_4858,N_4063);
xor U5640 (N_5640,N_4719,N_4241);
and U5641 (N_5641,N_4702,N_4544);
nor U5642 (N_5642,N_4401,N_4611);
or U5643 (N_5643,N_4396,N_4025);
nand U5644 (N_5644,N_4408,N_4230);
nor U5645 (N_5645,N_4653,N_4801);
nand U5646 (N_5646,N_4306,N_4378);
nand U5647 (N_5647,N_4055,N_4079);
or U5648 (N_5648,N_4263,N_4398);
nor U5649 (N_5649,N_4303,N_4377);
nand U5650 (N_5650,N_4413,N_4238);
and U5651 (N_5651,N_4882,N_4417);
and U5652 (N_5652,N_4272,N_4873);
and U5653 (N_5653,N_4051,N_4971);
nand U5654 (N_5654,N_4595,N_4056);
nand U5655 (N_5655,N_4214,N_4760);
nand U5656 (N_5656,N_4308,N_4900);
and U5657 (N_5657,N_4704,N_4949);
nor U5658 (N_5658,N_4718,N_4762);
nand U5659 (N_5659,N_4757,N_4788);
nor U5660 (N_5660,N_4732,N_4682);
nor U5661 (N_5661,N_4321,N_4945);
nand U5662 (N_5662,N_4973,N_4160);
and U5663 (N_5663,N_4331,N_4321);
or U5664 (N_5664,N_4096,N_4049);
nand U5665 (N_5665,N_4422,N_4622);
nor U5666 (N_5666,N_4208,N_4199);
and U5667 (N_5667,N_4150,N_4553);
nor U5668 (N_5668,N_4565,N_4846);
or U5669 (N_5669,N_4255,N_4093);
and U5670 (N_5670,N_4832,N_4337);
nand U5671 (N_5671,N_4098,N_4686);
nand U5672 (N_5672,N_4602,N_4206);
or U5673 (N_5673,N_4499,N_4230);
nand U5674 (N_5674,N_4085,N_4707);
nor U5675 (N_5675,N_4105,N_4724);
nand U5676 (N_5676,N_4171,N_4391);
nand U5677 (N_5677,N_4486,N_4230);
nor U5678 (N_5678,N_4161,N_4867);
and U5679 (N_5679,N_4471,N_4630);
nand U5680 (N_5680,N_4506,N_4769);
and U5681 (N_5681,N_4439,N_4841);
and U5682 (N_5682,N_4934,N_4564);
nor U5683 (N_5683,N_4112,N_4554);
and U5684 (N_5684,N_4369,N_4330);
or U5685 (N_5685,N_4042,N_4568);
nand U5686 (N_5686,N_4411,N_4512);
nand U5687 (N_5687,N_4323,N_4365);
or U5688 (N_5688,N_4218,N_4038);
and U5689 (N_5689,N_4347,N_4788);
nand U5690 (N_5690,N_4125,N_4309);
and U5691 (N_5691,N_4537,N_4327);
nand U5692 (N_5692,N_4104,N_4124);
and U5693 (N_5693,N_4266,N_4470);
nand U5694 (N_5694,N_4797,N_4662);
nor U5695 (N_5695,N_4054,N_4244);
nand U5696 (N_5696,N_4243,N_4309);
nor U5697 (N_5697,N_4080,N_4861);
xnor U5698 (N_5698,N_4100,N_4757);
nor U5699 (N_5699,N_4639,N_4252);
nor U5700 (N_5700,N_4827,N_4975);
or U5701 (N_5701,N_4566,N_4199);
nor U5702 (N_5702,N_4792,N_4414);
and U5703 (N_5703,N_4094,N_4011);
or U5704 (N_5704,N_4464,N_4223);
nand U5705 (N_5705,N_4469,N_4956);
nand U5706 (N_5706,N_4775,N_4776);
nor U5707 (N_5707,N_4507,N_4227);
nand U5708 (N_5708,N_4615,N_4419);
and U5709 (N_5709,N_4017,N_4099);
nor U5710 (N_5710,N_4749,N_4402);
and U5711 (N_5711,N_4239,N_4440);
nand U5712 (N_5712,N_4982,N_4348);
nor U5713 (N_5713,N_4073,N_4881);
and U5714 (N_5714,N_4086,N_4047);
or U5715 (N_5715,N_4789,N_4741);
and U5716 (N_5716,N_4912,N_4581);
and U5717 (N_5717,N_4126,N_4155);
nor U5718 (N_5718,N_4234,N_4865);
nor U5719 (N_5719,N_4868,N_4512);
and U5720 (N_5720,N_4842,N_4927);
nor U5721 (N_5721,N_4783,N_4104);
or U5722 (N_5722,N_4554,N_4005);
or U5723 (N_5723,N_4071,N_4998);
or U5724 (N_5724,N_4161,N_4896);
nand U5725 (N_5725,N_4944,N_4970);
and U5726 (N_5726,N_4876,N_4367);
nand U5727 (N_5727,N_4840,N_4335);
nor U5728 (N_5728,N_4170,N_4772);
nor U5729 (N_5729,N_4346,N_4109);
and U5730 (N_5730,N_4822,N_4463);
or U5731 (N_5731,N_4733,N_4604);
and U5732 (N_5732,N_4495,N_4614);
nor U5733 (N_5733,N_4572,N_4060);
nand U5734 (N_5734,N_4000,N_4958);
nand U5735 (N_5735,N_4422,N_4584);
nand U5736 (N_5736,N_4841,N_4040);
nor U5737 (N_5737,N_4533,N_4563);
nand U5738 (N_5738,N_4178,N_4397);
nand U5739 (N_5739,N_4741,N_4681);
and U5740 (N_5740,N_4128,N_4140);
and U5741 (N_5741,N_4137,N_4861);
nor U5742 (N_5742,N_4123,N_4634);
nand U5743 (N_5743,N_4364,N_4244);
and U5744 (N_5744,N_4556,N_4237);
nor U5745 (N_5745,N_4662,N_4002);
and U5746 (N_5746,N_4453,N_4894);
or U5747 (N_5747,N_4518,N_4245);
or U5748 (N_5748,N_4544,N_4258);
and U5749 (N_5749,N_4601,N_4806);
or U5750 (N_5750,N_4846,N_4871);
nor U5751 (N_5751,N_4818,N_4007);
nor U5752 (N_5752,N_4226,N_4551);
nand U5753 (N_5753,N_4222,N_4893);
nand U5754 (N_5754,N_4572,N_4584);
nand U5755 (N_5755,N_4053,N_4443);
and U5756 (N_5756,N_4461,N_4984);
nor U5757 (N_5757,N_4407,N_4212);
and U5758 (N_5758,N_4407,N_4602);
nor U5759 (N_5759,N_4015,N_4470);
nand U5760 (N_5760,N_4394,N_4266);
or U5761 (N_5761,N_4836,N_4538);
and U5762 (N_5762,N_4406,N_4886);
and U5763 (N_5763,N_4547,N_4192);
and U5764 (N_5764,N_4678,N_4535);
nor U5765 (N_5765,N_4741,N_4180);
nor U5766 (N_5766,N_4022,N_4412);
nor U5767 (N_5767,N_4843,N_4560);
nand U5768 (N_5768,N_4383,N_4103);
and U5769 (N_5769,N_4022,N_4303);
xnor U5770 (N_5770,N_4217,N_4796);
nor U5771 (N_5771,N_4667,N_4500);
nand U5772 (N_5772,N_4380,N_4811);
nand U5773 (N_5773,N_4365,N_4289);
nand U5774 (N_5774,N_4792,N_4784);
or U5775 (N_5775,N_4218,N_4679);
or U5776 (N_5776,N_4364,N_4687);
and U5777 (N_5777,N_4959,N_4902);
or U5778 (N_5778,N_4578,N_4189);
nor U5779 (N_5779,N_4485,N_4101);
or U5780 (N_5780,N_4471,N_4566);
and U5781 (N_5781,N_4603,N_4386);
and U5782 (N_5782,N_4317,N_4235);
or U5783 (N_5783,N_4609,N_4907);
nor U5784 (N_5784,N_4251,N_4440);
nand U5785 (N_5785,N_4405,N_4182);
or U5786 (N_5786,N_4761,N_4445);
and U5787 (N_5787,N_4632,N_4118);
nand U5788 (N_5788,N_4658,N_4319);
nor U5789 (N_5789,N_4449,N_4376);
or U5790 (N_5790,N_4014,N_4929);
or U5791 (N_5791,N_4468,N_4907);
or U5792 (N_5792,N_4568,N_4074);
nand U5793 (N_5793,N_4063,N_4244);
nand U5794 (N_5794,N_4706,N_4276);
nor U5795 (N_5795,N_4795,N_4615);
nor U5796 (N_5796,N_4617,N_4425);
and U5797 (N_5797,N_4155,N_4879);
and U5798 (N_5798,N_4303,N_4237);
and U5799 (N_5799,N_4018,N_4932);
nand U5800 (N_5800,N_4826,N_4828);
or U5801 (N_5801,N_4247,N_4102);
nor U5802 (N_5802,N_4269,N_4636);
nor U5803 (N_5803,N_4086,N_4108);
nand U5804 (N_5804,N_4992,N_4680);
nor U5805 (N_5805,N_4767,N_4410);
or U5806 (N_5806,N_4348,N_4543);
nor U5807 (N_5807,N_4913,N_4022);
nor U5808 (N_5808,N_4610,N_4976);
nand U5809 (N_5809,N_4139,N_4515);
nand U5810 (N_5810,N_4523,N_4839);
and U5811 (N_5811,N_4839,N_4427);
nand U5812 (N_5812,N_4939,N_4778);
nand U5813 (N_5813,N_4691,N_4385);
nor U5814 (N_5814,N_4999,N_4083);
and U5815 (N_5815,N_4170,N_4389);
or U5816 (N_5816,N_4188,N_4179);
nor U5817 (N_5817,N_4312,N_4475);
nor U5818 (N_5818,N_4013,N_4007);
nand U5819 (N_5819,N_4504,N_4950);
and U5820 (N_5820,N_4770,N_4676);
nor U5821 (N_5821,N_4524,N_4577);
nor U5822 (N_5822,N_4647,N_4365);
and U5823 (N_5823,N_4792,N_4745);
and U5824 (N_5824,N_4812,N_4258);
and U5825 (N_5825,N_4919,N_4696);
nor U5826 (N_5826,N_4204,N_4780);
or U5827 (N_5827,N_4491,N_4345);
or U5828 (N_5828,N_4346,N_4638);
nand U5829 (N_5829,N_4334,N_4294);
and U5830 (N_5830,N_4181,N_4863);
or U5831 (N_5831,N_4444,N_4477);
nand U5832 (N_5832,N_4844,N_4541);
nand U5833 (N_5833,N_4347,N_4207);
nor U5834 (N_5834,N_4989,N_4318);
or U5835 (N_5835,N_4168,N_4132);
nand U5836 (N_5836,N_4995,N_4552);
or U5837 (N_5837,N_4552,N_4433);
nor U5838 (N_5838,N_4541,N_4099);
nand U5839 (N_5839,N_4138,N_4739);
nor U5840 (N_5840,N_4339,N_4903);
and U5841 (N_5841,N_4334,N_4322);
and U5842 (N_5842,N_4493,N_4880);
and U5843 (N_5843,N_4243,N_4596);
and U5844 (N_5844,N_4225,N_4493);
and U5845 (N_5845,N_4732,N_4744);
and U5846 (N_5846,N_4048,N_4462);
nand U5847 (N_5847,N_4573,N_4986);
nand U5848 (N_5848,N_4543,N_4014);
nor U5849 (N_5849,N_4460,N_4454);
and U5850 (N_5850,N_4662,N_4506);
or U5851 (N_5851,N_4383,N_4180);
nor U5852 (N_5852,N_4612,N_4933);
nand U5853 (N_5853,N_4000,N_4293);
nand U5854 (N_5854,N_4293,N_4103);
nor U5855 (N_5855,N_4485,N_4880);
or U5856 (N_5856,N_4310,N_4116);
nand U5857 (N_5857,N_4656,N_4030);
nand U5858 (N_5858,N_4559,N_4296);
and U5859 (N_5859,N_4376,N_4014);
nand U5860 (N_5860,N_4895,N_4542);
or U5861 (N_5861,N_4183,N_4956);
nor U5862 (N_5862,N_4045,N_4657);
nor U5863 (N_5863,N_4805,N_4717);
or U5864 (N_5864,N_4588,N_4866);
and U5865 (N_5865,N_4365,N_4253);
and U5866 (N_5866,N_4025,N_4669);
nand U5867 (N_5867,N_4444,N_4183);
nand U5868 (N_5868,N_4621,N_4609);
and U5869 (N_5869,N_4147,N_4756);
and U5870 (N_5870,N_4139,N_4437);
nor U5871 (N_5871,N_4067,N_4242);
nand U5872 (N_5872,N_4816,N_4781);
nand U5873 (N_5873,N_4693,N_4179);
or U5874 (N_5874,N_4502,N_4129);
and U5875 (N_5875,N_4003,N_4239);
nor U5876 (N_5876,N_4411,N_4143);
or U5877 (N_5877,N_4683,N_4130);
nor U5878 (N_5878,N_4002,N_4424);
nor U5879 (N_5879,N_4591,N_4160);
or U5880 (N_5880,N_4249,N_4198);
nand U5881 (N_5881,N_4217,N_4437);
nand U5882 (N_5882,N_4096,N_4683);
nand U5883 (N_5883,N_4388,N_4403);
or U5884 (N_5884,N_4782,N_4655);
nand U5885 (N_5885,N_4202,N_4923);
or U5886 (N_5886,N_4987,N_4054);
or U5887 (N_5887,N_4867,N_4767);
and U5888 (N_5888,N_4431,N_4730);
nand U5889 (N_5889,N_4259,N_4562);
or U5890 (N_5890,N_4531,N_4003);
nand U5891 (N_5891,N_4014,N_4521);
nand U5892 (N_5892,N_4046,N_4888);
and U5893 (N_5893,N_4391,N_4550);
nor U5894 (N_5894,N_4062,N_4360);
or U5895 (N_5895,N_4470,N_4972);
nor U5896 (N_5896,N_4272,N_4203);
or U5897 (N_5897,N_4445,N_4627);
and U5898 (N_5898,N_4179,N_4569);
nor U5899 (N_5899,N_4159,N_4470);
nor U5900 (N_5900,N_4170,N_4604);
nor U5901 (N_5901,N_4462,N_4694);
and U5902 (N_5902,N_4227,N_4319);
or U5903 (N_5903,N_4996,N_4615);
nand U5904 (N_5904,N_4525,N_4521);
or U5905 (N_5905,N_4472,N_4126);
and U5906 (N_5906,N_4800,N_4963);
or U5907 (N_5907,N_4509,N_4914);
or U5908 (N_5908,N_4596,N_4258);
nand U5909 (N_5909,N_4142,N_4157);
and U5910 (N_5910,N_4744,N_4514);
nand U5911 (N_5911,N_4489,N_4448);
and U5912 (N_5912,N_4548,N_4761);
or U5913 (N_5913,N_4896,N_4169);
and U5914 (N_5914,N_4408,N_4883);
nand U5915 (N_5915,N_4954,N_4217);
nand U5916 (N_5916,N_4363,N_4394);
or U5917 (N_5917,N_4794,N_4317);
nor U5918 (N_5918,N_4820,N_4518);
or U5919 (N_5919,N_4598,N_4763);
or U5920 (N_5920,N_4932,N_4326);
nand U5921 (N_5921,N_4497,N_4301);
and U5922 (N_5922,N_4523,N_4344);
nor U5923 (N_5923,N_4512,N_4019);
nand U5924 (N_5924,N_4330,N_4992);
nor U5925 (N_5925,N_4839,N_4345);
or U5926 (N_5926,N_4822,N_4807);
nor U5927 (N_5927,N_4949,N_4145);
nor U5928 (N_5928,N_4831,N_4698);
or U5929 (N_5929,N_4164,N_4294);
and U5930 (N_5930,N_4215,N_4133);
nand U5931 (N_5931,N_4963,N_4295);
nor U5932 (N_5932,N_4604,N_4553);
nand U5933 (N_5933,N_4966,N_4135);
nor U5934 (N_5934,N_4045,N_4697);
nand U5935 (N_5935,N_4527,N_4403);
nor U5936 (N_5936,N_4950,N_4596);
or U5937 (N_5937,N_4822,N_4211);
and U5938 (N_5938,N_4303,N_4739);
nor U5939 (N_5939,N_4262,N_4273);
or U5940 (N_5940,N_4022,N_4083);
and U5941 (N_5941,N_4625,N_4042);
nand U5942 (N_5942,N_4478,N_4663);
nand U5943 (N_5943,N_4448,N_4862);
nor U5944 (N_5944,N_4140,N_4700);
nor U5945 (N_5945,N_4286,N_4795);
or U5946 (N_5946,N_4468,N_4432);
and U5947 (N_5947,N_4919,N_4852);
and U5948 (N_5948,N_4090,N_4274);
or U5949 (N_5949,N_4228,N_4979);
and U5950 (N_5950,N_4818,N_4686);
nand U5951 (N_5951,N_4910,N_4193);
or U5952 (N_5952,N_4110,N_4267);
or U5953 (N_5953,N_4676,N_4316);
nor U5954 (N_5954,N_4240,N_4608);
nand U5955 (N_5955,N_4668,N_4562);
nand U5956 (N_5956,N_4291,N_4461);
or U5957 (N_5957,N_4488,N_4372);
nand U5958 (N_5958,N_4786,N_4658);
and U5959 (N_5959,N_4294,N_4420);
nand U5960 (N_5960,N_4726,N_4614);
and U5961 (N_5961,N_4273,N_4337);
nor U5962 (N_5962,N_4030,N_4043);
and U5963 (N_5963,N_4377,N_4746);
and U5964 (N_5964,N_4380,N_4297);
nor U5965 (N_5965,N_4308,N_4625);
and U5966 (N_5966,N_4492,N_4723);
nand U5967 (N_5967,N_4106,N_4418);
nand U5968 (N_5968,N_4316,N_4110);
and U5969 (N_5969,N_4814,N_4372);
nor U5970 (N_5970,N_4171,N_4810);
and U5971 (N_5971,N_4788,N_4774);
and U5972 (N_5972,N_4489,N_4644);
or U5973 (N_5973,N_4123,N_4070);
nand U5974 (N_5974,N_4970,N_4745);
and U5975 (N_5975,N_4743,N_4675);
and U5976 (N_5976,N_4000,N_4309);
nand U5977 (N_5977,N_4992,N_4141);
nor U5978 (N_5978,N_4376,N_4873);
or U5979 (N_5979,N_4755,N_4220);
nand U5980 (N_5980,N_4995,N_4124);
nor U5981 (N_5981,N_4845,N_4624);
or U5982 (N_5982,N_4310,N_4456);
nor U5983 (N_5983,N_4986,N_4203);
or U5984 (N_5984,N_4109,N_4303);
nand U5985 (N_5985,N_4746,N_4745);
nor U5986 (N_5986,N_4603,N_4906);
nand U5987 (N_5987,N_4438,N_4445);
and U5988 (N_5988,N_4222,N_4704);
and U5989 (N_5989,N_4453,N_4540);
or U5990 (N_5990,N_4031,N_4842);
nor U5991 (N_5991,N_4043,N_4591);
nand U5992 (N_5992,N_4473,N_4233);
and U5993 (N_5993,N_4485,N_4725);
nand U5994 (N_5994,N_4602,N_4591);
nor U5995 (N_5995,N_4021,N_4988);
and U5996 (N_5996,N_4863,N_4071);
nor U5997 (N_5997,N_4346,N_4965);
nor U5998 (N_5998,N_4675,N_4349);
nor U5999 (N_5999,N_4641,N_4428);
nor U6000 (N_6000,N_5708,N_5989);
nor U6001 (N_6001,N_5481,N_5260);
nand U6002 (N_6002,N_5460,N_5316);
nor U6003 (N_6003,N_5727,N_5298);
and U6004 (N_6004,N_5326,N_5006);
nand U6005 (N_6005,N_5485,N_5158);
nand U6006 (N_6006,N_5056,N_5586);
or U6007 (N_6007,N_5574,N_5254);
nor U6008 (N_6008,N_5930,N_5129);
or U6009 (N_6009,N_5855,N_5279);
or U6010 (N_6010,N_5303,N_5300);
nor U6011 (N_6011,N_5729,N_5691);
or U6012 (N_6012,N_5422,N_5933);
nor U6013 (N_6013,N_5712,N_5513);
and U6014 (N_6014,N_5951,N_5847);
and U6015 (N_6015,N_5700,N_5709);
or U6016 (N_6016,N_5366,N_5264);
or U6017 (N_6017,N_5236,N_5957);
nor U6018 (N_6018,N_5868,N_5807);
or U6019 (N_6019,N_5151,N_5331);
or U6020 (N_6020,N_5813,N_5530);
and U6021 (N_6021,N_5580,N_5737);
and U6022 (N_6022,N_5561,N_5535);
or U6023 (N_6023,N_5613,N_5378);
nand U6024 (N_6024,N_5549,N_5314);
nand U6025 (N_6025,N_5541,N_5131);
xnor U6026 (N_6026,N_5084,N_5423);
nor U6027 (N_6027,N_5520,N_5754);
nor U6028 (N_6028,N_5845,N_5836);
and U6029 (N_6029,N_5653,N_5221);
or U6030 (N_6030,N_5685,N_5942);
xnor U6031 (N_6031,N_5698,N_5041);
nor U6032 (N_6032,N_5648,N_5705);
nor U6033 (N_6033,N_5343,N_5462);
or U6034 (N_6034,N_5826,N_5628);
nor U6035 (N_6035,N_5852,N_5644);
and U6036 (N_6036,N_5514,N_5843);
and U6037 (N_6037,N_5308,N_5089);
or U6038 (N_6038,N_5229,N_5101);
or U6039 (N_6039,N_5220,N_5658);
nor U6040 (N_6040,N_5878,N_5529);
and U6041 (N_6041,N_5725,N_5287);
nor U6042 (N_6042,N_5562,N_5367);
nor U6043 (N_6043,N_5039,N_5266);
nor U6044 (N_6044,N_5295,N_5659);
and U6045 (N_6045,N_5002,N_5200);
nand U6046 (N_6046,N_5823,N_5127);
nand U6047 (N_6047,N_5860,N_5392);
or U6048 (N_6048,N_5243,N_5251);
and U6049 (N_6049,N_5110,N_5741);
nor U6050 (N_6050,N_5450,N_5998);
or U6051 (N_6051,N_5456,N_5497);
and U6052 (N_6052,N_5978,N_5862);
nor U6053 (N_6053,N_5591,N_5111);
or U6054 (N_6054,N_5435,N_5437);
nand U6055 (N_6055,N_5160,N_5687);
or U6056 (N_6056,N_5502,N_5386);
and U6057 (N_6057,N_5067,N_5176);
and U6058 (N_6058,N_5155,N_5371);
nor U6059 (N_6059,N_5352,N_5442);
nand U6060 (N_6060,N_5947,N_5233);
nor U6061 (N_6061,N_5738,N_5771);
nor U6062 (N_6062,N_5184,N_5461);
nand U6063 (N_6063,N_5987,N_5165);
and U6064 (N_6064,N_5025,N_5595);
and U6065 (N_6065,N_5390,N_5969);
or U6066 (N_6066,N_5203,N_5364);
or U6067 (N_6067,N_5795,N_5861);
or U6068 (N_6068,N_5752,N_5802);
nand U6069 (N_6069,N_5894,N_5805);
or U6070 (N_6070,N_5003,N_5865);
or U6071 (N_6071,N_5936,N_5692);
nand U6072 (N_6072,N_5032,N_5268);
or U6073 (N_6073,N_5672,N_5666);
or U6074 (N_6074,N_5249,N_5822);
nand U6075 (N_6075,N_5699,N_5052);
and U6076 (N_6076,N_5743,N_5915);
nand U6077 (N_6077,N_5693,N_5985);
or U6078 (N_6078,N_5825,N_5026);
or U6079 (N_6079,N_5139,N_5647);
or U6080 (N_6080,N_5408,N_5244);
nor U6081 (N_6081,N_5714,N_5001);
and U6082 (N_6082,N_5179,N_5726);
or U6083 (N_6083,N_5100,N_5590);
nor U6084 (N_6084,N_5385,N_5850);
nor U6085 (N_6085,N_5370,N_5059);
and U6086 (N_6086,N_5286,N_5546);
nor U6087 (N_6087,N_5926,N_5169);
nand U6088 (N_6088,N_5764,N_5810);
nor U6089 (N_6089,N_5500,N_5818);
nand U6090 (N_6090,N_5080,N_5950);
or U6091 (N_6091,N_5465,N_5539);
or U6092 (N_6092,N_5064,N_5660);
and U6093 (N_6093,N_5381,N_5769);
nand U6094 (N_6094,N_5469,N_5128);
or U6095 (N_6095,N_5479,N_5047);
nand U6096 (N_6096,N_5828,N_5763);
nor U6097 (N_6097,N_5216,N_5282);
nand U6098 (N_6098,N_5866,N_5716);
and U6099 (N_6099,N_5225,N_5528);
nand U6100 (N_6100,N_5887,N_5911);
nor U6101 (N_6101,N_5191,N_5452);
or U6102 (N_6102,N_5411,N_5831);
nand U6103 (N_6103,N_5309,N_5929);
or U6104 (N_6104,N_5154,N_5639);
nor U6105 (N_6105,N_5748,N_5811);
and U6106 (N_6106,N_5982,N_5046);
and U6107 (N_6107,N_5710,N_5339);
nand U6108 (N_6108,N_5388,N_5044);
nor U6109 (N_6109,N_5271,N_5182);
nand U6110 (N_6110,N_5227,N_5173);
nand U6111 (N_6111,N_5917,N_5324);
nand U6112 (N_6112,N_5554,N_5076);
or U6113 (N_6113,N_5839,N_5609);
and U6114 (N_6114,N_5416,N_5816);
nand U6115 (N_6115,N_5990,N_5360);
nand U6116 (N_6116,N_5108,N_5099);
nand U6117 (N_6117,N_5149,N_5035);
nor U6118 (N_6118,N_5401,N_5317);
nor U6119 (N_6119,N_5780,N_5731);
and U6120 (N_6120,N_5820,N_5621);
and U6121 (N_6121,N_5235,N_5143);
or U6122 (N_6122,N_5397,N_5877);
nand U6123 (N_6123,N_5570,N_5890);
or U6124 (N_6124,N_5328,N_5923);
nand U6125 (N_6125,N_5453,N_5728);
nand U6126 (N_6126,N_5842,N_5956);
nand U6127 (N_6127,N_5840,N_5174);
or U6128 (N_6128,N_5185,N_5694);
and U6129 (N_6129,N_5637,N_5965);
nand U6130 (N_6130,N_5740,N_5602);
nor U6131 (N_6131,N_5292,N_5993);
and U6132 (N_6132,N_5796,N_5019);
and U6133 (N_6133,N_5622,N_5893);
nor U6134 (N_6134,N_5419,N_5794);
and U6135 (N_6135,N_5038,N_5278);
or U6136 (N_6136,N_5338,N_5848);
xor U6137 (N_6137,N_5955,N_5082);
nand U6138 (N_6138,N_5208,N_5130);
nor U6139 (N_6139,N_5967,N_5593);
nor U6140 (N_6140,N_5997,N_5121);
nand U6141 (N_6141,N_5575,N_5104);
nor U6142 (N_6142,N_5405,N_5856);
nor U6143 (N_6143,N_5272,N_5373);
and U6144 (N_6144,N_5302,N_5899);
nor U6145 (N_6145,N_5787,N_5567);
and U6146 (N_6146,N_5074,N_5635);
nor U6147 (N_6147,N_5719,N_5161);
or U6148 (N_6148,N_5582,N_5194);
or U6149 (N_6149,N_5318,N_5629);
and U6150 (N_6150,N_5237,N_5667);
nand U6151 (N_6151,N_5147,N_5142);
nand U6152 (N_6152,N_5234,N_5515);
and U6153 (N_6153,N_5902,N_5885);
and U6154 (N_6154,N_5336,N_5171);
nor U6155 (N_6155,N_5946,N_5977);
nand U6156 (N_6156,N_5106,N_5578);
nor U6157 (N_6157,N_5276,N_5480);
nor U6158 (N_6158,N_5070,N_5310);
and U6159 (N_6159,N_5913,N_5772);
nand U6160 (N_6160,N_5062,N_5673);
or U6161 (N_6161,N_5141,N_5132);
xnor U6162 (N_6162,N_5626,N_5471);
nand U6163 (N_6163,N_5550,N_5784);
nand U6164 (N_6164,N_5651,N_5472);
or U6165 (N_6165,N_5611,N_5410);
or U6166 (N_6166,N_5320,N_5501);
or U6167 (N_6167,N_5511,N_5995);
or U6168 (N_6168,N_5614,N_5572);
or U6169 (N_6169,N_5928,N_5706);
and U6170 (N_6170,N_5542,N_5674);
nor U6171 (N_6171,N_5724,N_5863);
nor U6172 (N_6172,N_5844,N_5421);
nand U6173 (N_6173,N_5544,N_5778);
and U6174 (N_6174,N_5113,N_5183);
and U6175 (N_6175,N_5322,N_5376);
nand U6176 (N_6176,N_5555,N_5833);
and U6177 (N_6177,N_5975,N_5342);
nor U6178 (N_6178,N_5464,N_5333);
nand U6179 (N_6179,N_5652,N_5808);
nor U6180 (N_6180,N_5896,N_5892);
or U6181 (N_6181,N_5841,N_5349);
or U6182 (N_6182,N_5873,N_5092);
xnor U6183 (N_6183,N_5558,N_5157);
and U6184 (N_6184,N_5536,N_5301);
and U6185 (N_6185,N_5350,N_5812);
xor U6186 (N_6186,N_5832,N_5164);
nor U6187 (N_6187,N_5396,N_5897);
xor U6188 (N_6188,N_5252,N_5988);
and U6189 (N_6189,N_5016,N_5400);
xnor U6190 (N_6190,N_5238,N_5087);
nand U6191 (N_6191,N_5023,N_5766);
nor U6192 (N_6192,N_5524,N_5145);
nor U6193 (N_6193,N_5077,N_5525);
and U6194 (N_6194,N_5334,N_5585);
or U6195 (N_6195,N_5703,N_5362);
or U6196 (N_6196,N_5283,N_5478);
or U6197 (N_6197,N_5526,N_5008);
nand U6198 (N_6198,N_5938,N_5009);
and U6199 (N_6199,N_5207,N_5224);
nand U6200 (N_6200,N_5718,N_5259);
nand U6201 (N_6201,N_5905,N_5623);
nand U6202 (N_6202,N_5284,N_5053);
or U6203 (N_6203,N_5455,N_5888);
and U6204 (N_6204,N_5918,N_5109);
nor U6205 (N_6205,N_5305,N_5230);
and U6206 (N_6206,N_5940,N_5323);
nand U6207 (N_6207,N_5196,N_5846);
nand U6208 (N_6208,N_5167,N_5968);
nor U6209 (N_6209,N_5085,N_5617);
xnor U6210 (N_6210,N_5270,N_5488);
nand U6211 (N_6211,N_5944,N_5199);
or U6212 (N_6212,N_5935,N_5922);
nand U6213 (N_6213,N_5215,N_5715);
nor U6214 (N_6214,N_5600,N_5296);
nand U6215 (N_6215,N_5767,N_5809);
or U6216 (N_6216,N_5246,N_5311);
nor U6217 (N_6217,N_5697,N_5914);
and U6218 (N_6218,N_5159,N_5656);
nor U6219 (N_6219,N_5289,N_5393);
and U6220 (N_6220,N_5800,N_5218);
nor U6221 (N_6221,N_5081,N_5049);
and U6222 (N_6222,N_5248,N_5152);
and U6223 (N_6223,N_5949,N_5886);
nand U6224 (N_6224,N_5912,N_5180);
nor U6225 (N_6225,N_5882,N_5739);
and U6226 (N_6226,N_5624,N_5186);
or U6227 (N_6227,N_5124,N_5557);
nor U6228 (N_6228,N_5730,N_5007);
nor U6229 (N_6229,N_5904,N_5854);
or U6230 (N_6230,N_5448,N_5680);
nand U6231 (N_6231,N_5347,N_5496);
nor U6232 (N_6232,N_5083,N_5432);
nor U6233 (N_6233,N_5773,N_5020);
and U6234 (N_6234,N_5701,N_5596);
nor U6235 (N_6235,N_5948,N_5753);
and U6236 (N_6236,N_5040,N_5118);
nand U6237 (N_6237,N_5239,N_5758);
or U6238 (N_6238,N_5636,N_5189);
nand U6239 (N_6239,N_5153,N_5615);
and U6240 (N_6240,N_5677,N_5190);
nor U6241 (N_6241,N_5201,N_5655);
or U6242 (N_6242,N_5060,N_5332);
and U6243 (N_6243,N_5664,N_5241);
or U6244 (N_6244,N_5503,N_5610);
nor U6245 (N_6245,N_5671,N_5906);
nor U6246 (N_6246,N_5799,N_5499);
and U6247 (N_6247,N_5090,N_5304);
nor U6248 (N_6248,N_5919,N_5420);
nor U6249 (N_6249,N_5434,N_5369);
nor U6250 (N_6250,N_5869,N_5365);
nor U6251 (N_6251,N_5732,N_5981);
nor U6252 (N_6252,N_5093,N_5195);
or U6253 (N_6253,N_5625,N_5983);
or U6254 (N_6254,N_5105,N_5711);
or U6255 (N_6255,N_5964,N_5924);
nor U6256 (N_6256,N_5379,N_5954);
nor U6257 (N_6257,N_5489,N_5538);
nor U6258 (N_6258,N_5454,N_5073);
nand U6259 (N_6259,N_5927,N_5872);
nor U6260 (N_6260,N_5690,N_5398);
nand U6261 (N_6261,N_5148,N_5315);
nor U6262 (N_6262,N_5493,N_5193);
or U6263 (N_6263,N_5353,N_5755);
or U6264 (N_6264,N_5556,N_5245);
nor U6265 (N_6265,N_5920,N_5116);
or U6266 (N_6266,N_5908,N_5181);
or U6267 (N_6267,N_5117,N_5441);
or U6268 (N_6268,N_5088,N_5330);
nand U6269 (N_6269,N_5058,N_5722);
or U6270 (N_6270,N_5150,N_5521);
nand U6271 (N_6271,N_5065,N_5290);
and U6272 (N_6272,N_5765,N_5681);
nor U6273 (N_6273,N_5669,N_5403);
nor U6274 (N_6274,N_5806,N_5140);
and U6275 (N_6275,N_5991,N_5280);
and U6276 (N_6276,N_5394,N_5518);
or U6277 (N_6277,N_5548,N_5688);
nor U6278 (N_6278,N_5354,N_5135);
nand U6279 (N_6279,N_5939,N_5391);
or U6280 (N_6280,N_5048,N_5146);
nand U6281 (N_6281,N_5783,N_5475);
nand U6282 (N_6282,N_5859,N_5592);
or U6283 (N_6283,N_5704,N_5382);
and U6284 (N_6284,N_5986,N_5976);
and U6285 (N_6285,N_5275,N_5683);
nor U6286 (N_6286,N_5774,N_5760);
nor U6287 (N_6287,N_5803,N_5895);
and U6288 (N_6288,N_5909,N_5013);
nand U6289 (N_6289,N_5576,N_5531);
and U6290 (N_6290,N_5086,N_5963);
or U6291 (N_6291,N_5258,N_5668);
nor U6292 (N_6292,N_5202,N_5830);
and U6293 (N_6293,N_5867,N_5492);
nor U6294 (N_6294,N_5356,N_5720);
nor U6295 (N_6295,N_5000,N_5075);
nor U6296 (N_6296,N_5407,N_5375);
and U6297 (N_6297,N_5430,N_5790);
or U6298 (N_6298,N_5770,N_5504);
or U6299 (N_6299,N_5584,N_5037);
or U6300 (N_6300,N_5126,N_5876);
or U6301 (N_6301,N_5785,N_5864);
nor U6302 (N_6302,N_5534,N_5506);
xor U6303 (N_6303,N_5319,N_5024);
or U6304 (N_6304,N_5545,N_5490);
or U6305 (N_6305,N_5214,N_5482);
and U6306 (N_6306,N_5979,N_5476);
and U6307 (N_6307,N_5115,N_5281);
nor U6308 (N_6308,N_5120,N_5027);
or U6309 (N_6309,N_5011,N_5022);
nand U6310 (N_6310,N_5446,N_5723);
nand U6311 (N_6311,N_5945,N_5066);
or U6312 (N_6312,N_5091,N_5903);
and U6313 (N_6313,N_5654,N_5829);
nand U6314 (N_6314,N_5566,N_5547);
xnor U6315 (N_6315,N_5607,N_5288);
and U6316 (N_6316,N_5695,N_5750);
nor U6317 (N_6317,N_5870,N_5910);
and U6318 (N_6318,N_5114,N_5491);
or U6319 (N_6319,N_5034,N_5449);
nand U6320 (N_6320,N_5177,N_5495);
or U6321 (N_6321,N_5533,N_5387);
nand U6322 (N_6322,N_5953,N_5368);
nor U6323 (N_6323,N_5606,N_5198);
or U6324 (N_6324,N_5033,N_5959);
nand U6325 (N_6325,N_5263,N_5267);
nand U6326 (N_6326,N_5507,N_5540);
nor U6327 (N_6327,N_5571,N_5222);
or U6328 (N_6328,N_5425,N_5851);
nor U6329 (N_6329,N_5634,N_5992);
nand U6330 (N_6330,N_5801,N_5791);
nor U6331 (N_6331,N_5605,N_5358);
nand U6332 (N_6332,N_5223,N_5473);
nor U6333 (N_6333,N_5916,N_5329);
nand U6334 (N_6334,N_5641,N_5247);
or U6335 (N_6335,N_5713,N_5451);
nor U6336 (N_6336,N_5262,N_5925);
and U6337 (N_6337,N_5028,N_5341);
nor U6338 (N_6338,N_5972,N_5068);
or U6339 (N_6339,N_5696,N_5657);
nor U6340 (N_6340,N_5071,N_5891);
nor U6341 (N_6341,N_5445,N_5344);
nor U6342 (N_6342,N_5178,N_5880);
nand U6343 (N_6343,N_5487,N_5523);
nor U6344 (N_6344,N_5036,N_5779);
nand U6345 (N_6345,N_5057,N_5686);
and U6346 (N_6346,N_5537,N_5678);
nor U6347 (N_6347,N_5431,N_5857);
nor U6348 (N_6348,N_5819,N_5406);
or U6349 (N_6349,N_5616,N_5608);
nand U6350 (N_6350,N_5901,N_5874);
and U6351 (N_6351,N_5505,N_5662);
nand U6352 (N_6352,N_5881,N_5166);
nor U6353 (N_6353,N_5751,N_5014);
and U6354 (N_6354,N_5119,N_5638);
and U6355 (N_6355,N_5340,N_5568);
nor U6356 (N_6356,N_5589,N_5072);
and U6357 (N_6357,N_5138,N_5588);
and U6358 (N_6358,N_5961,N_5426);
and U6359 (N_6359,N_5122,N_5351);
and U6360 (N_6360,N_5134,N_5594);
nor U6361 (N_6361,N_5745,N_5412);
and U6362 (N_6362,N_5941,N_5043);
or U6363 (N_6363,N_5389,N_5543);
or U6364 (N_6364,N_5458,N_5838);
nor U6365 (N_6365,N_5598,N_5879);
nor U6366 (N_6366,N_5642,N_5021);
nor U6367 (N_6367,N_5962,N_5508);
nor U6368 (N_6368,N_5670,N_5619);
or U6369 (N_6369,N_5675,N_5042);
nor U6370 (N_6370,N_5551,N_5439);
nor U6371 (N_6371,N_5418,N_5291);
and U6372 (N_6372,N_5684,N_5934);
or U6373 (N_6373,N_5834,N_5553);
and U6374 (N_6374,N_5374,N_5837);
nand U6375 (N_6375,N_5413,N_5232);
nor U6376 (N_6376,N_5966,N_5274);
and U6377 (N_6377,N_5597,N_5427);
and U6378 (N_6378,N_5098,N_5372);
or U6379 (N_6379,N_5971,N_5133);
and U6380 (N_6380,N_5815,N_5717);
or U6381 (N_6381,N_5477,N_5433);
nor U6382 (N_6382,N_5015,N_5633);
or U6383 (N_6383,N_5960,N_5261);
nand U6384 (N_6384,N_5383,N_5883);
nand U6385 (N_6385,N_5436,N_5197);
and U6386 (N_6386,N_5996,N_5294);
and U6387 (N_6387,N_5188,N_5733);
nand U6388 (N_6388,N_5483,N_5459);
and U6389 (N_6389,N_5835,N_5429);
nand U6390 (N_6390,N_5335,N_5853);
and U6391 (N_6391,N_5798,N_5577);
and U6392 (N_6392,N_5273,N_5463);
or U6393 (N_6393,N_5226,N_5587);
nor U6394 (N_6394,N_5564,N_5004);
nand U6395 (N_6395,N_5973,N_5984);
and U6396 (N_6396,N_5519,N_5095);
nor U6397 (N_6397,N_5631,N_5307);
and U6398 (N_6398,N_5620,N_5645);
nor U6399 (N_6399,N_5781,N_5559);
and U6400 (N_6400,N_5676,N_5399);
nor U6401 (N_6401,N_5030,N_5102);
nor U6402 (N_6402,N_5005,N_5522);
and U6403 (N_6403,N_5470,N_5438);
nor U6404 (N_6404,N_5156,N_5467);
nand U6405 (N_6405,N_5096,N_5395);
and U6406 (N_6406,N_5211,N_5630);
nor U6407 (N_6407,N_5974,N_5192);
nand U6408 (N_6408,N_5827,N_5797);
or U6409 (N_6409,N_5689,N_5516);
or U6410 (N_6410,N_5125,N_5205);
and U6411 (N_6411,N_5377,N_5123);
nor U6412 (N_6412,N_5168,N_5231);
nor U6413 (N_6413,N_5756,N_5494);
nor U6414 (N_6414,N_5943,N_5466);
nand U6415 (N_6415,N_5484,N_5665);
nor U6416 (N_6416,N_5170,N_5228);
or U6417 (N_6417,N_5618,N_5424);
or U6418 (N_6418,N_5632,N_5210);
or U6419 (N_6419,N_5257,N_5277);
and U6420 (N_6420,N_5612,N_5348);
nor U6421 (N_6421,N_5599,N_5579);
nand U6422 (N_6422,N_5649,N_5443);
or U6423 (N_6423,N_5824,N_5817);
nor U6424 (N_6424,N_5786,N_5643);
nand U6425 (N_6425,N_5162,N_5428);
nand U6426 (N_6426,N_5144,N_5012);
nor U6427 (N_6427,N_5734,N_5094);
nand U6428 (N_6428,N_5898,N_5137);
nand U6429 (N_6429,N_5415,N_5361);
nand U6430 (N_6430,N_5355,N_5363);
nand U6431 (N_6431,N_5517,N_5747);
nor U6432 (N_6432,N_5735,N_5849);
nand U6433 (N_6433,N_5889,N_5440);
xor U6434 (N_6434,N_5312,N_5107);
and U6435 (N_6435,N_5958,N_5097);
nand U6436 (N_6436,N_5468,N_5789);
nand U6437 (N_6437,N_5163,N_5414);
and U6438 (N_6438,N_5213,N_5079);
nand U6439 (N_6439,N_5017,N_5744);
nor U6440 (N_6440,N_5409,N_5931);
or U6441 (N_6441,N_5900,N_5661);
nor U6442 (N_6442,N_5560,N_5627);
nand U6443 (N_6443,N_5029,N_5907);
and U6444 (N_6444,N_5136,N_5736);
or U6445 (N_6445,N_5569,N_5782);
and U6446 (N_6446,N_5327,N_5474);
nand U6447 (N_6447,N_5788,N_5821);
or U6448 (N_6448,N_5253,N_5937);
and U6449 (N_6449,N_5884,N_5417);
nand U6450 (N_6450,N_5103,N_5209);
nor U6451 (N_6451,N_5775,N_5293);
and U6452 (N_6452,N_5804,N_5498);
nand U6453 (N_6453,N_5061,N_5357);
nor U6454 (N_6454,N_5583,N_5050);
and U6455 (N_6455,N_5952,N_5112);
and U6456 (N_6456,N_5250,N_5707);
or U6457 (N_6457,N_5325,N_5871);
nor U6458 (N_6458,N_5175,N_5762);
nor U6459 (N_6459,N_5646,N_5345);
and U6460 (N_6460,N_5980,N_5682);
nand U6461 (N_6461,N_5285,N_5742);
nand U6462 (N_6462,N_5814,N_5240);
nor U6463 (N_6463,N_5486,N_5206);
nand U6464 (N_6464,N_5078,N_5761);
nor U6465 (N_6465,N_5212,N_5759);
nand U6466 (N_6466,N_5217,N_5932);
nor U6467 (N_6467,N_5512,N_5402);
or U6468 (N_6468,N_5994,N_5702);
nand U6469 (N_6469,N_5601,N_5063);
and U6470 (N_6470,N_5242,N_5858);
nor U6471 (N_6471,N_5269,N_5970);
and U6472 (N_6472,N_5337,N_5999);
and U6473 (N_6473,N_5792,N_5777);
or U6474 (N_6474,N_5010,N_5380);
nand U6475 (N_6475,N_5297,N_5055);
nor U6476 (N_6476,N_5204,N_5527);
and U6477 (N_6477,N_5404,N_5444);
nor U6478 (N_6478,N_5757,N_5256);
and U6479 (N_6479,N_5603,N_5172);
or U6480 (N_6480,N_5650,N_5776);
nor U6481 (N_6481,N_5018,N_5359);
nor U6482 (N_6482,N_5663,N_5069);
xnor U6483 (N_6483,N_5187,N_5573);
nand U6484 (N_6484,N_5563,N_5510);
or U6485 (N_6485,N_5299,N_5255);
nor U6486 (N_6486,N_5346,N_5532);
or U6487 (N_6487,N_5581,N_5219);
xor U6488 (N_6488,N_5875,N_5051);
and U6489 (N_6489,N_5321,N_5265);
nor U6490 (N_6490,N_5509,N_5447);
or U6491 (N_6491,N_5384,N_5306);
nor U6492 (N_6492,N_5640,N_5746);
and U6493 (N_6493,N_5721,N_5457);
and U6494 (N_6494,N_5921,N_5768);
nor U6495 (N_6495,N_5749,N_5313);
and U6496 (N_6496,N_5565,N_5679);
or U6497 (N_6497,N_5552,N_5604);
and U6498 (N_6498,N_5054,N_5793);
or U6499 (N_6499,N_5031,N_5045);
nor U6500 (N_6500,N_5165,N_5051);
xnor U6501 (N_6501,N_5096,N_5586);
and U6502 (N_6502,N_5310,N_5571);
or U6503 (N_6503,N_5595,N_5281);
nand U6504 (N_6504,N_5574,N_5165);
nand U6505 (N_6505,N_5750,N_5125);
nor U6506 (N_6506,N_5400,N_5180);
nand U6507 (N_6507,N_5962,N_5413);
or U6508 (N_6508,N_5014,N_5883);
nand U6509 (N_6509,N_5457,N_5892);
and U6510 (N_6510,N_5911,N_5648);
nor U6511 (N_6511,N_5982,N_5853);
and U6512 (N_6512,N_5976,N_5847);
nand U6513 (N_6513,N_5594,N_5933);
or U6514 (N_6514,N_5642,N_5467);
and U6515 (N_6515,N_5289,N_5345);
or U6516 (N_6516,N_5898,N_5802);
nand U6517 (N_6517,N_5321,N_5205);
and U6518 (N_6518,N_5156,N_5157);
nand U6519 (N_6519,N_5764,N_5599);
nand U6520 (N_6520,N_5912,N_5184);
or U6521 (N_6521,N_5566,N_5349);
and U6522 (N_6522,N_5286,N_5095);
and U6523 (N_6523,N_5595,N_5971);
and U6524 (N_6524,N_5488,N_5683);
nand U6525 (N_6525,N_5683,N_5659);
and U6526 (N_6526,N_5035,N_5532);
nand U6527 (N_6527,N_5752,N_5573);
or U6528 (N_6528,N_5538,N_5464);
xnor U6529 (N_6529,N_5272,N_5092);
nor U6530 (N_6530,N_5339,N_5938);
or U6531 (N_6531,N_5436,N_5487);
nor U6532 (N_6532,N_5218,N_5799);
or U6533 (N_6533,N_5700,N_5356);
or U6534 (N_6534,N_5958,N_5882);
and U6535 (N_6535,N_5847,N_5458);
nor U6536 (N_6536,N_5355,N_5729);
or U6537 (N_6537,N_5398,N_5089);
and U6538 (N_6538,N_5660,N_5716);
and U6539 (N_6539,N_5128,N_5500);
nand U6540 (N_6540,N_5311,N_5767);
nor U6541 (N_6541,N_5769,N_5783);
and U6542 (N_6542,N_5550,N_5703);
nor U6543 (N_6543,N_5250,N_5003);
nand U6544 (N_6544,N_5596,N_5612);
nand U6545 (N_6545,N_5682,N_5478);
or U6546 (N_6546,N_5975,N_5280);
nand U6547 (N_6547,N_5034,N_5954);
nand U6548 (N_6548,N_5187,N_5262);
nor U6549 (N_6549,N_5334,N_5950);
nor U6550 (N_6550,N_5077,N_5319);
nor U6551 (N_6551,N_5217,N_5924);
or U6552 (N_6552,N_5556,N_5454);
nand U6553 (N_6553,N_5306,N_5739);
nand U6554 (N_6554,N_5066,N_5342);
or U6555 (N_6555,N_5853,N_5184);
nand U6556 (N_6556,N_5165,N_5597);
nand U6557 (N_6557,N_5138,N_5971);
nor U6558 (N_6558,N_5101,N_5320);
nand U6559 (N_6559,N_5698,N_5214);
or U6560 (N_6560,N_5330,N_5596);
nand U6561 (N_6561,N_5376,N_5541);
nor U6562 (N_6562,N_5465,N_5199);
nand U6563 (N_6563,N_5946,N_5950);
and U6564 (N_6564,N_5123,N_5964);
nor U6565 (N_6565,N_5300,N_5614);
or U6566 (N_6566,N_5746,N_5962);
or U6567 (N_6567,N_5449,N_5394);
nor U6568 (N_6568,N_5232,N_5113);
or U6569 (N_6569,N_5579,N_5874);
nor U6570 (N_6570,N_5920,N_5126);
and U6571 (N_6571,N_5965,N_5180);
nor U6572 (N_6572,N_5131,N_5539);
nor U6573 (N_6573,N_5083,N_5495);
nand U6574 (N_6574,N_5837,N_5857);
and U6575 (N_6575,N_5599,N_5169);
or U6576 (N_6576,N_5643,N_5237);
and U6577 (N_6577,N_5370,N_5504);
nor U6578 (N_6578,N_5135,N_5079);
and U6579 (N_6579,N_5531,N_5061);
nor U6580 (N_6580,N_5537,N_5432);
or U6581 (N_6581,N_5728,N_5557);
nand U6582 (N_6582,N_5324,N_5634);
and U6583 (N_6583,N_5126,N_5901);
or U6584 (N_6584,N_5660,N_5932);
or U6585 (N_6585,N_5765,N_5337);
or U6586 (N_6586,N_5292,N_5311);
nor U6587 (N_6587,N_5662,N_5878);
nand U6588 (N_6588,N_5377,N_5686);
and U6589 (N_6589,N_5673,N_5869);
nand U6590 (N_6590,N_5534,N_5029);
nand U6591 (N_6591,N_5910,N_5599);
xor U6592 (N_6592,N_5287,N_5772);
and U6593 (N_6593,N_5024,N_5478);
and U6594 (N_6594,N_5498,N_5636);
or U6595 (N_6595,N_5115,N_5097);
nand U6596 (N_6596,N_5542,N_5026);
nand U6597 (N_6597,N_5046,N_5048);
xor U6598 (N_6598,N_5390,N_5515);
nor U6599 (N_6599,N_5611,N_5315);
or U6600 (N_6600,N_5920,N_5903);
nor U6601 (N_6601,N_5816,N_5946);
or U6602 (N_6602,N_5894,N_5048);
nor U6603 (N_6603,N_5000,N_5057);
or U6604 (N_6604,N_5436,N_5259);
nand U6605 (N_6605,N_5866,N_5025);
or U6606 (N_6606,N_5101,N_5828);
and U6607 (N_6607,N_5421,N_5107);
or U6608 (N_6608,N_5609,N_5143);
and U6609 (N_6609,N_5876,N_5908);
nor U6610 (N_6610,N_5376,N_5007);
nand U6611 (N_6611,N_5575,N_5756);
nand U6612 (N_6612,N_5494,N_5323);
or U6613 (N_6613,N_5216,N_5752);
nand U6614 (N_6614,N_5155,N_5854);
and U6615 (N_6615,N_5784,N_5475);
or U6616 (N_6616,N_5142,N_5562);
or U6617 (N_6617,N_5618,N_5740);
or U6618 (N_6618,N_5226,N_5103);
nor U6619 (N_6619,N_5807,N_5419);
nand U6620 (N_6620,N_5864,N_5924);
nor U6621 (N_6621,N_5921,N_5701);
nand U6622 (N_6622,N_5835,N_5481);
or U6623 (N_6623,N_5004,N_5755);
nand U6624 (N_6624,N_5059,N_5274);
nand U6625 (N_6625,N_5042,N_5917);
or U6626 (N_6626,N_5548,N_5079);
or U6627 (N_6627,N_5088,N_5051);
nand U6628 (N_6628,N_5922,N_5806);
nor U6629 (N_6629,N_5257,N_5328);
nor U6630 (N_6630,N_5402,N_5116);
nor U6631 (N_6631,N_5740,N_5289);
or U6632 (N_6632,N_5863,N_5597);
nor U6633 (N_6633,N_5638,N_5939);
nor U6634 (N_6634,N_5809,N_5867);
nand U6635 (N_6635,N_5707,N_5166);
nor U6636 (N_6636,N_5491,N_5776);
nor U6637 (N_6637,N_5427,N_5975);
or U6638 (N_6638,N_5137,N_5241);
nor U6639 (N_6639,N_5245,N_5855);
nor U6640 (N_6640,N_5897,N_5976);
and U6641 (N_6641,N_5197,N_5056);
or U6642 (N_6642,N_5791,N_5674);
or U6643 (N_6643,N_5741,N_5556);
and U6644 (N_6644,N_5744,N_5881);
and U6645 (N_6645,N_5775,N_5852);
nor U6646 (N_6646,N_5768,N_5588);
and U6647 (N_6647,N_5801,N_5815);
nor U6648 (N_6648,N_5368,N_5992);
or U6649 (N_6649,N_5442,N_5121);
nand U6650 (N_6650,N_5668,N_5231);
and U6651 (N_6651,N_5908,N_5043);
and U6652 (N_6652,N_5969,N_5214);
or U6653 (N_6653,N_5156,N_5315);
or U6654 (N_6654,N_5001,N_5763);
xor U6655 (N_6655,N_5311,N_5263);
nor U6656 (N_6656,N_5789,N_5017);
nand U6657 (N_6657,N_5743,N_5732);
nand U6658 (N_6658,N_5924,N_5643);
nand U6659 (N_6659,N_5849,N_5243);
and U6660 (N_6660,N_5392,N_5126);
nor U6661 (N_6661,N_5434,N_5486);
and U6662 (N_6662,N_5004,N_5837);
nor U6663 (N_6663,N_5207,N_5494);
or U6664 (N_6664,N_5971,N_5520);
or U6665 (N_6665,N_5943,N_5119);
and U6666 (N_6666,N_5803,N_5917);
or U6667 (N_6667,N_5413,N_5070);
or U6668 (N_6668,N_5027,N_5692);
nor U6669 (N_6669,N_5086,N_5444);
and U6670 (N_6670,N_5505,N_5424);
or U6671 (N_6671,N_5029,N_5824);
or U6672 (N_6672,N_5844,N_5549);
and U6673 (N_6673,N_5706,N_5420);
nor U6674 (N_6674,N_5116,N_5756);
nor U6675 (N_6675,N_5379,N_5601);
and U6676 (N_6676,N_5274,N_5932);
and U6677 (N_6677,N_5386,N_5245);
and U6678 (N_6678,N_5144,N_5765);
or U6679 (N_6679,N_5591,N_5838);
nand U6680 (N_6680,N_5466,N_5932);
nand U6681 (N_6681,N_5661,N_5074);
nand U6682 (N_6682,N_5198,N_5281);
xor U6683 (N_6683,N_5922,N_5588);
and U6684 (N_6684,N_5066,N_5491);
nand U6685 (N_6685,N_5264,N_5492);
and U6686 (N_6686,N_5957,N_5972);
or U6687 (N_6687,N_5448,N_5381);
nor U6688 (N_6688,N_5953,N_5803);
and U6689 (N_6689,N_5813,N_5947);
nor U6690 (N_6690,N_5488,N_5362);
nand U6691 (N_6691,N_5937,N_5501);
nand U6692 (N_6692,N_5023,N_5463);
nor U6693 (N_6693,N_5481,N_5614);
nand U6694 (N_6694,N_5265,N_5250);
or U6695 (N_6695,N_5381,N_5203);
nor U6696 (N_6696,N_5338,N_5104);
nor U6697 (N_6697,N_5293,N_5621);
and U6698 (N_6698,N_5051,N_5350);
or U6699 (N_6699,N_5308,N_5217);
and U6700 (N_6700,N_5076,N_5618);
and U6701 (N_6701,N_5927,N_5036);
nand U6702 (N_6702,N_5036,N_5303);
nor U6703 (N_6703,N_5527,N_5118);
or U6704 (N_6704,N_5670,N_5721);
nand U6705 (N_6705,N_5843,N_5637);
nor U6706 (N_6706,N_5473,N_5305);
nor U6707 (N_6707,N_5507,N_5086);
or U6708 (N_6708,N_5505,N_5216);
or U6709 (N_6709,N_5926,N_5696);
and U6710 (N_6710,N_5096,N_5551);
nand U6711 (N_6711,N_5773,N_5959);
nand U6712 (N_6712,N_5849,N_5851);
and U6713 (N_6713,N_5931,N_5196);
xnor U6714 (N_6714,N_5405,N_5433);
and U6715 (N_6715,N_5289,N_5297);
nor U6716 (N_6716,N_5567,N_5232);
nand U6717 (N_6717,N_5569,N_5230);
nor U6718 (N_6718,N_5928,N_5192);
xnor U6719 (N_6719,N_5641,N_5647);
nor U6720 (N_6720,N_5989,N_5290);
or U6721 (N_6721,N_5230,N_5160);
or U6722 (N_6722,N_5718,N_5682);
nand U6723 (N_6723,N_5314,N_5527);
nor U6724 (N_6724,N_5530,N_5346);
and U6725 (N_6725,N_5244,N_5646);
or U6726 (N_6726,N_5770,N_5076);
and U6727 (N_6727,N_5002,N_5861);
and U6728 (N_6728,N_5664,N_5650);
nand U6729 (N_6729,N_5561,N_5516);
nor U6730 (N_6730,N_5429,N_5186);
and U6731 (N_6731,N_5384,N_5827);
nor U6732 (N_6732,N_5795,N_5271);
nand U6733 (N_6733,N_5057,N_5126);
or U6734 (N_6734,N_5013,N_5627);
nor U6735 (N_6735,N_5029,N_5009);
and U6736 (N_6736,N_5542,N_5968);
nor U6737 (N_6737,N_5320,N_5294);
nor U6738 (N_6738,N_5435,N_5768);
nor U6739 (N_6739,N_5367,N_5474);
or U6740 (N_6740,N_5589,N_5571);
or U6741 (N_6741,N_5269,N_5411);
and U6742 (N_6742,N_5636,N_5640);
or U6743 (N_6743,N_5172,N_5241);
and U6744 (N_6744,N_5446,N_5314);
or U6745 (N_6745,N_5201,N_5504);
nor U6746 (N_6746,N_5308,N_5837);
nand U6747 (N_6747,N_5742,N_5587);
nor U6748 (N_6748,N_5268,N_5862);
nand U6749 (N_6749,N_5461,N_5707);
and U6750 (N_6750,N_5331,N_5798);
or U6751 (N_6751,N_5045,N_5919);
nor U6752 (N_6752,N_5278,N_5868);
and U6753 (N_6753,N_5558,N_5567);
or U6754 (N_6754,N_5177,N_5831);
or U6755 (N_6755,N_5164,N_5173);
nand U6756 (N_6756,N_5095,N_5252);
or U6757 (N_6757,N_5116,N_5328);
nor U6758 (N_6758,N_5932,N_5572);
nor U6759 (N_6759,N_5429,N_5754);
or U6760 (N_6760,N_5851,N_5199);
and U6761 (N_6761,N_5790,N_5611);
and U6762 (N_6762,N_5978,N_5494);
nand U6763 (N_6763,N_5600,N_5447);
or U6764 (N_6764,N_5934,N_5267);
nand U6765 (N_6765,N_5668,N_5264);
or U6766 (N_6766,N_5173,N_5097);
nor U6767 (N_6767,N_5279,N_5305);
and U6768 (N_6768,N_5267,N_5285);
nand U6769 (N_6769,N_5961,N_5999);
nor U6770 (N_6770,N_5282,N_5493);
and U6771 (N_6771,N_5456,N_5301);
and U6772 (N_6772,N_5861,N_5145);
nand U6773 (N_6773,N_5144,N_5837);
and U6774 (N_6774,N_5585,N_5150);
or U6775 (N_6775,N_5994,N_5549);
or U6776 (N_6776,N_5506,N_5884);
nand U6777 (N_6777,N_5168,N_5988);
nor U6778 (N_6778,N_5361,N_5037);
nand U6779 (N_6779,N_5176,N_5562);
nand U6780 (N_6780,N_5728,N_5703);
nor U6781 (N_6781,N_5687,N_5680);
or U6782 (N_6782,N_5249,N_5645);
and U6783 (N_6783,N_5372,N_5030);
nor U6784 (N_6784,N_5704,N_5538);
nand U6785 (N_6785,N_5193,N_5208);
nor U6786 (N_6786,N_5002,N_5094);
nor U6787 (N_6787,N_5116,N_5082);
and U6788 (N_6788,N_5611,N_5952);
and U6789 (N_6789,N_5179,N_5876);
and U6790 (N_6790,N_5137,N_5974);
or U6791 (N_6791,N_5091,N_5881);
nor U6792 (N_6792,N_5220,N_5305);
nor U6793 (N_6793,N_5620,N_5661);
nand U6794 (N_6794,N_5559,N_5398);
nand U6795 (N_6795,N_5499,N_5400);
or U6796 (N_6796,N_5672,N_5486);
or U6797 (N_6797,N_5516,N_5188);
nand U6798 (N_6798,N_5031,N_5501);
nor U6799 (N_6799,N_5704,N_5304);
or U6800 (N_6800,N_5802,N_5730);
or U6801 (N_6801,N_5724,N_5617);
nor U6802 (N_6802,N_5284,N_5818);
nor U6803 (N_6803,N_5335,N_5495);
nand U6804 (N_6804,N_5699,N_5764);
or U6805 (N_6805,N_5291,N_5779);
nand U6806 (N_6806,N_5818,N_5791);
nand U6807 (N_6807,N_5103,N_5084);
nand U6808 (N_6808,N_5442,N_5876);
and U6809 (N_6809,N_5085,N_5121);
nor U6810 (N_6810,N_5106,N_5454);
and U6811 (N_6811,N_5458,N_5738);
or U6812 (N_6812,N_5790,N_5842);
or U6813 (N_6813,N_5629,N_5886);
or U6814 (N_6814,N_5009,N_5921);
nor U6815 (N_6815,N_5365,N_5575);
or U6816 (N_6816,N_5767,N_5861);
nand U6817 (N_6817,N_5537,N_5189);
nor U6818 (N_6818,N_5213,N_5645);
or U6819 (N_6819,N_5651,N_5406);
nor U6820 (N_6820,N_5495,N_5500);
or U6821 (N_6821,N_5389,N_5831);
nor U6822 (N_6822,N_5046,N_5388);
or U6823 (N_6823,N_5516,N_5443);
nand U6824 (N_6824,N_5701,N_5254);
and U6825 (N_6825,N_5267,N_5295);
nor U6826 (N_6826,N_5044,N_5243);
nor U6827 (N_6827,N_5142,N_5073);
nor U6828 (N_6828,N_5694,N_5350);
and U6829 (N_6829,N_5103,N_5581);
nor U6830 (N_6830,N_5909,N_5971);
and U6831 (N_6831,N_5192,N_5283);
and U6832 (N_6832,N_5583,N_5159);
nor U6833 (N_6833,N_5001,N_5603);
or U6834 (N_6834,N_5995,N_5400);
or U6835 (N_6835,N_5910,N_5902);
and U6836 (N_6836,N_5358,N_5437);
nand U6837 (N_6837,N_5188,N_5814);
nor U6838 (N_6838,N_5228,N_5560);
nand U6839 (N_6839,N_5562,N_5294);
nor U6840 (N_6840,N_5636,N_5425);
nor U6841 (N_6841,N_5121,N_5880);
nand U6842 (N_6842,N_5054,N_5418);
or U6843 (N_6843,N_5149,N_5673);
nand U6844 (N_6844,N_5811,N_5663);
nor U6845 (N_6845,N_5961,N_5125);
nor U6846 (N_6846,N_5849,N_5471);
nor U6847 (N_6847,N_5930,N_5804);
and U6848 (N_6848,N_5044,N_5011);
and U6849 (N_6849,N_5536,N_5183);
or U6850 (N_6850,N_5936,N_5622);
and U6851 (N_6851,N_5390,N_5481);
or U6852 (N_6852,N_5647,N_5098);
or U6853 (N_6853,N_5196,N_5609);
or U6854 (N_6854,N_5095,N_5475);
or U6855 (N_6855,N_5235,N_5268);
nand U6856 (N_6856,N_5393,N_5150);
and U6857 (N_6857,N_5588,N_5245);
nor U6858 (N_6858,N_5317,N_5873);
nand U6859 (N_6859,N_5493,N_5834);
and U6860 (N_6860,N_5400,N_5438);
or U6861 (N_6861,N_5781,N_5080);
and U6862 (N_6862,N_5589,N_5361);
and U6863 (N_6863,N_5190,N_5524);
and U6864 (N_6864,N_5023,N_5488);
nand U6865 (N_6865,N_5724,N_5702);
and U6866 (N_6866,N_5750,N_5026);
and U6867 (N_6867,N_5039,N_5163);
and U6868 (N_6868,N_5814,N_5175);
nand U6869 (N_6869,N_5663,N_5070);
nand U6870 (N_6870,N_5357,N_5439);
and U6871 (N_6871,N_5669,N_5861);
and U6872 (N_6872,N_5512,N_5154);
nand U6873 (N_6873,N_5189,N_5518);
and U6874 (N_6874,N_5439,N_5652);
nand U6875 (N_6875,N_5828,N_5488);
nor U6876 (N_6876,N_5003,N_5678);
and U6877 (N_6877,N_5779,N_5232);
or U6878 (N_6878,N_5341,N_5078);
nor U6879 (N_6879,N_5904,N_5894);
or U6880 (N_6880,N_5396,N_5513);
nand U6881 (N_6881,N_5801,N_5580);
nand U6882 (N_6882,N_5696,N_5409);
nor U6883 (N_6883,N_5738,N_5715);
or U6884 (N_6884,N_5662,N_5523);
nor U6885 (N_6885,N_5285,N_5088);
or U6886 (N_6886,N_5095,N_5452);
and U6887 (N_6887,N_5033,N_5041);
or U6888 (N_6888,N_5969,N_5055);
or U6889 (N_6889,N_5322,N_5268);
and U6890 (N_6890,N_5433,N_5766);
nor U6891 (N_6891,N_5976,N_5005);
nor U6892 (N_6892,N_5867,N_5438);
nand U6893 (N_6893,N_5169,N_5549);
nand U6894 (N_6894,N_5650,N_5165);
nor U6895 (N_6895,N_5253,N_5304);
and U6896 (N_6896,N_5595,N_5575);
nor U6897 (N_6897,N_5848,N_5793);
nand U6898 (N_6898,N_5619,N_5029);
or U6899 (N_6899,N_5423,N_5945);
or U6900 (N_6900,N_5001,N_5254);
or U6901 (N_6901,N_5541,N_5259);
nor U6902 (N_6902,N_5747,N_5002);
nand U6903 (N_6903,N_5397,N_5211);
nand U6904 (N_6904,N_5002,N_5634);
and U6905 (N_6905,N_5387,N_5053);
nand U6906 (N_6906,N_5055,N_5636);
and U6907 (N_6907,N_5620,N_5917);
nor U6908 (N_6908,N_5243,N_5407);
and U6909 (N_6909,N_5283,N_5230);
xor U6910 (N_6910,N_5784,N_5053);
nor U6911 (N_6911,N_5556,N_5242);
nor U6912 (N_6912,N_5240,N_5034);
and U6913 (N_6913,N_5181,N_5353);
or U6914 (N_6914,N_5585,N_5912);
or U6915 (N_6915,N_5784,N_5458);
or U6916 (N_6916,N_5219,N_5251);
nand U6917 (N_6917,N_5604,N_5092);
nand U6918 (N_6918,N_5743,N_5219);
or U6919 (N_6919,N_5404,N_5758);
and U6920 (N_6920,N_5503,N_5630);
nor U6921 (N_6921,N_5997,N_5244);
nand U6922 (N_6922,N_5389,N_5948);
and U6923 (N_6923,N_5639,N_5751);
or U6924 (N_6924,N_5736,N_5310);
nand U6925 (N_6925,N_5695,N_5225);
and U6926 (N_6926,N_5980,N_5758);
xor U6927 (N_6927,N_5745,N_5285);
and U6928 (N_6928,N_5491,N_5309);
nand U6929 (N_6929,N_5895,N_5687);
nor U6930 (N_6930,N_5541,N_5332);
or U6931 (N_6931,N_5632,N_5244);
nor U6932 (N_6932,N_5254,N_5268);
nor U6933 (N_6933,N_5271,N_5416);
and U6934 (N_6934,N_5715,N_5300);
and U6935 (N_6935,N_5804,N_5107);
nand U6936 (N_6936,N_5063,N_5760);
nor U6937 (N_6937,N_5390,N_5901);
and U6938 (N_6938,N_5863,N_5959);
or U6939 (N_6939,N_5441,N_5032);
nand U6940 (N_6940,N_5881,N_5612);
nand U6941 (N_6941,N_5978,N_5161);
nor U6942 (N_6942,N_5286,N_5555);
nor U6943 (N_6943,N_5283,N_5361);
nor U6944 (N_6944,N_5746,N_5156);
nor U6945 (N_6945,N_5512,N_5437);
nor U6946 (N_6946,N_5780,N_5774);
or U6947 (N_6947,N_5045,N_5617);
nand U6948 (N_6948,N_5510,N_5515);
or U6949 (N_6949,N_5384,N_5091);
nand U6950 (N_6950,N_5460,N_5130);
and U6951 (N_6951,N_5752,N_5461);
or U6952 (N_6952,N_5085,N_5901);
and U6953 (N_6953,N_5298,N_5501);
nor U6954 (N_6954,N_5117,N_5180);
and U6955 (N_6955,N_5705,N_5822);
and U6956 (N_6956,N_5608,N_5674);
or U6957 (N_6957,N_5274,N_5885);
nor U6958 (N_6958,N_5855,N_5535);
nand U6959 (N_6959,N_5312,N_5219);
nand U6960 (N_6960,N_5579,N_5373);
and U6961 (N_6961,N_5891,N_5216);
and U6962 (N_6962,N_5908,N_5764);
or U6963 (N_6963,N_5280,N_5029);
or U6964 (N_6964,N_5241,N_5091);
nor U6965 (N_6965,N_5375,N_5311);
nor U6966 (N_6966,N_5415,N_5422);
nor U6967 (N_6967,N_5286,N_5471);
nand U6968 (N_6968,N_5261,N_5717);
and U6969 (N_6969,N_5726,N_5982);
nand U6970 (N_6970,N_5943,N_5185);
nor U6971 (N_6971,N_5562,N_5161);
and U6972 (N_6972,N_5095,N_5396);
nand U6973 (N_6973,N_5718,N_5373);
and U6974 (N_6974,N_5271,N_5067);
nor U6975 (N_6975,N_5125,N_5381);
nand U6976 (N_6976,N_5127,N_5895);
nand U6977 (N_6977,N_5080,N_5722);
nand U6978 (N_6978,N_5596,N_5516);
and U6979 (N_6979,N_5604,N_5831);
or U6980 (N_6980,N_5998,N_5542);
and U6981 (N_6981,N_5800,N_5941);
or U6982 (N_6982,N_5326,N_5554);
and U6983 (N_6983,N_5827,N_5831);
and U6984 (N_6984,N_5658,N_5730);
nand U6985 (N_6985,N_5939,N_5270);
or U6986 (N_6986,N_5557,N_5648);
and U6987 (N_6987,N_5267,N_5962);
nor U6988 (N_6988,N_5692,N_5715);
nor U6989 (N_6989,N_5475,N_5750);
nand U6990 (N_6990,N_5128,N_5135);
or U6991 (N_6991,N_5783,N_5420);
or U6992 (N_6992,N_5254,N_5703);
and U6993 (N_6993,N_5573,N_5356);
and U6994 (N_6994,N_5692,N_5560);
nand U6995 (N_6995,N_5871,N_5141);
or U6996 (N_6996,N_5471,N_5762);
or U6997 (N_6997,N_5969,N_5505);
or U6998 (N_6998,N_5867,N_5682);
or U6999 (N_6999,N_5693,N_5050);
and U7000 (N_7000,N_6050,N_6914);
and U7001 (N_7001,N_6351,N_6236);
and U7002 (N_7002,N_6712,N_6445);
and U7003 (N_7003,N_6450,N_6662);
or U7004 (N_7004,N_6287,N_6444);
and U7005 (N_7005,N_6280,N_6491);
or U7006 (N_7006,N_6763,N_6912);
and U7007 (N_7007,N_6126,N_6362);
nand U7008 (N_7008,N_6890,N_6334);
or U7009 (N_7009,N_6277,N_6627);
nor U7010 (N_7010,N_6558,N_6534);
and U7011 (N_7011,N_6609,N_6123);
nor U7012 (N_7012,N_6632,N_6971);
or U7013 (N_7013,N_6306,N_6898);
nor U7014 (N_7014,N_6350,N_6948);
or U7015 (N_7015,N_6607,N_6060);
and U7016 (N_7016,N_6008,N_6330);
and U7017 (N_7017,N_6440,N_6465);
nand U7018 (N_7018,N_6459,N_6839);
nor U7019 (N_7019,N_6166,N_6681);
or U7020 (N_7020,N_6376,N_6652);
and U7021 (N_7021,N_6421,N_6292);
nor U7022 (N_7022,N_6992,N_6457);
nand U7023 (N_7023,N_6909,N_6594);
and U7024 (N_7024,N_6071,N_6380);
nand U7025 (N_7025,N_6369,N_6253);
nand U7026 (N_7026,N_6731,N_6694);
xnor U7027 (N_7027,N_6503,N_6939);
nor U7028 (N_7028,N_6677,N_6392);
nand U7029 (N_7029,N_6065,N_6022);
or U7030 (N_7030,N_6642,N_6940);
or U7031 (N_7031,N_6276,N_6713);
nand U7032 (N_7032,N_6499,N_6629);
and U7033 (N_7033,N_6090,N_6747);
and U7034 (N_7034,N_6782,N_6106);
xor U7035 (N_7035,N_6838,N_6866);
nor U7036 (N_7036,N_6266,N_6606);
nor U7037 (N_7037,N_6162,N_6476);
or U7038 (N_7038,N_6477,N_6025);
and U7039 (N_7039,N_6099,N_6636);
or U7040 (N_7040,N_6219,N_6274);
nand U7041 (N_7041,N_6846,N_6682);
nor U7042 (N_7042,N_6989,N_6107);
nand U7043 (N_7043,N_6868,N_6547);
or U7044 (N_7044,N_6225,N_6251);
and U7045 (N_7045,N_6168,N_6278);
or U7046 (N_7046,N_6834,N_6617);
nor U7047 (N_7047,N_6339,N_6319);
nor U7048 (N_7048,N_6341,N_6395);
nor U7049 (N_7049,N_6044,N_6064);
or U7050 (N_7050,N_6808,N_6154);
nand U7051 (N_7051,N_6938,N_6415);
or U7052 (N_7052,N_6686,N_6066);
or U7053 (N_7053,N_6222,N_6869);
and U7054 (N_7054,N_6772,N_6147);
nand U7055 (N_7055,N_6699,N_6180);
nand U7056 (N_7056,N_6666,N_6347);
and U7057 (N_7057,N_6411,N_6618);
nor U7058 (N_7058,N_6551,N_6344);
nand U7059 (N_7059,N_6608,N_6245);
and U7060 (N_7060,N_6806,N_6860);
nor U7061 (N_7061,N_6779,N_6648);
and U7062 (N_7062,N_6069,N_6270);
nand U7063 (N_7063,N_6286,N_6628);
nor U7064 (N_7064,N_6532,N_6078);
nand U7065 (N_7065,N_6262,N_6368);
or U7066 (N_7066,N_6439,N_6730);
nor U7067 (N_7067,N_6661,N_6974);
nand U7068 (N_7068,N_6564,N_6824);
nor U7069 (N_7069,N_6113,N_6563);
and U7070 (N_7070,N_6055,N_6175);
or U7071 (N_7071,N_6208,N_6619);
and U7072 (N_7072,N_6098,N_6934);
nand U7073 (N_7073,N_6058,N_6000);
and U7074 (N_7074,N_6194,N_6364);
nor U7075 (N_7075,N_6494,N_6927);
or U7076 (N_7076,N_6588,N_6878);
nor U7077 (N_7077,N_6358,N_6247);
or U7078 (N_7078,N_6237,N_6333);
nand U7079 (N_7079,N_6798,N_6243);
and U7080 (N_7080,N_6343,N_6036);
nor U7081 (N_7081,N_6216,N_6349);
nor U7082 (N_7082,N_6472,N_6031);
or U7083 (N_7083,N_6037,N_6488);
nor U7084 (N_7084,N_6127,N_6186);
or U7085 (N_7085,N_6603,N_6765);
and U7086 (N_7086,N_6794,N_6626);
nand U7087 (N_7087,N_6674,N_6787);
and U7088 (N_7088,N_6651,N_6665);
and U7089 (N_7089,N_6087,N_6531);
nor U7090 (N_7090,N_6998,N_6524);
nand U7091 (N_7091,N_6972,N_6460);
and U7092 (N_7092,N_6903,N_6643);
nand U7093 (N_7093,N_6673,N_6224);
or U7094 (N_7094,N_6508,N_6924);
and U7095 (N_7095,N_6359,N_6384);
nor U7096 (N_7096,N_6889,N_6511);
or U7097 (N_7097,N_6595,N_6057);
nor U7098 (N_7098,N_6404,N_6758);
xnor U7099 (N_7099,N_6049,N_6110);
or U7100 (N_7100,N_6767,N_6146);
nor U7101 (N_7101,N_6386,N_6716);
or U7102 (N_7102,N_6602,N_6176);
and U7103 (N_7103,N_6032,N_6814);
nand U7104 (N_7104,N_6610,N_6611);
nor U7105 (N_7105,N_6111,N_6753);
nor U7106 (N_7106,N_6843,N_6314);
nor U7107 (N_7107,N_6810,N_6687);
or U7108 (N_7108,N_6461,N_6128);
or U7109 (N_7109,N_6539,N_6373);
nand U7110 (N_7110,N_6235,N_6800);
or U7111 (N_7111,N_6118,N_6062);
nor U7112 (N_7112,N_6009,N_6668);
nand U7113 (N_7113,N_6275,N_6002);
and U7114 (N_7114,N_6569,N_6560);
or U7115 (N_7115,N_6954,N_6396);
nand U7116 (N_7116,N_6294,N_6596);
nor U7117 (N_7117,N_6452,N_6883);
and U7118 (N_7118,N_6536,N_6256);
nand U7119 (N_7119,N_6947,N_6241);
nor U7120 (N_7120,N_6300,N_6574);
and U7121 (N_7121,N_6955,N_6737);
and U7122 (N_7122,N_6148,N_6473);
or U7123 (N_7123,N_6298,N_6749);
nand U7124 (N_7124,N_6407,N_6259);
or U7125 (N_7125,N_6131,N_6430);
nor U7126 (N_7126,N_6405,N_6268);
nor U7127 (N_7127,N_6984,N_6733);
nor U7128 (N_7128,N_6248,N_6114);
and U7129 (N_7129,N_6513,N_6289);
nand U7130 (N_7130,N_6638,N_6310);
nor U7131 (N_7131,N_6757,N_6891);
nand U7132 (N_7132,N_6422,N_6074);
nand U7133 (N_7133,N_6550,N_6802);
nor U7134 (N_7134,N_6512,N_6052);
nand U7135 (N_7135,N_6228,N_6134);
nand U7136 (N_7136,N_6902,N_6656);
nand U7137 (N_7137,N_6417,N_6320);
xnor U7138 (N_7138,N_6023,N_6322);
or U7139 (N_7139,N_6719,N_6188);
and U7140 (N_7140,N_6139,N_6410);
or U7141 (N_7141,N_6826,N_6211);
and U7142 (N_7142,N_6515,N_6791);
xor U7143 (N_7143,N_6479,N_6013);
nor U7144 (N_7144,N_6095,N_6529);
and U7145 (N_7145,N_6635,N_6621);
or U7146 (N_7146,N_6953,N_6988);
nand U7147 (N_7147,N_6130,N_6525);
nand U7148 (N_7148,N_6841,N_6109);
nor U7149 (N_7149,N_6658,N_6520);
or U7150 (N_7150,N_6073,N_6004);
and U7151 (N_7151,N_6283,N_6068);
xor U7152 (N_7152,N_6246,N_6296);
nor U7153 (N_7153,N_6318,N_6533);
and U7154 (N_7154,N_6137,N_6391);
or U7155 (N_7155,N_6279,N_6418);
and U7156 (N_7156,N_6119,N_6209);
and U7157 (N_7157,N_6329,N_6084);
or U7158 (N_7158,N_6385,N_6640);
nor U7159 (N_7159,N_6093,N_6398);
or U7160 (N_7160,N_6762,N_6401);
or U7161 (N_7161,N_6876,N_6977);
nand U7162 (N_7162,N_6892,N_6535);
or U7163 (N_7163,N_6746,N_6414);
or U7164 (N_7164,N_6675,N_6260);
nor U7165 (N_7165,N_6580,N_6230);
nor U7166 (N_7166,N_6102,N_6265);
or U7167 (N_7167,N_6945,N_6865);
nand U7168 (N_7168,N_6308,N_6654);
and U7169 (N_7169,N_6432,N_6389);
nand U7170 (N_7170,N_6167,N_6683);
or U7171 (N_7171,N_6703,N_6151);
nor U7172 (N_7172,N_6173,N_6768);
and U7173 (N_7173,N_6925,N_6797);
nor U7174 (N_7174,N_6734,N_6101);
nor U7175 (N_7175,N_6647,N_6129);
nand U7176 (N_7176,N_6043,N_6233);
nand U7177 (N_7177,N_6091,N_6079);
nand U7178 (N_7178,N_6135,N_6795);
nand U7179 (N_7179,N_6553,N_6807);
nor U7180 (N_7180,N_6014,N_6848);
or U7181 (N_7181,N_6943,N_6773);
and U7182 (N_7182,N_6993,N_6315);
nor U7183 (N_7183,N_6451,N_6234);
nor U7184 (N_7184,N_6759,N_6083);
and U7185 (N_7185,N_6475,N_6170);
and U7186 (N_7186,N_6307,N_6431);
nand U7187 (N_7187,N_6498,N_6593);
or U7188 (N_7188,N_6631,N_6849);
nand U7189 (N_7189,N_6586,N_6141);
nand U7190 (N_7190,N_6156,N_6874);
nor U7191 (N_7191,N_6336,N_6152);
xnor U7192 (N_7192,N_6840,N_6738);
nor U7193 (N_7193,N_6867,N_6979);
or U7194 (N_7194,N_6342,N_6847);
nor U7195 (N_7195,N_6990,N_6858);
or U7196 (N_7196,N_6124,N_6736);
nor U7197 (N_7197,N_6149,N_6966);
and U7198 (N_7198,N_6671,N_6337);
nor U7199 (N_7199,N_6695,N_6857);
and U7200 (N_7200,N_6326,N_6830);
and U7201 (N_7201,N_6446,N_6669);
or U7202 (N_7202,N_6663,N_6585);
or U7203 (N_7203,N_6420,N_6781);
nand U7204 (N_7204,N_6873,N_6197);
nand U7205 (N_7205,N_6983,N_6899);
nor U7206 (N_7206,N_6360,N_6375);
or U7207 (N_7207,N_6085,N_6232);
nand U7208 (N_7208,N_6624,N_6584);
nand U7209 (N_7209,N_6252,N_6783);
nand U7210 (N_7210,N_6548,N_6557);
and U7211 (N_7211,N_6182,N_6019);
nand U7212 (N_7212,N_6922,N_6157);
nor U7213 (N_7213,N_6742,N_6698);
or U7214 (N_7214,N_6937,N_6637);
or U7215 (N_7215,N_6143,N_6901);
nor U7216 (N_7216,N_6115,N_6855);
and U7217 (N_7217,N_6076,N_6426);
nor U7218 (N_7218,N_6469,N_6965);
or U7219 (N_7219,N_6448,N_6996);
or U7220 (N_7220,N_6579,N_6519);
nand U7221 (N_7221,N_6975,N_6710);
nand U7222 (N_7222,N_6893,N_6213);
and U7223 (N_7223,N_6701,N_6165);
nor U7224 (N_7224,N_6919,N_6449);
and U7225 (N_7225,N_6163,N_6641);
and U7226 (N_7226,N_6054,N_6726);
nor U7227 (N_7227,N_6527,N_6545);
nand U7228 (N_7228,N_6960,N_6961);
nor U7229 (N_7229,N_6203,N_6456);
nand U7230 (N_7230,N_6305,N_6017);
and U7231 (N_7231,N_6220,N_6325);
nor U7232 (N_7232,N_6721,N_6041);
and U7233 (N_7233,N_6946,N_6010);
and U7234 (N_7234,N_6311,N_6549);
or U7235 (N_7235,N_6835,N_6026);
nand U7236 (N_7236,N_6427,N_6523);
and U7237 (N_7237,N_6577,N_6623);
or U7238 (N_7238,N_6309,N_6223);
and U7239 (N_7239,N_6226,N_6021);
nor U7240 (N_7240,N_6755,N_6600);
and U7241 (N_7241,N_6951,N_6818);
and U7242 (N_7242,N_6861,N_6863);
nor U7243 (N_7243,N_6471,N_6291);
nor U7244 (N_7244,N_6994,N_6900);
and U7245 (N_7245,N_6702,N_6438);
nor U7246 (N_7246,N_6212,N_6056);
or U7247 (N_7247,N_6504,N_6122);
nand U7248 (N_7248,N_6505,N_6756);
or U7249 (N_7249,N_6406,N_6896);
and U7250 (N_7250,N_6985,N_6352);
and U7251 (N_7251,N_6785,N_6968);
nand U7252 (N_7252,N_6086,N_6813);
or U7253 (N_7253,N_6480,N_6601);
and U7254 (N_7254,N_6112,N_6644);
and U7255 (N_7255,N_6443,N_6387);
and U7256 (N_7256,N_6917,N_6562);
nand U7257 (N_7257,N_6987,N_6633);
nand U7258 (N_7258,N_6447,N_6764);
nand U7259 (N_7259,N_6192,N_6711);
nor U7260 (N_7260,N_6048,N_6895);
xnor U7261 (N_7261,N_6489,N_6751);
nand U7262 (N_7262,N_6363,N_6852);
and U7263 (N_7263,N_6837,N_6374);
or U7264 (N_7264,N_6778,N_6522);
or U7265 (N_7265,N_6770,N_6853);
nor U7266 (N_7266,N_6024,N_6361);
nand U7267 (N_7267,N_6178,N_6570);
or U7268 (N_7268,N_6543,N_6214);
nand U7269 (N_7269,N_6189,N_6027);
or U7270 (N_7270,N_6200,N_6850);
nor U7271 (N_7271,N_6991,N_6070);
or U7272 (N_7272,N_6670,N_6202);
nand U7273 (N_7273,N_6204,N_6346);
nand U7274 (N_7274,N_6103,N_6589);
nand U7275 (N_7275,N_6664,N_6655);
nor U7276 (N_7276,N_6403,N_6267);
and U7277 (N_7277,N_6293,N_6717);
and U7278 (N_7278,N_6348,N_6120);
nand U7279 (N_7279,N_6567,N_6317);
and U7280 (N_7280,N_6018,N_6383);
nand U7281 (N_7281,N_6958,N_6038);
or U7282 (N_7282,N_6910,N_6572);
or U7283 (N_7283,N_6784,N_6371);
nor U7284 (N_7284,N_6367,N_6776);
nand U7285 (N_7285,N_6474,N_6382);
or U7286 (N_7286,N_6132,N_6125);
or U7287 (N_7287,N_6169,N_6541);
or U7288 (N_7288,N_6051,N_6831);
nor U7289 (N_7289,N_6324,N_6566);
and U7290 (N_7290,N_6497,N_6003);
nand U7291 (N_7291,N_6911,N_6517);
nor U7292 (N_7292,N_6882,N_6419);
or U7293 (N_7293,N_6886,N_6506);
nand U7294 (N_7294,N_6879,N_6926);
nand U7295 (N_7295,N_6880,N_6905);
nand U7296 (N_7296,N_6035,N_6752);
or U7297 (N_7297,N_6016,N_6928);
nand U7298 (N_7298,N_6030,N_6918);
nor U7299 (N_7299,N_6257,N_6780);
nand U7300 (N_7300,N_6487,N_6138);
nor U7301 (N_7301,N_6205,N_6575);
and U7302 (N_7302,N_6201,N_6179);
and U7303 (N_7303,N_6583,N_6526);
nor U7304 (N_7304,N_6788,N_6851);
or U7305 (N_7305,N_6920,N_6423);
or U7306 (N_7306,N_6705,N_6184);
or U7307 (N_7307,N_6092,N_6433);
nand U7308 (N_7308,N_6412,N_6366);
and U7309 (N_7309,N_6613,N_6425);
nand U7310 (N_7310,N_6356,N_6254);
nor U7311 (N_7311,N_6552,N_6281);
nand U7312 (N_7312,N_6587,N_6875);
or U7313 (N_7313,N_6688,N_6650);
or U7314 (N_7314,N_6081,N_6728);
nand U7315 (N_7315,N_6240,N_6789);
nor U7316 (N_7316,N_6832,N_6842);
and U7317 (N_7317,N_6921,N_6015);
nand U7318 (N_7318,N_6836,N_6136);
and U7319 (N_7319,N_6769,N_6484);
or U7320 (N_7320,N_6088,N_6408);
nor U7321 (N_7321,N_6269,N_6709);
nand U7322 (N_7322,N_6250,N_6967);
nand U7323 (N_7323,N_6142,N_6510);
nor U7324 (N_7324,N_6727,N_6261);
and U7325 (N_7325,N_6718,N_6799);
nor U7326 (N_7326,N_6931,N_6409);
nor U7327 (N_7327,N_6884,N_6273);
or U7328 (N_7328,N_6416,N_6227);
and U7329 (N_7329,N_6685,N_6316);
and U7330 (N_7330,N_6105,N_6462);
and U7331 (N_7331,N_6862,N_6775);
or U7332 (N_7332,N_6754,N_6238);
and U7333 (N_7333,N_6028,N_6297);
nor U7334 (N_7334,N_6453,N_6321);
nor U7335 (N_7335,N_6434,N_6741);
and U7336 (N_7336,N_6328,N_6011);
nand U7337 (N_7337,N_6812,N_6518);
and U7338 (N_7338,N_6885,N_6521);
nand U7339 (N_7339,N_6725,N_6516);
nand U7340 (N_7340,N_6467,N_6485);
and U7341 (N_7341,N_6047,N_6748);
and U7342 (N_7342,N_6684,N_6133);
nand U7343 (N_7343,N_6906,N_6740);
and U7344 (N_7344,N_6001,N_6986);
and U7345 (N_7345,N_6242,N_6796);
or U7346 (N_7346,N_6973,N_6645);
or U7347 (N_7347,N_6962,N_6935);
and U7348 (N_7348,N_6819,N_6809);
or U7349 (N_7349,N_6229,N_6823);
or U7350 (N_7350,N_6793,N_6639);
or U7351 (N_7351,N_6581,N_6653);
or U7352 (N_7352,N_6957,N_6397);
or U7353 (N_7353,N_6706,N_6390);
and U7354 (N_7354,N_6537,N_6714);
and U7355 (N_7355,N_6303,N_6715);
nor U7356 (N_7356,N_6659,N_6394);
or U7357 (N_7357,N_6542,N_6501);
and U7358 (N_7358,N_6458,N_6302);
and U7359 (N_7359,N_6210,N_6221);
nor U7360 (N_7360,N_6486,N_6672);
nor U7361 (N_7361,N_6218,N_6496);
and U7362 (N_7362,N_6108,N_6887);
and U7363 (N_7363,N_6195,N_6591);
or U7364 (N_7364,N_6492,N_6495);
and U7365 (N_7365,N_6915,N_6944);
nor U7366 (N_7366,N_6046,N_6708);
nor U7367 (N_7367,N_6978,N_6620);
nand U7368 (N_7368,N_6100,N_6872);
and U7369 (N_7369,N_6556,N_6077);
nor U7370 (N_7370,N_6082,N_6455);
and U7371 (N_7371,N_6304,N_6722);
or U7372 (N_7372,N_6691,N_6288);
and U7373 (N_7373,N_6576,N_6833);
nor U7374 (N_7374,N_6590,N_6264);
and U7375 (N_7375,N_6956,N_6828);
and U7376 (N_7376,N_6161,N_6821);
and U7377 (N_7377,N_6206,N_6089);
nor U7378 (N_7378,N_6429,N_6777);
and U7379 (N_7379,N_6441,N_6059);
nor U7380 (N_7380,N_6676,N_6870);
or U7381 (N_7381,N_6454,N_6171);
and U7382 (N_7382,N_6554,N_6528);
and U7383 (N_7383,N_6153,N_6413);
nand U7384 (N_7384,N_6981,N_6437);
nand U7385 (N_7385,N_6094,N_6530);
and U7386 (N_7386,N_6555,N_6908);
or U7387 (N_7387,N_6963,N_6700);
nand U7388 (N_7388,N_6097,N_6739);
nand U7389 (N_7389,N_6193,N_6854);
nor U7390 (N_7390,N_6612,N_6428);
and U7391 (N_7391,N_6766,N_6158);
and U7392 (N_7392,N_6258,N_6816);
or U7393 (N_7393,N_6040,N_6331);
nor U7394 (N_7394,N_6822,N_6950);
or U7395 (N_7395,N_6774,N_6907);
nor U7396 (N_7396,N_6913,N_6970);
or U7397 (N_7397,N_6573,N_6544);
and U7398 (N_7398,N_6982,N_6215);
and U7399 (N_7399,N_6692,N_6941);
nand U7400 (N_7400,N_6817,N_6295);
nor U7401 (N_7401,N_6466,N_6952);
and U7402 (N_7402,N_6061,N_6402);
and U7403 (N_7403,N_6424,N_6743);
nor U7404 (N_7404,N_6546,N_6185);
and U7405 (N_7405,N_6117,N_6801);
nand U7406 (N_7406,N_6353,N_6263);
nand U7407 (N_7407,N_6357,N_6904);
or U7408 (N_7408,N_6159,N_6005);
and U7409 (N_7409,N_6290,N_6696);
nand U7410 (N_7410,N_6881,N_6845);
nand U7411 (N_7411,N_6284,N_6299);
nand U7412 (N_7412,N_6646,N_6969);
or U7413 (N_7413,N_6976,N_6355);
nor U7414 (N_7414,N_6856,N_6436);
or U7415 (N_7415,N_6072,N_6231);
and U7416 (N_7416,N_6599,N_6500);
nand U7417 (N_7417,N_6622,N_6400);
or U7418 (N_7418,N_6121,N_6075);
nor U7419 (N_7419,N_6592,N_6388);
or U7420 (N_7420,N_6929,N_6301);
and U7421 (N_7421,N_6478,N_6198);
or U7422 (N_7422,N_6140,N_6680);
or U7423 (N_7423,N_6916,N_6820);
and U7424 (N_7424,N_6803,N_6285);
and U7425 (N_7425,N_6657,N_6615);
and U7426 (N_7426,N_6244,N_6249);
or U7427 (N_7427,N_6463,N_6217);
nor U7428 (N_7428,N_6568,N_6354);
nor U7429 (N_7429,N_6155,N_6335);
and U7430 (N_7430,N_6464,N_6177);
or U7431 (N_7431,N_6729,N_6145);
or U7432 (N_7432,N_6704,N_6897);
and U7433 (N_7433,N_6172,N_6690);
nand U7434 (N_7434,N_6745,N_6045);
and U7435 (N_7435,N_6864,N_6482);
nand U7436 (N_7436,N_6693,N_6805);
nor U7437 (N_7437,N_6160,N_6399);
nand U7438 (N_7438,N_6490,N_6894);
or U7439 (N_7439,N_6630,N_6006);
or U7440 (N_7440,N_6559,N_6829);
nor U7441 (N_7441,N_6507,N_6538);
nor U7442 (N_7442,N_6678,N_6790);
nand U7443 (N_7443,N_6012,N_6034);
nor U7444 (N_7444,N_6340,N_6381);
nor U7445 (N_7445,N_6735,N_6604);
nor U7446 (N_7446,N_6199,N_6771);
nand U7447 (N_7447,N_6365,N_6689);
nand U7448 (N_7448,N_6183,N_6732);
nand U7449 (N_7449,N_6571,N_6605);
nor U7450 (N_7450,N_6080,N_6104);
nor U7451 (N_7451,N_6660,N_6697);
and U7452 (N_7452,N_6561,N_6029);
nand U7453 (N_7453,N_6514,N_6679);
and U7454 (N_7454,N_6493,N_6877);
nand U7455 (N_7455,N_6191,N_6063);
or U7456 (N_7456,N_6483,N_6811);
nand U7457 (N_7457,N_6667,N_6007);
nor U7458 (N_7458,N_6634,N_6207);
nor U7459 (N_7459,N_6844,N_6723);
nor U7460 (N_7460,N_6053,N_6942);
nand U7461 (N_7461,N_6936,N_6239);
or U7462 (N_7462,N_6370,N_6379);
or U7463 (N_7463,N_6792,N_6442);
or U7464 (N_7464,N_6190,N_6323);
and U7465 (N_7465,N_6804,N_6150);
nand U7466 (N_7466,N_6378,N_6096);
or U7467 (N_7467,N_6949,N_6871);
nor U7468 (N_7468,N_6313,N_6859);
or U7469 (N_7469,N_6598,N_6327);
nor U7470 (N_7470,N_6750,N_6930);
and U7471 (N_7471,N_6181,N_6980);
and U7472 (N_7472,N_6345,N_6272);
nor U7473 (N_7473,N_6707,N_6164);
and U7474 (N_7474,N_6720,N_6372);
nand U7475 (N_7475,N_6020,N_6597);
and U7476 (N_7476,N_6625,N_6312);
nand U7477 (N_7477,N_6338,N_6509);
nand U7478 (N_7478,N_6888,N_6724);
or U7479 (N_7479,N_6377,N_6827);
and U7480 (N_7480,N_6786,N_6582);
and U7481 (N_7481,N_6540,N_6964);
nor U7482 (N_7482,N_6761,N_6932);
and U7483 (N_7483,N_6760,N_6042);
or U7484 (N_7484,N_6481,N_6997);
nand U7485 (N_7485,N_6174,N_6933);
nor U7486 (N_7486,N_6196,N_6144);
nor U7487 (N_7487,N_6995,N_6502);
and U7488 (N_7488,N_6271,N_6470);
nand U7489 (N_7489,N_6825,N_6999);
and U7490 (N_7490,N_6039,N_6959);
nand U7491 (N_7491,N_6649,N_6744);
nand U7492 (N_7492,N_6815,N_6616);
nand U7493 (N_7493,N_6614,N_6255);
or U7494 (N_7494,N_6282,N_6332);
nand U7495 (N_7495,N_6187,N_6923);
and U7496 (N_7496,N_6116,N_6033);
nor U7497 (N_7497,N_6468,N_6578);
nor U7498 (N_7498,N_6393,N_6067);
nor U7499 (N_7499,N_6565,N_6435);
or U7500 (N_7500,N_6936,N_6927);
or U7501 (N_7501,N_6806,N_6055);
nand U7502 (N_7502,N_6928,N_6182);
nand U7503 (N_7503,N_6813,N_6922);
xnor U7504 (N_7504,N_6783,N_6382);
and U7505 (N_7505,N_6626,N_6139);
nor U7506 (N_7506,N_6147,N_6335);
and U7507 (N_7507,N_6356,N_6793);
nand U7508 (N_7508,N_6502,N_6080);
nor U7509 (N_7509,N_6670,N_6767);
and U7510 (N_7510,N_6564,N_6918);
nor U7511 (N_7511,N_6286,N_6478);
and U7512 (N_7512,N_6795,N_6918);
and U7513 (N_7513,N_6635,N_6231);
nand U7514 (N_7514,N_6274,N_6825);
nor U7515 (N_7515,N_6427,N_6104);
or U7516 (N_7516,N_6946,N_6228);
and U7517 (N_7517,N_6784,N_6212);
nand U7518 (N_7518,N_6821,N_6036);
nand U7519 (N_7519,N_6859,N_6408);
or U7520 (N_7520,N_6377,N_6992);
or U7521 (N_7521,N_6644,N_6117);
nor U7522 (N_7522,N_6346,N_6255);
nor U7523 (N_7523,N_6425,N_6188);
and U7524 (N_7524,N_6866,N_6082);
and U7525 (N_7525,N_6466,N_6431);
nor U7526 (N_7526,N_6893,N_6817);
or U7527 (N_7527,N_6910,N_6043);
nand U7528 (N_7528,N_6061,N_6290);
or U7529 (N_7529,N_6051,N_6588);
nand U7530 (N_7530,N_6628,N_6209);
and U7531 (N_7531,N_6867,N_6757);
nor U7532 (N_7532,N_6877,N_6412);
or U7533 (N_7533,N_6246,N_6392);
nor U7534 (N_7534,N_6069,N_6824);
nand U7535 (N_7535,N_6114,N_6325);
nor U7536 (N_7536,N_6646,N_6451);
or U7537 (N_7537,N_6949,N_6762);
nor U7538 (N_7538,N_6772,N_6150);
nand U7539 (N_7539,N_6479,N_6857);
or U7540 (N_7540,N_6317,N_6826);
nor U7541 (N_7541,N_6558,N_6259);
and U7542 (N_7542,N_6793,N_6477);
and U7543 (N_7543,N_6942,N_6574);
nor U7544 (N_7544,N_6111,N_6586);
or U7545 (N_7545,N_6860,N_6933);
and U7546 (N_7546,N_6359,N_6323);
or U7547 (N_7547,N_6135,N_6270);
and U7548 (N_7548,N_6534,N_6363);
and U7549 (N_7549,N_6086,N_6802);
and U7550 (N_7550,N_6315,N_6717);
or U7551 (N_7551,N_6303,N_6855);
or U7552 (N_7552,N_6229,N_6306);
nor U7553 (N_7553,N_6702,N_6069);
nor U7554 (N_7554,N_6559,N_6509);
nor U7555 (N_7555,N_6538,N_6377);
nor U7556 (N_7556,N_6159,N_6101);
nor U7557 (N_7557,N_6424,N_6174);
or U7558 (N_7558,N_6124,N_6931);
nand U7559 (N_7559,N_6843,N_6205);
nand U7560 (N_7560,N_6218,N_6535);
or U7561 (N_7561,N_6885,N_6883);
and U7562 (N_7562,N_6221,N_6028);
nand U7563 (N_7563,N_6487,N_6176);
nor U7564 (N_7564,N_6102,N_6692);
nand U7565 (N_7565,N_6098,N_6331);
or U7566 (N_7566,N_6246,N_6763);
or U7567 (N_7567,N_6454,N_6786);
nand U7568 (N_7568,N_6853,N_6921);
or U7569 (N_7569,N_6861,N_6199);
or U7570 (N_7570,N_6938,N_6054);
and U7571 (N_7571,N_6852,N_6549);
and U7572 (N_7572,N_6625,N_6259);
nor U7573 (N_7573,N_6425,N_6455);
or U7574 (N_7574,N_6309,N_6803);
and U7575 (N_7575,N_6195,N_6612);
nand U7576 (N_7576,N_6439,N_6810);
and U7577 (N_7577,N_6386,N_6461);
nand U7578 (N_7578,N_6913,N_6844);
and U7579 (N_7579,N_6840,N_6051);
nand U7580 (N_7580,N_6303,N_6880);
nand U7581 (N_7581,N_6749,N_6777);
nand U7582 (N_7582,N_6967,N_6477);
or U7583 (N_7583,N_6461,N_6905);
nor U7584 (N_7584,N_6776,N_6162);
nand U7585 (N_7585,N_6837,N_6327);
and U7586 (N_7586,N_6432,N_6456);
or U7587 (N_7587,N_6348,N_6729);
and U7588 (N_7588,N_6749,N_6517);
and U7589 (N_7589,N_6301,N_6894);
nor U7590 (N_7590,N_6594,N_6917);
or U7591 (N_7591,N_6048,N_6995);
or U7592 (N_7592,N_6528,N_6691);
nand U7593 (N_7593,N_6595,N_6697);
nand U7594 (N_7594,N_6441,N_6872);
and U7595 (N_7595,N_6535,N_6157);
nand U7596 (N_7596,N_6128,N_6479);
or U7597 (N_7597,N_6848,N_6075);
and U7598 (N_7598,N_6741,N_6601);
nand U7599 (N_7599,N_6125,N_6094);
or U7600 (N_7600,N_6907,N_6439);
nor U7601 (N_7601,N_6339,N_6708);
or U7602 (N_7602,N_6585,N_6802);
and U7603 (N_7603,N_6240,N_6517);
nand U7604 (N_7604,N_6392,N_6546);
nand U7605 (N_7605,N_6013,N_6753);
xnor U7606 (N_7606,N_6881,N_6022);
nor U7607 (N_7607,N_6884,N_6969);
nand U7608 (N_7608,N_6186,N_6499);
or U7609 (N_7609,N_6601,N_6696);
nand U7610 (N_7610,N_6074,N_6675);
and U7611 (N_7611,N_6310,N_6618);
and U7612 (N_7612,N_6229,N_6265);
or U7613 (N_7613,N_6900,N_6983);
and U7614 (N_7614,N_6768,N_6259);
nand U7615 (N_7615,N_6304,N_6971);
and U7616 (N_7616,N_6971,N_6778);
nand U7617 (N_7617,N_6758,N_6257);
nand U7618 (N_7618,N_6964,N_6569);
nand U7619 (N_7619,N_6903,N_6267);
or U7620 (N_7620,N_6226,N_6106);
or U7621 (N_7621,N_6076,N_6462);
or U7622 (N_7622,N_6061,N_6982);
nor U7623 (N_7623,N_6941,N_6834);
nor U7624 (N_7624,N_6034,N_6414);
or U7625 (N_7625,N_6977,N_6894);
and U7626 (N_7626,N_6119,N_6082);
nand U7627 (N_7627,N_6231,N_6284);
and U7628 (N_7628,N_6935,N_6670);
or U7629 (N_7629,N_6936,N_6663);
or U7630 (N_7630,N_6478,N_6406);
nor U7631 (N_7631,N_6544,N_6073);
and U7632 (N_7632,N_6724,N_6736);
nor U7633 (N_7633,N_6720,N_6207);
or U7634 (N_7634,N_6791,N_6130);
nand U7635 (N_7635,N_6259,N_6029);
and U7636 (N_7636,N_6023,N_6308);
or U7637 (N_7637,N_6360,N_6651);
or U7638 (N_7638,N_6948,N_6321);
nor U7639 (N_7639,N_6338,N_6125);
and U7640 (N_7640,N_6983,N_6074);
nor U7641 (N_7641,N_6482,N_6164);
and U7642 (N_7642,N_6415,N_6564);
and U7643 (N_7643,N_6006,N_6305);
nand U7644 (N_7644,N_6669,N_6109);
and U7645 (N_7645,N_6127,N_6630);
or U7646 (N_7646,N_6932,N_6537);
or U7647 (N_7647,N_6304,N_6423);
or U7648 (N_7648,N_6396,N_6569);
or U7649 (N_7649,N_6400,N_6922);
nand U7650 (N_7650,N_6695,N_6779);
and U7651 (N_7651,N_6473,N_6863);
or U7652 (N_7652,N_6990,N_6094);
or U7653 (N_7653,N_6701,N_6205);
and U7654 (N_7654,N_6104,N_6809);
and U7655 (N_7655,N_6254,N_6367);
nand U7656 (N_7656,N_6061,N_6454);
or U7657 (N_7657,N_6585,N_6530);
and U7658 (N_7658,N_6339,N_6236);
nor U7659 (N_7659,N_6117,N_6373);
and U7660 (N_7660,N_6216,N_6678);
nor U7661 (N_7661,N_6928,N_6003);
and U7662 (N_7662,N_6301,N_6361);
nand U7663 (N_7663,N_6745,N_6708);
and U7664 (N_7664,N_6710,N_6526);
nor U7665 (N_7665,N_6607,N_6837);
nor U7666 (N_7666,N_6745,N_6155);
or U7667 (N_7667,N_6304,N_6791);
nand U7668 (N_7668,N_6910,N_6716);
nand U7669 (N_7669,N_6254,N_6074);
and U7670 (N_7670,N_6303,N_6781);
or U7671 (N_7671,N_6360,N_6131);
or U7672 (N_7672,N_6754,N_6114);
and U7673 (N_7673,N_6553,N_6559);
or U7674 (N_7674,N_6577,N_6738);
and U7675 (N_7675,N_6481,N_6558);
nand U7676 (N_7676,N_6832,N_6411);
nor U7677 (N_7677,N_6311,N_6727);
and U7678 (N_7678,N_6970,N_6164);
and U7679 (N_7679,N_6301,N_6189);
nand U7680 (N_7680,N_6994,N_6720);
or U7681 (N_7681,N_6389,N_6770);
and U7682 (N_7682,N_6879,N_6985);
and U7683 (N_7683,N_6508,N_6947);
or U7684 (N_7684,N_6153,N_6482);
nor U7685 (N_7685,N_6431,N_6261);
and U7686 (N_7686,N_6313,N_6749);
nand U7687 (N_7687,N_6246,N_6332);
and U7688 (N_7688,N_6793,N_6916);
nor U7689 (N_7689,N_6959,N_6860);
or U7690 (N_7690,N_6468,N_6252);
xnor U7691 (N_7691,N_6994,N_6580);
nor U7692 (N_7692,N_6836,N_6768);
and U7693 (N_7693,N_6340,N_6780);
nor U7694 (N_7694,N_6641,N_6294);
or U7695 (N_7695,N_6556,N_6409);
nand U7696 (N_7696,N_6784,N_6913);
nor U7697 (N_7697,N_6938,N_6617);
nor U7698 (N_7698,N_6833,N_6983);
nand U7699 (N_7699,N_6941,N_6438);
and U7700 (N_7700,N_6996,N_6129);
nand U7701 (N_7701,N_6232,N_6645);
and U7702 (N_7702,N_6984,N_6856);
nand U7703 (N_7703,N_6300,N_6881);
nor U7704 (N_7704,N_6439,N_6563);
nor U7705 (N_7705,N_6250,N_6210);
and U7706 (N_7706,N_6744,N_6542);
and U7707 (N_7707,N_6952,N_6710);
nor U7708 (N_7708,N_6496,N_6002);
or U7709 (N_7709,N_6075,N_6395);
nand U7710 (N_7710,N_6602,N_6878);
nand U7711 (N_7711,N_6137,N_6743);
nor U7712 (N_7712,N_6045,N_6699);
and U7713 (N_7713,N_6753,N_6378);
nand U7714 (N_7714,N_6960,N_6054);
or U7715 (N_7715,N_6244,N_6487);
nor U7716 (N_7716,N_6004,N_6919);
or U7717 (N_7717,N_6211,N_6364);
nor U7718 (N_7718,N_6760,N_6661);
nor U7719 (N_7719,N_6238,N_6198);
or U7720 (N_7720,N_6128,N_6218);
and U7721 (N_7721,N_6930,N_6786);
nand U7722 (N_7722,N_6407,N_6322);
nor U7723 (N_7723,N_6839,N_6922);
and U7724 (N_7724,N_6492,N_6247);
or U7725 (N_7725,N_6001,N_6783);
nor U7726 (N_7726,N_6794,N_6411);
nand U7727 (N_7727,N_6114,N_6176);
nand U7728 (N_7728,N_6079,N_6356);
or U7729 (N_7729,N_6932,N_6954);
nor U7730 (N_7730,N_6362,N_6772);
nand U7731 (N_7731,N_6123,N_6901);
or U7732 (N_7732,N_6503,N_6143);
or U7733 (N_7733,N_6190,N_6983);
nor U7734 (N_7734,N_6412,N_6620);
nand U7735 (N_7735,N_6665,N_6912);
nor U7736 (N_7736,N_6530,N_6058);
nand U7737 (N_7737,N_6897,N_6074);
nor U7738 (N_7738,N_6636,N_6649);
and U7739 (N_7739,N_6770,N_6958);
or U7740 (N_7740,N_6212,N_6207);
and U7741 (N_7741,N_6727,N_6935);
nor U7742 (N_7742,N_6753,N_6407);
nor U7743 (N_7743,N_6653,N_6890);
nand U7744 (N_7744,N_6265,N_6667);
nor U7745 (N_7745,N_6560,N_6427);
nor U7746 (N_7746,N_6759,N_6113);
nor U7747 (N_7747,N_6295,N_6836);
nor U7748 (N_7748,N_6681,N_6180);
nand U7749 (N_7749,N_6117,N_6196);
and U7750 (N_7750,N_6580,N_6774);
nor U7751 (N_7751,N_6162,N_6029);
and U7752 (N_7752,N_6315,N_6681);
and U7753 (N_7753,N_6624,N_6612);
nand U7754 (N_7754,N_6357,N_6100);
and U7755 (N_7755,N_6200,N_6145);
and U7756 (N_7756,N_6308,N_6909);
nand U7757 (N_7757,N_6918,N_6208);
nand U7758 (N_7758,N_6161,N_6177);
nor U7759 (N_7759,N_6543,N_6597);
or U7760 (N_7760,N_6131,N_6911);
nand U7761 (N_7761,N_6452,N_6284);
and U7762 (N_7762,N_6022,N_6728);
xor U7763 (N_7763,N_6014,N_6733);
nand U7764 (N_7764,N_6636,N_6702);
or U7765 (N_7765,N_6260,N_6036);
nand U7766 (N_7766,N_6159,N_6882);
nand U7767 (N_7767,N_6684,N_6938);
and U7768 (N_7768,N_6903,N_6334);
or U7769 (N_7769,N_6402,N_6215);
and U7770 (N_7770,N_6906,N_6513);
nor U7771 (N_7771,N_6406,N_6609);
nor U7772 (N_7772,N_6792,N_6560);
or U7773 (N_7773,N_6623,N_6221);
nor U7774 (N_7774,N_6398,N_6092);
nand U7775 (N_7775,N_6738,N_6866);
nand U7776 (N_7776,N_6003,N_6966);
nor U7777 (N_7777,N_6264,N_6791);
nand U7778 (N_7778,N_6212,N_6022);
and U7779 (N_7779,N_6793,N_6501);
or U7780 (N_7780,N_6127,N_6654);
nor U7781 (N_7781,N_6634,N_6848);
and U7782 (N_7782,N_6261,N_6095);
or U7783 (N_7783,N_6640,N_6158);
xor U7784 (N_7784,N_6466,N_6013);
nand U7785 (N_7785,N_6628,N_6929);
nand U7786 (N_7786,N_6475,N_6593);
or U7787 (N_7787,N_6709,N_6048);
and U7788 (N_7788,N_6993,N_6137);
or U7789 (N_7789,N_6557,N_6621);
nor U7790 (N_7790,N_6932,N_6417);
xnor U7791 (N_7791,N_6730,N_6014);
xnor U7792 (N_7792,N_6050,N_6479);
nand U7793 (N_7793,N_6232,N_6825);
and U7794 (N_7794,N_6413,N_6572);
nand U7795 (N_7795,N_6076,N_6999);
nor U7796 (N_7796,N_6671,N_6652);
nand U7797 (N_7797,N_6597,N_6500);
nor U7798 (N_7798,N_6700,N_6386);
nor U7799 (N_7799,N_6744,N_6668);
and U7800 (N_7800,N_6358,N_6370);
and U7801 (N_7801,N_6052,N_6771);
or U7802 (N_7802,N_6036,N_6317);
or U7803 (N_7803,N_6765,N_6972);
nand U7804 (N_7804,N_6673,N_6190);
and U7805 (N_7805,N_6355,N_6510);
and U7806 (N_7806,N_6049,N_6860);
nand U7807 (N_7807,N_6184,N_6926);
and U7808 (N_7808,N_6973,N_6487);
nand U7809 (N_7809,N_6077,N_6846);
or U7810 (N_7810,N_6070,N_6357);
nor U7811 (N_7811,N_6401,N_6796);
nor U7812 (N_7812,N_6636,N_6364);
nor U7813 (N_7813,N_6427,N_6723);
nor U7814 (N_7814,N_6610,N_6483);
nand U7815 (N_7815,N_6884,N_6674);
and U7816 (N_7816,N_6437,N_6377);
nand U7817 (N_7817,N_6221,N_6293);
or U7818 (N_7818,N_6487,N_6475);
nor U7819 (N_7819,N_6898,N_6177);
and U7820 (N_7820,N_6354,N_6265);
or U7821 (N_7821,N_6917,N_6507);
or U7822 (N_7822,N_6462,N_6193);
nor U7823 (N_7823,N_6989,N_6407);
and U7824 (N_7824,N_6292,N_6536);
and U7825 (N_7825,N_6319,N_6073);
or U7826 (N_7826,N_6569,N_6194);
nand U7827 (N_7827,N_6153,N_6508);
and U7828 (N_7828,N_6858,N_6474);
xnor U7829 (N_7829,N_6426,N_6595);
nand U7830 (N_7830,N_6195,N_6584);
nor U7831 (N_7831,N_6552,N_6616);
nand U7832 (N_7832,N_6100,N_6999);
or U7833 (N_7833,N_6370,N_6016);
nand U7834 (N_7834,N_6270,N_6879);
and U7835 (N_7835,N_6692,N_6312);
and U7836 (N_7836,N_6992,N_6243);
or U7837 (N_7837,N_6257,N_6144);
and U7838 (N_7838,N_6162,N_6730);
or U7839 (N_7839,N_6606,N_6461);
nor U7840 (N_7840,N_6218,N_6992);
and U7841 (N_7841,N_6683,N_6187);
or U7842 (N_7842,N_6698,N_6155);
nor U7843 (N_7843,N_6642,N_6992);
nor U7844 (N_7844,N_6828,N_6816);
nand U7845 (N_7845,N_6808,N_6927);
nor U7846 (N_7846,N_6836,N_6204);
and U7847 (N_7847,N_6593,N_6005);
nor U7848 (N_7848,N_6925,N_6802);
and U7849 (N_7849,N_6696,N_6964);
or U7850 (N_7850,N_6461,N_6045);
nand U7851 (N_7851,N_6518,N_6883);
nor U7852 (N_7852,N_6590,N_6161);
nor U7853 (N_7853,N_6316,N_6429);
nand U7854 (N_7854,N_6388,N_6838);
and U7855 (N_7855,N_6644,N_6822);
and U7856 (N_7856,N_6381,N_6750);
and U7857 (N_7857,N_6499,N_6704);
nor U7858 (N_7858,N_6594,N_6043);
and U7859 (N_7859,N_6741,N_6398);
nor U7860 (N_7860,N_6773,N_6108);
nor U7861 (N_7861,N_6977,N_6907);
and U7862 (N_7862,N_6112,N_6832);
and U7863 (N_7863,N_6132,N_6832);
and U7864 (N_7864,N_6058,N_6539);
nor U7865 (N_7865,N_6789,N_6762);
and U7866 (N_7866,N_6188,N_6277);
or U7867 (N_7867,N_6738,N_6000);
nand U7868 (N_7868,N_6068,N_6010);
and U7869 (N_7869,N_6154,N_6371);
or U7870 (N_7870,N_6294,N_6287);
and U7871 (N_7871,N_6510,N_6900);
nand U7872 (N_7872,N_6017,N_6410);
or U7873 (N_7873,N_6238,N_6907);
and U7874 (N_7874,N_6552,N_6060);
nor U7875 (N_7875,N_6679,N_6551);
xnor U7876 (N_7876,N_6070,N_6178);
nand U7877 (N_7877,N_6986,N_6077);
or U7878 (N_7878,N_6088,N_6635);
or U7879 (N_7879,N_6314,N_6258);
nor U7880 (N_7880,N_6662,N_6454);
nand U7881 (N_7881,N_6190,N_6916);
and U7882 (N_7882,N_6452,N_6862);
or U7883 (N_7883,N_6460,N_6768);
and U7884 (N_7884,N_6214,N_6536);
or U7885 (N_7885,N_6546,N_6248);
nor U7886 (N_7886,N_6746,N_6193);
and U7887 (N_7887,N_6839,N_6967);
and U7888 (N_7888,N_6236,N_6338);
nand U7889 (N_7889,N_6784,N_6686);
nand U7890 (N_7890,N_6600,N_6337);
or U7891 (N_7891,N_6343,N_6546);
nand U7892 (N_7892,N_6456,N_6416);
nor U7893 (N_7893,N_6219,N_6615);
nand U7894 (N_7894,N_6069,N_6227);
or U7895 (N_7895,N_6157,N_6061);
and U7896 (N_7896,N_6174,N_6364);
or U7897 (N_7897,N_6275,N_6717);
and U7898 (N_7898,N_6148,N_6110);
or U7899 (N_7899,N_6221,N_6525);
and U7900 (N_7900,N_6838,N_6449);
and U7901 (N_7901,N_6060,N_6353);
nor U7902 (N_7902,N_6216,N_6335);
nand U7903 (N_7903,N_6640,N_6210);
nand U7904 (N_7904,N_6583,N_6575);
xnor U7905 (N_7905,N_6013,N_6275);
or U7906 (N_7906,N_6975,N_6405);
or U7907 (N_7907,N_6768,N_6150);
nand U7908 (N_7908,N_6901,N_6410);
nor U7909 (N_7909,N_6481,N_6775);
and U7910 (N_7910,N_6616,N_6389);
or U7911 (N_7911,N_6326,N_6209);
nand U7912 (N_7912,N_6847,N_6701);
and U7913 (N_7913,N_6925,N_6909);
nand U7914 (N_7914,N_6500,N_6361);
nor U7915 (N_7915,N_6520,N_6635);
or U7916 (N_7916,N_6076,N_6390);
nor U7917 (N_7917,N_6614,N_6195);
nor U7918 (N_7918,N_6525,N_6969);
and U7919 (N_7919,N_6479,N_6127);
nand U7920 (N_7920,N_6881,N_6430);
xor U7921 (N_7921,N_6079,N_6527);
and U7922 (N_7922,N_6998,N_6860);
nand U7923 (N_7923,N_6949,N_6865);
and U7924 (N_7924,N_6161,N_6016);
or U7925 (N_7925,N_6070,N_6246);
nand U7926 (N_7926,N_6512,N_6029);
and U7927 (N_7927,N_6519,N_6534);
xnor U7928 (N_7928,N_6594,N_6671);
nand U7929 (N_7929,N_6035,N_6241);
or U7930 (N_7930,N_6696,N_6526);
and U7931 (N_7931,N_6391,N_6338);
and U7932 (N_7932,N_6341,N_6415);
nand U7933 (N_7933,N_6332,N_6067);
nand U7934 (N_7934,N_6886,N_6764);
nand U7935 (N_7935,N_6285,N_6139);
nand U7936 (N_7936,N_6156,N_6573);
nor U7937 (N_7937,N_6954,N_6454);
nor U7938 (N_7938,N_6960,N_6248);
nor U7939 (N_7939,N_6753,N_6614);
nor U7940 (N_7940,N_6903,N_6633);
and U7941 (N_7941,N_6189,N_6719);
or U7942 (N_7942,N_6218,N_6807);
or U7943 (N_7943,N_6495,N_6360);
nor U7944 (N_7944,N_6134,N_6365);
nor U7945 (N_7945,N_6685,N_6456);
nand U7946 (N_7946,N_6713,N_6126);
nor U7947 (N_7947,N_6110,N_6850);
nor U7948 (N_7948,N_6656,N_6189);
and U7949 (N_7949,N_6900,N_6815);
nand U7950 (N_7950,N_6368,N_6846);
nand U7951 (N_7951,N_6563,N_6390);
nor U7952 (N_7952,N_6117,N_6977);
or U7953 (N_7953,N_6181,N_6380);
nand U7954 (N_7954,N_6458,N_6845);
or U7955 (N_7955,N_6140,N_6385);
nor U7956 (N_7956,N_6072,N_6997);
or U7957 (N_7957,N_6402,N_6222);
and U7958 (N_7958,N_6684,N_6763);
nand U7959 (N_7959,N_6037,N_6298);
or U7960 (N_7960,N_6091,N_6117);
nor U7961 (N_7961,N_6942,N_6650);
or U7962 (N_7962,N_6554,N_6438);
nand U7963 (N_7963,N_6596,N_6807);
or U7964 (N_7964,N_6945,N_6681);
nor U7965 (N_7965,N_6581,N_6260);
and U7966 (N_7966,N_6136,N_6696);
nor U7967 (N_7967,N_6371,N_6676);
or U7968 (N_7968,N_6222,N_6234);
and U7969 (N_7969,N_6491,N_6587);
nor U7970 (N_7970,N_6237,N_6123);
nand U7971 (N_7971,N_6777,N_6598);
and U7972 (N_7972,N_6010,N_6626);
or U7973 (N_7973,N_6806,N_6149);
nand U7974 (N_7974,N_6269,N_6888);
nor U7975 (N_7975,N_6677,N_6676);
nor U7976 (N_7976,N_6793,N_6678);
nor U7977 (N_7977,N_6110,N_6952);
nor U7978 (N_7978,N_6814,N_6933);
nor U7979 (N_7979,N_6291,N_6932);
nand U7980 (N_7980,N_6919,N_6673);
and U7981 (N_7981,N_6991,N_6015);
nand U7982 (N_7982,N_6269,N_6726);
nor U7983 (N_7983,N_6354,N_6804);
nor U7984 (N_7984,N_6844,N_6645);
nor U7985 (N_7985,N_6170,N_6110);
and U7986 (N_7986,N_6168,N_6316);
nor U7987 (N_7987,N_6945,N_6868);
or U7988 (N_7988,N_6377,N_6322);
xnor U7989 (N_7989,N_6289,N_6051);
nor U7990 (N_7990,N_6346,N_6685);
nand U7991 (N_7991,N_6027,N_6004);
or U7992 (N_7992,N_6101,N_6650);
and U7993 (N_7993,N_6763,N_6564);
and U7994 (N_7994,N_6889,N_6570);
and U7995 (N_7995,N_6726,N_6738);
or U7996 (N_7996,N_6877,N_6196);
nor U7997 (N_7997,N_6435,N_6797);
and U7998 (N_7998,N_6321,N_6553);
nor U7999 (N_7999,N_6950,N_6400);
or U8000 (N_8000,N_7833,N_7528);
and U8001 (N_8001,N_7429,N_7614);
and U8002 (N_8002,N_7876,N_7825);
or U8003 (N_8003,N_7423,N_7730);
and U8004 (N_8004,N_7484,N_7097);
and U8005 (N_8005,N_7347,N_7225);
nor U8006 (N_8006,N_7633,N_7164);
and U8007 (N_8007,N_7741,N_7805);
or U8008 (N_8008,N_7778,N_7682);
nand U8009 (N_8009,N_7773,N_7177);
and U8010 (N_8010,N_7385,N_7068);
and U8011 (N_8011,N_7259,N_7257);
nand U8012 (N_8012,N_7529,N_7989);
nor U8013 (N_8013,N_7443,N_7731);
nor U8014 (N_8014,N_7502,N_7724);
nand U8015 (N_8015,N_7265,N_7692);
and U8016 (N_8016,N_7624,N_7428);
nor U8017 (N_8017,N_7238,N_7698);
nor U8018 (N_8018,N_7509,N_7954);
nand U8019 (N_8019,N_7699,N_7290);
nor U8020 (N_8020,N_7223,N_7754);
nor U8021 (N_8021,N_7104,N_7186);
or U8022 (N_8022,N_7439,N_7887);
nor U8023 (N_8023,N_7664,N_7233);
or U8024 (N_8024,N_7365,N_7878);
and U8025 (N_8025,N_7372,N_7222);
nor U8026 (N_8026,N_7626,N_7732);
nor U8027 (N_8027,N_7888,N_7143);
or U8028 (N_8028,N_7601,N_7487);
nand U8029 (N_8029,N_7471,N_7140);
nand U8030 (N_8030,N_7062,N_7415);
and U8031 (N_8031,N_7038,N_7941);
nand U8032 (N_8032,N_7437,N_7519);
nor U8033 (N_8033,N_7670,N_7100);
or U8034 (N_8034,N_7031,N_7786);
nor U8035 (N_8035,N_7102,N_7524);
nand U8036 (N_8036,N_7348,N_7974);
and U8037 (N_8037,N_7420,N_7854);
nor U8038 (N_8038,N_7880,N_7148);
or U8039 (N_8039,N_7351,N_7119);
nor U8040 (N_8040,N_7214,N_7976);
or U8041 (N_8041,N_7046,N_7053);
nand U8042 (N_8042,N_7149,N_7934);
or U8043 (N_8043,N_7714,N_7334);
or U8044 (N_8044,N_7340,N_7460);
or U8045 (N_8045,N_7433,N_7526);
and U8046 (N_8046,N_7708,N_7693);
nand U8047 (N_8047,N_7758,N_7281);
or U8048 (N_8048,N_7826,N_7820);
or U8049 (N_8049,N_7644,N_7126);
or U8050 (N_8050,N_7459,N_7444);
nor U8051 (N_8051,N_7364,N_7333);
nand U8052 (N_8052,N_7517,N_7554);
nand U8053 (N_8053,N_7915,N_7092);
nor U8054 (N_8054,N_7877,N_7268);
nand U8055 (N_8055,N_7435,N_7606);
or U8056 (N_8056,N_7921,N_7246);
nand U8057 (N_8057,N_7740,N_7330);
nand U8058 (N_8058,N_7011,N_7098);
nand U8059 (N_8059,N_7173,N_7962);
nor U8060 (N_8060,N_7811,N_7094);
or U8061 (N_8061,N_7118,N_7522);
nand U8062 (N_8062,N_7605,N_7386);
nand U8063 (N_8063,N_7367,N_7231);
and U8064 (N_8064,N_7065,N_7061);
or U8065 (N_8065,N_7768,N_7926);
nor U8066 (N_8066,N_7319,N_7288);
nor U8067 (N_8067,N_7586,N_7760);
nand U8068 (N_8068,N_7729,N_7360);
nand U8069 (N_8069,N_7623,N_7393);
and U8070 (N_8070,N_7870,N_7631);
nand U8071 (N_8071,N_7599,N_7668);
and U8072 (N_8072,N_7252,N_7142);
or U8073 (N_8073,N_7205,N_7906);
nor U8074 (N_8074,N_7822,N_7597);
nor U8075 (N_8075,N_7950,N_7085);
or U8076 (N_8076,N_7379,N_7841);
or U8077 (N_8077,N_7882,N_7520);
or U8078 (N_8078,N_7442,N_7852);
nor U8079 (N_8079,N_7331,N_7516);
nor U8080 (N_8080,N_7696,N_7553);
xnor U8081 (N_8081,N_7910,N_7803);
and U8082 (N_8082,N_7918,N_7325);
nand U8083 (N_8083,N_7530,N_7305);
nor U8084 (N_8084,N_7078,N_7132);
and U8085 (N_8085,N_7979,N_7397);
or U8086 (N_8086,N_7669,N_7712);
nand U8087 (N_8087,N_7680,N_7781);
nand U8088 (N_8088,N_7909,N_7081);
nor U8089 (N_8089,N_7609,N_7534);
or U8090 (N_8090,N_7258,N_7230);
nand U8091 (N_8091,N_7055,N_7001);
nor U8092 (N_8092,N_7799,N_7790);
or U8093 (N_8093,N_7480,N_7141);
or U8094 (N_8094,N_7335,N_7581);
nor U8095 (N_8095,N_7309,N_7616);
nor U8096 (N_8096,N_7892,N_7550);
and U8097 (N_8097,N_7017,N_7253);
nor U8098 (N_8098,N_7076,N_7184);
and U8099 (N_8099,N_7042,N_7172);
nor U8100 (N_8100,N_7855,N_7112);
nand U8101 (N_8101,N_7815,N_7776);
nor U8102 (N_8102,N_7703,N_7843);
and U8103 (N_8103,N_7720,N_7646);
and U8104 (N_8104,N_7908,N_7084);
or U8105 (N_8105,N_7717,N_7189);
and U8106 (N_8106,N_7679,N_7168);
and U8107 (N_8107,N_7861,N_7987);
nand U8108 (N_8108,N_7795,N_7774);
nand U8109 (N_8109,N_7035,N_7551);
nand U8110 (N_8110,N_7713,N_7536);
nor U8111 (N_8111,N_7206,N_7090);
nand U8112 (N_8112,N_7198,N_7697);
and U8113 (N_8113,N_7127,N_7959);
nand U8114 (N_8114,N_7337,N_7949);
and U8115 (N_8115,N_7845,N_7951);
nand U8116 (N_8116,N_7557,N_7492);
nand U8117 (N_8117,N_7326,N_7207);
and U8118 (N_8118,N_7371,N_7596);
nand U8119 (N_8119,N_7229,N_7436);
and U8120 (N_8120,N_7812,N_7525);
and U8121 (N_8121,N_7511,N_7802);
and U8122 (N_8122,N_7817,N_7830);
nand U8123 (N_8123,N_7508,N_7834);
and U8124 (N_8124,N_7036,N_7568);
nor U8125 (N_8125,N_7838,N_7899);
nor U8126 (N_8126,N_7089,N_7277);
nor U8127 (N_8127,N_7515,N_7975);
nand U8128 (N_8128,N_7985,N_7220);
or U8129 (N_8129,N_7647,N_7706);
or U8130 (N_8130,N_7789,N_7872);
nor U8131 (N_8131,N_7642,N_7700);
nor U8132 (N_8132,N_7737,N_7294);
nor U8133 (N_8133,N_7014,N_7472);
or U8134 (N_8134,N_7757,N_7973);
nor U8135 (N_8135,N_7124,N_7441);
and U8136 (N_8136,N_7864,N_7868);
nor U8137 (N_8137,N_7953,N_7398);
or U8138 (N_8138,N_7968,N_7945);
nor U8139 (N_8139,N_7159,N_7339);
nor U8140 (N_8140,N_7082,N_7312);
nor U8141 (N_8141,N_7702,N_7010);
or U8142 (N_8142,N_7327,N_7577);
nand U8143 (N_8143,N_7542,N_7400);
nor U8144 (N_8144,N_7659,N_7044);
nand U8145 (N_8145,N_7146,N_7376);
nor U8146 (N_8146,N_7565,N_7373);
nand U8147 (N_8147,N_7948,N_7448);
nor U8148 (N_8148,N_7540,N_7590);
and U8149 (N_8149,N_7637,N_7734);
nor U8150 (N_8150,N_7719,N_7675);
and U8151 (N_8151,N_7070,N_7662);
nor U8152 (N_8152,N_7282,N_7363);
nor U8153 (N_8153,N_7514,N_7005);
or U8154 (N_8154,N_7167,N_7969);
nor U8155 (N_8155,N_7176,N_7285);
and U8156 (N_8156,N_7871,N_7598);
nor U8157 (N_8157,N_7928,N_7671);
nand U8158 (N_8158,N_7937,N_7547);
or U8159 (N_8159,N_7978,N_7728);
or U8160 (N_8160,N_7279,N_7869);
or U8161 (N_8161,N_7162,N_7136);
nor U8162 (N_8162,N_7344,N_7762);
nor U8163 (N_8163,N_7504,N_7970);
nor U8164 (N_8164,N_7473,N_7286);
or U8165 (N_8165,N_7684,N_7401);
and U8166 (N_8166,N_7851,N_7410);
or U8167 (N_8167,N_7897,N_7125);
and U8168 (N_8168,N_7865,N_7071);
nor U8169 (N_8169,N_7602,N_7984);
or U8170 (N_8170,N_7656,N_7993);
and U8171 (N_8171,N_7007,N_7863);
or U8172 (N_8172,N_7801,N_7893);
nand U8173 (N_8173,N_7109,N_7254);
and U8174 (N_8174,N_7578,N_7711);
nand U8175 (N_8175,N_7414,N_7823);
or U8176 (N_8176,N_7224,N_7208);
or U8177 (N_8177,N_7181,N_7242);
and U8178 (N_8178,N_7287,N_7579);
nand U8179 (N_8179,N_7715,N_7583);
nand U8180 (N_8180,N_7391,N_7913);
nand U8181 (N_8181,N_7328,N_7532);
or U8182 (N_8182,N_7292,N_7678);
nor U8183 (N_8183,N_7635,N_7756);
nor U8184 (N_8184,N_7029,N_7408);
nand U8185 (N_8185,N_7641,N_7827);
or U8186 (N_8186,N_7636,N_7625);
nand U8187 (N_8187,N_7710,N_7063);
or U8188 (N_8188,N_7981,N_7990);
nand U8189 (N_8189,N_7034,N_7705);
nand U8190 (N_8190,N_7828,N_7170);
nand U8191 (N_8191,N_7936,N_7831);
nand U8192 (N_8192,N_7957,N_7383);
nor U8193 (N_8193,N_7153,N_7483);
nor U8194 (N_8194,N_7867,N_7160);
and U8195 (N_8195,N_7751,N_7311);
nand U8196 (N_8196,N_7417,N_7932);
nor U8197 (N_8197,N_7019,N_7824);
and U8198 (N_8198,N_7411,N_7133);
nand U8199 (N_8199,N_7537,N_7341);
nor U8200 (N_8200,N_7195,N_7800);
nor U8201 (N_8201,N_7667,N_7427);
nor U8202 (N_8202,N_7057,N_7556);
nand U8203 (N_8203,N_7559,N_7938);
nand U8204 (N_8204,N_7091,N_7180);
and U8205 (N_8205,N_7308,N_7901);
nor U8206 (N_8206,N_7192,N_7849);
and U8207 (N_8207,N_7779,N_7390);
or U8208 (N_8208,N_7298,N_7512);
nand U8209 (N_8209,N_7545,N_7021);
or U8210 (N_8210,N_7002,N_7507);
and U8211 (N_8211,N_7485,N_7748);
and U8212 (N_8212,N_7501,N_7307);
nand U8213 (N_8213,N_7389,N_7612);
nor U8214 (N_8214,N_7155,N_7174);
or U8215 (N_8215,N_7025,N_7235);
nand U8216 (N_8216,N_7110,N_7267);
or U8217 (N_8217,N_7182,N_7873);
and U8218 (N_8218,N_7709,N_7301);
nand U8219 (N_8219,N_7128,N_7505);
nand U8220 (N_8220,N_7016,N_7197);
nor U8221 (N_8221,N_7481,N_7818);
nor U8222 (N_8222,N_7695,N_7573);
nand U8223 (N_8223,N_7875,N_7278);
nor U8224 (N_8224,N_7560,N_7771);
nor U8225 (N_8225,N_7380,N_7083);
nor U8226 (N_8226,N_7617,N_7966);
and U8227 (N_8227,N_7458,N_7366);
or U8228 (N_8228,N_7353,N_7593);
xor U8229 (N_8229,N_7722,N_7881);
and U8230 (N_8230,N_7402,N_7388);
nor U8231 (N_8231,N_7093,N_7900);
nand U8232 (N_8232,N_7169,N_7850);
nor U8233 (N_8233,N_7660,N_7213);
nor U8234 (N_8234,N_7461,N_7039);
and U8235 (N_8235,N_7561,N_7199);
nand U8236 (N_8236,N_7270,N_7704);
nand U8237 (N_8237,N_7289,N_7156);
nand U8238 (N_8238,N_7359,N_7611);
and U8239 (N_8239,N_7067,N_7627);
nor U8240 (N_8240,N_7686,N_7580);
nor U8241 (N_8241,N_7368,N_7964);
or U8242 (N_8242,N_7193,N_7651);
nand U8243 (N_8243,N_7080,N_7009);
or U8244 (N_8244,N_7387,N_7432);
nor U8245 (N_8245,N_7217,N_7320);
or U8246 (N_8246,N_7058,N_7465);
and U8247 (N_8247,N_7582,N_7665);
nor U8248 (N_8248,N_7891,N_7994);
nor U8249 (N_8249,N_7295,N_7563);
or U8250 (N_8250,N_7707,N_7917);
and U8251 (N_8251,N_7269,N_7462);
nand U8252 (N_8252,N_7570,N_7054);
and U8253 (N_8253,N_7594,N_7629);
or U8254 (N_8254,N_7632,N_7299);
nand U8255 (N_8255,N_7761,N_7384);
nor U8256 (N_8256,N_7535,N_7056);
nor U8257 (N_8257,N_7575,N_7588);
or U8258 (N_8258,N_7099,N_7120);
nor U8259 (N_8259,N_7047,N_7455);
or U8260 (N_8260,N_7211,N_7293);
or U8261 (N_8261,N_7163,N_7933);
or U8262 (N_8262,N_7772,N_7382);
nand U8263 (N_8263,N_7450,N_7947);
nor U8264 (N_8264,N_7572,N_7694);
nand U8265 (N_8265,N_7188,N_7129);
or U8266 (N_8266,N_7832,N_7266);
nor U8267 (N_8267,N_7256,N_7321);
nor U8268 (N_8268,N_7610,N_7077);
and U8269 (N_8269,N_7316,N_7260);
and U8270 (N_8270,N_7451,N_7468);
and U8271 (N_8271,N_7890,N_7904);
and U8272 (N_8272,N_7490,N_7356);
nor U8273 (N_8273,N_7095,N_7944);
nand U8274 (N_8274,N_7381,N_7794);
and U8275 (N_8275,N_7226,N_7315);
or U8276 (N_8276,N_7131,N_7069);
or U8277 (N_8277,N_7343,N_7121);
nor U8278 (N_8278,N_7604,N_7958);
nor U8279 (N_8279,N_7555,N_7589);
or U8280 (N_8280,N_7105,N_7374);
nor U8281 (N_8281,N_7569,N_7539);
or U8282 (N_8282,N_7352,N_7809);
nand U8283 (N_8283,N_7621,N_7470);
nor U8284 (N_8284,N_7362,N_7350);
nor U8285 (N_8285,N_7424,N_7777);
nand U8286 (N_8286,N_7227,N_7988);
nor U8287 (N_8287,N_7785,N_7752);
nor U8288 (N_8288,N_7497,N_7767);
or U8289 (N_8289,N_7894,N_7237);
nor U8290 (N_8290,N_7543,N_7488);
nor U8291 (N_8291,N_7418,N_7718);
or U8292 (N_8292,N_7716,N_7775);
nand U8293 (N_8293,N_7615,N_7248);
or U8294 (N_8294,N_7187,N_7860);
nand U8295 (N_8295,N_7300,N_7840);
or U8296 (N_8296,N_7178,N_7123);
nor U8297 (N_8297,N_7619,N_7592);
nand U8298 (N_8298,N_7469,N_7920);
and U8299 (N_8299,N_7879,N_7049);
or U8300 (N_8300,N_7907,N_7313);
nand U8301 (N_8301,N_7464,N_7783);
or U8302 (N_8302,N_7037,N_7283);
or U8303 (N_8303,N_7232,N_7370);
or U8304 (N_8304,N_7422,N_7006);
nor U8305 (N_8305,N_7190,N_7276);
and U8306 (N_8306,N_7101,N_7902);
or U8307 (N_8307,N_7456,N_7073);
or U8308 (N_8308,N_7404,N_7243);
nor U8309 (N_8309,N_7438,N_7486);
nor U8310 (N_8310,N_7051,N_7796);
nand U8311 (N_8311,N_7275,N_7701);
nand U8312 (N_8312,N_7247,N_7130);
nand U8313 (N_8313,N_7527,N_7349);
and U8314 (N_8314,N_7329,N_7336);
or U8315 (N_8315,N_7273,N_7134);
and U8316 (N_8316,N_7640,N_7788);
or U8317 (N_8317,N_7262,N_7158);
xnor U8318 (N_8318,N_7804,N_7638);
nor U8319 (N_8319,N_7765,N_7430);
nand U8320 (N_8320,N_7690,N_7961);
nand U8321 (N_8321,N_7216,N_7332);
nand U8322 (N_8322,N_7079,N_7482);
nand U8323 (N_8323,N_7806,N_7000);
nor U8324 (N_8324,N_7986,N_7942);
and U8325 (N_8325,N_7952,N_7956);
nor U8326 (N_8326,N_7209,N_7033);
nor U8327 (N_8327,N_7742,N_7030);
and U8328 (N_8328,N_7249,N_7980);
nor U8329 (N_8329,N_7793,N_7658);
and U8330 (N_8330,N_7495,N_7191);
nor U8331 (N_8331,N_7735,N_7856);
nor U8332 (N_8332,N_7620,N_7013);
nand U8333 (N_8333,N_7999,N_7240);
xnor U8334 (N_8334,N_7323,N_7821);
nand U8335 (N_8335,N_7960,N_7466);
or U8336 (N_8336,N_7541,N_7060);
or U8337 (N_8337,N_7736,N_7144);
and U8338 (N_8338,N_7358,N_7296);
nand U8339 (N_8339,N_7903,N_7498);
nand U8340 (N_8340,N_7171,N_7396);
or U8341 (N_8341,N_7940,N_7674);
nor U8342 (N_8342,N_7784,N_7725);
and U8343 (N_8343,N_7585,N_7613);
or U8344 (N_8344,N_7607,N_7883);
and U8345 (N_8345,N_7816,N_7463);
nor U8346 (N_8346,N_7426,N_7139);
nand U8347 (N_8347,N_7489,N_7666);
nor U8348 (N_8348,N_7685,N_7244);
and U8349 (N_8349,N_7997,N_7431);
and U8350 (N_8350,N_7780,N_7965);
or U8351 (N_8351,N_7506,N_7836);
nand U8352 (N_8352,N_7221,N_7272);
nor U8353 (N_8353,N_7745,N_7531);
nand U8354 (N_8354,N_7064,N_7457);
and U8355 (N_8355,N_7923,N_7791);
or U8356 (N_8356,N_7683,N_7814);
nand U8357 (N_8357,N_7317,N_7755);
or U8358 (N_8358,N_7115,N_7819);
or U8359 (N_8359,N_7074,N_7835);
nor U8360 (N_8360,N_7931,N_7263);
nand U8361 (N_8361,N_7291,N_7407);
nor U8362 (N_8362,N_7150,N_7546);
xor U8363 (N_8363,N_7066,N_7770);
or U8364 (N_8364,N_7808,N_7212);
or U8365 (N_8365,N_7538,N_7653);
or U8366 (N_8366,N_7859,N_7510);
and U8367 (N_8367,N_7558,N_7759);
or U8368 (N_8368,N_7911,N_7043);
or U8369 (N_8369,N_7691,N_7261);
nor U8370 (N_8370,N_7677,N_7008);
nand U8371 (N_8371,N_7884,N_7727);
nor U8372 (N_8372,N_7346,N_7318);
nand U8373 (N_8373,N_7399,N_7750);
or U8374 (N_8374,N_7369,N_7764);
xor U8375 (N_8375,N_7518,N_7533);
or U8376 (N_8376,N_7354,N_7314);
and U8377 (N_8377,N_7255,N_7251);
or U8378 (N_8378,N_7655,N_7087);
nor U8379 (N_8379,N_7927,N_7147);
or U8380 (N_8380,N_7591,N_7274);
and U8381 (N_8381,N_7375,N_7419);
and U8382 (N_8382,N_7304,N_7322);
nor U8383 (N_8383,N_7412,N_7643);
or U8384 (N_8384,N_7107,N_7403);
nand U8385 (N_8385,N_7595,N_7858);
nand U8386 (N_8386,N_7652,N_7421);
or U8387 (N_8387,N_7500,N_7338);
or U8388 (N_8388,N_7241,N_7929);
or U8389 (N_8389,N_7434,N_7912);
and U8390 (N_8390,N_7681,N_7491);
nor U8391 (N_8391,N_7842,N_7072);
nand U8392 (N_8392,N_7574,N_7012);
and U8393 (N_8393,N_7185,N_7874);
nand U8394 (N_8394,N_7474,N_7452);
or U8395 (N_8395,N_7744,N_7862);
and U8396 (N_8396,N_7955,N_7250);
and U8397 (N_8397,N_7998,N_7648);
or U8398 (N_8398,N_7673,N_7145);
or U8399 (N_8399,N_7041,N_7991);
and U8400 (N_8400,N_7151,N_7889);
or U8401 (N_8401,N_7792,N_7446);
or U8402 (N_8402,N_7027,N_7165);
nor U8403 (N_8403,N_7924,N_7914);
nand U8404 (N_8404,N_7494,N_7797);
or U8405 (N_8405,N_7478,N_7117);
or U8406 (N_8406,N_7045,N_7857);
and U8407 (N_8407,N_7239,N_7634);
nand U8408 (N_8408,N_7161,N_7116);
nand U8409 (N_8409,N_7271,N_7608);
nand U8410 (N_8410,N_7747,N_7218);
and U8411 (N_8411,N_7245,N_7234);
nor U8412 (N_8412,N_7284,N_7630);
nor U8413 (N_8413,N_7023,N_7166);
nor U8414 (N_8414,N_7493,N_7848);
nor U8415 (N_8415,N_7086,N_7963);
and U8416 (N_8416,N_7687,N_7024);
or U8417 (N_8417,N_7749,N_7201);
or U8418 (N_8418,N_7739,N_7544);
or U8419 (N_8419,N_7576,N_7983);
nand U8420 (N_8420,N_7303,N_7813);
nor U8421 (N_8421,N_7015,N_7467);
and U8422 (N_8422,N_7114,N_7618);
nand U8423 (N_8423,N_7236,N_7584);
and U8424 (N_8424,N_7280,N_7440);
and U8425 (N_8425,N_7726,N_7088);
nor U8426 (N_8426,N_7183,N_7895);
nor U8427 (N_8427,N_7477,N_7106);
or U8428 (N_8428,N_7103,N_7196);
and U8429 (N_8429,N_7549,N_7721);
xor U8430 (N_8430,N_7919,N_7204);
and U8431 (N_8431,N_7154,N_7040);
nor U8432 (N_8432,N_7925,N_7743);
xor U8433 (N_8433,N_7971,N_7622);
and U8434 (N_8434,N_7122,N_7310);
nand U8435 (N_8435,N_7048,N_7769);
or U8436 (N_8436,N_7394,N_7137);
or U8437 (N_8437,N_7075,N_7898);
or U8438 (N_8438,N_7905,N_7676);
nor U8439 (N_8439,N_7567,N_7847);
and U8440 (N_8440,N_7175,N_7866);
nand U8441 (N_8441,N_7409,N_7406);
nor U8442 (N_8442,N_7967,N_7654);
or U8443 (N_8443,N_7157,N_7454);
nand U8444 (N_8444,N_7052,N_7059);
or U8445 (N_8445,N_7628,N_7521);
nor U8446 (N_8446,N_7499,N_7548);
and U8447 (N_8447,N_7324,N_7361);
nand U8448 (N_8448,N_7977,N_7829);
nor U8449 (N_8449,N_7004,N_7837);
or U8450 (N_8450,N_7787,N_7746);
xor U8451 (N_8451,N_7202,N_7203);
nand U8452 (N_8452,N_7113,N_7228);
or U8453 (N_8453,N_7566,N_7342);
nor U8454 (N_8454,N_7672,N_7453);
nand U8455 (N_8455,N_7302,N_7733);
nor U8456 (N_8456,N_7026,N_7523);
nor U8457 (N_8457,N_7723,N_7844);
and U8458 (N_8458,N_7810,N_7378);
and U8459 (N_8459,N_7603,N_7896);
and U8460 (N_8460,N_7395,N_7020);
or U8461 (N_8461,N_7946,N_7916);
and U8462 (N_8462,N_7886,N_7661);
or U8463 (N_8463,N_7416,N_7445);
and U8464 (N_8464,N_7306,N_7152);
or U8465 (N_8465,N_7688,N_7475);
nand U8466 (N_8466,N_7853,N_7018);
nor U8467 (N_8467,N_7972,N_7689);
and U8468 (N_8468,N_7476,N_7003);
or U8469 (N_8469,N_7210,N_7639);
nor U8470 (N_8470,N_7807,N_7111);
nor U8471 (N_8471,N_7405,N_7413);
nor U8472 (N_8472,N_7738,N_7377);
nand U8473 (N_8473,N_7885,N_7297);
nor U8474 (N_8474,N_7600,N_7447);
and U8475 (N_8475,N_7571,N_7552);
or U8476 (N_8476,N_7357,N_7930);
or U8477 (N_8477,N_7219,N_7846);
or U8478 (N_8478,N_7028,N_7513);
nor U8479 (N_8479,N_7650,N_7564);
nor U8480 (N_8480,N_7264,N_7345);
nor U8481 (N_8481,N_7392,N_7645);
nor U8482 (N_8482,N_7939,N_7200);
and U8483 (N_8483,N_7479,N_7649);
and U8484 (N_8484,N_7782,N_7503);
or U8485 (N_8485,N_7138,N_7425);
nor U8486 (N_8486,N_7032,N_7992);
and U8487 (N_8487,N_7935,N_7587);
nand U8488 (N_8488,N_7996,N_7022);
nand U8489 (N_8489,N_7766,N_7194);
or U8490 (N_8490,N_7562,N_7657);
nor U8491 (N_8491,N_7982,N_7995);
and U8492 (N_8492,N_7179,N_7050);
nor U8493 (N_8493,N_7922,N_7943);
nor U8494 (N_8494,N_7135,N_7215);
and U8495 (N_8495,N_7763,N_7663);
nor U8496 (N_8496,N_7108,N_7839);
and U8497 (N_8497,N_7496,N_7798);
or U8498 (N_8498,N_7096,N_7355);
nor U8499 (N_8499,N_7753,N_7449);
nand U8500 (N_8500,N_7456,N_7139);
or U8501 (N_8501,N_7860,N_7214);
or U8502 (N_8502,N_7435,N_7410);
nand U8503 (N_8503,N_7509,N_7764);
and U8504 (N_8504,N_7697,N_7405);
nand U8505 (N_8505,N_7531,N_7779);
nand U8506 (N_8506,N_7243,N_7948);
or U8507 (N_8507,N_7946,N_7619);
or U8508 (N_8508,N_7426,N_7561);
and U8509 (N_8509,N_7612,N_7788);
nand U8510 (N_8510,N_7895,N_7894);
nand U8511 (N_8511,N_7555,N_7541);
and U8512 (N_8512,N_7638,N_7206);
nand U8513 (N_8513,N_7415,N_7843);
or U8514 (N_8514,N_7651,N_7384);
nor U8515 (N_8515,N_7977,N_7476);
nand U8516 (N_8516,N_7827,N_7010);
nor U8517 (N_8517,N_7525,N_7825);
nor U8518 (N_8518,N_7477,N_7234);
nand U8519 (N_8519,N_7915,N_7978);
or U8520 (N_8520,N_7471,N_7644);
nand U8521 (N_8521,N_7323,N_7798);
nand U8522 (N_8522,N_7000,N_7543);
nand U8523 (N_8523,N_7096,N_7170);
nor U8524 (N_8524,N_7385,N_7349);
and U8525 (N_8525,N_7646,N_7551);
or U8526 (N_8526,N_7843,N_7033);
or U8527 (N_8527,N_7730,N_7474);
or U8528 (N_8528,N_7218,N_7532);
and U8529 (N_8529,N_7156,N_7638);
nand U8530 (N_8530,N_7107,N_7984);
or U8531 (N_8531,N_7252,N_7580);
nand U8532 (N_8532,N_7526,N_7290);
nor U8533 (N_8533,N_7166,N_7541);
nor U8534 (N_8534,N_7247,N_7470);
and U8535 (N_8535,N_7807,N_7064);
nand U8536 (N_8536,N_7877,N_7706);
and U8537 (N_8537,N_7836,N_7996);
nand U8538 (N_8538,N_7239,N_7664);
nor U8539 (N_8539,N_7663,N_7794);
or U8540 (N_8540,N_7091,N_7218);
or U8541 (N_8541,N_7495,N_7541);
nand U8542 (N_8542,N_7097,N_7810);
nand U8543 (N_8543,N_7003,N_7124);
xor U8544 (N_8544,N_7729,N_7026);
and U8545 (N_8545,N_7085,N_7590);
nor U8546 (N_8546,N_7776,N_7469);
or U8547 (N_8547,N_7109,N_7926);
and U8548 (N_8548,N_7814,N_7404);
nand U8549 (N_8549,N_7446,N_7559);
nor U8550 (N_8550,N_7739,N_7353);
nand U8551 (N_8551,N_7560,N_7908);
or U8552 (N_8552,N_7736,N_7411);
or U8553 (N_8553,N_7755,N_7689);
or U8554 (N_8554,N_7872,N_7972);
and U8555 (N_8555,N_7971,N_7352);
nand U8556 (N_8556,N_7860,N_7747);
and U8557 (N_8557,N_7179,N_7632);
nor U8558 (N_8558,N_7786,N_7643);
and U8559 (N_8559,N_7487,N_7845);
nand U8560 (N_8560,N_7679,N_7968);
nand U8561 (N_8561,N_7756,N_7902);
or U8562 (N_8562,N_7192,N_7461);
nand U8563 (N_8563,N_7045,N_7469);
nor U8564 (N_8564,N_7878,N_7299);
xnor U8565 (N_8565,N_7845,N_7357);
and U8566 (N_8566,N_7711,N_7055);
nand U8567 (N_8567,N_7993,N_7237);
nor U8568 (N_8568,N_7371,N_7224);
nand U8569 (N_8569,N_7294,N_7566);
nand U8570 (N_8570,N_7880,N_7000);
or U8571 (N_8571,N_7845,N_7289);
nand U8572 (N_8572,N_7235,N_7849);
or U8573 (N_8573,N_7131,N_7306);
and U8574 (N_8574,N_7840,N_7328);
xor U8575 (N_8575,N_7496,N_7520);
nand U8576 (N_8576,N_7693,N_7333);
or U8577 (N_8577,N_7940,N_7111);
or U8578 (N_8578,N_7844,N_7110);
or U8579 (N_8579,N_7822,N_7775);
nand U8580 (N_8580,N_7845,N_7198);
or U8581 (N_8581,N_7816,N_7527);
and U8582 (N_8582,N_7810,N_7223);
nand U8583 (N_8583,N_7655,N_7451);
nand U8584 (N_8584,N_7126,N_7667);
and U8585 (N_8585,N_7534,N_7265);
or U8586 (N_8586,N_7424,N_7659);
or U8587 (N_8587,N_7035,N_7082);
nand U8588 (N_8588,N_7288,N_7771);
nand U8589 (N_8589,N_7322,N_7769);
or U8590 (N_8590,N_7260,N_7590);
nor U8591 (N_8591,N_7396,N_7702);
xnor U8592 (N_8592,N_7861,N_7411);
nand U8593 (N_8593,N_7795,N_7275);
or U8594 (N_8594,N_7648,N_7729);
nand U8595 (N_8595,N_7376,N_7829);
or U8596 (N_8596,N_7852,N_7232);
nand U8597 (N_8597,N_7714,N_7409);
and U8598 (N_8598,N_7371,N_7826);
nand U8599 (N_8599,N_7205,N_7229);
nand U8600 (N_8600,N_7201,N_7577);
or U8601 (N_8601,N_7514,N_7315);
and U8602 (N_8602,N_7390,N_7826);
nor U8603 (N_8603,N_7705,N_7505);
nand U8604 (N_8604,N_7085,N_7962);
or U8605 (N_8605,N_7357,N_7016);
nand U8606 (N_8606,N_7063,N_7191);
or U8607 (N_8607,N_7295,N_7304);
and U8608 (N_8608,N_7753,N_7018);
and U8609 (N_8609,N_7030,N_7863);
nor U8610 (N_8610,N_7498,N_7683);
nand U8611 (N_8611,N_7547,N_7897);
or U8612 (N_8612,N_7956,N_7524);
and U8613 (N_8613,N_7366,N_7899);
and U8614 (N_8614,N_7554,N_7716);
nand U8615 (N_8615,N_7946,N_7112);
nand U8616 (N_8616,N_7824,N_7150);
and U8617 (N_8617,N_7558,N_7375);
and U8618 (N_8618,N_7911,N_7066);
nor U8619 (N_8619,N_7391,N_7837);
nand U8620 (N_8620,N_7112,N_7900);
or U8621 (N_8621,N_7074,N_7659);
nand U8622 (N_8622,N_7681,N_7782);
and U8623 (N_8623,N_7286,N_7222);
nor U8624 (N_8624,N_7944,N_7765);
nor U8625 (N_8625,N_7108,N_7202);
nand U8626 (N_8626,N_7007,N_7129);
and U8627 (N_8627,N_7662,N_7708);
nor U8628 (N_8628,N_7316,N_7896);
or U8629 (N_8629,N_7174,N_7851);
nand U8630 (N_8630,N_7575,N_7822);
and U8631 (N_8631,N_7745,N_7297);
and U8632 (N_8632,N_7792,N_7794);
or U8633 (N_8633,N_7165,N_7135);
and U8634 (N_8634,N_7003,N_7095);
nand U8635 (N_8635,N_7044,N_7863);
or U8636 (N_8636,N_7692,N_7839);
or U8637 (N_8637,N_7507,N_7548);
nand U8638 (N_8638,N_7994,N_7375);
nor U8639 (N_8639,N_7997,N_7400);
and U8640 (N_8640,N_7291,N_7377);
and U8641 (N_8641,N_7951,N_7461);
nor U8642 (N_8642,N_7248,N_7510);
or U8643 (N_8643,N_7217,N_7073);
and U8644 (N_8644,N_7814,N_7820);
nor U8645 (N_8645,N_7220,N_7868);
nor U8646 (N_8646,N_7771,N_7078);
nand U8647 (N_8647,N_7703,N_7848);
or U8648 (N_8648,N_7981,N_7038);
nor U8649 (N_8649,N_7471,N_7405);
and U8650 (N_8650,N_7984,N_7517);
and U8651 (N_8651,N_7404,N_7739);
nand U8652 (N_8652,N_7051,N_7104);
nand U8653 (N_8653,N_7178,N_7547);
nor U8654 (N_8654,N_7417,N_7840);
nand U8655 (N_8655,N_7923,N_7753);
nor U8656 (N_8656,N_7931,N_7151);
and U8657 (N_8657,N_7181,N_7793);
or U8658 (N_8658,N_7824,N_7661);
nand U8659 (N_8659,N_7115,N_7877);
or U8660 (N_8660,N_7632,N_7068);
and U8661 (N_8661,N_7408,N_7664);
nor U8662 (N_8662,N_7169,N_7708);
nand U8663 (N_8663,N_7490,N_7506);
or U8664 (N_8664,N_7494,N_7560);
nor U8665 (N_8665,N_7991,N_7431);
nand U8666 (N_8666,N_7654,N_7182);
nand U8667 (N_8667,N_7925,N_7096);
nand U8668 (N_8668,N_7008,N_7861);
or U8669 (N_8669,N_7268,N_7851);
or U8670 (N_8670,N_7919,N_7914);
nand U8671 (N_8671,N_7510,N_7417);
or U8672 (N_8672,N_7776,N_7893);
nand U8673 (N_8673,N_7138,N_7293);
nor U8674 (N_8674,N_7530,N_7901);
or U8675 (N_8675,N_7707,N_7155);
nand U8676 (N_8676,N_7495,N_7690);
and U8677 (N_8677,N_7510,N_7916);
nor U8678 (N_8678,N_7423,N_7207);
nand U8679 (N_8679,N_7251,N_7628);
or U8680 (N_8680,N_7350,N_7547);
and U8681 (N_8681,N_7113,N_7198);
nand U8682 (N_8682,N_7897,N_7703);
or U8683 (N_8683,N_7210,N_7091);
or U8684 (N_8684,N_7301,N_7353);
or U8685 (N_8685,N_7543,N_7127);
and U8686 (N_8686,N_7639,N_7084);
or U8687 (N_8687,N_7974,N_7154);
or U8688 (N_8688,N_7917,N_7980);
nand U8689 (N_8689,N_7001,N_7953);
and U8690 (N_8690,N_7942,N_7789);
nor U8691 (N_8691,N_7785,N_7715);
nor U8692 (N_8692,N_7672,N_7953);
nor U8693 (N_8693,N_7557,N_7803);
nor U8694 (N_8694,N_7795,N_7216);
nor U8695 (N_8695,N_7078,N_7526);
or U8696 (N_8696,N_7854,N_7249);
nand U8697 (N_8697,N_7703,N_7614);
nor U8698 (N_8698,N_7995,N_7229);
nor U8699 (N_8699,N_7430,N_7697);
or U8700 (N_8700,N_7755,N_7567);
nor U8701 (N_8701,N_7143,N_7131);
nor U8702 (N_8702,N_7679,N_7160);
nor U8703 (N_8703,N_7250,N_7555);
nand U8704 (N_8704,N_7980,N_7173);
or U8705 (N_8705,N_7675,N_7533);
nor U8706 (N_8706,N_7063,N_7423);
nand U8707 (N_8707,N_7648,N_7455);
and U8708 (N_8708,N_7471,N_7306);
and U8709 (N_8709,N_7568,N_7280);
and U8710 (N_8710,N_7542,N_7833);
and U8711 (N_8711,N_7795,N_7136);
xor U8712 (N_8712,N_7729,N_7348);
nand U8713 (N_8713,N_7146,N_7622);
and U8714 (N_8714,N_7191,N_7561);
or U8715 (N_8715,N_7496,N_7222);
nand U8716 (N_8716,N_7390,N_7766);
nor U8717 (N_8717,N_7112,N_7200);
nand U8718 (N_8718,N_7387,N_7629);
nand U8719 (N_8719,N_7949,N_7901);
nor U8720 (N_8720,N_7999,N_7055);
nand U8721 (N_8721,N_7799,N_7854);
and U8722 (N_8722,N_7489,N_7911);
and U8723 (N_8723,N_7648,N_7337);
and U8724 (N_8724,N_7601,N_7354);
nor U8725 (N_8725,N_7332,N_7410);
nand U8726 (N_8726,N_7354,N_7024);
nand U8727 (N_8727,N_7386,N_7134);
and U8728 (N_8728,N_7433,N_7270);
nor U8729 (N_8729,N_7356,N_7047);
nor U8730 (N_8730,N_7385,N_7643);
nand U8731 (N_8731,N_7670,N_7204);
and U8732 (N_8732,N_7888,N_7300);
and U8733 (N_8733,N_7862,N_7205);
nand U8734 (N_8734,N_7898,N_7637);
and U8735 (N_8735,N_7190,N_7778);
or U8736 (N_8736,N_7275,N_7343);
nand U8737 (N_8737,N_7993,N_7072);
nand U8738 (N_8738,N_7673,N_7622);
or U8739 (N_8739,N_7527,N_7263);
nor U8740 (N_8740,N_7094,N_7841);
and U8741 (N_8741,N_7766,N_7610);
nand U8742 (N_8742,N_7945,N_7318);
nand U8743 (N_8743,N_7445,N_7264);
or U8744 (N_8744,N_7160,N_7934);
and U8745 (N_8745,N_7826,N_7131);
nand U8746 (N_8746,N_7061,N_7680);
nor U8747 (N_8747,N_7471,N_7507);
nor U8748 (N_8748,N_7682,N_7366);
and U8749 (N_8749,N_7741,N_7174);
and U8750 (N_8750,N_7008,N_7641);
nor U8751 (N_8751,N_7249,N_7103);
nand U8752 (N_8752,N_7223,N_7981);
nor U8753 (N_8753,N_7270,N_7061);
and U8754 (N_8754,N_7649,N_7406);
or U8755 (N_8755,N_7983,N_7522);
and U8756 (N_8756,N_7774,N_7728);
xnor U8757 (N_8757,N_7048,N_7708);
nand U8758 (N_8758,N_7624,N_7506);
and U8759 (N_8759,N_7727,N_7161);
nand U8760 (N_8760,N_7660,N_7423);
and U8761 (N_8761,N_7009,N_7226);
and U8762 (N_8762,N_7841,N_7227);
and U8763 (N_8763,N_7550,N_7079);
nor U8764 (N_8764,N_7338,N_7822);
or U8765 (N_8765,N_7301,N_7125);
or U8766 (N_8766,N_7672,N_7030);
nor U8767 (N_8767,N_7765,N_7370);
or U8768 (N_8768,N_7940,N_7750);
nor U8769 (N_8769,N_7214,N_7310);
nor U8770 (N_8770,N_7162,N_7805);
nand U8771 (N_8771,N_7727,N_7802);
nand U8772 (N_8772,N_7968,N_7715);
nand U8773 (N_8773,N_7198,N_7760);
and U8774 (N_8774,N_7289,N_7146);
nand U8775 (N_8775,N_7214,N_7513);
nand U8776 (N_8776,N_7946,N_7869);
or U8777 (N_8777,N_7219,N_7590);
nor U8778 (N_8778,N_7962,N_7386);
nand U8779 (N_8779,N_7142,N_7530);
nor U8780 (N_8780,N_7499,N_7607);
nand U8781 (N_8781,N_7870,N_7002);
or U8782 (N_8782,N_7636,N_7345);
nand U8783 (N_8783,N_7160,N_7060);
nand U8784 (N_8784,N_7861,N_7729);
nand U8785 (N_8785,N_7899,N_7948);
and U8786 (N_8786,N_7527,N_7746);
nand U8787 (N_8787,N_7086,N_7258);
and U8788 (N_8788,N_7758,N_7490);
nor U8789 (N_8789,N_7889,N_7389);
nor U8790 (N_8790,N_7594,N_7412);
and U8791 (N_8791,N_7230,N_7452);
nand U8792 (N_8792,N_7962,N_7969);
or U8793 (N_8793,N_7492,N_7723);
or U8794 (N_8794,N_7950,N_7268);
and U8795 (N_8795,N_7413,N_7938);
nor U8796 (N_8796,N_7617,N_7934);
and U8797 (N_8797,N_7404,N_7866);
nand U8798 (N_8798,N_7569,N_7222);
nor U8799 (N_8799,N_7942,N_7409);
nand U8800 (N_8800,N_7848,N_7112);
nor U8801 (N_8801,N_7430,N_7053);
nand U8802 (N_8802,N_7797,N_7782);
nand U8803 (N_8803,N_7688,N_7960);
nor U8804 (N_8804,N_7156,N_7811);
or U8805 (N_8805,N_7774,N_7480);
nand U8806 (N_8806,N_7960,N_7829);
or U8807 (N_8807,N_7185,N_7446);
nand U8808 (N_8808,N_7035,N_7279);
and U8809 (N_8809,N_7055,N_7312);
or U8810 (N_8810,N_7619,N_7219);
nand U8811 (N_8811,N_7396,N_7730);
or U8812 (N_8812,N_7153,N_7493);
or U8813 (N_8813,N_7388,N_7058);
and U8814 (N_8814,N_7475,N_7737);
nor U8815 (N_8815,N_7437,N_7448);
nand U8816 (N_8816,N_7136,N_7053);
nor U8817 (N_8817,N_7075,N_7449);
or U8818 (N_8818,N_7082,N_7896);
and U8819 (N_8819,N_7477,N_7802);
nand U8820 (N_8820,N_7732,N_7343);
and U8821 (N_8821,N_7655,N_7119);
or U8822 (N_8822,N_7194,N_7639);
or U8823 (N_8823,N_7952,N_7707);
or U8824 (N_8824,N_7105,N_7600);
nor U8825 (N_8825,N_7428,N_7787);
nand U8826 (N_8826,N_7842,N_7383);
or U8827 (N_8827,N_7222,N_7919);
and U8828 (N_8828,N_7963,N_7097);
or U8829 (N_8829,N_7570,N_7230);
nor U8830 (N_8830,N_7915,N_7208);
nand U8831 (N_8831,N_7887,N_7480);
or U8832 (N_8832,N_7562,N_7909);
nor U8833 (N_8833,N_7288,N_7494);
or U8834 (N_8834,N_7155,N_7979);
nor U8835 (N_8835,N_7881,N_7165);
nand U8836 (N_8836,N_7344,N_7876);
and U8837 (N_8837,N_7898,N_7747);
nor U8838 (N_8838,N_7384,N_7999);
and U8839 (N_8839,N_7056,N_7651);
nand U8840 (N_8840,N_7495,N_7282);
or U8841 (N_8841,N_7813,N_7754);
nor U8842 (N_8842,N_7877,N_7669);
and U8843 (N_8843,N_7516,N_7547);
or U8844 (N_8844,N_7965,N_7910);
or U8845 (N_8845,N_7204,N_7615);
and U8846 (N_8846,N_7879,N_7034);
nand U8847 (N_8847,N_7219,N_7847);
nand U8848 (N_8848,N_7481,N_7730);
nor U8849 (N_8849,N_7977,N_7613);
and U8850 (N_8850,N_7849,N_7034);
or U8851 (N_8851,N_7636,N_7041);
nand U8852 (N_8852,N_7947,N_7794);
or U8853 (N_8853,N_7165,N_7651);
and U8854 (N_8854,N_7611,N_7239);
and U8855 (N_8855,N_7964,N_7826);
and U8856 (N_8856,N_7738,N_7056);
nor U8857 (N_8857,N_7586,N_7026);
or U8858 (N_8858,N_7572,N_7836);
nand U8859 (N_8859,N_7751,N_7498);
nor U8860 (N_8860,N_7372,N_7051);
or U8861 (N_8861,N_7707,N_7987);
nor U8862 (N_8862,N_7231,N_7167);
nand U8863 (N_8863,N_7787,N_7942);
or U8864 (N_8864,N_7194,N_7719);
or U8865 (N_8865,N_7017,N_7373);
nor U8866 (N_8866,N_7691,N_7672);
nor U8867 (N_8867,N_7931,N_7934);
nand U8868 (N_8868,N_7818,N_7572);
or U8869 (N_8869,N_7979,N_7585);
nand U8870 (N_8870,N_7960,N_7041);
nor U8871 (N_8871,N_7104,N_7287);
nand U8872 (N_8872,N_7294,N_7875);
nor U8873 (N_8873,N_7926,N_7090);
nand U8874 (N_8874,N_7396,N_7897);
and U8875 (N_8875,N_7774,N_7553);
and U8876 (N_8876,N_7172,N_7069);
nor U8877 (N_8877,N_7733,N_7568);
or U8878 (N_8878,N_7168,N_7735);
or U8879 (N_8879,N_7721,N_7278);
nand U8880 (N_8880,N_7663,N_7009);
and U8881 (N_8881,N_7758,N_7358);
or U8882 (N_8882,N_7063,N_7381);
and U8883 (N_8883,N_7940,N_7214);
or U8884 (N_8884,N_7297,N_7425);
or U8885 (N_8885,N_7461,N_7665);
or U8886 (N_8886,N_7769,N_7484);
nor U8887 (N_8887,N_7241,N_7297);
and U8888 (N_8888,N_7600,N_7986);
nor U8889 (N_8889,N_7119,N_7945);
nand U8890 (N_8890,N_7888,N_7786);
or U8891 (N_8891,N_7267,N_7171);
nor U8892 (N_8892,N_7154,N_7269);
nor U8893 (N_8893,N_7247,N_7633);
or U8894 (N_8894,N_7103,N_7750);
or U8895 (N_8895,N_7745,N_7130);
or U8896 (N_8896,N_7669,N_7933);
and U8897 (N_8897,N_7614,N_7256);
nand U8898 (N_8898,N_7367,N_7585);
and U8899 (N_8899,N_7725,N_7398);
or U8900 (N_8900,N_7849,N_7854);
or U8901 (N_8901,N_7216,N_7630);
nand U8902 (N_8902,N_7360,N_7768);
or U8903 (N_8903,N_7175,N_7355);
nand U8904 (N_8904,N_7593,N_7580);
nor U8905 (N_8905,N_7897,N_7967);
or U8906 (N_8906,N_7139,N_7641);
or U8907 (N_8907,N_7901,N_7555);
and U8908 (N_8908,N_7292,N_7261);
nand U8909 (N_8909,N_7175,N_7164);
or U8910 (N_8910,N_7467,N_7806);
nand U8911 (N_8911,N_7423,N_7123);
or U8912 (N_8912,N_7668,N_7817);
or U8913 (N_8913,N_7945,N_7905);
nand U8914 (N_8914,N_7590,N_7542);
xor U8915 (N_8915,N_7961,N_7785);
and U8916 (N_8916,N_7926,N_7977);
nand U8917 (N_8917,N_7756,N_7049);
or U8918 (N_8918,N_7570,N_7984);
nor U8919 (N_8919,N_7336,N_7250);
or U8920 (N_8920,N_7905,N_7552);
nand U8921 (N_8921,N_7254,N_7497);
xor U8922 (N_8922,N_7168,N_7146);
or U8923 (N_8923,N_7337,N_7861);
nand U8924 (N_8924,N_7965,N_7696);
nand U8925 (N_8925,N_7987,N_7705);
nor U8926 (N_8926,N_7929,N_7302);
and U8927 (N_8927,N_7428,N_7563);
or U8928 (N_8928,N_7225,N_7452);
or U8929 (N_8929,N_7832,N_7669);
and U8930 (N_8930,N_7807,N_7754);
nor U8931 (N_8931,N_7166,N_7210);
nor U8932 (N_8932,N_7421,N_7031);
and U8933 (N_8933,N_7284,N_7539);
and U8934 (N_8934,N_7314,N_7454);
and U8935 (N_8935,N_7841,N_7735);
or U8936 (N_8936,N_7803,N_7227);
and U8937 (N_8937,N_7245,N_7567);
or U8938 (N_8938,N_7610,N_7322);
nor U8939 (N_8939,N_7910,N_7082);
and U8940 (N_8940,N_7265,N_7122);
and U8941 (N_8941,N_7960,N_7679);
nor U8942 (N_8942,N_7534,N_7884);
nor U8943 (N_8943,N_7932,N_7416);
or U8944 (N_8944,N_7225,N_7078);
nor U8945 (N_8945,N_7174,N_7961);
or U8946 (N_8946,N_7209,N_7795);
or U8947 (N_8947,N_7540,N_7976);
nor U8948 (N_8948,N_7345,N_7722);
or U8949 (N_8949,N_7841,N_7843);
or U8950 (N_8950,N_7394,N_7722);
or U8951 (N_8951,N_7477,N_7807);
and U8952 (N_8952,N_7944,N_7990);
nand U8953 (N_8953,N_7668,N_7368);
or U8954 (N_8954,N_7535,N_7498);
xor U8955 (N_8955,N_7518,N_7960);
and U8956 (N_8956,N_7055,N_7342);
or U8957 (N_8957,N_7385,N_7476);
and U8958 (N_8958,N_7038,N_7617);
nor U8959 (N_8959,N_7651,N_7465);
nor U8960 (N_8960,N_7813,N_7322);
and U8961 (N_8961,N_7461,N_7673);
nand U8962 (N_8962,N_7116,N_7461);
and U8963 (N_8963,N_7326,N_7476);
and U8964 (N_8964,N_7889,N_7498);
nor U8965 (N_8965,N_7500,N_7532);
nand U8966 (N_8966,N_7903,N_7247);
or U8967 (N_8967,N_7330,N_7111);
nor U8968 (N_8968,N_7905,N_7459);
nand U8969 (N_8969,N_7725,N_7105);
nor U8970 (N_8970,N_7632,N_7160);
nand U8971 (N_8971,N_7465,N_7079);
nand U8972 (N_8972,N_7129,N_7273);
and U8973 (N_8973,N_7426,N_7286);
or U8974 (N_8974,N_7663,N_7085);
nand U8975 (N_8975,N_7848,N_7882);
and U8976 (N_8976,N_7327,N_7641);
nor U8977 (N_8977,N_7276,N_7658);
or U8978 (N_8978,N_7005,N_7582);
nor U8979 (N_8979,N_7105,N_7154);
or U8980 (N_8980,N_7071,N_7900);
nand U8981 (N_8981,N_7932,N_7640);
nand U8982 (N_8982,N_7880,N_7040);
or U8983 (N_8983,N_7636,N_7194);
nand U8984 (N_8984,N_7489,N_7233);
nor U8985 (N_8985,N_7095,N_7765);
nand U8986 (N_8986,N_7224,N_7444);
or U8987 (N_8987,N_7257,N_7809);
or U8988 (N_8988,N_7834,N_7012);
or U8989 (N_8989,N_7889,N_7345);
and U8990 (N_8990,N_7818,N_7561);
nand U8991 (N_8991,N_7863,N_7198);
or U8992 (N_8992,N_7535,N_7472);
or U8993 (N_8993,N_7413,N_7928);
or U8994 (N_8994,N_7975,N_7665);
or U8995 (N_8995,N_7229,N_7034);
nor U8996 (N_8996,N_7715,N_7931);
and U8997 (N_8997,N_7911,N_7393);
and U8998 (N_8998,N_7257,N_7315);
or U8999 (N_8999,N_7934,N_7001);
nor U9000 (N_9000,N_8506,N_8888);
and U9001 (N_9001,N_8213,N_8793);
nor U9002 (N_9002,N_8267,N_8776);
nand U9003 (N_9003,N_8202,N_8934);
or U9004 (N_9004,N_8984,N_8307);
and U9005 (N_9005,N_8653,N_8309);
nor U9006 (N_9006,N_8334,N_8559);
nand U9007 (N_9007,N_8060,N_8633);
or U9008 (N_9008,N_8374,N_8482);
nand U9009 (N_9009,N_8408,N_8567);
nand U9010 (N_9010,N_8388,N_8375);
or U9011 (N_9011,N_8448,N_8881);
nand U9012 (N_9012,N_8400,N_8150);
nor U9013 (N_9013,N_8623,N_8702);
and U9014 (N_9014,N_8657,N_8674);
and U9015 (N_9015,N_8279,N_8704);
or U9016 (N_9016,N_8049,N_8873);
nand U9017 (N_9017,N_8689,N_8666);
and U9018 (N_9018,N_8502,N_8092);
nand U9019 (N_9019,N_8869,N_8410);
or U9020 (N_9020,N_8921,N_8248);
and U9021 (N_9021,N_8014,N_8968);
or U9022 (N_9022,N_8350,N_8018);
nand U9023 (N_9023,N_8789,N_8361);
and U9024 (N_9024,N_8537,N_8211);
and U9025 (N_9025,N_8942,N_8097);
nand U9026 (N_9026,N_8056,N_8964);
or U9027 (N_9027,N_8719,N_8113);
or U9028 (N_9028,N_8883,N_8103);
nor U9029 (N_9029,N_8223,N_8868);
nand U9030 (N_9030,N_8333,N_8054);
nor U9031 (N_9031,N_8499,N_8855);
nor U9032 (N_9032,N_8144,N_8886);
and U9033 (N_9033,N_8534,N_8677);
nor U9034 (N_9034,N_8997,N_8458);
nor U9035 (N_9035,N_8960,N_8532);
and U9036 (N_9036,N_8165,N_8777);
nand U9037 (N_9037,N_8624,N_8336);
and U9038 (N_9038,N_8325,N_8008);
or U9039 (N_9039,N_8805,N_8221);
nand U9040 (N_9040,N_8667,N_8412);
and U9041 (N_9041,N_8194,N_8969);
or U9042 (N_9042,N_8076,N_8425);
nand U9043 (N_9043,N_8876,N_8987);
and U9044 (N_9044,N_8763,N_8439);
or U9045 (N_9045,N_8693,N_8233);
nor U9046 (N_9046,N_8580,N_8570);
and U9047 (N_9047,N_8321,N_8716);
nand U9048 (N_9048,N_8940,N_8906);
and U9049 (N_9049,N_8077,N_8440);
nor U9050 (N_9050,N_8038,N_8290);
nand U9051 (N_9051,N_8668,N_8444);
or U9052 (N_9052,N_8117,N_8293);
nand U9053 (N_9053,N_8685,N_8127);
nor U9054 (N_9054,N_8012,N_8265);
or U9055 (N_9055,N_8787,N_8630);
nand U9056 (N_9056,N_8414,N_8315);
nor U9057 (N_9057,N_8220,N_8814);
and U9058 (N_9058,N_8938,N_8579);
nor U9059 (N_9059,N_8671,N_8428);
or U9060 (N_9060,N_8149,N_8790);
and U9061 (N_9061,N_8151,N_8882);
nor U9062 (N_9062,N_8188,N_8652);
nor U9063 (N_9063,N_8714,N_8779);
nand U9064 (N_9064,N_8945,N_8919);
nand U9065 (N_9065,N_8295,N_8856);
nand U9066 (N_9066,N_8010,N_8759);
and U9067 (N_9067,N_8083,N_8650);
nor U9068 (N_9068,N_8470,N_8956);
or U9069 (N_9069,N_8516,N_8943);
nand U9070 (N_9070,N_8454,N_8132);
and U9071 (N_9071,N_8507,N_8746);
or U9072 (N_9072,N_8123,N_8583);
nor U9073 (N_9073,N_8420,N_8700);
nor U9074 (N_9074,N_8765,N_8898);
or U9075 (N_9075,N_8087,N_8550);
nand U9076 (N_9076,N_8783,N_8792);
nand U9077 (N_9077,N_8492,N_8398);
or U9078 (N_9078,N_8736,N_8187);
nand U9079 (N_9079,N_8015,N_8072);
or U9080 (N_9080,N_8246,N_8201);
nand U9081 (N_9081,N_8370,N_8781);
nor U9082 (N_9082,N_8493,N_8529);
and U9083 (N_9083,N_8585,N_8244);
nor U9084 (N_9084,N_8182,N_8903);
and U9085 (N_9085,N_8241,N_8118);
nor U9086 (N_9086,N_8287,N_8166);
nand U9087 (N_9087,N_8552,N_8939);
or U9088 (N_9088,N_8926,N_8277);
nand U9089 (N_9089,N_8344,N_8124);
nor U9090 (N_9090,N_8199,N_8638);
nand U9091 (N_9091,N_8933,N_8059);
or U9092 (N_9092,N_8218,N_8298);
or U9093 (N_9093,N_8718,N_8613);
nor U9094 (N_9094,N_8708,N_8864);
nor U9095 (N_9095,N_8498,N_8802);
nor U9096 (N_9096,N_8331,N_8270);
or U9097 (N_9097,N_8185,N_8680);
or U9098 (N_9098,N_8588,N_8356);
or U9099 (N_9099,N_8027,N_8542);
nand U9100 (N_9100,N_8831,N_8378);
nand U9101 (N_9101,N_8465,N_8706);
nor U9102 (N_9102,N_8067,N_8601);
or U9103 (N_9103,N_8569,N_8044);
nand U9104 (N_9104,N_8941,N_8462);
and U9105 (N_9105,N_8073,N_8819);
or U9106 (N_9106,N_8108,N_8197);
nand U9107 (N_9107,N_8691,N_8937);
and U9108 (N_9108,N_8701,N_8683);
and U9109 (N_9109,N_8639,N_8345);
nand U9110 (N_9110,N_8606,N_8399);
nand U9111 (N_9111,N_8730,N_8167);
or U9112 (N_9112,N_8100,N_8604);
or U9113 (N_9113,N_8810,N_8429);
or U9114 (N_9114,N_8391,N_8982);
nor U9115 (N_9115,N_8724,N_8477);
and U9116 (N_9116,N_8016,N_8426);
nand U9117 (N_9117,N_8446,N_8435);
or U9118 (N_9118,N_8139,N_8163);
or U9119 (N_9119,N_8406,N_8261);
nor U9120 (N_9120,N_8627,N_8026);
and U9121 (N_9121,N_8860,N_8929);
nand U9122 (N_9122,N_8091,N_8389);
nand U9123 (N_9123,N_8846,N_8515);
and U9124 (N_9124,N_8469,N_8324);
nor U9125 (N_9125,N_8705,N_8153);
and U9126 (N_9126,N_8467,N_8582);
or U9127 (N_9127,N_8296,N_8234);
nor U9128 (N_9128,N_8734,N_8184);
and U9129 (N_9129,N_8935,N_8335);
nor U9130 (N_9130,N_8847,N_8973);
and U9131 (N_9131,N_8803,N_8158);
or U9132 (N_9132,N_8670,N_8557);
and U9133 (N_9133,N_8208,N_8055);
nand U9134 (N_9134,N_8843,N_8093);
nor U9135 (N_9135,N_8731,N_8129);
nand U9136 (N_9136,N_8955,N_8541);
and U9137 (N_9137,N_8160,N_8602);
nor U9138 (N_9138,N_8180,N_8156);
and U9139 (N_9139,N_8824,N_8827);
nand U9140 (N_9140,N_8216,N_8382);
nor U9141 (N_9141,N_8033,N_8880);
or U9142 (N_9142,N_8205,N_8979);
xor U9143 (N_9143,N_8147,N_8319);
nand U9144 (N_9144,N_8249,N_8744);
nor U9145 (N_9145,N_8676,N_8312);
or U9146 (N_9146,N_8978,N_8751);
nor U9147 (N_9147,N_8082,N_8822);
and U9148 (N_9148,N_8256,N_8571);
or U9149 (N_9149,N_8183,N_8452);
and U9150 (N_9150,N_8795,N_8577);
xor U9151 (N_9151,N_8481,N_8480);
or U9152 (N_9152,N_8599,N_8584);
nand U9153 (N_9153,N_8707,N_8192);
or U9154 (N_9154,N_8917,N_8381);
and U9155 (N_9155,N_8999,N_8275);
xor U9156 (N_9156,N_8998,N_8057);
or U9157 (N_9157,N_8556,N_8696);
nand U9158 (N_9158,N_8005,N_8102);
or U9159 (N_9159,N_8517,N_8301);
nor U9160 (N_9160,N_8815,N_8423);
or U9161 (N_9161,N_8750,N_8817);
and U9162 (N_9162,N_8215,N_8304);
or U9163 (N_9163,N_8280,N_8581);
nor U9164 (N_9164,N_8145,N_8635);
or U9165 (N_9165,N_8871,N_8383);
or U9166 (N_9166,N_8445,N_8225);
nand U9167 (N_9167,N_8173,N_8189);
nand U9168 (N_9168,N_8514,N_8833);
or U9169 (N_9169,N_8314,N_8020);
or U9170 (N_9170,N_8046,N_8369);
or U9171 (N_9171,N_8832,N_8995);
nand U9172 (N_9172,N_8812,N_8434);
nand U9173 (N_9173,N_8755,N_8628);
xnor U9174 (N_9174,N_8954,N_8548);
and U9175 (N_9175,N_8328,N_8140);
nor U9176 (N_9176,N_8640,N_8258);
nor U9177 (N_9177,N_8340,N_8196);
nor U9178 (N_9178,N_8263,N_8608);
nor U9179 (N_9179,N_8422,N_8157);
or U9180 (N_9180,N_8840,N_8152);
and U9181 (N_9181,N_8713,N_8836);
nand U9182 (N_9182,N_8424,N_8901);
nand U9183 (N_9183,N_8566,N_8555);
or U9184 (N_9184,N_8828,N_8028);
nand U9185 (N_9185,N_8830,N_8456);
or U9186 (N_9186,N_8904,N_8593);
xor U9187 (N_9187,N_8509,N_8957);
nand U9188 (N_9188,N_8634,N_8510);
and U9189 (N_9189,N_8786,N_8587);
xnor U9190 (N_9190,N_8084,N_8379);
and U9191 (N_9191,N_8910,N_8154);
and U9192 (N_9192,N_8722,N_8308);
and U9193 (N_9193,N_8338,N_8226);
and U9194 (N_9194,N_8250,N_8455);
and U9195 (N_9195,N_8495,N_8808);
and U9196 (N_9196,N_8891,N_8266);
or U9197 (N_9197,N_8767,N_8339);
and U9198 (N_9198,N_8862,N_8362);
nor U9199 (N_9199,N_8743,N_8013);
or U9200 (N_9200,N_8141,N_8430);
nor U9201 (N_9201,N_8169,N_8447);
nor U9202 (N_9202,N_8521,N_8774);
nor U9203 (N_9203,N_8436,N_8981);
nor U9204 (N_9204,N_8519,N_8936);
nand U9205 (N_9205,N_8678,N_8944);
and U9206 (N_9206,N_8752,N_8992);
nor U9207 (N_9207,N_8172,N_8468);
nor U9208 (N_9208,N_8889,N_8007);
nand U9209 (N_9209,N_8130,N_8385);
and U9210 (N_9210,N_8377,N_8075);
nor U9211 (N_9211,N_8952,N_8190);
or U9212 (N_9212,N_8114,N_8665);
or U9213 (N_9213,N_8181,N_8897);
xnor U9214 (N_9214,N_8451,N_8051);
nand U9215 (N_9215,N_8159,N_8682);
and U9216 (N_9216,N_8659,N_8006);
xor U9217 (N_9217,N_8031,N_8273);
and U9218 (N_9218,N_8971,N_8053);
nor U9219 (N_9219,N_8745,N_8980);
or U9220 (N_9220,N_8305,N_8329);
nor U9221 (N_9221,N_8303,N_8487);
and U9222 (N_9222,N_8540,N_8632);
nor U9223 (N_9223,N_8065,N_8427);
or U9224 (N_9224,N_8850,N_8155);
nand U9225 (N_9225,N_8741,N_8648);
and U9226 (N_9226,N_8905,N_8642);
or U9227 (N_9227,N_8528,N_8255);
or U9228 (N_9228,N_8245,N_8484);
nor U9229 (N_9229,N_8526,N_8739);
or U9230 (N_9230,N_8863,N_8291);
nand U9231 (N_9231,N_8351,N_8219);
or U9232 (N_9232,N_8717,N_8923);
nand U9233 (N_9233,N_8254,N_8224);
nand U9234 (N_9234,N_8578,N_8967);
and U9235 (N_9235,N_8276,N_8186);
or U9236 (N_9236,N_8431,N_8364);
nand U9237 (N_9237,N_8035,N_8021);
nand U9238 (N_9238,N_8654,N_8094);
or U9239 (N_9239,N_8782,N_8384);
or U9240 (N_9240,N_8523,N_8829);
xor U9241 (N_9241,N_8457,N_8710);
or U9242 (N_9242,N_8620,N_8214);
nor U9243 (N_9243,N_8471,N_8317);
and U9244 (N_9244,N_8679,N_8925);
or U9245 (N_9245,N_8558,N_8212);
nor U9246 (N_9246,N_8614,N_8658);
and U9247 (N_9247,N_8848,N_8844);
nor U9248 (N_9248,N_8611,N_8721);
nand U9249 (N_9249,N_8081,N_8116);
nand U9250 (N_9250,N_8991,N_8994);
or U9251 (N_9251,N_8052,N_8066);
nand U9252 (N_9252,N_8612,N_8797);
or U9253 (N_9253,N_8373,N_8703);
or U9254 (N_9254,N_8209,N_8622);
and U9255 (N_9255,N_8545,N_8656);
nor U9256 (N_9256,N_8449,N_8965);
nand U9257 (N_9257,N_8358,N_8442);
nor U9258 (N_9258,N_8546,N_8775);
nor U9259 (N_9259,N_8547,N_8697);
and U9260 (N_9260,N_8915,N_8101);
nand U9261 (N_9261,N_8009,N_8040);
nand U9262 (N_9262,N_8788,N_8017);
and U9263 (N_9263,N_8737,N_8931);
nor U9264 (N_9264,N_8128,N_8441);
and U9265 (N_9265,N_8064,N_8958);
nand U9266 (N_9266,N_8095,N_8522);
or U9267 (N_9267,N_8762,N_8834);
or U9268 (N_9268,N_8918,N_8800);
nand U9269 (N_9269,N_8894,N_8003);
or U9270 (N_9270,N_8402,N_8404);
nand U9271 (N_9271,N_8643,N_8343);
and U9272 (N_9272,N_8306,N_8872);
and U9273 (N_9273,N_8845,N_8437);
nor U9274 (N_9274,N_8663,N_8433);
nand U9275 (N_9275,N_8753,N_8337);
nand U9276 (N_9276,N_8228,N_8371);
or U9277 (N_9277,N_8109,N_8088);
or U9278 (N_9278,N_8191,N_8323);
nand U9279 (N_9279,N_8394,N_8178);
nand U9280 (N_9280,N_8796,N_8176);
or U9281 (N_9281,N_8137,N_8136);
and U9282 (N_9282,N_8773,N_8951);
nor U9283 (N_9283,N_8047,N_8857);
or U9284 (N_9284,N_8911,N_8754);
or U9285 (N_9285,N_8791,N_8135);
nand U9286 (N_9286,N_8294,N_8625);
nand U9287 (N_9287,N_8988,N_8063);
or U9288 (N_9288,N_8518,N_8607);
nand U9289 (N_9289,N_8885,N_8207);
nand U9290 (N_9290,N_8924,N_8330);
or U9291 (N_9291,N_8948,N_8615);
or U9292 (N_9292,N_8576,N_8022);
or U9293 (N_9293,N_8177,N_8133);
nand U9294 (N_9294,N_8111,N_8074);
nand U9295 (N_9295,N_8393,N_8227);
nand U9296 (N_9296,N_8396,N_8596);
xnor U9297 (N_9297,N_8511,N_8970);
nor U9298 (N_9298,N_8148,N_8799);
and U9299 (N_9299,N_8242,N_8043);
nor U9300 (N_9300,N_8835,N_8080);
nand U9301 (N_9301,N_8645,N_8086);
and U9302 (N_9302,N_8501,N_8500);
nand U9303 (N_9303,N_8036,N_8210);
and U9304 (N_9304,N_8875,N_8839);
nand U9305 (N_9305,N_8974,N_8852);
and U9306 (N_9306,N_8568,N_8453);
nand U9307 (N_9307,N_8853,N_8669);
and U9308 (N_9308,N_8896,N_8479);
nand U9309 (N_9309,N_8461,N_8878);
nand U9310 (N_9310,N_8251,N_8977);
nand U9311 (N_9311,N_8575,N_8332);
and U9312 (N_9312,N_8616,N_8605);
and U9313 (N_9313,N_8297,N_8161);
nor U9314 (N_9314,N_8143,N_8617);
nand U9315 (N_9315,N_8972,N_8349);
nor U9316 (N_9316,N_8195,N_8825);
and U9317 (N_9317,N_8068,N_8784);
and U9318 (N_9318,N_8491,N_8748);
nor U9319 (N_9319,N_8203,N_8347);
nand U9320 (N_9320,N_8586,N_8125);
or U9321 (N_9321,N_8363,N_8694);
or U9322 (N_9322,N_8460,N_8895);
or U9323 (N_9323,N_8252,N_8079);
or U9324 (N_9324,N_8887,N_8646);
nor U9325 (N_9325,N_8818,N_8684);
or U9326 (N_9326,N_8728,N_8711);
and U9327 (N_9327,N_8747,N_8171);
nand U9328 (N_9328,N_8281,N_8284);
and U9329 (N_9329,N_8231,N_8908);
nor U9330 (N_9330,N_8473,N_8914);
and U9331 (N_9331,N_8078,N_8264);
and U9332 (N_9332,N_8342,N_8289);
or U9333 (N_9333,N_8572,N_8174);
and U9334 (N_9334,N_8070,N_8749);
or U9335 (N_9335,N_8168,N_8961);
nand U9336 (N_9336,N_8990,N_8866);
or U9337 (N_9337,N_8947,N_8397);
nor U9338 (N_9338,N_8692,N_8320);
nor U9339 (N_9339,N_8804,N_8346);
nor U9340 (N_9340,N_8041,N_8483);
nor U9341 (N_9341,N_8380,N_8771);
nand U9342 (N_9342,N_8574,N_8520);
nor U9343 (N_9343,N_8641,N_8912);
and U9344 (N_9344,N_8551,N_8235);
nand U9345 (N_9345,N_8348,N_8801);
nand U9346 (N_9346,N_8313,N_8681);
nand U9347 (N_9347,N_8772,N_8386);
and U9348 (N_9348,N_8727,N_8372);
or U9349 (N_9349,N_8411,N_8916);
nand U9350 (N_9350,N_8472,N_8401);
or U9351 (N_9351,N_8761,N_8989);
nand U9352 (N_9352,N_8239,N_8821);
nor U9353 (N_9353,N_8104,N_8354);
or U9354 (N_9354,N_8417,N_8024);
or U9355 (N_9355,N_8619,N_8131);
or U9356 (N_9356,N_8170,N_8061);
and U9357 (N_9357,N_8533,N_8352);
nand U9358 (N_9358,N_8950,N_8206);
or U9359 (N_9359,N_8976,N_8932);
and U9360 (N_9360,N_8413,N_8890);
xor U9361 (N_9361,N_8553,N_8770);
nor U9362 (N_9362,N_8816,N_8096);
or U9363 (N_9363,N_8664,N_8922);
nor U9364 (N_9364,N_8524,N_8403);
or U9365 (N_9365,N_8048,N_8565);
and U9366 (N_9366,N_8536,N_8419);
nand U9367 (N_9367,N_8310,N_8858);
nand U9368 (N_9368,N_8913,N_8563);
nor U9369 (N_9369,N_8288,N_8760);
nand U9370 (N_9370,N_8877,N_8900);
and U9371 (N_9371,N_8365,N_8134);
or U9372 (N_9372,N_8037,N_8806);
nand U9373 (N_9373,N_8610,N_8421);
nor U9374 (N_9374,N_8490,N_8661);
nor U9375 (N_9375,N_8660,N_8302);
nor U9376 (N_9376,N_8637,N_8766);
nor U9377 (N_9377,N_8841,N_8820);
or U9378 (N_9378,N_8268,N_8089);
and U9379 (N_9379,N_8278,N_8962);
nor U9380 (N_9380,N_8740,N_8723);
and U9381 (N_9381,N_8655,N_8311);
nand U9382 (N_9382,N_8709,N_8621);
and U9383 (N_9383,N_8376,N_8859);
or U9384 (N_9384,N_8949,N_8907);
nor U9385 (N_9385,N_8023,N_8164);
nor U9386 (N_9386,N_8230,N_8618);
nand U9387 (N_9387,N_8854,N_8497);
and U9388 (N_9388,N_8032,N_8042);
nor U9389 (N_9389,N_8513,N_8823);
or U9390 (N_9390,N_8318,N_8549);
and U9391 (N_9391,N_8651,N_8539);
or U9392 (N_9392,N_8757,N_8985);
or U9393 (N_9393,N_8649,N_8126);
and U9394 (N_9394,N_8395,N_8029);
nand U9395 (N_9395,N_8591,N_8699);
or U9396 (N_9396,N_8899,N_8930);
or U9397 (N_9397,N_8272,N_8243);
nor U9398 (N_9398,N_8418,N_8271);
nor U9399 (N_9399,N_8884,N_8626);
and U9400 (N_9400,N_8496,N_8690);
or U9401 (N_9401,N_8778,N_8769);
nor U9402 (N_9402,N_8341,N_8927);
or U9403 (N_9403,N_8756,N_8387);
or U9404 (N_9404,N_8715,N_8851);
nand U9405 (N_9405,N_8966,N_8368);
nand U9406 (N_9406,N_8920,N_8240);
nor U9407 (N_9407,N_8011,N_8768);
and U9408 (N_9408,N_8099,N_8867);
nor U9409 (N_9409,N_8438,N_8809);
nor U9410 (N_9410,N_8121,N_8554);
or U9411 (N_9411,N_8355,N_8098);
or U9412 (N_9412,N_8531,N_8030);
and U9413 (N_9413,N_8598,N_8001);
nand U9414 (N_9414,N_8508,N_8959);
and U9415 (N_9415,N_8459,N_8415);
or U9416 (N_9416,N_8636,N_8687);
or U9417 (N_9417,N_8589,N_8733);
and U9418 (N_9418,N_8780,N_8592);
and U9419 (N_9419,N_8726,N_8474);
or U9420 (N_9420,N_8909,N_8544);
and U9421 (N_9421,N_8476,N_8300);
or U9422 (N_9422,N_8292,N_8071);
nor U9423 (N_9423,N_8327,N_8409);
or U9424 (N_9424,N_8019,N_8198);
and U9425 (N_9425,N_8561,N_8600);
or U9426 (N_9426,N_8316,N_8179);
or U9427 (N_9427,N_8742,N_8735);
nor U9428 (N_9428,N_8902,N_8504);
nor U9429 (N_9429,N_8893,N_8257);
nand U9430 (N_9430,N_8259,N_8527);
nand U9431 (N_9431,N_8450,N_8603);
xnor U9432 (N_9432,N_8432,N_8486);
xor U9433 (N_9433,N_8720,N_8512);
or U9434 (N_9434,N_8120,N_8283);
and U9435 (N_9435,N_8253,N_8112);
or U9436 (N_9436,N_8353,N_8085);
nor U9437 (N_9437,N_8573,N_8861);
nand U9438 (N_9438,N_8050,N_8146);
and U9439 (N_9439,N_8996,N_8229);
nand U9440 (N_9440,N_8688,N_8002);
nand U9441 (N_9441,N_8237,N_8983);
nand U9442 (N_9442,N_8392,N_8590);
nor U9443 (N_9443,N_8672,N_8217);
nand U9444 (N_9444,N_8811,N_8986);
nor U9445 (N_9445,N_8758,N_8122);
nor U9446 (N_9446,N_8647,N_8115);
nand U9447 (N_9447,N_8946,N_8200);
nor U9448 (N_9448,N_8785,N_8838);
nor U9449 (N_9449,N_8090,N_8162);
or U9450 (N_9450,N_8119,N_8360);
nor U9451 (N_9451,N_8039,N_8466);
nor U9452 (N_9452,N_8000,N_8644);
nor U9453 (N_9453,N_8975,N_8738);
or U9454 (N_9454,N_8826,N_8874);
nor U9455 (N_9455,N_8069,N_8564);
and U9456 (N_9456,N_8106,N_8058);
or U9457 (N_9457,N_8142,N_8538);
or U9458 (N_9458,N_8475,N_8357);
nand U9459 (N_9459,N_8390,N_8807);
or U9460 (N_9460,N_8494,N_8594);
or U9461 (N_9461,N_8407,N_8928);
and U9462 (N_9462,N_8262,N_8204);
or U9463 (N_9463,N_8110,N_8963);
nor U9464 (N_9464,N_8485,N_8175);
nand U9465 (N_9465,N_8359,N_8629);
and U9466 (N_9466,N_8443,N_8543);
and U9467 (N_9467,N_8595,N_8236);
nor U9468 (N_9468,N_8597,N_8837);
nand U9469 (N_9469,N_8464,N_8562);
nor U9470 (N_9470,N_8138,N_8535);
nand U9471 (N_9471,N_8489,N_8695);
nor U9472 (N_9472,N_8794,N_8732);
nand U9473 (N_9473,N_8530,N_8260);
and U9474 (N_9474,N_8322,N_8503);
or U9475 (N_9475,N_8366,N_8367);
and U9476 (N_9476,N_8247,N_8865);
or U9477 (N_9477,N_8953,N_8892);
and U9478 (N_9478,N_8285,N_8045);
or U9479 (N_9479,N_8269,N_8870);
xor U9480 (N_9480,N_8193,N_8105);
nor U9481 (N_9481,N_8274,N_8405);
and U9482 (N_9482,N_8798,N_8560);
or U9483 (N_9483,N_8488,N_8686);
nor U9484 (N_9484,N_8673,N_8729);
nor U9485 (N_9485,N_8609,N_8662);
nand U9486 (N_9486,N_8107,N_8849);
nand U9487 (N_9487,N_8725,N_8282);
and U9488 (N_9488,N_8525,N_8463);
nand U9489 (N_9489,N_8238,N_8675);
nand U9490 (N_9490,N_8712,N_8004);
or U9491 (N_9491,N_8813,N_8879);
or U9492 (N_9492,N_8299,N_8416);
nor U9493 (N_9493,N_8062,N_8698);
or U9494 (N_9494,N_8993,N_8505);
and U9495 (N_9495,N_8326,N_8222);
nor U9496 (N_9496,N_8034,N_8478);
and U9497 (N_9497,N_8025,N_8842);
and U9498 (N_9498,N_8232,N_8764);
nor U9499 (N_9499,N_8631,N_8286);
nor U9500 (N_9500,N_8806,N_8846);
nand U9501 (N_9501,N_8644,N_8288);
nor U9502 (N_9502,N_8540,N_8509);
and U9503 (N_9503,N_8275,N_8862);
and U9504 (N_9504,N_8252,N_8284);
and U9505 (N_9505,N_8920,N_8449);
and U9506 (N_9506,N_8625,N_8770);
nand U9507 (N_9507,N_8283,N_8726);
and U9508 (N_9508,N_8578,N_8982);
or U9509 (N_9509,N_8509,N_8558);
and U9510 (N_9510,N_8541,N_8140);
nand U9511 (N_9511,N_8304,N_8850);
or U9512 (N_9512,N_8647,N_8204);
nand U9513 (N_9513,N_8435,N_8429);
or U9514 (N_9514,N_8127,N_8531);
or U9515 (N_9515,N_8323,N_8212);
and U9516 (N_9516,N_8468,N_8247);
or U9517 (N_9517,N_8332,N_8576);
and U9518 (N_9518,N_8344,N_8519);
or U9519 (N_9519,N_8771,N_8908);
or U9520 (N_9520,N_8178,N_8705);
nand U9521 (N_9521,N_8597,N_8701);
nor U9522 (N_9522,N_8538,N_8031);
or U9523 (N_9523,N_8711,N_8073);
and U9524 (N_9524,N_8491,N_8035);
nor U9525 (N_9525,N_8833,N_8868);
nand U9526 (N_9526,N_8836,N_8603);
nand U9527 (N_9527,N_8854,N_8710);
nor U9528 (N_9528,N_8745,N_8139);
and U9529 (N_9529,N_8091,N_8252);
and U9530 (N_9530,N_8877,N_8258);
nand U9531 (N_9531,N_8185,N_8208);
and U9532 (N_9532,N_8040,N_8055);
or U9533 (N_9533,N_8913,N_8947);
or U9534 (N_9534,N_8217,N_8847);
or U9535 (N_9535,N_8352,N_8412);
and U9536 (N_9536,N_8910,N_8898);
and U9537 (N_9537,N_8130,N_8956);
and U9538 (N_9538,N_8471,N_8239);
nor U9539 (N_9539,N_8794,N_8757);
and U9540 (N_9540,N_8910,N_8132);
nor U9541 (N_9541,N_8772,N_8866);
nand U9542 (N_9542,N_8910,N_8367);
and U9543 (N_9543,N_8932,N_8617);
or U9544 (N_9544,N_8270,N_8486);
nand U9545 (N_9545,N_8600,N_8092);
and U9546 (N_9546,N_8160,N_8620);
nand U9547 (N_9547,N_8947,N_8061);
or U9548 (N_9548,N_8703,N_8337);
nand U9549 (N_9549,N_8739,N_8568);
nand U9550 (N_9550,N_8052,N_8502);
nor U9551 (N_9551,N_8024,N_8914);
or U9552 (N_9552,N_8870,N_8382);
or U9553 (N_9553,N_8506,N_8443);
or U9554 (N_9554,N_8943,N_8974);
nor U9555 (N_9555,N_8192,N_8329);
or U9556 (N_9556,N_8074,N_8241);
or U9557 (N_9557,N_8539,N_8806);
nand U9558 (N_9558,N_8821,N_8709);
and U9559 (N_9559,N_8153,N_8947);
or U9560 (N_9560,N_8453,N_8488);
nand U9561 (N_9561,N_8787,N_8805);
nor U9562 (N_9562,N_8682,N_8063);
nand U9563 (N_9563,N_8584,N_8016);
nor U9564 (N_9564,N_8238,N_8604);
nor U9565 (N_9565,N_8691,N_8013);
nand U9566 (N_9566,N_8414,N_8385);
and U9567 (N_9567,N_8434,N_8679);
and U9568 (N_9568,N_8468,N_8444);
nand U9569 (N_9569,N_8001,N_8512);
or U9570 (N_9570,N_8882,N_8319);
xnor U9571 (N_9571,N_8167,N_8479);
or U9572 (N_9572,N_8191,N_8117);
and U9573 (N_9573,N_8216,N_8723);
and U9574 (N_9574,N_8214,N_8927);
or U9575 (N_9575,N_8781,N_8517);
and U9576 (N_9576,N_8633,N_8557);
nand U9577 (N_9577,N_8336,N_8038);
nand U9578 (N_9578,N_8662,N_8022);
and U9579 (N_9579,N_8318,N_8452);
nand U9580 (N_9580,N_8429,N_8185);
nor U9581 (N_9581,N_8172,N_8114);
or U9582 (N_9582,N_8544,N_8575);
and U9583 (N_9583,N_8749,N_8576);
nand U9584 (N_9584,N_8918,N_8231);
xor U9585 (N_9585,N_8291,N_8613);
nand U9586 (N_9586,N_8240,N_8545);
or U9587 (N_9587,N_8520,N_8653);
and U9588 (N_9588,N_8747,N_8694);
nand U9589 (N_9589,N_8938,N_8915);
nor U9590 (N_9590,N_8261,N_8762);
or U9591 (N_9591,N_8483,N_8338);
nand U9592 (N_9592,N_8142,N_8422);
nand U9593 (N_9593,N_8678,N_8609);
nor U9594 (N_9594,N_8138,N_8897);
and U9595 (N_9595,N_8983,N_8127);
nand U9596 (N_9596,N_8483,N_8203);
or U9597 (N_9597,N_8003,N_8209);
or U9598 (N_9598,N_8350,N_8443);
and U9599 (N_9599,N_8429,N_8046);
or U9600 (N_9600,N_8279,N_8431);
nand U9601 (N_9601,N_8756,N_8700);
or U9602 (N_9602,N_8442,N_8975);
and U9603 (N_9603,N_8532,N_8353);
or U9604 (N_9604,N_8358,N_8255);
nand U9605 (N_9605,N_8169,N_8659);
or U9606 (N_9606,N_8900,N_8716);
nor U9607 (N_9607,N_8380,N_8851);
nor U9608 (N_9608,N_8850,N_8827);
and U9609 (N_9609,N_8126,N_8008);
nor U9610 (N_9610,N_8401,N_8072);
or U9611 (N_9611,N_8301,N_8594);
nor U9612 (N_9612,N_8580,N_8605);
nor U9613 (N_9613,N_8810,N_8084);
or U9614 (N_9614,N_8440,N_8128);
nand U9615 (N_9615,N_8699,N_8566);
or U9616 (N_9616,N_8326,N_8848);
nand U9617 (N_9617,N_8479,N_8104);
or U9618 (N_9618,N_8982,N_8741);
or U9619 (N_9619,N_8307,N_8417);
or U9620 (N_9620,N_8397,N_8223);
or U9621 (N_9621,N_8911,N_8475);
and U9622 (N_9622,N_8640,N_8977);
or U9623 (N_9623,N_8104,N_8274);
or U9624 (N_9624,N_8307,N_8435);
nand U9625 (N_9625,N_8038,N_8660);
or U9626 (N_9626,N_8946,N_8965);
or U9627 (N_9627,N_8577,N_8047);
nand U9628 (N_9628,N_8975,N_8521);
nor U9629 (N_9629,N_8375,N_8549);
nor U9630 (N_9630,N_8906,N_8571);
nor U9631 (N_9631,N_8213,N_8647);
nand U9632 (N_9632,N_8780,N_8525);
nor U9633 (N_9633,N_8656,N_8099);
and U9634 (N_9634,N_8878,N_8767);
nor U9635 (N_9635,N_8171,N_8198);
or U9636 (N_9636,N_8789,N_8137);
or U9637 (N_9637,N_8736,N_8366);
nand U9638 (N_9638,N_8157,N_8642);
nand U9639 (N_9639,N_8590,N_8422);
nand U9640 (N_9640,N_8543,N_8261);
nand U9641 (N_9641,N_8101,N_8761);
and U9642 (N_9642,N_8434,N_8840);
or U9643 (N_9643,N_8699,N_8043);
nand U9644 (N_9644,N_8974,N_8277);
nor U9645 (N_9645,N_8516,N_8473);
nand U9646 (N_9646,N_8067,N_8464);
nand U9647 (N_9647,N_8494,N_8935);
nor U9648 (N_9648,N_8214,N_8898);
or U9649 (N_9649,N_8913,N_8283);
and U9650 (N_9650,N_8353,N_8974);
and U9651 (N_9651,N_8396,N_8056);
and U9652 (N_9652,N_8298,N_8642);
nand U9653 (N_9653,N_8569,N_8745);
and U9654 (N_9654,N_8334,N_8155);
or U9655 (N_9655,N_8432,N_8146);
nand U9656 (N_9656,N_8916,N_8978);
nor U9657 (N_9657,N_8588,N_8983);
nand U9658 (N_9658,N_8933,N_8325);
nor U9659 (N_9659,N_8667,N_8542);
nor U9660 (N_9660,N_8053,N_8480);
and U9661 (N_9661,N_8887,N_8653);
nor U9662 (N_9662,N_8170,N_8190);
or U9663 (N_9663,N_8114,N_8696);
and U9664 (N_9664,N_8056,N_8511);
nand U9665 (N_9665,N_8067,N_8904);
and U9666 (N_9666,N_8016,N_8225);
or U9667 (N_9667,N_8878,N_8164);
and U9668 (N_9668,N_8184,N_8312);
or U9669 (N_9669,N_8242,N_8545);
nor U9670 (N_9670,N_8441,N_8768);
nor U9671 (N_9671,N_8921,N_8849);
and U9672 (N_9672,N_8791,N_8542);
or U9673 (N_9673,N_8646,N_8787);
nand U9674 (N_9674,N_8214,N_8849);
nor U9675 (N_9675,N_8639,N_8112);
and U9676 (N_9676,N_8162,N_8004);
nand U9677 (N_9677,N_8556,N_8552);
nand U9678 (N_9678,N_8073,N_8445);
and U9679 (N_9679,N_8108,N_8500);
and U9680 (N_9680,N_8134,N_8472);
and U9681 (N_9681,N_8260,N_8746);
or U9682 (N_9682,N_8874,N_8149);
nor U9683 (N_9683,N_8240,N_8661);
or U9684 (N_9684,N_8018,N_8360);
xor U9685 (N_9685,N_8136,N_8365);
nand U9686 (N_9686,N_8108,N_8405);
or U9687 (N_9687,N_8421,N_8765);
nor U9688 (N_9688,N_8485,N_8267);
or U9689 (N_9689,N_8123,N_8644);
or U9690 (N_9690,N_8434,N_8049);
nand U9691 (N_9691,N_8543,N_8822);
nand U9692 (N_9692,N_8970,N_8726);
and U9693 (N_9693,N_8976,N_8333);
nor U9694 (N_9694,N_8068,N_8755);
nor U9695 (N_9695,N_8649,N_8262);
or U9696 (N_9696,N_8714,N_8482);
or U9697 (N_9697,N_8132,N_8517);
nor U9698 (N_9698,N_8394,N_8596);
xor U9699 (N_9699,N_8445,N_8492);
and U9700 (N_9700,N_8508,N_8122);
nand U9701 (N_9701,N_8824,N_8612);
and U9702 (N_9702,N_8142,N_8280);
xnor U9703 (N_9703,N_8017,N_8494);
nand U9704 (N_9704,N_8202,N_8312);
or U9705 (N_9705,N_8371,N_8668);
or U9706 (N_9706,N_8183,N_8738);
nor U9707 (N_9707,N_8244,N_8678);
nand U9708 (N_9708,N_8932,N_8425);
nand U9709 (N_9709,N_8392,N_8670);
or U9710 (N_9710,N_8385,N_8975);
and U9711 (N_9711,N_8553,N_8098);
or U9712 (N_9712,N_8558,N_8498);
or U9713 (N_9713,N_8523,N_8300);
and U9714 (N_9714,N_8667,N_8012);
and U9715 (N_9715,N_8463,N_8435);
nand U9716 (N_9716,N_8960,N_8922);
nor U9717 (N_9717,N_8125,N_8306);
or U9718 (N_9718,N_8207,N_8806);
or U9719 (N_9719,N_8245,N_8365);
or U9720 (N_9720,N_8973,N_8083);
or U9721 (N_9721,N_8547,N_8287);
nor U9722 (N_9722,N_8858,N_8416);
nor U9723 (N_9723,N_8915,N_8110);
nand U9724 (N_9724,N_8077,N_8254);
or U9725 (N_9725,N_8590,N_8676);
or U9726 (N_9726,N_8281,N_8202);
and U9727 (N_9727,N_8056,N_8680);
and U9728 (N_9728,N_8234,N_8406);
or U9729 (N_9729,N_8495,N_8802);
nor U9730 (N_9730,N_8585,N_8300);
nand U9731 (N_9731,N_8756,N_8755);
or U9732 (N_9732,N_8317,N_8925);
nor U9733 (N_9733,N_8608,N_8875);
nand U9734 (N_9734,N_8941,N_8082);
nand U9735 (N_9735,N_8947,N_8123);
nor U9736 (N_9736,N_8592,N_8572);
nor U9737 (N_9737,N_8189,N_8828);
or U9738 (N_9738,N_8429,N_8651);
nand U9739 (N_9739,N_8422,N_8003);
nor U9740 (N_9740,N_8646,N_8254);
nor U9741 (N_9741,N_8380,N_8782);
and U9742 (N_9742,N_8603,N_8068);
nand U9743 (N_9743,N_8283,N_8947);
or U9744 (N_9744,N_8569,N_8466);
or U9745 (N_9745,N_8039,N_8907);
nand U9746 (N_9746,N_8776,N_8270);
and U9747 (N_9747,N_8750,N_8920);
and U9748 (N_9748,N_8519,N_8780);
or U9749 (N_9749,N_8188,N_8844);
and U9750 (N_9750,N_8758,N_8494);
xnor U9751 (N_9751,N_8591,N_8864);
nor U9752 (N_9752,N_8744,N_8634);
nand U9753 (N_9753,N_8548,N_8692);
nor U9754 (N_9754,N_8822,N_8550);
and U9755 (N_9755,N_8458,N_8741);
nor U9756 (N_9756,N_8369,N_8498);
or U9757 (N_9757,N_8271,N_8180);
or U9758 (N_9758,N_8330,N_8146);
nand U9759 (N_9759,N_8265,N_8619);
nand U9760 (N_9760,N_8976,N_8677);
nand U9761 (N_9761,N_8706,N_8749);
and U9762 (N_9762,N_8941,N_8253);
nand U9763 (N_9763,N_8329,N_8051);
or U9764 (N_9764,N_8407,N_8560);
and U9765 (N_9765,N_8747,N_8101);
nor U9766 (N_9766,N_8807,N_8583);
and U9767 (N_9767,N_8840,N_8824);
or U9768 (N_9768,N_8855,N_8028);
nand U9769 (N_9769,N_8958,N_8662);
nor U9770 (N_9770,N_8844,N_8386);
or U9771 (N_9771,N_8209,N_8018);
nand U9772 (N_9772,N_8434,N_8536);
nor U9773 (N_9773,N_8611,N_8307);
and U9774 (N_9774,N_8765,N_8953);
nor U9775 (N_9775,N_8860,N_8252);
or U9776 (N_9776,N_8710,N_8246);
or U9777 (N_9777,N_8452,N_8613);
nand U9778 (N_9778,N_8441,N_8189);
or U9779 (N_9779,N_8197,N_8146);
nor U9780 (N_9780,N_8647,N_8456);
and U9781 (N_9781,N_8073,N_8002);
nand U9782 (N_9782,N_8338,N_8579);
and U9783 (N_9783,N_8219,N_8933);
or U9784 (N_9784,N_8291,N_8554);
or U9785 (N_9785,N_8386,N_8311);
nand U9786 (N_9786,N_8586,N_8614);
and U9787 (N_9787,N_8245,N_8169);
nand U9788 (N_9788,N_8492,N_8738);
nand U9789 (N_9789,N_8927,N_8675);
or U9790 (N_9790,N_8867,N_8726);
nor U9791 (N_9791,N_8686,N_8074);
and U9792 (N_9792,N_8511,N_8231);
or U9793 (N_9793,N_8323,N_8711);
and U9794 (N_9794,N_8391,N_8823);
nand U9795 (N_9795,N_8874,N_8314);
nand U9796 (N_9796,N_8004,N_8054);
nand U9797 (N_9797,N_8085,N_8007);
or U9798 (N_9798,N_8063,N_8568);
or U9799 (N_9799,N_8631,N_8920);
and U9800 (N_9800,N_8057,N_8875);
and U9801 (N_9801,N_8479,N_8252);
nor U9802 (N_9802,N_8383,N_8376);
nor U9803 (N_9803,N_8398,N_8286);
nor U9804 (N_9804,N_8179,N_8126);
nor U9805 (N_9805,N_8435,N_8221);
nand U9806 (N_9806,N_8429,N_8101);
or U9807 (N_9807,N_8681,N_8489);
or U9808 (N_9808,N_8339,N_8134);
nor U9809 (N_9809,N_8290,N_8137);
xnor U9810 (N_9810,N_8894,N_8690);
or U9811 (N_9811,N_8520,N_8426);
or U9812 (N_9812,N_8380,N_8859);
or U9813 (N_9813,N_8840,N_8210);
nand U9814 (N_9814,N_8119,N_8103);
nand U9815 (N_9815,N_8340,N_8165);
or U9816 (N_9816,N_8698,N_8959);
and U9817 (N_9817,N_8155,N_8091);
and U9818 (N_9818,N_8686,N_8145);
and U9819 (N_9819,N_8413,N_8471);
nand U9820 (N_9820,N_8760,N_8134);
nand U9821 (N_9821,N_8109,N_8851);
nand U9822 (N_9822,N_8123,N_8454);
and U9823 (N_9823,N_8066,N_8299);
nand U9824 (N_9824,N_8403,N_8659);
or U9825 (N_9825,N_8895,N_8504);
and U9826 (N_9826,N_8061,N_8702);
nand U9827 (N_9827,N_8679,N_8078);
or U9828 (N_9828,N_8250,N_8644);
nor U9829 (N_9829,N_8913,N_8688);
and U9830 (N_9830,N_8279,N_8273);
or U9831 (N_9831,N_8288,N_8525);
and U9832 (N_9832,N_8824,N_8467);
and U9833 (N_9833,N_8767,N_8178);
and U9834 (N_9834,N_8819,N_8147);
xnor U9835 (N_9835,N_8093,N_8871);
nor U9836 (N_9836,N_8630,N_8925);
or U9837 (N_9837,N_8973,N_8446);
and U9838 (N_9838,N_8773,N_8441);
nand U9839 (N_9839,N_8519,N_8433);
nor U9840 (N_9840,N_8948,N_8684);
and U9841 (N_9841,N_8228,N_8100);
and U9842 (N_9842,N_8136,N_8768);
nor U9843 (N_9843,N_8674,N_8921);
nand U9844 (N_9844,N_8018,N_8015);
and U9845 (N_9845,N_8945,N_8371);
and U9846 (N_9846,N_8096,N_8486);
and U9847 (N_9847,N_8344,N_8504);
or U9848 (N_9848,N_8167,N_8809);
nor U9849 (N_9849,N_8724,N_8297);
nor U9850 (N_9850,N_8462,N_8685);
nor U9851 (N_9851,N_8184,N_8886);
and U9852 (N_9852,N_8365,N_8994);
or U9853 (N_9853,N_8394,N_8857);
nor U9854 (N_9854,N_8901,N_8452);
and U9855 (N_9855,N_8071,N_8861);
nand U9856 (N_9856,N_8915,N_8077);
or U9857 (N_9857,N_8084,N_8671);
and U9858 (N_9858,N_8679,N_8416);
nor U9859 (N_9859,N_8233,N_8306);
or U9860 (N_9860,N_8407,N_8648);
or U9861 (N_9861,N_8177,N_8750);
nand U9862 (N_9862,N_8030,N_8829);
nand U9863 (N_9863,N_8055,N_8621);
nor U9864 (N_9864,N_8671,N_8893);
nor U9865 (N_9865,N_8102,N_8728);
nor U9866 (N_9866,N_8786,N_8610);
and U9867 (N_9867,N_8796,N_8213);
nor U9868 (N_9868,N_8035,N_8464);
nor U9869 (N_9869,N_8691,N_8712);
nor U9870 (N_9870,N_8306,N_8608);
nand U9871 (N_9871,N_8740,N_8539);
or U9872 (N_9872,N_8170,N_8615);
nor U9873 (N_9873,N_8126,N_8504);
and U9874 (N_9874,N_8925,N_8936);
nand U9875 (N_9875,N_8637,N_8411);
or U9876 (N_9876,N_8726,N_8100);
nor U9877 (N_9877,N_8248,N_8182);
or U9878 (N_9878,N_8139,N_8983);
and U9879 (N_9879,N_8800,N_8321);
and U9880 (N_9880,N_8167,N_8457);
nor U9881 (N_9881,N_8743,N_8069);
or U9882 (N_9882,N_8640,N_8023);
nor U9883 (N_9883,N_8930,N_8129);
nor U9884 (N_9884,N_8424,N_8839);
nor U9885 (N_9885,N_8402,N_8277);
nand U9886 (N_9886,N_8907,N_8448);
or U9887 (N_9887,N_8759,N_8669);
nor U9888 (N_9888,N_8597,N_8447);
and U9889 (N_9889,N_8533,N_8291);
or U9890 (N_9890,N_8270,N_8332);
nor U9891 (N_9891,N_8494,N_8727);
nor U9892 (N_9892,N_8638,N_8479);
nor U9893 (N_9893,N_8983,N_8404);
and U9894 (N_9894,N_8302,N_8943);
nor U9895 (N_9895,N_8374,N_8383);
nand U9896 (N_9896,N_8138,N_8730);
or U9897 (N_9897,N_8670,N_8100);
nor U9898 (N_9898,N_8131,N_8590);
xnor U9899 (N_9899,N_8079,N_8189);
or U9900 (N_9900,N_8669,N_8533);
nor U9901 (N_9901,N_8744,N_8772);
and U9902 (N_9902,N_8701,N_8061);
nor U9903 (N_9903,N_8712,N_8095);
nor U9904 (N_9904,N_8347,N_8074);
and U9905 (N_9905,N_8640,N_8423);
and U9906 (N_9906,N_8827,N_8029);
nor U9907 (N_9907,N_8963,N_8526);
or U9908 (N_9908,N_8913,N_8706);
nor U9909 (N_9909,N_8252,N_8247);
or U9910 (N_9910,N_8330,N_8056);
or U9911 (N_9911,N_8150,N_8369);
nor U9912 (N_9912,N_8229,N_8752);
or U9913 (N_9913,N_8966,N_8267);
and U9914 (N_9914,N_8709,N_8488);
or U9915 (N_9915,N_8611,N_8546);
or U9916 (N_9916,N_8405,N_8523);
or U9917 (N_9917,N_8510,N_8218);
and U9918 (N_9918,N_8777,N_8919);
nand U9919 (N_9919,N_8928,N_8330);
nor U9920 (N_9920,N_8420,N_8455);
nor U9921 (N_9921,N_8342,N_8133);
or U9922 (N_9922,N_8945,N_8765);
or U9923 (N_9923,N_8413,N_8816);
nand U9924 (N_9924,N_8796,N_8788);
nor U9925 (N_9925,N_8315,N_8279);
or U9926 (N_9926,N_8828,N_8165);
nor U9927 (N_9927,N_8870,N_8144);
xor U9928 (N_9928,N_8342,N_8643);
or U9929 (N_9929,N_8860,N_8745);
and U9930 (N_9930,N_8367,N_8442);
nor U9931 (N_9931,N_8074,N_8129);
nor U9932 (N_9932,N_8228,N_8323);
and U9933 (N_9933,N_8340,N_8679);
nor U9934 (N_9934,N_8277,N_8293);
or U9935 (N_9935,N_8072,N_8275);
nor U9936 (N_9936,N_8645,N_8540);
or U9937 (N_9937,N_8853,N_8332);
or U9938 (N_9938,N_8176,N_8412);
nand U9939 (N_9939,N_8027,N_8111);
or U9940 (N_9940,N_8270,N_8555);
and U9941 (N_9941,N_8847,N_8061);
and U9942 (N_9942,N_8501,N_8228);
nor U9943 (N_9943,N_8563,N_8838);
and U9944 (N_9944,N_8086,N_8275);
nor U9945 (N_9945,N_8648,N_8805);
or U9946 (N_9946,N_8150,N_8292);
or U9947 (N_9947,N_8684,N_8517);
or U9948 (N_9948,N_8161,N_8992);
or U9949 (N_9949,N_8937,N_8466);
or U9950 (N_9950,N_8593,N_8938);
nor U9951 (N_9951,N_8752,N_8179);
nor U9952 (N_9952,N_8109,N_8541);
and U9953 (N_9953,N_8851,N_8659);
and U9954 (N_9954,N_8745,N_8897);
nor U9955 (N_9955,N_8642,N_8450);
nor U9956 (N_9956,N_8707,N_8615);
and U9957 (N_9957,N_8623,N_8848);
nor U9958 (N_9958,N_8784,N_8361);
and U9959 (N_9959,N_8176,N_8718);
nor U9960 (N_9960,N_8085,N_8465);
or U9961 (N_9961,N_8639,N_8362);
nand U9962 (N_9962,N_8632,N_8239);
nand U9963 (N_9963,N_8697,N_8567);
nor U9964 (N_9964,N_8837,N_8217);
nand U9965 (N_9965,N_8800,N_8749);
nor U9966 (N_9966,N_8803,N_8945);
nor U9967 (N_9967,N_8817,N_8793);
and U9968 (N_9968,N_8578,N_8733);
nand U9969 (N_9969,N_8578,N_8245);
nand U9970 (N_9970,N_8291,N_8497);
nor U9971 (N_9971,N_8521,N_8702);
or U9972 (N_9972,N_8390,N_8861);
nand U9973 (N_9973,N_8375,N_8927);
or U9974 (N_9974,N_8909,N_8249);
nor U9975 (N_9975,N_8692,N_8308);
nand U9976 (N_9976,N_8046,N_8057);
and U9977 (N_9977,N_8369,N_8739);
nor U9978 (N_9978,N_8094,N_8889);
nand U9979 (N_9979,N_8217,N_8091);
nor U9980 (N_9980,N_8632,N_8286);
and U9981 (N_9981,N_8678,N_8725);
nand U9982 (N_9982,N_8609,N_8344);
and U9983 (N_9983,N_8213,N_8403);
and U9984 (N_9984,N_8040,N_8015);
nor U9985 (N_9985,N_8476,N_8474);
nand U9986 (N_9986,N_8870,N_8446);
and U9987 (N_9987,N_8736,N_8944);
and U9988 (N_9988,N_8630,N_8872);
and U9989 (N_9989,N_8849,N_8524);
nand U9990 (N_9990,N_8193,N_8571);
xnor U9991 (N_9991,N_8977,N_8901);
nand U9992 (N_9992,N_8959,N_8759);
and U9993 (N_9993,N_8363,N_8964);
or U9994 (N_9994,N_8407,N_8894);
nor U9995 (N_9995,N_8935,N_8970);
nand U9996 (N_9996,N_8552,N_8518);
nor U9997 (N_9997,N_8801,N_8364);
or U9998 (N_9998,N_8245,N_8273);
nor U9999 (N_9999,N_8228,N_8169);
nand UO_0 (O_0,N_9747,N_9331);
and UO_1 (O_1,N_9300,N_9072);
and UO_2 (O_2,N_9507,N_9479);
or UO_3 (O_3,N_9898,N_9235);
or UO_4 (O_4,N_9208,N_9036);
nand UO_5 (O_5,N_9639,N_9729);
and UO_6 (O_6,N_9324,N_9715);
and UO_7 (O_7,N_9003,N_9238);
and UO_8 (O_8,N_9470,N_9179);
nand UO_9 (O_9,N_9708,N_9837);
and UO_10 (O_10,N_9304,N_9906);
or UO_11 (O_11,N_9123,N_9915);
or UO_12 (O_12,N_9356,N_9981);
nand UO_13 (O_13,N_9372,N_9600);
nor UO_14 (O_14,N_9537,N_9211);
and UO_15 (O_15,N_9969,N_9526);
nor UO_16 (O_16,N_9484,N_9261);
nand UO_17 (O_17,N_9416,N_9452);
and UO_18 (O_18,N_9277,N_9247);
nor UO_19 (O_19,N_9485,N_9571);
nand UO_20 (O_20,N_9978,N_9861);
nand UO_21 (O_21,N_9840,N_9750);
nor UO_22 (O_22,N_9045,N_9189);
nor UO_23 (O_23,N_9995,N_9174);
nor UO_24 (O_24,N_9017,N_9332);
and UO_25 (O_25,N_9946,N_9581);
nor UO_26 (O_26,N_9051,N_9401);
nand UO_27 (O_27,N_9895,N_9322);
nand UO_28 (O_28,N_9568,N_9472);
or UO_29 (O_29,N_9585,N_9027);
nor UO_30 (O_30,N_9628,N_9414);
or UO_31 (O_31,N_9904,N_9831);
nand UO_32 (O_32,N_9403,N_9949);
nand UO_33 (O_33,N_9445,N_9902);
nor UO_34 (O_34,N_9375,N_9091);
or UO_35 (O_35,N_9303,N_9534);
nor UO_36 (O_36,N_9766,N_9287);
and UO_37 (O_37,N_9250,N_9762);
and UO_38 (O_38,N_9905,N_9097);
nand UO_39 (O_39,N_9741,N_9199);
nand UO_40 (O_40,N_9482,N_9162);
and UO_41 (O_41,N_9043,N_9626);
nor UO_42 (O_42,N_9835,N_9483);
or UO_43 (O_43,N_9578,N_9426);
nand UO_44 (O_44,N_9694,N_9810);
nand UO_45 (O_45,N_9712,N_9551);
and UO_46 (O_46,N_9623,N_9757);
nor UO_47 (O_47,N_9340,N_9848);
nor UO_48 (O_48,N_9703,N_9961);
and UO_49 (O_49,N_9925,N_9887);
nand UO_50 (O_50,N_9153,N_9746);
or UO_51 (O_51,N_9013,N_9115);
or UO_52 (O_52,N_9138,N_9522);
and UO_53 (O_53,N_9935,N_9592);
or UO_54 (O_54,N_9632,N_9075);
nand UO_55 (O_55,N_9275,N_9054);
and UO_56 (O_56,N_9201,N_9214);
and UO_57 (O_57,N_9582,N_9266);
nand UO_58 (O_58,N_9148,N_9099);
nand UO_59 (O_59,N_9548,N_9425);
and UO_60 (O_60,N_9874,N_9755);
nand UO_61 (O_61,N_9293,N_9910);
and UO_62 (O_62,N_9631,N_9279);
or UO_63 (O_63,N_9386,N_9731);
nand UO_64 (O_64,N_9643,N_9413);
nor UO_65 (O_65,N_9559,N_9020);
and UO_66 (O_66,N_9767,N_9845);
or UO_67 (O_67,N_9140,N_9907);
and UO_68 (O_68,N_9360,N_9506);
nand UO_69 (O_69,N_9866,N_9113);
nor UO_70 (O_70,N_9602,N_9418);
nor UO_71 (O_71,N_9489,N_9922);
or UO_72 (O_72,N_9224,N_9371);
nor UO_73 (O_73,N_9430,N_9310);
nor UO_74 (O_74,N_9794,N_9941);
or UO_75 (O_75,N_9180,N_9500);
and UO_76 (O_76,N_9771,N_9979);
and UO_77 (O_77,N_9696,N_9251);
nor UO_78 (O_78,N_9081,N_9352);
nand UO_79 (O_79,N_9010,N_9016);
nor UO_80 (O_80,N_9921,N_9753);
nor UO_81 (O_81,N_9319,N_9624);
nand UO_82 (O_82,N_9241,N_9101);
and UO_83 (O_83,N_9095,N_9187);
nand UO_84 (O_84,N_9955,N_9454);
or UO_85 (O_85,N_9583,N_9282);
or UO_86 (O_86,N_9885,N_9812);
or UO_87 (O_87,N_9052,N_9960);
nand UO_88 (O_88,N_9449,N_9351);
nand UO_89 (O_89,N_9131,N_9704);
nand UO_90 (O_90,N_9744,N_9496);
nor UO_91 (O_91,N_9157,N_9475);
and UO_92 (O_92,N_9620,N_9248);
nor UO_93 (O_93,N_9030,N_9650);
nand UO_94 (O_94,N_9543,N_9367);
nand UO_95 (O_95,N_9897,N_9385);
and UO_96 (O_96,N_9085,N_9209);
nand UO_97 (O_97,N_9665,N_9862);
and UO_98 (O_98,N_9685,N_9533);
nor UO_99 (O_99,N_9892,N_9836);
or UO_100 (O_100,N_9073,N_9383);
nand UO_101 (O_101,N_9673,N_9552);
or UO_102 (O_102,N_9181,N_9082);
nor UO_103 (O_103,N_9337,N_9029);
or UO_104 (O_104,N_9876,N_9005);
nor UO_105 (O_105,N_9575,N_9756);
nand UO_106 (O_106,N_9688,N_9523);
or UO_107 (O_107,N_9787,N_9071);
nor UO_108 (O_108,N_9871,N_9108);
and UO_109 (O_109,N_9038,N_9557);
nor UO_110 (O_110,N_9839,N_9727);
nor UO_111 (O_111,N_9121,N_9151);
nand UO_112 (O_112,N_9312,N_9999);
nor UO_113 (O_113,N_9598,N_9347);
nand UO_114 (O_114,N_9993,N_9384);
xor UO_115 (O_115,N_9570,N_9284);
nor UO_116 (O_116,N_9693,N_9613);
and UO_117 (O_117,N_9527,N_9843);
nand UO_118 (O_118,N_9333,N_9374);
nor UO_119 (O_119,N_9627,N_9675);
and UO_120 (O_120,N_9278,N_9358);
nand UO_121 (O_121,N_9461,N_9743);
nor UO_122 (O_122,N_9311,N_9008);
or UO_123 (O_123,N_9381,N_9429);
nor UO_124 (O_124,N_9652,N_9361);
nand UO_125 (O_125,N_9674,N_9677);
nand UO_126 (O_126,N_9320,N_9451);
nor UO_127 (O_127,N_9804,N_9074);
or UO_128 (O_128,N_9307,N_9612);
or UO_129 (O_129,N_9460,N_9658);
or UO_130 (O_130,N_9210,N_9359);
nor UO_131 (O_131,N_9368,N_9163);
nor UO_132 (O_132,N_9926,N_9574);
and UO_133 (O_133,N_9701,N_9257);
or UO_134 (O_134,N_9263,N_9634);
nand UO_135 (O_135,N_9448,N_9160);
nor UO_136 (O_136,N_9125,N_9591);
nand UO_137 (O_137,N_9988,N_9761);
or UO_138 (O_138,N_9745,N_9657);
or UO_139 (O_139,N_9059,N_9725);
nand UO_140 (O_140,N_9858,N_9962);
nand UO_141 (O_141,N_9034,N_9119);
nand UO_142 (O_142,N_9134,N_9923);
nand UO_143 (O_143,N_9531,N_9107);
nor UO_144 (O_144,N_9009,N_9481);
nor UO_145 (O_145,N_9509,N_9308);
or UO_146 (O_146,N_9102,N_9272);
nand UO_147 (O_147,N_9459,N_9388);
and UO_148 (O_148,N_9328,N_9130);
nand UO_149 (O_149,N_9580,N_9492);
or UO_150 (O_150,N_9649,N_9764);
nor UO_151 (O_151,N_9525,N_9689);
or UO_152 (O_152,N_9778,N_9023);
nor UO_153 (O_153,N_9667,N_9930);
and UO_154 (O_154,N_9900,N_9439);
nand UO_155 (O_155,N_9503,N_9722);
and UO_156 (O_156,N_9289,N_9851);
nor UO_157 (O_157,N_9239,N_9195);
nand UO_158 (O_158,N_9982,N_9560);
nor UO_159 (O_159,N_9989,N_9219);
and UO_160 (O_160,N_9058,N_9398);
or UO_161 (O_161,N_9830,N_9321);
nor UO_162 (O_162,N_9407,N_9774);
nor UO_163 (O_163,N_9477,N_9630);
or UO_164 (O_164,N_9517,N_9409);
nor UO_165 (O_165,N_9220,N_9234);
nand UO_166 (O_166,N_9641,N_9957);
nor UO_167 (O_167,N_9149,N_9264);
nand UO_168 (O_168,N_9716,N_9669);
and UO_169 (O_169,N_9589,N_9640);
nand UO_170 (O_170,N_9387,N_9122);
and UO_171 (O_171,N_9884,N_9141);
or UO_172 (O_172,N_9825,N_9518);
and UO_173 (O_173,N_9648,N_9958);
nand UO_174 (O_174,N_9883,N_9330);
or UO_175 (O_175,N_9490,N_9928);
and UO_176 (O_176,N_9026,N_9572);
nor UO_177 (O_177,N_9948,N_9903);
and UO_178 (O_178,N_9186,N_9408);
and UO_179 (O_179,N_9480,N_9563);
or UO_180 (O_180,N_9050,N_9267);
or UO_181 (O_181,N_9882,N_9080);
or UO_182 (O_182,N_9734,N_9083);
nand UO_183 (O_183,N_9400,N_9909);
or UO_184 (O_184,N_9815,N_9127);
or UO_185 (O_185,N_9348,N_9061);
nor UO_186 (O_186,N_9811,N_9879);
or UO_187 (O_187,N_9854,N_9539);
or UO_188 (O_188,N_9827,N_9818);
nor UO_189 (O_189,N_9856,N_9393);
nand UO_190 (O_190,N_9867,N_9939);
or UO_191 (O_191,N_9645,N_9139);
nor UO_192 (O_192,N_9881,N_9035);
nor UO_193 (O_193,N_9901,N_9644);
nor UO_194 (O_194,N_9914,N_9032);
nor UO_195 (O_195,N_9671,N_9512);
and UO_196 (O_196,N_9309,N_9037);
or UO_197 (O_197,N_9450,N_9159);
or UO_198 (O_198,N_9002,N_9863);
and UO_199 (O_199,N_9795,N_9281);
nand UO_200 (O_200,N_9659,N_9967);
nor UO_201 (O_201,N_9748,N_9007);
nor UO_202 (O_202,N_9126,N_9350);
nor UO_203 (O_203,N_9975,N_9775);
or UO_204 (O_204,N_9864,N_9520);
or UO_205 (O_205,N_9524,N_9555);
nand UO_206 (O_206,N_9614,N_9182);
nor UO_207 (O_207,N_9370,N_9198);
or UO_208 (O_208,N_9912,N_9584);
nand UO_209 (O_209,N_9891,N_9446);
nor UO_210 (O_210,N_9514,N_9440);
nor UO_211 (O_211,N_9633,N_9169);
and UO_212 (O_212,N_9937,N_9576);
nand UO_213 (O_213,N_9110,N_9803);
nand UO_214 (O_214,N_9154,N_9120);
nor UO_215 (O_215,N_9116,N_9323);
or UO_216 (O_216,N_9919,N_9977);
nand UO_217 (O_217,N_9814,N_9114);
and UO_218 (O_218,N_9200,N_9341);
nor UO_219 (O_219,N_9406,N_9676);
and UO_220 (O_220,N_9516,N_9824);
or UO_221 (O_221,N_9754,N_9093);
or UO_222 (O_222,N_9653,N_9604);
nand UO_223 (O_223,N_9012,N_9687);
and UO_224 (O_224,N_9713,N_9342);
or UO_225 (O_225,N_9391,N_9783);
nand UO_226 (O_226,N_9809,N_9699);
nand UO_227 (O_227,N_9390,N_9782);
nand UO_228 (O_228,N_9991,N_9178);
and UO_229 (O_229,N_9164,N_9362);
or UO_230 (O_230,N_9588,N_9684);
nor UO_231 (O_231,N_9338,N_9031);
nand UO_232 (O_232,N_9954,N_9730);
or UO_233 (O_233,N_9956,N_9098);
nor UO_234 (O_234,N_9702,N_9536);
nand UO_235 (O_235,N_9196,N_9111);
nand UO_236 (O_236,N_9807,N_9396);
nor UO_237 (O_237,N_9992,N_9672);
nor UO_238 (O_238,N_9252,N_9270);
nand UO_239 (O_239,N_9066,N_9670);
nand UO_240 (O_240,N_9916,N_9682);
or UO_241 (O_241,N_9192,N_9510);
nand UO_242 (O_242,N_9964,N_9380);
and UO_243 (O_243,N_9695,N_9805);
nand UO_244 (O_244,N_9103,N_9104);
nand UO_245 (O_245,N_9899,N_9339);
nor UO_246 (O_246,N_9711,N_9143);
and UO_247 (O_247,N_9273,N_9661);
and UO_248 (O_248,N_9474,N_9022);
nand UO_249 (O_249,N_9217,N_9049);
nor UO_250 (O_250,N_9647,N_9457);
nor UO_251 (O_251,N_9752,N_9285);
nand UO_252 (O_252,N_9816,N_9505);
or UO_253 (O_253,N_9942,N_9618);
nor UO_254 (O_254,N_9253,N_9732);
nor UO_255 (O_255,N_9412,N_9299);
and UO_256 (O_256,N_9132,N_9924);
or UO_257 (O_257,N_9420,N_9046);
nand UO_258 (O_258,N_9497,N_9959);
or UO_259 (O_259,N_9889,N_9599);
and UO_260 (O_260,N_9541,N_9760);
and UO_261 (O_261,N_9128,N_9222);
and UO_262 (O_262,N_9859,N_9929);
nor UO_263 (O_263,N_9172,N_9467);
nand UO_264 (O_264,N_9297,N_9152);
nor UO_265 (O_265,N_9048,N_9316);
nand UO_266 (O_266,N_9215,N_9232);
or UO_267 (O_267,N_9611,N_9796);
nand UO_268 (O_268,N_9044,N_9053);
nand UO_269 (O_269,N_9519,N_9155);
or UO_270 (O_270,N_9436,N_9822);
and UO_271 (O_271,N_9410,N_9262);
or UO_272 (O_272,N_9369,N_9759);
or UO_273 (O_273,N_9938,N_9972);
nand UO_274 (O_274,N_9343,N_9718);
or UO_275 (O_275,N_9313,N_9268);
or UO_276 (O_276,N_9076,N_9206);
nand UO_277 (O_277,N_9088,N_9158);
and UO_278 (O_278,N_9039,N_9817);
or UO_279 (O_279,N_9094,N_9786);
or UO_280 (O_280,N_9880,N_9985);
and UO_281 (O_281,N_9996,N_9271);
nor UO_282 (O_282,N_9586,N_9092);
and UO_283 (O_283,N_9736,N_9869);
or UO_284 (O_284,N_9984,N_9422);
and UO_285 (O_285,N_9055,N_9417);
nor UO_286 (O_286,N_9717,N_9276);
and UO_287 (O_287,N_9288,N_9784);
or UO_288 (O_288,N_9932,N_9502);
nor UO_289 (O_289,N_9011,N_9737);
or UO_290 (O_290,N_9549,N_9515);
nand UO_291 (O_291,N_9680,N_9465);
nand UO_292 (O_292,N_9968,N_9852);
or UO_293 (O_293,N_9965,N_9109);
nand UO_294 (O_294,N_9493,N_9453);
nor UO_295 (O_295,N_9770,N_9015);
nand UO_296 (O_296,N_9714,N_9184);
and UO_297 (O_297,N_9243,N_9875);
nor UO_298 (O_298,N_9553,N_9573);
nand UO_299 (O_299,N_9473,N_9260);
nand UO_300 (O_300,N_9236,N_9664);
nand UO_301 (O_301,N_9823,N_9364);
nor UO_302 (O_302,N_9742,N_9888);
and UO_303 (O_303,N_9167,N_9806);
or UO_304 (O_304,N_9917,N_9019);
nor UO_305 (O_305,N_9118,N_9980);
nand UO_306 (O_306,N_9399,N_9723);
or UO_307 (O_307,N_9443,N_9820);
nand UO_308 (O_308,N_9000,N_9190);
nand UO_309 (O_309,N_9014,N_9833);
and UO_310 (O_310,N_9908,N_9057);
nand UO_311 (O_311,N_9587,N_9637);
xor UO_312 (O_312,N_9462,N_9018);
and UO_313 (O_313,N_9792,N_9606);
and UO_314 (O_314,N_9763,N_9577);
and UO_315 (O_315,N_9228,N_9793);
and UO_316 (O_316,N_9678,N_9433);
nor UO_317 (O_317,N_9561,N_9245);
and UO_318 (O_318,N_9491,N_9934);
and UO_319 (O_319,N_9062,N_9963);
or UO_320 (O_320,N_9890,N_9305);
nand UO_321 (O_321,N_9683,N_9857);
nand UO_322 (O_322,N_9068,N_9668);
nand UO_323 (O_323,N_9435,N_9006);
nand UO_324 (O_324,N_9596,N_9302);
nor UO_325 (O_325,N_9161,N_9799);
nor UO_326 (O_326,N_9511,N_9679);
nand UO_327 (O_327,N_9933,N_9495);
or UO_328 (O_328,N_9797,N_9565);
nand UO_329 (O_329,N_9028,N_9535);
or UO_330 (O_330,N_9117,N_9137);
and UO_331 (O_331,N_9135,N_9705);
or UO_332 (O_332,N_9404,N_9601);
and UO_333 (O_333,N_9078,N_9376);
nand UO_334 (O_334,N_9204,N_9720);
nand UO_335 (O_335,N_9629,N_9064);
nand UO_336 (O_336,N_9878,N_9735);
and UO_337 (O_337,N_9004,N_9089);
and UO_338 (O_338,N_9545,N_9681);
nand UO_339 (O_339,N_9772,N_9758);
nand UO_340 (O_340,N_9202,N_9697);
nor UO_341 (O_341,N_9168,N_9041);
nor UO_342 (O_342,N_9920,N_9379);
nand UO_343 (O_343,N_9233,N_9306);
nand UO_344 (O_344,N_9998,N_9415);
or UO_345 (O_345,N_9176,N_9100);
nand UO_346 (O_346,N_9504,N_9144);
nand UO_347 (O_347,N_9529,N_9655);
xnor UO_348 (O_348,N_9700,N_9773);
and UO_349 (O_349,N_9240,N_9691);
nor UO_350 (O_350,N_9147,N_9710);
and UO_351 (O_351,N_9444,N_9544);
and UO_352 (O_352,N_9334,N_9619);
and UO_353 (O_353,N_9185,N_9855);
or UO_354 (O_354,N_9256,N_9301);
nor UO_355 (O_355,N_9944,N_9096);
or UO_356 (O_356,N_9471,N_9974);
or UO_357 (O_357,N_9488,N_9296);
nor UO_358 (O_358,N_9269,N_9721);
nor UO_359 (O_359,N_9458,N_9540);
nand UO_360 (O_360,N_9849,N_9090);
and UO_361 (O_361,N_9494,N_9175);
nor UO_362 (O_362,N_9254,N_9651);
and UO_363 (O_363,N_9590,N_9378);
nor UO_364 (O_364,N_9846,N_9150);
nand UO_365 (O_365,N_9171,N_9063);
nor UO_366 (O_366,N_9389,N_9419);
or UO_367 (O_367,N_9365,N_9298);
and UO_368 (O_368,N_9801,N_9616);
and UO_369 (O_369,N_9791,N_9437);
and UO_370 (O_370,N_9853,N_9777);
or UO_371 (O_371,N_9521,N_9327);
nor UO_372 (O_372,N_9749,N_9870);
nor UO_373 (O_373,N_9728,N_9283);
nand UO_374 (O_374,N_9976,N_9781);
or UO_375 (O_375,N_9244,N_9986);
nand UO_376 (O_376,N_9547,N_9397);
nor UO_377 (O_377,N_9079,N_9911);
and UO_378 (O_378,N_9556,N_9569);
or UO_379 (O_379,N_9405,N_9112);
and UO_380 (O_380,N_9751,N_9047);
nor UO_381 (O_381,N_9850,N_9105);
nor UO_382 (O_382,N_9530,N_9382);
nor UO_383 (O_383,N_9841,N_9001);
nor UO_384 (O_384,N_9971,N_9146);
nor UO_385 (O_385,N_9987,N_9086);
and UO_386 (O_386,N_9564,N_9021);
nor UO_387 (O_387,N_9084,N_9646);
or UO_388 (O_388,N_9819,N_9325);
nor UO_389 (O_389,N_9558,N_9318);
nor UO_390 (O_390,N_9625,N_9077);
nand UO_391 (O_391,N_9225,N_9615);
or UO_392 (O_392,N_9466,N_9290);
nand UO_393 (O_393,N_9617,N_9789);
or UO_394 (O_394,N_9872,N_9698);
nand UO_395 (O_395,N_9595,N_9326);
nand UO_396 (O_396,N_9428,N_9441);
nand UO_397 (O_397,N_9173,N_9255);
xor UO_398 (O_398,N_9945,N_9834);
and UO_399 (O_399,N_9597,N_9973);
nand UO_400 (O_400,N_9242,N_9860);
nor UO_401 (O_401,N_9145,N_9357);
and UO_402 (O_402,N_9124,N_9469);
nor UO_403 (O_403,N_9528,N_9508);
and UO_404 (O_404,N_9218,N_9424);
and UO_405 (O_405,N_9315,N_9868);
nand UO_406 (O_406,N_9994,N_9366);
nor UO_407 (O_407,N_9183,N_9070);
xor UO_408 (O_408,N_9970,N_9478);
or UO_409 (O_409,N_9203,N_9274);
nor UO_410 (O_410,N_9230,N_9636);
xor UO_411 (O_411,N_9724,N_9194);
nor UO_412 (O_412,N_9067,N_9893);
or UO_413 (O_413,N_9431,N_9069);
nor UO_414 (O_414,N_9554,N_9769);
and UO_415 (O_415,N_9546,N_9191);
or UO_416 (O_416,N_9780,N_9213);
nand UO_417 (O_417,N_9886,N_9106);
or UO_418 (O_418,N_9821,N_9550);
nor UO_419 (O_419,N_9726,N_9768);
or UO_420 (O_420,N_9345,N_9603);
or UO_421 (O_421,N_9662,N_9377);
and UO_422 (O_422,N_9918,N_9392);
nand UO_423 (O_423,N_9464,N_9142);
or UO_424 (O_424,N_9813,N_9193);
and UO_425 (O_425,N_9779,N_9231);
nor UO_426 (O_426,N_9798,N_9065);
nand UO_427 (O_427,N_9802,N_9566);
nor UO_428 (O_428,N_9719,N_9286);
and UO_429 (O_429,N_9579,N_9567);
or UO_430 (O_430,N_9024,N_9249);
and UO_431 (O_431,N_9188,N_9660);
or UO_432 (O_432,N_9785,N_9808);
and UO_433 (O_433,N_9896,N_9136);
nor UO_434 (O_434,N_9476,N_9776);
or UO_435 (O_435,N_9706,N_9156);
or UO_436 (O_436,N_9983,N_9442);
nor UO_437 (O_437,N_9609,N_9790);
or UO_438 (O_438,N_9501,N_9966);
nand UO_439 (O_439,N_9468,N_9291);
and UO_440 (O_440,N_9344,N_9894);
or UO_441 (O_441,N_9943,N_9947);
nor UO_442 (O_442,N_9170,N_9692);
nor UO_443 (O_443,N_9056,N_9487);
or UO_444 (O_444,N_9940,N_9788);
nor UO_445 (O_445,N_9226,N_9395);
or UO_446 (O_446,N_9363,N_9844);
and UO_447 (O_447,N_9353,N_9740);
or UO_448 (O_448,N_9423,N_9336);
nor UO_449 (O_449,N_9087,N_9133);
nand UO_450 (O_450,N_9455,N_9656);
or UO_451 (O_451,N_9654,N_9532);
or UO_452 (O_452,N_9562,N_9280);
nand UO_453 (O_453,N_9292,N_9593);
nand UO_454 (O_454,N_9258,N_9642);
and UO_455 (O_455,N_9950,N_9621);
or UO_456 (O_456,N_9355,N_9438);
nor UO_457 (O_457,N_9738,N_9739);
nand UO_458 (O_458,N_9040,N_9207);
nand UO_459 (O_459,N_9707,N_9456);
or UO_460 (O_460,N_9499,N_9394);
nor UO_461 (O_461,N_9177,N_9265);
nand UO_462 (O_462,N_9873,N_9294);
nand UO_463 (O_463,N_9237,N_9605);
nor UO_464 (O_464,N_9166,N_9594);
and UO_465 (O_465,N_9427,N_9447);
or UO_466 (O_466,N_9329,N_9229);
xnor UO_467 (O_467,N_9829,N_9877);
or UO_468 (O_468,N_9842,N_9295);
nor UO_469 (O_469,N_9335,N_9838);
or UO_470 (O_470,N_9666,N_9865);
nor UO_471 (O_471,N_9463,N_9638);
nand UO_472 (O_472,N_9610,N_9608);
or UO_473 (O_473,N_9421,N_9033);
or UO_474 (O_474,N_9663,N_9826);
nor UO_475 (O_475,N_9025,N_9542);
nand UO_476 (O_476,N_9733,N_9227);
nand UO_477 (O_477,N_9197,N_9373);
nand UO_478 (O_478,N_9690,N_9952);
nor UO_479 (O_479,N_9212,N_9765);
nand UO_480 (O_480,N_9246,N_9349);
or UO_481 (O_481,N_9913,N_9314);
nor UO_482 (O_482,N_9317,N_9538);
nand UO_483 (O_483,N_9953,N_9060);
and UO_484 (O_484,N_9607,N_9165);
or UO_485 (O_485,N_9709,N_9486);
and UO_486 (O_486,N_9259,N_9990);
or UO_487 (O_487,N_9129,N_9216);
or UO_488 (O_488,N_9221,N_9434);
and UO_489 (O_489,N_9622,N_9927);
nor UO_490 (O_490,N_9832,N_9402);
nand UO_491 (O_491,N_9936,N_9828);
nand UO_492 (O_492,N_9498,N_9411);
nand UO_493 (O_493,N_9847,N_9951);
nor UO_494 (O_494,N_9686,N_9432);
or UO_495 (O_495,N_9635,N_9346);
nor UO_496 (O_496,N_9205,N_9354);
or UO_497 (O_497,N_9800,N_9223);
and UO_498 (O_498,N_9931,N_9997);
nor UO_499 (O_499,N_9042,N_9513);
nand UO_500 (O_500,N_9576,N_9051);
and UO_501 (O_501,N_9287,N_9998);
nand UO_502 (O_502,N_9991,N_9868);
or UO_503 (O_503,N_9494,N_9499);
nand UO_504 (O_504,N_9642,N_9521);
and UO_505 (O_505,N_9860,N_9857);
and UO_506 (O_506,N_9733,N_9275);
nor UO_507 (O_507,N_9890,N_9620);
or UO_508 (O_508,N_9873,N_9115);
or UO_509 (O_509,N_9302,N_9061);
and UO_510 (O_510,N_9437,N_9293);
and UO_511 (O_511,N_9689,N_9931);
and UO_512 (O_512,N_9003,N_9315);
or UO_513 (O_513,N_9973,N_9099);
nor UO_514 (O_514,N_9301,N_9351);
nand UO_515 (O_515,N_9828,N_9278);
nand UO_516 (O_516,N_9894,N_9814);
and UO_517 (O_517,N_9099,N_9733);
nand UO_518 (O_518,N_9204,N_9621);
nor UO_519 (O_519,N_9329,N_9684);
nor UO_520 (O_520,N_9442,N_9985);
nor UO_521 (O_521,N_9941,N_9383);
nand UO_522 (O_522,N_9561,N_9345);
nor UO_523 (O_523,N_9671,N_9007);
nand UO_524 (O_524,N_9020,N_9279);
nor UO_525 (O_525,N_9670,N_9971);
nor UO_526 (O_526,N_9942,N_9902);
xnor UO_527 (O_527,N_9158,N_9146);
nand UO_528 (O_528,N_9819,N_9715);
or UO_529 (O_529,N_9371,N_9078);
nor UO_530 (O_530,N_9757,N_9962);
nand UO_531 (O_531,N_9717,N_9488);
nand UO_532 (O_532,N_9335,N_9649);
and UO_533 (O_533,N_9415,N_9290);
nand UO_534 (O_534,N_9695,N_9627);
or UO_535 (O_535,N_9228,N_9852);
or UO_536 (O_536,N_9349,N_9075);
or UO_537 (O_537,N_9779,N_9369);
nand UO_538 (O_538,N_9357,N_9169);
nand UO_539 (O_539,N_9451,N_9118);
or UO_540 (O_540,N_9038,N_9664);
or UO_541 (O_541,N_9430,N_9947);
nor UO_542 (O_542,N_9870,N_9509);
and UO_543 (O_543,N_9763,N_9843);
nor UO_544 (O_544,N_9229,N_9001);
nand UO_545 (O_545,N_9304,N_9157);
nor UO_546 (O_546,N_9966,N_9839);
or UO_547 (O_547,N_9963,N_9221);
and UO_548 (O_548,N_9338,N_9772);
or UO_549 (O_549,N_9524,N_9337);
nand UO_550 (O_550,N_9470,N_9383);
and UO_551 (O_551,N_9202,N_9394);
nor UO_552 (O_552,N_9464,N_9568);
or UO_553 (O_553,N_9528,N_9953);
or UO_554 (O_554,N_9054,N_9600);
nand UO_555 (O_555,N_9551,N_9292);
and UO_556 (O_556,N_9356,N_9665);
or UO_557 (O_557,N_9825,N_9734);
and UO_558 (O_558,N_9202,N_9907);
nand UO_559 (O_559,N_9094,N_9359);
nor UO_560 (O_560,N_9196,N_9571);
and UO_561 (O_561,N_9957,N_9520);
and UO_562 (O_562,N_9236,N_9442);
or UO_563 (O_563,N_9377,N_9163);
and UO_564 (O_564,N_9875,N_9731);
and UO_565 (O_565,N_9380,N_9257);
or UO_566 (O_566,N_9101,N_9420);
or UO_567 (O_567,N_9636,N_9530);
or UO_568 (O_568,N_9804,N_9315);
nand UO_569 (O_569,N_9441,N_9219);
nand UO_570 (O_570,N_9380,N_9183);
or UO_571 (O_571,N_9657,N_9355);
nand UO_572 (O_572,N_9926,N_9444);
xnor UO_573 (O_573,N_9510,N_9292);
or UO_574 (O_574,N_9733,N_9908);
nand UO_575 (O_575,N_9120,N_9295);
and UO_576 (O_576,N_9473,N_9723);
nor UO_577 (O_577,N_9840,N_9984);
or UO_578 (O_578,N_9653,N_9722);
and UO_579 (O_579,N_9659,N_9835);
nand UO_580 (O_580,N_9881,N_9339);
nor UO_581 (O_581,N_9395,N_9231);
and UO_582 (O_582,N_9727,N_9174);
nand UO_583 (O_583,N_9498,N_9852);
nand UO_584 (O_584,N_9945,N_9987);
nor UO_585 (O_585,N_9132,N_9166);
nand UO_586 (O_586,N_9651,N_9709);
nand UO_587 (O_587,N_9019,N_9838);
nand UO_588 (O_588,N_9907,N_9841);
nor UO_589 (O_589,N_9755,N_9878);
or UO_590 (O_590,N_9514,N_9564);
nand UO_591 (O_591,N_9672,N_9582);
nand UO_592 (O_592,N_9860,N_9865);
nand UO_593 (O_593,N_9903,N_9448);
or UO_594 (O_594,N_9333,N_9156);
or UO_595 (O_595,N_9126,N_9380);
or UO_596 (O_596,N_9997,N_9685);
and UO_597 (O_597,N_9202,N_9313);
or UO_598 (O_598,N_9493,N_9177);
and UO_599 (O_599,N_9961,N_9668);
and UO_600 (O_600,N_9621,N_9904);
nand UO_601 (O_601,N_9918,N_9152);
or UO_602 (O_602,N_9690,N_9029);
or UO_603 (O_603,N_9990,N_9300);
and UO_604 (O_604,N_9793,N_9130);
nand UO_605 (O_605,N_9987,N_9378);
nor UO_606 (O_606,N_9523,N_9552);
or UO_607 (O_607,N_9876,N_9316);
nand UO_608 (O_608,N_9143,N_9684);
nand UO_609 (O_609,N_9392,N_9988);
nor UO_610 (O_610,N_9219,N_9575);
nand UO_611 (O_611,N_9230,N_9956);
and UO_612 (O_612,N_9345,N_9850);
nor UO_613 (O_613,N_9954,N_9440);
nor UO_614 (O_614,N_9943,N_9873);
nand UO_615 (O_615,N_9895,N_9801);
and UO_616 (O_616,N_9516,N_9180);
and UO_617 (O_617,N_9269,N_9021);
nor UO_618 (O_618,N_9242,N_9666);
nor UO_619 (O_619,N_9244,N_9459);
nor UO_620 (O_620,N_9874,N_9016);
or UO_621 (O_621,N_9854,N_9525);
nand UO_622 (O_622,N_9853,N_9140);
nand UO_623 (O_623,N_9300,N_9762);
or UO_624 (O_624,N_9037,N_9748);
xnor UO_625 (O_625,N_9255,N_9126);
nor UO_626 (O_626,N_9368,N_9550);
and UO_627 (O_627,N_9104,N_9707);
and UO_628 (O_628,N_9117,N_9864);
and UO_629 (O_629,N_9579,N_9833);
nor UO_630 (O_630,N_9188,N_9386);
or UO_631 (O_631,N_9147,N_9617);
nand UO_632 (O_632,N_9417,N_9020);
nor UO_633 (O_633,N_9544,N_9098);
nand UO_634 (O_634,N_9154,N_9459);
nor UO_635 (O_635,N_9032,N_9258);
nor UO_636 (O_636,N_9918,N_9224);
nand UO_637 (O_637,N_9773,N_9145);
and UO_638 (O_638,N_9301,N_9142);
nor UO_639 (O_639,N_9941,N_9181);
nor UO_640 (O_640,N_9483,N_9878);
and UO_641 (O_641,N_9039,N_9802);
and UO_642 (O_642,N_9980,N_9432);
and UO_643 (O_643,N_9268,N_9490);
or UO_644 (O_644,N_9003,N_9433);
xor UO_645 (O_645,N_9577,N_9635);
and UO_646 (O_646,N_9999,N_9471);
or UO_647 (O_647,N_9775,N_9147);
and UO_648 (O_648,N_9536,N_9047);
and UO_649 (O_649,N_9657,N_9958);
nor UO_650 (O_650,N_9882,N_9756);
and UO_651 (O_651,N_9872,N_9188);
nand UO_652 (O_652,N_9861,N_9944);
and UO_653 (O_653,N_9967,N_9495);
and UO_654 (O_654,N_9046,N_9494);
nor UO_655 (O_655,N_9227,N_9071);
or UO_656 (O_656,N_9344,N_9297);
nand UO_657 (O_657,N_9990,N_9273);
or UO_658 (O_658,N_9475,N_9976);
and UO_659 (O_659,N_9974,N_9488);
nand UO_660 (O_660,N_9096,N_9544);
nor UO_661 (O_661,N_9285,N_9282);
nor UO_662 (O_662,N_9259,N_9223);
nand UO_663 (O_663,N_9903,N_9073);
or UO_664 (O_664,N_9526,N_9547);
or UO_665 (O_665,N_9314,N_9654);
or UO_666 (O_666,N_9584,N_9017);
nand UO_667 (O_667,N_9675,N_9014);
or UO_668 (O_668,N_9570,N_9219);
nand UO_669 (O_669,N_9986,N_9163);
nor UO_670 (O_670,N_9465,N_9988);
nand UO_671 (O_671,N_9847,N_9261);
and UO_672 (O_672,N_9691,N_9849);
nor UO_673 (O_673,N_9523,N_9499);
nand UO_674 (O_674,N_9398,N_9262);
or UO_675 (O_675,N_9101,N_9511);
nand UO_676 (O_676,N_9481,N_9497);
or UO_677 (O_677,N_9439,N_9116);
or UO_678 (O_678,N_9011,N_9527);
nand UO_679 (O_679,N_9916,N_9713);
nor UO_680 (O_680,N_9504,N_9084);
nor UO_681 (O_681,N_9441,N_9937);
nand UO_682 (O_682,N_9174,N_9186);
and UO_683 (O_683,N_9912,N_9718);
and UO_684 (O_684,N_9373,N_9328);
or UO_685 (O_685,N_9413,N_9261);
nand UO_686 (O_686,N_9042,N_9812);
nand UO_687 (O_687,N_9596,N_9546);
and UO_688 (O_688,N_9828,N_9668);
nand UO_689 (O_689,N_9429,N_9491);
nor UO_690 (O_690,N_9972,N_9245);
nor UO_691 (O_691,N_9501,N_9681);
and UO_692 (O_692,N_9587,N_9356);
nand UO_693 (O_693,N_9486,N_9312);
or UO_694 (O_694,N_9443,N_9306);
nor UO_695 (O_695,N_9859,N_9712);
or UO_696 (O_696,N_9290,N_9891);
and UO_697 (O_697,N_9965,N_9140);
and UO_698 (O_698,N_9722,N_9795);
nor UO_699 (O_699,N_9374,N_9074);
and UO_700 (O_700,N_9026,N_9333);
and UO_701 (O_701,N_9841,N_9560);
and UO_702 (O_702,N_9559,N_9619);
and UO_703 (O_703,N_9000,N_9843);
or UO_704 (O_704,N_9468,N_9300);
nor UO_705 (O_705,N_9225,N_9662);
and UO_706 (O_706,N_9095,N_9338);
xor UO_707 (O_707,N_9789,N_9501);
nor UO_708 (O_708,N_9693,N_9653);
nand UO_709 (O_709,N_9605,N_9511);
and UO_710 (O_710,N_9878,N_9300);
nand UO_711 (O_711,N_9025,N_9615);
xnor UO_712 (O_712,N_9189,N_9456);
nand UO_713 (O_713,N_9059,N_9302);
nand UO_714 (O_714,N_9478,N_9490);
or UO_715 (O_715,N_9765,N_9071);
nor UO_716 (O_716,N_9590,N_9449);
nor UO_717 (O_717,N_9442,N_9479);
and UO_718 (O_718,N_9914,N_9718);
and UO_719 (O_719,N_9706,N_9302);
nand UO_720 (O_720,N_9342,N_9772);
or UO_721 (O_721,N_9388,N_9307);
nor UO_722 (O_722,N_9982,N_9129);
or UO_723 (O_723,N_9800,N_9817);
nand UO_724 (O_724,N_9536,N_9833);
or UO_725 (O_725,N_9837,N_9277);
nand UO_726 (O_726,N_9534,N_9089);
and UO_727 (O_727,N_9623,N_9404);
or UO_728 (O_728,N_9020,N_9927);
nor UO_729 (O_729,N_9283,N_9226);
and UO_730 (O_730,N_9226,N_9641);
or UO_731 (O_731,N_9276,N_9914);
nand UO_732 (O_732,N_9849,N_9879);
nor UO_733 (O_733,N_9029,N_9886);
and UO_734 (O_734,N_9936,N_9124);
and UO_735 (O_735,N_9736,N_9616);
nand UO_736 (O_736,N_9252,N_9599);
xnor UO_737 (O_737,N_9591,N_9518);
nor UO_738 (O_738,N_9301,N_9618);
nand UO_739 (O_739,N_9406,N_9570);
nand UO_740 (O_740,N_9008,N_9408);
nor UO_741 (O_741,N_9404,N_9196);
or UO_742 (O_742,N_9017,N_9342);
or UO_743 (O_743,N_9092,N_9501);
nand UO_744 (O_744,N_9074,N_9357);
or UO_745 (O_745,N_9900,N_9501);
nand UO_746 (O_746,N_9820,N_9781);
xor UO_747 (O_747,N_9073,N_9774);
nor UO_748 (O_748,N_9846,N_9694);
or UO_749 (O_749,N_9627,N_9895);
and UO_750 (O_750,N_9093,N_9811);
or UO_751 (O_751,N_9391,N_9380);
or UO_752 (O_752,N_9157,N_9263);
nor UO_753 (O_753,N_9783,N_9436);
nand UO_754 (O_754,N_9032,N_9038);
or UO_755 (O_755,N_9399,N_9721);
nor UO_756 (O_756,N_9944,N_9802);
nand UO_757 (O_757,N_9741,N_9238);
and UO_758 (O_758,N_9926,N_9856);
nor UO_759 (O_759,N_9514,N_9689);
nand UO_760 (O_760,N_9831,N_9311);
or UO_761 (O_761,N_9871,N_9581);
nand UO_762 (O_762,N_9907,N_9388);
or UO_763 (O_763,N_9623,N_9290);
nand UO_764 (O_764,N_9350,N_9987);
nor UO_765 (O_765,N_9284,N_9561);
or UO_766 (O_766,N_9127,N_9716);
nand UO_767 (O_767,N_9961,N_9919);
or UO_768 (O_768,N_9681,N_9273);
and UO_769 (O_769,N_9905,N_9972);
nand UO_770 (O_770,N_9750,N_9809);
or UO_771 (O_771,N_9053,N_9332);
nor UO_772 (O_772,N_9622,N_9975);
or UO_773 (O_773,N_9442,N_9730);
nand UO_774 (O_774,N_9018,N_9938);
or UO_775 (O_775,N_9849,N_9274);
xor UO_776 (O_776,N_9359,N_9616);
nor UO_777 (O_777,N_9333,N_9817);
or UO_778 (O_778,N_9367,N_9997);
and UO_779 (O_779,N_9231,N_9666);
and UO_780 (O_780,N_9141,N_9679);
nand UO_781 (O_781,N_9584,N_9824);
nor UO_782 (O_782,N_9906,N_9971);
or UO_783 (O_783,N_9954,N_9790);
nand UO_784 (O_784,N_9646,N_9187);
xor UO_785 (O_785,N_9363,N_9953);
and UO_786 (O_786,N_9834,N_9391);
nor UO_787 (O_787,N_9411,N_9945);
nand UO_788 (O_788,N_9271,N_9965);
nor UO_789 (O_789,N_9358,N_9571);
or UO_790 (O_790,N_9556,N_9861);
nand UO_791 (O_791,N_9500,N_9521);
and UO_792 (O_792,N_9219,N_9207);
and UO_793 (O_793,N_9239,N_9809);
nand UO_794 (O_794,N_9000,N_9737);
nand UO_795 (O_795,N_9022,N_9613);
and UO_796 (O_796,N_9058,N_9919);
or UO_797 (O_797,N_9290,N_9301);
or UO_798 (O_798,N_9577,N_9525);
and UO_799 (O_799,N_9354,N_9560);
or UO_800 (O_800,N_9239,N_9027);
nor UO_801 (O_801,N_9668,N_9101);
nor UO_802 (O_802,N_9869,N_9126);
and UO_803 (O_803,N_9546,N_9490);
and UO_804 (O_804,N_9957,N_9708);
nor UO_805 (O_805,N_9516,N_9644);
xnor UO_806 (O_806,N_9047,N_9197);
nor UO_807 (O_807,N_9747,N_9129);
and UO_808 (O_808,N_9280,N_9140);
nor UO_809 (O_809,N_9831,N_9674);
or UO_810 (O_810,N_9839,N_9190);
nand UO_811 (O_811,N_9587,N_9483);
nand UO_812 (O_812,N_9670,N_9922);
or UO_813 (O_813,N_9415,N_9436);
and UO_814 (O_814,N_9719,N_9157);
nand UO_815 (O_815,N_9437,N_9366);
nor UO_816 (O_816,N_9754,N_9284);
or UO_817 (O_817,N_9128,N_9929);
or UO_818 (O_818,N_9894,N_9505);
nand UO_819 (O_819,N_9285,N_9519);
nor UO_820 (O_820,N_9306,N_9974);
nor UO_821 (O_821,N_9022,N_9759);
xnor UO_822 (O_822,N_9347,N_9880);
nor UO_823 (O_823,N_9168,N_9098);
nand UO_824 (O_824,N_9361,N_9431);
and UO_825 (O_825,N_9834,N_9752);
and UO_826 (O_826,N_9102,N_9439);
and UO_827 (O_827,N_9254,N_9846);
nand UO_828 (O_828,N_9443,N_9262);
and UO_829 (O_829,N_9470,N_9427);
or UO_830 (O_830,N_9380,N_9430);
nand UO_831 (O_831,N_9928,N_9574);
or UO_832 (O_832,N_9534,N_9997);
or UO_833 (O_833,N_9293,N_9816);
or UO_834 (O_834,N_9445,N_9478);
and UO_835 (O_835,N_9743,N_9829);
or UO_836 (O_836,N_9463,N_9320);
or UO_837 (O_837,N_9050,N_9250);
and UO_838 (O_838,N_9058,N_9576);
xor UO_839 (O_839,N_9526,N_9340);
nand UO_840 (O_840,N_9649,N_9060);
and UO_841 (O_841,N_9841,N_9116);
or UO_842 (O_842,N_9464,N_9279);
nand UO_843 (O_843,N_9053,N_9109);
or UO_844 (O_844,N_9779,N_9953);
or UO_845 (O_845,N_9923,N_9257);
and UO_846 (O_846,N_9577,N_9594);
or UO_847 (O_847,N_9278,N_9436);
nand UO_848 (O_848,N_9997,N_9631);
and UO_849 (O_849,N_9065,N_9986);
nor UO_850 (O_850,N_9040,N_9582);
or UO_851 (O_851,N_9901,N_9643);
and UO_852 (O_852,N_9632,N_9680);
nand UO_853 (O_853,N_9685,N_9104);
and UO_854 (O_854,N_9991,N_9832);
or UO_855 (O_855,N_9425,N_9779);
or UO_856 (O_856,N_9375,N_9271);
or UO_857 (O_857,N_9535,N_9439);
nor UO_858 (O_858,N_9969,N_9437);
nor UO_859 (O_859,N_9553,N_9714);
and UO_860 (O_860,N_9660,N_9533);
and UO_861 (O_861,N_9600,N_9011);
and UO_862 (O_862,N_9123,N_9555);
and UO_863 (O_863,N_9326,N_9083);
nor UO_864 (O_864,N_9192,N_9662);
or UO_865 (O_865,N_9298,N_9867);
nor UO_866 (O_866,N_9878,N_9463);
and UO_867 (O_867,N_9334,N_9174);
and UO_868 (O_868,N_9831,N_9881);
and UO_869 (O_869,N_9837,N_9707);
or UO_870 (O_870,N_9685,N_9031);
nand UO_871 (O_871,N_9593,N_9740);
nand UO_872 (O_872,N_9984,N_9232);
nor UO_873 (O_873,N_9048,N_9711);
or UO_874 (O_874,N_9360,N_9848);
nand UO_875 (O_875,N_9278,N_9681);
nand UO_876 (O_876,N_9506,N_9179);
and UO_877 (O_877,N_9868,N_9544);
nor UO_878 (O_878,N_9992,N_9991);
nor UO_879 (O_879,N_9434,N_9906);
nor UO_880 (O_880,N_9284,N_9052);
or UO_881 (O_881,N_9815,N_9644);
nand UO_882 (O_882,N_9171,N_9101);
nand UO_883 (O_883,N_9524,N_9017);
or UO_884 (O_884,N_9781,N_9435);
nand UO_885 (O_885,N_9137,N_9939);
or UO_886 (O_886,N_9749,N_9707);
nand UO_887 (O_887,N_9239,N_9660);
and UO_888 (O_888,N_9815,N_9831);
nor UO_889 (O_889,N_9920,N_9068);
nand UO_890 (O_890,N_9013,N_9435);
or UO_891 (O_891,N_9955,N_9054);
nand UO_892 (O_892,N_9629,N_9502);
nand UO_893 (O_893,N_9288,N_9939);
nand UO_894 (O_894,N_9179,N_9001);
nand UO_895 (O_895,N_9551,N_9776);
nor UO_896 (O_896,N_9763,N_9124);
nand UO_897 (O_897,N_9740,N_9451);
and UO_898 (O_898,N_9905,N_9729);
nor UO_899 (O_899,N_9419,N_9903);
nand UO_900 (O_900,N_9340,N_9566);
nor UO_901 (O_901,N_9487,N_9375);
nor UO_902 (O_902,N_9719,N_9177);
nor UO_903 (O_903,N_9289,N_9911);
or UO_904 (O_904,N_9618,N_9048);
nor UO_905 (O_905,N_9639,N_9778);
nand UO_906 (O_906,N_9111,N_9433);
or UO_907 (O_907,N_9274,N_9563);
nand UO_908 (O_908,N_9071,N_9499);
or UO_909 (O_909,N_9698,N_9741);
and UO_910 (O_910,N_9064,N_9363);
and UO_911 (O_911,N_9900,N_9949);
nor UO_912 (O_912,N_9159,N_9215);
nor UO_913 (O_913,N_9693,N_9232);
and UO_914 (O_914,N_9531,N_9817);
or UO_915 (O_915,N_9597,N_9659);
and UO_916 (O_916,N_9532,N_9839);
and UO_917 (O_917,N_9652,N_9806);
or UO_918 (O_918,N_9867,N_9403);
or UO_919 (O_919,N_9625,N_9558);
and UO_920 (O_920,N_9651,N_9444);
and UO_921 (O_921,N_9219,N_9749);
and UO_922 (O_922,N_9177,N_9240);
or UO_923 (O_923,N_9791,N_9370);
and UO_924 (O_924,N_9231,N_9244);
nand UO_925 (O_925,N_9235,N_9435);
nand UO_926 (O_926,N_9250,N_9658);
nand UO_927 (O_927,N_9368,N_9631);
xnor UO_928 (O_928,N_9952,N_9870);
nand UO_929 (O_929,N_9436,N_9940);
or UO_930 (O_930,N_9793,N_9646);
nand UO_931 (O_931,N_9650,N_9232);
or UO_932 (O_932,N_9133,N_9254);
or UO_933 (O_933,N_9554,N_9213);
nand UO_934 (O_934,N_9300,N_9490);
nand UO_935 (O_935,N_9664,N_9353);
or UO_936 (O_936,N_9299,N_9915);
and UO_937 (O_937,N_9920,N_9745);
and UO_938 (O_938,N_9234,N_9653);
nand UO_939 (O_939,N_9346,N_9059);
and UO_940 (O_940,N_9391,N_9428);
nand UO_941 (O_941,N_9224,N_9447);
and UO_942 (O_942,N_9859,N_9954);
or UO_943 (O_943,N_9197,N_9272);
nand UO_944 (O_944,N_9569,N_9577);
and UO_945 (O_945,N_9762,N_9916);
and UO_946 (O_946,N_9662,N_9983);
nor UO_947 (O_947,N_9397,N_9333);
nand UO_948 (O_948,N_9675,N_9895);
and UO_949 (O_949,N_9849,N_9461);
or UO_950 (O_950,N_9862,N_9537);
or UO_951 (O_951,N_9754,N_9321);
nor UO_952 (O_952,N_9910,N_9360);
and UO_953 (O_953,N_9698,N_9571);
nand UO_954 (O_954,N_9630,N_9940);
or UO_955 (O_955,N_9157,N_9905);
nand UO_956 (O_956,N_9413,N_9585);
or UO_957 (O_957,N_9343,N_9459);
nand UO_958 (O_958,N_9009,N_9791);
nor UO_959 (O_959,N_9669,N_9186);
xnor UO_960 (O_960,N_9685,N_9398);
and UO_961 (O_961,N_9517,N_9235);
nand UO_962 (O_962,N_9503,N_9717);
nor UO_963 (O_963,N_9460,N_9723);
nor UO_964 (O_964,N_9455,N_9138);
and UO_965 (O_965,N_9173,N_9363);
nand UO_966 (O_966,N_9661,N_9684);
and UO_967 (O_967,N_9912,N_9306);
and UO_968 (O_968,N_9895,N_9018);
nor UO_969 (O_969,N_9695,N_9661);
nand UO_970 (O_970,N_9213,N_9023);
nand UO_971 (O_971,N_9756,N_9897);
or UO_972 (O_972,N_9930,N_9564);
nor UO_973 (O_973,N_9711,N_9997);
and UO_974 (O_974,N_9472,N_9831);
nand UO_975 (O_975,N_9623,N_9765);
or UO_976 (O_976,N_9149,N_9443);
and UO_977 (O_977,N_9435,N_9487);
nand UO_978 (O_978,N_9427,N_9953);
nand UO_979 (O_979,N_9401,N_9612);
or UO_980 (O_980,N_9390,N_9714);
nand UO_981 (O_981,N_9014,N_9275);
and UO_982 (O_982,N_9186,N_9244);
nor UO_983 (O_983,N_9912,N_9374);
nand UO_984 (O_984,N_9006,N_9215);
and UO_985 (O_985,N_9745,N_9604);
nor UO_986 (O_986,N_9762,N_9494);
or UO_987 (O_987,N_9064,N_9038);
and UO_988 (O_988,N_9323,N_9767);
nand UO_989 (O_989,N_9591,N_9653);
or UO_990 (O_990,N_9447,N_9099);
nor UO_991 (O_991,N_9175,N_9272);
or UO_992 (O_992,N_9098,N_9494);
nand UO_993 (O_993,N_9531,N_9053);
and UO_994 (O_994,N_9357,N_9867);
nand UO_995 (O_995,N_9197,N_9901);
nor UO_996 (O_996,N_9537,N_9394);
nand UO_997 (O_997,N_9743,N_9846);
nand UO_998 (O_998,N_9053,N_9032);
nand UO_999 (O_999,N_9137,N_9562);
or UO_1000 (O_1000,N_9294,N_9085);
nand UO_1001 (O_1001,N_9291,N_9663);
or UO_1002 (O_1002,N_9456,N_9275);
nor UO_1003 (O_1003,N_9422,N_9627);
or UO_1004 (O_1004,N_9697,N_9240);
and UO_1005 (O_1005,N_9982,N_9262);
nor UO_1006 (O_1006,N_9344,N_9982);
and UO_1007 (O_1007,N_9747,N_9268);
and UO_1008 (O_1008,N_9986,N_9286);
or UO_1009 (O_1009,N_9439,N_9134);
nand UO_1010 (O_1010,N_9181,N_9763);
and UO_1011 (O_1011,N_9060,N_9143);
or UO_1012 (O_1012,N_9490,N_9663);
and UO_1013 (O_1013,N_9294,N_9541);
nand UO_1014 (O_1014,N_9989,N_9418);
nor UO_1015 (O_1015,N_9594,N_9831);
or UO_1016 (O_1016,N_9608,N_9821);
nand UO_1017 (O_1017,N_9591,N_9108);
nand UO_1018 (O_1018,N_9252,N_9107);
or UO_1019 (O_1019,N_9069,N_9353);
nor UO_1020 (O_1020,N_9451,N_9028);
and UO_1021 (O_1021,N_9274,N_9881);
nor UO_1022 (O_1022,N_9031,N_9067);
or UO_1023 (O_1023,N_9505,N_9165);
nand UO_1024 (O_1024,N_9107,N_9951);
nand UO_1025 (O_1025,N_9131,N_9228);
and UO_1026 (O_1026,N_9870,N_9488);
nand UO_1027 (O_1027,N_9747,N_9125);
or UO_1028 (O_1028,N_9157,N_9755);
nand UO_1029 (O_1029,N_9370,N_9092);
nand UO_1030 (O_1030,N_9549,N_9958);
nor UO_1031 (O_1031,N_9203,N_9703);
nor UO_1032 (O_1032,N_9283,N_9561);
or UO_1033 (O_1033,N_9888,N_9224);
xnor UO_1034 (O_1034,N_9132,N_9351);
nor UO_1035 (O_1035,N_9041,N_9485);
nand UO_1036 (O_1036,N_9740,N_9123);
nand UO_1037 (O_1037,N_9887,N_9084);
xnor UO_1038 (O_1038,N_9064,N_9927);
nand UO_1039 (O_1039,N_9848,N_9226);
nor UO_1040 (O_1040,N_9658,N_9837);
or UO_1041 (O_1041,N_9790,N_9966);
nor UO_1042 (O_1042,N_9919,N_9480);
and UO_1043 (O_1043,N_9621,N_9195);
nand UO_1044 (O_1044,N_9975,N_9475);
nand UO_1045 (O_1045,N_9448,N_9073);
and UO_1046 (O_1046,N_9335,N_9465);
nand UO_1047 (O_1047,N_9391,N_9305);
nor UO_1048 (O_1048,N_9650,N_9356);
or UO_1049 (O_1049,N_9733,N_9377);
nand UO_1050 (O_1050,N_9077,N_9659);
or UO_1051 (O_1051,N_9004,N_9156);
and UO_1052 (O_1052,N_9049,N_9897);
nor UO_1053 (O_1053,N_9223,N_9198);
xnor UO_1054 (O_1054,N_9836,N_9767);
and UO_1055 (O_1055,N_9157,N_9012);
nor UO_1056 (O_1056,N_9909,N_9032);
nand UO_1057 (O_1057,N_9727,N_9764);
or UO_1058 (O_1058,N_9062,N_9506);
nor UO_1059 (O_1059,N_9108,N_9808);
nor UO_1060 (O_1060,N_9721,N_9022);
nand UO_1061 (O_1061,N_9463,N_9438);
nand UO_1062 (O_1062,N_9703,N_9494);
nand UO_1063 (O_1063,N_9233,N_9414);
or UO_1064 (O_1064,N_9807,N_9256);
nor UO_1065 (O_1065,N_9218,N_9687);
nor UO_1066 (O_1066,N_9514,N_9814);
or UO_1067 (O_1067,N_9005,N_9291);
nor UO_1068 (O_1068,N_9550,N_9187);
nor UO_1069 (O_1069,N_9764,N_9993);
nand UO_1070 (O_1070,N_9107,N_9288);
nand UO_1071 (O_1071,N_9143,N_9678);
nor UO_1072 (O_1072,N_9572,N_9865);
nand UO_1073 (O_1073,N_9448,N_9503);
or UO_1074 (O_1074,N_9996,N_9380);
or UO_1075 (O_1075,N_9036,N_9562);
or UO_1076 (O_1076,N_9507,N_9490);
or UO_1077 (O_1077,N_9852,N_9071);
and UO_1078 (O_1078,N_9729,N_9877);
nand UO_1079 (O_1079,N_9707,N_9954);
or UO_1080 (O_1080,N_9782,N_9451);
and UO_1081 (O_1081,N_9941,N_9608);
nand UO_1082 (O_1082,N_9718,N_9198);
and UO_1083 (O_1083,N_9922,N_9014);
nor UO_1084 (O_1084,N_9569,N_9504);
nand UO_1085 (O_1085,N_9135,N_9992);
and UO_1086 (O_1086,N_9048,N_9041);
nand UO_1087 (O_1087,N_9161,N_9699);
or UO_1088 (O_1088,N_9489,N_9459);
or UO_1089 (O_1089,N_9692,N_9766);
nor UO_1090 (O_1090,N_9297,N_9267);
nand UO_1091 (O_1091,N_9782,N_9431);
and UO_1092 (O_1092,N_9573,N_9075);
nand UO_1093 (O_1093,N_9323,N_9454);
nor UO_1094 (O_1094,N_9252,N_9448);
nor UO_1095 (O_1095,N_9192,N_9813);
nand UO_1096 (O_1096,N_9543,N_9065);
and UO_1097 (O_1097,N_9629,N_9842);
nand UO_1098 (O_1098,N_9063,N_9585);
or UO_1099 (O_1099,N_9274,N_9380);
nor UO_1100 (O_1100,N_9792,N_9680);
and UO_1101 (O_1101,N_9525,N_9210);
and UO_1102 (O_1102,N_9320,N_9309);
and UO_1103 (O_1103,N_9946,N_9821);
or UO_1104 (O_1104,N_9115,N_9314);
or UO_1105 (O_1105,N_9859,N_9345);
and UO_1106 (O_1106,N_9803,N_9964);
nor UO_1107 (O_1107,N_9862,N_9209);
and UO_1108 (O_1108,N_9822,N_9549);
nand UO_1109 (O_1109,N_9595,N_9954);
or UO_1110 (O_1110,N_9921,N_9728);
nand UO_1111 (O_1111,N_9617,N_9206);
nor UO_1112 (O_1112,N_9333,N_9040);
nand UO_1113 (O_1113,N_9373,N_9504);
and UO_1114 (O_1114,N_9050,N_9158);
and UO_1115 (O_1115,N_9000,N_9630);
nor UO_1116 (O_1116,N_9022,N_9789);
nor UO_1117 (O_1117,N_9928,N_9337);
nand UO_1118 (O_1118,N_9717,N_9672);
and UO_1119 (O_1119,N_9100,N_9132);
and UO_1120 (O_1120,N_9860,N_9504);
and UO_1121 (O_1121,N_9823,N_9250);
nand UO_1122 (O_1122,N_9572,N_9674);
nand UO_1123 (O_1123,N_9213,N_9106);
and UO_1124 (O_1124,N_9131,N_9192);
nor UO_1125 (O_1125,N_9321,N_9636);
or UO_1126 (O_1126,N_9295,N_9533);
or UO_1127 (O_1127,N_9639,N_9223);
and UO_1128 (O_1128,N_9858,N_9879);
nor UO_1129 (O_1129,N_9694,N_9593);
nor UO_1130 (O_1130,N_9917,N_9381);
nor UO_1131 (O_1131,N_9617,N_9937);
nor UO_1132 (O_1132,N_9996,N_9676);
nor UO_1133 (O_1133,N_9784,N_9372);
nor UO_1134 (O_1134,N_9690,N_9325);
or UO_1135 (O_1135,N_9627,N_9763);
and UO_1136 (O_1136,N_9303,N_9602);
nand UO_1137 (O_1137,N_9671,N_9604);
nor UO_1138 (O_1138,N_9105,N_9531);
nand UO_1139 (O_1139,N_9468,N_9658);
or UO_1140 (O_1140,N_9303,N_9008);
or UO_1141 (O_1141,N_9301,N_9644);
nand UO_1142 (O_1142,N_9105,N_9346);
and UO_1143 (O_1143,N_9914,N_9692);
nand UO_1144 (O_1144,N_9210,N_9743);
or UO_1145 (O_1145,N_9479,N_9550);
and UO_1146 (O_1146,N_9537,N_9713);
nor UO_1147 (O_1147,N_9363,N_9401);
nor UO_1148 (O_1148,N_9938,N_9444);
nor UO_1149 (O_1149,N_9554,N_9124);
or UO_1150 (O_1150,N_9088,N_9978);
and UO_1151 (O_1151,N_9784,N_9543);
nand UO_1152 (O_1152,N_9223,N_9289);
and UO_1153 (O_1153,N_9051,N_9342);
and UO_1154 (O_1154,N_9178,N_9927);
or UO_1155 (O_1155,N_9103,N_9131);
or UO_1156 (O_1156,N_9521,N_9826);
or UO_1157 (O_1157,N_9104,N_9326);
nor UO_1158 (O_1158,N_9333,N_9412);
and UO_1159 (O_1159,N_9280,N_9955);
nand UO_1160 (O_1160,N_9675,N_9428);
nor UO_1161 (O_1161,N_9329,N_9666);
nor UO_1162 (O_1162,N_9670,N_9490);
or UO_1163 (O_1163,N_9208,N_9151);
nor UO_1164 (O_1164,N_9119,N_9608);
or UO_1165 (O_1165,N_9944,N_9515);
nor UO_1166 (O_1166,N_9462,N_9794);
or UO_1167 (O_1167,N_9608,N_9076);
and UO_1168 (O_1168,N_9273,N_9060);
or UO_1169 (O_1169,N_9842,N_9103);
or UO_1170 (O_1170,N_9756,N_9840);
nand UO_1171 (O_1171,N_9394,N_9651);
or UO_1172 (O_1172,N_9114,N_9428);
and UO_1173 (O_1173,N_9067,N_9058);
and UO_1174 (O_1174,N_9535,N_9928);
nor UO_1175 (O_1175,N_9264,N_9286);
or UO_1176 (O_1176,N_9968,N_9396);
and UO_1177 (O_1177,N_9767,N_9066);
nor UO_1178 (O_1178,N_9188,N_9168);
and UO_1179 (O_1179,N_9583,N_9283);
and UO_1180 (O_1180,N_9235,N_9066);
and UO_1181 (O_1181,N_9816,N_9450);
nand UO_1182 (O_1182,N_9019,N_9172);
and UO_1183 (O_1183,N_9552,N_9159);
nand UO_1184 (O_1184,N_9128,N_9541);
nand UO_1185 (O_1185,N_9729,N_9163);
nand UO_1186 (O_1186,N_9888,N_9030);
and UO_1187 (O_1187,N_9074,N_9413);
nor UO_1188 (O_1188,N_9956,N_9456);
nand UO_1189 (O_1189,N_9379,N_9882);
nor UO_1190 (O_1190,N_9609,N_9631);
nor UO_1191 (O_1191,N_9160,N_9699);
or UO_1192 (O_1192,N_9120,N_9340);
nand UO_1193 (O_1193,N_9972,N_9772);
or UO_1194 (O_1194,N_9586,N_9469);
nor UO_1195 (O_1195,N_9659,N_9656);
or UO_1196 (O_1196,N_9167,N_9375);
and UO_1197 (O_1197,N_9860,N_9636);
nand UO_1198 (O_1198,N_9878,N_9214);
or UO_1199 (O_1199,N_9340,N_9430);
nor UO_1200 (O_1200,N_9086,N_9757);
or UO_1201 (O_1201,N_9138,N_9015);
or UO_1202 (O_1202,N_9181,N_9732);
nand UO_1203 (O_1203,N_9000,N_9824);
or UO_1204 (O_1204,N_9622,N_9477);
nor UO_1205 (O_1205,N_9854,N_9808);
nor UO_1206 (O_1206,N_9437,N_9884);
and UO_1207 (O_1207,N_9056,N_9216);
or UO_1208 (O_1208,N_9857,N_9188);
nor UO_1209 (O_1209,N_9653,N_9314);
nand UO_1210 (O_1210,N_9455,N_9383);
nor UO_1211 (O_1211,N_9931,N_9051);
and UO_1212 (O_1212,N_9794,N_9556);
and UO_1213 (O_1213,N_9765,N_9960);
or UO_1214 (O_1214,N_9911,N_9585);
and UO_1215 (O_1215,N_9017,N_9528);
and UO_1216 (O_1216,N_9851,N_9803);
nor UO_1217 (O_1217,N_9458,N_9838);
nand UO_1218 (O_1218,N_9870,N_9500);
nor UO_1219 (O_1219,N_9419,N_9091);
nor UO_1220 (O_1220,N_9283,N_9881);
nor UO_1221 (O_1221,N_9310,N_9040);
nor UO_1222 (O_1222,N_9905,N_9018);
nand UO_1223 (O_1223,N_9235,N_9117);
or UO_1224 (O_1224,N_9503,N_9355);
and UO_1225 (O_1225,N_9153,N_9097);
and UO_1226 (O_1226,N_9718,N_9337);
or UO_1227 (O_1227,N_9864,N_9914);
and UO_1228 (O_1228,N_9279,N_9979);
nand UO_1229 (O_1229,N_9858,N_9235);
nor UO_1230 (O_1230,N_9276,N_9520);
and UO_1231 (O_1231,N_9883,N_9062);
and UO_1232 (O_1232,N_9487,N_9186);
or UO_1233 (O_1233,N_9057,N_9568);
nor UO_1234 (O_1234,N_9591,N_9577);
and UO_1235 (O_1235,N_9886,N_9221);
nand UO_1236 (O_1236,N_9630,N_9255);
or UO_1237 (O_1237,N_9872,N_9614);
nor UO_1238 (O_1238,N_9858,N_9318);
nand UO_1239 (O_1239,N_9867,N_9599);
or UO_1240 (O_1240,N_9938,N_9319);
and UO_1241 (O_1241,N_9730,N_9667);
or UO_1242 (O_1242,N_9779,N_9846);
or UO_1243 (O_1243,N_9128,N_9647);
nor UO_1244 (O_1244,N_9937,N_9099);
nand UO_1245 (O_1245,N_9808,N_9048);
nor UO_1246 (O_1246,N_9499,N_9261);
nand UO_1247 (O_1247,N_9605,N_9502);
or UO_1248 (O_1248,N_9357,N_9409);
nand UO_1249 (O_1249,N_9698,N_9720);
nand UO_1250 (O_1250,N_9159,N_9329);
nor UO_1251 (O_1251,N_9211,N_9908);
nand UO_1252 (O_1252,N_9002,N_9579);
nor UO_1253 (O_1253,N_9348,N_9610);
or UO_1254 (O_1254,N_9490,N_9892);
nor UO_1255 (O_1255,N_9455,N_9874);
or UO_1256 (O_1256,N_9053,N_9711);
and UO_1257 (O_1257,N_9672,N_9374);
nor UO_1258 (O_1258,N_9842,N_9753);
nand UO_1259 (O_1259,N_9204,N_9209);
or UO_1260 (O_1260,N_9992,N_9711);
nand UO_1261 (O_1261,N_9849,N_9308);
or UO_1262 (O_1262,N_9300,N_9123);
and UO_1263 (O_1263,N_9864,N_9787);
and UO_1264 (O_1264,N_9730,N_9092);
and UO_1265 (O_1265,N_9089,N_9074);
or UO_1266 (O_1266,N_9206,N_9272);
nand UO_1267 (O_1267,N_9000,N_9157);
and UO_1268 (O_1268,N_9078,N_9593);
or UO_1269 (O_1269,N_9379,N_9945);
nand UO_1270 (O_1270,N_9816,N_9296);
nand UO_1271 (O_1271,N_9255,N_9929);
and UO_1272 (O_1272,N_9941,N_9621);
or UO_1273 (O_1273,N_9376,N_9217);
nand UO_1274 (O_1274,N_9279,N_9001);
nor UO_1275 (O_1275,N_9112,N_9653);
nand UO_1276 (O_1276,N_9182,N_9374);
or UO_1277 (O_1277,N_9509,N_9372);
and UO_1278 (O_1278,N_9940,N_9777);
nor UO_1279 (O_1279,N_9302,N_9196);
and UO_1280 (O_1280,N_9889,N_9335);
nand UO_1281 (O_1281,N_9269,N_9033);
nor UO_1282 (O_1282,N_9524,N_9370);
or UO_1283 (O_1283,N_9156,N_9731);
nand UO_1284 (O_1284,N_9814,N_9258);
and UO_1285 (O_1285,N_9054,N_9644);
or UO_1286 (O_1286,N_9981,N_9474);
nor UO_1287 (O_1287,N_9801,N_9337);
nor UO_1288 (O_1288,N_9016,N_9329);
and UO_1289 (O_1289,N_9547,N_9694);
nor UO_1290 (O_1290,N_9586,N_9539);
nand UO_1291 (O_1291,N_9342,N_9508);
and UO_1292 (O_1292,N_9821,N_9908);
or UO_1293 (O_1293,N_9507,N_9130);
nand UO_1294 (O_1294,N_9425,N_9540);
and UO_1295 (O_1295,N_9661,N_9083);
and UO_1296 (O_1296,N_9764,N_9771);
and UO_1297 (O_1297,N_9190,N_9842);
or UO_1298 (O_1298,N_9257,N_9276);
and UO_1299 (O_1299,N_9576,N_9233);
or UO_1300 (O_1300,N_9385,N_9129);
and UO_1301 (O_1301,N_9902,N_9155);
nand UO_1302 (O_1302,N_9165,N_9523);
or UO_1303 (O_1303,N_9550,N_9211);
and UO_1304 (O_1304,N_9572,N_9001);
and UO_1305 (O_1305,N_9555,N_9638);
nor UO_1306 (O_1306,N_9436,N_9676);
and UO_1307 (O_1307,N_9198,N_9867);
nand UO_1308 (O_1308,N_9448,N_9420);
or UO_1309 (O_1309,N_9826,N_9536);
nand UO_1310 (O_1310,N_9864,N_9323);
nand UO_1311 (O_1311,N_9759,N_9603);
and UO_1312 (O_1312,N_9114,N_9981);
or UO_1313 (O_1313,N_9637,N_9272);
and UO_1314 (O_1314,N_9346,N_9180);
nand UO_1315 (O_1315,N_9188,N_9110);
nor UO_1316 (O_1316,N_9781,N_9700);
or UO_1317 (O_1317,N_9831,N_9988);
or UO_1318 (O_1318,N_9223,N_9764);
and UO_1319 (O_1319,N_9727,N_9600);
or UO_1320 (O_1320,N_9694,N_9800);
and UO_1321 (O_1321,N_9034,N_9393);
or UO_1322 (O_1322,N_9744,N_9769);
nor UO_1323 (O_1323,N_9280,N_9580);
and UO_1324 (O_1324,N_9971,N_9729);
or UO_1325 (O_1325,N_9227,N_9826);
nor UO_1326 (O_1326,N_9240,N_9816);
and UO_1327 (O_1327,N_9876,N_9549);
or UO_1328 (O_1328,N_9376,N_9303);
or UO_1329 (O_1329,N_9470,N_9685);
nand UO_1330 (O_1330,N_9356,N_9313);
nor UO_1331 (O_1331,N_9977,N_9770);
or UO_1332 (O_1332,N_9070,N_9906);
nor UO_1333 (O_1333,N_9270,N_9528);
or UO_1334 (O_1334,N_9003,N_9767);
nand UO_1335 (O_1335,N_9507,N_9378);
nand UO_1336 (O_1336,N_9496,N_9934);
nand UO_1337 (O_1337,N_9761,N_9039);
and UO_1338 (O_1338,N_9441,N_9189);
and UO_1339 (O_1339,N_9593,N_9531);
or UO_1340 (O_1340,N_9895,N_9723);
or UO_1341 (O_1341,N_9560,N_9133);
nor UO_1342 (O_1342,N_9549,N_9483);
and UO_1343 (O_1343,N_9606,N_9406);
or UO_1344 (O_1344,N_9431,N_9002);
xnor UO_1345 (O_1345,N_9143,N_9255);
nand UO_1346 (O_1346,N_9289,N_9130);
or UO_1347 (O_1347,N_9844,N_9842);
or UO_1348 (O_1348,N_9105,N_9584);
nor UO_1349 (O_1349,N_9387,N_9835);
nor UO_1350 (O_1350,N_9645,N_9706);
and UO_1351 (O_1351,N_9190,N_9248);
or UO_1352 (O_1352,N_9302,N_9722);
nor UO_1353 (O_1353,N_9815,N_9100);
nor UO_1354 (O_1354,N_9320,N_9310);
or UO_1355 (O_1355,N_9694,N_9367);
and UO_1356 (O_1356,N_9836,N_9510);
nor UO_1357 (O_1357,N_9295,N_9004);
or UO_1358 (O_1358,N_9529,N_9324);
nand UO_1359 (O_1359,N_9978,N_9788);
nor UO_1360 (O_1360,N_9694,N_9967);
and UO_1361 (O_1361,N_9420,N_9277);
nand UO_1362 (O_1362,N_9289,N_9208);
nand UO_1363 (O_1363,N_9082,N_9169);
or UO_1364 (O_1364,N_9782,N_9462);
and UO_1365 (O_1365,N_9757,N_9184);
nand UO_1366 (O_1366,N_9081,N_9061);
or UO_1367 (O_1367,N_9271,N_9764);
or UO_1368 (O_1368,N_9090,N_9365);
nand UO_1369 (O_1369,N_9327,N_9137);
or UO_1370 (O_1370,N_9947,N_9232);
nor UO_1371 (O_1371,N_9073,N_9740);
nor UO_1372 (O_1372,N_9538,N_9214);
and UO_1373 (O_1373,N_9361,N_9785);
nor UO_1374 (O_1374,N_9552,N_9339);
nand UO_1375 (O_1375,N_9204,N_9604);
nand UO_1376 (O_1376,N_9823,N_9523);
nand UO_1377 (O_1377,N_9999,N_9751);
nand UO_1378 (O_1378,N_9483,N_9111);
nor UO_1379 (O_1379,N_9865,N_9917);
nor UO_1380 (O_1380,N_9140,N_9646);
nand UO_1381 (O_1381,N_9229,N_9891);
or UO_1382 (O_1382,N_9146,N_9507);
or UO_1383 (O_1383,N_9223,N_9213);
or UO_1384 (O_1384,N_9862,N_9223);
nor UO_1385 (O_1385,N_9177,N_9312);
or UO_1386 (O_1386,N_9587,N_9764);
and UO_1387 (O_1387,N_9982,N_9727);
nand UO_1388 (O_1388,N_9024,N_9904);
or UO_1389 (O_1389,N_9695,N_9111);
and UO_1390 (O_1390,N_9304,N_9922);
nand UO_1391 (O_1391,N_9873,N_9595);
nor UO_1392 (O_1392,N_9615,N_9952);
nand UO_1393 (O_1393,N_9301,N_9371);
nor UO_1394 (O_1394,N_9229,N_9609);
nor UO_1395 (O_1395,N_9291,N_9238);
nand UO_1396 (O_1396,N_9605,N_9961);
nor UO_1397 (O_1397,N_9427,N_9936);
and UO_1398 (O_1398,N_9751,N_9237);
nor UO_1399 (O_1399,N_9822,N_9159);
and UO_1400 (O_1400,N_9377,N_9467);
or UO_1401 (O_1401,N_9461,N_9781);
nand UO_1402 (O_1402,N_9346,N_9802);
and UO_1403 (O_1403,N_9594,N_9698);
nor UO_1404 (O_1404,N_9776,N_9416);
xor UO_1405 (O_1405,N_9204,N_9375);
or UO_1406 (O_1406,N_9682,N_9729);
nand UO_1407 (O_1407,N_9680,N_9917);
and UO_1408 (O_1408,N_9937,N_9982);
nand UO_1409 (O_1409,N_9400,N_9462);
nor UO_1410 (O_1410,N_9414,N_9504);
nand UO_1411 (O_1411,N_9678,N_9679);
nand UO_1412 (O_1412,N_9569,N_9403);
or UO_1413 (O_1413,N_9849,N_9533);
or UO_1414 (O_1414,N_9437,N_9944);
nor UO_1415 (O_1415,N_9558,N_9223);
nor UO_1416 (O_1416,N_9886,N_9395);
nor UO_1417 (O_1417,N_9508,N_9098);
nand UO_1418 (O_1418,N_9188,N_9097);
nor UO_1419 (O_1419,N_9974,N_9985);
nand UO_1420 (O_1420,N_9584,N_9143);
or UO_1421 (O_1421,N_9072,N_9447);
xor UO_1422 (O_1422,N_9375,N_9660);
and UO_1423 (O_1423,N_9287,N_9650);
nand UO_1424 (O_1424,N_9076,N_9926);
nor UO_1425 (O_1425,N_9912,N_9078);
and UO_1426 (O_1426,N_9412,N_9020);
nand UO_1427 (O_1427,N_9712,N_9240);
nor UO_1428 (O_1428,N_9982,N_9448);
nand UO_1429 (O_1429,N_9945,N_9096);
nand UO_1430 (O_1430,N_9422,N_9650);
and UO_1431 (O_1431,N_9538,N_9872);
nand UO_1432 (O_1432,N_9195,N_9858);
nor UO_1433 (O_1433,N_9695,N_9092);
and UO_1434 (O_1434,N_9220,N_9319);
or UO_1435 (O_1435,N_9088,N_9725);
and UO_1436 (O_1436,N_9327,N_9560);
and UO_1437 (O_1437,N_9525,N_9996);
nor UO_1438 (O_1438,N_9675,N_9008);
or UO_1439 (O_1439,N_9828,N_9978);
and UO_1440 (O_1440,N_9092,N_9762);
nor UO_1441 (O_1441,N_9521,N_9238);
or UO_1442 (O_1442,N_9952,N_9083);
and UO_1443 (O_1443,N_9124,N_9722);
and UO_1444 (O_1444,N_9452,N_9266);
nand UO_1445 (O_1445,N_9114,N_9972);
nor UO_1446 (O_1446,N_9819,N_9272);
nor UO_1447 (O_1447,N_9310,N_9599);
nand UO_1448 (O_1448,N_9094,N_9376);
or UO_1449 (O_1449,N_9709,N_9300);
nand UO_1450 (O_1450,N_9710,N_9074);
or UO_1451 (O_1451,N_9729,N_9935);
nand UO_1452 (O_1452,N_9470,N_9777);
or UO_1453 (O_1453,N_9010,N_9949);
nor UO_1454 (O_1454,N_9545,N_9291);
or UO_1455 (O_1455,N_9155,N_9324);
and UO_1456 (O_1456,N_9089,N_9836);
nor UO_1457 (O_1457,N_9799,N_9917);
nand UO_1458 (O_1458,N_9458,N_9345);
nand UO_1459 (O_1459,N_9697,N_9309);
nand UO_1460 (O_1460,N_9834,N_9031);
and UO_1461 (O_1461,N_9947,N_9023);
or UO_1462 (O_1462,N_9390,N_9960);
nor UO_1463 (O_1463,N_9077,N_9154);
or UO_1464 (O_1464,N_9747,N_9208);
xor UO_1465 (O_1465,N_9250,N_9383);
and UO_1466 (O_1466,N_9763,N_9249);
nand UO_1467 (O_1467,N_9007,N_9018);
or UO_1468 (O_1468,N_9028,N_9307);
nor UO_1469 (O_1469,N_9321,N_9394);
xor UO_1470 (O_1470,N_9620,N_9703);
or UO_1471 (O_1471,N_9145,N_9910);
nor UO_1472 (O_1472,N_9518,N_9476);
and UO_1473 (O_1473,N_9873,N_9911);
nor UO_1474 (O_1474,N_9763,N_9217);
or UO_1475 (O_1475,N_9525,N_9617);
nor UO_1476 (O_1476,N_9905,N_9611);
or UO_1477 (O_1477,N_9438,N_9979);
or UO_1478 (O_1478,N_9978,N_9235);
nor UO_1479 (O_1479,N_9300,N_9062);
nand UO_1480 (O_1480,N_9906,N_9733);
nor UO_1481 (O_1481,N_9565,N_9209);
nand UO_1482 (O_1482,N_9299,N_9560);
nor UO_1483 (O_1483,N_9815,N_9395);
and UO_1484 (O_1484,N_9797,N_9033);
nand UO_1485 (O_1485,N_9575,N_9182);
or UO_1486 (O_1486,N_9709,N_9250);
nand UO_1487 (O_1487,N_9847,N_9322);
nor UO_1488 (O_1488,N_9222,N_9233);
and UO_1489 (O_1489,N_9816,N_9484);
nor UO_1490 (O_1490,N_9054,N_9052);
and UO_1491 (O_1491,N_9037,N_9560);
nor UO_1492 (O_1492,N_9381,N_9630);
or UO_1493 (O_1493,N_9788,N_9843);
and UO_1494 (O_1494,N_9105,N_9625);
nor UO_1495 (O_1495,N_9475,N_9039);
nand UO_1496 (O_1496,N_9536,N_9813);
nand UO_1497 (O_1497,N_9345,N_9754);
and UO_1498 (O_1498,N_9736,N_9688);
nor UO_1499 (O_1499,N_9673,N_9748);
endmodule