module basic_3000_30000_3500_25_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_2900,In_2178);
or U1 (N_1,In_1990,In_579);
and U2 (N_2,In_722,In_891);
and U3 (N_3,In_578,In_2384);
nand U4 (N_4,In_2672,In_1014);
nor U5 (N_5,In_2229,In_501);
nand U6 (N_6,In_2017,In_623);
and U7 (N_7,In_1433,In_1785);
and U8 (N_8,In_2508,In_2997);
nand U9 (N_9,In_2046,In_2744);
xor U10 (N_10,In_365,In_1517);
nor U11 (N_11,In_947,In_1415);
and U12 (N_12,In_2954,In_1260);
xnor U13 (N_13,In_1833,In_2398);
nor U14 (N_14,In_1632,In_1993);
and U15 (N_15,In_1252,In_1406);
and U16 (N_16,In_2291,In_2628);
nor U17 (N_17,In_2801,In_2994);
nand U18 (N_18,In_1427,In_1533);
nor U19 (N_19,In_2743,In_435);
nand U20 (N_20,In_702,In_1503);
nor U21 (N_21,In_2352,In_360);
nand U22 (N_22,In_2147,In_325);
xor U23 (N_23,In_1642,In_1808);
xor U24 (N_24,In_212,In_2258);
nand U25 (N_25,In_405,In_1047);
xnor U26 (N_26,In_1732,In_362);
or U27 (N_27,In_616,In_843);
and U28 (N_28,In_204,In_606);
nand U29 (N_29,In_2941,In_709);
nand U30 (N_30,In_2251,In_402);
nand U31 (N_31,In_628,In_163);
or U32 (N_32,In_15,In_460);
or U33 (N_33,In_1128,In_525);
xnor U34 (N_34,In_1112,In_368);
or U35 (N_35,In_1222,In_2795);
or U36 (N_36,In_1444,In_2572);
nor U37 (N_37,In_1970,In_1582);
and U38 (N_38,In_775,In_965);
and U39 (N_39,In_1174,In_1940);
nand U40 (N_40,In_1836,In_1566);
nand U41 (N_41,In_230,In_2759);
or U42 (N_42,In_776,In_1861);
and U43 (N_43,In_1109,In_1914);
nor U44 (N_44,In_1819,In_2632);
xor U45 (N_45,In_2138,In_109);
and U46 (N_46,In_189,In_2089);
and U47 (N_47,In_1285,In_2326);
or U48 (N_48,In_737,In_608);
or U49 (N_49,In_2282,In_651);
nor U50 (N_50,In_1609,In_1719);
and U51 (N_51,In_206,In_1775);
or U52 (N_52,In_2956,In_152);
and U53 (N_53,In_428,In_2187);
xor U54 (N_54,In_1324,In_2818);
nand U55 (N_55,In_619,In_2085);
nor U56 (N_56,In_2880,In_763);
nor U57 (N_57,In_1410,In_1391);
and U58 (N_58,In_2630,In_139);
or U59 (N_59,In_2652,In_626);
or U60 (N_60,In_71,In_994);
xnor U61 (N_61,In_2848,In_1598);
xnor U62 (N_62,In_2431,In_65);
nand U63 (N_63,In_1113,In_1188);
xor U64 (N_64,In_2543,In_2819);
xnor U65 (N_65,In_2936,In_2365);
and U66 (N_66,In_129,In_2532);
or U67 (N_67,In_423,In_1089);
or U68 (N_68,In_2295,In_1825);
nor U69 (N_69,In_1245,In_2617);
xnor U70 (N_70,In_770,In_1382);
and U71 (N_71,In_1064,In_2175);
or U72 (N_72,In_1526,In_505);
nand U73 (N_73,In_2306,In_1308);
or U74 (N_74,In_1803,In_794);
xnor U75 (N_75,In_2338,In_2739);
nor U76 (N_76,In_581,In_1232);
and U77 (N_77,In_1122,In_2377);
and U78 (N_78,In_1700,In_1886);
and U79 (N_79,In_1067,In_599);
xnor U80 (N_80,In_157,In_2664);
nand U81 (N_81,In_2287,In_2101);
nand U82 (N_82,In_2613,In_340);
xor U83 (N_83,In_2981,In_986);
or U84 (N_84,In_2144,In_827);
or U85 (N_85,In_2717,In_2845);
and U86 (N_86,In_1053,In_614);
or U87 (N_87,In_749,In_231);
or U88 (N_88,In_2515,In_2719);
nor U89 (N_89,In_2885,In_1054);
or U90 (N_90,In_1066,In_2053);
xnor U91 (N_91,In_2953,In_1393);
or U92 (N_92,In_2931,In_2857);
nand U93 (N_93,In_2914,In_1076);
and U94 (N_94,In_2180,In_429);
nor U95 (N_95,In_2789,In_633);
nor U96 (N_96,In_264,In_2191);
and U97 (N_97,In_1622,In_2689);
or U98 (N_98,In_507,In_558);
nand U99 (N_99,In_2999,In_130);
xor U100 (N_100,In_1627,In_318);
xor U101 (N_101,In_876,In_1579);
xor U102 (N_102,In_1491,In_1860);
nand U103 (N_103,In_1906,In_1556);
xnor U104 (N_104,In_1593,In_22);
and U105 (N_105,In_2260,In_2292);
nor U106 (N_106,In_1866,In_1704);
or U107 (N_107,In_312,In_458);
or U108 (N_108,In_2776,In_297);
nand U109 (N_109,In_2124,In_2627);
nor U110 (N_110,In_2379,In_2971);
or U111 (N_111,In_1212,In_2247);
xnor U112 (N_112,In_2786,In_495);
nand U113 (N_113,In_25,In_2127);
xnor U114 (N_114,In_2206,In_2047);
xnor U115 (N_115,In_2351,In_1639);
nor U116 (N_116,In_2596,In_2711);
nand U117 (N_117,In_1399,In_2509);
or U118 (N_118,In_474,In_2182);
nor U119 (N_119,In_1062,In_2959);
nand U120 (N_120,In_693,In_942);
nor U121 (N_121,In_1253,In_2582);
xor U122 (N_122,In_132,In_2902);
xor U123 (N_123,In_506,In_2969);
nor U124 (N_124,In_1030,In_669);
nor U125 (N_125,In_1500,In_1000);
nand U126 (N_126,In_2575,In_295);
or U127 (N_127,In_1121,In_82);
xor U128 (N_128,In_1226,In_1730);
and U129 (N_129,In_2561,In_2858);
or U130 (N_130,In_420,In_2346);
or U131 (N_131,In_2807,In_149);
or U132 (N_132,In_470,In_1304);
and U133 (N_133,In_1978,In_2335);
nand U134 (N_134,In_1981,In_1681);
or U135 (N_135,In_1110,In_1896);
nor U136 (N_136,In_1799,In_2141);
xor U137 (N_137,In_145,In_2656);
or U138 (N_138,In_2761,In_85);
or U139 (N_139,In_2299,In_2502);
xor U140 (N_140,In_92,In_2531);
xor U141 (N_141,In_728,In_418);
nand U142 (N_142,In_427,In_2771);
or U143 (N_143,In_1265,In_2074);
xor U144 (N_144,In_1046,In_1138);
and U145 (N_145,In_24,In_1839);
or U146 (N_146,In_896,In_530);
xor U147 (N_147,In_807,In_2076);
nor U148 (N_148,In_989,In_2951);
nand U149 (N_149,In_1498,In_1216);
nand U150 (N_150,In_851,In_1810);
xnor U151 (N_151,In_1457,In_609);
nor U152 (N_152,In_1220,In_1354);
nor U153 (N_153,In_1247,In_198);
or U154 (N_154,In_2888,In_670);
and U155 (N_155,In_2906,In_1045);
or U156 (N_156,In_1327,In_1079);
nor U157 (N_157,In_2010,In_2469);
nand U158 (N_158,In_2750,In_91);
nand U159 (N_159,In_567,In_2232);
nand U160 (N_160,In_2773,In_2334);
nor U161 (N_161,In_2648,In_1348);
and U162 (N_162,In_2035,In_1150);
or U163 (N_163,In_2444,In_1152);
nand U164 (N_164,In_2714,In_1596);
xnor U165 (N_165,In_821,In_238);
xnor U166 (N_166,In_2005,In_1873);
nor U167 (N_167,In_16,In_945);
or U168 (N_168,In_1749,In_921);
nor U169 (N_169,In_354,In_371);
and U170 (N_170,In_269,In_2043);
or U171 (N_171,In_1256,In_115);
xor U172 (N_172,In_419,In_1326);
or U173 (N_173,In_1543,In_1346);
nand U174 (N_174,In_755,In_2654);
or U175 (N_175,In_4,In_836);
xor U176 (N_176,In_2257,In_1548);
or U177 (N_177,In_2489,In_2310);
nand U178 (N_178,In_1040,In_298);
and U179 (N_179,In_2945,In_2174);
nand U180 (N_180,In_1276,In_1359);
nand U181 (N_181,In_1287,In_1170);
and U182 (N_182,In_2546,In_1300);
and U183 (N_183,In_216,In_188);
nor U184 (N_184,In_200,In_1698);
nor U185 (N_185,In_1997,In_2983);
nand U186 (N_186,In_1653,In_1360);
xnor U187 (N_187,In_1065,In_2115);
and U188 (N_188,In_2383,In_2316);
nand U189 (N_189,In_1384,In_2840);
and U190 (N_190,In_2006,In_2782);
and U191 (N_191,In_23,In_2219);
nor U192 (N_192,In_2021,In_485);
or U193 (N_193,In_2712,In_484);
and U194 (N_194,In_736,In_2146);
nor U195 (N_195,In_2143,In_158);
or U196 (N_196,In_1646,In_676);
or U197 (N_197,In_1025,In_476);
and U198 (N_198,In_1712,In_2312);
or U199 (N_199,In_2849,In_2638);
nor U200 (N_200,In_1036,In_475);
xnor U201 (N_201,In_1760,In_950);
nor U202 (N_202,In_2430,In_2152);
nand U203 (N_203,In_33,In_2909);
nor U204 (N_204,In_1599,In_1342);
nor U205 (N_205,In_1806,In_1830);
or U206 (N_206,In_124,In_125);
nor U207 (N_207,In_723,In_2121);
nor U208 (N_208,In_2093,In_1280);
or U209 (N_209,In_2067,In_834);
and U210 (N_210,In_1194,In_1388);
and U211 (N_211,In_607,In_2723);
and U212 (N_212,In_161,In_2498);
nor U213 (N_213,In_1716,In_746);
xor U214 (N_214,In_560,In_1748);
nand U215 (N_215,In_2249,In_2783);
and U216 (N_216,In_2978,In_1137);
or U217 (N_217,In_2420,In_1883);
nand U218 (N_218,In_744,In_1507);
nand U219 (N_219,In_2393,In_1925);
and U220 (N_220,In_1920,In_769);
nand U221 (N_221,In_1602,In_27);
nand U222 (N_222,In_2539,In_398);
xnor U223 (N_223,In_374,In_816);
and U224 (N_224,In_1394,In_1032);
nor U225 (N_225,In_454,In_642);
nand U226 (N_226,In_1288,In_2262);
nor U227 (N_227,In_1186,In_147);
nand U228 (N_228,In_1330,In_462);
and U229 (N_229,In_1196,In_1837);
xnor U230 (N_230,In_2185,In_1571);
nor U231 (N_231,In_399,In_281);
and U232 (N_232,In_2580,In_2687);
or U233 (N_233,In_1910,In_829);
nor U234 (N_234,In_2039,In_814);
nor U235 (N_235,In_520,In_2374);
nor U236 (N_236,In_293,In_1888);
or U237 (N_237,In_894,In_1262);
nor U238 (N_238,In_1984,In_1950);
nand U239 (N_239,In_881,In_688);
and U240 (N_240,In_1518,In_972);
xor U241 (N_241,In_548,In_1558);
nor U242 (N_242,In_856,In_2946);
nand U243 (N_243,In_639,In_1044);
nand U244 (N_244,In_98,In_2401);
nor U245 (N_245,In_1481,In_1091);
and U246 (N_246,In_596,In_1017);
xnor U247 (N_247,In_2296,In_2872);
xor U248 (N_248,In_2423,In_1553);
and U249 (N_249,In_2943,In_960);
or U250 (N_250,In_2566,In_394);
xor U251 (N_251,In_654,In_2002);
or U252 (N_252,In_2903,In_2955);
and U253 (N_253,In_2390,In_1859);
or U254 (N_254,In_602,In_378);
nor U255 (N_255,In_2032,In_1647);
nor U256 (N_256,In_1721,In_1880);
xnor U257 (N_257,In_2504,In_234);
nand U258 (N_258,In_760,In_445);
nand U259 (N_259,In_557,In_438);
nor U260 (N_260,In_1502,In_1012);
and U261 (N_261,In_317,In_1705);
or U262 (N_262,In_90,In_2988);
or U263 (N_263,In_267,In_659);
and U264 (N_264,In_1258,In_1419);
and U265 (N_265,In_1244,In_1001);
or U266 (N_266,In_1477,In_1918);
nand U267 (N_267,In_1977,In_2844);
nor U268 (N_268,In_215,In_1691);
nor U269 (N_269,In_1772,In_1878);
nand U270 (N_270,In_364,In_933);
nand U271 (N_271,In_931,In_251);
nor U272 (N_272,In_2547,In_1103);
and U273 (N_273,In_1926,In_1205);
xnor U274 (N_274,In_2403,In_1009);
xnor U275 (N_275,In_2441,In_146);
or U276 (N_276,In_1395,In_1960);
xor U277 (N_277,In_1461,In_575);
and U278 (N_278,In_652,In_2164);
or U279 (N_279,In_1497,In_201);
or U280 (N_280,In_2796,In_1423);
nor U281 (N_281,In_2195,In_2462);
xor U282 (N_282,In_235,In_672);
nand U283 (N_283,In_847,In_237);
or U284 (N_284,In_375,In_2438);
nand U285 (N_285,In_143,In_486);
nand U286 (N_286,In_2803,In_202);
nand U287 (N_287,In_2658,In_912);
and U288 (N_288,In_2137,In_291);
and U289 (N_289,In_860,In_1147);
nand U290 (N_290,In_2736,In_1532);
or U291 (N_291,In_2072,In_2019);
nand U292 (N_292,In_96,In_2594);
and U293 (N_293,In_561,In_2813);
and U294 (N_294,In_1093,In_1488);
and U295 (N_295,In_1398,In_1962);
and U296 (N_296,In_1893,In_753);
nor U297 (N_297,In_1356,In_2491);
or U298 (N_298,In_2823,In_1132);
or U299 (N_299,In_2563,In_2449);
nand U300 (N_300,In_2530,In_1104);
or U301 (N_301,In_1658,In_1235);
nor U302 (N_302,In_153,In_2995);
nor U303 (N_303,In_2330,In_2173);
nand U304 (N_304,In_186,In_1277);
and U305 (N_305,In_2843,In_667);
and U306 (N_306,In_636,In_1190);
nor U307 (N_307,In_2912,In_840);
xor U308 (N_308,In_439,In_1329);
nand U309 (N_309,In_1297,In_1915);
xnor U310 (N_310,In_1052,In_2402);
and U311 (N_311,In_1849,In_2757);
nand U312 (N_312,In_1303,In_1504);
and U313 (N_313,In_8,In_275);
and U314 (N_314,In_958,In_254);
nor U315 (N_315,In_1745,In_2192);
nand U316 (N_316,In_1793,In_1086);
and U317 (N_317,In_2935,In_94);
nor U318 (N_318,In_762,In_2079);
nand U319 (N_319,In_2694,In_2741);
nand U320 (N_320,In_696,In_1968);
nand U321 (N_321,In_845,In_1248);
nand U322 (N_322,In_612,In_338);
nand U323 (N_323,In_219,In_761);
xnor U324 (N_324,In_2463,In_1299);
nor U325 (N_325,In_1015,In_1733);
or U326 (N_326,In_349,In_1027);
nand U327 (N_327,In_694,In_2184);
or U328 (N_328,In_2389,In_2125);
and U329 (N_329,In_895,In_1161);
and U330 (N_330,In_617,In_2356);
nand U331 (N_331,In_2114,In_819);
or U332 (N_332,In_629,In_1416);
xor U333 (N_333,In_2339,In_1219);
or U334 (N_334,In_1075,In_882);
nor U335 (N_335,In_2060,In_552);
nor U336 (N_336,In_2298,In_593);
xnor U337 (N_337,In_514,In_1542);
or U338 (N_338,In_1637,In_893);
nand U339 (N_339,In_590,In_2793);
or U340 (N_340,In_1856,In_1355);
and U341 (N_341,In_1126,In_1770);
nand U342 (N_342,In_2871,In_2998);
nand U343 (N_343,In_2070,In_1870);
nor U344 (N_344,In_2418,In_2081);
and U345 (N_345,In_1955,In_1757);
or U346 (N_346,In_592,In_2371);
nand U347 (N_347,In_2932,In_2183);
or U348 (N_348,In_1845,In_757);
or U349 (N_349,In_2745,In_711);
or U350 (N_350,In_1520,In_1350);
or U351 (N_351,In_1016,In_366);
or U352 (N_352,In_527,In_1272);
nor U353 (N_353,In_1117,In_1595);
and U354 (N_354,In_180,In_333);
or U355 (N_355,In_1453,In_2023);
and U356 (N_356,In_1315,In_535);
or U357 (N_357,In_1485,In_2618);
nand U358 (N_358,In_1885,In_2601);
nand U359 (N_359,In_2920,In_313);
nand U360 (N_360,In_2243,In_1451);
xor U361 (N_361,In_1679,In_1411);
nand U362 (N_362,In_1335,In_1494);
xnor U363 (N_363,In_1051,In_1428);
or U364 (N_364,In_1751,In_1546);
xor U365 (N_365,In_2804,In_1165);
nor U366 (N_366,In_1209,In_388);
or U367 (N_367,In_77,In_2369);
xor U368 (N_368,In_565,In_2753);
nand U369 (N_369,In_2841,In_2241);
or U370 (N_370,In_492,In_1999);
nor U371 (N_371,In_2859,In_1203);
or U372 (N_372,In_1264,In_862);
and U373 (N_373,In_2160,In_1816);
or U374 (N_374,In_2036,In_2685);
xnor U375 (N_375,In_1992,In_334);
nor U376 (N_376,In_546,In_1710);
or U377 (N_377,In_467,In_885);
or U378 (N_378,In_1765,In_1690);
nand U379 (N_379,In_2140,In_1921);
nor U380 (N_380,In_1929,In_308);
or U381 (N_381,In_1241,In_2421);
or U382 (N_382,In_955,In_2790);
nand U383 (N_383,In_220,In_2105);
or U384 (N_384,In_222,In_2751);
xnor U385 (N_385,In_1515,In_1077);
xnor U386 (N_386,In_2011,In_2817);
or U387 (N_387,In_710,In_745);
nand U388 (N_388,In_613,In_2478);
or U389 (N_389,In_766,In_1641);
nor U390 (N_390,In_961,In_1208);
and U391 (N_391,In_825,In_2944);
nand U392 (N_392,In_2386,In_60);
nand U393 (N_393,In_2680,In_585);
and U394 (N_394,In_2993,In_2025);
nor U395 (N_395,In_526,In_1207);
and U396 (N_396,In_1414,In_857);
or U397 (N_397,In_1460,In_101);
xor U398 (N_398,In_1928,In_2308);
nor U399 (N_399,In_1363,In_321);
and U400 (N_400,In_866,In_409);
nand U401 (N_401,In_1635,In_2647);
nand U402 (N_402,In_1843,In_793);
xor U403 (N_403,In_302,In_57);
xnor U404 (N_404,In_1200,In_1204);
or U405 (N_405,In_936,In_647);
nand U406 (N_406,In_1796,In_957);
xor U407 (N_407,In_2448,In_724);
nor U408 (N_408,In_1358,In_2758);
nand U409 (N_409,In_2791,In_566);
and U410 (N_410,In_1787,In_1662);
or U411 (N_411,In_523,In_1167);
nand U412 (N_412,In_214,In_270);
nand U413 (N_413,In_2977,In_880);
and U414 (N_414,In_2474,In_1286);
nand U415 (N_415,In_2281,In_690);
or U416 (N_416,In_343,In_1755);
or U417 (N_417,In_2847,In_977);
nor U418 (N_418,In_1357,In_2194);
and U419 (N_419,In_30,In_240);
or U420 (N_420,In_311,In_2106);
xnor U421 (N_421,In_49,In_2128);
or U422 (N_422,In_2715,In_2240);
nor U423 (N_423,In_1740,In_964);
and U424 (N_424,In_2787,In_1344);
or U425 (N_425,In_352,In_446);
nor U426 (N_426,In_1597,In_2304);
nand U427 (N_427,In_2446,In_292);
xor U428 (N_428,In_2550,In_1474);
nor U429 (N_429,In_1743,In_1448);
and U430 (N_430,In_2354,In_1364);
or U431 (N_431,In_2865,In_1580);
nor U432 (N_432,In_1935,In_1851);
xnor U433 (N_433,In_226,In_195);
nor U434 (N_434,In_512,In_841);
nor U435 (N_435,In_1664,In_1169);
nor U436 (N_436,In_1043,In_1100);
nor U437 (N_437,In_1058,In_2022);
or U438 (N_438,In_729,In_1549);
nand U439 (N_439,In_2086,In_2591);
or U440 (N_440,In_1055,In_2684);
nor U441 (N_441,In_634,In_2533);
nand U442 (N_442,In_940,In_2815);
or U443 (N_443,In_871,In_2831);
nand U444 (N_444,In_1123,In_2838);
or U445 (N_445,In_1447,In_2661);
nor U446 (N_446,In_1754,In_284);
and U447 (N_447,In_2666,In_1007);
or U448 (N_448,In_2657,In_2230);
nand U449 (N_449,In_441,In_1413);
and U450 (N_450,In_779,In_73);
xnor U451 (N_451,In_2333,In_213);
and U452 (N_452,In_2641,In_1302);
nand U453 (N_453,In_1496,In_1547);
and U454 (N_454,In_1080,In_2792);
nand U455 (N_455,In_2690,In_1758);
and U456 (N_456,In_416,In_2560);
xor U457 (N_457,In_2785,In_516);
nand U458 (N_458,In_781,In_2899);
xnor U459 (N_459,In_20,In_2742);
or U460 (N_460,In_2511,In_2863);
and U461 (N_461,In_232,In_2860);
nor U462 (N_462,In_1701,In_582);
nor U463 (N_463,In_2665,In_183);
nor U464 (N_464,In_949,In_2397);
nor U465 (N_465,In_2579,In_778);
xnor U466 (N_466,In_1848,In_2604);
nand U467 (N_467,In_517,In_1724);
or U468 (N_468,In_353,In_389);
xnor U469 (N_469,In_925,In_598);
or U470 (N_470,In_2810,In_2486);
nor U471 (N_471,In_2145,In_531);
nor U472 (N_472,In_1750,In_245);
nor U473 (N_473,In_498,In_69);
or U474 (N_474,In_2487,In_1088);
xor U475 (N_475,In_2842,In_286);
nor U476 (N_476,In_1236,In_1270);
xnor U477 (N_477,In_1107,In_2827);
nand U478 (N_478,In_417,In_2189);
nor U479 (N_479,In_1636,In_828);
or U480 (N_480,In_1096,In_534);
nand U481 (N_481,In_1116,In_1901);
and U482 (N_482,In_2698,In_837);
and U483 (N_483,In_946,In_1242);
nand U484 (N_484,In_1267,In_2571);
xor U485 (N_485,In_2907,In_2479);
nor U486 (N_486,In_1835,In_2405);
and U487 (N_487,In_2001,In_1035);
nand U488 (N_488,In_190,In_1390);
and U489 (N_489,In_255,In_2557);
nor U490 (N_490,In_773,In_2974);
and U491 (N_491,In_1971,In_1687);
nand U492 (N_492,In_2780,In_2378);
nand U493 (N_493,In_1889,In_2166);
nand U494 (N_494,In_330,In_1033);
or U495 (N_495,In_2452,In_2718);
nor U496 (N_496,In_547,In_2967);
nor U497 (N_497,In_1604,In_1155);
nand U498 (N_498,In_663,In_2014);
xnor U499 (N_499,In_1590,In_310);
and U500 (N_500,In_545,In_2204);
nor U501 (N_501,In_2426,In_2904);
nand U502 (N_502,In_1289,In_357);
nand U503 (N_503,In_2372,In_1470);
xnor U504 (N_504,In_971,In_635);
nand U505 (N_505,In_2467,In_2190);
or U506 (N_506,In_2524,In_2455);
xnor U507 (N_507,In_1969,In_1269);
nor U508 (N_508,In_2307,In_1162);
xor U509 (N_509,In_914,In_2197);
xnor U510 (N_510,In_1613,In_155);
nor U511 (N_511,In_849,In_2443);
or U512 (N_512,In_1631,In_621);
xor U513 (N_513,In_2024,In_483);
and U514 (N_514,In_2850,In_256);
nor U515 (N_515,In_2669,In_941);
nor U516 (N_516,In_2071,In_1587);
nor U517 (N_517,In_1818,In_369);
xnor U518 (N_518,In_119,In_733);
nand U519 (N_519,In_1311,In_1605);
or U520 (N_520,In_296,In_391);
and U521 (N_521,In_407,In_2208);
nand U522 (N_522,In_865,In_1625);
xnor U523 (N_523,In_1290,In_861);
nand U524 (N_524,In_1656,In_1373);
nor U525 (N_525,In_1916,In_777);
nand U526 (N_526,In_1156,In_2921);
nand U527 (N_527,In_1811,In_2427);
and U528 (N_528,In_385,In_2061);
nor U529 (N_529,In_11,In_1961);
nand U530 (N_530,In_2054,In_2225);
and U531 (N_531,In_2624,In_764);
nand U532 (N_532,In_2327,In_2088);
and U533 (N_533,In_1168,In_2068);
nor U534 (N_534,In_2324,In_252);
or U535 (N_535,In_167,In_289);
xnor U536 (N_536,In_1805,In_2481);
nand U537 (N_537,In_2623,In_2595);
xor U538 (N_538,In_301,In_846);
and U539 (N_539,In_450,In_2480);
xnor U540 (N_540,In_521,In_122);
xor U541 (N_541,In_1829,In_1259);
nand U542 (N_542,In_2942,In_181);
nand U543 (N_543,In_344,In_2839);
xor U544 (N_544,In_2158,In_1430);
or U545 (N_545,In_2678,In_1567);
or U546 (N_546,In_1184,In_1469);
nor U547 (N_547,In_2413,In_1588);
nand U548 (N_548,In_2118,In_1643);
xor U549 (N_549,In_1817,In_2439);
or U550 (N_550,In_348,In_2768);
and U551 (N_551,In_2492,In_2825);
nor U552 (N_552,In_2535,In_89);
nand U553 (N_553,In_524,In_2037);
or U554 (N_554,In_1004,In_1897);
and U555 (N_555,In_983,In_300);
nor U556 (N_556,In_36,In_191);
and U557 (N_557,In_1367,In_1953);
nor U558 (N_558,In_995,In_236);
xnor U559 (N_559,In_2910,In_1307);
nor U560 (N_560,In_2490,In_1557);
xnor U561 (N_561,In_586,In_1171);
nand U562 (N_562,In_1900,In_67);
or U563 (N_563,In_1694,In_2873);
and U564 (N_564,In_1240,In_997);
and U565 (N_565,In_499,In_2692);
nor U566 (N_566,In_1924,In_1336);
nand U567 (N_567,In_184,In_2012);
or U568 (N_568,In_2055,In_1783);
nand U569 (N_569,In_2248,In_2679);
or U570 (N_570,In_1366,In_2970);
nand U571 (N_571,In_465,In_455);
and U572 (N_572,In_2933,In_782);
or U573 (N_573,In_1437,In_396);
or U574 (N_574,In_414,In_453);
xnor U575 (N_575,In_1099,In_2433);
and U576 (N_576,In_1191,In_2254);
or U577 (N_577,In_488,In_532);
nor U578 (N_578,In_2821,In_2040);
nand U579 (N_579,In_2976,In_2824);
nor U580 (N_580,In_768,In_1943);
nand U581 (N_581,In_641,In_2349);
nand U582 (N_582,In_1487,In_2673);
or U583 (N_583,In_2364,In_1529);
xor U584 (N_584,In_187,In_156);
nor U585 (N_585,In_897,In_1401);
and U586 (N_586,In_1251,In_1478);
nand U587 (N_587,In_350,In_144);
or U588 (N_588,In_2784,In_1446);
or U589 (N_589,In_2056,In_2883);
or U590 (N_590,In_1822,In_2737);
and U591 (N_591,In_1884,In_2422);
or U592 (N_592,In_1957,In_2457);
nor U593 (N_593,In_1050,In_2341);
or U594 (N_594,In_2133,In_2517);
and U595 (N_595,In_1037,In_1141);
nor U596 (N_596,In_655,In_1381);
or U597 (N_597,In_2979,In_1365);
or U598 (N_598,In_1559,In_320);
xnor U599 (N_599,In_2130,In_142);
xor U600 (N_600,In_2930,In_2836);
xor U601 (N_601,In_315,In_41);
nand U602 (N_602,In_888,In_1229);
nor U603 (N_603,In_2551,In_954);
or U604 (N_604,In_393,In_1741);
or U605 (N_605,In_2724,In_1442);
or U606 (N_606,In_2392,In_2642);
or U607 (N_607,In_1183,In_877);
xnor U608 (N_608,In_1143,In_1139);
and U609 (N_609,In_100,In_459);
nand U610 (N_610,In_1024,In_1585);
xor U611 (N_611,In_1111,In_2179);
nor U612 (N_612,In_1118,In_2637);
nand U613 (N_613,In_835,In_2470);
nor U614 (N_614,In_830,In_1490);
or U615 (N_615,In_790,In_2752);
nand U616 (N_616,In_1671,In_345);
and U617 (N_617,In_1946,In_1372);
and U618 (N_618,In_2205,In_1225);
nor U619 (N_619,In_601,In_1792);
nand U620 (N_620,In_241,In_2279);
xor U621 (N_621,In_1407,In_1185);
nor U622 (N_622,In_194,In_2777);
nor U623 (N_623,In_173,In_266);
or U624 (N_624,In_2778,In_2075);
nor U625 (N_625,In_2313,In_351);
nand U626 (N_626,In_1692,In_1257);
xor U627 (N_627,In_261,In_262);
or U628 (N_628,In_471,In_2756);
nand U629 (N_629,In_1341,In_2259);
or U630 (N_630,In_2607,In_886);
xnor U631 (N_631,In_1923,In_1215);
nor U632 (N_632,In_2529,In_1629);
xnor U633 (N_633,In_2963,In_336);
nand U634 (N_634,In_2097,In_1742);
nor U635 (N_635,In_928,In_1931);
or U636 (N_636,In_674,In_1345);
nand U637 (N_637,In_2332,In_2317);
xor U638 (N_638,In_1815,In_346);
nand U639 (N_639,In_2982,In_2830);
nand U640 (N_640,In_2155,In_2980);
xnor U641 (N_641,In_1630,In_2171);
or U642 (N_642,In_382,In_699);
xnor U643 (N_643,In_1351,In_1759);
or U644 (N_644,In_1397,In_842);
or U645 (N_645,In_1092,In_913);
xor U646 (N_646,In_244,In_2992);
nor U647 (N_647,In_556,In_2940);
nor U648 (N_648,In_2454,In_2794);
and U649 (N_649,In_786,In_1368);
xor U650 (N_650,In_500,In_2519);
and U651 (N_651,In_1163,In_2414);
xnor U652 (N_652,In_1198,In_653);
xnor U653 (N_653,In_1606,In_1246);
xnor U654 (N_654,In_2170,In_2495);
xor U655 (N_655,In_1070,In_1941);
or U656 (N_656,In_799,In_1508);
xnor U657 (N_657,In_656,In_756);
and U658 (N_658,In_171,In_1573);
nand U659 (N_659,In_451,In_700);
or U660 (N_660,In_2476,In_1292);
or U661 (N_661,In_2224,In_2406);
or U662 (N_662,In_1791,In_1695);
and U663 (N_663,In_1462,In_2425);
nand U664 (N_664,In_2196,In_1621);
or U665 (N_665,In_1458,In_2198);
and U666 (N_666,In_785,In_2004);
xor U667 (N_667,In_595,In_870);
xor U668 (N_668,In_123,In_1389);
nand U669 (N_669,In_1083,In_56);
nand U670 (N_670,In_332,In_951);
nand U671 (N_671,In_1283,In_2201);
nor U672 (N_672,In_2226,In_864);
nand U673 (N_673,In_1426,In_2588);
nand U674 (N_674,In_1723,In_2749);
xor U675 (N_675,In_999,In_2193);
nand U676 (N_676,In_2852,In_2385);
and U677 (N_677,In_1676,In_570);
xor U678 (N_678,In_1982,In_1224);
nor U679 (N_679,In_844,In_2747);
nand U680 (N_680,In_1180,In_2587);
or U681 (N_681,In_2927,In_1144);
or U682 (N_682,In_2699,In_2344);
and U683 (N_683,In_1693,In_2968);
and U684 (N_684,In_1789,In_2122);
and U685 (N_685,In_1904,In_299);
and U686 (N_686,In_689,In_133);
nand U687 (N_687,In_2030,In_179);
nor U688 (N_688,In_304,In_1640);
and U689 (N_689,In_1048,In_2861);
xor U690 (N_690,In_478,In_2266);
nor U691 (N_691,In_1263,In_917);
or U692 (N_692,In_35,In_2798);
and U693 (N_693,In_2616,In_2228);
nand U694 (N_694,In_2884,In_610);
and U695 (N_695,In_32,In_1218);
or U696 (N_696,In_550,In_1313);
nand U697 (N_697,In_2301,In_2828);
xor U698 (N_698,In_774,In_918);
nor U699 (N_699,In_466,In_1591);
xnor U700 (N_700,In_2542,In_2464);
nand U701 (N_701,In_367,In_2537);
nor U702 (N_702,In_2355,In_1951);
and U703 (N_703,In_1660,In_2303);
or U704 (N_704,In_2400,In_1973);
or U705 (N_705,In_791,In_1939);
and U706 (N_706,In_2018,In_1688);
and U707 (N_707,In_415,In_2553);
or U708 (N_708,In_1255,In_141);
nor U709 (N_709,In_68,In_1068);
and U710 (N_710,In_411,In_1273);
nand U711 (N_711,In_372,In_1744);
xor U712 (N_712,In_1160,In_203);
nand U713 (N_713,In_701,In_1129);
xnor U714 (N_714,In_1081,In_984);
nor U715 (N_715,In_1895,In_497);
nor U716 (N_716,In_83,In_1275);
or U717 (N_717,In_2293,In_615);
nor U718 (N_718,In_739,In_1175);
or U719 (N_719,In_1057,In_2619);
and U720 (N_720,In_2428,In_677);
or U721 (N_721,In_666,In_2987);
nand U722 (N_722,In_1353,In_1624);
and U723 (N_723,In_990,In_1776);
nor U724 (N_724,In_2049,In_1022);
nor U725 (N_725,In_185,In_2236);
nand U726 (N_726,In_2267,In_1784);
and U727 (N_727,In_605,In_463);
and U728 (N_728,In_1094,In_2309);
nor U729 (N_729,In_583,In_140);
xor U730 (N_730,In_2725,In_2746);
nand U731 (N_731,In_832,In_2700);
xnor U732 (N_732,In_1312,In_788);
or U733 (N_733,In_2337,In_2416);
nand U734 (N_734,In_2387,In_1864);
and U735 (N_735,In_1376,In_713);
and U736 (N_736,In_538,In_1858);
and U737 (N_737,In_1179,In_1584);
nor U738 (N_738,In_1841,In_685);
nand U739 (N_739,In_2069,In_627);
and U740 (N_740,In_1002,In_704);
or U741 (N_741,In_373,In_962);
xor U742 (N_742,In_1432,In_1298);
or U743 (N_743,In_2788,In_555);
or U744 (N_744,In_1120,In_2458);
and U745 (N_745,In_1663,In_1887);
and U746 (N_746,In_2928,In_681);
or U747 (N_747,In_2926,In_1347);
nor U748 (N_748,In_363,In_695);
and U749 (N_749,In_1431,In_1445);
xnor U750 (N_750,In_1134,In_1424);
and U751 (N_751,In_716,In_2323);
or U752 (N_752,In_1696,In_2139);
or U753 (N_753,In_2890,In_2098);
or U754 (N_754,In_1600,In_2826);
nor U755 (N_755,In_2347,In_0);
and U756 (N_756,In_2536,In_2353);
nand U757 (N_757,In_469,In_892);
xor U758 (N_758,In_1512,In_2417);
and U759 (N_759,In_468,In_138);
xnor U760 (N_760,In_2603,In_905);
nand U761 (N_761,In_979,In_337);
nor U762 (N_762,In_970,In_1133);
or U763 (N_763,In_2218,In_384);
xor U764 (N_764,In_1131,In_2050);
nor U765 (N_765,In_993,In_632);
xor U766 (N_766,In_2134,In_81);
and U767 (N_767,In_2703,In_174);
or U768 (N_768,In_2556,In_1675);
or U769 (N_769,In_2668,In_114);
nand U770 (N_770,In_2367,In_1441);
and U771 (N_771,In_305,In_742);
nand U772 (N_772,In_2829,In_5);
and U773 (N_773,In_2985,In_2876);
and U774 (N_774,In_1638,In_529);
nand U775 (N_775,In_513,In_1838);
nand U776 (N_776,In_1964,In_1778);
nand U777 (N_777,In_1454,In_2854);
xnor U778 (N_778,In_2210,In_1149);
nand U779 (N_779,In_1734,In_1334);
and U780 (N_780,In_1979,In_718);
and U781 (N_781,In_1634,In_1824);
and U782 (N_782,In_907,In_154);
nand U783 (N_783,In_1510,In_1933);
or U784 (N_784,In_1686,In_2611);
nor U785 (N_785,In_1493,In_2477);
or U786 (N_786,In_508,In_2154);
nor U787 (N_787,In_1544,In_1039);
nor U788 (N_788,In_1321,In_1465);
nor U789 (N_789,In_2221,In_923);
nor U790 (N_790,In_2820,In_1231);
or U791 (N_791,In_1578,In_564);
nor U792 (N_792,In_1586,In_1988);
and U793 (N_793,In_2567,In_2520);
or U794 (N_794,In_572,In_392);
or U795 (N_795,In_2442,In_2233);
and U796 (N_796,In_387,In_1736);
or U797 (N_797,In_2066,In_1812);
nand U798 (N_798,In_2222,In_1146);
xnor U799 (N_799,In_2261,In_2682);
and U800 (N_800,In_687,In_1581);
nor U801 (N_801,In_397,In_2186);
nor U802 (N_802,In_1795,In_347);
nor U803 (N_803,In_2577,In_2505);
xnor U804 (N_804,In_2325,In_1877);
nand U805 (N_805,In_1589,In_2319);
xor U806 (N_806,In_784,In_1735);
nor U807 (N_807,In_890,In_2095);
or U808 (N_808,In_1576,In_1223);
nor U809 (N_809,In_1711,In_2117);
nor U810 (N_810,In_2265,In_1189);
nand U811 (N_811,In_2659,In_2586);
and U812 (N_812,In_2754,In_2966);
nor U813 (N_813,In_727,In_2605);
or U814 (N_814,In_2925,In_1782);
nand U815 (N_815,In_539,In_839);
nor U816 (N_816,In_2135,In_1301);
nand U817 (N_817,In_853,In_1651);
and U818 (N_818,In_1539,In_493);
nand U819 (N_819,In_1570,In_973);
nor U820 (N_820,In_294,In_456);
and U821 (N_821,In_509,In_2459);
nor U822 (N_822,In_2870,In_1752);
or U823 (N_823,In_464,In_400);
or U824 (N_824,In_754,In_854);
xnor U825 (N_825,In_645,In_708);
nand U826 (N_826,In_1439,In_2688);
nand U827 (N_827,In_1857,In_588);
xnor U828 (N_828,In_1239,In_249);
xnor U829 (N_829,In_1339,In_2937);
nand U830 (N_830,In_2033,In_2227);
xnor U831 (N_831,In_2643,In_1005);
nor U832 (N_832,In_172,In_2770);
and U833 (N_833,In_2461,In_1254);
xor U834 (N_834,In_698,In_1338);
or U835 (N_835,In_919,In_533);
nand U836 (N_836,In_2314,In_242);
xor U837 (N_837,In_2584,In_2380);
nand U838 (N_838,In_74,In_1907);
nor U839 (N_839,In_2597,In_2234);
and U840 (N_840,In_75,In_1972);
or U841 (N_841,In_1618,In_1677);
nor U842 (N_842,In_996,In_1429);
and U843 (N_843,In_1142,In_1905);
nand U844 (N_844,In_1101,In_1797);
or U845 (N_845,In_852,In_1482);
nor U846 (N_846,In_1617,In_735);
nand U847 (N_847,In_2031,In_1059);
and U848 (N_848,In_2270,In_2092);
xnor U849 (N_849,In_106,In_2318);
xnor U850 (N_850,In_2705,In_421);
nand U851 (N_851,In_1463,In_767);
and U852 (N_852,In_1102,In_2728);
nand U853 (N_853,In_2887,In_279);
or U854 (N_854,In_2808,In_935);
xnor U855 (N_855,In_1377,In_2894);
nor U856 (N_856,In_924,In_47);
nand U857 (N_857,In_2382,In_481);
xor U858 (N_858,In_120,In_449);
nor U859 (N_859,In_2832,In_2762);
or U860 (N_860,In_288,In_314);
xnor U861 (N_861,In_1614,In_741);
nor U862 (N_862,In_518,In_568);
nand U863 (N_863,In_944,In_1234);
and U864 (N_864,In_1563,In_2895);
xor U865 (N_865,In_2058,In_2767);
or U866 (N_866,In_2924,In_1769);
xnor U867 (N_867,In_2691,In_715);
or U868 (N_868,In_664,In_1535);
xor U869 (N_869,In_2635,In_1703);
or U870 (N_870,In_2358,In_2671);
nor U871 (N_871,In_1867,In_1863);
xnor U872 (N_872,In_2159,In_2908);
and U873 (N_873,In_780,In_2456);
nor U874 (N_874,In_2451,In_1418);
and U875 (N_875,In_1823,In_1790);
nand U876 (N_876,In_1097,In_657);
xor U877 (N_877,In_2521,In_948);
or U878 (N_878,In_217,In_309);
xor U879 (N_879,In_6,In_1221);
and U880 (N_880,In_2704,In_2131);
and U881 (N_881,In_1678,In_1966);
nand U882 (N_882,In_985,In_969);
and U883 (N_883,In_1119,In_1564);
and U884 (N_884,In_2424,In_798);
and U885 (N_885,In_178,In_1157);
or U886 (N_886,In_808,In_379);
and U887 (N_887,In_1361,In_2835);
nor U888 (N_888,In_412,In_2702);
xnor U889 (N_889,In_934,In_2516);
nand U890 (N_890,In_2029,In_2598);
and U891 (N_891,In_1443,In_2949);
and U892 (N_892,In_1528,In_2846);
nand U893 (N_893,In_2116,In_1932);
and U894 (N_894,In_1164,In_1991);
or U895 (N_895,In_611,In_2552);
and U896 (N_896,In_1998,In_822);
or U897 (N_897,In_2294,In_1271);
or U898 (N_898,In_1124,In_1473);
and U899 (N_899,In_165,In_537);
and U900 (N_900,In_2733,In_1464);
xor U901 (N_901,In_1832,In_662);
nand U902 (N_902,In_2990,In_1176);
nor U903 (N_903,In_448,In_576);
nor U904 (N_904,In_2051,In_2957);
and U905 (N_905,In_1879,In_2713);
nor U906 (N_906,In_1659,In_1763);
and U907 (N_907,In_247,In_1728);
nand U908 (N_908,In_544,In_2947);
nand U909 (N_909,In_2207,In_2274);
xnor U910 (N_910,In_2237,In_589);
nand U911 (N_911,In_1945,In_686);
xnor U912 (N_912,In_730,In_932);
nor U913 (N_913,In_1831,In_2290);
nor U914 (N_914,In_959,In_1738);
nor U915 (N_915,In_1854,In_1771);
nand U916 (N_916,In_64,In_2167);
and U917 (N_917,In_2112,In_1781);
xor U918 (N_918,In_649,In_442);
and U919 (N_919,In_1513,In_661);
nand U920 (N_920,In_976,In_2484);
and U921 (N_921,In_1206,In_342);
or U922 (N_922,In_2450,In_227);
nand U923 (N_923,In_802,In_2636);
nand U924 (N_924,In_966,In_2496);
or U925 (N_925,In_875,In_1777);
nor U926 (N_926,In_553,In_2559);
nor U927 (N_927,In_712,In_2297);
and U928 (N_928,In_2730,In_2142);
xnor U929 (N_929,In_1610,In_2110);
nand U930 (N_930,In_673,In_1291);
and U931 (N_931,In_1404,In_2731);
and U932 (N_932,In_1919,In_573);
or U933 (N_933,In_2534,In_370);
nor U934 (N_934,In_562,In_116);
and U935 (N_935,In_307,In_2343);
nand U936 (N_936,In_2581,In_2726);
or U937 (N_937,In_801,In_603);
nor U938 (N_938,In_2275,In_1522);
nor U939 (N_939,In_2429,In_2091);
nand U940 (N_940,In_2562,In_2599);
and U941 (N_941,In_1420,In_490);
or U942 (N_942,In_1402,In_903);
xnor U943 (N_943,In_2453,In_2862);
nor U944 (N_944,In_1780,In_1319);
nor U945 (N_945,In_62,In_1949);
nand U946 (N_946,In_1087,In_1475);
or U947 (N_947,In_2812,In_2527);
nor U948 (N_948,In_2020,In_26);
and U949 (N_949,In_135,In_2864);
and U950 (N_950,In_1018,In_900);
nor U951 (N_951,In_443,In_2650);
and U952 (N_952,In_2200,In_1718);
or U953 (N_953,In_1654,In_2896);
nor U954 (N_954,In_1452,In_2345);
and U955 (N_955,In_205,In_1800);
or U956 (N_956,In_1495,In_404);
nand U957 (N_957,In_872,In_978);
xnor U958 (N_958,In_797,In_1337);
or U959 (N_959,In_2329,In_869);
or U960 (N_960,In_1560,In_2695);
nor U961 (N_961,In_66,In_2640);
or U962 (N_962,In_2612,In_2881);
nand U963 (N_963,In_2042,In_1944);
xnor U964 (N_964,In_1927,In_128);
xnor U965 (N_965,In_335,In_177);
nor U966 (N_966,In_1028,In_1725);
and U967 (N_967,In_1316,In_1847);
xor U968 (N_968,In_2615,In_1814);
xor U969 (N_969,In_818,In_2639);
and U970 (N_970,In_2677,In_956);
nor U971 (N_971,In_2412,In_1685);
or U972 (N_972,In_211,In_12);
or U973 (N_973,In_1492,In_2015);
xnor U974 (N_974,In_1855,In_2500);
nand U975 (N_975,In_1661,In_597);
xor U976 (N_976,In_1296,In_1592);
nor U977 (N_977,In_1158,In_2172);
xnor U978 (N_978,In_2289,In_721);
xor U979 (N_979,In_510,In_1479);
nor U980 (N_980,In_2962,In_2973);
nor U981 (N_981,In_278,In_1616);
nand U982 (N_982,In_2080,In_440);
nor U983 (N_983,In_1060,In_2506);
or U984 (N_984,In_2336,In_2589);
nand U985 (N_985,In_1154,In_927);
nand U986 (N_986,In_1213,In_2889);
xnor U987 (N_987,In_902,In_2868);
xor U988 (N_988,In_1813,In_1821);
or U989 (N_989,In_273,In_2246);
and U990 (N_990,In_1436,In_991);
nand U991 (N_991,In_1029,In_34);
xnor U992 (N_992,In_1530,In_395);
or U993 (N_993,In_2602,In_358);
xor U994 (N_994,In_2359,In_196);
and U995 (N_995,In_943,In_111);
xnor U996 (N_996,In_2108,In_1195);
nor U997 (N_997,In_1041,In_1869);
or U998 (N_998,In_1937,In_1417);
xnor U999 (N_999,In_2235,In_1942);
or U1000 (N_1000,In_750,In_233);
nand U1001 (N_1001,In_2084,In_1975);
and U1002 (N_1002,In_1534,In_2361);
or U1003 (N_1003,In_324,In_848);
xnor U1004 (N_1004,In_1568,In_922);
or U1005 (N_1005,In_740,In_2494);
nand U1006 (N_1006,In_640,In_1726);
nand U1007 (N_1007,In_1182,In_1125);
nand U1008 (N_1008,In_591,In_820);
xnor U1009 (N_1009,In_1708,In_2755);
nand U1010 (N_1010,In_1197,In_31);
nor U1011 (N_1011,In_1844,In_2168);
nor U1012 (N_1012,In_1909,In_574);
or U1013 (N_1013,In_1011,In_1405);
and U1014 (N_1014,In_2161,In_1840);
xor U1015 (N_1015,In_2720,In_747);
or U1016 (N_1016,In_97,In_1976);
nand U1017 (N_1017,In_431,In_1320);
or U1018 (N_1018,In_2203,In_1989);
xnor U1019 (N_1019,In_660,In_671);
and U1020 (N_1020,In_759,In_644);
nand U1021 (N_1021,In_168,In_2853);
or U1022 (N_1022,In_1762,In_1408);
nand U1023 (N_1023,In_2538,In_2781);
nor U1024 (N_1024,In_327,In_2833);
xnor U1025 (N_1025,In_1767,In_2162);
or U1026 (N_1026,In_1702,In_472);
nor U1027 (N_1027,In_1963,In_1827);
and U1028 (N_1028,In_39,In_2952);
nand U1029 (N_1029,In_1562,In_2891);
nand U1030 (N_1030,In_2216,In_175);
nand U1031 (N_1031,In_1008,In_719);
nand U1032 (N_1032,In_432,In_703);
nor U1033 (N_1033,In_2766,In_2583);
xnor U1034 (N_1034,In_2811,In_915);
and U1035 (N_1035,In_909,In_2608);
xnor U1036 (N_1036,In_528,In_855);
nand U1037 (N_1037,In_1227,In_1649);
nand U1038 (N_1038,In_2764,In_1865);
and U1039 (N_1039,In_2948,In_831);
and U1040 (N_1040,In_341,In_127);
nand U1041 (N_1041,In_339,In_815);
and U1042 (N_1042,In_79,In_1994);
xor U1043 (N_1043,In_631,In_2163);
nand U1044 (N_1044,In_1456,In_1332);
nand U1045 (N_1045,In_42,In_2165);
nor U1046 (N_1046,In_1318,In_2727);
nand U1047 (N_1047,In_804,In_1409);
nand U1048 (N_1048,In_1369,In_2564);
and U1049 (N_1049,In_1903,In_2368);
and U1050 (N_1050,In_1435,In_2814);
nand U1051 (N_1051,In_1370,In_29);
nand U1052 (N_1052,In_569,In_361);
nand U1053 (N_1053,In_2003,In_1514);
nor U1054 (N_1054,In_1536,In_197);
or U1055 (N_1055,In_2681,In_2918);
and U1056 (N_1056,In_2350,In_2721);
xnor U1057 (N_1057,In_2499,In_482);
or U1058 (N_1058,In_1551,In_2683);
nand U1059 (N_1059,In_2917,In_863);
nor U1060 (N_1060,In_37,In_920);
and U1061 (N_1061,In_682,In_1135);
xor U1062 (N_1062,In_926,In_2181);
and U1063 (N_1063,In_2238,In_424);
nor U1064 (N_1064,In_2503,In_584);
xnor U1065 (N_1065,In_1756,In_1934);
nand U1066 (N_1066,In_1714,In_86);
or U1067 (N_1067,In_789,In_515);
or U1068 (N_1068,In_1042,In_1181);
nor U1069 (N_1069,In_2150,In_2381);
nand U1070 (N_1070,In_904,In_2548);
nor U1071 (N_1071,In_2960,In_1306);
xor U1072 (N_1072,In_1550,In_2574);
and U1073 (N_1073,In_806,In_2834);
xnor U1074 (N_1074,In_2760,In_2027);
or U1075 (N_1075,In_1826,In_2528);
or U1076 (N_1076,In_1056,In_980);
nand U1077 (N_1077,In_889,In_199);
nand U1078 (N_1078,In_1666,In_1707);
nand U1079 (N_1079,In_2357,In_1722);
xnor U1080 (N_1080,In_540,In_2396);
and U1081 (N_1081,In_1930,In_812);
and U1082 (N_1082,In_668,In_1385);
or U1083 (N_1083,In_1820,In_2244);
and U1084 (N_1084,In_887,In_504);
nor U1085 (N_1085,In_967,In_1467);
and U1086 (N_1086,In_287,In_577);
or U1087 (N_1087,In_2875,In_1801);
or U1088 (N_1088,In_910,In_218);
nand U1089 (N_1089,In_2148,In_159);
nor U1090 (N_1090,In_1317,In_2497);
nand U1091 (N_1091,In_2735,In_519);
xor U1092 (N_1092,In_637,In_263);
xor U1093 (N_1093,In_738,In_182);
nand U1094 (N_1094,In_1038,In_2468);
nor U1095 (N_1095,In_2555,In_2286);
or U1096 (N_1096,In_898,In_9);
nand U1097 (N_1097,In_2631,In_1697);
nor U1098 (N_1098,In_2273,In_1766);
nand U1099 (N_1099,In_1807,In_878);
xor U1100 (N_1100,In_1019,In_2972);
or U1101 (N_1101,In_2410,In_1153);
nand U1102 (N_1102,In_406,In_1069);
or U1103 (N_1103,In_1106,In_2328);
and U1104 (N_1104,In_2245,In_2614);
xnor U1105 (N_1105,In_734,In_638);
xor U1106 (N_1106,In_107,In_1323);
nand U1107 (N_1107,In_2435,In_1959);
or U1108 (N_1108,In_2209,In_643);
nand U1109 (N_1109,In_2722,In_381);
or U1110 (N_1110,In_2026,In_2083);
nor U1111 (N_1111,In_2886,In_2609);
nor U1112 (N_1112,In_1683,In_176);
or U1113 (N_1113,In_2472,In_873);
nand U1114 (N_1114,In_2169,In_1295);
and U1115 (N_1115,In_1114,In_408);
and U1116 (N_1116,In_1872,In_2645);
xor U1117 (N_1117,In_50,In_1034);
xor U1118 (N_1118,In_2388,In_2800);
or U1119 (N_1119,In_487,In_1387);
nor U1120 (N_1120,In_2674,In_2253);
xor U1121 (N_1121,In_680,In_2211);
nor U1122 (N_1122,In_2625,In_246);
or U1123 (N_1123,In_2929,In_95);
or U1124 (N_1124,In_1908,In_2272);
and U1125 (N_1125,In_1746,In_988);
and U1126 (N_1126,In_1995,In_1608);
xor U1127 (N_1127,In_2709,In_2087);
nand U1128 (N_1128,In_61,In_879);
nor U1129 (N_1129,In_2634,In_803);
nand U1130 (N_1130,In_2,In_1136);
nor U1131 (N_1131,In_1917,In_1527);
nor U1132 (N_1132,In_2436,In_63);
or U1133 (N_1133,In_2028,In_426);
nor U1134 (N_1134,In_1166,In_743);
or U1135 (N_1135,In_758,In_604);
xor U1136 (N_1136,In_208,In_2473);
xnor U1137 (N_1137,In_787,In_1468);
xnor U1138 (N_1138,In_1545,In_1061);
xor U1139 (N_1139,In_87,In_783);
and U1140 (N_1140,In_99,In_1010);
or U1141 (N_1141,In_952,In_322);
or U1142 (N_1142,In_1108,In_401);
and U1143 (N_1143,In_554,In_1309);
xnor U1144 (N_1144,In_1911,In_2763);
nor U1145 (N_1145,In_2157,In_1250);
and U1146 (N_1146,In_1201,In_2514);
or U1147 (N_1147,In_1987,In_2898);
or U1148 (N_1148,In_2268,In_697);
and U1149 (N_1149,In_126,In_380);
nor U1150 (N_1150,In_319,In_1349);
nor U1151 (N_1151,In_2212,In_2471);
and U1152 (N_1152,In_2376,In_326);
nor U1153 (N_1153,In_2063,In_2590);
and U1154 (N_1154,In_901,In_2153);
and U1155 (N_1155,In_2620,In_899);
or U1156 (N_1156,In_53,In_1466);
nand U1157 (N_1157,In_503,In_2573);
nand U1158 (N_1158,In_502,In_772);
and U1159 (N_1159,In_2311,In_1565);
and U1160 (N_1160,In_253,In_2231);
nor U1161 (N_1161,In_21,In_2302);
or U1162 (N_1162,In_1974,In_1652);
xnor U1163 (N_1163,In_1371,In_2593);
or U1164 (N_1164,In_1809,In_2250);
or U1165 (N_1165,In_809,In_2769);
xor U1166 (N_1166,In_229,In_1233);
nand U1167 (N_1167,In_2911,In_1552);
nor U1168 (N_1168,In_2629,In_2626);
nor U1169 (N_1169,In_630,In_2415);
nand U1170 (N_1170,In_1980,In_765);
nor U1171 (N_1171,In_1450,In_1774);
or U1172 (N_1172,In_1561,In_3);
nand U1173 (N_1173,In_118,In_1594);
xnor U1174 (N_1174,In_1669,In_916);
nand U1175 (N_1175,In_2283,In_2269);
and U1176 (N_1176,In_2600,In_1145);
xnor U1177 (N_1177,In_2802,In_422);
nor U1178 (N_1178,In_2102,In_2078);
or U1179 (N_1179,In_2915,In_2621);
and U1180 (N_1180,In_2950,In_2965);
or U1181 (N_1181,In_102,In_303);
xor U1182 (N_1182,In_1178,In_228);
or U1183 (N_1183,In_2120,In_2797);
nand U1184 (N_1184,In_1689,In_2554);
and U1185 (N_1185,In_2923,In_1611);
xnor U1186 (N_1186,In_2882,In_44);
nand U1187 (N_1187,In_1601,In_963);
nor U1188 (N_1188,In_1278,In_2855);
and U1189 (N_1189,In_2107,In_1731);
or U1190 (N_1190,In_477,In_113);
or U1191 (N_1191,In_796,In_1352);
nor U1192 (N_1192,In_2082,In_1913);
nand U1193 (N_1193,In_433,In_2738);
or U1194 (N_1194,In_151,In_771);
nor U1195 (N_1195,In_1362,In_1471);
nand U1196 (N_1196,In_2096,In_136);
or U1197 (N_1197,In_1249,In_1392);
xor U1198 (N_1198,In_2558,In_2331);
nor U1199 (N_1199,In_1650,In_975);
or U1200 (N_1200,N_217,N_648);
nor U1201 (N_1201,N_122,In_1615);
nand U1202 (N_1202,In_1331,N_457);
nor U1203 (N_1203,In_705,In_1737);
xnor U1204 (N_1204,N_975,In_2321);
and U1205 (N_1205,In_2523,N_596);
xor U1206 (N_1206,In_1572,In_306);
or U1207 (N_1207,N_1110,In_1031);
nand U1208 (N_1208,N_759,N_821);
nor U1209 (N_1209,In_1523,N_281);
xnor U1210 (N_1210,N_338,N_516);
or U1211 (N_1211,N_904,N_198);
nand U1212 (N_1212,N_674,In_2975);
nand U1213 (N_1213,In_2447,N_827);
nand U1214 (N_1214,N_453,N_951);
or U1215 (N_1215,N_91,N_1014);
and U1216 (N_1216,N_195,N_1061);
or U1217 (N_1217,N_1147,N_780);
or U1218 (N_1218,In_2708,N_947);
and U1219 (N_1219,In_1082,In_536);
nand U1220 (N_1220,N_162,In_447);
and U1221 (N_1221,In_1538,In_810);
and U1222 (N_1222,In_1509,N_844);
nand U1223 (N_1223,N_983,N_929);
nand U1224 (N_1224,In_276,N_540);
and U1225 (N_1225,N_661,In_403);
xor U1226 (N_1226,N_801,In_78);
nand U1227 (N_1227,N_660,N_455);
nand U1228 (N_1228,N_541,In_2466);
nor U1229 (N_1229,N_1097,N_1131);
or U1230 (N_1230,In_110,N_78);
nand U1231 (N_1231,In_1130,In_1049);
or U1232 (N_1232,N_477,N_118);
and U1233 (N_1233,In_2394,N_467);
nor U1234 (N_1234,N_852,N_279);
nand U1235 (N_1235,In_2315,N_1134);
nand U1236 (N_1236,In_88,In_2867);
nand U1237 (N_1237,N_546,N_610);
nand U1238 (N_1238,N_111,N_501);
nand U1239 (N_1239,N_5,In_169);
or U1240 (N_1240,N_524,N_518);
xnor U1241 (N_1241,N_845,N_726);
nor U1242 (N_1242,N_26,N_617);
and U1243 (N_1243,In_265,N_1133);
nor U1244 (N_1244,N_377,N_642);
nor U1245 (N_1245,In_2578,N_877);
nor U1246 (N_1246,N_421,N_689);
nor U1247 (N_1247,In_1383,N_62);
nand U1248 (N_1248,N_38,N_312);
and U1249 (N_1249,In_1607,N_552);
nand U1250 (N_1250,N_720,In_1846);
or U1251 (N_1251,N_743,In_1794);
xnor U1252 (N_1252,N_741,N_861);
or U1253 (N_1253,N_503,N_1064);
and U1254 (N_1254,N_156,N_1186);
xor U1255 (N_1255,In_282,N_795);
nand U1256 (N_1256,N_739,N_1025);
and U1257 (N_1257,N_749,In_2090);
nand U1258 (N_1258,N_276,In_410);
or U1259 (N_1259,N_487,In_726);
nor U1260 (N_1260,N_45,N_1066);
xnor U1261 (N_1261,N_478,N_371);
and U1262 (N_1262,N_245,In_646);
nor U1263 (N_1263,N_108,In_2363);
xnor U1264 (N_1264,N_102,N_637);
nand U1265 (N_1265,In_2252,N_1105);
nand U1266 (N_1266,N_623,N_635);
or U1267 (N_1267,In_2104,N_1163);
and U1268 (N_1268,N_482,N_737);
nor U1269 (N_1269,N_578,N_1160);
nor U1270 (N_1270,N_1137,N_125);
nand U1271 (N_1271,N_410,N_711);
nor U1272 (N_1272,N_681,N_567);
or U1273 (N_1273,N_978,In_2123);
nor U1274 (N_1274,N_90,N_1135);
nand U1275 (N_1275,N_562,In_1020);
xnor U1276 (N_1276,N_563,In_600);
nor U1277 (N_1277,N_130,In_377);
nor U1278 (N_1278,N_543,N_317);
and U1279 (N_1279,N_892,N_1195);
nand U1280 (N_1280,In_1294,N_753);
or U1281 (N_1281,N_1121,N_79);
xnor U1282 (N_1282,N_598,In_1956);
nor U1283 (N_1283,N_764,N_906);
nor U1284 (N_1284,N_183,N_778);
and U1285 (N_1285,N_843,N_1079);
nand U1286 (N_1286,In_2048,N_422);
xnor U1287 (N_1287,In_1899,In_1603);
nor U1288 (N_1288,N_1102,N_1113);
nor U1289 (N_1289,In_2009,N_744);
nand U1290 (N_1290,In_982,In_1400);
nand U1291 (N_1291,N_17,N_806);
nand U1292 (N_1292,In_17,N_256);
nand U1293 (N_1293,In_210,N_246);
xnor U1294 (N_1294,N_858,N_776);
or U1295 (N_1295,N_902,N_556);
or U1296 (N_1296,N_592,N_51);
and U1297 (N_1297,N_220,N_257);
and U1298 (N_1298,N_577,N_134);
nor U1299 (N_1299,In_1852,In_938);
or U1300 (N_1300,In_1095,N_885);
xor U1301 (N_1301,In_1013,N_177);
and U1302 (N_1302,N_29,In_1322);
and U1303 (N_1303,N_564,N_504);
nand U1304 (N_1304,In_209,In_1105);
xnor U1305 (N_1305,N_926,N_31);
nand U1306 (N_1306,N_211,N_119);
xnor U1307 (N_1307,N_890,N_553);
nor U1308 (N_1308,N_182,N_944);
nand U1309 (N_1309,In_2276,N_83);
xor U1310 (N_1310,In_1505,N_1187);
and U1311 (N_1311,N_344,N_1086);
nor U1312 (N_1312,In_937,In_1644);
and U1313 (N_1313,N_494,In_813);
nor U1314 (N_1314,In_1237,In_1519);
xor U1315 (N_1315,N_520,N_908);
nor U1316 (N_1316,N_1067,In_2264);
xor U1317 (N_1317,N_638,N_862);
nor U1318 (N_1318,N_247,N_917);
or U1319 (N_1319,N_462,In_1531);
and U1320 (N_1320,N_857,N_591);
and U1321 (N_1321,N_1142,N_872);
nor U1322 (N_1322,N_1056,In_1422);
and U1323 (N_1323,N_252,N_1048);
nand U1324 (N_1324,In_274,In_2816);
xor U1325 (N_1325,N_653,N_842);
nor U1326 (N_1326,N_1174,N_417);
nand U1327 (N_1327,N_172,N_1164);
and U1328 (N_1328,In_1674,N_527);
or U1329 (N_1329,N_1183,N_408);
xnor U1330 (N_1330,In_2177,N_777);
nor U1331 (N_1331,In_692,N_302);
or U1332 (N_1332,In_2916,N_701);
xor U1333 (N_1333,In_1090,N_530);
xor U1334 (N_1334,N_785,In_444);
nor U1335 (N_1335,In_436,In_250);
and U1336 (N_1336,N_1181,In_277);
xnor U1337 (N_1337,N_307,N_675);
nor U1338 (N_1338,N_173,In_1894);
or U1339 (N_1339,In_1727,N_479);
xnor U1340 (N_1340,N_85,In_1078);
xnor U1341 (N_1341,N_242,N_870);
or U1342 (N_1342,In_833,In_1667);
or U1343 (N_1343,N_52,N_1150);
or U1344 (N_1344,In_80,In_148);
xnor U1345 (N_1345,In_2342,In_679);
xor U1346 (N_1346,In_1673,N_115);
xor U1347 (N_1347,In_1459,N_565);
or U1348 (N_1348,N_355,N_706);
or U1349 (N_1349,In_1192,N_448);
and U1350 (N_1350,N_224,N_407);
xor U1351 (N_1351,N_155,N_1176);
nand U1352 (N_1352,N_499,N_1023);
xnor U1353 (N_1353,In_2136,N_221);
or U1354 (N_1354,N_533,In_413);
xor U1355 (N_1355,N_960,In_121);
xnor U1356 (N_1356,In_2242,N_1009);
or U1357 (N_1357,N_698,In_675);
and U1358 (N_1358,N_121,N_71);
and U1359 (N_1359,In_1620,N_1199);
or U1360 (N_1360,In_2362,In_2869);
and U1361 (N_1361,In_1983,N_879);
or U1362 (N_1362,N_77,N_425);
and U1363 (N_1363,N_1035,N_1065);
xnor U1364 (N_1364,N_234,N_47);
nand U1365 (N_1365,N_92,In_257);
and U1366 (N_1366,N_1045,N_1098);
and U1367 (N_1367,N_846,In_2434);
or U1368 (N_1368,N_684,N_656);
and U1369 (N_1369,N_424,N_914);
xor U1370 (N_1370,In_2285,In_911);
nor U1371 (N_1371,In_998,N_296);
and U1372 (N_1372,N_1044,N_320);
xnor U1373 (N_1373,N_659,N_995);
and U1374 (N_1374,N_668,N_672);
or U1375 (N_1375,In_2255,N_1083);
or U1376 (N_1376,N_537,N_70);
nand U1377 (N_1377,In_2034,N_1015);
xnor U1378 (N_1378,N_814,In_2633);
nand U1379 (N_1379,In_105,In_2653);
nor U1380 (N_1380,N_412,N_287);
or U1381 (N_1381,N_36,N_1177);
nand U1382 (N_1382,In_2395,N_943);
nor U1383 (N_1383,In_2675,In_2073);
nand U1384 (N_1384,N_771,N_465);
nor U1385 (N_1385,In_248,In_2774);
xnor U1386 (N_1386,N_1159,N_998);
or U1387 (N_1387,N_64,N_900);
xor U1388 (N_1388,N_856,In_2407);
nand U1389 (N_1389,N_1081,N_416);
nand U1390 (N_1390,N_517,In_1293);
and U1391 (N_1391,N_394,N_688);
xor U1392 (N_1392,N_306,N_523);
nand U1393 (N_1393,N_971,In_543);
xnor U1394 (N_1394,N_210,N_61);
xor U1395 (N_1395,N_324,N_586);
nor U1396 (N_1396,N_282,In_2008);
and U1397 (N_1397,N_717,In_1747);
nand U1398 (N_1398,N_889,In_2465);
nand U1399 (N_1399,N_869,N_191);
or U1400 (N_1400,N_295,N_631);
nor U1401 (N_1401,N_807,N_670);
xnor U1402 (N_1402,In_2288,In_2263);
and U1403 (N_1403,N_142,N_1027);
nor U1404 (N_1404,In_1374,In_620);
and U1405 (N_1405,N_473,N_486);
xor U1406 (N_1406,N_969,N_59);
or U1407 (N_1407,In_376,In_571);
xnor U1408 (N_1408,In_2501,N_243);
or U1409 (N_1409,In_290,N_101);
nand U1410 (N_1410,N_539,In_2440);
nand U1411 (N_1411,In_225,N_16);
xnor U1412 (N_1412,N_587,In_1525);
and U1413 (N_1413,N_214,N_1034);
and U1414 (N_1414,N_934,In_1668);
xnor U1415 (N_1415,In_2411,In_131);
nor U1416 (N_1416,In_1521,N_152);
xnor U1417 (N_1417,In_1842,N_981);
or U1418 (N_1418,N_963,N_285);
nand U1419 (N_1419,In_2280,In_2103);
nand U1420 (N_1420,In_2874,N_464);
and U1421 (N_1421,N_141,N_230);
and U1422 (N_1422,In_2851,In_1440);
nor U1423 (N_1423,In_2340,In_859);
nor U1424 (N_1424,N_216,N_608);
nor U1425 (N_1425,N_622,N_54);
nand U1426 (N_1426,N_614,In_2892);
nand U1427 (N_1427,N_131,N_447);
nand U1428 (N_1428,N_472,N_415);
nor U1429 (N_1429,N_1037,N_992);
and U1430 (N_1430,N_912,N_611);
nor U1431 (N_1431,N_525,N_269);
nand U1432 (N_1432,In_359,N_1170);
xor U1433 (N_1433,In_1425,N_233);
xnor U1434 (N_1434,N_1109,N_167);
xor U1435 (N_1435,N_1193,N_14);
nor U1436 (N_1436,In_868,N_350);
nor U1437 (N_1437,In_2239,N_788);
nor U1438 (N_1438,N_933,In_316);
nand U1439 (N_1439,N_342,N_909);
xor U1440 (N_1440,N_1114,In_691);
nor U1441 (N_1441,N_962,N_755);
nand U1442 (N_1442,N_313,N_199);
or U1443 (N_1443,In_549,In_1773);
xnor U1444 (N_1444,In_437,N_431);
and U1445 (N_1445,N_942,N_124);
xnor U1446 (N_1446,In_2320,N_1082);
nand U1447 (N_1447,N_1101,N_208);
nand U1448 (N_1448,In_1948,In_2809);
and U1449 (N_1449,N_1008,N_748);
nand U1450 (N_1450,In_1511,In_331);
nor U1451 (N_1451,In_1645,N_87);
xor U1452 (N_1452,N_50,N_826);
and U1453 (N_1453,N_345,N_498);
nor U1454 (N_1454,N_323,N_791);
nand U1455 (N_1455,N_171,In_1151);
xnor U1456 (N_1456,In_2651,In_1073);
nand U1457 (N_1457,N_278,N_789);
nor U1458 (N_1458,In_551,N_497);
or U1459 (N_1459,In_1325,In_2964);
nor U1460 (N_1460,N_116,In_2271);
or U1461 (N_1461,N_1184,N_288);
and U1462 (N_1462,N_67,N_1020);
xor U1463 (N_1463,In_720,In_2707);
xnor U1464 (N_1464,In_1850,In_1922);
or U1465 (N_1465,N_1012,In_2592);
xnor U1466 (N_1466,N_190,N_333);
xnor U1467 (N_1467,N_314,N_1062);
nor U1468 (N_1468,N_542,In_1455);
nor U1469 (N_1469,In_1713,In_1583);
nor U1470 (N_1470,In_59,N_1072);
nand U1471 (N_1471,N_96,N_72);
and U1472 (N_1472,In_1554,N_28);
nand U1473 (N_1473,In_2094,In_2129);
and U1474 (N_1474,N_207,N_1070);
or U1475 (N_1475,N_831,N_910);
nand U1476 (N_1476,N_328,N_363);
and U1477 (N_1477,In_258,N_531);
or U1478 (N_1478,N_1029,N_174);
or U1479 (N_1479,N_761,N_1146);
nand U1480 (N_1480,N_897,In_491);
xor U1481 (N_1481,N_569,In_1684);
or U1482 (N_1482,N_1161,N_649);
and U1483 (N_1483,N_228,N_10);
xnor U1484 (N_1484,N_106,N_273);
nand U1485 (N_1485,N_700,In_2569);
xor U1486 (N_1486,In_2099,In_1375);
or U1487 (N_1487,In_2585,In_1084);
or U1488 (N_1488,N_946,N_646);
nand U1489 (N_1489,N_959,N_936);
or U1490 (N_1490,In_1006,In_522);
nand U1491 (N_1491,N_918,In_2119);
nand U1492 (N_1492,In_2305,N_1173);
xnor U1493 (N_1493,N_480,In_1516);
xnor U1494 (N_1494,N_80,N_379);
xnor U1495 (N_1495,N_809,N_583);
and U1496 (N_1496,In_150,N_321);
or U1497 (N_1497,In_939,N_213);
xor U1498 (N_1498,In_706,In_2662);
nor U1499 (N_1499,In_707,N_830);
or U1500 (N_1500,N_952,N_794);
or U1501 (N_1501,N_607,N_386);
nand U1502 (N_1502,N_441,In_1898);
and U1503 (N_1503,N_7,In_1506);
nor U1504 (N_1504,N_996,N_766);
or U1505 (N_1505,N_443,N_388);
and U1506 (N_1506,In_1438,N_255);
or U1507 (N_1507,N_270,In_2660);
nor U1508 (N_1508,N_620,N_267);
or U1509 (N_1509,N_24,N_702);
and U1510 (N_1510,In_2277,N_200);
and U1511 (N_1511,N_81,N_817);
nand U1512 (N_1512,N_931,N_1047);
nand U1513 (N_1513,N_341,In_725);
and U1514 (N_1514,N_375,N_429);
xor U1515 (N_1515,In_2693,N_715);
xnor U1516 (N_1516,N_1104,N_718);
and U1517 (N_1517,N_203,N_949);
and U1518 (N_1518,N_522,N_89);
and U1519 (N_1519,In_2622,In_1483);
or U1520 (N_1520,In_1187,In_2570);
or U1521 (N_1521,N_997,In_930);
or U1522 (N_1522,In_192,N_404);
nand U1523 (N_1523,In_1199,N_1084);
or U1524 (N_1524,N_1179,N_948);
nand U1525 (N_1525,N_358,N_148);
nor U1526 (N_1526,In_1657,N_33);
xor U1527 (N_1527,N_471,N_905);
xor U1528 (N_1528,In_1788,N_236);
or U1529 (N_1529,In_103,In_1214);
and U1530 (N_1530,N_239,N_6);
or U1531 (N_1531,N_813,N_489);
nor U1532 (N_1532,N_348,N_250);
nor U1533 (N_1533,In_2878,N_633);
and U1534 (N_1534,N_645,N_1116);
xnor U1535 (N_1535,In_883,N_193);
and U1536 (N_1536,In_1115,N_665);
nand U1537 (N_1537,N_1112,N_571);
and U1538 (N_1538,In_72,N_264);
or U1539 (N_1539,In_166,N_751);
nand U1540 (N_1540,N_9,In_1274);
nor U1541 (N_1541,In_1484,In_2360);
and U1542 (N_1542,N_1182,N_515);
nor U1543 (N_1543,N_1130,In_13);
nand U1544 (N_1544,N_128,In_1072);
or U1545 (N_1545,N_500,N_460);
nand U1546 (N_1546,N_957,N_368);
or U1547 (N_1547,N_402,N_939);
and U1548 (N_1548,N_859,In_1063);
xor U1549 (N_1549,N_169,N_1030);
nor U1550 (N_1550,N_366,N_994);
nor U1551 (N_1551,In_2059,N_1167);
or U1552 (N_1552,N_227,N_298);
or U1553 (N_1553,N_991,In_1261);
and U1554 (N_1554,N_1145,In_2057);
nand U1555 (N_1555,N_627,In_1148);
nor U1556 (N_1556,N_444,In_658);
nand U1557 (N_1557,In_2322,N_812);
nor U1558 (N_1558,N_851,N_164);
or U1559 (N_1559,In_2565,N_837);
nor U1560 (N_1560,N_535,N_356);
and U1561 (N_1561,In_1230,N_37);
and U1562 (N_1562,N_428,N_374);
and U1563 (N_1563,N_625,In_1952);
nor U1564 (N_1564,N_367,N_340);
nor U1565 (N_1565,N_223,N_1124);
nor U1566 (N_1566,N_663,N_937);
or U1567 (N_1567,N_626,In_170);
nand U1568 (N_1568,N_742,N_738);
nor U1569 (N_1569,In_58,In_14);
xnor U1570 (N_1570,N_529,N_1013);
or U1571 (N_1571,N_604,N_463);
and U1572 (N_1572,N_205,In_1266);
and U1573 (N_1573,In_2375,N_265);
and U1574 (N_1574,N_143,N_370);
and U1575 (N_1575,In_684,N_836);
nand U1576 (N_1576,In_2038,N_526);
xnor U1577 (N_1577,N_120,N_1190);
nand U1578 (N_1578,N_397,In_2697);
nand U1579 (N_1579,N_964,N_300);
nor U1580 (N_1580,N_1050,N_1144);
nand U1581 (N_1581,N_1000,N_385);
xor U1582 (N_1582,In_1882,In_48);
nor U1583 (N_1583,N_112,N_630);
and U1584 (N_1584,N_797,N_512);
and U1585 (N_1585,In_134,N_437);
and U1586 (N_1586,N_730,N_414);
or U1587 (N_1587,In_748,N_318);
nor U1588 (N_1588,N_928,N_335);
or U1589 (N_1589,N_1018,In_457);
nor U1590 (N_1590,N_832,N_1007);
xor U1591 (N_1591,In_2729,N_599);
and U1592 (N_1592,N_982,N_1063);
and U1593 (N_1593,N_669,N_584);
nor U1594 (N_1594,N_724,N_362);
xor U1595 (N_1595,N_1068,N_781);
and U1596 (N_1596,N_380,In_2568);
and U1597 (N_1597,In_1938,N_883);
or U1598 (N_1598,In_2475,N_1128);
or U1599 (N_1599,N_707,N_286);
or U1600 (N_1600,N_1055,N_572);
nand U1601 (N_1601,In_1386,N_735);
and U1602 (N_1602,In_1282,N_796);
nand U1603 (N_1603,N_644,N_153);
xor U1604 (N_1604,In_7,N_1122);
nor U1605 (N_1605,In_1380,N_792);
and U1606 (N_1606,In_1874,N_1149);
or U1607 (N_1607,In_1706,N_887);
or U1608 (N_1608,N_882,In_2176);
nor U1609 (N_1609,In_93,In_1026);
nor U1610 (N_1610,N_158,N_574);
nor U1611 (N_1611,In_2199,N_815);
xor U1612 (N_1612,N_808,N_495);
xor U1613 (N_1613,In_2432,In_2483);
or U1614 (N_1614,N_554,N_590);
or U1615 (N_1615,N_432,N_621);
nand U1616 (N_1616,In_2214,N_768);
and U1617 (N_1617,N_1024,N_582);
nor U1618 (N_1618,N_1197,N_202);
nand U1619 (N_1619,N_657,In_1489);
or U1620 (N_1620,N_19,N_439);
xnor U1621 (N_1621,N_206,N_888);
and U1622 (N_1622,In_329,N_197);
nor U1623 (N_1623,N_413,N_722);
and U1624 (N_1624,N_732,In_795);
nor U1625 (N_1625,N_272,N_454);
or U1626 (N_1626,In_2541,N_691);
xnor U1627 (N_1627,N_721,N_1123);
and U1628 (N_1628,N_880,N_218);
and U1629 (N_1629,N_509,N_74);
and U1630 (N_1630,In_1343,In_1876);
or U1631 (N_1631,N_1157,In_2989);
nor U1632 (N_1632,N_919,In_70);
and U1633 (N_1633,In_479,N_828);
xnor U1634 (N_1634,In_2300,N_434);
nor U1635 (N_1635,N_260,N_418);
nor U1636 (N_1636,N_95,N_274);
nor U1637 (N_1637,In_751,N_474);
and U1638 (N_1638,N_513,N_990);
nor U1639 (N_1639,N_597,In_328);
or U1640 (N_1640,N_873,N_907);
or U1641 (N_1641,In_2991,N_56);
nand U1642 (N_1642,N_647,In_108);
nand U1643 (N_1643,In_2370,N_671);
and U1644 (N_1644,N_435,N_1169);
nor U1645 (N_1645,In_1172,N_876);
nand U1646 (N_1646,N_1051,N_1021);
xnor U1647 (N_1647,In_1717,In_28);
or U1648 (N_1648,N_1156,In_2856);
xor U1649 (N_1649,N_27,N_48);
or U1650 (N_1650,In_858,N_557);
or U1651 (N_1651,N_746,N_337);
or U1652 (N_1652,N_259,In_867);
nand U1653 (N_1653,N_506,N_579);
xnor U1654 (N_1654,N_865,N_373);
nand U1655 (N_1655,In_1501,N_15);
or U1656 (N_1656,In_207,N_60);
or U1657 (N_1657,In_2732,In_38);
xor U1658 (N_1658,N_212,N_941);
or U1659 (N_1659,In_2507,In_164);
xor U1660 (N_1660,N_1143,In_2710);
nor U1661 (N_1661,N_787,N_979);
or U1662 (N_1662,N_450,In_1665);
and U1663 (N_1663,In_2897,N_1198);
or U1664 (N_1664,N_798,N_387);
nor U1665 (N_1665,N_168,In_1648);
and U1666 (N_1666,N_58,N_1138);
xnor U1667 (N_1667,N_745,N_1074);
nand U1668 (N_1668,N_528,In_594);
or U1669 (N_1669,In_2958,N_716);
and U1670 (N_1670,N_690,N_894);
or U1671 (N_1671,N_251,N_891);
and U1672 (N_1672,In_2151,N_551);
nand U1673 (N_1673,N_863,In_383);
xnor U1674 (N_1674,N_229,N_1196);
nor U1675 (N_1675,N_989,N_483);
and U1676 (N_1676,In_1655,N_570);
or U1677 (N_1677,In_824,N_209);
nor U1678 (N_1678,In_1985,N_752);
and U1679 (N_1679,In_805,N_987);
or U1680 (N_1680,N_1057,In_1753);
xor U1681 (N_1681,N_927,N_290);
xnor U1682 (N_1682,In_2919,In_1284);
nand U1683 (N_1683,N_18,In_1403);
nand U1684 (N_1684,N_445,In_874);
or U1685 (N_1685,N_634,N_855);
xnor U1686 (N_1686,In_355,In_1912);
nor U1687 (N_1687,In_2041,N_68);
or U1688 (N_1688,In_1434,N_1060);
and U1689 (N_1689,In_223,In_1729);
and U1690 (N_1690,In_461,N_481);
nand U1691 (N_1691,N_588,N_938);
and U1692 (N_1692,N_733,N_322);
or U1693 (N_1693,N_32,N_248);
nor U1694 (N_1694,N_999,In_2544);
xnor U1695 (N_1695,N_560,In_1228);
or U1696 (N_1696,In_1633,N_100);
nand U1697 (N_1697,N_973,In_908);
nand U1698 (N_1698,N_871,N_1185);
nor U1699 (N_1699,N_581,N_452);
nor U1700 (N_1700,N_820,N_176);
xnor U1701 (N_1701,In_280,N_170);
xnor U1702 (N_1702,N_651,In_162);
or U1703 (N_1703,N_349,N_364);
nand U1704 (N_1704,N_816,N_466);
xnor U1705 (N_1705,In_1217,N_580);
or U1706 (N_1706,N_1077,In_1421);
nand U1707 (N_1707,In_2837,N_652);
or U1708 (N_1708,In_1891,In_1211);
nor U1709 (N_1709,N_896,N_961);
and U1710 (N_1710,N_762,In_1892);
xor U1711 (N_1711,In_678,In_1305);
xnor U1712 (N_1712,In_1890,N_284);
xnor U1713 (N_1713,In_968,N_258);
and U1714 (N_1714,N_219,In_1074);
nand U1715 (N_1715,N_369,N_57);
or U1716 (N_1716,In_981,N_3);
or U1717 (N_1717,N_920,N_619);
xor U1718 (N_1718,N_186,N_357);
nor U1719 (N_1719,N_184,N_1091);
nor U1720 (N_1720,In_1739,In_1085);
nand U1721 (N_1721,N_1162,N_521);
xnor U1722 (N_1722,N_723,N_157);
or U1723 (N_1723,N_685,In_2901);
or U1724 (N_1724,N_507,N_756);
nand U1725 (N_1725,In_850,N_811);
nor U1726 (N_1726,N_25,N_1075);
and U1727 (N_1727,N_1125,N_163);
nor U1728 (N_1728,N_825,In_1021);
and U1729 (N_1729,N_1026,N_84);
or U1730 (N_1730,In_1480,N_126);
or U1731 (N_1731,In_1967,In_2765);
nand U1732 (N_1732,N_829,N_1141);
nor U1733 (N_1733,In_1577,In_1486);
and U1734 (N_1734,In_2663,N_1092);
and U1735 (N_1735,N_271,N_53);
nand U1736 (N_1736,N_618,N_316);
nor U1737 (N_1737,N_1006,In_792);
nor U1738 (N_1738,N_823,N_382);
nor U1739 (N_1739,In_2513,N_442);
or U1740 (N_1740,In_2905,N_696);
nor U1741 (N_1741,N_315,N_993);
nand U1742 (N_1742,N_8,N_175);
nand U1743 (N_1743,In_1314,In_1626);
nor U1744 (N_1744,N_1073,N_332);
or U1745 (N_1745,N_329,In_1575);
or U1746 (N_1746,In_19,N_1155);
and U1747 (N_1747,N_146,In_1159);
nand U1748 (N_1748,N_654,In_2202);
and U1749 (N_1749,N_1175,N_866);
nand U1750 (N_1750,N_734,N_1085);
nor U1751 (N_1751,N_107,In_2391);
or U1752 (N_1752,N_758,In_18);
or U1753 (N_1753,N_304,N_400);
nor U1754 (N_1754,In_992,N_226);
xor U1755 (N_1755,N_103,N_679);
nor U1756 (N_1756,In_1310,N_468);
or U1757 (N_1757,N_166,In_2996);
and U1758 (N_1758,In_2409,N_266);
xor U1759 (N_1759,N_409,N_488);
nor U1760 (N_1760,N_144,N_133);
and U1761 (N_1761,In_1540,N_549);
nand U1762 (N_1762,In_1098,N_773);
nor U1763 (N_1763,In_2007,N_46);
or U1764 (N_1764,In_1834,In_2667);
nor U1765 (N_1765,In_1623,N_976);
and U1766 (N_1766,N_1099,In_2408);
nor U1767 (N_1767,N_360,In_648);
xnor U1768 (N_1768,In_1670,In_811);
nor U1769 (N_1769,N_1151,N_782);
and U1770 (N_1770,In_2649,In_2062);
nand U1771 (N_1771,In_987,N_319);
nand U1772 (N_1772,N_1118,N_129);
and U1773 (N_1773,In_2934,N_1090);
nor U1774 (N_1774,N_1129,In_1764);
nor U1775 (N_1775,In_906,In_1524);
and U1776 (N_1776,In_1210,N_1115);
nand U1777 (N_1777,N_215,N_511);
and U1778 (N_1778,N_765,In_2482);
or U1779 (N_1779,N_405,In_624);
or U1780 (N_1780,N_641,In_2045);
nor U1781 (N_1781,N_23,N_151);
or U1782 (N_1782,N_783,N_676);
and U1783 (N_1783,N_705,N_343);
nand U1784 (N_1784,N_268,In_587);
nand U1785 (N_1785,N_1005,N_519);
and U1786 (N_1786,N_616,N_383);
xnor U1787 (N_1787,N_1166,N_673);
nand U1788 (N_1788,N_1094,In_1140);
or U1789 (N_1789,In_1786,In_2806);
or U1790 (N_1790,N_775,N_1001);
and U1791 (N_1791,N_180,In_2111);
xor U1792 (N_1792,N_339,N_712);
and U1793 (N_1793,In_1768,N_82);
and U1794 (N_1794,N_1103,N_336);
and U1795 (N_1795,N_280,N_66);
xnor U1796 (N_1796,N_93,N_1088);
nor U1797 (N_1797,N_779,In_650);
nor U1798 (N_1798,In_2077,N_179);
nand U1799 (N_1799,N_73,N_824);
and U1800 (N_1800,In_1202,N_760);
nor U1801 (N_1801,N_725,In_2986);
or U1802 (N_1802,N_898,N_94);
nand U1803 (N_1803,N_254,N_955);
or U1804 (N_1804,N_548,N_351);
xor U1805 (N_1805,N_678,N_160);
or U1806 (N_1806,N_436,N_984);
nand U1807 (N_1807,N_916,In_2938);
nand U1808 (N_1808,N_461,In_1193);
and U1809 (N_1809,N_42,In_1499);
nor U1810 (N_1810,N_1087,In_2126);
and U1811 (N_1811,In_1802,N_958);
and U1812 (N_1812,N_804,N_568);
nand U1813 (N_1813,N_113,N_114);
nor U1814 (N_1814,N_297,N_849);
nand U1815 (N_1815,N_613,N_1058);
nor U1816 (N_1816,In_2220,N_49);
xnor U1817 (N_1817,N_555,In_2646);
nand U1818 (N_1818,In_2149,N_878);
nand U1819 (N_1819,In_2013,N_704);
xnor U1820 (N_1820,N_932,N_922);
or U1821 (N_1821,In_1871,N_310);
nand U1822 (N_1822,In_2493,N_575);
or U1823 (N_1823,N_1017,N_662);
and U1824 (N_1824,N_361,N_903);
or U1825 (N_1825,In_625,N_834);
nand U1826 (N_1826,N_729,In_622);
or U1827 (N_1827,N_740,N_615);
and U1828 (N_1828,N_1148,N_41);
nor U1829 (N_1829,N_231,N_493);
and U1830 (N_1830,N_677,N_980);
nand U1831 (N_1831,N_767,In_1003);
nand U1832 (N_1832,N_605,N_277);
xor U1833 (N_1833,In_1281,N_65);
nor U1834 (N_1834,N_12,N_799);
nor U1835 (N_1835,In_1902,N_544);
nor U1836 (N_1836,N_1031,N_628);
nand U1837 (N_1837,N_833,N_491);
or U1838 (N_1838,N_612,In_2701);
nor U1839 (N_1839,In_2488,N_692);
nand U1840 (N_1840,N_594,In_480);
nor U1841 (N_1841,N_790,In_817);
and U1842 (N_1842,N_770,In_1173);
or U1843 (N_1843,In_2437,In_430);
and U1844 (N_1844,N_1096,In_2866);
and U1845 (N_1845,N_1004,In_2100);
nor U1846 (N_1846,N_240,In_40);
nand U1847 (N_1847,N_354,In_2156);
nor U1848 (N_1848,N_20,N_1002);
and U1849 (N_1849,N_75,In_2922);
nor U1850 (N_1850,In_1875,N_1107);
and U1851 (N_1851,N_573,In_496);
or U1852 (N_1852,In_54,N_884);
and U1853 (N_1853,In_1023,In_386);
nor U1854 (N_1854,In_2399,N_1178);
or U1855 (N_1855,N_365,In_1628);
and U1856 (N_1856,N_1032,N_1158);
xnor U1857 (N_1857,N_187,In_929);
nand U1858 (N_1858,In_2065,N_406);
xnor U1859 (N_1859,N_1078,In_2000);
nand U1860 (N_1860,N_1053,In_2893);
nand U1861 (N_1861,N_1069,N_602);
xnor U1862 (N_1862,N_140,N_1040);
nor U1863 (N_1863,N_389,N_1011);
xnor U1864 (N_1864,N_459,In_2512);
xor U1865 (N_1865,In_51,N_1093);
nand U1866 (N_1866,N_353,N_786);
nor U1867 (N_1867,N_532,In_618);
nand U1868 (N_1868,In_2132,In_1268);
nand U1869 (N_1869,N_576,In_323);
xnor U1870 (N_1870,N_915,N_132);
nor U1871 (N_1871,In_434,N_1106);
and U1872 (N_1872,N_968,In_2215);
and U1873 (N_1873,N_867,N_433);
and U1874 (N_1874,In_2518,In_559);
nor U1875 (N_1875,N_1168,N_727);
nor U1876 (N_1876,N_127,N_105);
or U1877 (N_1877,N_393,N_104);
and U1878 (N_1878,In_2805,N_430);
or U1879 (N_1879,N_881,In_1328);
or U1880 (N_1880,In_260,N_110);
xnor U1881 (N_1881,N_536,N_117);
xor U1882 (N_1882,N_275,In_2877);
xnor U1883 (N_1883,N_585,In_731);
nand U1884 (N_1884,In_1881,In_489);
and U1885 (N_1885,N_1028,N_299);
and U1886 (N_1886,N_840,N_854);
or U1887 (N_1887,N_1120,In_2256);
and U1888 (N_1888,N_376,In_1672);
nand U1889 (N_1889,N_534,N_423);
or U1890 (N_1890,N_728,N_40);
and U1891 (N_1891,N_346,N_185);
or U1892 (N_1892,N_97,In_2373);
and U1893 (N_1893,N_1117,N_593);
and U1894 (N_1894,In_2223,In_2696);
xor U1895 (N_1895,In_1862,N_710);
xnor U1896 (N_1896,N_1153,In_974);
or U1897 (N_1897,N_1132,N_476);
xor U1898 (N_1898,N_403,In_193);
xnor U1899 (N_1899,N_149,N_55);
and U1900 (N_1900,N_860,In_2525);
nor U1901 (N_1901,N_640,N_589);
and U1902 (N_1902,N_558,In_272);
xnor U1903 (N_1903,In_1680,In_10);
or U1904 (N_1904,N_945,N_1191);
nand U1905 (N_1905,In_2686,N_1019);
and U1906 (N_1906,In_259,N_950);
xor U1907 (N_1907,N_305,In_1804);
nand U1908 (N_1908,N_1100,In_1868);
nor U1909 (N_1909,N_326,In_1619);
nor U1910 (N_1910,In_2213,N_847);
nand U1911 (N_1911,N_1194,N_398);
and U1912 (N_1912,N_159,N_595);
xor U1913 (N_1913,N_292,N_750);
nor U1914 (N_1914,In_823,In_1071);
or U1915 (N_1915,N_774,In_2655);
or U1916 (N_1916,In_1279,N_913);
or U1917 (N_1917,In_1965,N_803);
nor U1918 (N_1918,N_713,In_52);
nor U1919 (N_1919,N_427,In_2460);
and U1920 (N_1920,In_1396,N_655);
or U1921 (N_1921,N_99,In_1761);
or U1922 (N_1922,In_2879,In_2113);
xor U1923 (N_1923,N_154,In_511);
and U1924 (N_1924,In_271,N_496);
xnor U1925 (N_1925,N_189,N_283);
nor U1926 (N_1926,N_1108,N_666);
nor U1927 (N_1927,N_309,In_2740);
xnor U1928 (N_1928,N_1080,In_45);
nor U1929 (N_1929,N_708,N_147);
and U1930 (N_1930,N_547,N_303);
or U1931 (N_1931,N_1036,In_714);
nor U1932 (N_1932,N_311,N_261);
and U1933 (N_1933,In_243,N_1192);
or U1934 (N_1934,N_458,In_2748);
nand U1935 (N_1935,N_492,In_1853);
or U1936 (N_1936,N_1154,N_137);
nand U1937 (N_1937,N_970,N_490);
nor U1938 (N_1938,In_800,In_838);
or U1939 (N_1939,In_717,In_1954);
xor U1940 (N_1940,N_664,N_868);
xor U1941 (N_1941,N_1127,In_1986);
or U1942 (N_1942,N_399,N_440);
and U1943 (N_1943,N_853,N_456);
and U1944 (N_1944,N_39,N_819);
xor U1945 (N_1945,In_2822,In_1238);
nor U1946 (N_1946,N_4,In_1699);
nor U1947 (N_1947,In_1537,N_334);
xor U1948 (N_1948,In_224,N_325);
xnor U1949 (N_1949,N_237,N_893);
and U1950 (N_1950,In_1333,N_1022);
or U1951 (N_1951,N_0,N_451);
nor U1952 (N_1952,N_449,In_2064);
nor U1953 (N_1953,N_192,N_249);
and U1954 (N_1954,In_2734,N_835);
or U1955 (N_1955,N_1119,N_757);
nor U1956 (N_1956,In_2549,N_1180);
nor U1957 (N_1957,N_985,In_1243);
and U1958 (N_1958,In_2485,In_239);
nor U1959 (N_1959,N_395,In_541);
nand U1960 (N_1960,N_1043,N_967);
nand U1961 (N_1961,N_135,In_2545);
xor U1962 (N_1962,In_752,N_954);
xor U1963 (N_1963,N_291,In_2419);
or U1964 (N_1964,N_35,N_639);
nor U1965 (N_1965,N_850,N_475);
and U1966 (N_1966,In_2606,N_138);
nand U1967 (N_1967,N_165,In_2676);
and U1968 (N_1968,N_510,N_330);
xor U1969 (N_1969,N_1089,In_221);
nand U1970 (N_1970,N_538,In_2404);
or U1971 (N_1971,N_754,N_1016);
nor U1972 (N_1972,In_390,N_331);
xnor U1973 (N_1973,N_643,N_697);
nor U1974 (N_1974,In_2109,N_545);
or U1975 (N_1975,In_76,N_680);
and U1976 (N_1976,N_658,N_396);
nor U1977 (N_1977,N_238,N_136);
xnor U1978 (N_1978,N_352,N_139);
nor U1979 (N_1979,In_356,In_1340);
xor U1980 (N_1980,N_561,N_194);
nor U1981 (N_1981,N_2,N_13);
and U1982 (N_1982,N_30,N_601);
or U1983 (N_1983,N_293,In_1720);
and U1984 (N_1984,N_411,N_1049);
and U1985 (N_1985,N_1189,N_875);
nor U1986 (N_1986,N_986,In_580);
nand U1987 (N_1987,In_2052,N_505);
and U1988 (N_1988,N_1003,N_235);
or U1989 (N_1989,N_378,In_1709);
or U1990 (N_1990,In_1378,N_693);
nand U1991 (N_1991,N_925,N_1010);
xor U1992 (N_1992,N_145,N_484);
and U1993 (N_1993,N_699,N_650);
or U1994 (N_1994,N_244,N_805);
nand U1995 (N_1995,N_966,N_606);
or U1996 (N_1996,In_84,In_1541);
and U1997 (N_1997,In_2775,N_1041);
or U1998 (N_1998,N_1139,N_629);
and U1999 (N_1999,N_44,In_112);
or U2000 (N_2000,In_268,N_924);
nor U2001 (N_2001,In_1936,N_784);
nand U2002 (N_2002,In_43,N_769);
nand U2003 (N_2003,In_494,N_772);
nand U2004 (N_2004,N_1095,In_1);
nor U2005 (N_2005,N_895,In_1476);
xnor U2006 (N_2006,N_632,In_1574);
and U2007 (N_2007,N_1188,N_508);
xor U2008 (N_2008,N_1140,In_1612);
nand U2009 (N_2009,N_1052,N_253);
xor U2010 (N_2010,N_624,In_1715);
xor U2011 (N_2011,In_2044,N_381);
and U2012 (N_2012,N_188,N_485);
or U2013 (N_2013,In_1127,In_2913);
xnor U2014 (N_2014,In_1996,In_2772);
nor U2015 (N_2015,N_822,N_818);
xor U2016 (N_2016,N_682,In_137);
nand U2017 (N_2017,N_886,N_953);
xor U2018 (N_2018,N_793,N_848);
or U2019 (N_2019,N_123,N_1165);
nor U2020 (N_2020,In_2526,In_2716);
nor U2021 (N_2021,In_2016,N_600);
nor U2022 (N_2022,In_1177,N_86);
xor U2023 (N_2023,N_1059,In_1449);
nor U2024 (N_2024,N_372,N_731);
nor U2025 (N_2025,In_452,N_709);
nor U2026 (N_2026,In_2610,In_2284);
nor U2027 (N_2027,N_514,In_104);
nor U2028 (N_2028,N_686,In_285);
xnor U2029 (N_2029,N_695,N_714);
and U2030 (N_2030,N_384,N_1038);
and U2031 (N_2031,N_420,N_178);
and U2032 (N_2032,N_559,In_2540);
or U2033 (N_2033,In_2576,In_2278);
nand U2034 (N_2034,In_2445,N_470);
and U2035 (N_2035,N_308,N_935);
nand U2036 (N_2036,In_2961,N_703);
nand U2037 (N_2037,In_2522,In_1569);
xor U2038 (N_2038,N_839,In_55);
xnor U2039 (N_2039,N_347,N_438);
xor U2040 (N_2040,N_225,N_1076);
and U2041 (N_2041,N_864,N_289);
or U2042 (N_2042,N_940,N_566);
xor U2043 (N_2043,N_222,In_732);
xnor U2044 (N_2044,N_1042,N_687);
nand U2045 (N_2045,N_694,N_636);
and U2046 (N_2046,In_46,In_1379);
and U2047 (N_2047,In_563,N_294);
nand U2048 (N_2048,N_1046,N_1126);
nor U2049 (N_2049,N_965,In_1828);
nor U2050 (N_2050,In_2510,In_665);
or U2051 (N_2051,N_232,N_930);
nand U2052 (N_2052,N_401,N_800);
nor U2053 (N_2053,N_1071,In_2706);
and U2054 (N_2054,In_683,N_1111);
nand U2055 (N_2055,In_2217,In_2984);
or U2056 (N_2056,N_327,N_390);
xor U2057 (N_2057,N_426,N_1136);
or U2058 (N_2058,In_826,N_446);
or U2059 (N_2059,N_899,N_88);
xor U2060 (N_2060,N_972,N_301);
xor U2061 (N_2061,N_974,N_956);
nor U2062 (N_2062,N_419,In_1779);
nor U2063 (N_2063,In_1412,N_392);
and U2064 (N_2064,In_884,N_34);
or U2065 (N_2065,In_2779,In_2939);
xnor U2066 (N_2066,N_719,N_22);
nand U2067 (N_2067,N_201,N_550);
or U2068 (N_2068,N_98,N_359);
nand U2069 (N_2069,N_901,N_977);
nor U2070 (N_2070,In_1798,N_802);
or U2071 (N_2071,In_953,N_43);
nor U2072 (N_2072,In_2188,N_204);
and U2073 (N_2073,N_262,N_667);
nor U2074 (N_2074,In_1947,N_11);
nand U2075 (N_2075,In_542,N_1);
nand U2076 (N_2076,In_117,N_391);
nor U2077 (N_2077,N_263,In_473);
or U2078 (N_2078,N_747,In_160);
nand U2079 (N_2079,In_1958,N_161);
nand U2080 (N_2080,In_425,N_1171);
nor U2081 (N_2081,In_2366,N_810);
or U2082 (N_2082,In_283,N_911);
nor U2083 (N_2083,N_150,N_109);
nand U2084 (N_2084,In_2670,N_69);
nand U2085 (N_2085,N_469,N_923);
xor U2086 (N_2086,In_2799,N_609);
nor U2087 (N_2087,N_988,N_683);
xor U2088 (N_2088,N_63,N_1172);
nand U2089 (N_2089,N_921,N_1152);
xnor U2090 (N_2090,N_181,N_763);
nand U2091 (N_2091,N_838,N_21);
xor U2092 (N_2092,N_76,N_196);
nand U2093 (N_2093,In_1555,N_502);
nor U2094 (N_2094,In_1472,N_841);
and U2095 (N_2095,In_2348,N_603);
xnor U2096 (N_2096,N_1039,N_736);
nor U2097 (N_2097,N_1033,In_1682);
nand U2098 (N_2098,N_1054,N_874);
nand U2099 (N_2099,In_2644,N_241);
or U2100 (N_2100,N_1085,N_694);
nor U2101 (N_2101,In_1898,In_103);
nand U2102 (N_2102,In_906,In_2156);
xor U2103 (N_2103,N_160,N_89);
and U2104 (N_2104,N_676,In_2913);
xnor U2105 (N_2105,N_294,N_292);
xnor U2106 (N_2106,N_193,N_899);
or U2107 (N_2107,N_333,In_1555);
xnor U2108 (N_2108,N_958,N_818);
or U2109 (N_2109,N_830,N_949);
nor U2110 (N_2110,N_953,N_557);
xnor U2111 (N_2111,N_680,In_1396);
nor U2112 (N_2112,N_12,N_740);
xnor U2113 (N_2113,N_685,N_43);
nand U2114 (N_2114,N_619,N_681);
or U2115 (N_2115,N_419,N_581);
and U2116 (N_2116,In_646,In_1871);
nand U2117 (N_2117,N_1186,N_861);
nand U2118 (N_2118,In_2434,In_2404);
xor U2119 (N_2119,N_564,N_828);
nor U2120 (N_2120,N_417,In_2706);
nor U2121 (N_2121,N_210,N_1165);
xor U2122 (N_2122,N_1096,N_1022);
nor U2123 (N_2123,N_308,In_43);
or U2124 (N_2124,In_2202,N_223);
nor U2125 (N_2125,N_499,In_2215);
xnor U2126 (N_2126,N_520,N_333);
xnor U2127 (N_2127,In_2545,N_1094);
or U2128 (N_2128,N_858,N_902);
or U2129 (N_2129,N_796,N_961);
xnor U2130 (N_2130,N_879,N_496);
nand U2131 (N_2131,N_798,N_29);
nor U2132 (N_2132,In_1455,N_198);
and U2133 (N_2133,N_463,N_793);
and U2134 (N_2134,N_192,In_1882);
nand U2135 (N_2135,N_675,N_790);
xnor U2136 (N_2136,N_805,N_343);
nor U2137 (N_2137,In_1305,N_935);
or U2138 (N_2138,N_677,N_783);
xnor U2139 (N_2139,N_13,N_1012);
and U2140 (N_2140,N_642,N_793);
nand U2141 (N_2141,In_981,In_2633);
and U2142 (N_2142,In_1554,In_987);
and U2143 (N_2143,In_166,N_990);
and U2144 (N_2144,N_9,N_1056);
or U2145 (N_2145,In_2879,N_681);
xor U2146 (N_2146,N_476,N_233);
nand U2147 (N_2147,N_624,In_679);
and U2148 (N_2148,N_450,N_1191);
or U2149 (N_2149,N_180,N_1133);
or U2150 (N_2150,In_792,N_1066);
xnor U2151 (N_2151,N_628,In_1804);
and U2152 (N_2152,N_749,N_768);
and U2153 (N_2153,In_1882,N_598);
xnor U2154 (N_2154,In_2549,N_141);
or U2155 (N_2155,N_760,In_18);
nor U2156 (N_2156,N_177,In_78);
and U2157 (N_2157,N_827,N_880);
or U2158 (N_2158,In_221,N_898);
or U2159 (N_2159,N_672,In_2708);
or U2160 (N_2160,N_811,N_109);
xnor U2161 (N_2161,In_1952,N_1020);
nor U2162 (N_2162,N_381,In_1523);
or U2163 (N_2163,N_467,N_1181);
nor U2164 (N_2164,In_795,N_905);
nor U2165 (N_2165,N_1162,N_1165);
nor U2166 (N_2166,N_492,N_630);
and U2167 (N_2167,N_417,N_293);
and U2168 (N_2168,In_1013,N_955);
or U2169 (N_2169,In_134,In_536);
xnor U2170 (N_2170,N_748,N_244);
nor U2171 (N_2171,N_646,N_824);
xnor U2172 (N_2172,N_678,N_478);
and U2173 (N_2173,N_430,In_1266);
nand U2174 (N_2174,N_471,In_706);
nand U2175 (N_2175,In_2320,N_649);
nand U2176 (N_2176,N_413,N_21);
xor U2177 (N_2177,N_476,N_633);
and U2178 (N_2178,N_1126,N_78);
and U2179 (N_2179,N_187,In_54);
nand U2180 (N_2180,In_1715,In_55);
xor U2181 (N_2181,In_134,N_487);
nand U2182 (N_2182,N_144,In_2568);
or U2183 (N_2183,N_427,N_1175);
nor U2184 (N_2184,In_2242,In_248);
or U2185 (N_2185,In_1148,In_752);
nand U2186 (N_2186,In_1325,In_2062);
nand U2187 (N_2187,In_2732,N_677);
nor U2188 (N_2188,N_174,In_1834);
nor U2189 (N_2189,N_488,N_809);
nor U2190 (N_2190,In_1328,In_542);
xnor U2191 (N_2191,N_418,In_2057);
xor U2192 (N_2192,N_155,N_379);
xnor U2193 (N_2193,N_837,N_20);
nor U2194 (N_2194,N_1090,N_562);
xor U2195 (N_2195,In_93,N_654);
and U2196 (N_2196,N_152,In_2576);
nand U2197 (N_2197,N_912,N_1102);
or U2198 (N_2198,N_1161,In_355);
and U2199 (N_2199,In_224,In_2707);
nand U2200 (N_2200,In_2391,N_360);
or U2201 (N_2201,N_410,N_889);
and U2202 (N_2202,In_824,N_660);
xnor U2203 (N_2203,In_2653,In_2445);
nand U2204 (N_2204,N_1119,N_824);
and U2205 (N_2205,N_1192,N_229);
nor U2206 (N_2206,N_835,N_361);
or U2207 (N_2207,In_2321,N_913);
nor U2208 (N_2208,In_1438,In_2322);
or U2209 (N_2209,N_1066,N_771);
nand U2210 (N_2210,N_1147,N_989);
xnor U2211 (N_2211,N_898,N_1178);
and U2212 (N_2212,N_144,In_268);
nand U2213 (N_2213,N_1177,N_110);
xnor U2214 (N_2214,N_297,In_2775);
nor U2215 (N_2215,N_80,In_2570);
or U2216 (N_2216,N_376,N_228);
and U2217 (N_2217,N_642,In_2708);
xor U2218 (N_2218,N_140,In_1340);
xor U2219 (N_2219,N_88,In_2526);
or U2220 (N_2220,N_136,N_422);
xor U2221 (N_2221,In_1912,N_1014);
or U2222 (N_2222,In_675,N_239);
nand U2223 (N_2223,N_747,N_1180);
nor U2224 (N_2224,In_2395,In_2526);
or U2225 (N_2225,N_114,N_618);
and U2226 (N_2226,N_468,N_771);
or U2227 (N_2227,N_313,N_270);
or U2228 (N_2228,In_1645,N_950);
xor U2229 (N_2229,N_40,In_1082);
nor U2230 (N_2230,N_729,In_1127);
nand U2231 (N_2231,In_1773,N_322);
xnor U2232 (N_2232,In_1525,N_425);
nand U2233 (N_2233,N_972,N_293);
nor U2234 (N_2234,N_727,In_329);
or U2235 (N_2235,In_939,N_987);
or U2236 (N_2236,N_800,N_443);
xnor U2237 (N_2237,In_103,N_150);
or U2238 (N_2238,N_64,N_416);
nand U2239 (N_2239,N_147,In_282);
and U2240 (N_2240,N_709,In_1331);
nor U2241 (N_2241,N_58,N_33);
and U2242 (N_2242,In_1577,In_1958);
xnor U2243 (N_2243,N_99,N_307);
nor U2244 (N_2244,N_897,N_321);
or U2245 (N_2245,N_725,In_563);
and U2246 (N_2246,In_58,N_638);
or U2247 (N_2247,In_410,N_53);
nand U2248 (N_2248,N_1134,N_476);
xor U2249 (N_2249,N_667,In_1378);
or U2250 (N_2250,In_1325,In_1148);
xor U2251 (N_2251,N_295,N_1001);
and U2252 (N_2252,N_191,N_777);
or U2253 (N_2253,N_868,N_650);
xnor U2254 (N_2254,In_1983,In_265);
xor U2255 (N_2255,N_821,N_363);
nor U2256 (N_2256,N_354,In_280);
and U2257 (N_2257,In_1228,N_915);
xnor U2258 (N_2258,N_437,N_940);
nor U2259 (N_2259,N_634,In_2513);
and U2260 (N_2260,N_371,N_746);
and U2261 (N_2261,In_2373,N_920);
or U2262 (N_2262,In_1074,N_181);
xor U2263 (N_2263,In_1238,N_518);
xor U2264 (N_2264,N_1006,In_2123);
and U2265 (N_2265,N_806,N_319);
xnor U2266 (N_2266,In_2278,In_1673);
nand U2267 (N_2267,In_2214,N_1132);
nor U2268 (N_2268,N_918,N_114);
nand U2269 (N_2269,In_551,In_2765);
nor U2270 (N_2270,N_574,N_120);
nor U2271 (N_2271,In_1798,In_1177);
or U2272 (N_2272,N_354,N_779);
and U2273 (N_2273,N_324,N_1049);
xor U2274 (N_2274,N_1116,In_84);
xor U2275 (N_2275,N_1196,N_984);
nor U2276 (N_2276,N_964,In_1105);
and U2277 (N_2277,In_2188,In_684);
and U2278 (N_2278,N_895,N_905);
and U2279 (N_2279,In_706,N_376);
and U2280 (N_2280,In_1644,In_2501);
or U2281 (N_2281,N_651,N_646);
nor U2282 (N_2282,In_2215,In_164);
or U2283 (N_2283,In_805,N_1166);
xnor U2284 (N_2284,N_487,N_236);
xor U2285 (N_2285,In_2488,N_1093);
nor U2286 (N_2286,N_652,N_970);
xnor U2287 (N_2287,N_409,In_17);
xnor U2288 (N_2288,N_528,N_584);
and U2289 (N_2289,In_1874,N_1166);
xor U2290 (N_2290,In_795,In_1031);
xor U2291 (N_2291,In_1130,In_2867);
nor U2292 (N_2292,N_333,N_106);
or U2293 (N_2293,N_1163,N_213);
nor U2294 (N_2294,N_92,N_835);
and U2295 (N_2295,N_572,In_1177);
xor U2296 (N_2296,N_1069,N_801);
and U2297 (N_2297,N_1012,N_54);
nand U2298 (N_2298,N_191,In_148);
xor U2299 (N_2299,In_1486,In_1440);
and U2300 (N_2300,N_547,In_489);
or U2301 (N_2301,N_1109,N_970);
xnor U2302 (N_2302,In_2676,In_1720);
or U2303 (N_2303,In_2252,N_23);
and U2304 (N_2304,N_1159,N_652);
nor U2305 (N_2305,In_1891,N_1094);
and U2306 (N_2306,N_246,N_288);
or U2307 (N_2307,N_630,N_467);
or U2308 (N_2308,N_918,N_138);
or U2309 (N_2309,N_1105,N_306);
or U2310 (N_2310,N_337,In_838);
or U2311 (N_2311,In_622,N_81);
or U2312 (N_2312,N_758,In_2321);
nand U2313 (N_2313,N_853,N_55);
xor U2314 (N_2314,In_2901,N_942);
xor U2315 (N_2315,N_423,In_1871);
or U2316 (N_2316,N_548,N_204);
xor U2317 (N_2317,In_1343,In_792);
and U2318 (N_2318,N_99,N_189);
and U2319 (N_2319,N_818,N_508);
xnor U2320 (N_2320,In_2136,N_932);
nand U2321 (N_2321,N_259,In_2675);
xor U2322 (N_2322,N_853,N_643);
or U2323 (N_2323,In_2278,N_1067);
or U2324 (N_2324,N_551,In_494);
nand U2325 (N_2325,In_2034,N_1148);
nor U2326 (N_2326,N_701,N_466);
and U2327 (N_2327,N_1019,N_926);
and U2328 (N_2328,N_971,N_1111);
and U2329 (N_2329,N_776,N_385);
xnor U2330 (N_2330,N_118,N_61);
and U2331 (N_2331,In_850,N_441);
or U2332 (N_2332,N_710,N_321);
or U2333 (N_2333,N_610,N_1090);
xnor U2334 (N_2334,In_1202,In_1540);
nand U2335 (N_2335,In_479,N_826);
or U2336 (N_2336,In_2585,In_2525);
nand U2337 (N_2337,In_2772,N_602);
xnor U2338 (N_2338,N_651,N_548);
or U2339 (N_2339,In_929,N_292);
nand U2340 (N_2340,N_932,N_399);
nand U2341 (N_2341,N_251,N_43);
and U2342 (N_2342,N_1163,N_655);
nand U2343 (N_2343,N_1014,In_1890);
xnor U2344 (N_2344,In_88,N_708);
nor U2345 (N_2345,N_883,N_1146);
nand U2346 (N_2346,N_841,N_938);
xor U2347 (N_2347,N_30,In_2188);
and U2348 (N_2348,In_511,N_866);
nor U2349 (N_2349,N_993,N_1017);
xor U2350 (N_2350,In_1328,N_977);
or U2351 (N_2351,In_480,N_169);
xnor U2352 (N_2352,N_381,N_176);
and U2353 (N_2353,In_10,N_1018);
and U2354 (N_2354,N_678,In_1794);
or U2355 (N_2355,In_48,In_2869);
nand U2356 (N_2356,N_57,N_271);
nand U2357 (N_2357,N_548,N_11);
nor U2358 (N_2358,N_1094,N_601);
xor U2359 (N_2359,In_386,N_20);
nand U2360 (N_2360,In_541,In_2407);
nor U2361 (N_2361,N_46,In_1230);
and U2362 (N_2362,N_68,In_1644);
nand U2363 (N_2363,N_1030,In_1612);
and U2364 (N_2364,N_812,In_2223);
nand U2365 (N_2365,N_295,N_647);
nor U2366 (N_2366,N_822,In_2111);
or U2367 (N_2367,N_89,In_277);
nor U2368 (N_2368,N_449,N_229);
nor U2369 (N_2369,N_617,N_555);
or U2370 (N_2370,In_1682,In_1912);
nor U2371 (N_2371,N_98,N_40);
or U2372 (N_2372,N_138,In_587);
or U2373 (N_2373,In_1727,In_2188);
or U2374 (N_2374,N_54,N_951);
and U2375 (N_2375,N_95,In_2360);
or U2376 (N_2376,N_363,N_530);
and U2377 (N_2377,N_389,In_2016);
xnor U2378 (N_2378,N_297,N_163);
xnor U2379 (N_2379,N_966,N_274);
xor U2380 (N_2380,In_2893,N_435);
nor U2381 (N_2381,In_1680,N_32);
and U2382 (N_2382,N_553,N_555);
nand U2383 (N_2383,N_561,N_1155);
or U2384 (N_2384,In_908,In_2565);
xor U2385 (N_2385,N_839,In_2649);
nand U2386 (N_2386,In_2996,N_255);
and U2387 (N_2387,In_811,N_213);
xor U2388 (N_2388,N_253,N_466);
nor U2389 (N_2389,N_794,In_2300);
nand U2390 (N_2390,In_1293,N_956);
nor U2391 (N_2391,N_101,In_2772);
xor U2392 (N_2392,In_1786,N_317);
xor U2393 (N_2393,In_1871,N_63);
nand U2394 (N_2394,N_204,N_429);
nor U2395 (N_2395,N_341,N_26);
nor U2396 (N_2396,In_684,N_853);
nor U2397 (N_2397,N_403,N_526);
nor U2398 (N_2398,In_987,N_550);
and U2399 (N_2399,In_1619,N_17);
nor U2400 (N_2400,N_1808,N_1279);
or U2401 (N_2401,N_1696,N_2066);
and U2402 (N_2402,N_2004,N_1304);
nand U2403 (N_2403,N_1705,N_1989);
and U2404 (N_2404,N_1425,N_1249);
nor U2405 (N_2405,N_2165,N_2217);
or U2406 (N_2406,N_2195,N_1883);
xor U2407 (N_2407,N_1708,N_1536);
nor U2408 (N_2408,N_1202,N_1839);
and U2409 (N_2409,N_1450,N_1684);
or U2410 (N_2410,N_2152,N_1353);
nor U2411 (N_2411,N_1558,N_2189);
or U2412 (N_2412,N_1618,N_2353);
or U2413 (N_2413,N_1910,N_2269);
nand U2414 (N_2414,N_2324,N_2090);
or U2415 (N_2415,N_2164,N_1465);
xor U2416 (N_2416,N_2247,N_2027);
nor U2417 (N_2417,N_1607,N_1673);
or U2418 (N_2418,N_1683,N_1534);
or U2419 (N_2419,N_2369,N_2373);
and U2420 (N_2420,N_1965,N_1832);
nand U2421 (N_2421,N_1755,N_2289);
and U2422 (N_2422,N_1648,N_1357);
and U2423 (N_2423,N_1571,N_2378);
nor U2424 (N_2424,N_2239,N_2209);
nand U2425 (N_2425,N_2257,N_1524);
and U2426 (N_2426,N_1897,N_1994);
xnor U2427 (N_2427,N_1819,N_2030);
xor U2428 (N_2428,N_1938,N_1513);
and U2429 (N_2429,N_1221,N_1688);
or U2430 (N_2430,N_2042,N_1235);
or U2431 (N_2431,N_1596,N_1500);
nor U2432 (N_2432,N_2077,N_1733);
xnor U2433 (N_2433,N_1559,N_1468);
or U2434 (N_2434,N_1506,N_2229);
and U2435 (N_2435,N_2120,N_1763);
nor U2436 (N_2436,N_1740,N_1486);
nor U2437 (N_2437,N_1981,N_1805);
nor U2438 (N_2438,N_2387,N_1544);
nand U2439 (N_2439,N_1416,N_2376);
xor U2440 (N_2440,N_2351,N_1514);
nor U2441 (N_2441,N_1713,N_1384);
and U2442 (N_2442,N_1459,N_1622);
nand U2443 (N_2443,N_1937,N_1847);
xnor U2444 (N_2444,N_1973,N_1380);
or U2445 (N_2445,N_1282,N_1944);
and U2446 (N_2446,N_1511,N_1549);
nor U2447 (N_2447,N_2395,N_1519);
and U2448 (N_2448,N_1849,N_1901);
nand U2449 (N_2449,N_1369,N_1855);
or U2450 (N_2450,N_2226,N_1941);
and U2451 (N_2451,N_1592,N_2242);
xnor U2452 (N_2452,N_1766,N_1335);
or U2453 (N_2453,N_2287,N_2001);
and U2454 (N_2454,N_1890,N_1798);
xor U2455 (N_2455,N_1846,N_1390);
nor U2456 (N_2456,N_2026,N_2052);
nor U2457 (N_2457,N_1619,N_1631);
nand U2458 (N_2458,N_1389,N_1757);
nand U2459 (N_2459,N_1480,N_1344);
and U2460 (N_2460,N_1496,N_2106);
nor U2461 (N_2461,N_2051,N_2199);
nand U2462 (N_2462,N_1200,N_2285);
and U2463 (N_2463,N_1617,N_1752);
nor U2464 (N_2464,N_1709,N_1430);
nor U2465 (N_2465,N_2187,N_2200);
nand U2466 (N_2466,N_1780,N_2315);
and U2467 (N_2467,N_1328,N_2291);
nor U2468 (N_2468,N_1347,N_2197);
and U2469 (N_2469,N_1546,N_1322);
nand U2470 (N_2470,N_1358,N_1845);
xnor U2471 (N_2471,N_1676,N_1306);
xnor U2472 (N_2472,N_1966,N_1820);
or U2473 (N_2473,N_1783,N_1552);
nand U2474 (N_2474,N_1632,N_1640);
nor U2475 (N_2475,N_1262,N_2091);
xor U2476 (N_2476,N_2254,N_2363);
nor U2477 (N_2477,N_2274,N_1442);
nor U2478 (N_2478,N_1630,N_1972);
nand U2479 (N_2479,N_2244,N_1414);
nor U2480 (N_2480,N_1257,N_1287);
or U2481 (N_2481,N_1641,N_1576);
nand U2482 (N_2482,N_2270,N_2080);
nand U2483 (N_2483,N_2009,N_1472);
xor U2484 (N_2484,N_1356,N_1337);
and U2485 (N_2485,N_2006,N_2007);
and U2486 (N_2486,N_1204,N_2109);
xnor U2487 (N_2487,N_1214,N_1542);
or U2488 (N_2488,N_1332,N_1577);
and U2489 (N_2489,N_1499,N_2172);
or U2490 (N_2490,N_1916,N_2010);
xor U2491 (N_2491,N_1624,N_1557);
nand U2492 (N_2492,N_1428,N_2029);
nor U2493 (N_2493,N_2094,N_1244);
nor U2494 (N_2494,N_1403,N_1764);
xor U2495 (N_2495,N_1889,N_2379);
or U2496 (N_2496,N_1875,N_1361);
or U2497 (N_2497,N_1957,N_1762);
and U2498 (N_2498,N_2215,N_1907);
or U2499 (N_2499,N_1949,N_1302);
nand U2500 (N_2500,N_1867,N_1217);
nand U2501 (N_2501,N_1948,N_1674);
nor U2502 (N_2502,N_1610,N_1888);
or U2503 (N_2503,N_2138,N_1288);
and U2504 (N_2504,N_2156,N_2390);
and U2505 (N_2505,N_1754,N_2345);
and U2506 (N_2506,N_2268,N_2064);
nor U2507 (N_2507,N_1788,N_1990);
nor U2508 (N_2508,N_1575,N_1609);
and U2509 (N_2509,N_2313,N_1869);
or U2510 (N_2510,N_2394,N_2129);
nor U2511 (N_2511,N_2063,N_1971);
or U2512 (N_2512,N_1354,N_1921);
nor U2513 (N_2513,N_1457,N_1427);
and U2514 (N_2514,N_2277,N_1809);
xor U2515 (N_2515,N_2035,N_2374);
and U2516 (N_2516,N_1939,N_2075);
xnor U2517 (N_2517,N_2320,N_1914);
nor U2518 (N_2518,N_2162,N_2005);
xor U2519 (N_2519,N_1848,N_1532);
nand U2520 (N_2520,N_1378,N_1580);
and U2521 (N_2521,N_1717,N_1697);
and U2522 (N_2522,N_1293,N_1738);
nand U2523 (N_2523,N_1995,N_1877);
xor U2524 (N_2524,N_1586,N_2062);
or U2525 (N_2525,N_2074,N_1613);
or U2526 (N_2526,N_1870,N_1979);
and U2527 (N_2527,N_1554,N_1926);
nor U2528 (N_2528,N_2155,N_1872);
xnor U2529 (N_2529,N_1386,N_1658);
nand U2530 (N_2530,N_1963,N_2382);
nand U2531 (N_2531,N_1844,N_1829);
nand U2532 (N_2532,N_2233,N_2208);
or U2533 (N_2533,N_1518,N_1765);
xnor U2534 (N_2534,N_2136,N_2015);
xnor U2535 (N_2535,N_1821,N_1647);
or U2536 (N_2536,N_1311,N_1290);
or U2537 (N_2537,N_1718,N_2142);
xnor U2538 (N_2538,N_2347,N_1635);
or U2539 (N_2539,N_1321,N_1999);
or U2540 (N_2540,N_1842,N_1746);
or U2541 (N_2541,N_2107,N_1993);
nand U2542 (N_2542,N_1315,N_1372);
nor U2543 (N_2543,N_1387,N_1258);
nor U2544 (N_2544,N_1953,N_1810);
xor U2545 (N_2545,N_1970,N_1830);
xnor U2546 (N_2546,N_1651,N_1538);
xor U2547 (N_2547,N_1227,N_2144);
and U2548 (N_2548,N_1209,N_1785);
or U2549 (N_2549,N_1976,N_1983);
and U2550 (N_2550,N_1878,N_2275);
nor U2551 (N_2551,N_1594,N_1233);
nor U2552 (N_2552,N_2216,N_2262);
or U2553 (N_2553,N_1621,N_1815);
or U2554 (N_2554,N_1736,N_1417);
and U2555 (N_2555,N_1539,N_1681);
and U2556 (N_2556,N_1439,N_1404);
and U2557 (N_2557,N_1488,N_1352);
xnor U2558 (N_2558,N_2218,N_1327);
nor U2559 (N_2559,N_1528,N_1634);
and U2560 (N_2560,N_1495,N_1769);
nand U2561 (N_2561,N_1894,N_2076);
nor U2562 (N_2562,N_1723,N_1779);
or U2563 (N_2563,N_1230,N_2352);
nand U2564 (N_2564,N_1961,N_1711);
xnor U2565 (N_2565,N_1716,N_1947);
nand U2566 (N_2566,N_1413,N_1350);
xor U2567 (N_2567,N_1261,N_2097);
or U2568 (N_2568,N_2253,N_1215);
or U2569 (N_2569,N_1366,N_1420);
or U2570 (N_2570,N_1286,N_1278);
and U2571 (N_2571,N_1929,N_2251);
nor U2572 (N_2572,N_1678,N_1461);
or U2573 (N_2573,N_2024,N_1260);
nor U2574 (N_2574,N_1374,N_1871);
nand U2575 (N_2575,N_1476,N_2178);
xnor U2576 (N_2576,N_1370,N_2204);
nor U2577 (N_2577,N_2058,N_2067);
nor U2578 (N_2578,N_2264,N_1301);
xnor U2579 (N_2579,N_1643,N_1323);
nor U2580 (N_2580,N_1873,N_1923);
or U2581 (N_2581,N_1501,N_1945);
or U2582 (N_2582,N_2196,N_1886);
xnor U2583 (N_2583,N_1656,N_1911);
or U2584 (N_2584,N_1750,N_1263);
nor U2585 (N_2585,N_1507,N_1469);
or U2586 (N_2586,N_1714,N_2334);
nand U2587 (N_2587,N_1774,N_1393);
or U2588 (N_2588,N_2084,N_1280);
nor U2589 (N_2589,N_1608,N_1671);
and U2590 (N_2590,N_2300,N_1454);
or U2591 (N_2591,N_2128,N_1969);
nor U2592 (N_2592,N_1653,N_2392);
xor U2593 (N_2593,N_2317,N_2248);
nor U2594 (N_2594,N_1857,N_1355);
xnor U2595 (N_2595,N_2055,N_1767);
or U2596 (N_2596,N_1955,N_1781);
nand U2597 (N_2597,N_1447,N_2013);
or U2598 (N_2598,N_1952,N_2327);
or U2599 (N_2599,N_1578,N_1320);
xnor U2600 (N_2600,N_1463,N_2114);
or U2601 (N_2601,N_1606,N_1456);
and U2602 (N_2602,N_1410,N_2223);
nor U2603 (N_2603,N_1602,N_1707);
nand U2604 (N_2604,N_1568,N_1589);
xnor U2605 (N_2605,N_1884,N_2349);
and U2606 (N_2606,N_1564,N_1529);
xnor U2607 (N_2607,N_2160,N_1704);
xor U2608 (N_2608,N_1803,N_1412);
nand U2609 (N_2609,N_2366,N_1930);
and U2610 (N_2610,N_2322,N_1865);
xor U2611 (N_2611,N_2117,N_2284);
nor U2612 (N_2612,N_1229,N_1487);
and U2613 (N_2613,N_1466,N_2098);
nor U2614 (N_2614,N_1383,N_1595);
and U2615 (N_2615,N_1368,N_1625);
or U2616 (N_2616,N_1626,N_1960);
or U2617 (N_2617,N_2070,N_1980);
and U2618 (N_2618,N_1636,N_2231);
or U2619 (N_2619,N_2143,N_1715);
nor U2620 (N_2620,N_1724,N_1822);
xnor U2621 (N_2621,N_2371,N_1770);
nor U2622 (N_2622,N_1893,N_1446);
xnor U2623 (N_2623,N_2103,N_2367);
or U2624 (N_2624,N_1359,N_1943);
nor U2625 (N_2625,N_1903,N_2056);
nand U2626 (N_2626,N_1494,N_2263);
and U2627 (N_2627,N_1591,N_1840);
nor U2628 (N_2628,N_1411,N_2060);
xor U2629 (N_2629,N_1246,N_1462);
or U2630 (N_2630,N_2053,N_1334);
or U2631 (N_2631,N_2017,N_1652);
or U2632 (N_2632,N_1207,N_1912);
or U2633 (N_2633,N_2225,N_1931);
nand U2634 (N_2634,N_1730,N_1240);
nand U2635 (N_2635,N_2238,N_1816);
nand U2636 (N_2636,N_2082,N_1213);
xnor U2637 (N_2637,N_1693,N_1789);
or U2638 (N_2638,N_1238,N_1598);
or U2639 (N_2639,N_2296,N_1218);
or U2640 (N_2640,N_1208,N_1216);
xor U2641 (N_2641,N_1802,N_1792);
xnor U2642 (N_2642,N_1504,N_2297);
xnor U2643 (N_2643,N_1579,N_1997);
nor U2644 (N_2644,N_1786,N_1206);
or U2645 (N_2645,N_1541,N_1706);
nor U2646 (N_2646,N_1772,N_2286);
xnor U2647 (N_2647,N_1933,N_1695);
nor U2648 (N_2648,N_1483,N_2360);
nand U2649 (N_2649,N_1799,N_1614);
and U2650 (N_2650,N_1722,N_2140);
or U2651 (N_2651,N_1881,N_1232);
nand U2652 (N_2652,N_1795,N_2279);
nand U2653 (N_2653,N_2110,N_2354);
and U2654 (N_2654,N_2377,N_2278);
nor U2655 (N_2655,N_2167,N_1719);
nor U2656 (N_2656,N_1771,N_2047);
and U2657 (N_2657,N_2230,N_2180);
or U2658 (N_2658,N_2381,N_2210);
nor U2659 (N_2659,N_1909,N_1269);
xnor U2660 (N_2660,N_1396,N_2383);
nand U2661 (N_2661,N_1502,N_2306);
nand U2662 (N_2662,N_2149,N_2193);
nand U2663 (N_2663,N_1690,N_1475);
and U2664 (N_2664,N_1545,N_1913);
nor U2665 (N_2665,N_1954,N_2331);
nand U2666 (N_2666,N_1588,N_1560);
xor U2667 (N_2667,N_1484,N_2171);
xor U2668 (N_2668,N_2012,N_1904);
nor U2669 (N_2669,N_1566,N_1932);
xor U2670 (N_2670,N_1737,N_2391);
nor U2671 (N_2671,N_2161,N_1859);
or U2672 (N_2672,N_1827,N_1892);
nand U2673 (N_2673,N_1649,N_1562);
xnor U2674 (N_2674,N_1276,N_2272);
or U2675 (N_2675,N_1556,N_1272);
and U2676 (N_2676,N_2163,N_1784);
and U2677 (N_2677,N_2232,N_1868);
nor U2678 (N_2678,N_1982,N_1837);
nand U2679 (N_2679,N_2086,N_1753);
and U2680 (N_2680,N_1398,N_1267);
xnor U2681 (N_2681,N_1680,N_1418);
xor U2682 (N_2682,N_1956,N_1988);
or U2683 (N_2683,N_1925,N_1807);
or U2684 (N_2684,N_2294,N_1677);
nand U2685 (N_2685,N_2301,N_1751);
or U2686 (N_2686,N_2069,N_1497);
nor U2687 (N_2687,N_1547,N_1241);
xor U2688 (N_2688,N_1977,N_1406);
xnor U2689 (N_2689,N_1646,N_2258);
nand U2690 (N_2690,N_1927,N_1312);
and U2691 (N_2691,N_1834,N_1721);
xnor U2692 (N_2692,N_1485,N_1303);
nand U2693 (N_2693,N_2057,N_1567);
nand U2694 (N_2694,N_1974,N_1838);
nor U2695 (N_2695,N_2266,N_1285);
xor U2696 (N_2696,N_2113,N_1399);
and U2697 (N_2697,N_2108,N_1314);
xnor U2698 (N_2698,N_2183,N_2177);
xnor U2699 (N_2699,N_2150,N_1522);
xor U2700 (N_2700,N_2050,N_1599);
and U2701 (N_2701,N_1756,N_1408);
nor U2702 (N_2702,N_1419,N_2252);
nor U2703 (N_2703,N_2388,N_2328);
or U2704 (N_2704,N_2151,N_2089);
nor U2705 (N_2705,N_2043,N_1407);
or U2706 (N_2706,N_1409,N_1936);
nor U2707 (N_2707,N_1629,N_1385);
nand U2708 (N_2708,N_1228,N_1265);
xor U2709 (N_2709,N_1512,N_2083);
nor U2710 (N_2710,N_2095,N_1503);
xor U2711 (N_2711,N_1345,N_2227);
or U2712 (N_2712,N_1448,N_2314);
nand U2713 (N_2713,N_1432,N_1274);
nor U2714 (N_2714,N_1759,N_1453);
or U2715 (N_2715,N_1700,N_1563);
nand U2716 (N_2716,N_1902,N_2093);
or U2717 (N_2717,N_2222,N_2166);
xor U2718 (N_2718,N_1382,N_1525);
xor U2719 (N_2719,N_1467,N_1394);
xor U2720 (N_2720,N_1470,N_1898);
and U2721 (N_2721,N_1800,N_2190);
or U2722 (N_2722,N_2330,N_1222);
xor U2723 (N_2723,N_2037,N_2112);
nand U2724 (N_2724,N_2329,N_1231);
or U2725 (N_2725,N_1268,N_2137);
nor U2726 (N_2726,N_1778,N_1555);
xnor U2727 (N_2727,N_2116,N_1402);
nor U2728 (N_2728,N_1679,N_1823);
nor U2729 (N_2729,N_1437,N_1604);
and U2730 (N_2730,N_2359,N_2021);
nand U2731 (N_2731,N_2348,N_2040);
and U2732 (N_2732,N_1210,N_1864);
xnor U2733 (N_2733,N_1729,N_2041);
or U2734 (N_2734,N_1685,N_1998);
and U2735 (N_2735,N_1252,N_1236);
nand U2736 (N_2736,N_1694,N_1318);
and U2737 (N_2737,N_2224,N_1585);
and U2738 (N_2738,N_2308,N_1710);
nand U2739 (N_2739,N_1339,N_1642);
nand U2740 (N_2740,N_1367,N_1429);
or U2741 (N_2741,N_1259,N_2246);
nand U2742 (N_2742,N_1537,N_2159);
xnor U2743 (N_2743,N_2393,N_1825);
or U2744 (N_2744,N_1379,N_1573);
or U2745 (N_2745,N_1203,N_2341);
nand U2746 (N_2746,N_2337,N_2398);
xor U2747 (N_2747,N_1482,N_2356);
xnor U2748 (N_2748,N_2122,N_1794);
nor U2749 (N_2749,N_1551,N_1491);
xor U2750 (N_2750,N_1922,N_1300);
nor U2751 (N_2751,N_1289,N_1951);
nand U2752 (N_2752,N_1401,N_2170);
and U2753 (N_2753,N_1317,N_1831);
or U2754 (N_2754,N_2174,N_1876);
xnor U2755 (N_2755,N_2350,N_1942);
nor U2756 (N_2756,N_1623,N_2380);
xor U2757 (N_2757,N_1985,N_2250);
nand U2758 (N_2758,N_1313,N_2335);
or U2759 (N_2759,N_2338,N_2061);
nand U2760 (N_2760,N_2022,N_1860);
or U2761 (N_2761,N_1874,N_1841);
nor U2762 (N_2762,N_2234,N_1360);
or U2763 (N_2763,N_2292,N_1908);
nand U2764 (N_2764,N_1742,N_1987);
and U2765 (N_2765,N_1761,N_1728);
xor U2766 (N_2766,N_2265,N_1935);
and U2767 (N_2767,N_2186,N_1284);
xnor U2768 (N_2768,N_2214,N_1224);
nand U2769 (N_2769,N_1324,N_2134);
nand U2770 (N_2770,N_1431,N_2243);
xor U2771 (N_2771,N_2185,N_2121);
or U2772 (N_2772,N_1330,N_2111);
nand U2773 (N_2773,N_1583,N_1699);
and U2774 (N_2774,N_2281,N_1391);
or U2775 (N_2775,N_2261,N_2293);
xor U2776 (N_2776,N_1880,N_2344);
or U2777 (N_2777,N_1958,N_2105);
nor U2778 (N_2778,N_1515,N_1277);
nand U2779 (N_2779,N_1283,N_1307);
and U2780 (N_2780,N_1275,N_1295);
nor U2781 (N_2781,N_1516,N_2000);
nand U2782 (N_2782,N_2201,N_1310);
and U2783 (N_2783,N_2323,N_2326);
nor U2784 (N_2784,N_2290,N_2020);
and U2785 (N_2785,N_1388,N_2228);
or U2786 (N_2786,N_1639,N_2085);
nor U2787 (N_2787,N_1239,N_2008);
xnor U2788 (N_2788,N_2221,N_1791);
xnor U2789 (N_2789,N_2318,N_1818);
xnor U2790 (N_2790,N_1308,N_2219);
nand U2791 (N_2791,N_2298,N_2375);
and U2792 (N_2792,N_2032,N_2065);
xor U2793 (N_2793,N_1309,N_1319);
and U2794 (N_2794,N_1248,N_1734);
and U2795 (N_2795,N_2249,N_2175);
and U2796 (N_2796,N_1743,N_2276);
nand U2797 (N_2797,N_2202,N_2319);
and U2798 (N_2798,N_1508,N_1666);
or U2799 (N_2799,N_1601,N_1587);
nand U2800 (N_2800,N_1242,N_1490);
nand U2801 (N_2801,N_1615,N_2059);
or U2802 (N_2802,N_1959,N_2036);
nor U2803 (N_2803,N_2169,N_1325);
nand U2804 (N_2804,N_1667,N_1612);
nor U2805 (N_2805,N_1243,N_2311);
xnor U2806 (N_2806,N_1481,N_1664);
nor U2807 (N_2807,N_1918,N_1928);
or U2808 (N_2808,N_1984,N_1220);
nor U2809 (N_2809,N_1531,N_2124);
or U2810 (N_2810,N_2245,N_1804);
xor U2811 (N_2811,N_2316,N_1801);
nand U2812 (N_2812,N_1686,N_1895);
nor U2813 (N_2813,N_1211,N_1991);
xnor U2814 (N_2814,N_2126,N_1441);
nor U2815 (N_2815,N_1620,N_1782);
and U2816 (N_2816,N_1748,N_1341);
nor U2817 (N_2817,N_2141,N_2158);
and U2818 (N_2818,N_1776,N_2299);
nand U2819 (N_2819,N_1254,N_1297);
nand U2820 (N_2820,N_1768,N_1689);
and U2821 (N_2821,N_2325,N_1343);
nand U2822 (N_2822,N_2220,N_1727);
xnor U2823 (N_2823,N_1251,N_1205);
xor U2824 (N_2824,N_1659,N_1294);
nand U2825 (N_2825,N_1509,N_1540);
or U2826 (N_2826,N_2304,N_2385);
or U2827 (N_2827,N_1661,N_2191);
or U2828 (N_2828,N_2255,N_2132);
or U2829 (N_2829,N_1731,N_1266);
xnor U2830 (N_2830,N_1814,N_1896);
xnor U2831 (N_2831,N_2372,N_1826);
and U2832 (N_2832,N_2034,N_1424);
nand U2833 (N_2833,N_1917,N_2039);
nor U2834 (N_2834,N_2295,N_1811);
or U2835 (N_2835,N_2355,N_2397);
nor U2836 (N_2836,N_1520,N_1296);
and U2837 (N_2837,N_1668,N_1226);
nand U2838 (N_2838,N_2148,N_1682);
nor U2839 (N_2839,N_1663,N_1854);
nand U2840 (N_2840,N_1237,N_1253);
nand U2841 (N_2841,N_1720,N_2240);
or U2842 (N_2842,N_2176,N_1375);
and U2843 (N_2843,N_1436,N_1331);
nand U2844 (N_2844,N_2119,N_1856);
nor U2845 (N_2845,N_1299,N_1858);
and U2846 (N_2846,N_1600,N_1915);
xor U2847 (N_2847,N_1650,N_1445);
or U2848 (N_2848,N_1245,N_2365);
nor U2849 (N_2849,N_2023,N_2305);
xnor U2850 (N_2850,N_1364,N_2203);
and U2851 (N_2851,N_2342,N_1660);
nor U2852 (N_2852,N_1291,N_2181);
and U2853 (N_2853,N_2362,N_2307);
xor U2854 (N_2854,N_1793,N_1247);
or U2855 (N_2855,N_1478,N_1934);
or U2856 (N_2856,N_1745,N_2192);
nand U2857 (N_2857,N_1861,N_2396);
nor U2858 (N_2858,N_1256,N_1900);
or U2859 (N_2859,N_1813,N_1395);
nor U2860 (N_2860,N_1505,N_2025);
nor U2861 (N_2861,N_2054,N_1381);
or U2862 (N_2862,N_1305,N_1455);
and U2863 (N_2863,N_1806,N_1530);
or U2864 (N_2864,N_1726,N_2198);
and U2865 (N_2865,N_2282,N_1866);
xnor U2866 (N_2866,N_1940,N_2092);
xnor U2867 (N_2867,N_2309,N_1924);
nand U2868 (N_2868,N_1775,N_2131);
or U2869 (N_2869,N_2071,N_1458);
or U2870 (N_2870,N_2073,N_2099);
xor U2871 (N_2871,N_1739,N_1603);
nor U2872 (N_2872,N_2087,N_1787);
and U2873 (N_2873,N_1316,N_1443);
and U2874 (N_2874,N_1565,N_1986);
and U2875 (N_2875,N_1996,N_1692);
or U2876 (N_2876,N_1628,N_1654);
nand U2877 (N_2877,N_2019,N_2115);
nor U2878 (N_2878,N_1670,N_1906);
or U2879 (N_2879,N_1712,N_2157);
nand U2880 (N_2880,N_1234,N_2357);
xor U2881 (N_2881,N_1964,N_1438);
nor U2882 (N_2882,N_1271,N_1572);
and U2883 (N_2883,N_1250,N_1590);
nand U2884 (N_2884,N_1797,N_1665);
nor U2885 (N_2885,N_1550,N_2049);
or U2886 (N_2886,N_2358,N_1392);
xor U2887 (N_2887,N_2361,N_1891);
and U2888 (N_2888,N_1645,N_2368);
xor U2889 (N_2889,N_2280,N_1703);
nor U2890 (N_2890,N_1835,N_2127);
or U2891 (N_2891,N_1879,N_1887);
or U2892 (N_2892,N_1255,N_1812);
nor U2893 (N_2893,N_2139,N_1662);
and U2894 (N_2894,N_2211,N_1451);
and U2895 (N_2895,N_1517,N_2241);
xor U2896 (N_2896,N_1899,N_1346);
or U2897 (N_2897,N_1967,N_1336);
xnor U2898 (N_2898,N_1582,N_1843);
nor U2899 (N_2899,N_1975,N_1400);
or U2900 (N_2900,N_2147,N_2168);
or U2901 (N_2901,N_1526,N_2273);
nand U2902 (N_2902,N_1611,N_1326);
xor U2903 (N_2903,N_1850,N_2135);
or U2904 (N_2904,N_2133,N_1460);
or U2905 (N_2905,N_1992,N_1828);
and U2906 (N_2906,N_1348,N_1489);
nand U2907 (N_2907,N_2271,N_2088);
nand U2908 (N_2908,N_2237,N_1479);
and U2909 (N_2909,N_2389,N_1444);
nand U2910 (N_2910,N_1452,N_1223);
xor U2911 (N_2911,N_1365,N_1477);
nand U2912 (N_2912,N_2102,N_2081);
or U2913 (N_2913,N_2018,N_2003);
xor U2914 (N_2914,N_1270,N_1644);
and U2915 (N_2915,N_1616,N_1672);
and U2916 (N_2916,N_2346,N_1919);
nand U2917 (N_2917,N_1363,N_2179);
and U2918 (N_2918,N_1543,N_2333);
xnor U2919 (N_2919,N_1493,N_2048);
nand U2920 (N_2920,N_1362,N_1535);
and U2921 (N_2921,N_1824,N_1434);
xnor U2922 (N_2922,N_1422,N_1377);
nor U2923 (N_2923,N_1397,N_2207);
nand U2924 (N_2924,N_1373,N_2384);
xor U2925 (N_2925,N_1920,N_1735);
and U2926 (N_2926,N_2033,N_1510);
or U2927 (N_2927,N_1449,N_2370);
nand U2928 (N_2928,N_2031,N_1885);
nand U2929 (N_2929,N_1338,N_2153);
or U2930 (N_2930,N_1669,N_2236);
or U2931 (N_2931,N_1597,N_1747);
and U2932 (N_2932,N_2146,N_1691);
or U2933 (N_2933,N_1527,N_1201);
nor U2934 (N_2934,N_1836,N_1329);
nand U2935 (N_2935,N_2212,N_1638);
or U2936 (N_2936,N_1421,N_1637);
or U2937 (N_2937,N_1905,N_2173);
nor U2938 (N_2938,N_1749,N_1333);
nand U2939 (N_2939,N_2343,N_2188);
nand U2940 (N_2940,N_1657,N_2259);
xor U2941 (N_2941,N_2100,N_1570);
nor U2942 (N_2942,N_2184,N_1687);
nor U2943 (N_2943,N_2364,N_1548);
xnor U2944 (N_2944,N_1593,N_1561);
nor U2945 (N_2945,N_2028,N_2312);
xnor U2946 (N_2946,N_1569,N_1574);
nor U2947 (N_2947,N_2130,N_1292);
and U2948 (N_2948,N_1760,N_1581);
and U2949 (N_2949,N_2038,N_2145);
or U2950 (N_2950,N_2332,N_1773);
xor U2951 (N_2951,N_1471,N_2072);
nand U2952 (N_2952,N_1435,N_1633);
nor U2953 (N_2953,N_1523,N_2016);
nor U2954 (N_2954,N_1732,N_2011);
and U2955 (N_2955,N_1882,N_1584);
and U2956 (N_2956,N_1741,N_2321);
xnor U2957 (N_2957,N_1340,N_2096);
and U2958 (N_2958,N_2205,N_1349);
and U2959 (N_2959,N_1273,N_1376);
or U2960 (N_2960,N_1851,N_1426);
xor U2961 (N_2961,N_1962,N_1744);
and U2962 (N_2962,N_2046,N_1225);
or U2963 (N_2963,N_2045,N_1702);
xor U2964 (N_2964,N_1415,N_1701);
and U2965 (N_2965,N_1725,N_2399);
nor U2966 (N_2966,N_1553,N_1474);
nand U2967 (N_2967,N_2267,N_1863);
or U2968 (N_2968,N_1758,N_1978);
or U2969 (N_2969,N_1946,N_2078);
nand U2970 (N_2970,N_1371,N_2340);
xnor U2971 (N_2971,N_1212,N_1796);
and U2972 (N_2972,N_2154,N_2339);
xor U2973 (N_2973,N_1790,N_2194);
or U2974 (N_2974,N_2044,N_1405);
nor U2975 (N_2975,N_1950,N_2068);
xor U2976 (N_2976,N_2256,N_1968);
xor U2977 (N_2977,N_2118,N_1521);
nor U2978 (N_2978,N_1440,N_1464);
or U2979 (N_2979,N_2123,N_2260);
and U2980 (N_2980,N_2386,N_2182);
or U2981 (N_2981,N_1351,N_1533);
or U2982 (N_2982,N_2002,N_2303);
and U2983 (N_2983,N_1852,N_2213);
xor U2984 (N_2984,N_2101,N_1833);
and U2985 (N_2985,N_1498,N_1264);
xnor U2986 (N_2986,N_1817,N_2336);
and U2987 (N_2987,N_1298,N_2288);
nor U2988 (N_2988,N_2206,N_1492);
and U2989 (N_2989,N_1698,N_1777);
nor U2990 (N_2990,N_2079,N_2014);
and U2991 (N_2991,N_1605,N_1627);
nor U2992 (N_2992,N_1423,N_1655);
nand U2993 (N_2993,N_1473,N_1342);
nand U2994 (N_2994,N_1219,N_2310);
and U2995 (N_2995,N_1675,N_1862);
or U2996 (N_2996,N_2302,N_2104);
and U2997 (N_2997,N_1433,N_2125);
and U2998 (N_2998,N_1281,N_1853);
and U2999 (N_2999,N_2283,N_2235);
and U3000 (N_3000,N_1763,N_2319);
xor U3001 (N_3001,N_2205,N_1835);
or U3002 (N_3002,N_1336,N_2234);
or U3003 (N_3003,N_1408,N_1533);
nor U3004 (N_3004,N_1749,N_2248);
or U3005 (N_3005,N_1830,N_1272);
xor U3006 (N_3006,N_2047,N_1961);
or U3007 (N_3007,N_1403,N_2005);
and U3008 (N_3008,N_1346,N_1670);
xor U3009 (N_3009,N_1558,N_2262);
nor U3010 (N_3010,N_2250,N_1240);
or U3011 (N_3011,N_1772,N_1350);
nand U3012 (N_3012,N_1676,N_2042);
and U3013 (N_3013,N_1914,N_2192);
or U3014 (N_3014,N_2007,N_1685);
nor U3015 (N_3015,N_1648,N_1627);
or U3016 (N_3016,N_2047,N_2086);
and U3017 (N_3017,N_2218,N_1888);
or U3018 (N_3018,N_2037,N_1492);
or U3019 (N_3019,N_1464,N_1597);
and U3020 (N_3020,N_2276,N_2061);
xor U3021 (N_3021,N_1304,N_2188);
nor U3022 (N_3022,N_2235,N_2359);
or U3023 (N_3023,N_1358,N_1286);
and U3024 (N_3024,N_1465,N_2061);
nand U3025 (N_3025,N_2077,N_2142);
or U3026 (N_3026,N_2187,N_1204);
xnor U3027 (N_3027,N_2212,N_2368);
nor U3028 (N_3028,N_1378,N_1739);
nor U3029 (N_3029,N_2145,N_2049);
or U3030 (N_3030,N_1926,N_2358);
and U3031 (N_3031,N_2192,N_2246);
nand U3032 (N_3032,N_2077,N_1289);
nor U3033 (N_3033,N_2113,N_1948);
nand U3034 (N_3034,N_2017,N_2184);
nand U3035 (N_3035,N_1579,N_1337);
nor U3036 (N_3036,N_2185,N_2343);
nand U3037 (N_3037,N_1530,N_2340);
xnor U3038 (N_3038,N_2103,N_1421);
or U3039 (N_3039,N_1637,N_1873);
or U3040 (N_3040,N_1711,N_2335);
or U3041 (N_3041,N_2313,N_1788);
xnor U3042 (N_3042,N_1959,N_2028);
or U3043 (N_3043,N_2301,N_1602);
nand U3044 (N_3044,N_2394,N_2194);
nand U3045 (N_3045,N_1554,N_1925);
xor U3046 (N_3046,N_1970,N_1722);
nand U3047 (N_3047,N_1269,N_1259);
xnor U3048 (N_3048,N_2073,N_1486);
or U3049 (N_3049,N_1237,N_1899);
xor U3050 (N_3050,N_1504,N_1981);
and U3051 (N_3051,N_1934,N_1395);
xor U3052 (N_3052,N_2042,N_2120);
nor U3053 (N_3053,N_2113,N_1367);
xor U3054 (N_3054,N_2173,N_1200);
nor U3055 (N_3055,N_1864,N_1986);
xnor U3056 (N_3056,N_2184,N_1290);
nand U3057 (N_3057,N_2109,N_1947);
xor U3058 (N_3058,N_2297,N_2331);
and U3059 (N_3059,N_2363,N_2190);
xnor U3060 (N_3060,N_1235,N_2114);
xor U3061 (N_3061,N_1535,N_1243);
nor U3062 (N_3062,N_1477,N_1756);
or U3063 (N_3063,N_1811,N_1899);
or U3064 (N_3064,N_1554,N_1386);
nor U3065 (N_3065,N_1986,N_1656);
xnor U3066 (N_3066,N_1321,N_2126);
nor U3067 (N_3067,N_2157,N_1850);
xor U3068 (N_3068,N_1335,N_1331);
nand U3069 (N_3069,N_2166,N_1407);
or U3070 (N_3070,N_1647,N_1691);
and U3071 (N_3071,N_1984,N_2182);
and U3072 (N_3072,N_2359,N_1734);
xor U3073 (N_3073,N_1638,N_1588);
nor U3074 (N_3074,N_2382,N_1288);
xor U3075 (N_3075,N_2231,N_1320);
nor U3076 (N_3076,N_2162,N_1549);
or U3077 (N_3077,N_1218,N_1560);
nor U3078 (N_3078,N_2314,N_1670);
and U3079 (N_3079,N_2075,N_1248);
or U3080 (N_3080,N_1527,N_1972);
and U3081 (N_3081,N_1886,N_2383);
and U3082 (N_3082,N_1939,N_1874);
nand U3083 (N_3083,N_1837,N_2079);
xor U3084 (N_3084,N_1707,N_1254);
nand U3085 (N_3085,N_1490,N_2074);
and U3086 (N_3086,N_1445,N_1828);
nand U3087 (N_3087,N_2282,N_2051);
nand U3088 (N_3088,N_2363,N_1815);
and U3089 (N_3089,N_1442,N_1806);
nor U3090 (N_3090,N_2360,N_1810);
xor U3091 (N_3091,N_1557,N_2358);
nor U3092 (N_3092,N_1470,N_2318);
or U3093 (N_3093,N_2218,N_2100);
or U3094 (N_3094,N_1416,N_1827);
nand U3095 (N_3095,N_2065,N_1284);
nor U3096 (N_3096,N_1618,N_1700);
nor U3097 (N_3097,N_1891,N_2067);
and U3098 (N_3098,N_1603,N_2114);
xor U3099 (N_3099,N_2168,N_1489);
and U3100 (N_3100,N_2088,N_1660);
and U3101 (N_3101,N_1754,N_1800);
nand U3102 (N_3102,N_1887,N_2198);
nor U3103 (N_3103,N_2240,N_1247);
nor U3104 (N_3104,N_1201,N_2075);
nand U3105 (N_3105,N_2295,N_1574);
and U3106 (N_3106,N_2017,N_1834);
and U3107 (N_3107,N_2240,N_1664);
xor U3108 (N_3108,N_1588,N_2281);
nand U3109 (N_3109,N_1994,N_2244);
nand U3110 (N_3110,N_1660,N_1690);
or U3111 (N_3111,N_2005,N_1204);
or U3112 (N_3112,N_2364,N_2344);
nor U3113 (N_3113,N_2354,N_1470);
or U3114 (N_3114,N_2271,N_1474);
xor U3115 (N_3115,N_1225,N_1971);
or U3116 (N_3116,N_2178,N_2191);
nor U3117 (N_3117,N_2376,N_2217);
xor U3118 (N_3118,N_2061,N_1200);
or U3119 (N_3119,N_2183,N_1797);
nor U3120 (N_3120,N_1215,N_1798);
nor U3121 (N_3121,N_1945,N_1638);
nand U3122 (N_3122,N_1302,N_1624);
nor U3123 (N_3123,N_2188,N_2375);
nand U3124 (N_3124,N_1980,N_1752);
or U3125 (N_3125,N_1276,N_1735);
nand U3126 (N_3126,N_1878,N_1665);
and U3127 (N_3127,N_2058,N_1710);
or U3128 (N_3128,N_1904,N_1854);
nor U3129 (N_3129,N_1978,N_2094);
xnor U3130 (N_3130,N_1873,N_2369);
nand U3131 (N_3131,N_2337,N_1606);
nor U3132 (N_3132,N_2249,N_1749);
nand U3133 (N_3133,N_2244,N_1446);
nand U3134 (N_3134,N_1727,N_1383);
nand U3135 (N_3135,N_1466,N_1981);
nor U3136 (N_3136,N_2157,N_1453);
nor U3137 (N_3137,N_1892,N_1778);
and U3138 (N_3138,N_1443,N_1820);
and U3139 (N_3139,N_1269,N_1454);
xor U3140 (N_3140,N_1576,N_1534);
nand U3141 (N_3141,N_1818,N_1504);
and U3142 (N_3142,N_1870,N_1640);
or U3143 (N_3143,N_1503,N_1372);
nor U3144 (N_3144,N_2279,N_1489);
nor U3145 (N_3145,N_1531,N_1793);
xor U3146 (N_3146,N_1778,N_1532);
or U3147 (N_3147,N_2016,N_2174);
or U3148 (N_3148,N_2247,N_1605);
and U3149 (N_3149,N_1514,N_2109);
xor U3150 (N_3150,N_2309,N_1926);
and U3151 (N_3151,N_1828,N_2326);
nand U3152 (N_3152,N_1563,N_1829);
nor U3153 (N_3153,N_1484,N_2313);
or U3154 (N_3154,N_1513,N_1580);
nor U3155 (N_3155,N_1543,N_1600);
nand U3156 (N_3156,N_1365,N_1413);
xor U3157 (N_3157,N_2300,N_2056);
nor U3158 (N_3158,N_1758,N_2232);
or U3159 (N_3159,N_2279,N_1625);
nor U3160 (N_3160,N_1790,N_1611);
and U3161 (N_3161,N_1715,N_1864);
nor U3162 (N_3162,N_1873,N_2072);
or U3163 (N_3163,N_1522,N_2015);
nand U3164 (N_3164,N_1648,N_2244);
and U3165 (N_3165,N_1802,N_1393);
nand U3166 (N_3166,N_2242,N_1541);
or U3167 (N_3167,N_1701,N_1202);
nor U3168 (N_3168,N_1611,N_2322);
or U3169 (N_3169,N_1827,N_2259);
nand U3170 (N_3170,N_1838,N_1975);
nor U3171 (N_3171,N_1949,N_2057);
and U3172 (N_3172,N_2013,N_1799);
and U3173 (N_3173,N_1768,N_1245);
nor U3174 (N_3174,N_1371,N_2182);
and U3175 (N_3175,N_2261,N_2129);
or U3176 (N_3176,N_1932,N_2396);
xor U3177 (N_3177,N_1288,N_1994);
nor U3178 (N_3178,N_1970,N_1435);
or U3179 (N_3179,N_2082,N_1841);
nand U3180 (N_3180,N_1587,N_1570);
xor U3181 (N_3181,N_2215,N_2182);
and U3182 (N_3182,N_2383,N_2161);
xnor U3183 (N_3183,N_1387,N_2065);
or U3184 (N_3184,N_2137,N_1542);
xor U3185 (N_3185,N_1900,N_1946);
nand U3186 (N_3186,N_2233,N_1813);
xor U3187 (N_3187,N_1616,N_1725);
xnor U3188 (N_3188,N_1839,N_2117);
or U3189 (N_3189,N_1658,N_1936);
xnor U3190 (N_3190,N_1226,N_2026);
or U3191 (N_3191,N_2001,N_2199);
xor U3192 (N_3192,N_2001,N_2216);
xnor U3193 (N_3193,N_1213,N_1570);
nor U3194 (N_3194,N_1227,N_1914);
nor U3195 (N_3195,N_2399,N_2051);
and U3196 (N_3196,N_2210,N_1236);
nor U3197 (N_3197,N_1441,N_1884);
nor U3198 (N_3198,N_1628,N_1975);
and U3199 (N_3199,N_2224,N_1314);
or U3200 (N_3200,N_2326,N_2089);
nor U3201 (N_3201,N_2362,N_2063);
nand U3202 (N_3202,N_1330,N_1956);
nand U3203 (N_3203,N_2080,N_1469);
xnor U3204 (N_3204,N_2357,N_1349);
nor U3205 (N_3205,N_2316,N_2037);
nand U3206 (N_3206,N_1523,N_1689);
nor U3207 (N_3207,N_2051,N_1947);
nor U3208 (N_3208,N_1724,N_1720);
or U3209 (N_3209,N_2218,N_2031);
or U3210 (N_3210,N_2083,N_1244);
nand U3211 (N_3211,N_1748,N_2330);
or U3212 (N_3212,N_1375,N_1667);
or U3213 (N_3213,N_1353,N_2043);
nor U3214 (N_3214,N_1682,N_1663);
or U3215 (N_3215,N_1420,N_2282);
nor U3216 (N_3216,N_1740,N_1985);
and U3217 (N_3217,N_1268,N_1552);
and U3218 (N_3218,N_1231,N_1855);
xor U3219 (N_3219,N_2066,N_2060);
xor U3220 (N_3220,N_2309,N_1846);
nand U3221 (N_3221,N_2108,N_1961);
or U3222 (N_3222,N_1982,N_2019);
nor U3223 (N_3223,N_1909,N_1469);
or U3224 (N_3224,N_1435,N_2235);
or U3225 (N_3225,N_1591,N_1582);
nand U3226 (N_3226,N_1751,N_2121);
nor U3227 (N_3227,N_1901,N_1895);
or U3228 (N_3228,N_1756,N_1939);
and U3229 (N_3229,N_1911,N_2233);
nand U3230 (N_3230,N_1551,N_2278);
nor U3231 (N_3231,N_1640,N_1892);
and U3232 (N_3232,N_1853,N_2106);
nand U3233 (N_3233,N_2394,N_2254);
or U3234 (N_3234,N_1556,N_1925);
or U3235 (N_3235,N_1585,N_1747);
or U3236 (N_3236,N_2072,N_2132);
nand U3237 (N_3237,N_1750,N_2196);
nand U3238 (N_3238,N_1885,N_2397);
nand U3239 (N_3239,N_1672,N_2066);
nand U3240 (N_3240,N_2003,N_2030);
nor U3241 (N_3241,N_1776,N_1449);
or U3242 (N_3242,N_1970,N_1774);
xor U3243 (N_3243,N_2147,N_2066);
nand U3244 (N_3244,N_1239,N_1590);
and U3245 (N_3245,N_1978,N_2233);
or U3246 (N_3246,N_1374,N_1665);
xor U3247 (N_3247,N_2242,N_1910);
nor U3248 (N_3248,N_1597,N_2288);
nand U3249 (N_3249,N_2039,N_1553);
nand U3250 (N_3250,N_1706,N_1552);
nand U3251 (N_3251,N_1988,N_1994);
nand U3252 (N_3252,N_2380,N_1358);
and U3253 (N_3253,N_2030,N_1236);
or U3254 (N_3254,N_1288,N_1506);
nor U3255 (N_3255,N_1807,N_2312);
and U3256 (N_3256,N_2032,N_1897);
nor U3257 (N_3257,N_2158,N_2188);
xnor U3258 (N_3258,N_1729,N_1599);
and U3259 (N_3259,N_1896,N_2053);
and U3260 (N_3260,N_1674,N_2387);
xor U3261 (N_3261,N_2163,N_1594);
nand U3262 (N_3262,N_1453,N_1451);
and U3263 (N_3263,N_1904,N_1740);
nand U3264 (N_3264,N_2117,N_2232);
xor U3265 (N_3265,N_1379,N_2390);
and U3266 (N_3266,N_1982,N_2160);
xor U3267 (N_3267,N_1755,N_2320);
or U3268 (N_3268,N_2367,N_1938);
or U3269 (N_3269,N_1629,N_1678);
xor U3270 (N_3270,N_1843,N_1498);
xor U3271 (N_3271,N_1890,N_1513);
nand U3272 (N_3272,N_1516,N_1622);
or U3273 (N_3273,N_1317,N_1898);
or U3274 (N_3274,N_1651,N_1601);
or U3275 (N_3275,N_2370,N_2169);
xnor U3276 (N_3276,N_1245,N_1786);
nor U3277 (N_3277,N_1717,N_2013);
and U3278 (N_3278,N_1248,N_2269);
or U3279 (N_3279,N_2227,N_1956);
and U3280 (N_3280,N_1966,N_1822);
or U3281 (N_3281,N_1369,N_1846);
and U3282 (N_3282,N_2124,N_1390);
xor U3283 (N_3283,N_2205,N_1485);
nor U3284 (N_3284,N_1260,N_1270);
xor U3285 (N_3285,N_1976,N_2277);
nor U3286 (N_3286,N_1644,N_2386);
or U3287 (N_3287,N_2134,N_2294);
nor U3288 (N_3288,N_1239,N_2340);
and U3289 (N_3289,N_1844,N_2293);
or U3290 (N_3290,N_1499,N_1853);
xnor U3291 (N_3291,N_2310,N_1721);
nand U3292 (N_3292,N_2376,N_1639);
xnor U3293 (N_3293,N_1680,N_2204);
and U3294 (N_3294,N_1546,N_1258);
nor U3295 (N_3295,N_2073,N_1758);
and U3296 (N_3296,N_2096,N_2087);
or U3297 (N_3297,N_1360,N_2080);
or U3298 (N_3298,N_1605,N_2317);
and U3299 (N_3299,N_2199,N_2363);
nand U3300 (N_3300,N_1722,N_1962);
nor U3301 (N_3301,N_1715,N_1549);
nor U3302 (N_3302,N_1972,N_2257);
xnor U3303 (N_3303,N_1272,N_2392);
or U3304 (N_3304,N_1414,N_2107);
xor U3305 (N_3305,N_1862,N_2160);
or U3306 (N_3306,N_1298,N_2304);
nand U3307 (N_3307,N_1689,N_1787);
and U3308 (N_3308,N_1776,N_2244);
or U3309 (N_3309,N_2121,N_1565);
nand U3310 (N_3310,N_1941,N_1262);
and U3311 (N_3311,N_1897,N_2243);
and U3312 (N_3312,N_2317,N_1367);
xor U3313 (N_3313,N_1897,N_1237);
xor U3314 (N_3314,N_2292,N_1494);
nor U3315 (N_3315,N_1808,N_1511);
or U3316 (N_3316,N_2160,N_1306);
or U3317 (N_3317,N_2233,N_2275);
nor U3318 (N_3318,N_2141,N_1782);
and U3319 (N_3319,N_2247,N_2324);
and U3320 (N_3320,N_2195,N_1922);
and U3321 (N_3321,N_1919,N_1250);
and U3322 (N_3322,N_1667,N_1387);
and U3323 (N_3323,N_1490,N_2395);
nand U3324 (N_3324,N_1203,N_2164);
or U3325 (N_3325,N_2306,N_1864);
xnor U3326 (N_3326,N_1412,N_2399);
xnor U3327 (N_3327,N_1664,N_2333);
or U3328 (N_3328,N_2085,N_2155);
or U3329 (N_3329,N_2048,N_2190);
nand U3330 (N_3330,N_1670,N_2108);
or U3331 (N_3331,N_1706,N_1368);
xor U3332 (N_3332,N_1462,N_1966);
and U3333 (N_3333,N_1659,N_1342);
or U3334 (N_3334,N_1960,N_1707);
xnor U3335 (N_3335,N_2238,N_1678);
nor U3336 (N_3336,N_1786,N_2070);
xnor U3337 (N_3337,N_1388,N_2143);
xnor U3338 (N_3338,N_1526,N_2141);
nor U3339 (N_3339,N_1280,N_2009);
xnor U3340 (N_3340,N_2091,N_1992);
nand U3341 (N_3341,N_2055,N_1232);
or U3342 (N_3342,N_1277,N_1809);
and U3343 (N_3343,N_1724,N_1988);
nand U3344 (N_3344,N_2080,N_2006);
nor U3345 (N_3345,N_1551,N_1513);
nor U3346 (N_3346,N_1646,N_2200);
or U3347 (N_3347,N_1400,N_1996);
nand U3348 (N_3348,N_1650,N_1732);
nand U3349 (N_3349,N_2184,N_1721);
or U3350 (N_3350,N_1378,N_1465);
nand U3351 (N_3351,N_2087,N_1279);
or U3352 (N_3352,N_2105,N_1495);
and U3353 (N_3353,N_1603,N_2189);
nand U3354 (N_3354,N_2032,N_1272);
xnor U3355 (N_3355,N_2369,N_1933);
or U3356 (N_3356,N_1341,N_2317);
nand U3357 (N_3357,N_1663,N_2328);
or U3358 (N_3358,N_1499,N_2389);
and U3359 (N_3359,N_1764,N_2313);
or U3360 (N_3360,N_1333,N_1543);
nor U3361 (N_3361,N_1851,N_1565);
xnor U3362 (N_3362,N_1244,N_1392);
nor U3363 (N_3363,N_1803,N_2012);
nand U3364 (N_3364,N_1873,N_1794);
nor U3365 (N_3365,N_2288,N_1972);
nor U3366 (N_3366,N_1709,N_1331);
nand U3367 (N_3367,N_2336,N_2203);
and U3368 (N_3368,N_1402,N_2307);
and U3369 (N_3369,N_1472,N_2036);
and U3370 (N_3370,N_2235,N_1401);
xor U3371 (N_3371,N_1637,N_2284);
nand U3372 (N_3372,N_1441,N_1606);
or U3373 (N_3373,N_1951,N_1358);
or U3374 (N_3374,N_1755,N_2044);
or U3375 (N_3375,N_2333,N_2225);
nor U3376 (N_3376,N_1842,N_1720);
and U3377 (N_3377,N_1438,N_1881);
nand U3378 (N_3378,N_1937,N_1997);
xnor U3379 (N_3379,N_1536,N_1676);
nand U3380 (N_3380,N_1721,N_1672);
or U3381 (N_3381,N_2003,N_1918);
and U3382 (N_3382,N_1381,N_1290);
xor U3383 (N_3383,N_1538,N_2010);
and U3384 (N_3384,N_2165,N_2177);
or U3385 (N_3385,N_1889,N_2314);
nand U3386 (N_3386,N_1529,N_1293);
nand U3387 (N_3387,N_1388,N_1211);
nand U3388 (N_3388,N_2040,N_1912);
nand U3389 (N_3389,N_2040,N_2199);
xor U3390 (N_3390,N_1499,N_1470);
xnor U3391 (N_3391,N_1282,N_2296);
and U3392 (N_3392,N_1480,N_1602);
and U3393 (N_3393,N_2017,N_2109);
or U3394 (N_3394,N_2059,N_1314);
or U3395 (N_3395,N_2323,N_1236);
xor U3396 (N_3396,N_2123,N_2075);
nor U3397 (N_3397,N_1334,N_1604);
nor U3398 (N_3398,N_1688,N_1444);
or U3399 (N_3399,N_2186,N_1425);
or U3400 (N_3400,N_2238,N_1985);
nand U3401 (N_3401,N_2127,N_2048);
nand U3402 (N_3402,N_1357,N_1741);
nor U3403 (N_3403,N_2026,N_2250);
nand U3404 (N_3404,N_2373,N_2287);
and U3405 (N_3405,N_2022,N_1810);
nand U3406 (N_3406,N_2039,N_2211);
nor U3407 (N_3407,N_1555,N_2346);
nand U3408 (N_3408,N_2000,N_1601);
nor U3409 (N_3409,N_1240,N_1938);
nor U3410 (N_3410,N_1243,N_2316);
nor U3411 (N_3411,N_2155,N_1324);
nand U3412 (N_3412,N_1926,N_1669);
nand U3413 (N_3413,N_1403,N_1586);
nor U3414 (N_3414,N_1521,N_2126);
and U3415 (N_3415,N_1791,N_2059);
nand U3416 (N_3416,N_1843,N_1378);
nand U3417 (N_3417,N_1758,N_2371);
nand U3418 (N_3418,N_1486,N_2370);
nor U3419 (N_3419,N_1560,N_1593);
xnor U3420 (N_3420,N_1210,N_1226);
nor U3421 (N_3421,N_2052,N_1959);
nor U3422 (N_3422,N_1637,N_2147);
nor U3423 (N_3423,N_1839,N_1375);
nand U3424 (N_3424,N_1328,N_1414);
and U3425 (N_3425,N_1267,N_2189);
nand U3426 (N_3426,N_1598,N_2323);
or U3427 (N_3427,N_1347,N_1610);
or U3428 (N_3428,N_2390,N_1635);
nor U3429 (N_3429,N_1781,N_1821);
xnor U3430 (N_3430,N_1854,N_2171);
and U3431 (N_3431,N_2233,N_1403);
nor U3432 (N_3432,N_1724,N_1209);
nand U3433 (N_3433,N_1819,N_1986);
and U3434 (N_3434,N_1264,N_1331);
xnor U3435 (N_3435,N_1346,N_1354);
nor U3436 (N_3436,N_1779,N_2068);
or U3437 (N_3437,N_1644,N_1236);
and U3438 (N_3438,N_1547,N_1632);
xnor U3439 (N_3439,N_1502,N_2056);
nor U3440 (N_3440,N_1347,N_1534);
or U3441 (N_3441,N_2016,N_2205);
or U3442 (N_3442,N_1866,N_2150);
nand U3443 (N_3443,N_1719,N_1679);
nand U3444 (N_3444,N_1985,N_1237);
nor U3445 (N_3445,N_2293,N_2086);
nor U3446 (N_3446,N_2335,N_1727);
nor U3447 (N_3447,N_1378,N_1433);
nand U3448 (N_3448,N_1734,N_1386);
and U3449 (N_3449,N_1900,N_1514);
nand U3450 (N_3450,N_2248,N_1920);
nor U3451 (N_3451,N_1521,N_2163);
nor U3452 (N_3452,N_1583,N_2045);
and U3453 (N_3453,N_1207,N_1994);
and U3454 (N_3454,N_2169,N_1945);
nand U3455 (N_3455,N_2085,N_1304);
and U3456 (N_3456,N_2323,N_1326);
and U3457 (N_3457,N_1274,N_1994);
and U3458 (N_3458,N_1987,N_1355);
xnor U3459 (N_3459,N_1499,N_1736);
xor U3460 (N_3460,N_2031,N_1937);
nand U3461 (N_3461,N_1431,N_2317);
nand U3462 (N_3462,N_2080,N_1818);
xor U3463 (N_3463,N_2013,N_1816);
xnor U3464 (N_3464,N_1815,N_1350);
nor U3465 (N_3465,N_1604,N_1914);
and U3466 (N_3466,N_2201,N_1470);
nor U3467 (N_3467,N_1889,N_1325);
nor U3468 (N_3468,N_1965,N_1536);
or U3469 (N_3469,N_1365,N_2348);
nand U3470 (N_3470,N_2168,N_1428);
nor U3471 (N_3471,N_1540,N_2113);
nor U3472 (N_3472,N_1967,N_2198);
xor U3473 (N_3473,N_1627,N_1746);
or U3474 (N_3474,N_1782,N_2324);
and U3475 (N_3475,N_1405,N_2140);
or U3476 (N_3476,N_1558,N_2029);
nor U3477 (N_3477,N_2249,N_2183);
nand U3478 (N_3478,N_2025,N_2174);
nor U3479 (N_3479,N_1753,N_1721);
nor U3480 (N_3480,N_1344,N_2045);
xnor U3481 (N_3481,N_2338,N_1474);
and U3482 (N_3482,N_2360,N_2323);
xor U3483 (N_3483,N_2034,N_1975);
nor U3484 (N_3484,N_1200,N_1903);
and U3485 (N_3485,N_2316,N_1222);
and U3486 (N_3486,N_2297,N_1619);
nor U3487 (N_3487,N_2348,N_1407);
nand U3488 (N_3488,N_1654,N_1263);
or U3489 (N_3489,N_2327,N_1233);
nor U3490 (N_3490,N_1892,N_1410);
nand U3491 (N_3491,N_2114,N_1257);
xor U3492 (N_3492,N_2159,N_2172);
nor U3493 (N_3493,N_2246,N_1923);
and U3494 (N_3494,N_2157,N_1949);
nor U3495 (N_3495,N_2255,N_2318);
xnor U3496 (N_3496,N_1785,N_1672);
or U3497 (N_3497,N_1301,N_1314);
nor U3498 (N_3498,N_1219,N_1285);
nand U3499 (N_3499,N_2097,N_1683);
and U3500 (N_3500,N_1480,N_1694);
or U3501 (N_3501,N_1585,N_1978);
and U3502 (N_3502,N_2323,N_1361);
or U3503 (N_3503,N_2157,N_1954);
xnor U3504 (N_3504,N_1814,N_1377);
or U3505 (N_3505,N_1996,N_1708);
nor U3506 (N_3506,N_1455,N_1311);
xnor U3507 (N_3507,N_1288,N_1977);
nor U3508 (N_3508,N_2092,N_2347);
or U3509 (N_3509,N_1593,N_1416);
or U3510 (N_3510,N_2142,N_2297);
or U3511 (N_3511,N_2166,N_1769);
and U3512 (N_3512,N_1370,N_1609);
nor U3513 (N_3513,N_1734,N_2287);
xnor U3514 (N_3514,N_2292,N_1313);
or U3515 (N_3515,N_1558,N_1871);
nand U3516 (N_3516,N_1653,N_2126);
and U3517 (N_3517,N_2280,N_2101);
or U3518 (N_3518,N_1360,N_1307);
xor U3519 (N_3519,N_1604,N_1711);
xnor U3520 (N_3520,N_1708,N_2056);
or U3521 (N_3521,N_1473,N_1515);
xnor U3522 (N_3522,N_1887,N_2035);
nand U3523 (N_3523,N_1796,N_1836);
nor U3524 (N_3524,N_2284,N_1458);
xnor U3525 (N_3525,N_1474,N_1795);
xnor U3526 (N_3526,N_1254,N_1362);
nand U3527 (N_3527,N_1964,N_1752);
nor U3528 (N_3528,N_1290,N_2333);
and U3529 (N_3529,N_2155,N_1472);
nand U3530 (N_3530,N_1245,N_1520);
or U3531 (N_3531,N_1751,N_1698);
xor U3532 (N_3532,N_1654,N_1939);
nand U3533 (N_3533,N_2281,N_1747);
nand U3534 (N_3534,N_1284,N_1202);
nor U3535 (N_3535,N_1353,N_1833);
and U3536 (N_3536,N_2268,N_1758);
nand U3537 (N_3537,N_1559,N_2267);
nand U3538 (N_3538,N_1878,N_2213);
nor U3539 (N_3539,N_1742,N_1682);
and U3540 (N_3540,N_2293,N_2148);
nand U3541 (N_3541,N_2349,N_1929);
and U3542 (N_3542,N_2207,N_2198);
nand U3543 (N_3543,N_1386,N_1757);
xor U3544 (N_3544,N_1417,N_2340);
or U3545 (N_3545,N_1630,N_2074);
xnor U3546 (N_3546,N_2137,N_1271);
nand U3547 (N_3547,N_1297,N_1609);
and U3548 (N_3548,N_1738,N_2031);
and U3549 (N_3549,N_1953,N_1985);
xor U3550 (N_3550,N_1954,N_1964);
and U3551 (N_3551,N_1264,N_1770);
and U3552 (N_3552,N_1976,N_1461);
or U3553 (N_3553,N_2269,N_2133);
nand U3554 (N_3554,N_1511,N_2393);
nand U3555 (N_3555,N_2103,N_1217);
nor U3556 (N_3556,N_2050,N_1567);
nor U3557 (N_3557,N_1864,N_1200);
xnor U3558 (N_3558,N_2326,N_1375);
xor U3559 (N_3559,N_1821,N_2005);
nand U3560 (N_3560,N_2147,N_1991);
nand U3561 (N_3561,N_2339,N_2200);
or U3562 (N_3562,N_1277,N_1833);
and U3563 (N_3563,N_1800,N_1487);
nand U3564 (N_3564,N_1283,N_1599);
nor U3565 (N_3565,N_2366,N_1787);
nor U3566 (N_3566,N_2067,N_1682);
nand U3567 (N_3567,N_1337,N_2278);
nor U3568 (N_3568,N_1703,N_1687);
nor U3569 (N_3569,N_1588,N_2229);
nand U3570 (N_3570,N_1282,N_1697);
or U3571 (N_3571,N_1290,N_1429);
nand U3572 (N_3572,N_2353,N_2061);
nor U3573 (N_3573,N_2210,N_2024);
xnor U3574 (N_3574,N_2042,N_2183);
and U3575 (N_3575,N_1316,N_1839);
xnor U3576 (N_3576,N_1393,N_1463);
xor U3577 (N_3577,N_1590,N_1538);
or U3578 (N_3578,N_2140,N_1544);
nor U3579 (N_3579,N_1205,N_1349);
xnor U3580 (N_3580,N_1384,N_1862);
nand U3581 (N_3581,N_1808,N_1984);
and U3582 (N_3582,N_1740,N_2039);
and U3583 (N_3583,N_1333,N_1275);
or U3584 (N_3584,N_2108,N_1618);
nand U3585 (N_3585,N_1588,N_1756);
and U3586 (N_3586,N_1760,N_1998);
nor U3587 (N_3587,N_1584,N_2267);
or U3588 (N_3588,N_1713,N_1850);
nand U3589 (N_3589,N_2179,N_1271);
nor U3590 (N_3590,N_1637,N_2026);
nor U3591 (N_3591,N_1401,N_2088);
nand U3592 (N_3592,N_2133,N_2252);
nor U3593 (N_3593,N_1958,N_2082);
nand U3594 (N_3594,N_1741,N_2129);
xnor U3595 (N_3595,N_2198,N_1593);
and U3596 (N_3596,N_1417,N_1729);
nand U3597 (N_3597,N_2339,N_2014);
xnor U3598 (N_3598,N_1320,N_2391);
nand U3599 (N_3599,N_1247,N_2339);
or U3600 (N_3600,N_2798,N_3443);
xor U3601 (N_3601,N_3496,N_3262);
nand U3602 (N_3602,N_2990,N_3371);
xnor U3603 (N_3603,N_3154,N_3438);
nor U3604 (N_3604,N_3072,N_2501);
nand U3605 (N_3605,N_3383,N_3089);
xnor U3606 (N_3606,N_3551,N_2760);
nand U3607 (N_3607,N_3189,N_3097);
or U3608 (N_3608,N_3400,N_3251);
or U3609 (N_3609,N_3593,N_3521);
or U3610 (N_3610,N_3208,N_2742);
nor U3611 (N_3611,N_2673,N_2869);
xnor U3612 (N_3612,N_3148,N_3158);
or U3613 (N_3613,N_3488,N_3197);
xnor U3614 (N_3614,N_3152,N_3556);
nor U3615 (N_3615,N_3076,N_2774);
nor U3616 (N_3616,N_3368,N_2485);
xnor U3617 (N_3617,N_3357,N_3324);
nand U3618 (N_3618,N_3566,N_3479);
nand U3619 (N_3619,N_3423,N_2462);
and U3620 (N_3620,N_2625,N_3242);
xor U3621 (N_3621,N_3114,N_3524);
xnor U3622 (N_3622,N_2484,N_2675);
nand U3623 (N_3623,N_3062,N_3414);
or U3624 (N_3624,N_2792,N_2426);
nand U3625 (N_3625,N_3468,N_3255);
and U3626 (N_3626,N_2514,N_3265);
nor U3627 (N_3627,N_3598,N_2498);
and U3628 (N_3628,N_2654,N_2558);
nand U3629 (N_3629,N_3023,N_3536);
and U3630 (N_3630,N_2456,N_3178);
and U3631 (N_3631,N_3007,N_3366);
and U3632 (N_3632,N_2735,N_2598);
and U3633 (N_3633,N_2607,N_3012);
and U3634 (N_3634,N_2809,N_2812);
nor U3635 (N_3635,N_2852,N_3204);
nor U3636 (N_3636,N_2833,N_3247);
or U3637 (N_3637,N_3014,N_3388);
and U3638 (N_3638,N_2860,N_2994);
nand U3639 (N_3639,N_3080,N_2545);
nor U3640 (N_3640,N_2828,N_3191);
or U3641 (N_3641,N_3353,N_3585);
and U3642 (N_3642,N_3293,N_3385);
and U3643 (N_3643,N_2508,N_2608);
xnor U3644 (N_3644,N_2422,N_2695);
or U3645 (N_3645,N_3042,N_3253);
and U3646 (N_3646,N_3106,N_2929);
nor U3647 (N_3647,N_3446,N_3452);
xnor U3648 (N_3648,N_3431,N_3006);
or U3649 (N_3649,N_3436,N_2521);
nor U3650 (N_3650,N_2820,N_2698);
nor U3651 (N_3651,N_3445,N_3442);
and U3652 (N_3652,N_2414,N_2824);
nor U3653 (N_3653,N_2899,N_2767);
xnor U3654 (N_3654,N_2663,N_3369);
or U3655 (N_3655,N_2472,N_3416);
or U3656 (N_3656,N_3312,N_2800);
xnor U3657 (N_3657,N_2517,N_3546);
or U3658 (N_3658,N_3290,N_2580);
or U3659 (N_3659,N_3430,N_3311);
or U3660 (N_3660,N_3003,N_2609);
or U3661 (N_3661,N_3028,N_2400);
or U3662 (N_3662,N_2822,N_3466);
xnor U3663 (N_3663,N_3061,N_2579);
or U3664 (N_3664,N_2979,N_2638);
and U3665 (N_3665,N_2814,N_2984);
or U3666 (N_3666,N_2684,N_2629);
xnor U3667 (N_3667,N_3509,N_3026);
nand U3668 (N_3668,N_3422,N_2887);
nand U3669 (N_3669,N_3338,N_3111);
xnor U3670 (N_3670,N_3088,N_2790);
nand U3671 (N_3671,N_2952,N_3354);
nand U3672 (N_3672,N_3087,N_3054);
xor U3673 (N_3673,N_2652,N_3459);
and U3674 (N_3674,N_2620,N_3230);
and U3675 (N_3675,N_2420,N_3515);
xnor U3676 (N_3676,N_2796,N_3548);
and U3677 (N_3677,N_2585,N_2593);
nand U3678 (N_3678,N_2779,N_3339);
nand U3679 (N_3679,N_3565,N_3123);
and U3680 (N_3680,N_2881,N_2572);
and U3681 (N_3681,N_3126,N_3395);
and U3682 (N_3682,N_2565,N_3108);
xor U3683 (N_3683,N_3561,N_3075);
xnor U3684 (N_3684,N_3011,N_3024);
xor U3685 (N_3685,N_2996,N_3182);
nand U3686 (N_3686,N_3522,N_3124);
nor U3687 (N_3687,N_3033,N_3199);
nand U3688 (N_3688,N_3306,N_3505);
nor U3689 (N_3689,N_2861,N_2591);
or U3690 (N_3690,N_3211,N_3579);
xnor U3691 (N_3691,N_2478,N_2702);
xor U3692 (N_3692,N_3508,N_2910);
nand U3693 (N_3693,N_2540,N_2449);
nor U3694 (N_3694,N_2440,N_2448);
and U3695 (N_3695,N_2885,N_2917);
nor U3696 (N_3696,N_2576,N_2537);
or U3697 (N_3697,N_2575,N_3387);
nand U3698 (N_3698,N_2407,N_2884);
xnor U3699 (N_3699,N_2592,N_2936);
nand U3700 (N_3700,N_3584,N_2908);
nor U3701 (N_3701,N_3346,N_3381);
or U3702 (N_3702,N_2965,N_2487);
nand U3703 (N_3703,N_2804,N_2436);
and U3704 (N_3704,N_3105,N_2795);
nand U3705 (N_3705,N_2443,N_2474);
nor U3706 (N_3706,N_2689,N_3065);
nand U3707 (N_3707,N_2639,N_2586);
nand U3708 (N_3708,N_2644,N_3577);
and U3709 (N_3709,N_3279,N_3491);
and U3710 (N_3710,N_3044,N_2883);
or U3711 (N_3711,N_2835,N_3470);
nor U3712 (N_3712,N_2787,N_3254);
nand U3713 (N_3713,N_3454,N_3038);
nand U3714 (N_3714,N_2534,N_2612);
nor U3715 (N_3715,N_3564,N_2811);
or U3716 (N_3716,N_2476,N_2511);
nor U3717 (N_3717,N_2909,N_2801);
or U3718 (N_3718,N_3529,N_3348);
nand U3719 (N_3719,N_2648,N_2749);
nor U3720 (N_3720,N_3037,N_2988);
nand U3721 (N_3721,N_3205,N_3483);
or U3722 (N_3722,N_3334,N_2458);
and U3723 (N_3723,N_2692,N_2481);
nor U3724 (N_3724,N_2865,N_2408);
xnor U3725 (N_3725,N_3081,N_2710);
xor U3726 (N_3726,N_2678,N_3147);
nor U3727 (N_3727,N_2816,N_2739);
xor U3728 (N_3728,N_3296,N_3035);
xor U3729 (N_3729,N_3399,N_3016);
or U3730 (N_3730,N_2997,N_3489);
or U3731 (N_3731,N_3153,N_3294);
xor U3732 (N_3732,N_2959,N_2913);
and U3733 (N_3733,N_2653,N_2621);
or U3734 (N_3734,N_2606,N_3250);
and U3735 (N_3735,N_2859,N_3025);
or U3736 (N_3736,N_2830,N_3288);
or U3737 (N_3737,N_3453,N_3228);
and U3738 (N_3738,N_3240,N_2759);
nand U3739 (N_3739,N_3372,N_3352);
nor U3740 (N_3740,N_2552,N_2890);
and U3741 (N_3741,N_2791,N_2601);
or U3742 (N_3742,N_2571,N_2748);
or U3743 (N_3743,N_3163,N_2687);
nand U3744 (N_3744,N_2978,N_3404);
nor U3745 (N_3745,N_2630,N_3527);
nand U3746 (N_3746,N_3307,N_3068);
or U3747 (N_3747,N_3428,N_2457);
or U3748 (N_3748,N_3193,N_2868);
and U3749 (N_3749,N_2752,N_2584);
or U3750 (N_3750,N_3020,N_2421);
or U3751 (N_3751,N_3592,N_2789);
or U3752 (N_3752,N_3393,N_2529);
or U3753 (N_3753,N_2533,N_3444);
or U3754 (N_3754,N_2793,N_3005);
and U3755 (N_3755,N_2943,N_3241);
nor U3756 (N_3756,N_3109,N_2506);
and U3757 (N_3757,N_2619,N_3289);
and U3758 (N_3758,N_3467,N_2488);
nor U3759 (N_3759,N_2982,N_3526);
or U3760 (N_3760,N_2966,N_2999);
nor U3761 (N_3761,N_2623,N_3375);
xnor U3762 (N_3762,N_3272,N_3258);
and U3763 (N_3763,N_3116,N_2761);
nor U3764 (N_3764,N_3560,N_3164);
or U3765 (N_3765,N_3341,N_2963);
xnor U3766 (N_3766,N_2751,N_2797);
and U3767 (N_3767,N_3233,N_3532);
nor U3768 (N_3768,N_2855,N_2465);
xnor U3769 (N_3769,N_2717,N_2613);
xnor U3770 (N_3770,N_2496,N_3408);
xnor U3771 (N_3771,N_2627,N_3046);
or U3772 (N_3772,N_2526,N_2803);
nor U3773 (N_3773,N_3326,N_3567);
and U3774 (N_3774,N_2986,N_2668);
and U3775 (N_3775,N_3209,N_2515);
xor U3776 (N_3776,N_3083,N_3215);
nor U3777 (N_3777,N_2546,N_3297);
nor U3778 (N_3778,N_3520,N_3538);
xor U3779 (N_3779,N_3224,N_3175);
or U3780 (N_3780,N_3058,N_3170);
nand U3781 (N_3781,N_2562,N_2723);
and U3782 (N_3782,N_3079,N_2681);
and U3783 (N_3783,N_2660,N_2412);
nand U3784 (N_3784,N_3122,N_3327);
nor U3785 (N_3785,N_2581,N_3409);
and U3786 (N_3786,N_2904,N_2956);
nand U3787 (N_3787,N_2479,N_3500);
nor U3788 (N_3788,N_3426,N_3207);
nor U3789 (N_3789,N_2903,N_2446);
xor U3790 (N_3790,N_2991,N_2856);
or U3791 (N_3791,N_2998,N_3367);
nand U3792 (N_3792,N_2772,N_3214);
nor U3793 (N_3793,N_2734,N_3319);
xor U3794 (N_3794,N_3476,N_2799);
xnor U3795 (N_3795,N_3583,N_3000);
or U3796 (N_3796,N_2777,N_3473);
or U3797 (N_3797,N_3402,N_3464);
or U3798 (N_3798,N_3516,N_2682);
nand U3799 (N_3799,N_3456,N_2905);
or U3800 (N_3800,N_2950,N_2507);
and U3801 (N_3801,N_3517,N_2520);
and U3802 (N_3802,N_3173,N_3051);
nor U3803 (N_3803,N_2649,N_2564);
or U3804 (N_3804,N_3130,N_3425);
nand U3805 (N_3805,N_2543,N_2719);
xor U3806 (N_3806,N_3528,N_3303);
and U3807 (N_3807,N_3474,N_3135);
nor U3808 (N_3808,N_2510,N_2722);
xnor U3809 (N_3809,N_3499,N_3273);
nor U3810 (N_3810,N_3301,N_3162);
xnor U3811 (N_3811,N_3386,N_2872);
nand U3812 (N_3812,N_2522,N_2403);
and U3813 (N_3813,N_2582,N_3047);
nor U3814 (N_3814,N_3142,N_3340);
or U3815 (N_3815,N_3523,N_2486);
and U3816 (N_3816,N_3413,N_3554);
xnor U3817 (N_3817,N_3321,N_2844);
xnor U3818 (N_3818,N_2753,N_3139);
or U3819 (N_3819,N_2504,N_2813);
xnor U3820 (N_3820,N_2926,N_2974);
xnor U3821 (N_3821,N_3156,N_3085);
and U3822 (N_3822,N_2785,N_3120);
or U3823 (N_3823,N_2490,N_3417);
nand U3824 (N_3824,N_2473,N_2976);
nor U3825 (N_3825,N_3384,N_2667);
or U3826 (N_3826,N_2938,N_3292);
nand U3827 (N_3827,N_2688,N_3314);
xnor U3828 (N_3828,N_2524,N_2875);
nor U3829 (N_3829,N_2771,N_3394);
xor U3830 (N_3830,N_2895,N_2736);
and U3831 (N_3831,N_3295,N_2831);
nor U3832 (N_3832,N_3008,N_2808);
nor U3833 (N_3833,N_3181,N_3355);
or U3834 (N_3834,N_3506,N_2461);
and U3835 (N_3835,N_3298,N_3485);
nand U3836 (N_3836,N_3271,N_3285);
and U3837 (N_3837,N_3392,N_2642);
nor U3838 (N_3838,N_3218,N_2437);
nor U3839 (N_3839,N_2445,N_3542);
nand U3840 (N_3840,N_3370,N_2631);
nand U3841 (N_3841,N_3107,N_3276);
xor U3842 (N_3842,N_2889,N_2658);
nor U3843 (N_3843,N_3418,N_3389);
or U3844 (N_3844,N_2964,N_3013);
and U3845 (N_3845,N_3433,N_3493);
nand U3846 (N_3846,N_2781,N_2829);
or U3847 (N_3847,N_3513,N_2637);
and U3848 (N_3848,N_3378,N_3531);
nor U3849 (N_3849,N_3235,N_3343);
or U3850 (N_3850,N_3451,N_3225);
or U3851 (N_3851,N_3084,N_2622);
xor U3852 (N_3852,N_3570,N_3465);
nor U3853 (N_3853,N_2746,N_2941);
and U3854 (N_3854,N_2706,N_2589);
or U3855 (N_3855,N_3057,N_3305);
or U3856 (N_3856,N_3447,N_3568);
xor U3857 (N_3857,N_2857,N_3210);
xnor U3858 (N_3858,N_2815,N_2876);
nand U3859 (N_3859,N_2893,N_3264);
xor U3860 (N_3860,N_3270,N_3141);
nor U3861 (N_3861,N_3283,N_2972);
nor U3862 (N_3862,N_3201,N_3450);
or U3863 (N_3863,N_3512,N_3421);
nand U3864 (N_3864,N_3091,N_2651);
nor U3865 (N_3865,N_3406,N_2786);
xor U3866 (N_3866,N_3086,N_3263);
nand U3867 (N_3867,N_3463,N_2776);
nor U3868 (N_3868,N_2993,N_3304);
or U3869 (N_3869,N_2834,N_2676);
nor U3870 (N_3870,N_2617,N_2728);
nand U3871 (N_3871,N_3501,N_3510);
nand U3872 (N_3872,N_2961,N_3015);
and U3873 (N_3873,N_3186,N_2674);
and U3874 (N_3874,N_3238,N_2432);
and U3875 (N_3875,N_3547,N_3177);
xor U3876 (N_3876,N_2823,N_3525);
nor U3877 (N_3877,N_2519,N_3236);
and U3878 (N_3878,N_2670,N_2764);
nand U3879 (N_3879,N_3535,N_2907);
xnor U3880 (N_3880,N_2467,N_3274);
and U3881 (N_3881,N_3115,N_2602);
nand U3882 (N_3882,N_2873,N_3458);
or U3883 (N_3883,N_3415,N_2902);
nor U3884 (N_3884,N_2453,N_3149);
nor U3885 (N_3885,N_2442,N_2699);
and U3886 (N_3886,N_2664,N_2704);
xor U3887 (N_3887,N_2709,N_2891);
nand U3888 (N_3888,N_3335,N_3071);
nor U3889 (N_3889,N_2531,N_2628);
or U3890 (N_3890,N_3492,N_3239);
and U3891 (N_3891,N_3138,N_2578);
xor U3892 (N_3892,N_3581,N_2817);
nand U3893 (N_3893,N_3027,N_2934);
nor U3894 (N_3894,N_3266,N_3403);
or U3895 (N_3895,N_2518,N_3518);
nand U3896 (N_3896,N_2957,N_3096);
nand U3897 (N_3897,N_2770,N_3101);
xor U3898 (N_3898,N_2845,N_2570);
xor U3899 (N_3899,N_2599,N_2928);
or U3900 (N_3900,N_2877,N_3259);
nand U3901 (N_3901,N_3481,N_2731);
or U3902 (N_3902,N_2842,N_2741);
nor U3903 (N_3903,N_2662,N_2724);
xnor U3904 (N_3904,N_3195,N_3471);
nor U3905 (N_3905,N_3377,N_3477);
nand U3906 (N_3906,N_2864,N_2583);
xnor U3907 (N_3907,N_3336,N_2766);
and U3908 (N_3908,N_3475,N_3132);
xor U3909 (N_3909,N_2512,N_3229);
or U3910 (N_3910,N_3498,N_2756);
and U3911 (N_3911,N_3318,N_3316);
nor U3912 (N_3912,N_3432,N_2509);
or U3913 (N_3913,N_2841,N_2794);
or U3914 (N_3914,N_2897,N_2683);
nor U3915 (N_3915,N_2549,N_2880);
xor U3916 (N_3916,N_2843,N_2464);
xnor U3917 (N_3917,N_3144,N_2419);
and U3918 (N_3918,N_2563,N_3202);
nand U3919 (N_3919,N_3179,N_2661);
and U3920 (N_3920,N_3519,N_3244);
and U3921 (N_3921,N_3494,N_2947);
nand U3922 (N_3922,N_2973,N_3364);
or U3923 (N_3923,N_2714,N_3420);
or U3924 (N_3924,N_2655,N_2497);
xnor U3925 (N_3925,N_3486,N_2825);
xnor U3926 (N_3926,N_3010,N_3009);
nand U3927 (N_3927,N_2666,N_3587);
or U3928 (N_3928,N_2680,N_3398);
or U3929 (N_3929,N_2945,N_2919);
nand U3930 (N_3930,N_3104,N_2755);
xor U3931 (N_3931,N_3143,N_3165);
and U3932 (N_3932,N_2922,N_2995);
nand U3933 (N_3933,N_2503,N_3249);
and U3934 (N_3934,N_3070,N_3441);
or U3935 (N_3935,N_3373,N_2541);
xnor U3936 (N_3936,N_2901,N_2451);
or U3937 (N_3937,N_3543,N_2677);
nor U3938 (N_3938,N_3039,N_2551);
and U3939 (N_3939,N_3300,N_3212);
and U3940 (N_3940,N_2747,N_3376);
or U3941 (N_3941,N_2611,N_3419);
nand U3942 (N_3942,N_3559,N_2685);
nor U3943 (N_3943,N_3308,N_2784);
nor U3944 (N_3944,N_2513,N_2523);
nor U3945 (N_3945,N_3462,N_2989);
nor U3946 (N_3946,N_2624,N_3030);
and U3947 (N_3947,N_3232,N_2435);
xor U3948 (N_3948,N_2836,N_2696);
and U3949 (N_3949,N_3150,N_2587);
nand U3950 (N_3950,N_2807,N_2444);
or U3951 (N_3951,N_3439,N_2559);
nand U3952 (N_3952,N_3576,N_2818);
nor U3953 (N_3953,N_2939,N_2441);
and U3954 (N_3954,N_3053,N_2650);
nor U3955 (N_3955,N_2775,N_3333);
xor U3956 (N_3956,N_2713,N_3050);
nor U3957 (N_3957,N_3129,N_3280);
nor U3958 (N_3958,N_2615,N_3045);
or U3959 (N_3959,N_2953,N_2433);
nor U3960 (N_3960,N_3365,N_3206);
nor U3961 (N_3961,N_3455,N_3216);
or U3962 (N_3962,N_3243,N_3379);
and U3963 (N_3963,N_2425,N_2635);
and U3964 (N_3964,N_3599,N_2935);
nor U3965 (N_3965,N_2577,N_3222);
nor U3966 (N_3966,N_3572,N_3449);
xnor U3967 (N_3967,N_3231,N_3220);
xor U3968 (N_3968,N_2733,N_2871);
or U3969 (N_3969,N_3102,N_2590);
or U3970 (N_3970,N_2574,N_2430);
or U3971 (N_3971,N_2505,N_3580);
or U3972 (N_3972,N_2940,N_2862);
and U3973 (N_3973,N_3256,N_2705);
or U3974 (N_3974,N_3017,N_2427);
xnor U3975 (N_3975,N_3268,N_3048);
and U3976 (N_3976,N_2553,N_3429);
or U3977 (N_3977,N_3412,N_2888);
or U3978 (N_3978,N_2700,N_3507);
or U3979 (N_3979,N_3582,N_3281);
and U3980 (N_3980,N_3261,N_3460);
and U3981 (N_3981,N_2482,N_3504);
or U3982 (N_3982,N_3069,N_2851);
xor U3983 (N_3983,N_2894,N_3555);
and U3984 (N_3984,N_2750,N_3345);
nand U3985 (N_3985,N_2404,N_3396);
nor U3986 (N_3986,N_3041,N_2914);
nand U3987 (N_3987,N_2434,N_2636);
or U3988 (N_3988,N_2532,N_3330);
and U3989 (N_3989,N_2566,N_2424);
or U3990 (N_3990,N_2968,N_2539);
and U3991 (N_3991,N_2886,N_3573);
xor U3992 (N_3992,N_3484,N_2805);
and U3993 (N_3993,N_2489,N_3029);
xnor U3994 (N_3994,N_3052,N_2827);
or U3995 (N_3995,N_3103,N_2931);
or U3996 (N_3996,N_2701,N_2491);
nor U3997 (N_3997,N_3134,N_2536);
nor U3998 (N_3998,N_3049,N_3284);
nand U3999 (N_3999,N_3131,N_3167);
nand U4000 (N_4000,N_2640,N_2874);
or U4001 (N_4001,N_2946,N_3176);
and U4002 (N_4002,N_2711,N_2405);
xnor U4003 (N_4003,N_2544,N_3502);
nand U4004 (N_4004,N_2921,N_2838);
nor U4005 (N_4005,N_3344,N_2900);
or U4006 (N_4006,N_2610,N_2821);
and U4007 (N_4007,N_2694,N_2431);
or U4008 (N_4008,N_3257,N_3128);
or U4009 (N_4009,N_3094,N_3213);
xnor U4010 (N_4010,N_3275,N_3155);
and U4011 (N_4011,N_2686,N_3064);
xor U4012 (N_4012,N_3363,N_2858);
xor U4013 (N_4013,N_2410,N_2826);
xor U4014 (N_4014,N_2768,N_3112);
nor U4015 (N_4015,N_2948,N_3328);
xor U4016 (N_4016,N_2460,N_3349);
xor U4017 (N_4017,N_3119,N_3350);
xor U4018 (N_4018,N_2542,N_3534);
nor U4019 (N_4019,N_3590,N_2415);
nor U4020 (N_4020,N_3185,N_3099);
xnor U4021 (N_4021,N_3480,N_3161);
and U4022 (N_4022,N_2530,N_2870);
nor U4023 (N_4023,N_3246,N_3411);
and U4024 (N_4024,N_3180,N_3435);
or U4025 (N_4025,N_2906,N_3067);
nand U4026 (N_4026,N_2614,N_2471);
nand U4027 (N_4027,N_2720,N_2715);
and U4028 (N_4028,N_2604,N_3332);
nor U4029 (N_4029,N_3427,N_3401);
nor U4030 (N_4030,N_3482,N_2616);
or U4031 (N_4031,N_3184,N_3077);
nand U4032 (N_4032,N_2960,N_3059);
or U4033 (N_4033,N_2712,N_3098);
or U4034 (N_4034,N_2454,N_3269);
nor U4035 (N_4035,N_2561,N_3034);
nor U4036 (N_4036,N_2892,N_2778);
nor U4037 (N_4037,N_2848,N_2573);
or U4038 (N_4038,N_3002,N_3503);
xor U4039 (N_4039,N_2878,N_2954);
xnor U4040 (N_4040,N_2925,N_3127);
or U4041 (N_4041,N_2762,N_2647);
and U4042 (N_4042,N_3495,N_2788);
xnor U4043 (N_4043,N_2810,N_2594);
nand U4044 (N_4044,N_2596,N_3313);
xnor U4045 (N_4045,N_2918,N_2665);
or U4046 (N_4046,N_2428,N_2763);
nand U4047 (N_4047,N_2516,N_2557);
nor U4048 (N_4048,N_2769,N_2927);
and U4049 (N_4049,N_2402,N_2896);
or U4050 (N_4050,N_3125,N_3074);
nand U4051 (N_4051,N_2937,N_3337);
nor U4052 (N_4052,N_3562,N_3198);
nand U4053 (N_4053,N_3021,N_3360);
nor U4054 (N_4054,N_2882,N_3157);
nand U4055 (N_4055,N_3168,N_2740);
and U4056 (N_4056,N_3248,N_3589);
or U4057 (N_4057,N_2757,N_2641);
xnor U4058 (N_4058,N_3252,N_2450);
xor U4059 (N_4059,N_3113,N_2477);
and U4060 (N_4060,N_2502,N_3032);
nor U4061 (N_4061,N_3457,N_2944);
xnor U4062 (N_4062,N_2981,N_3380);
or U4063 (N_4063,N_3056,N_3361);
xor U4064 (N_4064,N_3001,N_3171);
and U4065 (N_4065,N_2656,N_3203);
nand U4066 (N_4066,N_2932,N_3342);
and U4067 (N_4067,N_2765,N_2499);
nand U4068 (N_4068,N_2500,N_3036);
or U4069 (N_4069,N_2423,N_3558);
nor U4070 (N_4070,N_2949,N_2679);
or U4071 (N_4071,N_3018,N_3196);
or U4072 (N_4072,N_2560,N_2605);
and U4073 (N_4073,N_2725,N_3374);
nand U4074 (N_4074,N_2992,N_2847);
or U4075 (N_4075,N_3187,N_2550);
nor U4076 (N_4076,N_3060,N_3022);
or U4077 (N_4077,N_2463,N_3595);
xor U4078 (N_4078,N_3575,N_3390);
nor U4079 (N_4079,N_3424,N_3478);
nor U4080 (N_4080,N_3351,N_2853);
nor U4081 (N_4081,N_2554,N_3226);
or U4082 (N_4082,N_2690,N_3552);
and U4083 (N_4083,N_2406,N_3137);
or U4084 (N_4084,N_3286,N_2942);
nor U4085 (N_4085,N_3596,N_2923);
and U4086 (N_4086,N_3078,N_3530);
or U4087 (N_4087,N_2758,N_2951);
nor U4088 (N_4088,N_2911,N_2626);
or U4089 (N_4089,N_3391,N_2480);
nor U4090 (N_4090,N_3557,N_3121);
xnor U4091 (N_4091,N_2588,N_3092);
nand U4092 (N_4092,N_2975,N_2743);
nor U4093 (N_4093,N_3448,N_3310);
or U4094 (N_4094,N_3347,N_3299);
nor U4095 (N_4095,N_2691,N_2538);
nor U4096 (N_4096,N_3331,N_2737);
and U4097 (N_4097,N_2416,N_2567);
nand U4098 (N_4098,N_3472,N_3440);
xor U4099 (N_4099,N_3325,N_2738);
and U4100 (N_4100,N_3586,N_3317);
and U4101 (N_4101,N_2643,N_2915);
nand U4102 (N_4102,N_3063,N_2595);
nand U4103 (N_4103,N_2802,N_3591);
nand U4104 (N_4104,N_3574,N_3541);
xnor U4105 (N_4105,N_3329,N_3004);
and U4106 (N_4106,N_3140,N_2469);
or U4107 (N_4107,N_2971,N_2920);
and U4108 (N_4108,N_2879,N_2745);
and U4109 (N_4109,N_3260,N_3545);
or U4110 (N_4110,N_2840,N_2898);
and U4111 (N_4111,N_3183,N_2452);
nand U4112 (N_4112,N_2401,N_3497);
and U4113 (N_4113,N_2754,N_3055);
or U4114 (N_4114,N_3282,N_2555);
nand U4115 (N_4115,N_3594,N_3323);
or U4116 (N_4116,N_3302,N_2977);
xnor U4117 (N_4117,N_2849,N_2535);
nor U4118 (N_4118,N_3278,N_2730);
nor U4119 (N_4119,N_2547,N_2659);
or U4120 (N_4120,N_3553,N_3382);
nor U4121 (N_4121,N_2493,N_3227);
nand U4122 (N_4122,N_3159,N_3166);
nor U4123 (N_4123,N_2819,N_2568);
and U4124 (N_4124,N_2569,N_2707);
xnor U4125 (N_4125,N_3358,N_3405);
and U4126 (N_4126,N_3136,N_3194);
and U4127 (N_4127,N_3237,N_3550);
or U4128 (N_4128,N_2854,N_3192);
nor U4129 (N_4129,N_3200,N_3569);
nand U4130 (N_4130,N_2924,N_2438);
nor U4131 (N_4131,N_2867,N_2969);
nand U4132 (N_4132,N_3146,N_2744);
and U4133 (N_4133,N_3588,N_2773);
and U4134 (N_4134,N_2411,N_2556);
nand U4135 (N_4135,N_2470,N_3117);
xor U4136 (N_4136,N_3151,N_2603);
nor U4137 (N_4137,N_2409,N_3277);
xnor U4138 (N_4138,N_2703,N_3234);
or U4139 (N_4139,N_3217,N_3040);
and U4140 (N_4140,N_2447,N_2716);
xnor U4141 (N_4141,N_3043,N_2413);
or U4142 (N_4142,N_3571,N_3090);
nand U4143 (N_4143,N_2806,N_3287);
or U4144 (N_4144,N_3172,N_3533);
and U4145 (N_4145,N_3539,N_2930);
and U4146 (N_4146,N_2646,N_3190);
xnor U4147 (N_4147,N_2527,N_3461);
nand U4148 (N_4148,N_3145,N_3540);
nor U4149 (N_4149,N_2839,N_3514);
nand U4150 (N_4150,N_2863,N_2780);
or U4151 (N_4151,N_2468,N_2525);
and U4152 (N_4152,N_2429,N_2671);
or U4153 (N_4153,N_2912,N_3544);
nand U4154 (N_4154,N_3487,N_2618);
and U4155 (N_4155,N_3407,N_3309);
nand U4156 (N_4156,N_3093,N_2417);
xnor U4157 (N_4157,N_3578,N_2782);
and U4158 (N_4158,N_3095,N_2466);
or U4159 (N_4159,N_3073,N_3437);
nor U4160 (N_4160,N_3315,N_2832);
xor U4161 (N_4161,N_2727,N_3322);
nand U4162 (N_4162,N_2632,N_2933);
and U4163 (N_4163,N_3291,N_2528);
xor U4164 (N_4164,N_2726,N_3031);
nand U4165 (N_4165,N_2718,N_3133);
xor U4166 (N_4166,N_3469,N_3410);
and U4167 (N_4167,N_3219,N_2955);
nor U4168 (N_4168,N_2729,N_2657);
nand U4169 (N_4169,N_3019,N_3110);
nor U4170 (N_4170,N_2958,N_2721);
xor U4171 (N_4171,N_3223,N_2633);
nor U4172 (N_4172,N_2732,N_3490);
nand U4173 (N_4173,N_3174,N_2634);
xor U4174 (N_4174,N_2600,N_3100);
xnor U4175 (N_4175,N_3537,N_2494);
xnor U4176 (N_4176,N_2983,N_3188);
nor U4177 (N_4177,N_2783,N_3362);
or U4178 (N_4178,N_2970,N_3169);
nor U4179 (N_4179,N_3563,N_2495);
xnor U4180 (N_4180,N_2985,N_3320);
and U4181 (N_4181,N_3359,N_3356);
and U4182 (N_4182,N_2597,N_2455);
or U4183 (N_4183,N_3549,N_3082);
nor U4184 (N_4184,N_2987,N_3160);
or U4185 (N_4185,N_2846,N_3245);
nand U4186 (N_4186,N_2967,N_2645);
nor U4187 (N_4187,N_2669,N_3267);
nor U4188 (N_4188,N_3397,N_2916);
xor U4189 (N_4189,N_3434,N_3511);
nor U4190 (N_4190,N_2483,N_2850);
nor U4191 (N_4191,N_2672,N_3118);
nor U4192 (N_4192,N_2697,N_2439);
nor U4193 (N_4193,N_3221,N_3066);
or U4194 (N_4194,N_2492,N_2459);
or U4195 (N_4195,N_3597,N_2708);
and U4196 (N_4196,N_2980,N_2962);
xnor U4197 (N_4197,N_2837,N_2866);
or U4198 (N_4198,N_2475,N_2693);
nor U4199 (N_4199,N_2548,N_2418);
or U4200 (N_4200,N_3192,N_3066);
or U4201 (N_4201,N_2821,N_2856);
nand U4202 (N_4202,N_3478,N_3382);
xor U4203 (N_4203,N_3565,N_3185);
or U4204 (N_4204,N_2411,N_2788);
and U4205 (N_4205,N_3252,N_2538);
and U4206 (N_4206,N_2828,N_3533);
xor U4207 (N_4207,N_2567,N_2854);
or U4208 (N_4208,N_2842,N_2871);
or U4209 (N_4209,N_2907,N_3576);
and U4210 (N_4210,N_3508,N_3232);
and U4211 (N_4211,N_2803,N_3124);
and U4212 (N_4212,N_3050,N_3108);
nor U4213 (N_4213,N_3465,N_3308);
and U4214 (N_4214,N_2656,N_2691);
nor U4215 (N_4215,N_2414,N_3023);
or U4216 (N_4216,N_3011,N_3512);
nor U4217 (N_4217,N_3211,N_3561);
or U4218 (N_4218,N_2911,N_2716);
and U4219 (N_4219,N_3294,N_2995);
nand U4220 (N_4220,N_3297,N_2836);
or U4221 (N_4221,N_2739,N_3407);
nor U4222 (N_4222,N_2798,N_2468);
or U4223 (N_4223,N_3588,N_2701);
nand U4224 (N_4224,N_3483,N_3501);
xor U4225 (N_4225,N_2621,N_3400);
and U4226 (N_4226,N_2619,N_3164);
xnor U4227 (N_4227,N_2725,N_3361);
or U4228 (N_4228,N_3013,N_3340);
and U4229 (N_4229,N_3416,N_3190);
or U4230 (N_4230,N_3175,N_3284);
nor U4231 (N_4231,N_2626,N_3224);
nand U4232 (N_4232,N_3512,N_2803);
nor U4233 (N_4233,N_2768,N_2926);
xnor U4234 (N_4234,N_2507,N_3403);
or U4235 (N_4235,N_3273,N_3306);
nor U4236 (N_4236,N_2799,N_3270);
nor U4237 (N_4237,N_3588,N_2790);
and U4238 (N_4238,N_2515,N_2916);
xnor U4239 (N_4239,N_3029,N_3063);
xor U4240 (N_4240,N_3400,N_2730);
or U4241 (N_4241,N_2638,N_3014);
xor U4242 (N_4242,N_2813,N_2507);
nand U4243 (N_4243,N_3221,N_2486);
nor U4244 (N_4244,N_3367,N_3164);
nand U4245 (N_4245,N_3328,N_2756);
and U4246 (N_4246,N_3340,N_3471);
nor U4247 (N_4247,N_2535,N_3357);
or U4248 (N_4248,N_3459,N_2688);
nor U4249 (N_4249,N_3526,N_3349);
nand U4250 (N_4250,N_3557,N_2498);
nand U4251 (N_4251,N_3391,N_2562);
and U4252 (N_4252,N_3267,N_3422);
or U4253 (N_4253,N_3511,N_2914);
nand U4254 (N_4254,N_2494,N_3238);
nor U4255 (N_4255,N_2628,N_2826);
or U4256 (N_4256,N_3014,N_2609);
nand U4257 (N_4257,N_2506,N_3309);
nand U4258 (N_4258,N_3145,N_3281);
and U4259 (N_4259,N_3112,N_2520);
nand U4260 (N_4260,N_2542,N_3031);
xor U4261 (N_4261,N_2633,N_2867);
and U4262 (N_4262,N_2903,N_3251);
and U4263 (N_4263,N_3051,N_2868);
nor U4264 (N_4264,N_3540,N_3458);
xor U4265 (N_4265,N_2569,N_2551);
nor U4266 (N_4266,N_3528,N_2849);
nor U4267 (N_4267,N_3342,N_2963);
xnor U4268 (N_4268,N_3286,N_2435);
or U4269 (N_4269,N_2815,N_2968);
or U4270 (N_4270,N_3158,N_2891);
nor U4271 (N_4271,N_2801,N_2419);
nor U4272 (N_4272,N_2915,N_2817);
nor U4273 (N_4273,N_2788,N_3322);
xor U4274 (N_4274,N_3213,N_2629);
and U4275 (N_4275,N_3251,N_2987);
or U4276 (N_4276,N_3558,N_3369);
nand U4277 (N_4277,N_2791,N_3404);
nor U4278 (N_4278,N_2791,N_2531);
nor U4279 (N_4279,N_2767,N_3266);
nor U4280 (N_4280,N_3204,N_2877);
nand U4281 (N_4281,N_3169,N_2506);
nor U4282 (N_4282,N_3561,N_3220);
xor U4283 (N_4283,N_3414,N_3446);
nor U4284 (N_4284,N_3260,N_2409);
or U4285 (N_4285,N_2853,N_3059);
and U4286 (N_4286,N_2412,N_2432);
nor U4287 (N_4287,N_2699,N_2958);
nor U4288 (N_4288,N_3099,N_2632);
or U4289 (N_4289,N_2737,N_2645);
nor U4290 (N_4290,N_3596,N_3519);
xnor U4291 (N_4291,N_3325,N_2554);
xnor U4292 (N_4292,N_3508,N_3525);
or U4293 (N_4293,N_3051,N_3500);
and U4294 (N_4294,N_2840,N_2916);
nand U4295 (N_4295,N_2573,N_3562);
xor U4296 (N_4296,N_2964,N_3361);
or U4297 (N_4297,N_3479,N_3405);
nand U4298 (N_4298,N_3235,N_3303);
nand U4299 (N_4299,N_2969,N_3406);
and U4300 (N_4300,N_2749,N_2717);
nor U4301 (N_4301,N_2796,N_2898);
or U4302 (N_4302,N_2809,N_2659);
and U4303 (N_4303,N_2525,N_3131);
nand U4304 (N_4304,N_3188,N_2735);
xor U4305 (N_4305,N_2637,N_2613);
or U4306 (N_4306,N_3324,N_3599);
xor U4307 (N_4307,N_3537,N_2783);
nor U4308 (N_4308,N_3452,N_2783);
and U4309 (N_4309,N_2709,N_3043);
nand U4310 (N_4310,N_2464,N_3227);
nor U4311 (N_4311,N_2809,N_3341);
and U4312 (N_4312,N_2595,N_3005);
xnor U4313 (N_4313,N_3127,N_3020);
or U4314 (N_4314,N_3592,N_2606);
or U4315 (N_4315,N_3202,N_2452);
and U4316 (N_4316,N_3561,N_2961);
and U4317 (N_4317,N_3592,N_2410);
or U4318 (N_4318,N_2788,N_3269);
or U4319 (N_4319,N_3510,N_3132);
and U4320 (N_4320,N_2446,N_3498);
nor U4321 (N_4321,N_3533,N_3278);
or U4322 (N_4322,N_3542,N_3560);
nand U4323 (N_4323,N_3223,N_3228);
nor U4324 (N_4324,N_2573,N_2963);
xnor U4325 (N_4325,N_2567,N_2840);
nand U4326 (N_4326,N_3054,N_2858);
and U4327 (N_4327,N_2651,N_2873);
nor U4328 (N_4328,N_3018,N_3149);
or U4329 (N_4329,N_2977,N_3465);
xnor U4330 (N_4330,N_3092,N_3274);
and U4331 (N_4331,N_2937,N_3295);
xnor U4332 (N_4332,N_2667,N_3280);
xor U4333 (N_4333,N_2626,N_2656);
nand U4334 (N_4334,N_2661,N_3264);
nand U4335 (N_4335,N_2854,N_2958);
xnor U4336 (N_4336,N_2468,N_2943);
or U4337 (N_4337,N_3511,N_2450);
nand U4338 (N_4338,N_2957,N_2984);
xor U4339 (N_4339,N_2455,N_2702);
nand U4340 (N_4340,N_3471,N_2792);
or U4341 (N_4341,N_3097,N_2964);
xor U4342 (N_4342,N_2545,N_3346);
xor U4343 (N_4343,N_2425,N_2603);
or U4344 (N_4344,N_2496,N_3566);
nor U4345 (N_4345,N_3345,N_3463);
or U4346 (N_4346,N_2427,N_2692);
or U4347 (N_4347,N_3101,N_2657);
xnor U4348 (N_4348,N_2435,N_2466);
nand U4349 (N_4349,N_3205,N_2573);
nor U4350 (N_4350,N_2476,N_2520);
and U4351 (N_4351,N_3585,N_3139);
xor U4352 (N_4352,N_2921,N_2551);
nand U4353 (N_4353,N_3101,N_2852);
nand U4354 (N_4354,N_3107,N_3219);
or U4355 (N_4355,N_3441,N_2993);
xor U4356 (N_4356,N_2919,N_3315);
nor U4357 (N_4357,N_2525,N_3186);
or U4358 (N_4358,N_3032,N_2624);
or U4359 (N_4359,N_2702,N_2718);
nor U4360 (N_4360,N_3253,N_2842);
and U4361 (N_4361,N_2859,N_2635);
nor U4362 (N_4362,N_3375,N_2921);
or U4363 (N_4363,N_2611,N_3592);
nor U4364 (N_4364,N_2607,N_2691);
and U4365 (N_4365,N_2851,N_3586);
xor U4366 (N_4366,N_2680,N_2704);
or U4367 (N_4367,N_3124,N_3445);
nand U4368 (N_4368,N_3003,N_2794);
nor U4369 (N_4369,N_3389,N_3181);
or U4370 (N_4370,N_2500,N_3208);
nand U4371 (N_4371,N_2625,N_2527);
nor U4372 (N_4372,N_3110,N_3432);
xor U4373 (N_4373,N_2425,N_3100);
nand U4374 (N_4374,N_3210,N_2542);
and U4375 (N_4375,N_3562,N_2430);
nand U4376 (N_4376,N_3465,N_3409);
and U4377 (N_4377,N_2742,N_2875);
nor U4378 (N_4378,N_2855,N_3172);
or U4379 (N_4379,N_3239,N_3298);
or U4380 (N_4380,N_2533,N_3259);
or U4381 (N_4381,N_3199,N_3428);
nor U4382 (N_4382,N_2655,N_3358);
xor U4383 (N_4383,N_2865,N_3287);
xor U4384 (N_4384,N_3473,N_2874);
or U4385 (N_4385,N_2496,N_3060);
xnor U4386 (N_4386,N_2706,N_3331);
nand U4387 (N_4387,N_2899,N_2938);
or U4388 (N_4388,N_3346,N_3074);
or U4389 (N_4389,N_2637,N_3009);
nor U4390 (N_4390,N_3017,N_2661);
nand U4391 (N_4391,N_3157,N_2471);
nand U4392 (N_4392,N_2486,N_2627);
nor U4393 (N_4393,N_3533,N_2583);
or U4394 (N_4394,N_2688,N_3060);
nor U4395 (N_4395,N_3545,N_2585);
and U4396 (N_4396,N_3239,N_3165);
or U4397 (N_4397,N_2883,N_2937);
nor U4398 (N_4398,N_2559,N_2498);
and U4399 (N_4399,N_3438,N_3557);
and U4400 (N_4400,N_2871,N_3376);
xor U4401 (N_4401,N_2959,N_3511);
or U4402 (N_4402,N_3448,N_2675);
and U4403 (N_4403,N_2473,N_3168);
or U4404 (N_4404,N_2506,N_3399);
nor U4405 (N_4405,N_3336,N_2824);
nand U4406 (N_4406,N_2401,N_2429);
xnor U4407 (N_4407,N_2945,N_2586);
nand U4408 (N_4408,N_3071,N_3342);
nand U4409 (N_4409,N_2985,N_2504);
and U4410 (N_4410,N_3145,N_3432);
and U4411 (N_4411,N_2599,N_2977);
nor U4412 (N_4412,N_2586,N_2597);
nor U4413 (N_4413,N_2800,N_2643);
nor U4414 (N_4414,N_2672,N_2700);
nand U4415 (N_4415,N_3219,N_2577);
nand U4416 (N_4416,N_3559,N_2759);
and U4417 (N_4417,N_2632,N_3157);
nor U4418 (N_4418,N_3220,N_2470);
xor U4419 (N_4419,N_2582,N_3537);
or U4420 (N_4420,N_3160,N_2979);
nand U4421 (N_4421,N_2495,N_3260);
or U4422 (N_4422,N_2918,N_3216);
nand U4423 (N_4423,N_3116,N_2613);
or U4424 (N_4424,N_2422,N_3158);
or U4425 (N_4425,N_3187,N_3576);
xnor U4426 (N_4426,N_2669,N_3367);
and U4427 (N_4427,N_3020,N_2436);
and U4428 (N_4428,N_2843,N_3137);
and U4429 (N_4429,N_2722,N_2729);
xor U4430 (N_4430,N_3105,N_3325);
or U4431 (N_4431,N_2801,N_2510);
or U4432 (N_4432,N_3096,N_3042);
xor U4433 (N_4433,N_2997,N_3324);
nand U4434 (N_4434,N_2964,N_2811);
xor U4435 (N_4435,N_2675,N_3093);
xnor U4436 (N_4436,N_2876,N_2695);
nor U4437 (N_4437,N_3343,N_3040);
xor U4438 (N_4438,N_3472,N_3142);
nor U4439 (N_4439,N_2886,N_3001);
xor U4440 (N_4440,N_2580,N_2811);
or U4441 (N_4441,N_3501,N_3131);
or U4442 (N_4442,N_3200,N_3369);
nor U4443 (N_4443,N_2899,N_2657);
xnor U4444 (N_4444,N_3489,N_2482);
xor U4445 (N_4445,N_3159,N_2428);
and U4446 (N_4446,N_3035,N_3473);
nor U4447 (N_4447,N_2627,N_2728);
or U4448 (N_4448,N_2728,N_2858);
and U4449 (N_4449,N_3510,N_2584);
or U4450 (N_4450,N_2514,N_3486);
nand U4451 (N_4451,N_2905,N_3460);
or U4452 (N_4452,N_3132,N_2496);
nand U4453 (N_4453,N_3242,N_3574);
nand U4454 (N_4454,N_2789,N_2887);
or U4455 (N_4455,N_3035,N_3322);
and U4456 (N_4456,N_3255,N_2404);
or U4457 (N_4457,N_2695,N_2498);
nand U4458 (N_4458,N_2989,N_2592);
and U4459 (N_4459,N_3519,N_3065);
or U4460 (N_4460,N_3585,N_3281);
and U4461 (N_4461,N_3035,N_2404);
nor U4462 (N_4462,N_3579,N_3428);
nand U4463 (N_4463,N_2997,N_2434);
nor U4464 (N_4464,N_2970,N_3238);
or U4465 (N_4465,N_2452,N_3198);
xnor U4466 (N_4466,N_2444,N_2903);
or U4467 (N_4467,N_2912,N_3581);
xor U4468 (N_4468,N_3012,N_3370);
and U4469 (N_4469,N_2613,N_2777);
xnor U4470 (N_4470,N_3230,N_3267);
or U4471 (N_4471,N_2964,N_3321);
and U4472 (N_4472,N_2768,N_3380);
nand U4473 (N_4473,N_3503,N_3301);
or U4474 (N_4474,N_2442,N_3280);
or U4475 (N_4475,N_3366,N_3142);
xor U4476 (N_4476,N_2415,N_2742);
or U4477 (N_4477,N_3552,N_3542);
nand U4478 (N_4478,N_2492,N_2539);
nor U4479 (N_4479,N_2980,N_2981);
or U4480 (N_4480,N_3428,N_2439);
nand U4481 (N_4481,N_2501,N_2760);
nand U4482 (N_4482,N_2478,N_2773);
nand U4483 (N_4483,N_3305,N_2754);
xnor U4484 (N_4484,N_3019,N_2574);
xor U4485 (N_4485,N_3384,N_3048);
nand U4486 (N_4486,N_2863,N_2577);
xor U4487 (N_4487,N_2921,N_2641);
xnor U4488 (N_4488,N_2811,N_2570);
or U4489 (N_4489,N_2908,N_3439);
and U4490 (N_4490,N_2815,N_2447);
xnor U4491 (N_4491,N_3526,N_2670);
or U4492 (N_4492,N_3361,N_3059);
nand U4493 (N_4493,N_3174,N_3172);
nor U4494 (N_4494,N_2428,N_3027);
nand U4495 (N_4495,N_2563,N_2567);
nor U4496 (N_4496,N_3281,N_3334);
xnor U4497 (N_4497,N_3148,N_3457);
and U4498 (N_4498,N_3395,N_3462);
nor U4499 (N_4499,N_2962,N_2859);
and U4500 (N_4500,N_2772,N_2523);
nor U4501 (N_4501,N_3554,N_2753);
nand U4502 (N_4502,N_3195,N_3418);
or U4503 (N_4503,N_3435,N_2467);
xor U4504 (N_4504,N_2447,N_2632);
and U4505 (N_4505,N_2605,N_3184);
and U4506 (N_4506,N_2866,N_2425);
and U4507 (N_4507,N_3589,N_2705);
nand U4508 (N_4508,N_2980,N_2533);
and U4509 (N_4509,N_3580,N_2861);
and U4510 (N_4510,N_3446,N_2464);
xnor U4511 (N_4511,N_3300,N_2531);
nand U4512 (N_4512,N_2969,N_2614);
nor U4513 (N_4513,N_3236,N_3382);
nand U4514 (N_4514,N_3225,N_3251);
nor U4515 (N_4515,N_3290,N_2978);
xnor U4516 (N_4516,N_3280,N_3249);
or U4517 (N_4517,N_3423,N_2416);
or U4518 (N_4518,N_3366,N_2936);
xor U4519 (N_4519,N_3214,N_3137);
xnor U4520 (N_4520,N_2786,N_2582);
nand U4521 (N_4521,N_2708,N_2927);
and U4522 (N_4522,N_2731,N_3081);
nand U4523 (N_4523,N_2587,N_3394);
and U4524 (N_4524,N_3454,N_3042);
xor U4525 (N_4525,N_2966,N_2763);
nand U4526 (N_4526,N_3520,N_2779);
or U4527 (N_4527,N_3560,N_3275);
or U4528 (N_4528,N_2769,N_2519);
nor U4529 (N_4529,N_2438,N_3251);
or U4530 (N_4530,N_2452,N_2985);
and U4531 (N_4531,N_2778,N_3197);
or U4532 (N_4532,N_3439,N_2791);
and U4533 (N_4533,N_3518,N_3345);
or U4534 (N_4534,N_2568,N_3508);
xnor U4535 (N_4535,N_2759,N_3471);
xor U4536 (N_4536,N_2942,N_3420);
xnor U4537 (N_4537,N_3058,N_2461);
and U4538 (N_4538,N_2888,N_2804);
nor U4539 (N_4539,N_3560,N_2585);
nand U4540 (N_4540,N_3093,N_2916);
nor U4541 (N_4541,N_2666,N_2930);
nand U4542 (N_4542,N_2935,N_3146);
or U4543 (N_4543,N_3372,N_3073);
xnor U4544 (N_4544,N_2660,N_2447);
nor U4545 (N_4545,N_3044,N_3593);
nand U4546 (N_4546,N_2990,N_2778);
and U4547 (N_4547,N_2618,N_3452);
nor U4548 (N_4548,N_3130,N_2922);
nor U4549 (N_4549,N_2803,N_3368);
and U4550 (N_4550,N_2634,N_2631);
nor U4551 (N_4551,N_3564,N_3480);
or U4552 (N_4552,N_3030,N_2500);
nor U4553 (N_4553,N_3072,N_3205);
xnor U4554 (N_4554,N_2800,N_2582);
nand U4555 (N_4555,N_2518,N_2760);
or U4556 (N_4556,N_3171,N_3381);
or U4557 (N_4557,N_3506,N_3046);
or U4558 (N_4558,N_2792,N_2626);
or U4559 (N_4559,N_2423,N_3566);
nand U4560 (N_4560,N_2666,N_3254);
xnor U4561 (N_4561,N_2574,N_3582);
nor U4562 (N_4562,N_2572,N_2640);
xor U4563 (N_4563,N_2968,N_3166);
nor U4564 (N_4564,N_3592,N_2620);
xnor U4565 (N_4565,N_2594,N_3401);
or U4566 (N_4566,N_2409,N_2966);
nand U4567 (N_4567,N_2760,N_2831);
xor U4568 (N_4568,N_3275,N_2865);
nand U4569 (N_4569,N_2450,N_3094);
or U4570 (N_4570,N_3007,N_3551);
nand U4571 (N_4571,N_3484,N_2830);
or U4572 (N_4572,N_3432,N_2727);
nand U4573 (N_4573,N_2675,N_2746);
nor U4574 (N_4574,N_2608,N_3308);
or U4575 (N_4575,N_3381,N_2752);
and U4576 (N_4576,N_3583,N_2509);
or U4577 (N_4577,N_2658,N_2431);
and U4578 (N_4578,N_2570,N_3259);
and U4579 (N_4579,N_2774,N_3066);
or U4580 (N_4580,N_3105,N_2543);
nand U4581 (N_4581,N_2497,N_2677);
or U4582 (N_4582,N_2651,N_3254);
xnor U4583 (N_4583,N_3444,N_2951);
and U4584 (N_4584,N_3240,N_3500);
xnor U4585 (N_4585,N_2599,N_2727);
nor U4586 (N_4586,N_3134,N_3474);
or U4587 (N_4587,N_3405,N_2671);
and U4588 (N_4588,N_3447,N_2729);
nor U4589 (N_4589,N_2978,N_3527);
and U4590 (N_4590,N_3350,N_2926);
xor U4591 (N_4591,N_2825,N_3002);
xor U4592 (N_4592,N_2508,N_3367);
xor U4593 (N_4593,N_2477,N_2515);
or U4594 (N_4594,N_3227,N_3413);
xnor U4595 (N_4595,N_2475,N_3521);
and U4596 (N_4596,N_2784,N_2512);
nor U4597 (N_4597,N_2983,N_3117);
xor U4598 (N_4598,N_3581,N_3308);
xor U4599 (N_4599,N_3059,N_3223);
xor U4600 (N_4600,N_3550,N_3562);
or U4601 (N_4601,N_3291,N_3059);
nor U4602 (N_4602,N_2805,N_2826);
xnor U4603 (N_4603,N_2915,N_2627);
xnor U4604 (N_4604,N_2855,N_2762);
nand U4605 (N_4605,N_3033,N_2439);
or U4606 (N_4606,N_2554,N_2420);
xnor U4607 (N_4607,N_3532,N_2739);
nor U4608 (N_4608,N_3237,N_3542);
or U4609 (N_4609,N_2674,N_2862);
xor U4610 (N_4610,N_2767,N_3016);
nor U4611 (N_4611,N_3505,N_2562);
xor U4612 (N_4612,N_3114,N_3536);
nand U4613 (N_4613,N_3057,N_2791);
xor U4614 (N_4614,N_2897,N_3181);
nand U4615 (N_4615,N_3250,N_2737);
and U4616 (N_4616,N_2433,N_3324);
nor U4617 (N_4617,N_2616,N_2967);
or U4618 (N_4618,N_2622,N_2803);
and U4619 (N_4619,N_3377,N_2828);
nor U4620 (N_4620,N_2544,N_3558);
nor U4621 (N_4621,N_3299,N_2585);
or U4622 (N_4622,N_3321,N_2465);
and U4623 (N_4623,N_2556,N_3006);
or U4624 (N_4624,N_3171,N_3360);
xor U4625 (N_4625,N_2953,N_2971);
xnor U4626 (N_4626,N_2453,N_3168);
and U4627 (N_4627,N_3439,N_2534);
nor U4628 (N_4628,N_3480,N_2798);
and U4629 (N_4629,N_3217,N_2752);
and U4630 (N_4630,N_2572,N_2825);
xor U4631 (N_4631,N_3551,N_3173);
nand U4632 (N_4632,N_2726,N_2964);
or U4633 (N_4633,N_2531,N_2499);
and U4634 (N_4634,N_3028,N_3277);
xor U4635 (N_4635,N_3196,N_3560);
nand U4636 (N_4636,N_3165,N_2646);
or U4637 (N_4637,N_2669,N_3021);
nand U4638 (N_4638,N_2963,N_2755);
nor U4639 (N_4639,N_2562,N_2982);
and U4640 (N_4640,N_2836,N_2906);
or U4641 (N_4641,N_3019,N_3481);
and U4642 (N_4642,N_2701,N_3156);
or U4643 (N_4643,N_2411,N_2473);
and U4644 (N_4644,N_3193,N_3249);
nand U4645 (N_4645,N_3410,N_2464);
nand U4646 (N_4646,N_2943,N_2851);
nand U4647 (N_4647,N_3222,N_3346);
and U4648 (N_4648,N_2691,N_3253);
nand U4649 (N_4649,N_3128,N_2855);
or U4650 (N_4650,N_3438,N_2432);
and U4651 (N_4651,N_3059,N_3352);
nand U4652 (N_4652,N_3537,N_3357);
or U4653 (N_4653,N_3531,N_3212);
xnor U4654 (N_4654,N_2445,N_2917);
or U4655 (N_4655,N_3468,N_3360);
nand U4656 (N_4656,N_2751,N_2919);
nor U4657 (N_4657,N_3067,N_2497);
xnor U4658 (N_4658,N_2917,N_3597);
and U4659 (N_4659,N_2404,N_2750);
nor U4660 (N_4660,N_3514,N_2722);
or U4661 (N_4661,N_2774,N_2634);
nor U4662 (N_4662,N_2933,N_3044);
or U4663 (N_4663,N_3102,N_3586);
and U4664 (N_4664,N_2689,N_3584);
xor U4665 (N_4665,N_2536,N_3556);
xnor U4666 (N_4666,N_2974,N_3450);
and U4667 (N_4667,N_3269,N_2846);
or U4668 (N_4668,N_3252,N_3532);
xor U4669 (N_4669,N_2896,N_2974);
nor U4670 (N_4670,N_2509,N_3539);
and U4671 (N_4671,N_2781,N_3568);
nor U4672 (N_4672,N_2478,N_2608);
or U4673 (N_4673,N_3196,N_2621);
xor U4674 (N_4674,N_2501,N_2415);
nor U4675 (N_4675,N_3544,N_2489);
nor U4676 (N_4676,N_3300,N_2999);
nand U4677 (N_4677,N_3299,N_2402);
nand U4678 (N_4678,N_2833,N_3524);
xor U4679 (N_4679,N_3068,N_3351);
or U4680 (N_4680,N_3557,N_3151);
or U4681 (N_4681,N_3428,N_3333);
nor U4682 (N_4682,N_2455,N_3506);
xor U4683 (N_4683,N_3495,N_3218);
and U4684 (N_4684,N_3066,N_3298);
xnor U4685 (N_4685,N_3366,N_3511);
nor U4686 (N_4686,N_3477,N_3378);
xnor U4687 (N_4687,N_2636,N_3252);
nand U4688 (N_4688,N_2837,N_3482);
or U4689 (N_4689,N_2508,N_2414);
xnor U4690 (N_4690,N_3188,N_2937);
nor U4691 (N_4691,N_2720,N_2473);
xnor U4692 (N_4692,N_3573,N_2922);
or U4693 (N_4693,N_3124,N_2470);
or U4694 (N_4694,N_3553,N_3530);
nor U4695 (N_4695,N_2474,N_3175);
nand U4696 (N_4696,N_2806,N_2801);
nand U4697 (N_4697,N_3284,N_2915);
xnor U4698 (N_4698,N_2427,N_3503);
xnor U4699 (N_4699,N_2916,N_3230);
nor U4700 (N_4700,N_2720,N_3429);
and U4701 (N_4701,N_3347,N_3206);
or U4702 (N_4702,N_3370,N_3259);
or U4703 (N_4703,N_3494,N_3051);
nor U4704 (N_4704,N_3527,N_3337);
nand U4705 (N_4705,N_2483,N_3065);
nor U4706 (N_4706,N_3438,N_2727);
nand U4707 (N_4707,N_2458,N_3362);
and U4708 (N_4708,N_2554,N_2514);
nor U4709 (N_4709,N_3490,N_2916);
nand U4710 (N_4710,N_2442,N_3525);
and U4711 (N_4711,N_2786,N_2926);
nor U4712 (N_4712,N_3122,N_3415);
and U4713 (N_4713,N_3360,N_2698);
nor U4714 (N_4714,N_3544,N_2895);
xnor U4715 (N_4715,N_2841,N_2874);
nand U4716 (N_4716,N_2720,N_3551);
and U4717 (N_4717,N_2714,N_3565);
or U4718 (N_4718,N_3033,N_2577);
xor U4719 (N_4719,N_3053,N_2552);
or U4720 (N_4720,N_3251,N_3394);
and U4721 (N_4721,N_2887,N_3467);
xnor U4722 (N_4722,N_3423,N_3429);
nor U4723 (N_4723,N_3521,N_2675);
nor U4724 (N_4724,N_3205,N_3574);
nand U4725 (N_4725,N_3064,N_2651);
and U4726 (N_4726,N_2799,N_2977);
nor U4727 (N_4727,N_3438,N_2487);
or U4728 (N_4728,N_3332,N_3108);
and U4729 (N_4729,N_2606,N_3482);
or U4730 (N_4730,N_2635,N_2811);
nand U4731 (N_4731,N_2799,N_2454);
xnor U4732 (N_4732,N_2542,N_3014);
and U4733 (N_4733,N_3531,N_3559);
nor U4734 (N_4734,N_2524,N_3004);
or U4735 (N_4735,N_3237,N_3083);
nand U4736 (N_4736,N_3204,N_2991);
xor U4737 (N_4737,N_2628,N_2878);
xor U4738 (N_4738,N_3152,N_3203);
and U4739 (N_4739,N_3293,N_3432);
or U4740 (N_4740,N_2864,N_3432);
nor U4741 (N_4741,N_3319,N_3190);
or U4742 (N_4742,N_3131,N_2986);
nand U4743 (N_4743,N_3362,N_2680);
xnor U4744 (N_4744,N_3271,N_2834);
or U4745 (N_4745,N_3009,N_2901);
or U4746 (N_4746,N_2554,N_2593);
or U4747 (N_4747,N_3292,N_3027);
or U4748 (N_4748,N_3465,N_2705);
xor U4749 (N_4749,N_3022,N_2512);
or U4750 (N_4750,N_2682,N_2846);
and U4751 (N_4751,N_3079,N_2493);
xor U4752 (N_4752,N_3111,N_2461);
and U4753 (N_4753,N_3545,N_2779);
xor U4754 (N_4754,N_2826,N_3571);
or U4755 (N_4755,N_2600,N_2974);
or U4756 (N_4756,N_3129,N_2495);
nor U4757 (N_4757,N_2642,N_2514);
nor U4758 (N_4758,N_3311,N_2949);
nor U4759 (N_4759,N_3044,N_3179);
nor U4760 (N_4760,N_2923,N_2439);
nand U4761 (N_4761,N_3498,N_3097);
nor U4762 (N_4762,N_2970,N_3222);
nor U4763 (N_4763,N_3432,N_2648);
and U4764 (N_4764,N_3136,N_3389);
and U4765 (N_4765,N_2484,N_2570);
nor U4766 (N_4766,N_3414,N_2673);
nand U4767 (N_4767,N_2583,N_2905);
and U4768 (N_4768,N_2855,N_2997);
or U4769 (N_4769,N_3043,N_3544);
xor U4770 (N_4770,N_3097,N_2939);
or U4771 (N_4771,N_2642,N_3346);
or U4772 (N_4772,N_2448,N_2806);
or U4773 (N_4773,N_3361,N_2879);
or U4774 (N_4774,N_3130,N_3550);
xnor U4775 (N_4775,N_3051,N_2542);
nand U4776 (N_4776,N_2519,N_3547);
xnor U4777 (N_4777,N_2638,N_2604);
and U4778 (N_4778,N_3292,N_2425);
xnor U4779 (N_4779,N_3189,N_3568);
xnor U4780 (N_4780,N_3114,N_2417);
xor U4781 (N_4781,N_3165,N_2881);
or U4782 (N_4782,N_3382,N_2681);
and U4783 (N_4783,N_2408,N_3266);
nor U4784 (N_4784,N_2935,N_3388);
and U4785 (N_4785,N_2471,N_2401);
nand U4786 (N_4786,N_3364,N_2765);
nor U4787 (N_4787,N_2821,N_2625);
nor U4788 (N_4788,N_3292,N_2491);
xor U4789 (N_4789,N_3288,N_3209);
nor U4790 (N_4790,N_2917,N_3056);
and U4791 (N_4791,N_2749,N_2689);
nor U4792 (N_4792,N_2751,N_2997);
xnor U4793 (N_4793,N_3558,N_2918);
nor U4794 (N_4794,N_3239,N_2832);
nor U4795 (N_4795,N_3116,N_3213);
nor U4796 (N_4796,N_2802,N_2457);
and U4797 (N_4797,N_3108,N_2521);
nor U4798 (N_4798,N_3537,N_2817);
nor U4799 (N_4799,N_2891,N_3025);
xnor U4800 (N_4800,N_4493,N_4384);
and U4801 (N_4801,N_4551,N_4269);
nor U4802 (N_4802,N_4211,N_3754);
nand U4803 (N_4803,N_4739,N_3824);
nor U4804 (N_4804,N_3631,N_4499);
and U4805 (N_4805,N_3760,N_4520);
nor U4806 (N_4806,N_4653,N_4346);
nand U4807 (N_4807,N_4528,N_3625);
xnor U4808 (N_4808,N_4021,N_4446);
nor U4809 (N_4809,N_4102,N_4050);
and U4810 (N_4810,N_3646,N_4176);
xnor U4811 (N_4811,N_4659,N_3710);
nand U4812 (N_4812,N_4198,N_4578);
nand U4813 (N_4813,N_4027,N_3826);
nand U4814 (N_4814,N_3698,N_4227);
and U4815 (N_4815,N_3932,N_4416);
and U4816 (N_4816,N_3645,N_4015);
and U4817 (N_4817,N_3683,N_4078);
nand U4818 (N_4818,N_3636,N_4676);
nor U4819 (N_4819,N_4611,N_4468);
or U4820 (N_4820,N_4241,N_3835);
nand U4821 (N_4821,N_3753,N_3756);
xnor U4822 (N_4822,N_4434,N_3933);
nor U4823 (N_4823,N_4329,N_3984);
and U4824 (N_4824,N_4637,N_3612);
or U4825 (N_4825,N_4393,N_4461);
nand U4826 (N_4826,N_4340,N_4438);
nand U4827 (N_4827,N_4106,N_3627);
nand U4828 (N_4828,N_3998,N_4151);
nor U4829 (N_4829,N_4013,N_4402);
nor U4830 (N_4830,N_4382,N_4691);
nand U4831 (N_4831,N_3650,N_4391);
and U4832 (N_4832,N_4354,N_4268);
or U4833 (N_4833,N_4724,N_4479);
or U4834 (N_4834,N_3907,N_4463);
nand U4835 (N_4835,N_4649,N_4206);
nor U4836 (N_4836,N_4255,N_4126);
or U4837 (N_4837,N_4511,N_3622);
or U4838 (N_4838,N_4359,N_3891);
and U4839 (N_4839,N_4322,N_4726);
nor U4840 (N_4840,N_4639,N_4732);
nand U4841 (N_4841,N_4287,N_3973);
nand U4842 (N_4842,N_4593,N_4117);
nand U4843 (N_4843,N_3679,N_4740);
or U4844 (N_4844,N_3742,N_3670);
nor U4845 (N_4845,N_3740,N_3665);
and U4846 (N_4846,N_4041,N_4586);
nand U4847 (N_4847,N_4118,N_4383);
or U4848 (N_4848,N_3703,N_4708);
nand U4849 (N_4849,N_3803,N_3883);
xor U4850 (N_4850,N_4299,N_4624);
xnor U4851 (N_4851,N_3879,N_4533);
nor U4852 (N_4852,N_3800,N_4335);
nand U4853 (N_4853,N_4096,N_3709);
and U4854 (N_4854,N_4303,N_4609);
nand U4855 (N_4855,N_4664,N_4376);
nor U4856 (N_4856,N_4552,N_4454);
or U4857 (N_4857,N_3989,N_3987);
xnor U4858 (N_4858,N_4772,N_3841);
or U4859 (N_4859,N_3900,N_3678);
nand U4860 (N_4860,N_4143,N_4453);
xor U4861 (N_4861,N_4768,N_3635);
nor U4862 (N_4862,N_4625,N_4773);
and U4863 (N_4863,N_4066,N_3745);
and U4864 (N_4864,N_3818,N_4355);
or U4865 (N_4865,N_3948,N_3822);
nand U4866 (N_4866,N_4407,N_4471);
or U4867 (N_4867,N_3970,N_4228);
and U4868 (N_4868,N_3831,N_4422);
and U4869 (N_4869,N_4068,N_3674);
nor U4870 (N_4870,N_4314,N_4091);
xnor U4871 (N_4871,N_4719,N_3769);
nand U4872 (N_4872,N_3963,N_3807);
nor U4873 (N_4873,N_4642,N_3603);
or U4874 (N_4874,N_4425,N_4460);
or U4875 (N_4875,N_3974,N_4543);
nor U4876 (N_4876,N_4202,N_4309);
nand U4877 (N_4877,N_3884,N_3766);
nor U4878 (N_4878,N_3639,N_4364);
xor U4879 (N_4879,N_4709,N_3901);
or U4880 (N_4880,N_4785,N_3910);
xor U4881 (N_4881,N_3906,N_4620);
nand U4882 (N_4882,N_3787,N_4432);
and U4883 (N_4883,N_3684,N_4689);
nor U4884 (N_4884,N_4778,N_4009);
or U4885 (N_4885,N_4283,N_3934);
nor U4886 (N_4886,N_4686,N_4790);
and U4887 (N_4887,N_4403,N_4232);
nand U4888 (N_4888,N_3702,N_4475);
nor U4889 (N_4889,N_4555,N_4678);
and U4890 (N_4890,N_4690,N_3776);
xnor U4891 (N_4891,N_4749,N_4270);
xnor U4892 (N_4892,N_4224,N_4107);
or U4893 (N_4893,N_4782,N_4500);
or U4894 (N_4894,N_4447,N_4163);
nand U4895 (N_4895,N_3930,N_4249);
nand U4896 (N_4896,N_4683,N_4288);
or U4897 (N_4897,N_3726,N_3735);
and U4898 (N_4898,N_3793,N_4246);
and U4899 (N_4899,N_3915,N_4680);
xnor U4900 (N_4900,N_4750,N_3669);
nand U4901 (N_4901,N_4504,N_4065);
and U4902 (N_4902,N_4563,N_4131);
nand U4903 (N_4903,N_3940,N_4165);
or U4904 (N_4904,N_4099,N_4650);
xnor U4905 (N_4905,N_4527,N_3700);
nand U4906 (N_4906,N_4641,N_3997);
nand U4907 (N_4907,N_4644,N_3777);
or U4908 (N_4908,N_4368,N_4345);
or U4909 (N_4909,N_3617,N_4567);
nand U4910 (N_4910,N_4149,N_4305);
and U4911 (N_4911,N_4161,N_3959);
nor U4912 (N_4912,N_4164,N_4765);
nor U4913 (N_4913,N_4569,N_4497);
xor U4914 (N_4914,N_3782,N_4146);
nor U4915 (N_4915,N_4058,N_3601);
xor U4916 (N_4916,N_4754,N_3882);
or U4917 (N_4917,N_3964,N_3925);
and U4918 (N_4918,N_4697,N_3943);
and U4919 (N_4919,N_4579,N_4047);
nand U4920 (N_4920,N_3768,N_4252);
or U4921 (N_4921,N_3652,N_3994);
nor U4922 (N_4922,N_4159,N_3842);
nand U4923 (N_4923,N_4536,N_3648);
nor U4924 (N_4924,N_3770,N_3844);
or U4925 (N_4925,N_3764,N_4109);
and U4926 (N_4926,N_3881,N_4054);
or U4927 (N_4927,N_4408,N_4591);
or U4928 (N_4928,N_4170,N_4011);
or U4929 (N_4929,N_3653,N_3607);
or U4930 (N_4930,N_4052,N_4059);
xor U4931 (N_4931,N_4328,N_4127);
xnor U4932 (N_4932,N_4764,N_4597);
xnor U4933 (N_4933,N_4787,N_3682);
xnor U4934 (N_4934,N_4240,N_4779);
xor U4935 (N_4935,N_4729,N_4489);
nand U4936 (N_4936,N_3641,N_3672);
nand U4937 (N_4937,N_4038,N_4236);
nor U4938 (N_4938,N_4519,N_3899);
xor U4939 (N_4939,N_3729,N_4061);
or U4940 (N_4940,N_4745,N_4783);
nand U4941 (N_4941,N_3725,N_4512);
xnor U4942 (N_4942,N_4501,N_4072);
xor U4943 (N_4943,N_4646,N_4713);
xnor U4944 (N_4944,N_3849,N_4019);
or U4945 (N_4945,N_4168,N_4025);
or U4946 (N_4946,N_4141,N_4000);
and U4947 (N_4947,N_4286,N_4263);
nand U4948 (N_4948,N_4222,N_4743);
or U4949 (N_4949,N_4636,N_4123);
xnor U4950 (N_4950,N_4158,N_4049);
and U4951 (N_4951,N_3968,N_4367);
nand U4952 (N_4952,N_4427,N_3664);
or U4953 (N_4953,N_4156,N_4115);
xnor U4954 (N_4954,N_3867,N_4509);
or U4955 (N_4955,N_3657,N_3861);
nor U4956 (N_4956,N_4681,N_4744);
xnor U4957 (N_4957,N_3917,N_4484);
xnor U4958 (N_4958,N_3662,N_4560);
and U4959 (N_4959,N_4728,N_3732);
xnor U4960 (N_4960,N_3965,N_4244);
xnor U4961 (N_4961,N_3789,N_4296);
or U4962 (N_4962,N_3781,N_4024);
or U4963 (N_4963,N_4561,N_3696);
nor U4964 (N_4964,N_3628,N_4008);
and U4965 (N_4965,N_4456,N_4717);
nand U4966 (N_4966,N_4539,N_4698);
and U4967 (N_4967,N_4010,N_3676);
or U4968 (N_4968,N_4092,N_4445);
nand U4969 (N_4969,N_3720,N_4656);
nand U4970 (N_4970,N_4581,N_4397);
xor U4971 (N_4971,N_3937,N_4570);
xor U4972 (N_4972,N_3637,N_3847);
nand U4973 (N_4973,N_4332,N_3894);
or U4974 (N_4974,N_4325,N_4692);
nand U4975 (N_4975,N_4258,N_4221);
nand U4976 (N_4976,N_4317,N_4640);
and U4977 (N_4977,N_4351,N_4273);
and U4978 (N_4978,N_3748,N_4200);
nor U4979 (N_4979,N_3949,N_3909);
nand U4980 (N_4980,N_4515,N_4629);
and U4981 (N_4981,N_4747,N_4400);
or U4982 (N_4982,N_3921,N_3954);
nand U4983 (N_4983,N_4596,N_4542);
or U4984 (N_4984,N_4358,N_4183);
nor U4985 (N_4985,N_4239,N_4429);
nor U4986 (N_4986,N_3869,N_4795);
xnor U4987 (N_4987,N_4410,N_4290);
xor U4988 (N_4988,N_3784,N_4534);
and U4989 (N_4989,N_3751,N_4532);
nor U4990 (N_4990,N_4030,N_4214);
nand U4991 (N_4991,N_3995,N_4166);
or U4992 (N_4992,N_4181,N_4457);
xnor U4993 (N_4993,N_4420,N_4226);
and U4994 (N_4994,N_3680,N_4588);
xor U4995 (N_4995,N_4294,N_4084);
nand U4996 (N_4996,N_4621,N_3810);
nand U4997 (N_4997,N_4344,N_4139);
nand U4998 (N_4998,N_3815,N_4759);
or U4999 (N_4999,N_3922,N_4356);
nor U5000 (N_5000,N_3614,N_4231);
nor U5001 (N_5001,N_4120,N_4042);
or U5002 (N_5002,N_4544,N_4167);
nand U5003 (N_5003,N_4023,N_4067);
or U5004 (N_5004,N_4152,N_4748);
nand U5005 (N_5005,N_4459,N_4207);
and U5006 (N_5006,N_3850,N_4671);
and U5007 (N_5007,N_4399,N_4352);
or U5008 (N_5008,N_3902,N_4776);
nand U5009 (N_5009,N_4476,N_4350);
or U5010 (N_5010,N_4265,N_3673);
and U5011 (N_5011,N_4370,N_4613);
or U5012 (N_5012,N_4398,N_4148);
nor U5013 (N_5013,N_4796,N_3956);
and U5014 (N_5014,N_4213,N_3689);
nand U5015 (N_5015,N_4424,N_4606);
or U5016 (N_5016,N_3945,N_4046);
or U5017 (N_5017,N_3613,N_4134);
and U5018 (N_5018,N_4392,N_4114);
nor U5019 (N_5019,N_4074,N_3885);
nand U5020 (N_5020,N_4320,N_4710);
or U5021 (N_5021,N_4757,N_4274);
or U5022 (N_5022,N_3864,N_4366);
nand U5023 (N_5023,N_4132,N_4614);
xor U5024 (N_5024,N_4751,N_4205);
or U5025 (N_5025,N_3743,N_3982);
nand U5026 (N_5026,N_4297,N_4412);
nand U5027 (N_5027,N_4016,N_3685);
and U5028 (N_5028,N_4142,N_4669);
xor U5029 (N_5029,N_3852,N_4103);
xor U5030 (N_5030,N_4187,N_4572);
and U5031 (N_5031,N_4349,N_3830);
or U5032 (N_5032,N_4380,N_4057);
nand U5033 (N_5033,N_4219,N_4029);
nor U5034 (N_5034,N_3651,N_3991);
xor U5035 (N_5035,N_3983,N_4048);
or U5036 (N_5036,N_4298,N_4666);
nor U5037 (N_5037,N_3606,N_4464);
nand U5038 (N_5038,N_3744,N_3857);
xor U5039 (N_5039,N_3619,N_4760);
nor U5040 (N_5040,N_3695,N_3877);
and U5041 (N_5041,N_3659,N_4550);
and U5042 (N_5042,N_3693,N_4388);
or U5043 (N_5043,N_3758,N_4720);
or U5044 (N_5044,N_3977,N_3714);
nor U5045 (N_5045,N_4582,N_3878);
and U5046 (N_5046,N_4377,N_3871);
nand U5047 (N_5047,N_3611,N_4254);
xnor U5048 (N_5048,N_3999,N_4311);
and U5049 (N_5049,N_3905,N_3914);
nand U5050 (N_5050,N_4071,N_4051);
and U5051 (N_5051,N_4105,N_4062);
or U5052 (N_5052,N_3923,N_4365);
nand U5053 (N_5053,N_4571,N_3976);
nand U5054 (N_5054,N_3772,N_4558);
xor U5055 (N_5055,N_4448,N_3866);
and U5056 (N_5056,N_4409,N_3632);
nand U5057 (N_5057,N_4256,N_4124);
nand U5058 (N_5058,N_4341,N_4342);
nor U5059 (N_5059,N_3896,N_4481);
or U5060 (N_5060,N_3904,N_3752);
nand U5061 (N_5061,N_4259,N_4153);
and U5062 (N_5062,N_4630,N_3774);
nand U5063 (N_5063,N_3610,N_4343);
nor U5064 (N_5064,N_4670,N_3941);
and U5065 (N_5065,N_4705,N_4177);
nor U5066 (N_5066,N_4662,N_4353);
xnor U5067 (N_5067,N_3737,N_4327);
nand U5068 (N_5068,N_4701,N_4601);
or U5069 (N_5069,N_4291,N_4411);
and U5070 (N_5070,N_4261,N_3761);
nor U5071 (N_5071,N_4673,N_3813);
xnor U5072 (N_5072,N_3947,N_4251);
nor U5073 (N_5073,N_4474,N_3730);
nor U5074 (N_5074,N_4293,N_3715);
or U5075 (N_5075,N_3897,N_4079);
nand U5076 (N_5076,N_4069,N_4238);
nand U5077 (N_5077,N_3630,N_3868);
nor U5078 (N_5078,N_4703,N_4465);
nand U5079 (N_5079,N_4130,N_3931);
or U5080 (N_5080,N_4693,N_4264);
nand U5081 (N_5081,N_4375,N_4618);
and U5082 (N_5082,N_4337,N_4169);
or U5083 (N_5083,N_4138,N_3819);
nand U5084 (N_5084,N_3775,N_4752);
and U5085 (N_5085,N_4414,N_4111);
and U5086 (N_5086,N_4575,N_4304);
nor U5087 (N_5087,N_4070,N_4612);
nand U5088 (N_5088,N_3862,N_4180);
nand U5089 (N_5089,N_4711,N_3750);
and U5090 (N_5090,N_3724,N_4741);
xnor U5091 (N_5091,N_4635,N_3958);
nand U5092 (N_5092,N_4426,N_4490);
xor U5093 (N_5093,N_4573,N_4598);
xnor U5094 (N_5094,N_3920,N_4482);
nand U5095 (N_5095,N_3957,N_3895);
or U5096 (N_5096,N_3865,N_3739);
and U5097 (N_5097,N_4566,N_4727);
and U5098 (N_5098,N_4313,N_4699);
and U5099 (N_5099,N_4191,N_3706);
and U5100 (N_5100,N_4554,N_3747);
nor U5101 (N_5101,N_3778,N_4005);
nand U5102 (N_5102,N_3860,N_4530);
xnor U5103 (N_5103,N_4272,N_3623);
nor U5104 (N_5104,N_4508,N_3708);
and U5105 (N_5105,N_3690,N_4179);
xnor U5106 (N_5106,N_4516,N_4220);
and U5107 (N_5107,N_4178,N_4458);
nand U5108 (N_5108,N_4538,N_4546);
nand U5109 (N_5109,N_3890,N_3955);
nor U5110 (N_5110,N_4155,N_4610);
xnor U5111 (N_5111,N_4435,N_4562);
and U5112 (N_5112,N_3981,N_4044);
nor U5113 (N_5113,N_4326,N_4430);
or U5114 (N_5114,N_3853,N_4045);
and U5115 (N_5115,N_3616,N_4667);
nor U5116 (N_5116,N_3609,N_3771);
xnor U5117 (N_5117,N_4502,N_4233);
or U5118 (N_5118,N_3697,N_3944);
nor U5119 (N_5119,N_4758,N_3856);
nand U5120 (N_5120,N_4762,N_4083);
nor U5121 (N_5121,N_4001,N_4626);
nand U5122 (N_5122,N_4668,N_3738);
nand U5123 (N_5123,N_3805,N_4738);
or U5124 (N_5124,N_3661,N_4212);
nand U5125 (N_5125,N_3671,N_3838);
or U5126 (N_5126,N_4095,N_4372);
xnor U5127 (N_5127,N_4073,N_4250);
or U5128 (N_5128,N_4595,N_3663);
nor U5129 (N_5129,N_3855,N_3757);
nand U5130 (N_5130,N_3929,N_3794);
nor U5131 (N_5131,N_3858,N_4262);
and U5132 (N_5132,N_4529,N_4585);
nor U5133 (N_5133,N_4318,N_3655);
xor U5134 (N_5134,N_3886,N_4651);
and U5135 (N_5135,N_4734,N_4452);
nand U5136 (N_5136,N_4182,N_3692);
xor U5137 (N_5137,N_4746,N_3823);
nand U5138 (N_5138,N_4679,N_4089);
nand U5139 (N_5139,N_4524,N_4617);
nand U5140 (N_5140,N_3952,N_4040);
nand U5141 (N_5141,N_4136,N_3950);
nand U5142 (N_5142,N_4087,N_4210);
or U5143 (N_5143,N_4439,N_4682);
or U5144 (N_5144,N_4531,N_4470);
xor U5145 (N_5145,N_4147,N_4786);
and U5146 (N_5146,N_4282,N_3731);
or U5147 (N_5147,N_4129,N_4517);
xor U5148 (N_5148,N_4605,N_3681);
nor U5149 (N_5149,N_4135,N_4553);
nor U5150 (N_5150,N_4133,N_3797);
nor U5151 (N_5151,N_4753,N_3699);
and U5152 (N_5152,N_3600,N_4022);
nand U5153 (N_5153,N_4604,N_4633);
or U5154 (N_5154,N_4216,N_4731);
or U5155 (N_5155,N_3660,N_3916);
or U5156 (N_5156,N_4333,N_4654);
nand U5157 (N_5157,N_4162,N_3993);
xnor U5158 (N_5158,N_3654,N_4279);
nor U5159 (N_5159,N_4085,N_4483);
or U5160 (N_5160,N_3875,N_4535);
nor U5161 (N_5161,N_3666,N_4592);
xor U5162 (N_5162,N_4632,N_3908);
or U5163 (N_5163,N_4140,N_3780);
nand U5164 (N_5164,N_4685,N_3717);
and U5165 (N_5165,N_4781,N_3798);
nand U5166 (N_5166,N_3667,N_3605);
xnor U5167 (N_5167,N_4034,N_4736);
and U5168 (N_5168,N_4017,N_4033);
nor U5169 (N_5169,N_4184,N_3643);
xor U5170 (N_5170,N_4192,N_4525);
xnor U5171 (N_5171,N_4600,N_4473);
nand U5172 (N_5172,N_4623,N_3719);
or U5173 (N_5173,N_4714,N_4577);
nor U5174 (N_5174,N_4789,N_4631);
and U5175 (N_5175,N_3924,N_4390);
nor U5176 (N_5176,N_4003,N_3786);
or U5177 (N_5177,N_4406,N_4002);
xor U5178 (N_5178,N_3996,N_3918);
xor U5179 (N_5179,N_4518,N_3785);
nand U5180 (N_5180,N_3802,N_3969);
nor U5181 (N_5181,N_4599,N_4514);
nor U5182 (N_5182,N_3876,N_3953);
xnor U5183 (N_5183,N_4308,N_4607);
nand U5184 (N_5184,N_4761,N_4491);
or U5185 (N_5185,N_3779,N_4174);
xor U5186 (N_5186,N_3712,N_4310);
or U5187 (N_5187,N_4037,N_4253);
xor U5188 (N_5188,N_4721,N_4658);
xor U5189 (N_5189,N_4437,N_4401);
xnor U5190 (N_5190,N_3913,N_4674);
or U5191 (N_5191,N_3927,N_4235);
nor U5192 (N_5192,N_4396,N_4498);
nor U5193 (N_5193,N_4215,N_3978);
nand U5194 (N_5194,N_4035,N_4323);
nand U5195 (N_5195,N_4110,N_4204);
and U5196 (N_5196,N_3912,N_4075);
nand U5197 (N_5197,N_4793,N_3837);
nor U5198 (N_5198,N_3755,N_4229);
nor U5199 (N_5199,N_3846,N_4415);
or U5200 (N_5200,N_4797,N_4661);
xor U5201 (N_5201,N_3859,N_4324);
or U5202 (N_5202,N_4413,N_3903);
nand U5203 (N_5203,N_3618,N_4615);
nor U5204 (N_5204,N_3707,N_3640);
or U5205 (N_5205,N_4700,N_3615);
xor U5206 (N_5206,N_4431,N_3893);
and U5207 (N_5207,N_4302,N_4225);
or U5208 (N_5208,N_4039,N_4603);
or U5209 (N_5209,N_3668,N_4389);
and U5210 (N_5210,N_4196,N_4018);
nor U5211 (N_5211,N_4442,N_4675);
and U5212 (N_5212,N_3935,N_4108);
nor U5213 (N_5213,N_4113,N_3874);
nand U5214 (N_5214,N_4695,N_3626);
and U5215 (N_5215,N_3644,N_3647);
or U5216 (N_5216,N_3833,N_3898);
or U5217 (N_5217,N_4510,N_4094);
or U5218 (N_5218,N_4492,N_4418);
or U5219 (N_5219,N_4285,N_3975);
and U5220 (N_5220,N_4469,N_4373);
nor U5221 (N_5221,N_4557,N_4171);
nand U5222 (N_5222,N_4590,N_4766);
and U5223 (N_5223,N_3892,N_4245);
xnor U5224 (N_5224,N_4082,N_3961);
and U5225 (N_5225,N_4014,N_3808);
nor U5226 (N_5226,N_4730,N_3840);
xor U5227 (N_5227,N_4230,N_4742);
xnor U5228 (N_5228,N_4537,N_4660);
nand U5229 (N_5229,N_4289,N_4704);
nand U5230 (N_5230,N_4347,N_4379);
nand U5231 (N_5231,N_3691,N_3888);
or U5232 (N_5232,N_4417,N_4462);
or U5233 (N_5233,N_4576,N_4378);
nor U5234 (N_5234,N_4093,N_4712);
or U5235 (N_5235,N_4799,N_4199);
nor U5236 (N_5236,N_4716,N_3649);
nand U5237 (N_5237,N_4436,N_3716);
or U5238 (N_5238,N_4687,N_3806);
nor U5239 (N_5239,N_4487,N_4275);
nor U5240 (N_5240,N_4195,N_4619);
nand U5241 (N_5241,N_3656,N_4237);
nor U5242 (N_5242,N_4798,N_3990);
nand U5243 (N_5243,N_4394,N_4652);
or U5244 (N_5244,N_4549,N_4506);
nor U5245 (N_5245,N_4769,N_3809);
nor U5246 (N_5246,N_4257,N_4242);
and U5247 (N_5247,N_4004,N_4101);
nand U5248 (N_5248,N_4608,N_4548);
nor U5249 (N_5249,N_4478,N_4185);
and U5250 (N_5250,N_4319,N_3677);
xor U5251 (N_5251,N_4722,N_3939);
nor U5252 (N_5252,N_4443,N_4688);
and U5253 (N_5253,N_4485,N_3836);
xnor U5254 (N_5254,N_4568,N_3759);
and U5255 (N_5255,N_4718,N_4441);
nand U5256 (N_5256,N_4189,N_4580);
or U5257 (N_5257,N_4587,N_4193);
nor U5258 (N_5258,N_4503,N_4064);
or U5259 (N_5259,N_3829,N_4622);
and U5260 (N_5260,N_4006,N_4331);
xor U5261 (N_5261,N_4208,N_3911);
nor U5262 (N_5262,N_4077,N_4315);
nor U5263 (N_5263,N_4694,N_3624);
nand U5264 (N_5264,N_4565,N_4564);
nor U5265 (N_5265,N_4278,N_3701);
xor U5266 (N_5266,N_4763,N_4715);
xnor U5267 (N_5267,N_3790,N_3919);
nand U5268 (N_5268,N_3962,N_3992);
or U5269 (N_5269,N_4280,N_4203);
and U5270 (N_5270,N_3633,N_4647);
xnor U5271 (N_5271,N_4243,N_4186);
nand U5272 (N_5272,N_3642,N_4663);
and U5273 (N_5273,N_4137,N_4472);
and U5274 (N_5274,N_4433,N_3620);
or U5275 (N_5275,N_4770,N_3762);
xnor U5276 (N_5276,N_3851,N_3723);
nand U5277 (N_5277,N_3736,N_4360);
and U5278 (N_5278,N_4602,N_3799);
nand U5279 (N_5279,N_3936,N_3814);
nand U5280 (N_5280,N_4444,N_3733);
nand U5281 (N_5281,N_4556,N_4486);
and U5282 (N_5282,N_3811,N_4480);
xor U5283 (N_5283,N_3988,N_3870);
and U5284 (N_5284,N_3749,N_3741);
nand U5285 (N_5285,N_4173,N_3686);
nand U5286 (N_5286,N_4648,N_4197);
nor U5287 (N_5287,N_4767,N_4655);
xor U5288 (N_5288,N_4281,N_4540);
nor U5289 (N_5289,N_4404,N_4154);
nand U5290 (N_5290,N_3783,N_4755);
nand U5291 (N_5291,N_4513,N_3843);
and U5292 (N_5292,N_4369,N_3887);
or U5293 (N_5293,N_4450,N_4775);
xnor U5294 (N_5294,N_4055,N_4086);
or U5295 (N_5295,N_4494,N_4574);
xnor U5296 (N_5296,N_4247,N_4702);
or U5297 (N_5297,N_3951,N_4088);
or U5298 (N_5298,N_3889,N_3634);
nand U5299 (N_5299,N_4330,N_3926);
nor U5300 (N_5300,N_4547,N_4028);
nor U5301 (N_5301,N_3608,N_4036);
xor U5302 (N_5302,N_4706,N_4116);
nor U5303 (N_5303,N_4260,N_3820);
and U5304 (N_5304,N_4777,N_4321);
nor U5305 (N_5305,N_4144,N_3979);
or U5306 (N_5306,N_4784,N_4440);
nor U5307 (N_5307,N_4634,N_4467);
nor U5308 (N_5308,N_4098,N_4090);
nor U5309 (N_5309,N_3872,N_4336);
and U5310 (N_5310,N_4218,N_3763);
and U5311 (N_5311,N_4097,N_3621);
or U5312 (N_5312,N_4449,N_4362);
nand U5313 (N_5313,N_4387,N_3845);
nand U5314 (N_5314,N_4583,N_4119);
nand U5315 (N_5315,N_3711,N_3967);
and U5316 (N_5316,N_4791,N_4338);
nand U5317 (N_5317,N_4306,N_4295);
nand U5318 (N_5318,N_4312,N_4361);
nand U5319 (N_5319,N_4423,N_4419);
and U5320 (N_5320,N_3804,N_4160);
and U5321 (N_5321,N_3765,N_4194);
xnor U5322 (N_5322,N_4395,N_4725);
nand U5323 (N_5323,N_4012,N_3728);
and U5324 (N_5324,N_4122,N_4628);
and U5325 (N_5325,N_4007,N_4201);
and U5326 (N_5326,N_4060,N_3688);
nand U5327 (N_5327,N_3788,N_4112);
nor U5328 (N_5328,N_4526,N_4284);
or U5329 (N_5329,N_4348,N_4521);
and U5330 (N_5330,N_3604,N_3773);
nor U5331 (N_5331,N_4466,N_4672);
xnor U5332 (N_5332,N_4188,N_3863);
nor U5333 (N_5333,N_3687,N_3834);
nor U5334 (N_5334,N_4488,N_3817);
and U5335 (N_5335,N_4381,N_4032);
xnor U5336 (N_5336,N_3721,N_4627);
nand U5337 (N_5337,N_4780,N_4357);
nand U5338 (N_5338,N_4043,N_3938);
nor U5339 (N_5339,N_4300,N_4507);
nand U5340 (N_5340,N_4495,N_4792);
nor U5341 (N_5341,N_4496,N_4316);
or U5342 (N_5342,N_4223,N_3727);
nor U5343 (N_5343,N_4076,N_4723);
xnor U5344 (N_5344,N_3873,N_4421);
nand U5345 (N_5345,N_3880,N_4707);
nand U5346 (N_5346,N_4545,N_4774);
xor U5347 (N_5347,N_4234,N_4657);
and U5348 (N_5348,N_3928,N_4100);
or U5349 (N_5349,N_3675,N_4145);
nand U5350 (N_5350,N_3705,N_4386);
or U5351 (N_5351,N_3848,N_4505);
or U5352 (N_5352,N_3801,N_4737);
and U5353 (N_5353,N_4307,N_3694);
nand U5354 (N_5354,N_3986,N_3821);
xnor U5355 (N_5355,N_4209,N_3629);
xor U5356 (N_5356,N_4026,N_4266);
and U5357 (N_5357,N_3704,N_3966);
nor U5358 (N_5358,N_4594,N_4053);
xnor U5359 (N_5359,N_3971,N_4217);
and U5360 (N_5360,N_4638,N_4771);
nor U5361 (N_5361,N_4081,N_4267);
or U5362 (N_5362,N_4684,N_4788);
or U5363 (N_5363,N_4541,N_3746);
nor U5364 (N_5364,N_3718,N_4121);
nand U5365 (N_5365,N_4385,N_4334);
xor U5366 (N_5366,N_3795,N_3832);
and U5367 (N_5367,N_4190,N_3828);
nand U5368 (N_5368,N_4735,N_4374);
or U5369 (N_5369,N_3713,N_4125);
or U5370 (N_5370,N_4363,N_3946);
xnor U5371 (N_5371,N_4794,N_3827);
nor U5372 (N_5372,N_3980,N_4056);
or U5373 (N_5373,N_3722,N_4584);
or U5374 (N_5374,N_4616,N_3767);
nor U5375 (N_5375,N_3972,N_4665);
and U5376 (N_5376,N_4292,N_4339);
xnor U5377 (N_5377,N_4301,N_4523);
nand U5378 (N_5378,N_4477,N_4271);
xnor U5379 (N_5379,N_4405,N_4559);
xor U5380 (N_5380,N_3854,N_4455);
xnor U5381 (N_5381,N_3792,N_3960);
nand U5382 (N_5382,N_3602,N_4063);
and U5383 (N_5383,N_4104,N_3985);
nor U5384 (N_5384,N_3825,N_4157);
or U5385 (N_5385,N_3796,N_3734);
nand U5386 (N_5386,N_3812,N_4756);
xor U5387 (N_5387,N_3658,N_4645);
nor U5388 (N_5388,N_4172,N_4451);
or U5389 (N_5389,N_3839,N_4522);
xnor U5390 (N_5390,N_4696,N_4080);
and U5391 (N_5391,N_4128,N_4277);
xor U5392 (N_5392,N_4150,N_4428);
or U5393 (N_5393,N_3942,N_4020);
and U5394 (N_5394,N_4733,N_4276);
nor U5395 (N_5395,N_3791,N_4031);
or U5396 (N_5396,N_3816,N_4371);
or U5397 (N_5397,N_4589,N_4643);
or U5398 (N_5398,N_4175,N_4677);
nand U5399 (N_5399,N_3638,N_4248);
xnor U5400 (N_5400,N_4345,N_4545);
nand U5401 (N_5401,N_4300,N_4234);
and U5402 (N_5402,N_4374,N_4796);
nor U5403 (N_5403,N_4336,N_3790);
xnor U5404 (N_5404,N_4329,N_4192);
and U5405 (N_5405,N_4022,N_4386);
or U5406 (N_5406,N_4765,N_4460);
nand U5407 (N_5407,N_4028,N_4678);
or U5408 (N_5408,N_4017,N_4393);
nor U5409 (N_5409,N_4122,N_3968);
xor U5410 (N_5410,N_4539,N_4439);
xor U5411 (N_5411,N_4488,N_4268);
xor U5412 (N_5412,N_4013,N_4732);
nor U5413 (N_5413,N_4591,N_4153);
nor U5414 (N_5414,N_3966,N_3851);
or U5415 (N_5415,N_3761,N_4011);
and U5416 (N_5416,N_4788,N_4191);
xnor U5417 (N_5417,N_4511,N_3735);
or U5418 (N_5418,N_4442,N_4623);
or U5419 (N_5419,N_3673,N_3708);
and U5420 (N_5420,N_4370,N_4748);
xnor U5421 (N_5421,N_3744,N_4553);
or U5422 (N_5422,N_4772,N_3607);
nand U5423 (N_5423,N_4042,N_3935);
nor U5424 (N_5424,N_4004,N_4200);
or U5425 (N_5425,N_3697,N_4454);
nor U5426 (N_5426,N_3927,N_4282);
nand U5427 (N_5427,N_3847,N_4121);
xnor U5428 (N_5428,N_4037,N_4213);
nand U5429 (N_5429,N_4286,N_4599);
and U5430 (N_5430,N_4698,N_4344);
or U5431 (N_5431,N_3961,N_4682);
nor U5432 (N_5432,N_3725,N_4024);
nor U5433 (N_5433,N_3915,N_3932);
nand U5434 (N_5434,N_4724,N_4589);
xor U5435 (N_5435,N_3690,N_4641);
nor U5436 (N_5436,N_4492,N_4042);
nor U5437 (N_5437,N_4103,N_4230);
or U5438 (N_5438,N_4038,N_3745);
and U5439 (N_5439,N_3652,N_4639);
or U5440 (N_5440,N_4079,N_4603);
or U5441 (N_5441,N_4496,N_4502);
and U5442 (N_5442,N_4488,N_4074);
xnor U5443 (N_5443,N_4698,N_3605);
and U5444 (N_5444,N_4649,N_4284);
nor U5445 (N_5445,N_3906,N_4738);
nand U5446 (N_5446,N_4598,N_4215);
xor U5447 (N_5447,N_3689,N_3986);
xor U5448 (N_5448,N_3998,N_3763);
xnor U5449 (N_5449,N_4409,N_4063);
nor U5450 (N_5450,N_4435,N_4374);
or U5451 (N_5451,N_3640,N_4677);
and U5452 (N_5452,N_4163,N_4495);
and U5453 (N_5453,N_3988,N_4502);
and U5454 (N_5454,N_3887,N_4260);
or U5455 (N_5455,N_3852,N_3604);
nor U5456 (N_5456,N_4164,N_4540);
nand U5457 (N_5457,N_3631,N_4180);
or U5458 (N_5458,N_4656,N_4302);
xnor U5459 (N_5459,N_4387,N_3880);
nor U5460 (N_5460,N_3646,N_3787);
nor U5461 (N_5461,N_4670,N_3956);
xnor U5462 (N_5462,N_4554,N_4532);
nor U5463 (N_5463,N_3679,N_4457);
or U5464 (N_5464,N_4017,N_4564);
nand U5465 (N_5465,N_4444,N_4034);
or U5466 (N_5466,N_4079,N_4316);
xor U5467 (N_5467,N_4205,N_4605);
nand U5468 (N_5468,N_4638,N_3692);
xor U5469 (N_5469,N_4591,N_4791);
or U5470 (N_5470,N_3886,N_4683);
nand U5471 (N_5471,N_3804,N_3940);
nand U5472 (N_5472,N_4279,N_3942);
nand U5473 (N_5473,N_4002,N_3841);
xor U5474 (N_5474,N_4695,N_4033);
and U5475 (N_5475,N_4551,N_4624);
nand U5476 (N_5476,N_3943,N_3878);
nand U5477 (N_5477,N_3633,N_3989);
nor U5478 (N_5478,N_3739,N_4422);
or U5479 (N_5479,N_3688,N_3915);
nor U5480 (N_5480,N_4491,N_3835);
xor U5481 (N_5481,N_4787,N_4027);
nor U5482 (N_5482,N_4595,N_4512);
and U5483 (N_5483,N_4013,N_3799);
or U5484 (N_5484,N_4553,N_4636);
xnor U5485 (N_5485,N_3753,N_4297);
nand U5486 (N_5486,N_4463,N_4583);
nand U5487 (N_5487,N_4404,N_4071);
and U5488 (N_5488,N_4142,N_4754);
nand U5489 (N_5489,N_4250,N_3916);
and U5490 (N_5490,N_3810,N_4199);
and U5491 (N_5491,N_4207,N_3956);
nor U5492 (N_5492,N_4747,N_4577);
or U5493 (N_5493,N_4041,N_4777);
or U5494 (N_5494,N_3829,N_4303);
xnor U5495 (N_5495,N_3752,N_4097);
nand U5496 (N_5496,N_3740,N_3792);
or U5497 (N_5497,N_4411,N_3699);
or U5498 (N_5498,N_3807,N_3758);
or U5499 (N_5499,N_4246,N_4355);
xor U5500 (N_5500,N_3669,N_4157);
xor U5501 (N_5501,N_4120,N_4117);
nand U5502 (N_5502,N_4278,N_3986);
nand U5503 (N_5503,N_4589,N_4486);
nor U5504 (N_5504,N_3897,N_4565);
nor U5505 (N_5505,N_3693,N_3690);
nor U5506 (N_5506,N_4693,N_4405);
nand U5507 (N_5507,N_3986,N_3712);
and U5508 (N_5508,N_4601,N_4422);
and U5509 (N_5509,N_4599,N_4349);
nor U5510 (N_5510,N_3657,N_4104);
nand U5511 (N_5511,N_4280,N_4757);
xnor U5512 (N_5512,N_3668,N_3638);
or U5513 (N_5513,N_4301,N_4100);
xnor U5514 (N_5514,N_3866,N_4282);
or U5515 (N_5515,N_4631,N_4198);
and U5516 (N_5516,N_4690,N_4743);
xnor U5517 (N_5517,N_3640,N_4469);
and U5518 (N_5518,N_3685,N_3983);
nor U5519 (N_5519,N_4281,N_4787);
nand U5520 (N_5520,N_4465,N_4172);
xor U5521 (N_5521,N_4486,N_4733);
xor U5522 (N_5522,N_4509,N_4653);
nor U5523 (N_5523,N_4098,N_4352);
nor U5524 (N_5524,N_3660,N_3771);
and U5525 (N_5525,N_3768,N_4297);
and U5526 (N_5526,N_4179,N_4171);
or U5527 (N_5527,N_4123,N_3689);
nand U5528 (N_5528,N_4004,N_4388);
nand U5529 (N_5529,N_4773,N_4250);
and U5530 (N_5530,N_3943,N_3653);
or U5531 (N_5531,N_4532,N_4744);
nand U5532 (N_5532,N_3666,N_4429);
nand U5533 (N_5533,N_4793,N_4747);
nor U5534 (N_5534,N_4217,N_3724);
nand U5535 (N_5535,N_4678,N_4377);
and U5536 (N_5536,N_4774,N_4365);
xnor U5537 (N_5537,N_3775,N_4539);
and U5538 (N_5538,N_3793,N_4213);
nor U5539 (N_5539,N_3809,N_4148);
nand U5540 (N_5540,N_4755,N_4729);
xor U5541 (N_5541,N_3743,N_3796);
or U5542 (N_5542,N_4191,N_4745);
xnor U5543 (N_5543,N_4537,N_3640);
nand U5544 (N_5544,N_4552,N_4070);
and U5545 (N_5545,N_4512,N_4302);
and U5546 (N_5546,N_4586,N_4629);
and U5547 (N_5547,N_3784,N_4307);
nor U5548 (N_5548,N_4097,N_3670);
nand U5549 (N_5549,N_3973,N_4541);
and U5550 (N_5550,N_3983,N_4623);
xor U5551 (N_5551,N_4114,N_4237);
nand U5552 (N_5552,N_4259,N_4308);
nor U5553 (N_5553,N_4083,N_3950);
and U5554 (N_5554,N_4086,N_4507);
nand U5555 (N_5555,N_4378,N_3969);
nand U5556 (N_5556,N_3882,N_3649);
or U5557 (N_5557,N_4716,N_4441);
nor U5558 (N_5558,N_3682,N_4314);
nand U5559 (N_5559,N_3648,N_4717);
nand U5560 (N_5560,N_4160,N_3942);
nand U5561 (N_5561,N_3971,N_3615);
or U5562 (N_5562,N_4038,N_4112);
nand U5563 (N_5563,N_4761,N_4708);
nand U5564 (N_5564,N_4324,N_3601);
xnor U5565 (N_5565,N_4639,N_3836);
xnor U5566 (N_5566,N_3723,N_4782);
xnor U5567 (N_5567,N_4076,N_3681);
and U5568 (N_5568,N_4567,N_4746);
xnor U5569 (N_5569,N_4784,N_4582);
nor U5570 (N_5570,N_3869,N_4234);
nor U5571 (N_5571,N_3682,N_4626);
xor U5572 (N_5572,N_4467,N_4604);
or U5573 (N_5573,N_4307,N_4217);
or U5574 (N_5574,N_4665,N_4208);
nor U5575 (N_5575,N_3819,N_4412);
or U5576 (N_5576,N_4132,N_3604);
or U5577 (N_5577,N_3908,N_4617);
xnor U5578 (N_5578,N_4045,N_4778);
nor U5579 (N_5579,N_4383,N_3862);
and U5580 (N_5580,N_4695,N_4271);
nor U5581 (N_5581,N_4291,N_4150);
nor U5582 (N_5582,N_4213,N_4701);
or U5583 (N_5583,N_4578,N_3717);
or U5584 (N_5584,N_3717,N_4074);
or U5585 (N_5585,N_3845,N_3884);
xor U5586 (N_5586,N_3786,N_3790);
or U5587 (N_5587,N_3797,N_4456);
nor U5588 (N_5588,N_4286,N_3833);
nand U5589 (N_5589,N_3690,N_4260);
or U5590 (N_5590,N_3656,N_3916);
nand U5591 (N_5591,N_4570,N_3740);
or U5592 (N_5592,N_3874,N_4785);
or U5593 (N_5593,N_3777,N_4642);
nand U5594 (N_5594,N_4746,N_4170);
xnor U5595 (N_5595,N_4520,N_4444);
or U5596 (N_5596,N_3794,N_4174);
xnor U5597 (N_5597,N_4236,N_4455);
and U5598 (N_5598,N_4276,N_4649);
nand U5599 (N_5599,N_3933,N_4792);
nand U5600 (N_5600,N_4054,N_3794);
and U5601 (N_5601,N_4731,N_4763);
xor U5602 (N_5602,N_4662,N_4650);
xor U5603 (N_5603,N_3662,N_4517);
and U5604 (N_5604,N_3832,N_4127);
and U5605 (N_5605,N_3780,N_4305);
and U5606 (N_5606,N_4361,N_4465);
or U5607 (N_5607,N_4169,N_4205);
and U5608 (N_5608,N_4224,N_4798);
nor U5609 (N_5609,N_3912,N_4739);
or U5610 (N_5610,N_3805,N_4645);
nand U5611 (N_5611,N_4543,N_4480);
nor U5612 (N_5612,N_4191,N_4442);
or U5613 (N_5613,N_4654,N_4053);
nand U5614 (N_5614,N_4639,N_3629);
nand U5615 (N_5615,N_4545,N_3954);
or U5616 (N_5616,N_4325,N_4456);
nand U5617 (N_5617,N_4653,N_3922);
nor U5618 (N_5618,N_4642,N_3646);
and U5619 (N_5619,N_4414,N_4012);
nand U5620 (N_5620,N_4277,N_3890);
or U5621 (N_5621,N_4612,N_3875);
or U5622 (N_5622,N_4031,N_4592);
and U5623 (N_5623,N_4563,N_3993);
or U5624 (N_5624,N_4538,N_4203);
and U5625 (N_5625,N_4754,N_3984);
or U5626 (N_5626,N_4547,N_4737);
nor U5627 (N_5627,N_3888,N_3653);
or U5628 (N_5628,N_4625,N_4420);
or U5629 (N_5629,N_4374,N_3684);
or U5630 (N_5630,N_4230,N_4002);
or U5631 (N_5631,N_3619,N_3979);
nand U5632 (N_5632,N_3969,N_3665);
xor U5633 (N_5633,N_4694,N_3608);
nor U5634 (N_5634,N_3918,N_4248);
or U5635 (N_5635,N_4048,N_4229);
nand U5636 (N_5636,N_4395,N_4442);
and U5637 (N_5637,N_3729,N_4109);
nor U5638 (N_5638,N_3724,N_3819);
nor U5639 (N_5639,N_4706,N_4509);
nor U5640 (N_5640,N_4755,N_3643);
xor U5641 (N_5641,N_3600,N_3642);
or U5642 (N_5642,N_4290,N_4653);
nor U5643 (N_5643,N_4566,N_3964);
or U5644 (N_5644,N_4728,N_4532);
or U5645 (N_5645,N_3940,N_4282);
xor U5646 (N_5646,N_4085,N_3796);
or U5647 (N_5647,N_3772,N_3614);
xor U5648 (N_5648,N_3926,N_4492);
or U5649 (N_5649,N_3678,N_4014);
xnor U5650 (N_5650,N_3720,N_4493);
and U5651 (N_5651,N_4523,N_4772);
nor U5652 (N_5652,N_3689,N_3628);
and U5653 (N_5653,N_3907,N_4625);
xor U5654 (N_5654,N_4783,N_4247);
nand U5655 (N_5655,N_3896,N_4613);
or U5656 (N_5656,N_3674,N_4510);
nand U5657 (N_5657,N_4134,N_4776);
xor U5658 (N_5658,N_4740,N_4282);
nor U5659 (N_5659,N_4754,N_3912);
and U5660 (N_5660,N_3741,N_4736);
nor U5661 (N_5661,N_4139,N_4070);
nand U5662 (N_5662,N_4127,N_4605);
nor U5663 (N_5663,N_4106,N_3649);
nor U5664 (N_5664,N_3808,N_4421);
nand U5665 (N_5665,N_4260,N_4177);
nor U5666 (N_5666,N_4703,N_3920);
xnor U5667 (N_5667,N_4215,N_4741);
xnor U5668 (N_5668,N_4203,N_4635);
nand U5669 (N_5669,N_4638,N_4061);
or U5670 (N_5670,N_3651,N_3745);
nor U5671 (N_5671,N_4562,N_3969);
xor U5672 (N_5672,N_3962,N_4198);
nor U5673 (N_5673,N_4226,N_4601);
nand U5674 (N_5674,N_4501,N_3794);
nor U5675 (N_5675,N_3632,N_4418);
and U5676 (N_5676,N_4612,N_4698);
or U5677 (N_5677,N_4199,N_4654);
xor U5678 (N_5678,N_3688,N_4232);
xor U5679 (N_5679,N_4107,N_4500);
nand U5680 (N_5680,N_4185,N_4760);
xnor U5681 (N_5681,N_4052,N_4116);
xnor U5682 (N_5682,N_4589,N_4645);
or U5683 (N_5683,N_4024,N_4713);
xor U5684 (N_5684,N_4069,N_3780);
nor U5685 (N_5685,N_4704,N_3961);
or U5686 (N_5686,N_3816,N_3988);
and U5687 (N_5687,N_4543,N_4179);
nand U5688 (N_5688,N_3926,N_3838);
nor U5689 (N_5689,N_4799,N_3808);
and U5690 (N_5690,N_4360,N_3612);
nor U5691 (N_5691,N_3945,N_3666);
and U5692 (N_5692,N_4586,N_3826);
and U5693 (N_5693,N_4227,N_4063);
xor U5694 (N_5694,N_3611,N_4040);
nand U5695 (N_5695,N_4795,N_3989);
or U5696 (N_5696,N_4660,N_4533);
xnor U5697 (N_5697,N_4418,N_4715);
nand U5698 (N_5698,N_4730,N_4181);
or U5699 (N_5699,N_3864,N_4602);
or U5700 (N_5700,N_4114,N_3782);
xor U5701 (N_5701,N_4442,N_4093);
and U5702 (N_5702,N_4750,N_3789);
nand U5703 (N_5703,N_3779,N_4678);
xor U5704 (N_5704,N_3972,N_4463);
xor U5705 (N_5705,N_3996,N_4625);
xor U5706 (N_5706,N_3653,N_4319);
nor U5707 (N_5707,N_3664,N_4552);
and U5708 (N_5708,N_4083,N_4513);
nand U5709 (N_5709,N_3670,N_3674);
or U5710 (N_5710,N_4406,N_4760);
nand U5711 (N_5711,N_4300,N_4333);
and U5712 (N_5712,N_4183,N_4447);
nand U5713 (N_5713,N_4054,N_4665);
xor U5714 (N_5714,N_4688,N_4253);
nand U5715 (N_5715,N_4395,N_4390);
xor U5716 (N_5716,N_4238,N_3982);
nand U5717 (N_5717,N_4406,N_3673);
nor U5718 (N_5718,N_4745,N_4089);
nand U5719 (N_5719,N_4580,N_4150);
nand U5720 (N_5720,N_4688,N_3802);
nor U5721 (N_5721,N_4663,N_4178);
nor U5722 (N_5722,N_4502,N_4788);
or U5723 (N_5723,N_4649,N_4638);
nor U5724 (N_5724,N_4100,N_4556);
xnor U5725 (N_5725,N_3715,N_4194);
nor U5726 (N_5726,N_3712,N_4019);
or U5727 (N_5727,N_4732,N_4777);
and U5728 (N_5728,N_4773,N_4280);
or U5729 (N_5729,N_4136,N_3661);
and U5730 (N_5730,N_4256,N_4168);
and U5731 (N_5731,N_4626,N_4356);
nor U5732 (N_5732,N_3762,N_4062);
or U5733 (N_5733,N_4080,N_3751);
nand U5734 (N_5734,N_3728,N_3618);
nor U5735 (N_5735,N_4462,N_4742);
nand U5736 (N_5736,N_3660,N_4112);
nand U5737 (N_5737,N_3842,N_4551);
and U5738 (N_5738,N_3912,N_3779);
nor U5739 (N_5739,N_4085,N_3654);
and U5740 (N_5740,N_4442,N_4557);
and U5741 (N_5741,N_4359,N_4627);
nand U5742 (N_5742,N_3835,N_4170);
or U5743 (N_5743,N_4180,N_3752);
or U5744 (N_5744,N_4165,N_4009);
nand U5745 (N_5745,N_4748,N_4165);
and U5746 (N_5746,N_4401,N_4332);
nand U5747 (N_5747,N_4752,N_4014);
or U5748 (N_5748,N_4704,N_4658);
nand U5749 (N_5749,N_4516,N_3614);
nor U5750 (N_5750,N_3969,N_4436);
nand U5751 (N_5751,N_4553,N_4134);
nor U5752 (N_5752,N_4186,N_3771);
nor U5753 (N_5753,N_3903,N_3642);
nand U5754 (N_5754,N_3888,N_4523);
and U5755 (N_5755,N_4630,N_4716);
nor U5756 (N_5756,N_4234,N_3863);
or U5757 (N_5757,N_3659,N_3658);
nand U5758 (N_5758,N_4561,N_3923);
nand U5759 (N_5759,N_4676,N_4096);
or U5760 (N_5760,N_4066,N_4518);
xnor U5761 (N_5761,N_3757,N_4471);
and U5762 (N_5762,N_4536,N_4450);
and U5763 (N_5763,N_4660,N_3788);
or U5764 (N_5764,N_4285,N_4124);
nor U5765 (N_5765,N_3803,N_4103);
or U5766 (N_5766,N_4092,N_4355);
and U5767 (N_5767,N_3776,N_4271);
nand U5768 (N_5768,N_4324,N_4598);
and U5769 (N_5769,N_4380,N_3952);
and U5770 (N_5770,N_3815,N_3655);
nor U5771 (N_5771,N_4039,N_3639);
and U5772 (N_5772,N_4310,N_4257);
and U5773 (N_5773,N_3818,N_4206);
nand U5774 (N_5774,N_4793,N_4742);
or U5775 (N_5775,N_4398,N_4659);
nand U5776 (N_5776,N_4156,N_4082);
xor U5777 (N_5777,N_4739,N_3661);
and U5778 (N_5778,N_4630,N_3979);
or U5779 (N_5779,N_3716,N_3889);
nor U5780 (N_5780,N_3860,N_4105);
and U5781 (N_5781,N_4546,N_4191);
and U5782 (N_5782,N_4690,N_4598);
or U5783 (N_5783,N_3953,N_4332);
or U5784 (N_5784,N_4039,N_4375);
nor U5785 (N_5785,N_4319,N_4653);
nand U5786 (N_5786,N_4247,N_4227);
nand U5787 (N_5787,N_4337,N_4625);
or U5788 (N_5788,N_4216,N_4726);
nand U5789 (N_5789,N_3717,N_4780);
and U5790 (N_5790,N_3946,N_4045);
nand U5791 (N_5791,N_3676,N_3936);
nand U5792 (N_5792,N_3975,N_4588);
and U5793 (N_5793,N_4495,N_4461);
nand U5794 (N_5794,N_4127,N_3972);
nor U5795 (N_5795,N_4699,N_3781);
xnor U5796 (N_5796,N_4656,N_4682);
nor U5797 (N_5797,N_4086,N_4249);
and U5798 (N_5798,N_3654,N_3834);
nor U5799 (N_5799,N_4010,N_4475);
nand U5800 (N_5800,N_3788,N_4053);
and U5801 (N_5801,N_3702,N_4392);
and U5802 (N_5802,N_3649,N_3610);
and U5803 (N_5803,N_3700,N_4036);
nor U5804 (N_5804,N_3624,N_4495);
xnor U5805 (N_5805,N_4014,N_4147);
nand U5806 (N_5806,N_3920,N_3989);
nor U5807 (N_5807,N_3856,N_4240);
nand U5808 (N_5808,N_4057,N_4602);
nor U5809 (N_5809,N_3955,N_4420);
nor U5810 (N_5810,N_4495,N_4367);
xnor U5811 (N_5811,N_3949,N_4467);
and U5812 (N_5812,N_4241,N_4267);
or U5813 (N_5813,N_4789,N_3804);
nand U5814 (N_5814,N_3829,N_3973);
nor U5815 (N_5815,N_3900,N_3836);
or U5816 (N_5816,N_3878,N_3682);
xnor U5817 (N_5817,N_3961,N_4543);
xnor U5818 (N_5818,N_3728,N_3748);
xnor U5819 (N_5819,N_4124,N_4662);
and U5820 (N_5820,N_4544,N_4440);
nand U5821 (N_5821,N_3839,N_3946);
xnor U5822 (N_5822,N_4333,N_4757);
and U5823 (N_5823,N_4560,N_4760);
and U5824 (N_5824,N_4125,N_3859);
and U5825 (N_5825,N_4426,N_4261);
or U5826 (N_5826,N_4338,N_3950);
and U5827 (N_5827,N_3740,N_4199);
or U5828 (N_5828,N_3783,N_4277);
and U5829 (N_5829,N_4080,N_3891);
nand U5830 (N_5830,N_4180,N_3742);
nand U5831 (N_5831,N_3893,N_3638);
and U5832 (N_5832,N_4146,N_3823);
and U5833 (N_5833,N_4656,N_4770);
nor U5834 (N_5834,N_4535,N_4531);
nand U5835 (N_5835,N_4078,N_4669);
and U5836 (N_5836,N_4146,N_4101);
or U5837 (N_5837,N_3986,N_3979);
nand U5838 (N_5838,N_4058,N_4763);
nand U5839 (N_5839,N_4556,N_4063);
nand U5840 (N_5840,N_4060,N_3750);
nor U5841 (N_5841,N_3833,N_4674);
or U5842 (N_5842,N_4781,N_4484);
xnor U5843 (N_5843,N_3871,N_4150);
or U5844 (N_5844,N_4556,N_4188);
and U5845 (N_5845,N_4289,N_4216);
nand U5846 (N_5846,N_4276,N_4711);
xnor U5847 (N_5847,N_4112,N_4657);
xnor U5848 (N_5848,N_4249,N_4063);
nand U5849 (N_5849,N_3985,N_4690);
xor U5850 (N_5850,N_4521,N_4133);
or U5851 (N_5851,N_4400,N_4424);
xor U5852 (N_5852,N_4752,N_4353);
nor U5853 (N_5853,N_4796,N_3770);
nand U5854 (N_5854,N_4072,N_4552);
or U5855 (N_5855,N_4338,N_4662);
xor U5856 (N_5856,N_4038,N_4318);
nand U5857 (N_5857,N_4422,N_3734);
nand U5858 (N_5858,N_4039,N_4688);
nand U5859 (N_5859,N_4092,N_4055);
nor U5860 (N_5860,N_3610,N_4317);
xnor U5861 (N_5861,N_4458,N_4528);
or U5862 (N_5862,N_3843,N_3788);
and U5863 (N_5863,N_4233,N_4646);
xnor U5864 (N_5864,N_4176,N_4560);
xnor U5865 (N_5865,N_4768,N_4686);
and U5866 (N_5866,N_4374,N_4115);
or U5867 (N_5867,N_4355,N_3750);
or U5868 (N_5868,N_3905,N_4094);
nor U5869 (N_5869,N_3699,N_4296);
xor U5870 (N_5870,N_4414,N_3960);
xnor U5871 (N_5871,N_3922,N_4421);
and U5872 (N_5872,N_4445,N_4503);
nor U5873 (N_5873,N_4602,N_3683);
and U5874 (N_5874,N_3638,N_4523);
nand U5875 (N_5875,N_3805,N_4308);
nand U5876 (N_5876,N_4329,N_4788);
nor U5877 (N_5877,N_3623,N_3923);
or U5878 (N_5878,N_4238,N_4070);
nand U5879 (N_5879,N_4282,N_4593);
nor U5880 (N_5880,N_4151,N_3605);
nand U5881 (N_5881,N_4138,N_3787);
nor U5882 (N_5882,N_3623,N_4314);
nor U5883 (N_5883,N_4637,N_3762);
xor U5884 (N_5884,N_4735,N_4683);
and U5885 (N_5885,N_3935,N_4152);
and U5886 (N_5886,N_3913,N_3845);
nand U5887 (N_5887,N_4067,N_3600);
or U5888 (N_5888,N_3679,N_3981);
and U5889 (N_5889,N_4094,N_4570);
xnor U5890 (N_5890,N_4748,N_4606);
nand U5891 (N_5891,N_3848,N_4543);
xnor U5892 (N_5892,N_3975,N_4394);
nor U5893 (N_5893,N_3803,N_4273);
or U5894 (N_5894,N_4195,N_3990);
and U5895 (N_5895,N_4180,N_4159);
or U5896 (N_5896,N_4363,N_4128);
nor U5897 (N_5897,N_4468,N_4771);
nor U5898 (N_5898,N_3912,N_4514);
nor U5899 (N_5899,N_3606,N_4066);
nand U5900 (N_5900,N_4464,N_4376);
and U5901 (N_5901,N_4049,N_3918);
xnor U5902 (N_5902,N_3798,N_3983);
nor U5903 (N_5903,N_3871,N_4138);
or U5904 (N_5904,N_4727,N_4349);
nand U5905 (N_5905,N_3842,N_3900);
nor U5906 (N_5906,N_3989,N_3924);
nand U5907 (N_5907,N_4262,N_4575);
xor U5908 (N_5908,N_4093,N_4486);
or U5909 (N_5909,N_4579,N_3656);
or U5910 (N_5910,N_4562,N_4116);
nor U5911 (N_5911,N_4082,N_4511);
or U5912 (N_5912,N_4530,N_4560);
or U5913 (N_5913,N_3677,N_4158);
and U5914 (N_5914,N_4695,N_4588);
xnor U5915 (N_5915,N_4300,N_4082);
or U5916 (N_5916,N_4380,N_4659);
and U5917 (N_5917,N_4030,N_4111);
or U5918 (N_5918,N_4231,N_4053);
and U5919 (N_5919,N_3929,N_3824);
xor U5920 (N_5920,N_3937,N_4439);
and U5921 (N_5921,N_3634,N_3698);
nand U5922 (N_5922,N_4147,N_3952);
nor U5923 (N_5923,N_3880,N_4603);
and U5924 (N_5924,N_3616,N_4752);
or U5925 (N_5925,N_4270,N_4209);
nor U5926 (N_5926,N_3700,N_4628);
and U5927 (N_5927,N_4225,N_4220);
nand U5928 (N_5928,N_4573,N_4549);
nand U5929 (N_5929,N_4445,N_4276);
nand U5930 (N_5930,N_4054,N_3998);
xor U5931 (N_5931,N_3823,N_3699);
nand U5932 (N_5932,N_3988,N_4517);
nor U5933 (N_5933,N_3710,N_3755);
nor U5934 (N_5934,N_4473,N_4516);
nand U5935 (N_5935,N_3967,N_3892);
nor U5936 (N_5936,N_4252,N_4439);
and U5937 (N_5937,N_4253,N_4252);
nand U5938 (N_5938,N_4766,N_4109);
or U5939 (N_5939,N_3978,N_4401);
nand U5940 (N_5940,N_4569,N_4699);
or U5941 (N_5941,N_4454,N_4140);
or U5942 (N_5942,N_4303,N_4278);
or U5943 (N_5943,N_3680,N_3779);
nand U5944 (N_5944,N_3737,N_4603);
xor U5945 (N_5945,N_4788,N_3815);
xor U5946 (N_5946,N_3655,N_4593);
xnor U5947 (N_5947,N_4565,N_4725);
nor U5948 (N_5948,N_4590,N_4501);
and U5949 (N_5949,N_4188,N_4749);
nor U5950 (N_5950,N_4514,N_4387);
nand U5951 (N_5951,N_4263,N_4557);
nand U5952 (N_5952,N_4059,N_4101);
nand U5953 (N_5953,N_4410,N_4398);
or U5954 (N_5954,N_4710,N_4248);
nand U5955 (N_5955,N_4180,N_4134);
or U5956 (N_5956,N_3899,N_4044);
and U5957 (N_5957,N_4591,N_4556);
or U5958 (N_5958,N_4239,N_3979);
and U5959 (N_5959,N_3942,N_4473);
nor U5960 (N_5960,N_4421,N_3963);
xor U5961 (N_5961,N_3847,N_3841);
xnor U5962 (N_5962,N_4789,N_3633);
or U5963 (N_5963,N_3979,N_4761);
nand U5964 (N_5964,N_4020,N_4164);
nand U5965 (N_5965,N_3647,N_4512);
nor U5966 (N_5966,N_4798,N_4367);
nor U5967 (N_5967,N_4180,N_4219);
and U5968 (N_5968,N_4642,N_4300);
or U5969 (N_5969,N_4570,N_3919);
nand U5970 (N_5970,N_4595,N_4019);
and U5971 (N_5971,N_4332,N_4076);
nor U5972 (N_5972,N_4452,N_4751);
nor U5973 (N_5973,N_4063,N_4639);
and U5974 (N_5974,N_3647,N_3972);
nor U5975 (N_5975,N_3970,N_3974);
or U5976 (N_5976,N_3918,N_3885);
xor U5977 (N_5977,N_3708,N_4134);
and U5978 (N_5978,N_3820,N_4407);
xor U5979 (N_5979,N_4143,N_3733);
or U5980 (N_5980,N_4702,N_3948);
or U5981 (N_5981,N_4714,N_3881);
or U5982 (N_5982,N_3640,N_3741);
or U5983 (N_5983,N_4453,N_3968);
nand U5984 (N_5984,N_4702,N_4724);
nand U5985 (N_5985,N_3623,N_3739);
and U5986 (N_5986,N_4533,N_4506);
or U5987 (N_5987,N_4679,N_4305);
nor U5988 (N_5988,N_3737,N_4204);
and U5989 (N_5989,N_3673,N_4655);
xor U5990 (N_5990,N_3951,N_4181);
or U5991 (N_5991,N_4632,N_4249);
nor U5992 (N_5992,N_4496,N_3712);
nor U5993 (N_5993,N_4207,N_4398);
or U5994 (N_5994,N_3651,N_3806);
and U5995 (N_5995,N_3778,N_3609);
xnor U5996 (N_5996,N_4261,N_4323);
nand U5997 (N_5997,N_3767,N_4549);
xor U5998 (N_5998,N_3686,N_3734);
and U5999 (N_5999,N_3681,N_4268);
xnor U6000 (N_6000,N_5943,N_5475);
and U6001 (N_6001,N_4906,N_4995);
nor U6002 (N_6002,N_5073,N_5522);
and U6003 (N_6003,N_5589,N_5774);
nand U6004 (N_6004,N_5969,N_5361);
or U6005 (N_6005,N_5518,N_5819);
xnor U6006 (N_6006,N_4805,N_5516);
nand U6007 (N_6007,N_5906,N_5759);
nor U6008 (N_6008,N_5504,N_5473);
nor U6009 (N_6009,N_5862,N_4915);
nor U6010 (N_6010,N_4989,N_5183);
or U6011 (N_6011,N_5894,N_4821);
and U6012 (N_6012,N_5312,N_5338);
or U6013 (N_6013,N_5339,N_5793);
nand U6014 (N_6014,N_5854,N_5169);
nor U6015 (N_6015,N_5617,N_5344);
and U6016 (N_6016,N_5497,N_5388);
nor U6017 (N_6017,N_5807,N_5179);
nor U6018 (N_6018,N_5071,N_5374);
xnor U6019 (N_6019,N_5904,N_5148);
or U6020 (N_6020,N_4979,N_5562);
nand U6021 (N_6021,N_5709,N_5384);
and U6022 (N_6022,N_5353,N_5600);
or U6023 (N_6023,N_5653,N_5330);
and U6024 (N_6024,N_5279,N_5884);
xnor U6025 (N_6025,N_5947,N_5958);
nor U6026 (N_6026,N_5822,N_5735);
xor U6027 (N_6027,N_4991,N_5274);
and U6028 (N_6028,N_5983,N_5375);
and U6029 (N_6029,N_5980,N_5047);
and U6030 (N_6030,N_5424,N_5668);
nand U6031 (N_6031,N_5777,N_4985);
nand U6032 (N_6032,N_5354,N_5025);
nand U6033 (N_6033,N_5262,N_5520);
or U6034 (N_6034,N_5087,N_5283);
or U6035 (N_6035,N_5152,N_5981);
nand U6036 (N_6036,N_4828,N_5145);
or U6037 (N_6037,N_5769,N_5800);
xor U6038 (N_6038,N_5936,N_5010);
and U6039 (N_6039,N_5949,N_5515);
nand U6040 (N_6040,N_5242,N_5533);
nor U6041 (N_6041,N_5325,N_5125);
xor U6042 (N_6042,N_5260,N_5181);
or U6043 (N_6043,N_5607,N_5319);
nor U6044 (N_6044,N_5540,N_4822);
and U6045 (N_6045,N_5858,N_5123);
nand U6046 (N_6046,N_5840,N_4896);
and U6047 (N_6047,N_4964,N_4957);
nor U6048 (N_6048,N_5240,N_5397);
nand U6049 (N_6049,N_5965,N_5720);
nor U6050 (N_6050,N_5568,N_5514);
xor U6051 (N_6051,N_5824,N_4953);
or U6052 (N_6052,N_5147,N_5846);
or U6053 (N_6053,N_5491,N_4910);
and U6054 (N_6054,N_5622,N_5112);
nor U6055 (N_6055,N_5608,N_5068);
or U6056 (N_6056,N_4981,N_5582);
nand U6057 (N_6057,N_5650,N_5389);
nor U6058 (N_6058,N_5950,N_5027);
nor U6059 (N_6059,N_5198,N_5866);
nand U6060 (N_6060,N_5641,N_5869);
and U6061 (N_6061,N_5521,N_5892);
xnor U6062 (N_6062,N_5655,N_4983);
nor U6063 (N_6063,N_5511,N_5919);
and U6064 (N_6064,N_5215,N_4926);
xnor U6065 (N_6065,N_5646,N_5719);
nor U6066 (N_6066,N_5078,N_5470);
xnor U6067 (N_6067,N_5914,N_5923);
or U6068 (N_6068,N_5352,N_5435);
xor U6069 (N_6069,N_5953,N_5038);
nor U6070 (N_6070,N_4986,N_5150);
xnor U6071 (N_6071,N_5634,N_5432);
or U6072 (N_6072,N_4944,N_5941);
nor U6073 (N_6073,N_4950,N_5201);
nand U6074 (N_6074,N_5826,N_5626);
and U6075 (N_6075,N_5860,N_5924);
nand U6076 (N_6076,N_4952,N_5405);
nor U6077 (N_6077,N_5083,N_5539);
and U6078 (N_6078,N_5591,N_5697);
xor U6079 (N_6079,N_5736,N_5212);
nor U6080 (N_6080,N_5502,N_5080);
nand U6081 (N_6081,N_5391,N_4881);
nor U6082 (N_6082,N_4929,N_5633);
nand U6083 (N_6083,N_5954,N_5378);
nand U6084 (N_6084,N_5429,N_5844);
and U6085 (N_6085,N_5244,N_5452);
xor U6086 (N_6086,N_5088,N_5744);
or U6087 (N_6087,N_5086,N_4809);
and U6088 (N_6088,N_5509,N_5238);
xnor U6089 (N_6089,N_5368,N_5155);
or U6090 (N_6090,N_5531,N_5865);
and U6091 (N_6091,N_5098,N_5304);
and U6092 (N_6092,N_5971,N_5786);
or U6093 (N_6093,N_5792,N_5915);
and U6094 (N_6094,N_5801,N_4891);
xnor U6095 (N_6095,N_5692,N_5898);
and U6096 (N_6096,N_5265,N_4824);
xor U6097 (N_6097,N_5783,N_5340);
nor U6098 (N_6098,N_4988,N_5482);
nor U6099 (N_6099,N_5726,N_4912);
and U6100 (N_6100,N_5109,N_5929);
and U6101 (N_6101,N_5317,N_5925);
and U6102 (N_6102,N_5448,N_5507);
and U6103 (N_6103,N_5679,N_5610);
nor U6104 (N_6104,N_5615,N_5839);
or U6105 (N_6105,N_5479,N_4801);
xnor U6106 (N_6106,N_5671,N_5829);
or U6107 (N_6107,N_5111,N_5324);
or U6108 (N_6108,N_5072,N_5036);
nor U6109 (N_6109,N_5921,N_5146);
nor U6110 (N_6110,N_4997,N_5308);
and U6111 (N_6111,N_5237,N_5165);
nor U6112 (N_6112,N_5381,N_5657);
nand U6113 (N_6113,N_5398,N_5416);
xor U6114 (N_6114,N_4874,N_5439);
nand U6115 (N_6115,N_5296,N_5942);
xnor U6116 (N_6116,N_5833,N_5661);
nor U6117 (N_6117,N_4845,N_4954);
nor U6118 (N_6118,N_5253,N_5422);
xor U6119 (N_6119,N_5433,N_5842);
or U6120 (N_6120,N_5951,N_5673);
nor U6121 (N_6121,N_5138,N_4928);
xor U6122 (N_6122,N_5986,N_5809);
xor U6123 (N_6123,N_5306,N_5670);
nor U6124 (N_6124,N_5945,N_5816);
xnor U6125 (N_6125,N_5506,N_5908);
nand U6126 (N_6126,N_5289,N_4806);
nand U6127 (N_6127,N_5415,N_4897);
xnor U6128 (N_6128,N_5041,N_5498);
nand U6129 (N_6129,N_5042,N_4987);
or U6130 (N_6130,N_4931,N_5779);
nand U6131 (N_6131,N_4888,N_5016);
or U6132 (N_6132,N_5794,N_4898);
and U6133 (N_6133,N_5104,N_5838);
xor U6134 (N_6134,N_5367,N_5758);
xnor U6135 (N_6135,N_4917,N_5130);
nor U6136 (N_6136,N_5303,N_5040);
nand U6137 (N_6137,N_5191,N_5689);
or U6138 (N_6138,N_4834,N_5836);
nand U6139 (N_6139,N_5768,N_5402);
nand U6140 (N_6140,N_5233,N_5170);
nor U6141 (N_6141,N_5092,N_4977);
or U6142 (N_6142,N_4855,N_4992);
and U6143 (N_6143,N_5723,N_5747);
or U6144 (N_6144,N_5229,N_5024);
or U6145 (N_6145,N_5311,N_5246);
nor U6146 (N_6146,N_5117,N_5553);
nor U6147 (N_6147,N_5911,N_5300);
and U6148 (N_6148,N_5133,N_5992);
or U6149 (N_6149,N_5535,N_4866);
xnor U6150 (N_6150,N_5756,N_4930);
nor U6151 (N_6151,N_5820,N_5772);
and U6152 (N_6152,N_5210,N_4933);
or U6153 (N_6153,N_5458,N_5185);
xnor U6154 (N_6154,N_5815,N_4868);
or U6155 (N_6155,N_4965,N_5828);
and U6156 (N_6156,N_4894,N_5484);
and U6157 (N_6157,N_4826,N_4984);
nor U6158 (N_6158,N_5188,N_5619);
or U6159 (N_6159,N_5536,N_5857);
nor U6160 (N_6160,N_5206,N_5314);
xnor U6161 (N_6161,N_5285,N_5167);
xnor U6162 (N_6162,N_5970,N_4938);
nor U6163 (N_6163,N_5952,N_5910);
and U6164 (N_6164,N_4803,N_5392);
and U6165 (N_6165,N_5000,N_5383);
or U6166 (N_6166,N_5703,N_5849);
xor U6167 (N_6167,N_5213,N_5302);
nor U6168 (N_6168,N_5814,N_5868);
xor U6169 (N_6169,N_5767,N_5897);
xor U6170 (N_6170,N_5399,N_4859);
nand U6171 (N_6171,N_5879,N_4890);
and U6172 (N_6172,N_5499,N_5021);
or U6173 (N_6173,N_5032,N_5920);
nand U6174 (N_6174,N_4889,N_5594);
nand U6175 (N_6175,N_4836,N_4862);
nand U6176 (N_6176,N_5834,N_5883);
or U6177 (N_6177,N_5382,N_5065);
nor U6178 (N_6178,N_5343,N_5688);
nor U6179 (N_6179,N_4851,N_5550);
and U6180 (N_6180,N_4841,N_5139);
nor U6181 (N_6181,N_5575,N_5168);
nor U6182 (N_6182,N_5813,N_5691);
xnor U6183 (N_6183,N_5420,N_4852);
or U6184 (N_6184,N_5926,N_5160);
and U6185 (N_6185,N_5176,N_5494);
nor U6186 (N_6186,N_4942,N_5297);
or U6187 (N_6187,N_5293,N_5790);
or U6188 (N_6188,N_4902,N_4921);
xor U6189 (N_6189,N_5128,N_5707);
nand U6190 (N_6190,N_5284,N_5708);
or U6191 (N_6191,N_5364,N_5171);
nand U6192 (N_6192,N_5488,N_5644);
xor U6193 (N_6193,N_5856,N_5318);
or U6194 (N_6194,N_5269,N_5863);
nand U6195 (N_6195,N_5789,N_5802);
xnor U6196 (N_6196,N_5893,N_5593);
xor U6197 (N_6197,N_5075,N_5554);
or U6198 (N_6198,N_5292,N_4967);
nor U6199 (N_6199,N_5320,N_5525);
and U6200 (N_6200,N_5887,N_4849);
or U6201 (N_6201,N_5234,N_5738);
and U6202 (N_6202,N_5698,N_5453);
or U6203 (N_6203,N_4885,N_4839);
or U6204 (N_6204,N_5379,N_5564);
or U6205 (N_6205,N_5366,N_5418);
nor U6206 (N_6206,N_5326,N_4937);
and U6207 (N_6207,N_5408,N_5574);
xnor U6208 (N_6208,N_5806,N_5187);
nor U6209 (N_6209,N_5658,N_5103);
xor U6210 (N_6210,N_4951,N_4846);
nor U6211 (N_6211,N_5116,N_5276);
xor U6212 (N_6212,N_5063,N_5751);
or U6213 (N_6213,N_5180,N_4804);
and U6214 (N_6214,N_5172,N_5136);
nor U6215 (N_6215,N_5465,N_5226);
xnor U6216 (N_6216,N_5216,N_5775);
and U6217 (N_6217,N_5725,N_4811);
xnor U6218 (N_6218,N_5254,N_4800);
nor U6219 (N_6219,N_5323,N_5079);
nor U6220 (N_6220,N_5604,N_5939);
nand U6221 (N_6221,N_4895,N_4940);
and U6222 (N_6222,N_5263,N_5114);
xnor U6223 (N_6223,N_5282,N_5651);
or U6224 (N_6224,N_5766,N_5053);
nor U6225 (N_6225,N_5665,N_5876);
and U6226 (N_6226,N_5023,N_5870);
nand U6227 (N_6227,N_5606,N_5545);
nor U6228 (N_6228,N_5592,N_4999);
and U6229 (N_6229,N_5076,N_5144);
or U6230 (N_6230,N_5557,N_5596);
nor U6231 (N_6231,N_5818,N_5476);
xor U6232 (N_6232,N_5648,N_5695);
nand U6233 (N_6233,N_5649,N_5218);
nor U6234 (N_6234,N_4850,N_5446);
and U6235 (N_6235,N_5624,N_4923);
xnor U6236 (N_6236,N_5890,N_5044);
nor U6237 (N_6237,N_5249,N_5517);
nor U6238 (N_6238,N_5590,N_5985);
nor U6239 (N_6239,N_5734,N_4908);
xor U6240 (N_6240,N_5529,N_5852);
xnor U6241 (N_6241,N_5436,N_5636);
and U6242 (N_6242,N_5549,N_4990);
or U6243 (N_6243,N_5565,N_5154);
or U6244 (N_6244,N_5380,N_4878);
or U6245 (N_6245,N_5745,N_5472);
nand U6246 (N_6246,N_5528,N_5257);
or U6247 (N_6247,N_4945,N_5853);
xnor U6248 (N_6248,N_5960,N_5605);
and U6249 (N_6249,N_5683,N_5395);
nor U6250 (N_6250,N_5447,N_5552);
nor U6251 (N_6251,N_5483,N_5394);
xnor U6252 (N_6252,N_5752,N_5674);
nor U6253 (N_6253,N_5687,N_5107);
xnor U6254 (N_6254,N_5737,N_5390);
nand U6255 (N_6255,N_5578,N_5537);
nand U6256 (N_6256,N_5885,N_5938);
or U6257 (N_6257,N_5918,N_5310);
or U6258 (N_6258,N_5715,N_5640);
and U6259 (N_6259,N_5430,N_5749);
nor U6260 (N_6260,N_5055,N_4843);
xor U6261 (N_6261,N_5663,N_5696);
and U6262 (N_6262,N_5855,N_4970);
or U6263 (N_6263,N_5362,N_4971);
nor U6264 (N_6264,N_5933,N_5239);
nand U6265 (N_6265,N_5119,N_5827);
nor U6266 (N_6266,N_5110,N_4832);
nor U6267 (N_6267,N_5332,N_5355);
xnor U6268 (N_6268,N_5746,N_5232);
xor U6269 (N_6269,N_5175,N_5796);
and U6270 (N_6270,N_5159,N_5995);
nor U6271 (N_6271,N_5329,N_5990);
xor U6272 (N_6272,N_5327,N_5664);
nand U6273 (N_6273,N_5222,N_5837);
and U6274 (N_6274,N_5255,N_5486);
nor U6275 (N_6275,N_5204,N_4814);
xor U6276 (N_6276,N_5121,N_5930);
and U6277 (N_6277,N_5850,N_5157);
nand U6278 (N_6278,N_5984,N_5882);
and U6279 (N_6279,N_5008,N_5077);
and U6280 (N_6280,N_5654,N_4857);
nand U6281 (N_6281,N_4907,N_5230);
nor U6282 (N_6282,N_5621,N_5508);
nor U6283 (N_6283,N_5532,N_5106);
and U6284 (N_6284,N_5427,N_5916);
xor U6285 (N_6285,N_5357,N_4918);
nand U6286 (N_6286,N_4823,N_5443);
xor U6287 (N_6287,N_5988,N_5334);
nand U6288 (N_6288,N_5419,N_5294);
nand U6289 (N_6289,N_5195,N_5132);
or U6290 (N_6290,N_5645,N_5248);
xnor U6291 (N_6291,N_4949,N_5135);
or U6292 (N_6292,N_5421,N_5903);
xor U6293 (N_6293,N_5760,N_5100);
or U6294 (N_6294,N_5817,N_5880);
xor U6295 (N_6295,N_5753,N_5026);
or U6296 (N_6296,N_5156,N_5652);
or U6297 (N_6297,N_5825,N_5616);
and U6298 (N_6298,N_5444,N_4955);
nor U6299 (N_6299,N_4813,N_5001);
and U6300 (N_6300,N_5821,N_5888);
and U6301 (N_6301,N_5441,N_5987);
nand U6302 (N_6302,N_5740,N_5129);
and U6303 (N_6303,N_5174,N_5713);
and U6304 (N_6304,N_5913,N_5280);
xor U6305 (N_6305,N_5750,N_4830);
and U6306 (N_6306,N_5770,N_5886);
nor U6307 (N_6307,N_5561,N_5989);
nor U6308 (N_6308,N_4920,N_5700);
xnor U6309 (N_6309,N_5712,N_5084);
nand U6310 (N_6310,N_5909,N_5586);
or U6311 (N_6311,N_5396,N_5467);
and U6312 (N_6312,N_4833,N_4810);
xor U6313 (N_6313,N_5881,N_5754);
nand U6314 (N_6314,N_5702,N_5597);
nor U6315 (N_6315,N_5599,N_4922);
nand U6316 (N_6316,N_5523,N_5386);
xor U6317 (N_6317,N_5931,N_5957);
nand U6318 (N_6318,N_5048,N_4871);
xor U6319 (N_6319,N_5463,N_5051);
nor U6320 (N_6320,N_5228,N_4935);
nor U6321 (N_6321,N_5718,N_5336);
and U6322 (N_6322,N_5959,N_5823);
xnor U6323 (N_6323,N_5124,N_5406);
xor U6324 (N_6324,N_4876,N_4847);
and U6325 (N_6325,N_5351,N_5099);
and U6326 (N_6326,N_5315,N_5997);
nand U6327 (N_6327,N_5478,N_5322);
nor U6328 (N_6328,N_5546,N_5524);
or U6329 (N_6329,N_5050,N_5151);
nor U6330 (N_6330,N_5677,N_5808);
xor U6331 (N_6331,N_5773,N_4901);
nand U6332 (N_6332,N_5178,N_4972);
or U6333 (N_6333,N_5643,N_5804);
or U6334 (N_6334,N_4966,N_5118);
xnor U6335 (N_6335,N_4808,N_5035);
or U6336 (N_6336,N_5999,N_5601);
or U6337 (N_6337,N_5732,N_5140);
nor U6338 (N_6338,N_5991,N_5871);
xor U6339 (N_6339,N_5544,N_4960);
nor U6340 (N_6340,N_5012,N_5602);
nand U6341 (N_6341,N_5611,N_5681);
and U6342 (N_6342,N_5627,N_5143);
nor U6343 (N_6343,N_5481,N_5309);
or U6344 (N_6344,N_5895,N_5266);
and U6345 (N_6345,N_5328,N_5757);
xor U6346 (N_6346,N_5227,N_5678);
and U6347 (N_6347,N_5505,N_5457);
xnor U6348 (N_6348,N_4817,N_4816);
or U6349 (N_6349,N_5731,N_5363);
or U6350 (N_6350,N_4893,N_5031);
nor U6351 (N_6351,N_5542,N_4909);
nand U6352 (N_6352,N_5963,N_5037);
nor U6353 (N_6353,N_5161,N_4982);
xnor U6354 (N_6354,N_5131,N_5994);
or U6355 (N_6355,N_5434,N_5449);
or U6356 (N_6356,N_5716,N_5468);
or U6357 (N_6357,N_5928,N_5085);
xor U6358 (N_6358,N_5270,N_5094);
nand U6359 (N_6359,N_4975,N_5900);
xor U6360 (N_6360,N_4867,N_5799);
nor U6361 (N_6361,N_5975,N_5203);
nand U6362 (N_6362,N_5966,N_5376);
and U6363 (N_6363,N_5555,N_5462);
nand U6364 (N_6364,N_5584,N_4934);
and U6365 (N_6365,N_5638,N_5830);
nor U6366 (N_6366,N_5199,N_5305);
or U6367 (N_6367,N_5007,N_5291);
or U6368 (N_6368,N_4887,N_5207);
xor U6369 (N_6369,N_5243,N_5009);
nor U6370 (N_6370,N_5955,N_4870);
or U6371 (N_6371,N_5061,N_5872);
nand U6372 (N_6372,N_5074,N_5934);
or U6373 (N_6373,N_5487,N_5371);
nor U6374 (N_6374,N_5033,N_4860);
xor U6375 (N_6375,N_5360,N_5186);
xor U6376 (N_6376,N_5571,N_5637);
and U6377 (N_6377,N_5141,N_4827);
nor U6378 (N_6378,N_4853,N_5197);
xor U6379 (N_6379,N_5797,N_5058);
xnor U6380 (N_6380,N_4873,N_5579);
xnor U6381 (N_6381,N_5097,N_4820);
nor U6382 (N_6382,N_5414,N_5275);
nor U6383 (N_6383,N_5059,N_5847);
nand U6384 (N_6384,N_5469,N_5864);
xnor U6385 (N_6385,N_5445,N_4962);
nand U6386 (N_6386,N_4883,N_4911);
nor U6387 (N_6387,N_5935,N_4996);
nor U6388 (N_6388,N_5656,N_5543);
or U6389 (N_6389,N_5581,N_4969);
xnor U6390 (N_6390,N_5017,N_5460);
nand U6391 (N_6391,N_5019,N_5043);
or U6392 (N_6392,N_5425,N_5843);
xnor U6393 (N_6393,N_5787,N_5580);
and U6394 (N_6394,N_5845,N_5996);
or U6395 (N_6395,N_5451,N_5020);
nor U6396 (N_6396,N_5559,N_4924);
and U6397 (N_6397,N_5261,N_5417);
and U6398 (N_6398,N_5316,N_4872);
nor U6399 (N_6399,N_5192,N_5587);
xor U6400 (N_6400,N_5273,N_5729);
and U6401 (N_6401,N_5978,N_5630);
or U6402 (N_6402,N_5676,N_5937);
xor U6403 (N_6403,N_5173,N_5477);
nand U6404 (N_6404,N_5803,N_5742);
nand U6405 (N_6405,N_5002,N_5861);
nor U6406 (N_6406,N_5558,N_5224);
and U6407 (N_6407,N_5595,N_5538);
and U6408 (N_6408,N_5474,N_4858);
xor U6409 (N_6409,N_5321,N_5190);
nor U6410 (N_6410,N_4879,N_5685);
and U6411 (N_6411,N_5659,N_4815);
or U6412 (N_6412,N_5070,N_5899);
xor U6413 (N_6413,N_5049,N_5976);
or U6414 (N_6414,N_5454,N_5278);
nand U6415 (N_6415,N_5705,N_5917);
and U6416 (N_6416,N_5585,N_5346);
xor U6417 (N_6417,N_5603,N_4865);
xor U6418 (N_6418,N_5778,N_4829);
and U6419 (N_6419,N_5798,N_4914);
nand U6420 (N_6420,N_5003,N_5841);
nor U6421 (N_6421,N_5572,N_5295);
and U6422 (N_6422,N_5214,N_5831);
nand U6423 (N_6423,N_5795,N_5612);
xor U6424 (N_6424,N_5556,N_5231);
nand U6425 (N_6425,N_5200,N_5331);
and U6426 (N_6426,N_5307,N_5495);
nand U6427 (N_6427,N_5889,N_5301);
and U6428 (N_6428,N_5570,N_5788);
and U6429 (N_6429,N_5721,N_5961);
or U6430 (N_6430,N_4864,N_5694);
xor U6431 (N_6431,N_5387,N_5493);
nor U6432 (N_6432,N_4904,N_5534);
nor U6433 (N_6433,N_5287,N_4948);
nand U6434 (N_6434,N_5513,N_5771);
nor U6435 (N_6435,N_5905,N_5962);
xor U6436 (N_6436,N_5998,N_4825);
xnor U6437 (N_6437,N_5358,N_5193);
and U6438 (N_6438,N_5241,N_4869);
nand U6439 (N_6439,N_5902,N_5411);
nor U6440 (N_6440,N_5022,N_5877);
nor U6441 (N_6441,N_4974,N_5333);
and U6442 (N_6442,N_5781,N_5639);
nand U6443 (N_6443,N_5166,N_4959);
xor U6444 (N_6444,N_4886,N_5347);
xor U6445 (N_6445,N_4958,N_5034);
nand U6446 (N_6446,N_4875,N_4807);
and U6447 (N_6447,N_4963,N_5526);
and U6448 (N_6448,N_5632,N_5548);
xnor U6449 (N_6449,N_5583,N_5761);
xor U6450 (N_6450,N_5510,N_4941);
or U6451 (N_6451,N_5728,N_5625);
nor U6452 (N_6452,N_5972,N_4932);
nor U6453 (N_6453,N_4842,N_5805);
xnor U6454 (N_6454,N_5867,N_5496);
nor U6455 (N_6455,N_4905,N_5054);
or U6456 (N_6456,N_5205,N_5567);
xnor U6457 (N_6457,N_5973,N_5286);
nand U6458 (N_6458,N_5993,N_5219);
nor U6459 (N_6459,N_5052,N_5717);
nor U6460 (N_6460,N_5530,N_5979);
nand U6461 (N_6461,N_5456,N_5013);
nor U6462 (N_6462,N_5428,N_5202);
xnor U6463 (N_6463,N_5369,N_5250);
nand U6464 (N_6464,N_5182,N_4899);
xnor U6465 (N_6465,N_4946,N_5551);
nand U6466 (N_6466,N_5946,N_5089);
nand U6467 (N_6467,N_4802,N_5461);
nand U6468 (N_6468,N_5710,N_5810);
nor U6469 (N_6469,N_5722,N_4819);
or U6470 (N_6470,N_5006,N_4913);
nor U6471 (N_6471,N_5209,N_5335);
nor U6472 (N_6472,N_5404,N_5459);
xor U6473 (N_6473,N_5350,N_5512);
and U6474 (N_6474,N_4994,N_5045);
or U6475 (N_6475,N_5784,N_5113);
or U6476 (N_6476,N_5891,N_5785);
xnor U6477 (N_6477,N_5409,N_5137);
or U6478 (N_6478,N_5763,N_4861);
xnor U6479 (N_6479,N_4844,N_5851);
or U6480 (N_6480,N_5401,N_5039);
nand U6481 (N_6481,N_5609,N_5733);
and U6482 (N_6482,N_5848,N_5811);
or U6483 (N_6483,N_5741,N_5267);
nor U6484 (N_6484,N_5385,N_5503);
or U6485 (N_6485,N_4980,N_5588);
nand U6486 (N_6486,N_5056,N_5755);
nand U6487 (N_6487,N_5102,N_5480);
or U6488 (N_6488,N_5365,N_5245);
xor U6489 (N_6489,N_5256,N_5014);
nor U6490 (N_6490,N_5066,N_5356);
and U6491 (N_6491,N_5413,N_5873);
and U6492 (N_6492,N_5684,N_5944);
nor U6493 (N_6493,N_5057,N_5407);
and U6494 (N_6494,N_5901,N_5108);
nor U6495 (N_6495,N_5628,N_5948);
and U6496 (N_6496,N_4835,N_5127);
nand U6497 (N_6497,N_4840,N_5964);
nor U6498 (N_6498,N_5091,N_5563);
or U6499 (N_6499,N_4927,N_4812);
nand U6500 (N_6500,N_5120,N_5101);
xor U6501 (N_6501,N_4961,N_5667);
nor U6502 (N_6502,N_5560,N_4943);
nand U6503 (N_6503,N_4856,N_5922);
or U6504 (N_6504,N_5184,N_5372);
and U6505 (N_6505,N_4880,N_5598);
nor U6506 (N_6506,N_5686,N_5631);
xnor U6507 (N_6507,N_5153,N_5223);
xnor U6508 (N_6508,N_5450,N_5730);
and U6509 (N_6509,N_5666,N_5221);
or U6510 (N_6510,N_5765,N_5442);
and U6511 (N_6511,N_5464,N_5748);
nor U6512 (N_6512,N_5647,N_5455);
nor U6513 (N_6513,N_5015,N_5067);
xor U6514 (N_6514,N_5370,N_5440);
or U6515 (N_6515,N_5196,N_4936);
nand U6516 (N_6516,N_4956,N_5471);
nor U6517 (N_6517,N_5281,N_5134);
xnor U6518 (N_6518,N_5345,N_4998);
xnor U6519 (N_6519,N_5236,N_4877);
xor U6520 (N_6520,N_5438,N_5672);
nor U6521 (N_6521,N_4884,N_5743);
or U6522 (N_6522,N_5412,N_5377);
xnor U6523 (N_6523,N_5974,N_5977);
xor U6524 (N_6524,N_5149,N_5859);
xnor U6525 (N_6525,N_5874,N_5635);
xor U6526 (N_6526,N_4968,N_5431);
and U6527 (N_6527,N_5162,N_5069);
or U6528 (N_6528,N_5541,N_5251);
or U6529 (N_6529,N_5277,N_4837);
or U6530 (N_6530,N_5982,N_5082);
nand U6531 (N_6531,N_5062,N_5403);
nand U6532 (N_6532,N_4863,N_4973);
xor U6533 (N_6533,N_5268,N_5217);
nor U6534 (N_6534,N_5791,N_4976);
and U6535 (N_6535,N_5693,N_5095);
xnor U6536 (N_6536,N_5142,N_5706);
nand U6537 (N_6537,N_5349,N_5485);
or U6538 (N_6538,N_5573,N_5252);
xnor U6539 (N_6539,N_5122,N_5629);
xnor U6540 (N_6540,N_5623,N_5126);
xor U6541 (N_6541,N_5290,N_5235);
nor U6542 (N_6542,N_5400,N_4818);
and U6543 (N_6543,N_5690,N_5247);
xor U6544 (N_6544,N_5618,N_5029);
nand U6545 (N_6545,N_5437,N_5081);
nand U6546 (N_6546,N_4831,N_5714);
and U6547 (N_6547,N_5782,N_5342);
nand U6548 (N_6548,N_5927,N_5932);
xor U6549 (N_6549,N_5566,N_5762);
nand U6550 (N_6550,N_5519,N_5614);
nand U6551 (N_6551,N_5258,N_4854);
xor U6552 (N_6552,N_5500,N_5341);
or U6553 (N_6553,N_5064,N_5373);
xor U6554 (N_6554,N_5577,N_5466);
nand U6555 (N_6555,N_5832,N_5682);
nor U6556 (N_6556,N_4947,N_5660);
or U6557 (N_6557,N_5675,N_5211);
xor U6558 (N_6558,N_5613,N_5711);
xor U6559 (N_6559,N_5299,N_5426);
nand U6560 (N_6560,N_4978,N_5423);
or U6561 (N_6561,N_4900,N_5028);
and U6562 (N_6562,N_5547,N_5348);
or U6563 (N_6563,N_5940,N_5158);
or U6564 (N_6564,N_5812,N_5393);
nand U6565 (N_6565,N_4916,N_5298);
nor U6566 (N_6566,N_5492,N_5967);
and U6567 (N_6567,N_5096,N_5046);
and U6568 (N_6568,N_5724,N_5489);
and U6569 (N_6569,N_5105,N_5907);
and U6570 (N_6570,N_5527,N_5490);
nor U6571 (N_6571,N_5271,N_4892);
nand U6572 (N_6572,N_5163,N_5727);
nor U6573 (N_6573,N_4882,N_5264);
nor U6574 (N_6574,N_4838,N_5764);
xnor U6575 (N_6575,N_5875,N_5018);
and U6576 (N_6576,N_5288,N_5194);
nand U6577 (N_6577,N_5060,N_5177);
or U6578 (N_6578,N_4903,N_5569);
nor U6579 (N_6579,N_5501,N_5680);
nor U6580 (N_6580,N_5189,N_5313);
or U6581 (N_6581,N_5410,N_4993);
nor U6582 (N_6582,N_5220,N_5739);
and U6583 (N_6583,N_5359,N_5835);
xnor U6584 (N_6584,N_4939,N_5620);
or U6585 (N_6585,N_5776,N_5030);
nor U6586 (N_6586,N_5090,N_4848);
and U6587 (N_6587,N_5662,N_5896);
nand U6588 (N_6588,N_5208,N_5968);
or U6589 (N_6589,N_5164,N_5956);
nand U6590 (N_6590,N_5005,N_5669);
or U6591 (N_6591,N_5272,N_4919);
nand U6592 (N_6592,N_5225,N_5701);
or U6593 (N_6593,N_5642,N_4925);
and U6594 (N_6594,N_5878,N_5699);
and U6595 (N_6595,N_5576,N_5912);
nor U6596 (N_6596,N_5011,N_5093);
nor U6597 (N_6597,N_5337,N_5004);
xnor U6598 (N_6598,N_5115,N_5780);
and U6599 (N_6599,N_5704,N_5259);
xor U6600 (N_6600,N_5309,N_4921);
or U6601 (N_6601,N_5589,N_5563);
nand U6602 (N_6602,N_5186,N_4859);
nor U6603 (N_6603,N_5550,N_5111);
and U6604 (N_6604,N_5688,N_5578);
xor U6605 (N_6605,N_5169,N_4910);
or U6606 (N_6606,N_5372,N_5716);
nor U6607 (N_6607,N_5750,N_5097);
xor U6608 (N_6608,N_5700,N_5566);
xor U6609 (N_6609,N_4975,N_4806);
and U6610 (N_6610,N_5471,N_5869);
and U6611 (N_6611,N_4897,N_4812);
or U6612 (N_6612,N_4905,N_5717);
and U6613 (N_6613,N_5865,N_5511);
or U6614 (N_6614,N_5993,N_5877);
xor U6615 (N_6615,N_4916,N_5863);
or U6616 (N_6616,N_5880,N_5360);
and U6617 (N_6617,N_5463,N_4948);
nand U6618 (N_6618,N_5446,N_5110);
nand U6619 (N_6619,N_5807,N_5448);
xnor U6620 (N_6620,N_5820,N_4965);
nor U6621 (N_6621,N_5388,N_5074);
nand U6622 (N_6622,N_5185,N_5373);
xnor U6623 (N_6623,N_5564,N_5782);
or U6624 (N_6624,N_5864,N_5994);
nor U6625 (N_6625,N_5623,N_5563);
or U6626 (N_6626,N_5589,N_5517);
and U6627 (N_6627,N_5750,N_5224);
or U6628 (N_6628,N_5436,N_5840);
nand U6629 (N_6629,N_5551,N_5490);
xor U6630 (N_6630,N_5025,N_5915);
and U6631 (N_6631,N_5959,N_5804);
xor U6632 (N_6632,N_5126,N_4806);
and U6633 (N_6633,N_5827,N_5906);
or U6634 (N_6634,N_4871,N_5136);
nor U6635 (N_6635,N_5066,N_5266);
and U6636 (N_6636,N_5723,N_4952);
or U6637 (N_6637,N_5665,N_5724);
xnor U6638 (N_6638,N_5339,N_5666);
nand U6639 (N_6639,N_5064,N_5375);
and U6640 (N_6640,N_5159,N_5399);
nor U6641 (N_6641,N_5660,N_5263);
nand U6642 (N_6642,N_5434,N_5920);
xor U6643 (N_6643,N_5820,N_4850);
xor U6644 (N_6644,N_5747,N_5038);
nand U6645 (N_6645,N_5341,N_4885);
and U6646 (N_6646,N_5097,N_5548);
xor U6647 (N_6647,N_5068,N_5992);
xor U6648 (N_6648,N_5348,N_5540);
nand U6649 (N_6649,N_4811,N_4832);
nand U6650 (N_6650,N_5812,N_5870);
and U6651 (N_6651,N_5037,N_5268);
and U6652 (N_6652,N_5952,N_5624);
xnor U6653 (N_6653,N_5118,N_4908);
nor U6654 (N_6654,N_5110,N_5129);
xor U6655 (N_6655,N_5404,N_5574);
and U6656 (N_6656,N_4897,N_5599);
nor U6657 (N_6657,N_5531,N_4956);
nor U6658 (N_6658,N_5175,N_5587);
xor U6659 (N_6659,N_5801,N_5887);
and U6660 (N_6660,N_4819,N_4957);
or U6661 (N_6661,N_4865,N_5805);
nand U6662 (N_6662,N_5599,N_4841);
and U6663 (N_6663,N_5162,N_5748);
nor U6664 (N_6664,N_5969,N_5880);
nor U6665 (N_6665,N_5878,N_5283);
nor U6666 (N_6666,N_4930,N_5950);
and U6667 (N_6667,N_5936,N_5820);
nand U6668 (N_6668,N_5546,N_5861);
or U6669 (N_6669,N_5117,N_5951);
or U6670 (N_6670,N_4847,N_5859);
nor U6671 (N_6671,N_5283,N_5483);
nor U6672 (N_6672,N_5009,N_5171);
nand U6673 (N_6673,N_5650,N_5102);
nor U6674 (N_6674,N_5145,N_5707);
nor U6675 (N_6675,N_5255,N_5912);
nor U6676 (N_6676,N_5174,N_5853);
xnor U6677 (N_6677,N_5557,N_5649);
and U6678 (N_6678,N_5607,N_5960);
nor U6679 (N_6679,N_5732,N_5663);
nand U6680 (N_6680,N_5412,N_4805);
or U6681 (N_6681,N_5265,N_5743);
or U6682 (N_6682,N_4950,N_5801);
nand U6683 (N_6683,N_4830,N_5089);
nor U6684 (N_6684,N_5967,N_5664);
nand U6685 (N_6685,N_5198,N_5059);
nand U6686 (N_6686,N_4955,N_5126);
nor U6687 (N_6687,N_5938,N_5882);
or U6688 (N_6688,N_5524,N_5855);
nor U6689 (N_6689,N_5256,N_5236);
nor U6690 (N_6690,N_5209,N_5842);
nor U6691 (N_6691,N_5376,N_5080);
or U6692 (N_6692,N_5088,N_5076);
and U6693 (N_6693,N_4867,N_5537);
nor U6694 (N_6694,N_5414,N_5508);
nand U6695 (N_6695,N_4816,N_5110);
and U6696 (N_6696,N_5471,N_4833);
or U6697 (N_6697,N_4820,N_5695);
and U6698 (N_6698,N_5402,N_5977);
and U6699 (N_6699,N_5170,N_5303);
xor U6700 (N_6700,N_5147,N_5698);
nor U6701 (N_6701,N_5080,N_5764);
and U6702 (N_6702,N_5058,N_5485);
or U6703 (N_6703,N_5177,N_5758);
nor U6704 (N_6704,N_5935,N_5948);
and U6705 (N_6705,N_5743,N_5226);
or U6706 (N_6706,N_4956,N_5133);
nand U6707 (N_6707,N_5454,N_5674);
nor U6708 (N_6708,N_5688,N_5746);
nand U6709 (N_6709,N_5016,N_5166);
or U6710 (N_6710,N_5978,N_5197);
nor U6711 (N_6711,N_5732,N_4971);
xor U6712 (N_6712,N_5271,N_5562);
or U6713 (N_6713,N_5326,N_5359);
nand U6714 (N_6714,N_4966,N_5288);
nor U6715 (N_6715,N_5048,N_5293);
or U6716 (N_6716,N_5053,N_5099);
and U6717 (N_6717,N_4929,N_5583);
and U6718 (N_6718,N_5627,N_4853);
and U6719 (N_6719,N_4977,N_5055);
or U6720 (N_6720,N_4823,N_5576);
and U6721 (N_6721,N_5496,N_5717);
nand U6722 (N_6722,N_5824,N_4831);
nand U6723 (N_6723,N_5928,N_5771);
nand U6724 (N_6724,N_5176,N_5653);
or U6725 (N_6725,N_5691,N_5606);
nand U6726 (N_6726,N_5387,N_4882);
or U6727 (N_6727,N_5392,N_5291);
nand U6728 (N_6728,N_5957,N_5233);
nand U6729 (N_6729,N_5221,N_5907);
or U6730 (N_6730,N_5957,N_5604);
or U6731 (N_6731,N_5424,N_5723);
nand U6732 (N_6732,N_5253,N_5182);
xor U6733 (N_6733,N_5276,N_5047);
or U6734 (N_6734,N_5091,N_5074);
nor U6735 (N_6735,N_5583,N_5870);
xnor U6736 (N_6736,N_4819,N_5865);
or U6737 (N_6737,N_5549,N_5620);
and U6738 (N_6738,N_5656,N_4927);
nand U6739 (N_6739,N_5915,N_5880);
or U6740 (N_6740,N_5171,N_4905);
nand U6741 (N_6741,N_5752,N_5882);
xnor U6742 (N_6742,N_5682,N_5711);
and U6743 (N_6743,N_5325,N_4893);
or U6744 (N_6744,N_5252,N_5249);
nand U6745 (N_6745,N_5237,N_4927);
xnor U6746 (N_6746,N_5650,N_5653);
or U6747 (N_6747,N_4989,N_5209);
and U6748 (N_6748,N_5140,N_5117);
nor U6749 (N_6749,N_4871,N_5763);
nor U6750 (N_6750,N_5638,N_5903);
and U6751 (N_6751,N_5888,N_5936);
xor U6752 (N_6752,N_5766,N_5862);
or U6753 (N_6753,N_5077,N_5775);
nand U6754 (N_6754,N_5603,N_5218);
xor U6755 (N_6755,N_5372,N_5701);
nand U6756 (N_6756,N_5565,N_5399);
nor U6757 (N_6757,N_4978,N_5092);
nand U6758 (N_6758,N_5662,N_5408);
nand U6759 (N_6759,N_5583,N_5398);
xor U6760 (N_6760,N_5624,N_5429);
nor U6761 (N_6761,N_5807,N_4938);
and U6762 (N_6762,N_5989,N_4958);
or U6763 (N_6763,N_5136,N_5678);
or U6764 (N_6764,N_5154,N_5807);
and U6765 (N_6765,N_5160,N_5186);
or U6766 (N_6766,N_5452,N_4975);
and U6767 (N_6767,N_5390,N_4910);
and U6768 (N_6768,N_5779,N_4999);
and U6769 (N_6769,N_5076,N_5189);
xnor U6770 (N_6770,N_5599,N_5370);
nand U6771 (N_6771,N_4931,N_5816);
or U6772 (N_6772,N_5029,N_4983);
nand U6773 (N_6773,N_5566,N_5988);
and U6774 (N_6774,N_5871,N_5415);
or U6775 (N_6775,N_5949,N_5497);
and U6776 (N_6776,N_5155,N_5008);
and U6777 (N_6777,N_4921,N_5719);
or U6778 (N_6778,N_5567,N_5584);
xnor U6779 (N_6779,N_5016,N_5658);
xor U6780 (N_6780,N_5135,N_5166);
or U6781 (N_6781,N_5509,N_5828);
xnor U6782 (N_6782,N_5892,N_5355);
nor U6783 (N_6783,N_5221,N_5692);
nand U6784 (N_6784,N_4966,N_5865);
nor U6785 (N_6785,N_5620,N_5072);
or U6786 (N_6786,N_5042,N_5252);
nor U6787 (N_6787,N_5011,N_5998);
nor U6788 (N_6788,N_5489,N_5936);
nor U6789 (N_6789,N_5543,N_5591);
xor U6790 (N_6790,N_5438,N_5203);
xor U6791 (N_6791,N_5873,N_5143);
or U6792 (N_6792,N_4868,N_4936);
xor U6793 (N_6793,N_4943,N_5730);
or U6794 (N_6794,N_5010,N_5311);
or U6795 (N_6795,N_5398,N_4804);
xnor U6796 (N_6796,N_5459,N_5348);
and U6797 (N_6797,N_5860,N_5227);
and U6798 (N_6798,N_5953,N_5020);
xnor U6799 (N_6799,N_4938,N_5520);
and U6800 (N_6800,N_4952,N_5581);
and U6801 (N_6801,N_5851,N_5811);
nand U6802 (N_6802,N_5039,N_5546);
nand U6803 (N_6803,N_5144,N_5369);
and U6804 (N_6804,N_5068,N_5264);
xnor U6805 (N_6805,N_5796,N_5842);
nor U6806 (N_6806,N_5061,N_5489);
xor U6807 (N_6807,N_4820,N_4984);
nor U6808 (N_6808,N_5718,N_5260);
or U6809 (N_6809,N_5328,N_5249);
and U6810 (N_6810,N_5741,N_4813);
xor U6811 (N_6811,N_5970,N_5001);
nand U6812 (N_6812,N_4929,N_5054);
and U6813 (N_6813,N_5889,N_5876);
xor U6814 (N_6814,N_5721,N_5957);
and U6815 (N_6815,N_5691,N_4893);
or U6816 (N_6816,N_4977,N_4904);
or U6817 (N_6817,N_5199,N_5495);
nand U6818 (N_6818,N_4972,N_5432);
nor U6819 (N_6819,N_5203,N_4925);
nand U6820 (N_6820,N_5392,N_5209);
and U6821 (N_6821,N_5359,N_5275);
nand U6822 (N_6822,N_5446,N_5910);
nand U6823 (N_6823,N_5235,N_5755);
nand U6824 (N_6824,N_5613,N_4835);
xor U6825 (N_6825,N_5051,N_5529);
xor U6826 (N_6826,N_5429,N_5096);
nand U6827 (N_6827,N_5973,N_5674);
xnor U6828 (N_6828,N_5488,N_4808);
or U6829 (N_6829,N_5942,N_5922);
xnor U6830 (N_6830,N_4975,N_5665);
and U6831 (N_6831,N_4828,N_4818);
nand U6832 (N_6832,N_5930,N_5141);
and U6833 (N_6833,N_5878,N_4924);
nand U6834 (N_6834,N_5460,N_5641);
or U6835 (N_6835,N_5767,N_5276);
nand U6836 (N_6836,N_5004,N_5548);
nor U6837 (N_6837,N_5883,N_5517);
xor U6838 (N_6838,N_4819,N_5775);
nor U6839 (N_6839,N_5838,N_4902);
nand U6840 (N_6840,N_5514,N_5125);
xnor U6841 (N_6841,N_5206,N_4943);
nand U6842 (N_6842,N_5969,N_5038);
and U6843 (N_6843,N_5392,N_4985);
xor U6844 (N_6844,N_5160,N_5533);
or U6845 (N_6845,N_5770,N_4856);
and U6846 (N_6846,N_5872,N_5003);
nor U6847 (N_6847,N_5814,N_5891);
nor U6848 (N_6848,N_4892,N_5916);
nor U6849 (N_6849,N_4938,N_5358);
nor U6850 (N_6850,N_4807,N_5817);
nand U6851 (N_6851,N_5347,N_5108);
nand U6852 (N_6852,N_5651,N_5302);
or U6853 (N_6853,N_5340,N_5934);
nor U6854 (N_6854,N_5308,N_5300);
nor U6855 (N_6855,N_5697,N_5773);
nor U6856 (N_6856,N_5231,N_5702);
xor U6857 (N_6857,N_5975,N_5740);
or U6858 (N_6858,N_5896,N_5968);
nor U6859 (N_6859,N_4856,N_5453);
xor U6860 (N_6860,N_5315,N_5494);
or U6861 (N_6861,N_5933,N_5970);
and U6862 (N_6862,N_5719,N_5178);
or U6863 (N_6863,N_5587,N_5217);
nor U6864 (N_6864,N_5117,N_5770);
nor U6865 (N_6865,N_5583,N_5840);
nand U6866 (N_6866,N_5433,N_5084);
nand U6867 (N_6867,N_4885,N_4831);
nor U6868 (N_6868,N_5024,N_5596);
xor U6869 (N_6869,N_5867,N_5975);
nor U6870 (N_6870,N_5295,N_5175);
or U6871 (N_6871,N_5108,N_4889);
nor U6872 (N_6872,N_4987,N_5535);
xnor U6873 (N_6873,N_4897,N_5672);
xor U6874 (N_6874,N_4955,N_4879);
and U6875 (N_6875,N_5133,N_5367);
nand U6876 (N_6876,N_5319,N_5850);
nand U6877 (N_6877,N_5432,N_5849);
nand U6878 (N_6878,N_5008,N_5998);
xor U6879 (N_6879,N_5278,N_4910);
or U6880 (N_6880,N_5908,N_5485);
and U6881 (N_6881,N_5916,N_5773);
nand U6882 (N_6882,N_5161,N_5866);
xnor U6883 (N_6883,N_5810,N_4948);
and U6884 (N_6884,N_5160,N_5018);
or U6885 (N_6885,N_5989,N_5832);
nand U6886 (N_6886,N_5795,N_5432);
xor U6887 (N_6887,N_4838,N_5369);
and U6888 (N_6888,N_4987,N_5916);
or U6889 (N_6889,N_4920,N_5409);
xnor U6890 (N_6890,N_5637,N_5590);
or U6891 (N_6891,N_5185,N_5812);
nand U6892 (N_6892,N_4800,N_5706);
nor U6893 (N_6893,N_5976,N_5047);
xnor U6894 (N_6894,N_5714,N_5639);
xor U6895 (N_6895,N_4841,N_5987);
nand U6896 (N_6896,N_5872,N_5473);
or U6897 (N_6897,N_5146,N_5699);
nand U6898 (N_6898,N_5940,N_4907);
nand U6899 (N_6899,N_5810,N_5441);
xor U6900 (N_6900,N_5582,N_5329);
or U6901 (N_6901,N_5414,N_5956);
nor U6902 (N_6902,N_5561,N_5361);
nand U6903 (N_6903,N_5414,N_5142);
xnor U6904 (N_6904,N_5596,N_5379);
xnor U6905 (N_6905,N_5094,N_5737);
nor U6906 (N_6906,N_5827,N_5976);
xor U6907 (N_6907,N_5421,N_5074);
xnor U6908 (N_6908,N_5275,N_5471);
nand U6909 (N_6909,N_5266,N_5082);
xor U6910 (N_6910,N_5750,N_4815);
or U6911 (N_6911,N_5287,N_4827);
xor U6912 (N_6912,N_5840,N_5190);
and U6913 (N_6913,N_5767,N_5536);
nor U6914 (N_6914,N_5305,N_4863);
nand U6915 (N_6915,N_4879,N_5377);
nand U6916 (N_6916,N_5152,N_5393);
or U6917 (N_6917,N_5131,N_5391);
nand U6918 (N_6918,N_5495,N_5985);
nor U6919 (N_6919,N_5239,N_5554);
or U6920 (N_6920,N_5500,N_5397);
xnor U6921 (N_6921,N_5144,N_5547);
nor U6922 (N_6922,N_4938,N_5896);
xor U6923 (N_6923,N_5530,N_5955);
nor U6924 (N_6924,N_5128,N_5825);
nand U6925 (N_6925,N_5787,N_5073);
or U6926 (N_6926,N_5937,N_5686);
nor U6927 (N_6927,N_4996,N_5569);
nand U6928 (N_6928,N_5127,N_5073);
nor U6929 (N_6929,N_5431,N_5525);
xnor U6930 (N_6930,N_5580,N_5502);
xor U6931 (N_6931,N_5123,N_5790);
or U6932 (N_6932,N_5224,N_4835);
nand U6933 (N_6933,N_5324,N_5395);
and U6934 (N_6934,N_5744,N_5894);
xor U6935 (N_6935,N_5406,N_5353);
nand U6936 (N_6936,N_5455,N_4848);
or U6937 (N_6937,N_5973,N_5170);
nor U6938 (N_6938,N_5728,N_5246);
xor U6939 (N_6939,N_5783,N_4975);
and U6940 (N_6940,N_5803,N_5122);
and U6941 (N_6941,N_4841,N_5036);
xnor U6942 (N_6942,N_5998,N_5597);
and U6943 (N_6943,N_5641,N_5339);
and U6944 (N_6944,N_5709,N_4862);
or U6945 (N_6945,N_5408,N_5942);
xnor U6946 (N_6946,N_4838,N_5749);
nand U6947 (N_6947,N_5762,N_5564);
or U6948 (N_6948,N_4837,N_4868);
nand U6949 (N_6949,N_5560,N_4881);
xnor U6950 (N_6950,N_5753,N_5650);
xor U6951 (N_6951,N_5448,N_5053);
or U6952 (N_6952,N_5884,N_4933);
or U6953 (N_6953,N_5226,N_5789);
nand U6954 (N_6954,N_5454,N_5013);
nor U6955 (N_6955,N_5121,N_5895);
xor U6956 (N_6956,N_4936,N_5139);
or U6957 (N_6957,N_5501,N_5767);
xnor U6958 (N_6958,N_5189,N_5297);
xor U6959 (N_6959,N_5808,N_5135);
nand U6960 (N_6960,N_5154,N_5021);
nor U6961 (N_6961,N_5201,N_5231);
or U6962 (N_6962,N_5812,N_5201);
xnor U6963 (N_6963,N_5040,N_5589);
or U6964 (N_6964,N_5552,N_4961);
nand U6965 (N_6965,N_5028,N_5682);
nor U6966 (N_6966,N_5869,N_5787);
and U6967 (N_6967,N_5811,N_5552);
xnor U6968 (N_6968,N_5633,N_5416);
xor U6969 (N_6969,N_5869,N_5831);
or U6970 (N_6970,N_5321,N_5894);
or U6971 (N_6971,N_4911,N_5658);
and U6972 (N_6972,N_5551,N_4823);
nand U6973 (N_6973,N_5247,N_5559);
xnor U6974 (N_6974,N_5012,N_5051);
nor U6975 (N_6975,N_5807,N_5647);
or U6976 (N_6976,N_5783,N_5789);
nand U6977 (N_6977,N_5235,N_5912);
or U6978 (N_6978,N_5400,N_5074);
nand U6979 (N_6979,N_5929,N_5243);
or U6980 (N_6980,N_4970,N_5116);
and U6981 (N_6981,N_5929,N_5246);
xor U6982 (N_6982,N_5994,N_5112);
or U6983 (N_6983,N_5292,N_5753);
nand U6984 (N_6984,N_5555,N_5656);
or U6985 (N_6985,N_5088,N_4902);
and U6986 (N_6986,N_5657,N_5695);
nor U6987 (N_6987,N_5523,N_5995);
nor U6988 (N_6988,N_5830,N_5942);
nand U6989 (N_6989,N_5949,N_5456);
xnor U6990 (N_6990,N_5111,N_5594);
and U6991 (N_6991,N_5519,N_5664);
nand U6992 (N_6992,N_5314,N_5415);
or U6993 (N_6993,N_5749,N_5159);
xnor U6994 (N_6994,N_5770,N_5465);
nand U6995 (N_6995,N_5125,N_4931);
nand U6996 (N_6996,N_5208,N_5329);
xor U6997 (N_6997,N_5812,N_5694);
nor U6998 (N_6998,N_4850,N_5586);
and U6999 (N_6999,N_5171,N_5578);
nor U7000 (N_7000,N_5844,N_5369);
and U7001 (N_7001,N_5569,N_5078);
nand U7002 (N_7002,N_5195,N_5532);
and U7003 (N_7003,N_5232,N_5887);
or U7004 (N_7004,N_5647,N_5563);
and U7005 (N_7005,N_5165,N_4971);
and U7006 (N_7006,N_4839,N_5827);
and U7007 (N_7007,N_5864,N_5023);
nand U7008 (N_7008,N_5558,N_5597);
and U7009 (N_7009,N_5169,N_4895);
or U7010 (N_7010,N_5520,N_5906);
nor U7011 (N_7011,N_5526,N_5859);
nand U7012 (N_7012,N_4998,N_5240);
and U7013 (N_7013,N_4868,N_5181);
nor U7014 (N_7014,N_5091,N_4899);
nand U7015 (N_7015,N_4900,N_5876);
nand U7016 (N_7016,N_5838,N_4927);
and U7017 (N_7017,N_5170,N_5001);
nand U7018 (N_7018,N_5872,N_5236);
and U7019 (N_7019,N_4898,N_5785);
and U7020 (N_7020,N_4800,N_4945);
or U7021 (N_7021,N_5387,N_4947);
nor U7022 (N_7022,N_5537,N_5847);
xor U7023 (N_7023,N_5834,N_5381);
or U7024 (N_7024,N_5430,N_5457);
or U7025 (N_7025,N_5175,N_5475);
nor U7026 (N_7026,N_5696,N_5961);
or U7027 (N_7027,N_5302,N_5856);
xor U7028 (N_7028,N_4956,N_4983);
nor U7029 (N_7029,N_5259,N_5399);
nor U7030 (N_7030,N_5778,N_4843);
and U7031 (N_7031,N_5844,N_4926);
nand U7032 (N_7032,N_5823,N_5571);
and U7033 (N_7033,N_4943,N_5811);
and U7034 (N_7034,N_5575,N_5113);
nand U7035 (N_7035,N_5761,N_5393);
nor U7036 (N_7036,N_5427,N_5909);
xor U7037 (N_7037,N_4957,N_5866);
xor U7038 (N_7038,N_5660,N_5631);
xnor U7039 (N_7039,N_5778,N_5678);
or U7040 (N_7040,N_5439,N_5429);
xor U7041 (N_7041,N_4846,N_5797);
or U7042 (N_7042,N_5128,N_5833);
nor U7043 (N_7043,N_5520,N_5803);
xor U7044 (N_7044,N_5181,N_5324);
xor U7045 (N_7045,N_5582,N_5127);
xor U7046 (N_7046,N_4866,N_5978);
nor U7047 (N_7047,N_5089,N_5231);
nand U7048 (N_7048,N_5483,N_5472);
nor U7049 (N_7049,N_5203,N_5940);
nand U7050 (N_7050,N_4841,N_5956);
xnor U7051 (N_7051,N_5008,N_5588);
and U7052 (N_7052,N_5820,N_4990);
nand U7053 (N_7053,N_5193,N_5577);
nor U7054 (N_7054,N_5162,N_5461);
nand U7055 (N_7055,N_5176,N_4901);
nand U7056 (N_7056,N_5738,N_5227);
and U7057 (N_7057,N_5684,N_5870);
xnor U7058 (N_7058,N_5476,N_5356);
and U7059 (N_7059,N_5659,N_5737);
and U7060 (N_7060,N_4841,N_5054);
xnor U7061 (N_7061,N_5449,N_4841);
and U7062 (N_7062,N_5646,N_5178);
nand U7063 (N_7063,N_5611,N_5633);
nor U7064 (N_7064,N_5143,N_5447);
nand U7065 (N_7065,N_4811,N_5574);
and U7066 (N_7066,N_5781,N_4938);
nor U7067 (N_7067,N_5145,N_5579);
xnor U7068 (N_7068,N_5096,N_5568);
nor U7069 (N_7069,N_5304,N_4850);
xnor U7070 (N_7070,N_5837,N_5610);
or U7071 (N_7071,N_5578,N_5598);
or U7072 (N_7072,N_4952,N_5778);
and U7073 (N_7073,N_5317,N_5363);
nand U7074 (N_7074,N_5361,N_5603);
nand U7075 (N_7075,N_5058,N_5373);
xnor U7076 (N_7076,N_5985,N_5930);
nand U7077 (N_7077,N_5627,N_5680);
nand U7078 (N_7078,N_5439,N_5604);
or U7079 (N_7079,N_5708,N_5071);
or U7080 (N_7080,N_5501,N_5374);
nand U7081 (N_7081,N_5105,N_5128);
and U7082 (N_7082,N_4843,N_5629);
xor U7083 (N_7083,N_5467,N_5014);
xor U7084 (N_7084,N_5113,N_5026);
nor U7085 (N_7085,N_5364,N_5192);
nor U7086 (N_7086,N_5675,N_5462);
nand U7087 (N_7087,N_5469,N_5866);
nor U7088 (N_7088,N_5763,N_5052);
and U7089 (N_7089,N_5278,N_5273);
or U7090 (N_7090,N_5421,N_4885);
nand U7091 (N_7091,N_5823,N_5595);
nor U7092 (N_7092,N_5538,N_4833);
and U7093 (N_7093,N_5796,N_5740);
or U7094 (N_7094,N_5642,N_4970);
nor U7095 (N_7095,N_5553,N_5633);
xor U7096 (N_7096,N_4935,N_5310);
nor U7097 (N_7097,N_5052,N_5344);
nand U7098 (N_7098,N_5064,N_5518);
xnor U7099 (N_7099,N_5626,N_5288);
xnor U7100 (N_7100,N_5660,N_5361);
xor U7101 (N_7101,N_5701,N_5944);
nand U7102 (N_7102,N_5836,N_5549);
nand U7103 (N_7103,N_5225,N_5911);
or U7104 (N_7104,N_5872,N_5160);
or U7105 (N_7105,N_5683,N_5823);
and U7106 (N_7106,N_5783,N_4932);
or U7107 (N_7107,N_5398,N_5516);
and U7108 (N_7108,N_5220,N_5025);
xnor U7109 (N_7109,N_5096,N_5194);
xor U7110 (N_7110,N_5278,N_5263);
or U7111 (N_7111,N_5427,N_5833);
nand U7112 (N_7112,N_5446,N_4966);
nor U7113 (N_7113,N_5834,N_5291);
xor U7114 (N_7114,N_5095,N_5857);
and U7115 (N_7115,N_5879,N_4993);
and U7116 (N_7116,N_5697,N_5799);
xor U7117 (N_7117,N_5331,N_5842);
nand U7118 (N_7118,N_5959,N_5716);
xor U7119 (N_7119,N_5473,N_5954);
or U7120 (N_7120,N_5431,N_4912);
nand U7121 (N_7121,N_4946,N_5087);
nor U7122 (N_7122,N_5789,N_4972);
and U7123 (N_7123,N_4851,N_5946);
nand U7124 (N_7124,N_5144,N_4825);
nand U7125 (N_7125,N_5629,N_5369);
xnor U7126 (N_7126,N_5090,N_5598);
xor U7127 (N_7127,N_5253,N_5500);
xor U7128 (N_7128,N_5861,N_5236);
nand U7129 (N_7129,N_5726,N_4913);
xor U7130 (N_7130,N_5617,N_4983);
xor U7131 (N_7131,N_5607,N_5201);
nor U7132 (N_7132,N_5401,N_5090);
nor U7133 (N_7133,N_4983,N_5230);
nor U7134 (N_7134,N_5630,N_5292);
xnor U7135 (N_7135,N_5502,N_5521);
or U7136 (N_7136,N_5767,N_4843);
nand U7137 (N_7137,N_5496,N_5844);
and U7138 (N_7138,N_5362,N_5963);
nor U7139 (N_7139,N_5846,N_5522);
or U7140 (N_7140,N_5741,N_5461);
nand U7141 (N_7141,N_5925,N_5607);
and U7142 (N_7142,N_5677,N_5242);
or U7143 (N_7143,N_5788,N_5487);
or U7144 (N_7144,N_4877,N_5427);
nor U7145 (N_7145,N_5374,N_5836);
or U7146 (N_7146,N_5365,N_5911);
nand U7147 (N_7147,N_5320,N_5541);
nand U7148 (N_7148,N_5647,N_5823);
xor U7149 (N_7149,N_5813,N_5576);
and U7150 (N_7150,N_4942,N_5390);
or U7151 (N_7151,N_5748,N_5772);
nand U7152 (N_7152,N_5536,N_5941);
nor U7153 (N_7153,N_5696,N_5759);
xor U7154 (N_7154,N_5445,N_5877);
and U7155 (N_7155,N_4824,N_5714);
nor U7156 (N_7156,N_5213,N_5289);
nor U7157 (N_7157,N_5128,N_5210);
nand U7158 (N_7158,N_5648,N_5642);
and U7159 (N_7159,N_5993,N_5867);
nor U7160 (N_7160,N_5470,N_5782);
nand U7161 (N_7161,N_5227,N_4844);
xor U7162 (N_7162,N_5673,N_5838);
nor U7163 (N_7163,N_5869,N_5822);
xor U7164 (N_7164,N_5698,N_5953);
nor U7165 (N_7165,N_5902,N_5409);
nor U7166 (N_7166,N_5974,N_5583);
or U7167 (N_7167,N_4982,N_5743);
nand U7168 (N_7168,N_5371,N_5889);
or U7169 (N_7169,N_5472,N_5555);
nor U7170 (N_7170,N_5982,N_4862);
xnor U7171 (N_7171,N_5864,N_5435);
nor U7172 (N_7172,N_4934,N_5101);
or U7173 (N_7173,N_5781,N_5398);
or U7174 (N_7174,N_5803,N_5172);
nor U7175 (N_7175,N_5223,N_4934);
or U7176 (N_7176,N_5918,N_5019);
nor U7177 (N_7177,N_4970,N_5037);
or U7178 (N_7178,N_5219,N_5694);
nand U7179 (N_7179,N_5842,N_5269);
nor U7180 (N_7180,N_5117,N_5722);
nand U7181 (N_7181,N_5550,N_4808);
and U7182 (N_7182,N_5062,N_5282);
or U7183 (N_7183,N_5099,N_5874);
nand U7184 (N_7184,N_4998,N_4828);
nor U7185 (N_7185,N_5335,N_5584);
nor U7186 (N_7186,N_5253,N_5697);
xnor U7187 (N_7187,N_5538,N_5850);
nand U7188 (N_7188,N_5035,N_5330);
nor U7189 (N_7189,N_5050,N_5820);
and U7190 (N_7190,N_4841,N_5796);
and U7191 (N_7191,N_5135,N_4839);
nand U7192 (N_7192,N_5766,N_5637);
nand U7193 (N_7193,N_4989,N_5773);
and U7194 (N_7194,N_5796,N_4993);
or U7195 (N_7195,N_5429,N_5639);
nor U7196 (N_7196,N_5324,N_5722);
and U7197 (N_7197,N_5611,N_4800);
or U7198 (N_7198,N_4903,N_5799);
and U7199 (N_7199,N_5026,N_5885);
or U7200 (N_7200,N_7144,N_6825);
and U7201 (N_7201,N_6272,N_6288);
nor U7202 (N_7202,N_6932,N_6560);
or U7203 (N_7203,N_6928,N_6279);
nand U7204 (N_7204,N_6236,N_7030);
nor U7205 (N_7205,N_6814,N_6681);
nand U7206 (N_7206,N_6062,N_7063);
nor U7207 (N_7207,N_6790,N_6353);
and U7208 (N_7208,N_6076,N_7077);
and U7209 (N_7209,N_6225,N_7037);
or U7210 (N_7210,N_6401,N_6386);
nand U7211 (N_7211,N_6499,N_6303);
xor U7212 (N_7212,N_6100,N_6801);
or U7213 (N_7213,N_6833,N_6508);
nor U7214 (N_7214,N_6090,N_6187);
nand U7215 (N_7215,N_6041,N_7059);
or U7216 (N_7216,N_6102,N_6006);
and U7217 (N_7217,N_6764,N_6421);
nand U7218 (N_7218,N_6275,N_6974);
and U7219 (N_7219,N_6605,N_6824);
nor U7220 (N_7220,N_6648,N_6603);
or U7221 (N_7221,N_6740,N_6715);
or U7222 (N_7222,N_6767,N_6134);
xnor U7223 (N_7223,N_6354,N_6741);
nor U7224 (N_7224,N_6630,N_6297);
nand U7225 (N_7225,N_6578,N_6761);
xnor U7226 (N_7226,N_6523,N_6862);
and U7227 (N_7227,N_6116,N_7107);
and U7228 (N_7228,N_7174,N_7060);
xnor U7229 (N_7229,N_7054,N_6773);
nand U7230 (N_7230,N_6299,N_6185);
nand U7231 (N_7231,N_6848,N_6846);
nor U7232 (N_7232,N_6856,N_6398);
xor U7233 (N_7233,N_6947,N_6491);
nor U7234 (N_7234,N_6680,N_6336);
nor U7235 (N_7235,N_6831,N_6751);
and U7236 (N_7236,N_6598,N_6970);
or U7237 (N_7237,N_6564,N_6613);
xor U7238 (N_7238,N_6488,N_6362);
xor U7239 (N_7239,N_6101,N_6584);
xor U7240 (N_7240,N_6614,N_6432);
xnor U7241 (N_7241,N_6670,N_6069);
or U7242 (N_7242,N_6192,N_6416);
nor U7243 (N_7243,N_6057,N_6829);
nor U7244 (N_7244,N_6092,N_6608);
and U7245 (N_7245,N_6391,N_6794);
nor U7246 (N_7246,N_6513,N_6157);
and U7247 (N_7247,N_6669,N_6782);
or U7248 (N_7248,N_6242,N_6471);
and U7249 (N_7249,N_6325,N_6817);
xnor U7250 (N_7250,N_6477,N_7116);
nand U7251 (N_7251,N_6066,N_6646);
nor U7252 (N_7252,N_6440,N_7162);
or U7253 (N_7253,N_6379,N_6286);
xnor U7254 (N_7254,N_6063,N_7129);
nor U7255 (N_7255,N_6469,N_6688);
or U7256 (N_7256,N_6395,N_6196);
or U7257 (N_7257,N_6533,N_6504);
xnor U7258 (N_7258,N_6726,N_6166);
xor U7259 (N_7259,N_6203,N_6755);
nand U7260 (N_7260,N_6459,N_6569);
xor U7261 (N_7261,N_6691,N_6312);
or U7262 (N_7262,N_6855,N_6453);
nand U7263 (N_7263,N_6505,N_7148);
or U7264 (N_7264,N_6546,N_6094);
or U7265 (N_7265,N_6418,N_6800);
xor U7266 (N_7266,N_7120,N_6992);
xor U7267 (N_7267,N_6510,N_6624);
and U7268 (N_7268,N_7135,N_6022);
and U7269 (N_7269,N_6036,N_7114);
xor U7270 (N_7270,N_6876,N_6132);
xor U7271 (N_7271,N_6583,N_6599);
nor U7272 (N_7272,N_6254,N_6672);
and U7273 (N_7273,N_6202,N_7051);
xnor U7274 (N_7274,N_6543,N_6350);
xor U7275 (N_7275,N_7076,N_7078);
xor U7276 (N_7276,N_6650,N_6280);
or U7277 (N_7277,N_6870,N_6382);
and U7278 (N_7278,N_6285,N_6184);
and U7279 (N_7279,N_6219,N_7069);
nand U7280 (N_7280,N_6808,N_7040);
and U7281 (N_7281,N_6534,N_6333);
nand U7282 (N_7282,N_6934,N_7007);
nand U7283 (N_7283,N_6218,N_6926);
nand U7284 (N_7284,N_6212,N_7156);
nand U7285 (N_7285,N_6798,N_6204);
xor U7286 (N_7286,N_6082,N_6557);
and U7287 (N_7287,N_6052,N_6430);
xnor U7288 (N_7288,N_6652,N_6905);
nor U7289 (N_7289,N_6492,N_6699);
nand U7290 (N_7290,N_6540,N_6109);
nand U7291 (N_7291,N_6776,N_6832);
or U7292 (N_7292,N_6438,N_6886);
or U7293 (N_7293,N_6037,N_6337);
or U7294 (N_7294,N_6836,N_6916);
nand U7295 (N_7295,N_7191,N_7150);
nand U7296 (N_7296,N_6284,N_6189);
nor U7297 (N_7297,N_6732,N_6592);
xnor U7298 (N_7298,N_6507,N_6664);
nor U7299 (N_7299,N_6908,N_6526);
and U7300 (N_7300,N_6446,N_6892);
or U7301 (N_7301,N_6125,N_7009);
or U7302 (N_7302,N_6347,N_6002);
xor U7303 (N_7303,N_6207,N_6251);
nand U7304 (N_7304,N_6072,N_7016);
or U7305 (N_7305,N_6977,N_6525);
nand U7306 (N_7306,N_6611,N_6305);
and U7307 (N_7307,N_6826,N_6739);
nor U7308 (N_7308,N_7153,N_7021);
nand U7309 (N_7309,N_6497,N_6146);
nand U7310 (N_7310,N_6019,N_6566);
nand U7311 (N_7311,N_6213,N_6475);
xor U7312 (N_7312,N_7112,N_6186);
or U7313 (N_7313,N_6058,N_6230);
xnor U7314 (N_7314,N_6873,N_6768);
nand U7315 (N_7315,N_6665,N_6287);
xor U7316 (N_7316,N_6657,N_7055);
and U7317 (N_7317,N_6896,N_6946);
or U7318 (N_7318,N_7095,N_6858);
nand U7319 (N_7319,N_6594,N_6793);
nand U7320 (N_7320,N_6729,N_6404);
and U7321 (N_7321,N_6633,N_7041);
nand U7322 (N_7322,N_6442,N_6127);
or U7323 (N_7323,N_7057,N_7090);
xor U7324 (N_7324,N_6294,N_6621);
xnor U7325 (N_7325,N_6123,N_6509);
xor U7326 (N_7326,N_6241,N_6344);
or U7327 (N_7327,N_6417,N_6685);
nand U7328 (N_7328,N_6248,N_6035);
or U7329 (N_7329,N_6194,N_7137);
nand U7330 (N_7330,N_6056,N_6983);
nand U7331 (N_7331,N_6496,N_6677);
nor U7332 (N_7332,N_7047,N_6411);
and U7333 (N_7333,N_6004,N_6874);
nor U7334 (N_7334,N_6638,N_7071);
nand U7335 (N_7335,N_6880,N_6269);
nor U7336 (N_7336,N_6419,N_6465);
nor U7337 (N_7337,N_7104,N_6554);
or U7338 (N_7338,N_6747,N_6744);
xnor U7339 (N_7339,N_6175,N_6990);
xor U7340 (N_7340,N_6589,N_6257);
or U7341 (N_7341,N_6223,N_6812);
nor U7342 (N_7342,N_6885,N_7158);
nand U7343 (N_7343,N_7046,N_6541);
nand U7344 (N_7344,N_7151,N_6178);
nand U7345 (N_7345,N_7093,N_6228);
or U7346 (N_7346,N_6520,N_6324);
xnor U7347 (N_7347,N_6698,N_6258);
nor U7348 (N_7348,N_7119,N_7123);
nand U7349 (N_7349,N_6697,N_6647);
or U7350 (N_7350,N_6769,N_6070);
nor U7351 (N_7351,N_6360,N_6054);
or U7352 (N_7352,N_7159,N_7160);
xor U7353 (N_7353,N_6470,N_6635);
xor U7354 (N_7354,N_7102,N_6718);
nor U7355 (N_7355,N_6881,N_6179);
and U7356 (N_7356,N_6122,N_6821);
nor U7357 (N_7357,N_7115,N_6130);
nor U7358 (N_7358,N_6780,N_6850);
nand U7359 (N_7359,N_6849,N_6791);
nand U7360 (N_7360,N_6595,N_6075);
nand U7361 (N_7361,N_6950,N_6436);
xnor U7362 (N_7362,N_6556,N_6707);
nand U7363 (N_7363,N_6834,N_6724);
nand U7364 (N_7364,N_6443,N_6674);
or U7365 (N_7365,N_7122,N_6345);
xnor U7366 (N_7366,N_6064,N_6910);
or U7367 (N_7367,N_6572,N_6933);
nor U7368 (N_7368,N_7070,N_6893);
nand U7369 (N_7369,N_6609,N_6129);
or U7370 (N_7370,N_6167,N_6579);
xnor U7371 (N_7371,N_6806,N_6570);
xor U7372 (N_7372,N_6811,N_6679);
and U7373 (N_7373,N_6281,N_7117);
and U7374 (N_7374,N_6495,N_6632);
nor U7375 (N_7375,N_6091,N_6847);
and U7376 (N_7376,N_6040,N_6224);
nor U7377 (N_7377,N_6937,N_6183);
nor U7378 (N_7378,N_7183,N_6607);
and U7379 (N_7379,N_6929,N_6588);
nor U7380 (N_7380,N_6061,N_6593);
or U7381 (N_7381,N_6760,N_7029);
xnor U7382 (N_7382,N_6431,N_6323);
xnor U7383 (N_7383,N_6144,N_6696);
and U7384 (N_7384,N_7126,N_6877);
nand U7385 (N_7385,N_6898,N_6027);
and U7386 (N_7386,N_6244,N_6689);
nand U7387 (N_7387,N_6645,N_6340);
nor U7388 (N_7388,N_7085,N_6988);
xnor U7389 (N_7389,N_6349,N_7161);
nand U7390 (N_7390,N_7170,N_6270);
xnor U7391 (N_7391,N_6625,N_6433);
and U7392 (N_7392,N_6278,N_6200);
and U7393 (N_7393,N_6482,N_6103);
nor U7394 (N_7394,N_6169,N_6531);
xnor U7395 (N_7395,N_6128,N_6126);
and U7396 (N_7396,N_6924,N_6086);
or U7397 (N_7397,N_6799,N_6558);
xor U7398 (N_7398,N_6034,N_6766);
or U7399 (N_7399,N_7023,N_6455);
xor U7400 (N_7400,N_6752,N_6666);
and U7401 (N_7401,N_6919,N_6077);
nor U7402 (N_7402,N_6571,N_6567);
and U7403 (N_7403,N_6463,N_6911);
nand U7404 (N_7404,N_6622,N_6945);
xor U7405 (N_7405,N_6758,N_6296);
and U7406 (N_7406,N_7101,N_6964);
xnor U7407 (N_7407,N_6173,N_6756);
nor U7408 (N_7408,N_6237,N_6450);
nand U7409 (N_7409,N_7028,N_6610);
and U7410 (N_7410,N_6087,N_6882);
xnor U7411 (N_7411,N_6141,N_6402);
nand U7412 (N_7412,N_6394,N_6538);
and U7413 (N_7413,N_6262,N_6788);
nand U7414 (N_7414,N_6073,N_6046);
nand U7415 (N_7415,N_7176,N_6221);
or U7416 (N_7416,N_7019,N_6001);
or U7417 (N_7417,N_7141,N_6914);
nor U7418 (N_7418,N_6745,N_6804);
xor U7419 (N_7419,N_6373,N_6464);
or U7420 (N_7420,N_6981,N_7193);
nand U7421 (N_7421,N_7097,N_6883);
nand U7422 (N_7422,N_6795,N_6955);
and U7423 (N_7423,N_6445,N_6827);
nor U7424 (N_7424,N_6423,N_6243);
or U7425 (N_7425,N_6591,N_7039);
and U7426 (N_7426,N_6757,N_6449);
nor U7427 (N_7427,N_6348,N_7050);
or U7428 (N_7428,N_6409,N_6239);
and U7429 (N_7429,N_6511,N_6997);
and U7430 (N_7430,N_6452,N_6959);
or U7431 (N_7431,N_7044,N_6987);
xor U7432 (N_7432,N_6009,N_6261);
xor U7433 (N_7433,N_6967,N_6894);
and U7434 (N_7434,N_6642,N_6792);
nand U7435 (N_7435,N_6264,N_7125);
xor U7436 (N_7436,N_6921,N_7168);
xor U7437 (N_7437,N_6211,N_6013);
or U7438 (N_7438,N_6235,N_7147);
and U7439 (N_7439,N_6489,N_6338);
nand U7440 (N_7440,N_6887,N_7121);
and U7441 (N_7441,N_6923,N_6743);
nand U7442 (N_7442,N_6487,N_6042);
nor U7443 (N_7443,N_6840,N_6390);
or U7444 (N_7444,N_6568,N_6078);
xnor U7445 (N_7445,N_6003,N_6246);
xor U7446 (N_7446,N_6209,N_7194);
or U7447 (N_7447,N_6447,N_7049);
nand U7448 (N_7448,N_6011,N_6462);
or U7449 (N_7449,N_6500,N_6293);
or U7450 (N_7450,N_6982,N_6667);
and U7451 (N_7451,N_6807,N_7163);
nor U7452 (N_7452,N_6658,N_6138);
nand U7453 (N_7453,N_6902,N_6428);
nor U7454 (N_7454,N_6388,N_6434);
or U7455 (N_7455,N_7184,N_7127);
and U7456 (N_7456,N_6152,N_6118);
and U7457 (N_7457,N_6991,N_6942);
and U7458 (N_7458,N_6639,N_6180);
nand U7459 (N_7459,N_6121,N_6014);
xor U7460 (N_7460,N_6456,N_6931);
nor U7461 (N_7461,N_6097,N_6181);
nor U7462 (N_7462,N_6028,N_6922);
nand U7463 (N_7463,N_6781,N_6441);
nor U7464 (N_7464,N_7081,N_6326);
xnor U7465 (N_7465,N_6637,N_7014);
nor U7466 (N_7466,N_6309,N_6651);
and U7467 (N_7467,N_6722,N_6810);
xnor U7468 (N_7468,N_6518,N_6083);
xnor U7469 (N_7469,N_6466,N_6783);
nand U7470 (N_7470,N_7186,N_6984);
or U7471 (N_7471,N_7196,N_6370);
nor U7472 (N_7472,N_7038,N_7177);
and U7473 (N_7473,N_6749,N_6918);
nor U7474 (N_7474,N_6171,N_6429);
and U7475 (N_7475,N_6329,N_6335);
or U7476 (N_7476,N_6878,N_6662);
and U7477 (N_7477,N_6944,N_6484);
or U7478 (N_7478,N_6153,N_6841);
nand U7479 (N_7479,N_7027,N_7061);
or U7480 (N_7480,N_7167,N_6641);
nor U7481 (N_7481,N_6995,N_7092);
xnor U7482 (N_7482,N_6381,N_6112);
nand U7483 (N_7483,N_6364,N_6618);
xor U7484 (N_7484,N_6490,N_6620);
and U7485 (N_7485,N_6728,N_6039);
nor U7486 (N_7486,N_6208,N_6313);
nand U7487 (N_7487,N_6494,N_7036);
nand U7488 (N_7488,N_7074,N_6860);
xnor U7489 (N_7489,N_7011,N_6796);
nand U7490 (N_7490,N_6357,N_7072);
nor U7491 (N_7491,N_6871,N_6815);
or U7492 (N_7492,N_6392,N_7020);
nor U7493 (N_7493,N_6844,N_7111);
nor U7494 (N_7494,N_6602,N_6539);
nor U7495 (N_7495,N_7043,N_6195);
and U7496 (N_7496,N_6867,N_6414);
and U7497 (N_7497,N_6700,N_6396);
or U7498 (N_7498,N_6159,N_6994);
and U7499 (N_7499,N_6371,N_6580);
nor U7500 (N_7500,N_7058,N_6852);
nor U7501 (N_7501,N_6512,N_7082);
xnor U7502 (N_7502,N_7032,N_6188);
or U7503 (N_7503,N_6938,N_6080);
or U7504 (N_7504,N_7067,N_6655);
nand U7505 (N_7505,N_7103,N_6535);
or U7506 (N_7506,N_6133,N_6585);
or U7507 (N_7507,N_6822,N_6273);
or U7508 (N_7508,N_6839,N_6385);
nor U7509 (N_7509,N_6249,N_6735);
nand U7510 (N_7510,N_6366,N_6957);
or U7511 (N_7511,N_6703,N_6851);
nor U7512 (N_7512,N_6563,N_6716);
nand U7513 (N_7513,N_6474,N_7005);
nand U7514 (N_7514,N_6684,N_6634);
and U7515 (N_7515,N_6105,N_6170);
nor U7516 (N_7516,N_6425,N_6565);
and U7517 (N_7517,N_7096,N_6709);
xnor U7518 (N_7518,N_6835,N_7132);
and U7519 (N_7519,N_6256,N_6936);
xor U7520 (N_7520,N_6176,N_6522);
or U7521 (N_7521,N_6098,N_6330);
or U7522 (N_7522,N_6816,N_6252);
xnor U7523 (N_7523,N_6205,N_6820);
and U7524 (N_7524,N_6214,N_6079);
xor U7525 (N_7525,N_7175,N_6775);
xor U7526 (N_7526,N_6164,N_7088);
or U7527 (N_7527,N_6199,N_7133);
nand U7528 (N_7528,N_6142,N_6985);
and U7529 (N_7529,N_6032,N_6765);
nand U7530 (N_7530,N_7106,N_6427);
xnor U7531 (N_7531,N_6823,N_6912);
and U7532 (N_7532,N_6081,N_6163);
nor U7533 (N_7533,N_6005,N_7000);
xor U7534 (N_7534,N_6020,N_6746);
nor U7535 (N_7535,N_7087,N_6247);
or U7536 (N_7536,N_6038,N_6012);
and U7537 (N_7537,N_6972,N_6383);
nor U7538 (N_7538,N_6659,N_6177);
or U7539 (N_7539,N_6996,N_6193);
or U7540 (N_7540,N_6389,N_6777);
nand U7541 (N_7541,N_6139,N_6233);
nand U7542 (N_7542,N_6675,N_7199);
or U7543 (N_7543,N_6114,N_6161);
nand U7544 (N_7544,N_6107,N_6318);
xnor U7545 (N_7545,N_7031,N_6426);
nor U7546 (N_7546,N_6377,N_6060);
xnor U7547 (N_7547,N_7138,N_6606);
nand U7548 (N_7548,N_6889,N_6197);
nand U7549 (N_7549,N_6838,N_6267);
or U7550 (N_7550,N_6479,N_7192);
nor U7551 (N_7551,N_6590,N_6467);
nor U7552 (N_7552,N_6059,N_6640);
and U7553 (N_7553,N_6310,N_6542);
xnor U7554 (N_7554,N_6282,N_7169);
or U7555 (N_7555,N_7190,N_7118);
xor U7556 (N_7556,N_6380,N_7080);
xnor U7557 (N_7557,N_6015,N_7045);
xnor U7558 (N_7558,N_6577,N_6085);
nand U7559 (N_7559,N_7180,N_6708);
nand U7560 (N_7560,N_6730,N_6277);
and U7561 (N_7561,N_6375,N_6734);
nand U7562 (N_7562,N_6582,N_6151);
nand U7563 (N_7563,N_6485,N_6925);
nand U7564 (N_7564,N_7073,N_6292);
nor U7565 (N_7565,N_7128,N_6050);
nand U7566 (N_7566,N_6460,N_6530);
nand U7567 (N_7567,N_6899,N_6317);
nor U7568 (N_7568,N_6692,N_6424);
nor U7569 (N_7569,N_6245,N_6108);
nand U7570 (N_7570,N_6191,N_6891);
and U7571 (N_7571,N_6978,N_6155);
nand U7572 (N_7572,N_6444,N_6415);
nand U7573 (N_7573,N_6316,N_6864);
and U7574 (N_7574,N_6748,N_6909);
xor U7575 (N_7575,N_6096,N_7152);
nor U7576 (N_7576,N_7173,N_6927);
nand U7577 (N_7577,N_6514,N_7185);
nor U7578 (N_7578,N_6900,N_7075);
or U7579 (N_7579,N_6884,N_7083);
or U7580 (N_7580,N_6420,N_6227);
and U7581 (N_7581,N_7136,N_7026);
nand U7582 (N_7582,N_7164,N_6033);
nand U7583 (N_7583,N_6017,N_6963);
or U7584 (N_7584,N_6573,N_6327);
and U7585 (N_7585,N_6830,N_6457);
and U7586 (N_7586,N_7002,N_6023);
or U7587 (N_7587,N_6106,N_6631);
nor U7588 (N_7588,N_6930,N_6828);
nand U7589 (N_7589,N_6853,N_6965);
nor U7590 (N_7590,N_6516,N_6158);
and U7591 (N_7591,N_6055,N_6234);
nand U7592 (N_7592,N_6971,N_6628);
nand U7593 (N_7593,N_6263,N_6302);
xor U7594 (N_7594,N_6711,N_7048);
nor U7595 (N_7595,N_6216,N_6819);
and U7596 (N_7596,N_6407,N_6952);
and U7597 (N_7597,N_6615,N_6113);
or U7598 (N_7598,N_6953,N_6717);
and U7599 (N_7599,N_6030,N_6653);
or U7600 (N_7600,N_6481,N_6368);
xor U7601 (N_7601,N_7008,N_6879);
nor U7602 (N_7602,N_6154,N_6943);
nor U7603 (N_7603,N_6259,N_6682);
and U7604 (N_7604,N_6731,N_6049);
and U7605 (N_7605,N_6376,N_7013);
nand U7606 (N_7606,N_6727,N_6021);
nand U7607 (N_7607,N_6774,N_6559);
and U7608 (N_7608,N_6000,N_6182);
and U7609 (N_7609,N_6435,N_7006);
xor U7610 (N_7610,N_6369,N_6007);
xor U7611 (N_7611,N_6710,N_6948);
or U7612 (N_7612,N_6940,N_7089);
nand U7613 (N_7613,N_6478,N_6147);
nand U7614 (N_7614,N_6818,N_6686);
xor U7615 (N_7615,N_6623,N_6045);
xnor U7616 (N_7616,N_7015,N_6412);
or U7617 (N_7617,N_6754,N_6315);
or U7618 (N_7618,N_6156,N_6545);
nand U7619 (N_7619,N_6454,N_6863);
xnor U7620 (N_7620,N_7053,N_6053);
nand U7621 (N_7621,N_6374,N_6403);
and U7622 (N_7622,N_6544,N_7166);
nand U7623 (N_7623,N_7165,N_6311);
nor U7624 (N_7624,N_6738,N_6220);
nand U7625 (N_7625,N_6600,N_7179);
nand U7626 (N_7626,N_7098,N_6979);
nor U7627 (N_7627,N_6956,N_7091);
or U7628 (N_7628,N_6271,N_7139);
nand U7629 (N_7629,N_6561,N_6524);
and U7630 (N_7630,N_6869,N_6365);
nor U7631 (N_7631,N_6290,N_6586);
or U7632 (N_7632,N_6694,N_6702);
nand U7633 (N_7633,N_6695,N_6503);
nor U7634 (N_7634,N_6384,N_6552);
nor U7635 (N_7635,N_6319,N_6413);
nor U7636 (N_7636,N_6359,N_6581);
nand U7637 (N_7637,N_6016,N_6636);
and U7638 (N_7638,N_6010,N_6018);
and U7639 (N_7639,N_6029,N_6802);
nor U7640 (N_7640,N_7109,N_6548);
and U7641 (N_7641,N_7056,N_6136);
nor U7642 (N_7642,N_6966,N_6408);
or U7643 (N_7643,N_6110,N_7068);
nor U7644 (N_7644,N_6872,N_6068);
and U7645 (N_7645,N_6506,N_6663);
xor U7646 (N_7646,N_6253,N_6410);
and U7647 (N_7647,N_6145,N_6865);
xor U7648 (N_7648,N_6787,N_6701);
or U7649 (N_7649,N_6784,N_6084);
nand U7650 (N_7650,N_6939,N_6941);
nand U7651 (N_7651,N_6705,N_7084);
xnor U7652 (N_7652,N_6320,N_6875);
xnor U7653 (N_7653,N_6473,N_6448);
nand U7654 (N_7654,N_6260,N_6550);
nor U7655 (N_7655,N_6649,N_6342);
nor U7656 (N_7656,N_6976,N_6975);
or U7657 (N_7657,N_6809,N_6935);
or U7658 (N_7658,N_6148,N_6973);
nor U7659 (N_7659,N_6472,N_6498);
or U7660 (N_7660,N_7189,N_6683);
and U7661 (N_7661,N_6172,N_7003);
nand U7662 (N_7662,N_7010,N_6575);
or U7663 (N_7663,N_6321,N_7155);
and U7664 (N_7664,N_6866,N_6837);
nand U7665 (N_7665,N_6763,N_6240);
xor U7666 (N_7666,N_6387,N_6276);
nor U7667 (N_7667,N_6958,N_6993);
nor U7668 (N_7668,N_6678,N_6690);
or U7669 (N_7669,N_6355,N_6328);
and U7670 (N_7670,N_7188,N_6437);
or U7671 (N_7671,N_6307,N_6644);
nor U7672 (N_7672,N_6786,N_6174);
nor U7673 (N_7673,N_6845,N_6753);
and U7674 (N_7674,N_6289,N_6629);
nand U7675 (N_7675,N_6742,N_6736);
or U7676 (N_7676,N_6160,N_7181);
nor U7677 (N_7677,N_7110,N_7130);
nand U7678 (N_7678,N_6089,N_6890);
xor U7679 (N_7679,N_6406,N_6555);
nor U7680 (N_7680,N_6601,N_6547);
nand U7681 (N_7681,N_6719,N_6190);
or U7682 (N_7682,N_6797,N_6356);
nor U7683 (N_7683,N_6857,N_6527);
and U7684 (N_7684,N_6115,N_6458);
and U7685 (N_7685,N_6562,N_6759);
nor U7686 (N_7686,N_6117,N_7131);
nor U7687 (N_7687,N_6917,N_6206);
or U7688 (N_7688,N_6501,N_6162);
or U7689 (N_7689,N_6551,N_7124);
and U7690 (N_7690,N_6399,N_6250);
xnor U7691 (N_7691,N_6025,N_6951);
or U7692 (N_7692,N_6961,N_6378);
and U7693 (N_7693,N_6168,N_7149);
nand U7694 (N_7694,N_6616,N_6597);
xor U7695 (N_7695,N_6339,N_6150);
xnor U7696 (N_7696,N_6713,N_6989);
or U7697 (N_7697,N_6468,N_6119);
or U7698 (N_7698,N_6897,N_7012);
nor U7699 (N_7699,N_6779,N_6612);
and U7700 (N_7700,N_6626,N_6859);
or U7701 (N_7701,N_6676,N_6803);
and U7702 (N_7702,N_7086,N_7197);
and U7703 (N_7703,N_6198,N_7108);
nand U7704 (N_7704,N_6854,N_6274);
nand U7705 (N_7705,N_6044,N_6969);
and U7706 (N_7706,N_6008,N_7042);
nand U7707 (N_7707,N_6397,N_6131);
or U7708 (N_7708,N_6222,N_6904);
nand U7709 (N_7709,N_6067,N_6483);
or U7710 (N_7710,N_7022,N_6026);
and U7711 (N_7711,N_6047,N_6596);
and U7712 (N_7712,N_6532,N_6137);
or U7713 (N_7713,N_6226,N_6687);
or U7714 (N_7714,N_6367,N_6549);
and U7715 (N_7715,N_6915,N_6422);
and U7716 (N_7716,N_6704,N_6099);
or U7717 (N_7717,N_6231,N_6266);
nand U7718 (N_7718,N_6574,N_6451);
nand U7719 (N_7719,N_6372,N_6143);
or U7720 (N_7720,N_7140,N_7001);
nor U7721 (N_7721,N_6095,N_6813);
nand U7722 (N_7722,N_6901,N_6954);
or U7723 (N_7723,N_7035,N_6229);
and U7724 (N_7724,N_6232,N_7142);
xnor U7725 (N_7725,N_6673,N_6750);
nor U7726 (N_7726,N_6486,N_6331);
or U7727 (N_7727,N_6949,N_6088);
and U7728 (N_7728,N_6656,N_7033);
or U7729 (N_7729,N_6043,N_7172);
nor U7730 (N_7730,N_6352,N_7024);
and U7731 (N_7731,N_6627,N_6120);
or U7732 (N_7732,N_6706,N_6048);
nand U7733 (N_7733,N_6771,N_6268);
and U7734 (N_7734,N_6306,N_6093);
and U7735 (N_7735,N_6660,N_7146);
nor U7736 (N_7736,N_7171,N_6517);
xor U7737 (N_7737,N_6604,N_6439);
and U7738 (N_7738,N_6861,N_6671);
xor U7739 (N_7739,N_6217,N_6346);
nor U7740 (N_7740,N_6291,N_6351);
and U7741 (N_7741,N_6314,N_6733);
xnor U7742 (N_7742,N_7094,N_6210);
nor U7743 (N_7743,N_6308,N_6341);
and U7744 (N_7744,N_6619,N_7034);
nand U7745 (N_7745,N_6265,N_6770);
or U7746 (N_7746,N_6762,N_6968);
or U7747 (N_7747,N_6537,N_6515);
nor U7748 (N_7748,N_6998,N_7195);
and U7749 (N_7749,N_6712,N_6519);
nand U7750 (N_7750,N_7004,N_6587);
and U7751 (N_7751,N_6322,N_6668);
xor U7752 (N_7752,N_6693,N_6661);
and U7753 (N_7753,N_6283,N_7100);
nor U7754 (N_7754,N_6301,N_7066);
xor U7755 (N_7755,N_6361,N_6906);
and U7756 (N_7756,N_7182,N_6714);
xnor U7757 (N_7757,N_6720,N_6334);
or U7758 (N_7758,N_6962,N_6654);
nor U7759 (N_7759,N_7143,N_6476);
nand U7760 (N_7760,N_6051,N_6913);
or U7761 (N_7761,N_6405,N_6843);
nor U7762 (N_7762,N_6528,N_6980);
nor U7763 (N_7763,N_7145,N_6772);
nor U7764 (N_7764,N_6461,N_7157);
nor U7765 (N_7765,N_6165,N_7099);
nor U7766 (N_7766,N_6304,N_6502);
or U7767 (N_7767,N_6536,N_6576);
and U7768 (N_7768,N_6400,N_6960);
nand U7769 (N_7769,N_6725,N_6140);
nor U7770 (N_7770,N_7105,N_7018);
xnor U7771 (N_7771,N_6124,N_6135);
xor U7772 (N_7772,N_6920,N_6149);
or U7773 (N_7773,N_6842,N_6521);
nor U7774 (N_7774,N_6723,N_6358);
nand U7775 (N_7775,N_7052,N_6789);
nor U7776 (N_7776,N_6907,N_6343);
nand U7777 (N_7777,N_6778,N_6255);
xnor U7778 (N_7778,N_6300,N_6805);
nand U7779 (N_7779,N_6721,N_7025);
xor U7780 (N_7780,N_6024,N_6111);
and U7781 (N_7781,N_6643,N_6785);
or U7782 (N_7782,N_6031,N_6393);
xnor U7783 (N_7783,N_7154,N_7178);
and U7784 (N_7784,N_6104,N_7113);
xnor U7785 (N_7785,N_6737,N_6363);
and U7786 (N_7786,N_6903,N_6986);
or U7787 (N_7787,N_7062,N_6895);
xor U7788 (N_7788,N_6201,N_6298);
xnor U7789 (N_7789,N_6999,N_6238);
or U7790 (N_7790,N_7017,N_6868);
xnor U7791 (N_7791,N_6888,N_6295);
nor U7792 (N_7792,N_7134,N_7065);
xnor U7793 (N_7793,N_6529,N_6480);
or U7794 (N_7794,N_6215,N_6332);
nand U7795 (N_7795,N_6493,N_7079);
nand U7796 (N_7796,N_7198,N_6617);
and U7797 (N_7797,N_6553,N_7187);
or U7798 (N_7798,N_7064,N_6065);
nor U7799 (N_7799,N_6071,N_6074);
nand U7800 (N_7800,N_6813,N_7015);
nor U7801 (N_7801,N_7084,N_7042);
or U7802 (N_7802,N_6325,N_6980);
nand U7803 (N_7803,N_6556,N_6087);
nor U7804 (N_7804,N_6598,N_6321);
nand U7805 (N_7805,N_6488,N_7099);
nand U7806 (N_7806,N_6142,N_6493);
and U7807 (N_7807,N_7167,N_6403);
or U7808 (N_7808,N_6011,N_6038);
and U7809 (N_7809,N_6184,N_6004);
and U7810 (N_7810,N_6138,N_6285);
and U7811 (N_7811,N_7169,N_6810);
xnor U7812 (N_7812,N_6851,N_6887);
nor U7813 (N_7813,N_6619,N_6813);
or U7814 (N_7814,N_6258,N_6171);
xnor U7815 (N_7815,N_6667,N_6254);
and U7816 (N_7816,N_6537,N_7137);
or U7817 (N_7817,N_7181,N_6491);
or U7818 (N_7818,N_6111,N_6575);
xor U7819 (N_7819,N_6351,N_6401);
nor U7820 (N_7820,N_6173,N_6206);
xor U7821 (N_7821,N_6199,N_6681);
or U7822 (N_7822,N_6419,N_6518);
nand U7823 (N_7823,N_6108,N_6201);
nand U7824 (N_7824,N_6865,N_6481);
xor U7825 (N_7825,N_7067,N_6637);
and U7826 (N_7826,N_6107,N_6598);
and U7827 (N_7827,N_6799,N_6032);
xor U7828 (N_7828,N_6153,N_6212);
nand U7829 (N_7829,N_7040,N_6751);
and U7830 (N_7830,N_6394,N_6944);
nand U7831 (N_7831,N_7169,N_7148);
or U7832 (N_7832,N_6035,N_6282);
nand U7833 (N_7833,N_6080,N_7186);
and U7834 (N_7834,N_6443,N_7060);
nor U7835 (N_7835,N_6967,N_6263);
nor U7836 (N_7836,N_6059,N_6429);
nor U7837 (N_7837,N_6247,N_6121);
nand U7838 (N_7838,N_6720,N_6140);
xor U7839 (N_7839,N_6735,N_6596);
xor U7840 (N_7840,N_6253,N_6874);
nor U7841 (N_7841,N_6487,N_6912);
nand U7842 (N_7842,N_6584,N_6317);
nand U7843 (N_7843,N_6073,N_7151);
and U7844 (N_7844,N_7051,N_6880);
or U7845 (N_7845,N_6191,N_6616);
and U7846 (N_7846,N_7191,N_6885);
xnor U7847 (N_7847,N_6755,N_6431);
nand U7848 (N_7848,N_6569,N_6688);
and U7849 (N_7849,N_6540,N_6829);
xor U7850 (N_7850,N_6038,N_6820);
xor U7851 (N_7851,N_7197,N_6071);
and U7852 (N_7852,N_6694,N_6988);
nor U7853 (N_7853,N_6401,N_6560);
or U7854 (N_7854,N_6287,N_6366);
nand U7855 (N_7855,N_6140,N_6419);
or U7856 (N_7856,N_7164,N_6700);
xnor U7857 (N_7857,N_6245,N_6774);
xor U7858 (N_7858,N_7054,N_6934);
and U7859 (N_7859,N_6381,N_6841);
xnor U7860 (N_7860,N_6019,N_6368);
and U7861 (N_7861,N_6626,N_6468);
nand U7862 (N_7862,N_6188,N_6838);
or U7863 (N_7863,N_6225,N_6465);
nor U7864 (N_7864,N_7005,N_6615);
xor U7865 (N_7865,N_6326,N_6737);
or U7866 (N_7866,N_6277,N_6589);
nand U7867 (N_7867,N_6035,N_6121);
nor U7868 (N_7868,N_6153,N_6109);
xnor U7869 (N_7869,N_7128,N_6098);
nor U7870 (N_7870,N_6295,N_6296);
or U7871 (N_7871,N_6990,N_6205);
xnor U7872 (N_7872,N_6905,N_7053);
or U7873 (N_7873,N_6258,N_6937);
and U7874 (N_7874,N_6548,N_6108);
and U7875 (N_7875,N_6561,N_6440);
and U7876 (N_7876,N_7149,N_6563);
nand U7877 (N_7877,N_6569,N_6377);
nor U7878 (N_7878,N_6884,N_6676);
and U7879 (N_7879,N_6483,N_7124);
or U7880 (N_7880,N_6766,N_6750);
nand U7881 (N_7881,N_6440,N_6271);
or U7882 (N_7882,N_6020,N_6433);
and U7883 (N_7883,N_6281,N_6916);
xnor U7884 (N_7884,N_7187,N_6472);
nand U7885 (N_7885,N_6249,N_6062);
nor U7886 (N_7886,N_6619,N_6785);
and U7887 (N_7887,N_6505,N_7116);
nand U7888 (N_7888,N_6991,N_7109);
or U7889 (N_7889,N_7030,N_7004);
and U7890 (N_7890,N_7162,N_6776);
xnor U7891 (N_7891,N_6398,N_6519);
or U7892 (N_7892,N_6380,N_6931);
nand U7893 (N_7893,N_6647,N_6282);
xnor U7894 (N_7894,N_7089,N_7030);
xor U7895 (N_7895,N_6679,N_6572);
xnor U7896 (N_7896,N_6980,N_6480);
or U7897 (N_7897,N_6954,N_6113);
or U7898 (N_7898,N_6037,N_7100);
or U7899 (N_7899,N_6138,N_6424);
and U7900 (N_7900,N_6712,N_7039);
nor U7901 (N_7901,N_7111,N_7172);
or U7902 (N_7902,N_7163,N_6083);
xnor U7903 (N_7903,N_6711,N_6628);
and U7904 (N_7904,N_6276,N_6031);
nand U7905 (N_7905,N_6986,N_7129);
nor U7906 (N_7906,N_6683,N_6883);
nand U7907 (N_7907,N_6852,N_6588);
xnor U7908 (N_7908,N_6468,N_6126);
xor U7909 (N_7909,N_6563,N_6046);
or U7910 (N_7910,N_6389,N_6099);
nor U7911 (N_7911,N_6042,N_6528);
nand U7912 (N_7912,N_6014,N_6556);
xor U7913 (N_7913,N_6357,N_7016);
nand U7914 (N_7914,N_6992,N_6022);
xor U7915 (N_7915,N_6790,N_7116);
nor U7916 (N_7916,N_6662,N_6122);
xor U7917 (N_7917,N_6295,N_6927);
and U7918 (N_7918,N_6820,N_6019);
or U7919 (N_7919,N_6931,N_6975);
xnor U7920 (N_7920,N_7194,N_6968);
and U7921 (N_7921,N_6086,N_6075);
nor U7922 (N_7922,N_7099,N_7042);
xnor U7923 (N_7923,N_6195,N_6147);
nand U7924 (N_7924,N_7189,N_6560);
xnor U7925 (N_7925,N_6967,N_6235);
xor U7926 (N_7926,N_6456,N_7070);
nor U7927 (N_7927,N_6321,N_6245);
and U7928 (N_7928,N_6910,N_7095);
xnor U7929 (N_7929,N_7019,N_6604);
and U7930 (N_7930,N_6102,N_6662);
nor U7931 (N_7931,N_6679,N_7018);
nor U7932 (N_7932,N_6026,N_6798);
xnor U7933 (N_7933,N_6532,N_6659);
nor U7934 (N_7934,N_7124,N_6848);
xor U7935 (N_7935,N_6412,N_6159);
nand U7936 (N_7936,N_6019,N_6668);
xnor U7937 (N_7937,N_6898,N_6714);
and U7938 (N_7938,N_7165,N_6284);
or U7939 (N_7939,N_6020,N_6941);
and U7940 (N_7940,N_6876,N_6055);
nor U7941 (N_7941,N_6803,N_7167);
and U7942 (N_7942,N_7081,N_7126);
xnor U7943 (N_7943,N_6344,N_6994);
nor U7944 (N_7944,N_6665,N_6664);
xnor U7945 (N_7945,N_7176,N_6169);
nand U7946 (N_7946,N_6058,N_6445);
nor U7947 (N_7947,N_7094,N_6421);
nor U7948 (N_7948,N_6448,N_6553);
or U7949 (N_7949,N_6088,N_6268);
nand U7950 (N_7950,N_6409,N_6612);
or U7951 (N_7951,N_6296,N_6751);
and U7952 (N_7952,N_6149,N_6370);
or U7953 (N_7953,N_7010,N_6015);
xnor U7954 (N_7954,N_6393,N_6366);
xor U7955 (N_7955,N_6061,N_6416);
xor U7956 (N_7956,N_6101,N_6318);
and U7957 (N_7957,N_6820,N_7056);
and U7958 (N_7958,N_6370,N_6361);
or U7959 (N_7959,N_6967,N_7096);
and U7960 (N_7960,N_6257,N_6429);
or U7961 (N_7961,N_6370,N_6328);
nor U7962 (N_7962,N_6165,N_7048);
nor U7963 (N_7963,N_6734,N_6854);
or U7964 (N_7964,N_6004,N_6928);
xor U7965 (N_7965,N_7066,N_7166);
nand U7966 (N_7966,N_7005,N_6074);
xor U7967 (N_7967,N_6729,N_6107);
nor U7968 (N_7968,N_6995,N_7188);
nand U7969 (N_7969,N_6474,N_6576);
nor U7970 (N_7970,N_7025,N_6433);
and U7971 (N_7971,N_7159,N_6206);
or U7972 (N_7972,N_6022,N_6042);
and U7973 (N_7973,N_6445,N_6663);
and U7974 (N_7974,N_6388,N_6111);
xnor U7975 (N_7975,N_6846,N_6002);
nor U7976 (N_7976,N_6392,N_6106);
or U7977 (N_7977,N_6947,N_6165);
nor U7978 (N_7978,N_6128,N_6037);
xor U7979 (N_7979,N_6430,N_6795);
nand U7980 (N_7980,N_6823,N_6189);
nor U7981 (N_7981,N_6404,N_6707);
or U7982 (N_7982,N_7065,N_7121);
or U7983 (N_7983,N_6420,N_6636);
nand U7984 (N_7984,N_6601,N_6771);
xor U7985 (N_7985,N_7065,N_6000);
and U7986 (N_7986,N_6742,N_6527);
xor U7987 (N_7987,N_7153,N_6089);
and U7988 (N_7988,N_7045,N_6785);
nor U7989 (N_7989,N_6423,N_7188);
nor U7990 (N_7990,N_6716,N_6447);
nor U7991 (N_7991,N_7138,N_6241);
or U7992 (N_7992,N_7120,N_6953);
and U7993 (N_7993,N_6868,N_6238);
xnor U7994 (N_7994,N_6269,N_6313);
nand U7995 (N_7995,N_6726,N_6908);
nand U7996 (N_7996,N_6899,N_6803);
and U7997 (N_7997,N_6221,N_6117);
nand U7998 (N_7998,N_6634,N_7103);
and U7999 (N_7999,N_6475,N_6832);
or U8000 (N_8000,N_6009,N_7026);
nand U8001 (N_8001,N_6620,N_6260);
nor U8002 (N_8002,N_7167,N_6656);
xnor U8003 (N_8003,N_6162,N_6006);
and U8004 (N_8004,N_6656,N_6059);
nor U8005 (N_8005,N_6419,N_6338);
nor U8006 (N_8006,N_6781,N_6776);
and U8007 (N_8007,N_6471,N_6864);
or U8008 (N_8008,N_6322,N_6140);
nor U8009 (N_8009,N_7088,N_6501);
or U8010 (N_8010,N_7195,N_6630);
nand U8011 (N_8011,N_6757,N_6599);
nor U8012 (N_8012,N_6837,N_6593);
and U8013 (N_8013,N_7100,N_6344);
nand U8014 (N_8014,N_7021,N_6911);
and U8015 (N_8015,N_6329,N_6292);
or U8016 (N_8016,N_6415,N_7039);
and U8017 (N_8017,N_6531,N_6451);
nor U8018 (N_8018,N_6661,N_6309);
and U8019 (N_8019,N_6489,N_6183);
nand U8020 (N_8020,N_6488,N_6593);
nand U8021 (N_8021,N_7077,N_6473);
nand U8022 (N_8022,N_6794,N_6070);
xor U8023 (N_8023,N_6303,N_6170);
or U8024 (N_8024,N_7003,N_6171);
and U8025 (N_8025,N_6493,N_6671);
and U8026 (N_8026,N_6658,N_6837);
or U8027 (N_8027,N_7105,N_6280);
nand U8028 (N_8028,N_6773,N_6960);
nor U8029 (N_8029,N_6096,N_6911);
and U8030 (N_8030,N_6225,N_6025);
or U8031 (N_8031,N_6782,N_6497);
xnor U8032 (N_8032,N_6852,N_7041);
nand U8033 (N_8033,N_6056,N_6495);
or U8034 (N_8034,N_6000,N_7175);
nor U8035 (N_8035,N_6967,N_6342);
nor U8036 (N_8036,N_6529,N_6192);
nor U8037 (N_8037,N_7128,N_6522);
nand U8038 (N_8038,N_6871,N_6641);
nand U8039 (N_8039,N_7179,N_6629);
nor U8040 (N_8040,N_6319,N_6666);
or U8041 (N_8041,N_7178,N_6753);
xor U8042 (N_8042,N_6700,N_6453);
and U8043 (N_8043,N_7024,N_6490);
and U8044 (N_8044,N_7187,N_6850);
xnor U8045 (N_8045,N_6033,N_6922);
or U8046 (N_8046,N_6415,N_6443);
nor U8047 (N_8047,N_6701,N_6691);
nor U8048 (N_8048,N_6049,N_6554);
nor U8049 (N_8049,N_6124,N_6544);
nor U8050 (N_8050,N_6062,N_6285);
or U8051 (N_8051,N_6162,N_6533);
xor U8052 (N_8052,N_6894,N_6995);
nand U8053 (N_8053,N_6446,N_6942);
nor U8054 (N_8054,N_6765,N_6886);
or U8055 (N_8055,N_6002,N_6624);
or U8056 (N_8056,N_6282,N_6277);
nand U8057 (N_8057,N_6353,N_6196);
nand U8058 (N_8058,N_6898,N_6775);
and U8059 (N_8059,N_6114,N_6062);
nand U8060 (N_8060,N_7037,N_6601);
nand U8061 (N_8061,N_6657,N_6462);
nand U8062 (N_8062,N_7010,N_6654);
xor U8063 (N_8063,N_6941,N_6138);
or U8064 (N_8064,N_6672,N_6574);
xor U8065 (N_8065,N_6601,N_7196);
and U8066 (N_8066,N_6972,N_6869);
xnor U8067 (N_8067,N_6574,N_6745);
or U8068 (N_8068,N_7133,N_6569);
nor U8069 (N_8069,N_6356,N_6352);
xnor U8070 (N_8070,N_6686,N_6002);
xor U8071 (N_8071,N_7022,N_7136);
nand U8072 (N_8072,N_6230,N_6629);
nand U8073 (N_8073,N_6642,N_6340);
xor U8074 (N_8074,N_6289,N_7098);
xnor U8075 (N_8075,N_6082,N_6888);
nor U8076 (N_8076,N_6386,N_6169);
xor U8077 (N_8077,N_6276,N_6209);
nor U8078 (N_8078,N_6050,N_6695);
or U8079 (N_8079,N_6706,N_6344);
nor U8080 (N_8080,N_6303,N_6342);
nand U8081 (N_8081,N_6707,N_6538);
or U8082 (N_8082,N_6913,N_6058);
or U8083 (N_8083,N_6066,N_6971);
or U8084 (N_8084,N_6576,N_6733);
nand U8085 (N_8085,N_6846,N_6380);
or U8086 (N_8086,N_7127,N_7080);
or U8087 (N_8087,N_6542,N_6128);
and U8088 (N_8088,N_6058,N_6567);
nand U8089 (N_8089,N_6445,N_6473);
nor U8090 (N_8090,N_6349,N_6577);
nand U8091 (N_8091,N_6239,N_6195);
xnor U8092 (N_8092,N_6979,N_6099);
nand U8093 (N_8093,N_6269,N_6059);
nand U8094 (N_8094,N_6119,N_6931);
or U8095 (N_8095,N_6672,N_6422);
and U8096 (N_8096,N_6031,N_6390);
nand U8097 (N_8097,N_6941,N_7083);
or U8098 (N_8098,N_6632,N_7190);
xor U8099 (N_8099,N_6054,N_7061);
nand U8100 (N_8100,N_7183,N_6553);
nor U8101 (N_8101,N_6962,N_6065);
xnor U8102 (N_8102,N_7163,N_7013);
or U8103 (N_8103,N_6404,N_7153);
or U8104 (N_8104,N_6057,N_6583);
or U8105 (N_8105,N_6221,N_6904);
nor U8106 (N_8106,N_6706,N_7101);
xnor U8107 (N_8107,N_6404,N_6910);
and U8108 (N_8108,N_6641,N_6332);
or U8109 (N_8109,N_6113,N_6497);
and U8110 (N_8110,N_6522,N_6807);
or U8111 (N_8111,N_6481,N_6223);
nor U8112 (N_8112,N_6990,N_6436);
nand U8113 (N_8113,N_6666,N_6550);
nand U8114 (N_8114,N_7045,N_6228);
nand U8115 (N_8115,N_6548,N_6277);
and U8116 (N_8116,N_6678,N_6833);
xnor U8117 (N_8117,N_6498,N_6776);
and U8118 (N_8118,N_6449,N_6023);
nand U8119 (N_8119,N_6939,N_6977);
xor U8120 (N_8120,N_7130,N_6857);
or U8121 (N_8121,N_6593,N_6259);
xor U8122 (N_8122,N_6830,N_6376);
or U8123 (N_8123,N_6200,N_6695);
and U8124 (N_8124,N_6858,N_6343);
nand U8125 (N_8125,N_6089,N_7017);
nor U8126 (N_8126,N_6142,N_7177);
nor U8127 (N_8127,N_6944,N_6868);
and U8128 (N_8128,N_7161,N_6493);
and U8129 (N_8129,N_7151,N_6553);
nand U8130 (N_8130,N_6512,N_6936);
and U8131 (N_8131,N_6028,N_6983);
and U8132 (N_8132,N_6724,N_6529);
xor U8133 (N_8133,N_6849,N_6571);
or U8134 (N_8134,N_6730,N_6137);
nor U8135 (N_8135,N_6319,N_6396);
and U8136 (N_8136,N_6647,N_7160);
nand U8137 (N_8137,N_6390,N_6014);
nand U8138 (N_8138,N_6395,N_6336);
xor U8139 (N_8139,N_6695,N_6884);
nor U8140 (N_8140,N_6323,N_6573);
nor U8141 (N_8141,N_6588,N_6666);
xor U8142 (N_8142,N_6724,N_6582);
nand U8143 (N_8143,N_6587,N_6090);
or U8144 (N_8144,N_6648,N_6388);
nand U8145 (N_8145,N_6906,N_6232);
or U8146 (N_8146,N_7095,N_6914);
nor U8147 (N_8147,N_6489,N_7087);
xor U8148 (N_8148,N_6226,N_6981);
nand U8149 (N_8149,N_6775,N_6965);
xor U8150 (N_8150,N_6032,N_6453);
xnor U8151 (N_8151,N_6075,N_6354);
nor U8152 (N_8152,N_7092,N_6332);
or U8153 (N_8153,N_6709,N_6668);
nand U8154 (N_8154,N_6672,N_6071);
and U8155 (N_8155,N_7099,N_6318);
xnor U8156 (N_8156,N_7005,N_6954);
xor U8157 (N_8157,N_6521,N_6403);
nor U8158 (N_8158,N_6340,N_6286);
xnor U8159 (N_8159,N_7192,N_6226);
nand U8160 (N_8160,N_6115,N_7139);
nor U8161 (N_8161,N_6190,N_7031);
xor U8162 (N_8162,N_6291,N_6100);
and U8163 (N_8163,N_6204,N_6375);
nand U8164 (N_8164,N_6209,N_6406);
or U8165 (N_8165,N_7158,N_6778);
nand U8166 (N_8166,N_6912,N_6336);
xnor U8167 (N_8167,N_6212,N_6014);
xnor U8168 (N_8168,N_6843,N_6781);
and U8169 (N_8169,N_6189,N_7031);
xor U8170 (N_8170,N_6327,N_6827);
xor U8171 (N_8171,N_7195,N_6650);
and U8172 (N_8172,N_6975,N_7170);
and U8173 (N_8173,N_6477,N_6741);
or U8174 (N_8174,N_6577,N_6149);
nand U8175 (N_8175,N_6370,N_6123);
xnor U8176 (N_8176,N_6495,N_6033);
nand U8177 (N_8177,N_6117,N_6237);
nand U8178 (N_8178,N_6138,N_6866);
xnor U8179 (N_8179,N_6384,N_6704);
nand U8180 (N_8180,N_6008,N_6403);
xnor U8181 (N_8181,N_6816,N_6305);
or U8182 (N_8182,N_7108,N_6713);
nand U8183 (N_8183,N_6890,N_6389);
xor U8184 (N_8184,N_6457,N_6224);
nand U8185 (N_8185,N_6916,N_6274);
xor U8186 (N_8186,N_6276,N_6890);
xnor U8187 (N_8187,N_6520,N_6175);
or U8188 (N_8188,N_6367,N_6855);
nand U8189 (N_8189,N_6441,N_6501);
and U8190 (N_8190,N_6071,N_7095);
nand U8191 (N_8191,N_6366,N_6517);
nand U8192 (N_8192,N_6805,N_7088);
nor U8193 (N_8193,N_6464,N_6612);
and U8194 (N_8194,N_6875,N_6010);
xnor U8195 (N_8195,N_6208,N_6561);
and U8196 (N_8196,N_6908,N_6227);
or U8197 (N_8197,N_6451,N_6523);
or U8198 (N_8198,N_6822,N_6871);
or U8199 (N_8199,N_6467,N_6824);
nor U8200 (N_8200,N_6309,N_6524);
nand U8201 (N_8201,N_6812,N_6966);
or U8202 (N_8202,N_7121,N_6893);
or U8203 (N_8203,N_6655,N_6949);
and U8204 (N_8204,N_6408,N_7064);
or U8205 (N_8205,N_6544,N_6952);
or U8206 (N_8206,N_6082,N_6378);
nor U8207 (N_8207,N_7056,N_7109);
or U8208 (N_8208,N_7134,N_6940);
and U8209 (N_8209,N_6493,N_6342);
or U8210 (N_8210,N_6262,N_6149);
nand U8211 (N_8211,N_6845,N_6794);
nand U8212 (N_8212,N_6339,N_6575);
nor U8213 (N_8213,N_6030,N_6977);
nor U8214 (N_8214,N_6489,N_7162);
nor U8215 (N_8215,N_6284,N_6721);
nand U8216 (N_8216,N_6128,N_6033);
xnor U8217 (N_8217,N_6405,N_6508);
nor U8218 (N_8218,N_6418,N_6901);
nor U8219 (N_8219,N_6360,N_6856);
and U8220 (N_8220,N_6729,N_6211);
xor U8221 (N_8221,N_6194,N_6320);
nand U8222 (N_8222,N_6957,N_7017);
or U8223 (N_8223,N_6099,N_7143);
nand U8224 (N_8224,N_7174,N_6306);
nand U8225 (N_8225,N_6214,N_6792);
xor U8226 (N_8226,N_6437,N_6431);
and U8227 (N_8227,N_7097,N_6682);
and U8228 (N_8228,N_6577,N_6816);
nand U8229 (N_8229,N_6986,N_6327);
nand U8230 (N_8230,N_6495,N_6312);
xnor U8231 (N_8231,N_6151,N_6685);
nor U8232 (N_8232,N_6361,N_6772);
xor U8233 (N_8233,N_6447,N_6339);
nand U8234 (N_8234,N_6649,N_6938);
xor U8235 (N_8235,N_6668,N_6324);
or U8236 (N_8236,N_6011,N_6341);
nand U8237 (N_8237,N_6767,N_6214);
and U8238 (N_8238,N_6092,N_6100);
or U8239 (N_8239,N_6139,N_6501);
nand U8240 (N_8240,N_6443,N_6683);
xnor U8241 (N_8241,N_6660,N_6347);
xnor U8242 (N_8242,N_6206,N_6830);
xnor U8243 (N_8243,N_6861,N_6002);
nor U8244 (N_8244,N_6789,N_6849);
nor U8245 (N_8245,N_6283,N_6386);
xor U8246 (N_8246,N_6787,N_6981);
xor U8247 (N_8247,N_6916,N_6646);
and U8248 (N_8248,N_6771,N_6179);
or U8249 (N_8249,N_6979,N_7002);
and U8250 (N_8250,N_6878,N_6461);
or U8251 (N_8251,N_6616,N_6828);
xnor U8252 (N_8252,N_6982,N_7152);
nor U8253 (N_8253,N_6871,N_6165);
and U8254 (N_8254,N_7107,N_6841);
nor U8255 (N_8255,N_6497,N_6416);
nand U8256 (N_8256,N_6998,N_7176);
and U8257 (N_8257,N_6056,N_7131);
xnor U8258 (N_8258,N_6649,N_6311);
xnor U8259 (N_8259,N_6056,N_6261);
and U8260 (N_8260,N_6776,N_6701);
nor U8261 (N_8261,N_6190,N_6908);
or U8262 (N_8262,N_6108,N_6957);
and U8263 (N_8263,N_6933,N_7181);
xor U8264 (N_8264,N_6262,N_6298);
nand U8265 (N_8265,N_6846,N_6143);
nor U8266 (N_8266,N_6299,N_6511);
or U8267 (N_8267,N_6307,N_6887);
xor U8268 (N_8268,N_6502,N_6311);
nand U8269 (N_8269,N_7027,N_7012);
or U8270 (N_8270,N_6802,N_6143);
or U8271 (N_8271,N_6069,N_7107);
and U8272 (N_8272,N_6885,N_6730);
nor U8273 (N_8273,N_6808,N_6413);
or U8274 (N_8274,N_7082,N_6747);
and U8275 (N_8275,N_6868,N_7195);
and U8276 (N_8276,N_6283,N_6362);
or U8277 (N_8277,N_6329,N_6459);
nor U8278 (N_8278,N_6905,N_6489);
nand U8279 (N_8279,N_7110,N_7029);
nor U8280 (N_8280,N_6588,N_6524);
or U8281 (N_8281,N_6084,N_6179);
nor U8282 (N_8282,N_6810,N_6087);
or U8283 (N_8283,N_6700,N_6568);
or U8284 (N_8284,N_6385,N_6644);
or U8285 (N_8285,N_7190,N_7096);
nor U8286 (N_8286,N_6762,N_6210);
xnor U8287 (N_8287,N_6294,N_6213);
or U8288 (N_8288,N_6893,N_6560);
nand U8289 (N_8289,N_6810,N_6298);
or U8290 (N_8290,N_6629,N_6381);
nor U8291 (N_8291,N_6551,N_7150);
nand U8292 (N_8292,N_6595,N_6254);
nor U8293 (N_8293,N_6701,N_6940);
nor U8294 (N_8294,N_6204,N_6958);
xnor U8295 (N_8295,N_6627,N_6188);
and U8296 (N_8296,N_7117,N_7091);
nor U8297 (N_8297,N_7185,N_6928);
nor U8298 (N_8298,N_6912,N_6767);
nor U8299 (N_8299,N_6568,N_6445);
nand U8300 (N_8300,N_6529,N_6371);
or U8301 (N_8301,N_6427,N_6243);
xor U8302 (N_8302,N_6155,N_6723);
and U8303 (N_8303,N_7111,N_6692);
nor U8304 (N_8304,N_7190,N_7187);
or U8305 (N_8305,N_6844,N_7156);
nand U8306 (N_8306,N_6500,N_7077);
and U8307 (N_8307,N_7084,N_6792);
nor U8308 (N_8308,N_6245,N_7176);
and U8309 (N_8309,N_6406,N_6232);
and U8310 (N_8310,N_6984,N_6488);
nor U8311 (N_8311,N_6109,N_6965);
or U8312 (N_8312,N_6512,N_7193);
nor U8313 (N_8313,N_6018,N_6629);
nor U8314 (N_8314,N_6569,N_6417);
or U8315 (N_8315,N_6172,N_6044);
or U8316 (N_8316,N_6731,N_6450);
nand U8317 (N_8317,N_7078,N_7149);
or U8318 (N_8318,N_6324,N_6390);
nand U8319 (N_8319,N_6151,N_6916);
nand U8320 (N_8320,N_6514,N_6039);
xnor U8321 (N_8321,N_6552,N_6430);
and U8322 (N_8322,N_6145,N_7010);
nor U8323 (N_8323,N_6076,N_6999);
and U8324 (N_8324,N_6908,N_6202);
nor U8325 (N_8325,N_6989,N_7178);
or U8326 (N_8326,N_6647,N_6066);
nand U8327 (N_8327,N_6835,N_7103);
xor U8328 (N_8328,N_6732,N_6850);
nand U8329 (N_8329,N_7011,N_6572);
xnor U8330 (N_8330,N_6688,N_6086);
or U8331 (N_8331,N_7176,N_6717);
nand U8332 (N_8332,N_7062,N_7079);
nor U8333 (N_8333,N_7077,N_6560);
nand U8334 (N_8334,N_6740,N_7109);
nor U8335 (N_8335,N_7174,N_6764);
xnor U8336 (N_8336,N_6094,N_6931);
xor U8337 (N_8337,N_6001,N_7021);
or U8338 (N_8338,N_7124,N_6685);
nor U8339 (N_8339,N_6360,N_6565);
nand U8340 (N_8340,N_6766,N_6630);
xor U8341 (N_8341,N_6544,N_6475);
nor U8342 (N_8342,N_6747,N_6169);
and U8343 (N_8343,N_6883,N_6501);
xnor U8344 (N_8344,N_6385,N_6892);
and U8345 (N_8345,N_6150,N_6856);
nand U8346 (N_8346,N_6951,N_6315);
nor U8347 (N_8347,N_6994,N_6230);
and U8348 (N_8348,N_6247,N_6371);
and U8349 (N_8349,N_6954,N_6570);
and U8350 (N_8350,N_6971,N_6613);
or U8351 (N_8351,N_6243,N_7173);
nand U8352 (N_8352,N_6064,N_6048);
nor U8353 (N_8353,N_7011,N_6410);
xnor U8354 (N_8354,N_6899,N_6432);
or U8355 (N_8355,N_7101,N_6266);
nand U8356 (N_8356,N_6779,N_6795);
nor U8357 (N_8357,N_6781,N_6436);
xor U8358 (N_8358,N_6848,N_6862);
nand U8359 (N_8359,N_7103,N_6333);
and U8360 (N_8360,N_6201,N_6783);
xor U8361 (N_8361,N_6849,N_6804);
and U8362 (N_8362,N_7141,N_6507);
and U8363 (N_8363,N_6587,N_6688);
nor U8364 (N_8364,N_6632,N_6780);
and U8365 (N_8365,N_6607,N_7115);
and U8366 (N_8366,N_6027,N_6210);
and U8367 (N_8367,N_6615,N_6301);
or U8368 (N_8368,N_6689,N_6163);
nand U8369 (N_8369,N_6556,N_7017);
nor U8370 (N_8370,N_7009,N_7023);
or U8371 (N_8371,N_6913,N_6598);
xnor U8372 (N_8372,N_6602,N_7181);
xor U8373 (N_8373,N_6319,N_6887);
nor U8374 (N_8374,N_6502,N_6368);
or U8375 (N_8375,N_6531,N_6935);
nor U8376 (N_8376,N_6765,N_6366);
nor U8377 (N_8377,N_6181,N_6496);
or U8378 (N_8378,N_6151,N_6759);
or U8379 (N_8379,N_7047,N_6992);
and U8380 (N_8380,N_6422,N_6541);
or U8381 (N_8381,N_6378,N_6374);
xor U8382 (N_8382,N_7194,N_6464);
nor U8383 (N_8383,N_6229,N_6183);
nand U8384 (N_8384,N_6796,N_7027);
xor U8385 (N_8385,N_6433,N_6265);
and U8386 (N_8386,N_6372,N_6310);
and U8387 (N_8387,N_7023,N_6674);
and U8388 (N_8388,N_6769,N_7048);
nand U8389 (N_8389,N_6068,N_6679);
nand U8390 (N_8390,N_6138,N_6892);
and U8391 (N_8391,N_6931,N_6973);
xor U8392 (N_8392,N_7174,N_6431);
nor U8393 (N_8393,N_6665,N_6560);
nor U8394 (N_8394,N_6273,N_6524);
or U8395 (N_8395,N_6898,N_6450);
xor U8396 (N_8396,N_6379,N_6261);
xor U8397 (N_8397,N_6563,N_6264);
or U8398 (N_8398,N_6692,N_6410);
xor U8399 (N_8399,N_6472,N_6994);
or U8400 (N_8400,N_7787,N_7324);
or U8401 (N_8401,N_8064,N_8182);
and U8402 (N_8402,N_7322,N_8271);
and U8403 (N_8403,N_7482,N_7284);
nand U8404 (N_8404,N_7224,N_7936);
nor U8405 (N_8405,N_7659,N_8159);
nor U8406 (N_8406,N_7293,N_7361);
nor U8407 (N_8407,N_8050,N_7943);
nand U8408 (N_8408,N_7443,N_7635);
and U8409 (N_8409,N_7543,N_8371);
nor U8410 (N_8410,N_8038,N_7255);
nor U8411 (N_8411,N_7447,N_8367);
and U8412 (N_8412,N_7887,N_7473);
nor U8413 (N_8413,N_8336,N_8289);
nand U8414 (N_8414,N_8276,N_7474);
nor U8415 (N_8415,N_7963,N_8137);
nor U8416 (N_8416,N_7667,N_8356);
nor U8417 (N_8417,N_7258,N_7213);
or U8418 (N_8418,N_7750,N_7511);
nor U8419 (N_8419,N_7714,N_7535);
or U8420 (N_8420,N_7481,N_7939);
nor U8421 (N_8421,N_7432,N_8079);
or U8422 (N_8422,N_7625,N_8022);
or U8423 (N_8423,N_8178,N_7947);
and U8424 (N_8424,N_7825,N_7358);
or U8425 (N_8425,N_8049,N_7433);
xnor U8426 (N_8426,N_7412,N_8196);
nand U8427 (N_8427,N_7316,N_7982);
nand U8428 (N_8428,N_7927,N_7631);
xnor U8429 (N_8429,N_7405,N_7652);
or U8430 (N_8430,N_7634,N_8121);
and U8431 (N_8431,N_8136,N_7462);
xnor U8432 (N_8432,N_8353,N_7526);
or U8433 (N_8433,N_8036,N_7640);
xnor U8434 (N_8434,N_7704,N_8110);
nor U8435 (N_8435,N_7363,N_7458);
nor U8436 (N_8436,N_8335,N_8010);
and U8437 (N_8437,N_8295,N_8305);
xnor U8438 (N_8438,N_7669,N_7299);
nand U8439 (N_8439,N_7513,N_8005);
nor U8440 (N_8440,N_7344,N_8056);
or U8441 (N_8441,N_7238,N_7389);
and U8442 (N_8442,N_7239,N_7476);
and U8443 (N_8443,N_7710,N_8292);
or U8444 (N_8444,N_7990,N_7264);
and U8445 (N_8445,N_7368,N_7660);
nand U8446 (N_8446,N_8015,N_8372);
or U8447 (N_8447,N_7402,N_8157);
or U8448 (N_8448,N_8072,N_8177);
nor U8449 (N_8449,N_7451,N_7249);
xnor U8450 (N_8450,N_7833,N_8124);
nand U8451 (N_8451,N_8269,N_7510);
and U8452 (N_8452,N_8105,N_7338);
nand U8453 (N_8453,N_7556,N_8155);
xor U8454 (N_8454,N_8207,N_7973);
or U8455 (N_8455,N_8297,N_7257);
and U8456 (N_8456,N_8150,N_8008);
nor U8457 (N_8457,N_7904,N_7277);
nand U8458 (N_8458,N_7411,N_7618);
or U8459 (N_8459,N_8317,N_7487);
and U8460 (N_8460,N_7636,N_8054);
nor U8461 (N_8461,N_8166,N_7464);
nand U8462 (N_8462,N_7450,N_8384);
nor U8463 (N_8463,N_7656,N_7676);
nand U8464 (N_8464,N_8216,N_8218);
xor U8465 (N_8465,N_7657,N_7722);
xor U8466 (N_8466,N_8272,N_8252);
xor U8467 (N_8467,N_7522,N_7601);
nand U8468 (N_8468,N_8204,N_7680);
or U8469 (N_8469,N_7865,N_7502);
xor U8470 (N_8470,N_7350,N_7845);
nor U8471 (N_8471,N_7880,N_8299);
xnor U8472 (N_8472,N_7627,N_7665);
nand U8473 (N_8473,N_7839,N_7240);
and U8474 (N_8474,N_7414,N_7843);
and U8475 (N_8475,N_7568,N_7883);
nor U8476 (N_8476,N_8152,N_8045);
or U8477 (N_8477,N_8131,N_8115);
or U8478 (N_8478,N_7335,N_7427);
nor U8479 (N_8479,N_8030,N_7766);
or U8480 (N_8480,N_8173,N_8091);
and U8481 (N_8481,N_7615,N_7422);
nor U8482 (N_8482,N_7301,N_7546);
nand U8483 (N_8483,N_7811,N_7353);
nand U8484 (N_8484,N_7735,N_8326);
xnor U8485 (N_8485,N_8301,N_8311);
xor U8486 (N_8486,N_7649,N_7308);
nor U8487 (N_8487,N_8320,N_7800);
xor U8488 (N_8488,N_8026,N_8234);
or U8489 (N_8489,N_8338,N_7252);
xnor U8490 (N_8490,N_8314,N_7355);
and U8491 (N_8491,N_7746,N_7823);
and U8492 (N_8492,N_8241,N_7259);
xor U8493 (N_8493,N_7285,N_7337);
nand U8494 (N_8494,N_7767,N_7761);
nor U8495 (N_8495,N_8001,N_8349);
nor U8496 (N_8496,N_7648,N_7690);
nor U8497 (N_8497,N_7364,N_8130);
nor U8498 (N_8498,N_8307,N_7948);
xor U8499 (N_8499,N_7323,N_7393);
or U8500 (N_8500,N_7399,N_7668);
nand U8501 (N_8501,N_8151,N_8061);
and U8502 (N_8502,N_7595,N_8163);
xor U8503 (N_8503,N_8048,N_8189);
nor U8504 (N_8504,N_7609,N_7287);
xor U8505 (N_8505,N_8359,N_7849);
xnor U8506 (N_8506,N_8120,N_8215);
or U8507 (N_8507,N_7785,N_7897);
nand U8508 (N_8508,N_7744,N_7949);
xor U8509 (N_8509,N_7608,N_7431);
xor U8510 (N_8510,N_7586,N_7228);
nand U8511 (N_8511,N_7791,N_8341);
nor U8512 (N_8512,N_7540,N_7616);
nand U8513 (N_8513,N_7696,N_7330);
nand U8514 (N_8514,N_8098,N_7560);
or U8515 (N_8515,N_7260,N_8270);
and U8516 (N_8516,N_7452,N_7282);
and U8517 (N_8517,N_7349,N_8238);
xnor U8518 (N_8518,N_7694,N_7840);
or U8519 (N_8519,N_7396,N_7491);
nand U8520 (N_8520,N_7663,N_8065);
or U8521 (N_8521,N_7866,N_7573);
and U8522 (N_8522,N_7463,N_7569);
and U8523 (N_8523,N_8147,N_7279);
nand U8524 (N_8524,N_8334,N_8298);
nor U8525 (N_8525,N_7445,N_8290);
nor U8526 (N_8526,N_7242,N_7436);
xor U8527 (N_8527,N_7318,N_8073);
and U8528 (N_8528,N_8123,N_7995);
nor U8529 (N_8529,N_7553,N_7521);
nor U8530 (N_8530,N_7374,N_7759);
and U8531 (N_8531,N_7738,N_7524);
or U8532 (N_8532,N_8258,N_7468);
or U8533 (N_8533,N_8191,N_7327);
xnor U8534 (N_8534,N_8244,N_7698);
xnor U8535 (N_8535,N_8057,N_7333);
and U8536 (N_8536,N_7666,N_8192);
nor U8537 (N_8537,N_8236,N_7429);
nand U8538 (N_8538,N_8176,N_8232);
nand U8539 (N_8539,N_8351,N_7243);
nand U8540 (N_8540,N_7902,N_7769);
nand U8541 (N_8541,N_7864,N_7461);
nand U8542 (N_8542,N_7629,N_8145);
xor U8543 (N_8543,N_7517,N_7960);
nor U8544 (N_8544,N_7894,N_8169);
nor U8545 (N_8545,N_7886,N_8162);
nor U8546 (N_8546,N_7821,N_7419);
nor U8547 (N_8547,N_8394,N_8200);
xnor U8548 (N_8548,N_7380,N_7289);
or U8549 (N_8549,N_7362,N_8055);
nor U8550 (N_8550,N_7683,N_8245);
or U8551 (N_8551,N_7490,N_8278);
nor U8552 (N_8552,N_8085,N_7590);
nor U8553 (N_8553,N_8206,N_7533);
or U8554 (N_8554,N_8309,N_7415);
xor U8555 (N_8555,N_7876,N_7398);
and U8556 (N_8556,N_8190,N_7860);
xnor U8557 (N_8557,N_8275,N_7519);
or U8558 (N_8558,N_7575,N_7921);
and U8559 (N_8559,N_7945,N_7729);
nand U8560 (N_8560,N_8249,N_7600);
xnor U8561 (N_8561,N_7512,N_8285);
and U8562 (N_8562,N_7583,N_7717);
or U8563 (N_8563,N_8165,N_7888);
nor U8564 (N_8564,N_8369,N_8293);
and U8565 (N_8565,N_7976,N_7664);
nand U8566 (N_8566,N_7241,N_7449);
xor U8567 (N_8567,N_7745,N_7388);
xor U8568 (N_8568,N_7773,N_7699);
nor U8569 (N_8569,N_7373,N_7879);
or U8570 (N_8570,N_7713,N_7923);
nor U8571 (N_8571,N_7387,N_7971);
nand U8572 (N_8572,N_8254,N_7986);
xnor U8573 (N_8573,N_7806,N_7961);
xor U8574 (N_8574,N_7263,N_7911);
nand U8575 (N_8575,N_8257,N_7455);
nor U8576 (N_8576,N_7736,N_7807);
nand U8577 (N_8577,N_8199,N_7312);
nand U8578 (N_8578,N_7313,N_7742);
nor U8579 (N_8579,N_7547,N_8004);
xor U8580 (N_8580,N_7944,N_8081);
xor U8581 (N_8581,N_8323,N_8350);
and U8582 (N_8582,N_7917,N_7370);
and U8583 (N_8583,N_7441,N_7261);
nand U8584 (N_8584,N_7235,N_7734);
xor U8585 (N_8585,N_7805,N_7444);
and U8586 (N_8586,N_8087,N_8160);
and U8587 (N_8587,N_8108,N_7677);
or U8588 (N_8588,N_7267,N_7671);
nand U8589 (N_8589,N_7584,N_7222);
nor U8590 (N_8590,N_7296,N_7993);
xor U8591 (N_8591,N_8116,N_7715);
nor U8592 (N_8592,N_8067,N_7525);
nor U8593 (N_8593,N_7347,N_7813);
nand U8594 (N_8594,N_7689,N_7397);
nor U8595 (N_8595,N_7915,N_7326);
and U8596 (N_8596,N_7203,N_8223);
and U8597 (N_8597,N_7695,N_7996);
nor U8598 (N_8598,N_7246,N_7731);
and U8599 (N_8599,N_7930,N_8247);
xor U8600 (N_8600,N_7256,N_8329);
xor U8601 (N_8601,N_8063,N_7617);
xnor U8602 (N_8602,N_7214,N_7782);
nor U8603 (N_8603,N_8346,N_7765);
and U8604 (N_8604,N_8273,N_7647);
nor U8605 (N_8605,N_8397,N_8266);
nor U8606 (N_8606,N_7375,N_8167);
or U8607 (N_8607,N_7581,N_7220);
nor U8608 (N_8608,N_8071,N_7542);
or U8609 (N_8609,N_7612,N_7779);
or U8610 (N_8610,N_7899,N_7898);
and U8611 (N_8611,N_8377,N_7868);
or U8612 (N_8612,N_7937,N_7611);
or U8613 (N_8613,N_7691,N_7558);
and U8614 (N_8614,N_8093,N_7645);
nor U8615 (N_8615,N_8274,N_8313);
and U8616 (N_8616,N_7869,N_7622);
xor U8617 (N_8617,N_7651,N_7372);
and U8618 (N_8618,N_7837,N_7851);
nor U8619 (N_8619,N_7409,N_7836);
nor U8620 (N_8620,N_7774,N_8194);
nand U8621 (N_8621,N_8017,N_7549);
nand U8622 (N_8622,N_7489,N_7877);
and U8623 (N_8623,N_8186,N_7295);
or U8624 (N_8624,N_8066,N_7340);
or U8625 (N_8625,N_7391,N_8214);
or U8626 (N_8626,N_7200,N_8312);
or U8627 (N_8627,N_8128,N_7972);
xnor U8628 (N_8628,N_7795,N_7788);
or U8629 (N_8629,N_7217,N_7269);
nor U8630 (N_8630,N_8102,N_7733);
xor U8631 (N_8631,N_7410,N_7594);
xnor U8632 (N_8632,N_8043,N_7365);
and U8633 (N_8633,N_8154,N_7223);
or U8634 (N_8634,N_7237,N_8170);
nor U8635 (N_8635,N_8125,N_7968);
nand U8636 (N_8636,N_7933,N_7799);
nand U8637 (N_8637,N_7446,N_7751);
nand U8638 (N_8638,N_7529,N_7278);
or U8639 (N_8639,N_7830,N_7946);
nand U8640 (N_8640,N_8158,N_8304);
or U8641 (N_8641,N_8358,N_7254);
and U8642 (N_8642,N_7701,N_7245);
and U8643 (N_8643,N_7828,N_7764);
and U8644 (N_8644,N_7250,N_7369);
xnor U8645 (N_8645,N_8342,N_7570);
nand U8646 (N_8646,N_8264,N_7614);
and U8647 (N_8647,N_7824,N_7918);
nor U8648 (N_8648,N_7564,N_7354);
nor U8649 (N_8649,N_8226,N_8140);
nor U8650 (N_8650,N_8227,N_7628);
and U8651 (N_8651,N_7814,N_8046);
nor U8652 (N_8652,N_7928,N_7724);
nor U8653 (N_8653,N_7232,N_7501);
or U8654 (N_8654,N_7497,N_8197);
nand U8655 (N_8655,N_7720,N_7992);
xor U8656 (N_8656,N_7784,N_7802);
or U8657 (N_8657,N_7619,N_7924);
or U8658 (N_8658,N_7456,N_8282);
nand U8659 (N_8659,N_7857,N_7459);
and U8660 (N_8660,N_7827,N_7610);
nand U8661 (N_8661,N_8332,N_7233);
or U8662 (N_8662,N_7658,N_8279);
nor U8663 (N_8663,N_7748,N_7925);
nor U8664 (N_8664,N_7226,N_8246);
and U8665 (N_8665,N_8259,N_7320);
nand U8666 (N_8666,N_8094,N_8024);
nor U8667 (N_8667,N_7931,N_8181);
nand U8668 (N_8668,N_8229,N_7832);
nor U8669 (N_8669,N_8316,N_7752);
or U8670 (N_8670,N_7571,N_8149);
nand U8671 (N_8671,N_7721,N_8080);
nand U8672 (N_8672,N_7229,N_8347);
nand U8673 (N_8673,N_7777,N_7483);
nand U8674 (N_8674,N_7674,N_8062);
xor U8675 (N_8675,N_7906,N_7563);
and U8676 (N_8676,N_7567,N_8286);
or U8677 (N_8677,N_8075,N_7878);
xor U8678 (N_8678,N_7820,N_7826);
nand U8679 (N_8679,N_7938,N_7620);
xor U8680 (N_8680,N_7390,N_7498);
xnor U8681 (N_8681,N_7797,N_7465);
and U8682 (N_8682,N_7211,N_7808);
and U8683 (N_8683,N_7964,N_8357);
nand U8684 (N_8684,N_7273,N_7988);
or U8685 (N_8685,N_7528,N_7291);
or U8686 (N_8686,N_7381,N_8002);
nand U8687 (N_8687,N_7210,N_7884);
nor U8688 (N_8688,N_7951,N_7231);
xnor U8689 (N_8689,N_7896,N_8277);
nand U8690 (N_8690,N_7606,N_8374);
nor U8691 (N_8691,N_7321,N_7794);
and U8692 (N_8692,N_8378,N_7598);
or U8693 (N_8693,N_7440,N_8052);
and U8694 (N_8694,N_8156,N_7859);
and U8695 (N_8695,N_7585,N_7225);
xor U8696 (N_8696,N_8360,N_8039);
nand U8697 (N_8697,N_8396,N_8082);
nand U8698 (N_8698,N_7589,N_7379);
nor U8699 (N_8699,N_7418,N_7294);
nor U8700 (N_8700,N_8308,N_7934);
or U8701 (N_8701,N_7406,N_7726);
nand U8702 (N_8702,N_7219,N_7413);
xnor U8703 (N_8703,N_7711,N_7999);
xnor U8704 (N_8704,N_7780,N_7655);
or U8705 (N_8705,N_7514,N_8033);
xor U8706 (N_8706,N_7812,N_7435);
nor U8707 (N_8707,N_8393,N_8168);
xnor U8708 (N_8708,N_7965,N_7247);
xnor U8709 (N_8709,N_8348,N_7979);
nand U8710 (N_8710,N_7974,N_7508);
nor U8711 (N_8711,N_8090,N_8035);
xor U8712 (N_8712,N_7653,N_7216);
nand U8713 (N_8713,N_7856,N_8013);
nor U8714 (N_8714,N_7457,N_7378);
and U8715 (N_8715,N_7700,N_7343);
or U8716 (N_8716,N_7822,N_7817);
or U8717 (N_8717,N_7342,N_7500);
and U8718 (N_8718,N_7920,N_7728);
or U8719 (N_8719,N_8146,N_8250);
xor U8720 (N_8720,N_8325,N_8243);
or U8721 (N_8721,N_7309,N_7959);
nand U8722 (N_8722,N_8032,N_7719);
and U8723 (N_8723,N_8209,N_8122);
or U8724 (N_8724,N_7339,N_7985);
nor U8725 (N_8725,N_8319,N_7532);
nand U8726 (N_8726,N_7912,N_8034);
xor U8727 (N_8727,N_7204,N_8138);
nor U8728 (N_8728,N_8028,N_7329);
xnor U8729 (N_8729,N_7297,N_7493);
nor U8730 (N_8730,N_8132,N_8127);
nor U8731 (N_8731,N_8047,N_7919);
nor U8732 (N_8732,N_7492,N_8092);
or U8733 (N_8733,N_8179,N_7607);
and U8734 (N_8734,N_7408,N_7477);
nor U8735 (N_8735,N_8095,N_7940);
and U8736 (N_8736,N_7967,N_7360);
or U8737 (N_8737,N_8037,N_7395);
and U8738 (N_8738,N_8007,N_7809);
or U8739 (N_8739,N_7882,N_8175);
nor U8740 (N_8740,N_7420,N_7206);
nor U8741 (N_8741,N_8041,N_7212);
nand U8742 (N_8742,N_8231,N_8113);
or U8743 (N_8743,N_7305,N_8253);
nand U8744 (N_8744,N_7929,N_7834);
nand U8745 (N_8745,N_8172,N_8174);
nand U8746 (N_8746,N_7209,N_8315);
xnor U8747 (N_8747,N_8133,N_7819);
or U8748 (N_8748,N_7854,N_7956);
xnor U8749 (N_8749,N_8118,N_8361);
nand U8750 (N_8750,N_8228,N_7227);
nand U8751 (N_8751,N_7592,N_8042);
nor U8752 (N_8752,N_7311,N_7815);
and U8753 (N_8753,N_7386,N_8268);
nand U8754 (N_8754,N_7475,N_7861);
and U8755 (N_8755,N_7955,N_7875);
xor U8756 (N_8756,N_7266,N_7891);
nand U8757 (N_8757,N_8235,N_7470);
and U8758 (N_8758,N_8233,N_8280);
or U8759 (N_8759,N_7646,N_7778);
or U8760 (N_8760,N_7604,N_8211);
and U8761 (N_8761,N_8058,N_8016);
nor U8762 (N_8762,N_7684,N_7593);
and U8763 (N_8763,N_8018,N_8239);
nor U8764 (N_8764,N_8224,N_8382);
or U8765 (N_8765,N_7576,N_7234);
xnor U8766 (N_8766,N_7909,N_8070);
or U8767 (N_8767,N_7626,N_8345);
and U8768 (N_8768,N_8365,N_7872);
and U8769 (N_8769,N_8370,N_7536);
nand U8770 (N_8770,N_7692,N_7644);
and U8771 (N_8771,N_8184,N_7962);
nor U8772 (N_8772,N_8135,N_7681);
xor U8773 (N_8773,N_8077,N_8265);
or U8774 (N_8774,N_8106,N_7439);
and U8775 (N_8775,N_7613,N_7505);
xor U8776 (N_8776,N_7803,N_8027);
or U8777 (N_8777,N_7366,N_7907);
nand U8778 (N_8778,N_8213,N_8251);
xor U8779 (N_8779,N_8053,N_7471);
and U8780 (N_8780,N_8099,N_8139);
and U8781 (N_8781,N_7596,N_8129);
nor U8782 (N_8782,N_8281,N_7730);
and U8783 (N_8783,N_8104,N_8364);
xnor U8784 (N_8784,N_8389,N_7314);
nor U8785 (N_8785,N_7552,N_8019);
nand U8786 (N_8786,N_7509,N_7356);
nor U8787 (N_8787,N_7208,N_8386);
xor U8788 (N_8788,N_7417,N_7760);
xnor U8789 (N_8789,N_7376,N_7908);
and U8790 (N_8790,N_8153,N_7853);
or U8791 (N_8791,N_7587,N_7460);
or U8792 (N_8792,N_7518,N_7332);
nand U8793 (N_8793,N_8112,N_8217);
and U8794 (N_8794,N_7428,N_7466);
nand U8795 (N_8795,N_8387,N_8040);
xor U8796 (N_8796,N_8012,N_7863);
nor U8797 (N_8797,N_7969,N_7539);
or U8798 (N_8798,N_7977,N_7591);
and U8799 (N_8799,N_8328,N_7453);
xnor U8800 (N_8800,N_7550,N_7310);
nand U8801 (N_8801,N_7675,N_7281);
xor U8802 (N_8802,N_7424,N_8383);
and U8803 (N_8803,N_7978,N_8161);
nor U8804 (N_8804,N_8368,N_7580);
and U8805 (N_8805,N_7480,N_7952);
nand U8806 (N_8806,N_7958,N_8119);
nand U8807 (N_8807,N_7248,N_7672);
xnor U8808 (N_8808,N_7632,N_8084);
nor U8809 (N_8809,N_8171,N_7708);
or U8810 (N_8810,N_7303,N_8362);
xor U8811 (N_8811,N_7582,N_7989);
and U8812 (N_8812,N_8381,N_8388);
nand U8813 (N_8813,N_8020,N_7997);
nand U8814 (N_8814,N_7737,N_7987);
and U8815 (N_8815,N_8260,N_8310);
and U8816 (N_8816,N_7268,N_7957);
nand U8817 (N_8817,N_7633,N_7842);
and U8818 (N_8818,N_8202,N_7789);
nor U8819 (N_8819,N_8287,N_7838);
nand U8820 (N_8820,N_7251,N_7357);
or U8821 (N_8821,N_7472,N_7205);
or U8822 (N_8822,N_7437,N_8083);
nor U8823 (N_8823,N_7537,N_7871);
nor U8824 (N_8824,N_7743,N_7682);
nand U8825 (N_8825,N_7574,N_7981);
nor U8826 (N_8826,N_7538,N_7527);
nand U8827 (N_8827,N_8331,N_7913);
xor U8828 (N_8828,N_7740,N_8060);
or U8829 (N_8829,N_8222,N_7346);
nand U8830 (N_8830,N_7732,N_7603);
nor U8831 (N_8831,N_7499,N_7367);
nor U8832 (N_8832,N_8003,N_7793);
and U8833 (N_8833,N_7623,N_7341);
and U8834 (N_8834,N_7602,N_7716);
and U8835 (N_8835,N_7768,N_8375);
and U8836 (N_8836,N_7283,N_7597);
nor U8837 (N_8837,N_7816,N_7707);
nor U8838 (N_8838,N_8363,N_7848);
xor U8839 (N_8839,N_7855,N_7274);
xor U8840 (N_8840,N_7485,N_7705);
and U8841 (N_8841,N_7757,N_7926);
and U8842 (N_8842,N_7783,N_7516);
or U8843 (N_8843,N_7662,N_7221);
or U8844 (N_8844,N_7494,N_8248);
and U8845 (N_8845,N_8373,N_7300);
nor U8846 (N_8846,N_8343,N_7423);
xnor U8847 (N_8847,N_7551,N_8011);
nand U8848 (N_8848,N_7488,N_7434);
xnor U8849 (N_8849,N_7202,N_8126);
or U8850 (N_8850,N_7796,N_7290);
or U8851 (N_8851,N_7910,N_7272);
xnor U8852 (N_8852,N_8086,N_7565);
xor U8853 (N_8853,N_7306,N_7298);
or U8854 (N_8854,N_7776,N_7881);
or U8855 (N_8855,N_8069,N_8306);
nor U8856 (N_8856,N_7442,N_8107);
nor U8857 (N_8857,N_7831,N_8339);
or U8858 (N_8858,N_7236,N_7377);
and U8859 (N_8859,N_8031,N_7847);
nand U8860 (N_8860,N_7201,N_7630);
or U8861 (N_8861,N_8242,N_7970);
xor U8862 (N_8862,N_8294,N_7523);
and U8863 (N_8863,N_7382,N_7772);
xnor U8864 (N_8864,N_7621,N_7798);
xor U8865 (N_8865,N_7392,N_7846);
nor U8866 (N_8866,N_7345,N_7892);
nand U8867 (N_8867,N_7867,N_8263);
xnor U8868 (N_8868,N_8101,N_7495);
xnor U8869 (N_8869,N_7953,N_7544);
and U8870 (N_8870,N_7792,N_8256);
nor U8871 (N_8871,N_7942,N_8398);
and U8872 (N_8872,N_7207,N_7557);
nor U8873 (N_8873,N_8379,N_8240);
nand U8874 (N_8874,N_7302,N_7770);
xnor U8875 (N_8875,N_7984,N_8262);
or U8876 (N_8876,N_8142,N_8392);
xor U8877 (N_8877,N_7404,N_7901);
or U8878 (N_8878,N_8195,N_7753);
nand U8879 (N_8879,N_8076,N_8023);
nand U8880 (N_8880,N_7775,N_8230);
and U8881 (N_8881,N_8302,N_7914);
xnor U8882 (N_8882,N_8193,N_7966);
and U8883 (N_8883,N_8205,N_8183);
or U8884 (N_8884,N_7709,N_8114);
xor U8885 (N_8885,N_8009,N_8134);
and U8886 (N_8886,N_8143,N_8164);
nand U8887 (N_8887,N_7496,N_7230);
or U8888 (N_8888,N_8210,N_7755);
or U8889 (N_8889,N_7670,N_7276);
nand U8890 (N_8890,N_7661,N_7756);
or U8891 (N_8891,N_7504,N_8100);
xor U8892 (N_8892,N_7359,N_7638);
or U8893 (N_8893,N_7758,N_7588);
and U8894 (N_8894,N_8219,N_7407);
and U8895 (N_8895,N_8284,N_8078);
xor U8896 (N_8896,N_8203,N_7401);
and U8897 (N_8897,N_7394,N_8201);
or U8898 (N_8898,N_7253,N_8366);
or U8899 (N_8899,N_7637,N_8354);
xor U8900 (N_8900,N_7727,N_7693);
nor U8901 (N_8901,N_7548,N_7643);
or U8902 (N_8902,N_7706,N_8255);
nand U8903 (N_8903,N_7741,N_8021);
and U8904 (N_8904,N_8337,N_8187);
and U8905 (N_8905,N_7577,N_7288);
or U8906 (N_8906,N_7534,N_7555);
or U8907 (N_8907,N_7562,N_7818);
or U8908 (N_8908,N_7998,N_8088);
or U8909 (N_8909,N_8324,N_7678);
nand U8910 (N_8910,N_8330,N_8103);
or U8911 (N_8911,N_7336,N_7723);
or U8912 (N_8912,N_7467,N_7403);
nor U8913 (N_8913,N_8300,N_8399);
xnor U8914 (N_8914,N_7954,N_8068);
nor U8915 (N_8915,N_8380,N_7425);
xor U8916 (N_8916,N_7781,N_7950);
nor U8917 (N_8917,N_8340,N_7801);
nand U8918 (N_8918,N_8395,N_8180);
or U8919 (N_8919,N_8051,N_8148);
and U8920 (N_8920,N_7348,N_7317);
and U8921 (N_8921,N_7486,N_8117);
or U8922 (N_8922,N_7697,N_7448);
nand U8923 (N_8923,N_8385,N_7889);
nor U8924 (N_8924,N_8220,N_7639);
nor U8925 (N_8925,N_7762,N_8355);
or U8926 (N_8926,N_7835,N_7994);
or U8927 (N_8927,N_8212,N_7559);
nand U8928 (N_8928,N_7265,N_7438);
or U8929 (N_8929,N_7873,N_7506);
nor U8930 (N_8930,N_8044,N_7935);
or U8931 (N_8931,N_8109,N_8344);
and U8932 (N_8932,N_8391,N_7545);
nor U8933 (N_8933,N_7852,N_7975);
xor U8934 (N_8934,N_7850,N_7687);
and U8935 (N_8935,N_7605,N_7703);
nor U8936 (N_8936,N_8074,N_8352);
nor U8937 (N_8937,N_7905,N_7932);
nand U8938 (N_8938,N_8333,N_7725);
nand U8939 (N_8939,N_8288,N_8225);
nor U8940 (N_8940,N_7304,N_7579);
xnor U8941 (N_8941,N_7515,N_7307);
nand U8942 (N_8942,N_7702,N_7270);
or U8943 (N_8943,N_7244,N_7903);
or U8944 (N_8944,N_7810,N_8000);
xor U8945 (N_8945,N_8111,N_7712);
xnor U8946 (N_8946,N_7650,N_7858);
or U8947 (N_8947,N_8327,N_7578);
nand U8948 (N_8948,N_7351,N_7469);
xor U8949 (N_8949,N_7430,N_8089);
xnor U8950 (N_8950,N_8322,N_7385);
nand U8951 (N_8951,N_8296,N_8059);
or U8952 (N_8952,N_8208,N_7641);
nor U8953 (N_8953,N_8198,N_7983);
xor U8954 (N_8954,N_7900,N_7771);
and U8955 (N_8955,N_7454,N_7885);
and U8956 (N_8956,N_7786,N_7890);
and U8957 (N_8957,N_8303,N_7319);
and U8958 (N_8958,N_7941,N_8188);
xnor U8959 (N_8959,N_8097,N_7334);
nand U8960 (N_8960,N_8321,N_8014);
or U8961 (N_8961,N_8141,N_7328);
and U8962 (N_8962,N_7566,N_7421);
nor U8963 (N_8963,N_7688,N_7916);
xnor U8964 (N_8964,N_8185,N_7292);
or U8965 (N_8965,N_7654,N_8261);
and U8966 (N_8966,N_7371,N_7874);
or U8967 (N_8967,N_7844,N_7503);
xor U8968 (N_8968,N_7507,N_7980);
and U8969 (N_8969,N_7271,N_8006);
or U8970 (N_8970,N_7804,N_8096);
or U8971 (N_8971,N_7280,N_8144);
nor U8972 (N_8972,N_7624,N_7642);
and U8973 (N_8973,N_7679,N_7747);
nand U8974 (N_8974,N_7530,N_7218);
nor U8975 (N_8975,N_8029,N_7262);
nand U8976 (N_8976,N_8291,N_8390);
and U8977 (N_8977,N_7790,N_7685);
nor U8978 (N_8978,N_8221,N_7922);
xnor U8979 (N_8979,N_7599,N_7531);
xor U8980 (N_8980,N_7895,N_7352);
nand U8981 (N_8981,N_7400,N_7763);
or U8982 (N_8982,N_7572,N_7416);
nor U8983 (N_8983,N_8318,N_7384);
nor U8984 (N_8984,N_7841,N_7870);
and U8985 (N_8985,N_7718,N_7286);
xor U8986 (N_8986,N_7749,N_8267);
nand U8987 (N_8987,N_7331,N_7991);
xor U8988 (N_8988,N_7541,N_7520);
nand U8989 (N_8989,N_7754,N_7478);
nor U8990 (N_8990,N_8237,N_7686);
and U8991 (N_8991,N_7673,N_7215);
and U8992 (N_8992,N_7275,N_7479);
and U8993 (N_8993,N_7829,N_7383);
nand U8994 (N_8994,N_7315,N_7893);
nand U8995 (N_8995,N_8283,N_7561);
nand U8996 (N_8996,N_8376,N_7739);
nand U8997 (N_8997,N_7554,N_7484);
or U8998 (N_8998,N_7862,N_7426);
or U8999 (N_8999,N_8025,N_7325);
nand U9000 (N_9000,N_7614,N_8345);
or U9001 (N_9001,N_7262,N_7210);
xnor U9002 (N_9002,N_7293,N_7806);
xnor U9003 (N_9003,N_8200,N_7577);
and U9004 (N_9004,N_7383,N_7823);
or U9005 (N_9005,N_7968,N_8398);
nand U9006 (N_9006,N_8161,N_8297);
and U9007 (N_9007,N_7898,N_8059);
nor U9008 (N_9008,N_8273,N_7636);
and U9009 (N_9009,N_8128,N_8068);
xnor U9010 (N_9010,N_7932,N_7502);
and U9011 (N_9011,N_7464,N_7586);
and U9012 (N_9012,N_7848,N_8115);
or U9013 (N_9013,N_7847,N_7778);
nand U9014 (N_9014,N_8115,N_7661);
xor U9015 (N_9015,N_7629,N_8124);
nor U9016 (N_9016,N_7497,N_7253);
nor U9017 (N_9017,N_8397,N_8169);
and U9018 (N_9018,N_7754,N_7477);
and U9019 (N_9019,N_8041,N_7522);
or U9020 (N_9020,N_7434,N_8039);
or U9021 (N_9021,N_7883,N_7294);
nand U9022 (N_9022,N_7874,N_7221);
nand U9023 (N_9023,N_8377,N_8012);
xor U9024 (N_9024,N_7338,N_8141);
or U9025 (N_9025,N_8024,N_7375);
nand U9026 (N_9026,N_7974,N_7523);
nand U9027 (N_9027,N_8123,N_7456);
or U9028 (N_9028,N_7777,N_7716);
and U9029 (N_9029,N_8161,N_8394);
xor U9030 (N_9030,N_8319,N_8299);
or U9031 (N_9031,N_8219,N_8318);
nor U9032 (N_9032,N_8137,N_7248);
and U9033 (N_9033,N_8152,N_8155);
nor U9034 (N_9034,N_8235,N_7509);
or U9035 (N_9035,N_7559,N_7520);
nor U9036 (N_9036,N_7405,N_7613);
nand U9037 (N_9037,N_7863,N_7959);
and U9038 (N_9038,N_7648,N_7858);
or U9039 (N_9039,N_8211,N_7340);
or U9040 (N_9040,N_7325,N_7389);
nor U9041 (N_9041,N_8302,N_8113);
and U9042 (N_9042,N_8298,N_8184);
or U9043 (N_9043,N_7575,N_8167);
nand U9044 (N_9044,N_7868,N_7458);
and U9045 (N_9045,N_7997,N_8232);
nand U9046 (N_9046,N_8130,N_8333);
nand U9047 (N_9047,N_7882,N_7350);
xnor U9048 (N_9048,N_7908,N_8005);
xor U9049 (N_9049,N_8048,N_8058);
nand U9050 (N_9050,N_8382,N_8212);
or U9051 (N_9051,N_7617,N_7338);
and U9052 (N_9052,N_7377,N_8292);
or U9053 (N_9053,N_7638,N_7305);
nand U9054 (N_9054,N_7992,N_8169);
or U9055 (N_9055,N_8116,N_7221);
or U9056 (N_9056,N_7283,N_7702);
nand U9057 (N_9057,N_8331,N_7445);
nand U9058 (N_9058,N_8187,N_7315);
or U9059 (N_9059,N_7481,N_7474);
xnor U9060 (N_9060,N_7494,N_7402);
xor U9061 (N_9061,N_7435,N_7886);
and U9062 (N_9062,N_7917,N_7669);
nor U9063 (N_9063,N_7466,N_8322);
and U9064 (N_9064,N_7663,N_7423);
nand U9065 (N_9065,N_7836,N_8302);
nor U9066 (N_9066,N_8028,N_8347);
or U9067 (N_9067,N_7532,N_7655);
nor U9068 (N_9068,N_7224,N_7911);
or U9069 (N_9069,N_8317,N_8144);
xnor U9070 (N_9070,N_8092,N_7298);
nor U9071 (N_9071,N_7449,N_7777);
nor U9072 (N_9072,N_7509,N_7284);
xor U9073 (N_9073,N_7839,N_8010);
xor U9074 (N_9074,N_7279,N_7359);
nand U9075 (N_9075,N_7459,N_7563);
xnor U9076 (N_9076,N_7996,N_7424);
xor U9077 (N_9077,N_7885,N_7484);
nor U9078 (N_9078,N_7767,N_8257);
nand U9079 (N_9079,N_7466,N_7667);
and U9080 (N_9080,N_7764,N_8035);
xnor U9081 (N_9081,N_7304,N_7726);
nand U9082 (N_9082,N_7887,N_8386);
nand U9083 (N_9083,N_7860,N_7820);
xnor U9084 (N_9084,N_8176,N_8297);
nor U9085 (N_9085,N_7236,N_7489);
or U9086 (N_9086,N_8022,N_8151);
nand U9087 (N_9087,N_8332,N_8342);
nor U9088 (N_9088,N_7297,N_8051);
nor U9089 (N_9089,N_7696,N_7595);
xor U9090 (N_9090,N_7416,N_7365);
and U9091 (N_9091,N_7850,N_7336);
xnor U9092 (N_9092,N_7717,N_8313);
and U9093 (N_9093,N_7588,N_7663);
nand U9094 (N_9094,N_7334,N_7763);
or U9095 (N_9095,N_7294,N_7779);
nand U9096 (N_9096,N_8030,N_7451);
or U9097 (N_9097,N_7961,N_7299);
or U9098 (N_9098,N_7204,N_7209);
or U9099 (N_9099,N_7980,N_7844);
or U9100 (N_9100,N_8143,N_7588);
nand U9101 (N_9101,N_7510,N_7941);
nor U9102 (N_9102,N_8211,N_7305);
nor U9103 (N_9103,N_7305,N_8267);
or U9104 (N_9104,N_8107,N_8039);
nor U9105 (N_9105,N_8099,N_7247);
nor U9106 (N_9106,N_8198,N_8179);
nand U9107 (N_9107,N_8037,N_7409);
nand U9108 (N_9108,N_7319,N_7462);
nand U9109 (N_9109,N_8271,N_8026);
and U9110 (N_9110,N_8165,N_8336);
xnor U9111 (N_9111,N_8266,N_7239);
or U9112 (N_9112,N_7823,N_7886);
nand U9113 (N_9113,N_7547,N_7638);
nand U9114 (N_9114,N_7216,N_8390);
or U9115 (N_9115,N_7781,N_7886);
or U9116 (N_9116,N_7602,N_8082);
xor U9117 (N_9117,N_7371,N_8053);
or U9118 (N_9118,N_8331,N_7209);
nand U9119 (N_9119,N_7730,N_7841);
xor U9120 (N_9120,N_8247,N_7620);
and U9121 (N_9121,N_8106,N_7367);
or U9122 (N_9122,N_7593,N_7247);
and U9123 (N_9123,N_7492,N_8063);
nand U9124 (N_9124,N_7668,N_7418);
or U9125 (N_9125,N_7693,N_7362);
or U9126 (N_9126,N_7800,N_7395);
xnor U9127 (N_9127,N_7292,N_8111);
nor U9128 (N_9128,N_7697,N_8247);
and U9129 (N_9129,N_8047,N_7780);
and U9130 (N_9130,N_8208,N_7544);
or U9131 (N_9131,N_7866,N_7572);
nand U9132 (N_9132,N_7226,N_8177);
nand U9133 (N_9133,N_7246,N_7690);
or U9134 (N_9134,N_8291,N_7996);
xor U9135 (N_9135,N_7500,N_7847);
nand U9136 (N_9136,N_8349,N_7890);
nand U9137 (N_9137,N_8098,N_7267);
or U9138 (N_9138,N_8312,N_8048);
or U9139 (N_9139,N_8239,N_7648);
or U9140 (N_9140,N_7581,N_7295);
and U9141 (N_9141,N_8354,N_8287);
xor U9142 (N_9142,N_7597,N_8244);
xor U9143 (N_9143,N_8296,N_8240);
nand U9144 (N_9144,N_7243,N_7897);
nor U9145 (N_9145,N_7654,N_7720);
nand U9146 (N_9146,N_7908,N_7392);
xnor U9147 (N_9147,N_7859,N_7597);
xnor U9148 (N_9148,N_7689,N_8137);
xnor U9149 (N_9149,N_7471,N_7414);
or U9150 (N_9150,N_7833,N_8343);
or U9151 (N_9151,N_7391,N_7404);
nand U9152 (N_9152,N_7662,N_8226);
xor U9153 (N_9153,N_7764,N_7781);
or U9154 (N_9154,N_7508,N_8016);
xor U9155 (N_9155,N_8367,N_7520);
xor U9156 (N_9156,N_8037,N_7585);
nand U9157 (N_9157,N_8046,N_7557);
nand U9158 (N_9158,N_7467,N_8394);
nand U9159 (N_9159,N_7585,N_7363);
nand U9160 (N_9160,N_7584,N_8072);
and U9161 (N_9161,N_8324,N_8087);
xnor U9162 (N_9162,N_7385,N_7747);
and U9163 (N_9163,N_7631,N_7938);
xnor U9164 (N_9164,N_7414,N_7347);
nand U9165 (N_9165,N_7582,N_7659);
xor U9166 (N_9166,N_8102,N_8131);
and U9167 (N_9167,N_7415,N_7462);
or U9168 (N_9168,N_7707,N_7690);
or U9169 (N_9169,N_8282,N_7453);
xor U9170 (N_9170,N_7550,N_7440);
nor U9171 (N_9171,N_7882,N_8176);
nor U9172 (N_9172,N_7811,N_7301);
xnor U9173 (N_9173,N_7738,N_7296);
xnor U9174 (N_9174,N_8328,N_8028);
nor U9175 (N_9175,N_7612,N_8178);
nor U9176 (N_9176,N_7657,N_8076);
or U9177 (N_9177,N_7774,N_7703);
or U9178 (N_9178,N_7560,N_7832);
xnor U9179 (N_9179,N_7260,N_8203);
nand U9180 (N_9180,N_7477,N_7991);
and U9181 (N_9181,N_7432,N_7806);
and U9182 (N_9182,N_7778,N_7355);
nor U9183 (N_9183,N_7404,N_7872);
or U9184 (N_9184,N_7496,N_7239);
xnor U9185 (N_9185,N_7505,N_7577);
nor U9186 (N_9186,N_8241,N_7222);
or U9187 (N_9187,N_7605,N_7602);
nand U9188 (N_9188,N_7703,N_7319);
or U9189 (N_9189,N_7208,N_7533);
nand U9190 (N_9190,N_8392,N_8002);
nor U9191 (N_9191,N_7661,N_8194);
nand U9192 (N_9192,N_7740,N_7954);
xor U9193 (N_9193,N_7573,N_8218);
or U9194 (N_9194,N_7896,N_7213);
or U9195 (N_9195,N_7456,N_7231);
xor U9196 (N_9196,N_7336,N_7821);
xnor U9197 (N_9197,N_8247,N_8232);
nand U9198 (N_9198,N_7984,N_7458);
nor U9199 (N_9199,N_7238,N_8258);
nand U9200 (N_9200,N_7793,N_7688);
and U9201 (N_9201,N_7877,N_8268);
nor U9202 (N_9202,N_7870,N_8303);
xor U9203 (N_9203,N_7919,N_7451);
or U9204 (N_9204,N_8134,N_7737);
and U9205 (N_9205,N_7351,N_8333);
or U9206 (N_9206,N_7984,N_7731);
nor U9207 (N_9207,N_7633,N_7261);
or U9208 (N_9208,N_8050,N_7536);
nor U9209 (N_9209,N_7788,N_8269);
and U9210 (N_9210,N_7731,N_8002);
xnor U9211 (N_9211,N_7843,N_7882);
and U9212 (N_9212,N_7704,N_8075);
xor U9213 (N_9213,N_7204,N_7245);
nor U9214 (N_9214,N_7352,N_8245);
and U9215 (N_9215,N_7353,N_8223);
xnor U9216 (N_9216,N_8248,N_8095);
or U9217 (N_9217,N_7837,N_7786);
xnor U9218 (N_9218,N_7235,N_7515);
xor U9219 (N_9219,N_8399,N_8180);
nor U9220 (N_9220,N_8270,N_7402);
or U9221 (N_9221,N_7383,N_8005);
nor U9222 (N_9222,N_7710,N_8189);
nand U9223 (N_9223,N_8090,N_8169);
and U9224 (N_9224,N_8363,N_7241);
or U9225 (N_9225,N_8279,N_7530);
nor U9226 (N_9226,N_7527,N_7994);
nor U9227 (N_9227,N_8336,N_8221);
or U9228 (N_9228,N_7933,N_7428);
or U9229 (N_9229,N_7512,N_7842);
nor U9230 (N_9230,N_8032,N_7810);
or U9231 (N_9231,N_7558,N_7890);
nand U9232 (N_9232,N_8110,N_7261);
nor U9233 (N_9233,N_7218,N_7554);
or U9234 (N_9234,N_7826,N_7667);
nor U9235 (N_9235,N_8283,N_8140);
xnor U9236 (N_9236,N_8311,N_7489);
nand U9237 (N_9237,N_8316,N_7980);
nand U9238 (N_9238,N_7527,N_8383);
or U9239 (N_9239,N_7332,N_8243);
or U9240 (N_9240,N_7466,N_7268);
or U9241 (N_9241,N_7842,N_7981);
or U9242 (N_9242,N_7233,N_7755);
xnor U9243 (N_9243,N_7548,N_8071);
nor U9244 (N_9244,N_8349,N_8022);
and U9245 (N_9245,N_7967,N_7296);
nor U9246 (N_9246,N_7583,N_7739);
or U9247 (N_9247,N_7303,N_7253);
nor U9248 (N_9248,N_8287,N_7728);
xnor U9249 (N_9249,N_7577,N_7900);
or U9250 (N_9250,N_7495,N_8277);
nand U9251 (N_9251,N_8232,N_7233);
nand U9252 (N_9252,N_7860,N_7420);
xor U9253 (N_9253,N_7640,N_7443);
or U9254 (N_9254,N_7735,N_8344);
and U9255 (N_9255,N_7962,N_7446);
and U9256 (N_9256,N_7325,N_7730);
and U9257 (N_9257,N_7939,N_7253);
and U9258 (N_9258,N_7481,N_7663);
nor U9259 (N_9259,N_8163,N_7884);
nand U9260 (N_9260,N_7763,N_7607);
or U9261 (N_9261,N_7575,N_7556);
nand U9262 (N_9262,N_7702,N_7410);
and U9263 (N_9263,N_7831,N_7238);
or U9264 (N_9264,N_8166,N_8223);
nor U9265 (N_9265,N_8076,N_7458);
and U9266 (N_9266,N_7267,N_8241);
and U9267 (N_9267,N_8364,N_8342);
nand U9268 (N_9268,N_7430,N_7893);
and U9269 (N_9269,N_7671,N_7978);
nor U9270 (N_9270,N_8004,N_8386);
and U9271 (N_9271,N_7962,N_7603);
or U9272 (N_9272,N_7587,N_7483);
nor U9273 (N_9273,N_7538,N_8153);
nor U9274 (N_9274,N_8268,N_7268);
and U9275 (N_9275,N_7303,N_8282);
nand U9276 (N_9276,N_7800,N_7235);
or U9277 (N_9277,N_8357,N_7919);
nand U9278 (N_9278,N_7730,N_7525);
and U9279 (N_9279,N_7255,N_7201);
or U9280 (N_9280,N_7256,N_8000);
xnor U9281 (N_9281,N_8085,N_7706);
nand U9282 (N_9282,N_7818,N_7493);
nor U9283 (N_9283,N_7611,N_7881);
or U9284 (N_9284,N_7630,N_8260);
nand U9285 (N_9285,N_8334,N_7257);
and U9286 (N_9286,N_7682,N_7728);
and U9287 (N_9287,N_7488,N_8076);
and U9288 (N_9288,N_8358,N_7424);
nand U9289 (N_9289,N_7628,N_8279);
nand U9290 (N_9290,N_8301,N_8026);
and U9291 (N_9291,N_7592,N_7298);
nor U9292 (N_9292,N_7616,N_7260);
nand U9293 (N_9293,N_7448,N_7560);
xor U9294 (N_9294,N_7489,N_8148);
and U9295 (N_9295,N_7246,N_7374);
and U9296 (N_9296,N_7581,N_7554);
xor U9297 (N_9297,N_7278,N_8023);
or U9298 (N_9298,N_7886,N_7788);
xor U9299 (N_9299,N_8219,N_7362);
and U9300 (N_9300,N_7573,N_8378);
xnor U9301 (N_9301,N_8327,N_7507);
xnor U9302 (N_9302,N_7222,N_7616);
nand U9303 (N_9303,N_7990,N_7539);
xor U9304 (N_9304,N_7698,N_7502);
nand U9305 (N_9305,N_7204,N_7593);
nor U9306 (N_9306,N_7523,N_7495);
nor U9307 (N_9307,N_7211,N_8038);
nand U9308 (N_9308,N_7544,N_7992);
nand U9309 (N_9309,N_7719,N_7762);
nand U9310 (N_9310,N_8189,N_8171);
and U9311 (N_9311,N_8068,N_7763);
xnor U9312 (N_9312,N_8242,N_7357);
and U9313 (N_9313,N_7914,N_7844);
nor U9314 (N_9314,N_7928,N_8204);
or U9315 (N_9315,N_8379,N_7258);
or U9316 (N_9316,N_7266,N_7508);
xor U9317 (N_9317,N_7697,N_7772);
nor U9318 (N_9318,N_8147,N_7562);
nor U9319 (N_9319,N_7429,N_7486);
nor U9320 (N_9320,N_7910,N_7258);
or U9321 (N_9321,N_7603,N_7672);
nor U9322 (N_9322,N_8084,N_7654);
xor U9323 (N_9323,N_7518,N_7531);
and U9324 (N_9324,N_7748,N_7659);
nand U9325 (N_9325,N_8009,N_7282);
or U9326 (N_9326,N_7338,N_8340);
xor U9327 (N_9327,N_7272,N_7808);
nor U9328 (N_9328,N_7477,N_7446);
nand U9329 (N_9329,N_7866,N_8014);
and U9330 (N_9330,N_8377,N_8151);
nor U9331 (N_9331,N_7852,N_7204);
or U9332 (N_9332,N_8026,N_7494);
nand U9333 (N_9333,N_7377,N_7742);
nor U9334 (N_9334,N_7582,N_7952);
and U9335 (N_9335,N_7858,N_8004);
or U9336 (N_9336,N_8225,N_7280);
or U9337 (N_9337,N_7325,N_7864);
nand U9338 (N_9338,N_7944,N_8270);
nand U9339 (N_9339,N_7357,N_7845);
nor U9340 (N_9340,N_8250,N_8295);
xor U9341 (N_9341,N_7626,N_7543);
xnor U9342 (N_9342,N_7600,N_7812);
nor U9343 (N_9343,N_7744,N_7762);
xnor U9344 (N_9344,N_7380,N_8385);
xor U9345 (N_9345,N_7282,N_8189);
and U9346 (N_9346,N_7320,N_7637);
xor U9347 (N_9347,N_7339,N_7818);
or U9348 (N_9348,N_7335,N_8372);
xnor U9349 (N_9349,N_8136,N_7466);
or U9350 (N_9350,N_8308,N_7476);
nor U9351 (N_9351,N_7271,N_8356);
and U9352 (N_9352,N_8317,N_7274);
nor U9353 (N_9353,N_7241,N_7851);
nor U9354 (N_9354,N_7441,N_7801);
nand U9355 (N_9355,N_7330,N_7300);
nor U9356 (N_9356,N_8348,N_7205);
xor U9357 (N_9357,N_7809,N_7578);
nand U9358 (N_9358,N_8108,N_8192);
and U9359 (N_9359,N_8002,N_7285);
and U9360 (N_9360,N_7917,N_7919);
and U9361 (N_9361,N_8369,N_7717);
nand U9362 (N_9362,N_7696,N_7495);
and U9363 (N_9363,N_8377,N_7864);
and U9364 (N_9364,N_7746,N_7952);
nand U9365 (N_9365,N_8271,N_7900);
xnor U9366 (N_9366,N_7691,N_7320);
or U9367 (N_9367,N_8212,N_7859);
nor U9368 (N_9368,N_8211,N_7470);
and U9369 (N_9369,N_8048,N_8243);
nand U9370 (N_9370,N_8131,N_8074);
or U9371 (N_9371,N_7909,N_7607);
nor U9372 (N_9372,N_7488,N_8005);
and U9373 (N_9373,N_7705,N_8020);
and U9374 (N_9374,N_7373,N_7609);
nor U9375 (N_9375,N_7463,N_7786);
or U9376 (N_9376,N_7488,N_7590);
xor U9377 (N_9377,N_7253,N_7302);
nor U9378 (N_9378,N_7815,N_8260);
and U9379 (N_9379,N_8003,N_8225);
nor U9380 (N_9380,N_7517,N_7619);
or U9381 (N_9381,N_7439,N_7975);
or U9382 (N_9382,N_8265,N_8266);
nor U9383 (N_9383,N_7524,N_7801);
nand U9384 (N_9384,N_7751,N_7558);
and U9385 (N_9385,N_8262,N_8326);
or U9386 (N_9386,N_7697,N_8357);
and U9387 (N_9387,N_7647,N_8053);
nand U9388 (N_9388,N_8238,N_7672);
xnor U9389 (N_9389,N_7789,N_7447);
and U9390 (N_9390,N_8126,N_8208);
xnor U9391 (N_9391,N_7919,N_8144);
xnor U9392 (N_9392,N_7631,N_7366);
or U9393 (N_9393,N_8389,N_7454);
xor U9394 (N_9394,N_8168,N_8068);
xnor U9395 (N_9395,N_8354,N_7983);
nor U9396 (N_9396,N_7430,N_7568);
nor U9397 (N_9397,N_7566,N_7717);
nor U9398 (N_9398,N_8270,N_8081);
xor U9399 (N_9399,N_8387,N_7302);
or U9400 (N_9400,N_7906,N_8035);
nor U9401 (N_9401,N_7639,N_8256);
nor U9402 (N_9402,N_8127,N_7213);
nand U9403 (N_9403,N_7726,N_7778);
or U9404 (N_9404,N_7692,N_7717);
or U9405 (N_9405,N_7608,N_7951);
and U9406 (N_9406,N_7739,N_8016);
xnor U9407 (N_9407,N_7827,N_7288);
nand U9408 (N_9408,N_7800,N_7350);
nand U9409 (N_9409,N_8342,N_7827);
nand U9410 (N_9410,N_8178,N_7534);
or U9411 (N_9411,N_7697,N_8299);
xor U9412 (N_9412,N_7441,N_7479);
nand U9413 (N_9413,N_8203,N_7230);
or U9414 (N_9414,N_8093,N_7596);
or U9415 (N_9415,N_7217,N_8265);
and U9416 (N_9416,N_7703,N_7527);
xor U9417 (N_9417,N_8303,N_8330);
xnor U9418 (N_9418,N_8318,N_8141);
nor U9419 (N_9419,N_7225,N_8085);
and U9420 (N_9420,N_7595,N_7265);
nor U9421 (N_9421,N_7762,N_7583);
nor U9422 (N_9422,N_7897,N_7829);
nor U9423 (N_9423,N_7964,N_7458);
nor U9424 (N_9424,N_8002,N_8323);
and U9425 (N_9425,N_8321,N_7290);
or U9426 (N_9426,N_7863,N_7953);
nor U9427 (N_9427,N_8320,N_8280);
nand U9428 (N_9428,N_8022,N_7860);
or U9429 (N_9429,N_7310,N_8020);
or U9430 (N_9430,N_7426,N_7268);
nand U9431 (N_9431,N_7412,N_7829);
nand U9432 (N_9432,N_7358,N_7858);
nand U9433 (N_9433,N_7296,N_7513);
xor U9434 (N_9434,N_7765,N_7406);
and U9435 (N_9435,N_8118,N_7874);
and U9436 (N_9436,N_7423,N_8192);
xnor U9437 (N_9437,N_7937,N_7313);
or U9438 (N_9438,N_7406,N_7531);
or U9439 (N_9439,N_8035,N_8376);
and U9440 (N_9440,N_7796,N_7694);
nor U9441 (N_9441,N_7988,N_8284);
or U9442 (N_9442,N_7862,N_7673);
and U9443 (N_9443,N_7772,N_7963);
and U9444 (N_9444,N_7576,N_7480);
or U9445 (N_9445,N_7498,N_7619);
nor U9446 (N_9446,N_8068,N_7557);
nand U9447 (N_9447,N_7594,N_8139);
or U9448 (N_9448,N_7381,N_7393);
nor U9449 (N_9449,N_7954,N_7566);
nand U9450 (N_9450,N_8307,N_7930);
xor U9451 (N_9451,N_7751,N_8015);
or U9452 (N_9452,N_8037,N_8199);
and U9453 (N_9453,N_7300,N_7327);
nand U9454 (N_9454,N_7524,N_8121);
nor U9455 (N_9455,N_7302,N_8126);
and U9456 (N_9456,N_7891,N_7771);
or U9457 (N_9457,N_7620,N_7549);
nand U9458 (N_9458,N_7702,N_8342);
nor U9459 (N_9459,N_8179,N_7499);
nand U9460 (N_9460,N_8261,N_7944);
xor U9461 (N_9461,N_7241,N_7849);
nand U9462 (N_9462,N_7703,N_7968);
nor U9463 (N_9463,N_8385,N_8187);
nand U9464 (N_9464,N_7747,N_7692);
or U9465 (N_9465,N_7729,N_7924);
nand U9466 (N_9466,N_8052,N_7354);
xnor U9467 (N_9467,N_8359,N_7701);
nand U9468 (N_9468,N_7507,N_8118);
nor U9469 (N_9469,N_7502,N_7756);
or U9470 (N_9470,N_7315,N_7848);
nand U9471 (N_9471,N_7201,N_7358);
and U9472 (N_9472,N_7610,N_7450);
or U9473 (N_9473,N_8215,N_7315);
xnor U9474 (N_9474,N_7418,N_7316);
nand U9475 (N_9475,N_8136,N_7885);
nor U9476 (N_9476,N_7573,N_7353);
xnor U9477 (N_9477,N_8023,N_7441);
nand U9478 (N_9478,N_8373,N_7478);
xor U9479 (N_9479,N_7493,N_7925);
and U9480 (N_9480,N_8058,N_7564);
or U9481 (N_9481,N_8078,N_7464);
and U9482 (N_9482,N_8135,N_8104);
or U9483 (N_9483,N_8218,N_8282);
nand U9484 (N_9484,N_8341,N_7847);
nor U9485 (N_9485,N_8015,N_7383);
nor U9486 (N_9486,N_7296,N_7408);
or U9487 (N_9487,N_7831,N_7224);
or U9488 (N_9488,N_8054,N_7841);
xor U9489 (N_9489,N_7674,N_8376);
xor U9490 (N_9490,N_7615,N_7941);
xnor U9491 (N_9491,N_7680,N_8124);
nor U9492 (N_9492,N_7618,N_7297);
and U9493 (N_9493,N_7332,N_7721);
or U9494 (N_9494,N_7774,N_7275);
nor U9495 (N_9495,N_8203,N_7274);
nand U9496 (N_9496,N_7943,N_7737);
or U9497 (N_9497,N_7511,N_7849);
or U9498 (N_9498,N_7813,N_7788);
nand U9499 (N_9499,N_8305,N_7944);
xor U9500 (N_9500,N_8019,N_8010);
and U9501 (N_9501,N_8331,N_8110);
or U9502 (N_9502,N_8319,N_7955);
and U9503 (N_9503,N_7924,N_7750);
xor U9504 (N_9504,N_8176,N_7962);
or U9505 (N_9505,N_8289,N_8341);
nor U9506 (N_9506,N_8092,N_8276);
or U9507 (N_9507,N_7636,N_7308);
xnor U9508 (N_9508,N_7819,N_7798);
xor U9509 (N_9509,N_8087,N_8238);
or U9510 (N_9510,N_7931,N_7705);
or U9511 (N_9511,N_7951,N_7302);
nor U9512 (N_9512,N_8161,N_7949);
nand U9513 (N_9513,N_7613,N_8294);
xor U9514 (N_9514,N_7508,N_7544);
nand U9515 (N_9515,N_8190,N_7539);
xnor U9516 (N_9516,N_7696,N_7832);
nand U9517 (N_9517,N_8036,N_7910);
xor U9518 (N_9518,N_7863,N_8140);
or U9519 (N_9519,N_7790,N_8364);
xnor U9520 (N_9520,N_7889,N_7888);
xor U9521 (N_9521,N_8262,N_7702);
xnor U9522 (N_9522,N_8033,N_7941);
nand U9523 (N_9523,N_7263,N_7398);
nand U9524 (N_9524,N_7553,N_7242);
nor U9525 (N_9525,N_7657,N_7960);
or U9526 (N_9526,N_8141,N_7371);
and U9527 (N_9527,N_8267,N_8386);
nand U9528 (N_9528,N_8369,N_8198);
nand U9529 (N_9529,N_8370,N_8006);
nor U9530 (N_9530,N_7412,N_7394);
nand U9531 (N_9531,N_7378,N_7302);
nand U9532 (N_9532,N_8398,N_7271);
and U9533 (N_9533,N_7424,N_7993);
nand U9534 (N_9534,N_8259,N_8103);
nor U9535 (N_9535,N_8324,N_7843);
nor U9536 (N_9536,N_8200,N_8058);
nor U9537 (N_9537,N_8309,N_7850);
nor U9538 (N_9538,N_7405,N_7482);
nor U9539 (N_9539,N_8254,N_7842);
and U9540 (N_9540,N_7518,N_8330);
and U9541 (N_9541,N_8107,N_7496);
and U9542 (N_9542,N_7943,N_8122);
and U9543 (N_9543,N_7496,N_8281);
xnor U9544 (N_9544,N_7435,N_7312);
and U9545 (N_9545,N_8381,N_7474);
nor U9546 (N_9546,N_8263,N_7228);
nor U9547 (N_9547,N_8041,N_8308);
or U9548 (N_9548,N_7875,N_7356);
or U9549 (N_9549,N_7945,N_8200);
nor U9550 (N_9550,N_7220,N_7554);
or U9551 (N_9551,N_7655,N_7592);
or U9552 (N_9552,N_7907,N_7946);
or U9553 (N_9553,N_8086,N_7461);
nand U9554 (N_9554,N_8158,N_7797);
nor U9555 (N_9555,N_8220,N_8314);
xor U9556 (N_9556,N_8126,N_8363);
xor U9557 (N_9557,N_7645,N_7649);
or U9558 (N_9558,N_8277,N_8105);
xnor U9559 (N_9559,N_7286,N_8203);
nand U9560 (N_9560,N_7371,N_8257);
nand U9561 (N_9561,N_7549,N_7794);
or U9562 (N_9562,N_7734,N_8350);
or U9563 (N_9563,N_8392,N_7870);
xor U9564 (N_9564,N_8005,N_7482);
nor U9565 (N_9565,N_7727,N_7752);
nand U9566 (N_9566,N_7560,N_8038);
nand U9567 (N_9567,N_7899,N_8125);
xnor U9568 (N_9568,N_7443,N_7211);
nand U9569 (N_9569,N_8348,N_7616);
nand U9570 (N_9570,N_8262,N_8227);
and U9571 (N_9571,N_7830,N_7894);
nor U9572 (N_9572,N_8133,N_7955);
xnor U9573 (N_9573,N_8177,N_7335);
nor U9574 (N_9574,N_8012,N_7330);
and U9575 (N_9575,N_8063,N_8282);
or U9576 (N_9576,N_8153,N_7279);
nor U9577 (N_9577,N_8369,N_8264);
nor U9578 (N_9578,N_7253,N_7382);
nand U9579 (N_9579,N_7538,N_7413);
and U9580 (N_9580,N_8080,N_8061);
and U9581 (N_9581,N_8397,N_7550);
or U9582 (N_9582,N_8142,N_7283);
and U9583 (N_9583,N_7496,N_8256);
nor U9584 (N_9584,N_8374,N_7767);
or U9585 (N_9585,N_7562,N_8287);
and U9586 (N_9586,N_7707,N_7980);
or U9587 (N_9587,N_8029,N_8086);
nor U9588 (N_9588,N_7711,N_8061);
or U9589 (N_9589,N_8227,N_8253);
nand U9590 (N_9590,N_8304,N_8320);
or U9591 (N_9591,N_8211,N_7600);
nand U9592 (N_9592,N_7902,N_7775);
nand U9593 (N_9593,N_7544,N_8376);
nor U9594 (N_9594,N_7426,N_7851);
and U9595 (N_9595,N_7400,N_8071);
nand U9596 (N_9596,N_7534,N_7860);
and U9597 (N_9597,N_8272,N_8304);
nor U9598 (N_9598,N_8086,N_7950);
nor U9599 (N_9599,N_7232,N_7420);
and U9600 (N_9600,N_9461,N_9051);
nor U9601 (N_9601,N_8701,N_8617);
xor U9602 (N_9602,N_9441,N_9542);
nand U9603 (N_9603,N_8655,N_9075);
xor U9604 (N_9604,N_9270,N_9220);
or U9605 (N_9605,N_9264,N_9336);
or U9606 (N_9606,N_9546,N_9415);
or U9607 (N_9607,N_9295,N_9044);
xnor U9608 (N_9608,N_8431,N_8440);
nor U9609 (N_9609,N_9057,N_8918);
or U9610 (N_9610,N_8709,N_8848);
or U9611 (N_9611,N_8559,N_9133);
or U9612 (N_9612,N_9320,N_8909);
nand U9613 (N_9613,N_8621,N_9055);
nor U9614 (N_9614,N_8726,N_9413);
xor U9615 (N_9615,N_8411,N_8402);
nor U9616 (N_9616,N_9585,N_9377);
nand U9617 (N_9617,N_8523,N_8610);
nor U9618 (N_9618,N_9218,N_8419);
nor U9619 (N_9619,N_9189,N_8682);
nor U9620 (N_9620,N_8849,N_8647);
nor U9621 (N_9621,N_9383,N_9102);
nand U9622 (N_9622,N_8817,N_8512);
and U9623 (N_9623,N_8824,N_8988);
and U9624 (N_9624,N_8550,N_8683);
xnor U9625 (N_9625,N_9513,N_9175);
nor U9626 (N_9626,N_8977,N_9274);
and U9627 (N_9627,N_9293,N_9229);
xnor U9628 (N_9628,N_9346,N_9560);
or U9629 (N_9629,N_8964,N_9471);
nor U9630 (N_9630,N_8777,N_8873);
or U9631 (N_9631,N_8915,N_8519);
and U9632 (N_9632,N_9187,N_8775);
nor U9633 (N_9633,N_8906,N_9242);
and U9634 (N_9634,N_9458,N_8857);
and U9635 (N_9635,N_9532,N_9420);
and U9636 (N_9636,N_9540,N_8566);
xnor U9637 (N_9637,N_8955,N_9446);
or U9638 (N_9638,N_9043,N_9317);
xor U9639 (N_9639,N_8643,N_9314);
or U9640 (N_9640,N_8913,N_9036);
nand U9641 (N_9641,N_8724,N_8965);
xor U9642 (N_9642,N_9062,N_8416);
nand U9643 (N_9643,N_9160,N_9351);
xor U9644 (N_9644,N_8804,N_8876);
nor U9645 (N_9645,N_9076,N_9165);
or U9646 (N_9646,N_9506,N_8771);
or U9647 (N_9647,N_8920,N_9039);
or U9648 (N_9648,N_9168,N_9271);
or U9649 (N_9649,N_8493,N_8813);
and U9650 (N_9650,N_9490,N_8819);
nor U9651 (N_9651,N_9400,N_8469);
nor U9652 (N_9652,N_8535,N_8719);
nand U9653 (N_9653,N_8993,N_9027);
and U9654 (N_9654,N_9276,N_9502);
xnor U9655 (N_9655,N_9469,N_8592);
xnor U9656 (N_9656,N_8407,N_9308);
xor U9657 (N_9657,N_8596,N_8705);
and U9658 (N_9658,N_9111,N_9499);
nor U9659 (N_9659,N_9593,N_9553);
or U9660 (N_9660,N_8979,N_8880);
or U9661 (N_9661,N_8616,N_9018);
xnor U9662 (N_9662,N_8486,N_8805);
nand U9663 (N_9663,N_9578,N_9070);
and U9664 (N_9664,N_9121,N_9100);
or U9665 (N_9665,N_9065,N_9092);
and U9666 (N_9666,N_9485,N_9060);
xnor U9667 (N_9667,N_9564,N_8862);
nor U9668 (N_9668,N_9598,N_8738);
nor U9669 (N_9669,N_8432,N_8967);
nand U9670 (N_9670,N_9170,N_8676);
nor U9671 (N_9671,N_8941,N_8811);
and U9672 (N_9672,N_9365,N_8947);
and U9673 (N_9673,N_8867,N_8894);
or U9674 (N_9674,N_8501,N_9040);
and U9675 (N_9675,N_9211,N_9422);
and U9676 (N_9676,N_8445,N_9402);
nand U9677 (N_9677,N_8664,N_9522);
xnor U9678 (N_9678,N_8442,N_9486);
nor U9679 (N_9679,N_8450,N_9479);
and U9680 (N_9680,N_9209,N_9307);
nand U9681 (N_9681,N_9385,N_8842);
or U9682 (N_9682,N_8882,N_8496);
or U9683 (N_9683,N_8418,N_8905);
xor U9684 (N_9684,N_8956,N_9398);
or U9685 (N_9685,N_8879,N_9186);
nor U9686 (N_9686,N_8503,N_9073);
xnor U9687 (N_9687,N_8627,N_8716);
nand U9688 (N_9688,N_9436,N_9159);
nor U9689 (N_9689,N_8604,N_9541);
nand U9690 (N_9690,N_9219,N_8925);
nand U9691 (N_9691,N_9054,N_9419);
nand U9692 (N_9692,N_9200,N_9533);
nor U9693 (N_9693,N_9590,N_9334);
and U9694 (N_9694,N_8448,N_9306);
nand U9695 (N_9695,N_9266,N_9103);
nand U9696 (N_9696,N_8755,N_9529);
nor U9697 (N_9697,N_8723,N_9583);
nand U9698 (N_9698,N_8669,N_8489);
and U9699 (N_9699,N_9491,N_8721);
or U9700 (N_9700,N_8620,N_9562);
xnor U9701 (N_9701,N_8659,N_9496);
or U9702 (N_9702,N_9205,N_9514);
and U9703 (N_9703,N_8999,N_8573);
nor U9704 (N_9704,N_8498,N_9355);
and U9705 (N_9705,N_8679,N_8688);
and U9706 (N_9706,N_9114,N_8973);
nand U9707 (N_9707,N_8516,N_8495);
and U9708 (N_9708,N_8585,N_9592);
nor U9709 (N_9709,N_8533,N_9120);
or U9710 (N_9710,N_8983,N_8417);
nor U9711 (N_9711,N_9179,N_8969);
nor U9712 (N_9712,N_9025,N_8704);
or U9713 (N_9713,N_9528,N_9369);
and U9714 (N_9714,N_9580,N_9526);
and U9715 (N_9715,N_9575,N_9118);
nand U9716 (N_9716,N_9589,N_8991);
and U9717 (N_9717,N_9058,N_8549);
xnor U9718 (N_9718,N_8751,N_8608);
or U9719 (N_9719,N_8789,N_8995);
or U9720 (N_9720,N_9408,N_9428);
xor U9721 (N_9721,N_8644,N_9315);
nor U9722 (N_9722,N_8818,N_9232);
or U9723 (N_9723,N_8713,N_9136);
and U9724 (N_9724,N_8479,N_9344);
or U9725 (N_9725,N_8797,N_8639);
xnor U9726 (N_9726,N_9586,N_9239);
and U9727 (N_9727,N_8878,N_8695);
or U9728 (N_9728,N_8974,N_8544);
xor U9729 (N_9729,N_9341,N_8997);
nor U9730 (N_9730,N_9433,N_9374);
and U9731 (N_9731,N_9582,N_8808);
nand U9732 (N_9732,N_9228,N_8899);
and U9733 (N_9733,N_8594,N_9443);
xor U9734 (N_9734,N_8685,N_9156);
or U9735 (N_9735,N_8707,N_9566);
nor U9736 (N_9736,N_9366,N_9280);
and U9737 (N_9737,N_9152,N_9362);
or U9738 (N_9738,N_8600,N_8844);
or U9739 (N_9739,N_8574,N_8892);
nor U9740 (N_9740,N_9305,N_9390);
and U9741 (N_9741,N_9333,N_8746);
and U9742 (N_9742,N_8641,N_9403);
nor U9743 (N_9743,N_9157,N_8624);
and U9744 (N_9744,N_8992,N_8770);
nand U9745 (N_9745,N_8400,N_9448);
or U9746 (N_9746,N_8952,N_9524);
or U9747 (N_9747,N_9064,N_8891);
xor U9748 (N_9748,N_8959,N_8858);
or U9749 (N_9749,N_9534,N_8868);
nand U9750 (N_9750,N_8931,N_8401);
nand U9751 (N_9751,N_9131,N_9122);
nor U9752 (N_9752,N_9049,N_8658);
and U9753 (N_9753,N_9453,N_8437);
or U9754 (N_9754,N_8843,N_9337);
nand U9755 (N_9755,N_9389,N_8531);
and U9756 (N_9756,N_9031,N_8874);
nand U9757 (N_9757,N_8829,N_8485);
nor U9758 (N_9758,N_9345,N_8500);
xor U9759 (N_9759,N_8505,N_9154);
or U9760 (N_9760,N_8949,N_8917);
or U9761 (N_9761,N_9278,N_8452);
or U9762 (N_9762,N_9105,N_9263);
or U9763 (N_9763,N_9384,N_8927);
nor U9764 (N_9764,N_8403,N_8786);
xor U9765 (N_9765,N_9254,N_9097);
xor U9766 (N_9766,N_9370,N_9387);
nor U9767 (N_9767,N_8730,N_9304);
nand U9768 (N_9768,N_9032,N_9137);
nand U9769 (N_9769,N_9361,N_8727);
nor U9770 (N_9770,N_8904,N_9301);
and U9771 (N_9771,N_9193,N_9162);
or U9772 (N_9772,N_8473,N_8888);
nand U9773 (N_9773,N_8686,N_8565);
or U9774 (N_9774,N_8845,N_9382);
nor U9775 (N_9775,N_8853,N_8561);
nor U9776 (N_9776,N_8653,N_8657);
xnor U9777 (N_9777,N_9026,N_8762);
or U9778 (N_9778,N_8740,N_8532);
or U9779 (N_9779,N_8936,N_8546);
nand U9780 (N_9780,N_9584,N_9376);
xnor U9781 (N_9781,N_8663,N_9130);
and U9782 (N_9782,N_8728,N_8996);
nand U9783 (N_9783,N_9262,N_9392);
xnor U9784 (N_9784,N_9299,N_8856);
or U9785 (N_9785,N_9041,N_8515);
xor U9786 (N_9786,N_8924,N_9191);
nand U9787 (N_9787,N_8839,N_8788);
nor U9788 (N_9788,N_8636,N_9368);
xnor U9789 (N_9789,N_8687,N_8812);
nand U9790 (N_9790,N_8563,N_8773);
xor U9791 (N_9791,N_9116,N_8692);
and U9792 (N_9792,N_9017,N_8735);
xnor U9793 (N_9793,N_8816,N_8897);
nor U9794 (N_9794,N_8612,N_9451);
or U9795 (N_9795,N_8433,N_9466);
and U9796 (N_9796,N_9284,N_9520);
and U9797 (N_9797,N_8810,N_9285);
xor U9798 (N_9798,N_8926,N_8938);
xnor U9799 (N_9799,N_8932,N_9056);
and U9800 (N_9800,N_9255,N_9406);
nand U9801 (N_9801,N_8598,N_9570);
or U9802 (N_9802,N_8630,N_8711);
and U9803 (N_9803,N_8425,N_8739);
xnor U9804 (N_9804,N_8944,N_9321);
xnor U9805 (N_9805,N_8784,N_8722);
and U9806 (N_9806,N_9367,N_8801);
xor U9807 (N_9807,N_8534,N_8953);
or U9808 (N_9808,N_9016,N_8492);
xnor U9809 (N_9809,N_9573,N_8745);
or U9810 (N_9810,N_9082,N_8556);
nor U9811 (N_9811,N_9417,N_9350);
nand U9812 (N_9812,N_8741,N_9335);
nor U9813 (N_9813,N_8649,N_9201);
or U9814 (N_9814,N_9459,N_9343);
nand U9815 (N_9815,N_8970,N_9147);
nor U9816 (N_9816,N_8584,N_8677);
nor U9817 (N_9817,N_9005,N_8475);
nor U9818 (N_9818,N_8444,N_8852);
nor U9819 (N_9819,N_9177,N_8513);
nand U9820 (N_9820,N_9360,N_9099);
xnor U9821 (N_9821,N_8517,N_9158);
or U9822 (N_9822,N_8575,N_9429);
and U9823 (N_9823,N_8451,N_8424);
nor U9824 (N_9824,N_8483,N_8577);
or U9825 (N_9825,N_9525,N_9006);
xnor U9826 (N_9826,N_8459,N_9173);
and U9827 (N_9827,N_9038,N_8934);
and U9828 (N_9828,N_8468,N_8782);
and U9829 (N_9829,N_8465,N_8841);
and U9830 (N_9830,N_8539,N_9047);
xnor U9831 (N_9831,N_9576,N_8750);
xor U9832 (N_9832,N_9416,N_8968);
nand U9833 (N_9833,N_8971,N_8733);
xnor U9834 (N_9834,N_8869,N_9565);
nand U9835 (N_9835,N_9226,N_9591);
nand U9836 (N_9836,N_8521,N_8582);
and U9837 (N_9837,N_8910,N_8989);
and U9838 (N_9838,N_9543,N_9372);
and U9839 (N_9839,N_8860,N_9123);
xnor U9840 (N_9840,N_9080,N_8441);
nand U9841 (N_9841,N_9208,N_9569);
nand U9842 (N_9842,N_8802,N_9288);
nand U9843 (N_9843,N_9113,N_8760);
nor U9844 (N_9844,N_9164,N_9587);
xnor U9845 (N_9845,N_8435,N_8467);
nand U9846 (N_9846,N_8470,N_9077);
or U9847 (N_9847,N_8825,N_8903);
or U9848 (N_9848,N_9414,N_9045);
or U9849 (N_9849,N_9324,N_9110);
or U9850 (N_9850,N_8637,N_8461);
or U9851 (N_9851,N_8569,N_9431);
xor U9852 (N_9852,N_8962,N_8509);
nor U9853 (N_9853,N_8871,N_8564);
nand U9854 (N_9854,N_8607,N_9029);
nand U9855 (N_9855,N_9023,N_9011);
or U9856 (N_9856,N_8615,N_9236);
and U9857 (N_9857,N_8893,N_9518);
nand U9858 (N_9858,N_9440,N_8861);
nor U9859 (N_9859,N_8678,N_8651);
nand U9860 (N_9860,N_9238,N_8652);
and U9861 (N_9861,N_9125,N_9090);
xor U9862 (N_9862,N_8846,N_9151);
xor U9863 (N_9863,N_8806,N_8506);
nor U9864 (N_9864,N_8428,N_9203);
nand U9865 (N_9865,N_8912,N_8434);
nor U9866 (N_9866,N_9473,N_8420);
and U9867 (N_9867,N_9059,N_9316);
or U9868 (N_9868,N_9083,N_8954);
and U9869 (N_9869,N_9501,N_9096);
xnor U9870 (N_9870,N_9275,N_9223);
nor U9871 (N_9871,N_8737,N_9001);
nand U9872 (N_9872,N_9134,N_8712);
xnor U9873 (N_9873,N_8629,N_9225);
nand U9874 (N_9874,N_9445,N_9124);
nand U9875 (N_9875,N_9145,N_8866);
or U9876 (N_9876,N_9536,N_9396);
or U9877 (N_9877,N_8972,N_8886);
xnor U9878 (N_9878,N_9289,N_9129);
or U9879 (N_9879,N_8474,N_9181);
nand U9880 (N_9880,N_8725,N_8943);
or U9881 (N_9881,N_8587,N_8680);
and U9882 (N_9882,N_8628,N_9184);
nand U9883 (N_9883,N_8767,N_9290);
xnor U9884 (N_9884,N_9204,N_8530);
nor U9885 (N_9885,N_9030,N_9240);
or U9886 (N_9886,N_8581,N_8614);
or U9887 (N_9887,N_9310,N_8870);
xor U9888 (N_9888,N_8508,N_9438);
nand U9889 (N_9889,N_9237,N_8718);
nand U9890 (N_9890,N_8729,N_8985);
nor U9891 (N_9891,N_8487,N_8759);
or U9892 (N_9892,N_9128,N_8758);
and U9893 (N_9893,N_9405,N_9509);
or U9894 (N_9894,N_9022,N_8793);
nand U9895 (N_9895,N_8548,N_8776);
and U9896 (N_9896,N_9404,N_8601);
nand U9897 (N_9897,N_8422,N_9234);
or U9898 (N_9898,N_8514,N_9594);
and U9899 (N_9899,N_8491,N_8895);
and U9900 (N_9900,N_8527,N_8413);
and U9901 (N_9901,N_9331,N_9574);
nor U9902 (N_9902,N_9277,N_9439);
xnor U9903 (N_9903,N_9595,N_9019);
and U9904 (N_9904,N_9381,N_9206);
nand U9905 (N_9905,N_9303,N_9332);
xnor U9906 (N_9906,N_9550,N_9068);
nor U9907 (N_9907,N_9535,N_8700);
xor U9908 (N_9908,N_9063,N_9507);
or U9909 (N_9909,N_9388,N_9563);
nor U9910 (N_9910,N_8715,N_8580);
xnor U9911 (N_9911,N_8631,N_8887);
and U9912 (N_9912,N_8634,N_8619);
or U9913 (N_9913,N_8611,N_8822);
nand U9914 (N_9914,N_9008,N_9150);
and U9915 (N_9915,N_8982,N_8765);
or U9916 (N_9916,N_8720,N_9287);
nor U9917 (N_9917,N_9178,N_8734);
or U9918 (N_9918,N_8504,N_9511);
or U9919 (N_9919,N_9326,N_9207);
and U9920 (N_9920,N_8595,N_8976);
nor U9921 (N_9921,N_8691,N_9265);
nor U9922 (N_9922,N_9020,N_9493);
nor U9923 (N_9923,N_9117,N_8951);
xnor U9924 (N_9924,N_8850,N_8937);
nand U9925 (N_9925,N_8497,N_9329);
nor U9926 (N_9926,N_9050,N_8714);
and U9927 (N_9927,N_8613,N_9500);
and U9928 (N_9928,N_9425,N_9247);
or U9929 (N_9929,N_8638,N_9423);
nand U9930 (N_9930,N_8405,N_8590);
xnor U9931 (N_9931,N_8510,N_9286);
nor U9932 (N_9932,N_9450,N_9163);
and U9933 (N_9933,N_8935,N_8562);
nor U9934 (N_9934,N_8583,N_9363);
or U9935 (N_9935,N_8791,N_9475);
or U9936 (N_9936,N_9126,N_9169);
or U9937 (N_9937,N_8645,N_8698);
nor U9938 (N_9938,N_9002,N_9084);
nand U9939 (N_9939,N_8851,N_9581);
or U9940 (N_9940,N_9482,N_9464);
or U9941 (N_9941,N_9579,N_8490);
and U9942 (N_9942,N_8987,N_8436);
xnor U9943 (N_9943,N_9213,N_8787);
nor U9944 (N_9944,N_8499,N_9457);
nor U9945 (N_9945,N_8939,N_8537);
xnor U9946 (N_9946,N_9519,N_9003);
xnor U9947 (N_9947,N_8593,N_9246);
xnor U9948 (N_9948,N_9328,N_8749);
nor U9949 (N_9949,N_9476,N_8945);
xnor U9950 (N_9950,N_9000,N_8681);
nor U9951 (N_9951,N_9190,N_9268);
and U9952 (N_9952,N_9094,N_8558);
nor U9953 (N_9953,N_8911,N_8928);
xor U9954 (N_9954,N_8803,N_8702);
or U9955 (N_9955,N_8660,N_9089);
xnor U9956 (N_9956,N_9327,N_8980);
and U9957 (N_9957,N_9427,N_9078);
nor U9958 (N_9958,N_9460,N_9487);
and U9959 (N_9959,N_9244,N_9074);
nor U9960 (N_9960,N_9504,N_8706);
and U9961 (N_9961,N_9515,N_9407);
nor U9962 (N_9962,N_8553,N_8540);
or U9963 (N_9963,N_8412,N_8632);
and U9964 (N_9964,N_9087,N_8642);
nor U9965 (N_9965,N_8567,N_8547);
and U9966 (N_9966,N_8586,N_9508);
and U9967 (N_9967,N_9233,N_9139);
nor U9968 (N_9968,N_9272,N_9227);
nor U9969 (N_9969,N_8807,N_9222);
and U9970 (N_9970,N_9424,N_9069);
xnor U9971 (N_9971,N_8443,N_8579);
nor U9972 (N_9972,N_9259,N_8410);
xnor U9973 (N_9973,N_8963,N_8966);
and U9974 (N_9974,N_8650,N_8481);
nor U9975 (N_9975,N_8798,N_8673);
or U9976 (N_9976,N_8480,N_8482);
nand U9977 (N_9977,N_9283,N_8854);
nor U9978 (N_9978,N_8462,N_9323);
and U9979 (N_9979,N_9021,N_8752);
nand U9980 (N_9980,N_9282,N_8484);
nor U9981 (N_9981,N_9558,N_8990);
xor U9982 (N_9982,N_9221,N_9531);
nand U9983 (N_9983,N_8447,N_9495);
and U9984 (N_9984,N_8774,N_9599);
nor U9985 (N_9985,N_8785,N_8830);
nand U9986 (N_9986,N_9210,N_8415);
and U9987 (N_9987,N_9091,N_8648);
nand U9988 (N_9988,N_9538,N_8795);
xnor U9989 (N_9989,N_9281,N_9195);
or U9990 (N_9990,N_9391,N_8406);
and U9991 (N_9991,N_8840,N_8666);
nand U9992 (N_9992,N_8576,N_9554);
nor U9993 (N_9993,N_9061,N_9503);
nand U9994 (N_9994,N_8815,N_9248);
and U9995 (N_9995,N_8697,N_9375);
nand U9996 (N_9996,N_9048,N_8570);
xor U9997 (N_9997,N_9235,N_8466);
nand U9998 (N_9998,N_9397,N_9010);
or U9999 (N_9999,N_8900,N_8998);
xor U10000 (N_10000,N_8568,N_9449);
and U10001 (N_10001,N_9174,N_9401);
or U10002 (N_10002,N_9410,N_9498);
nor U10003 (N_10003,N_8828,N_8526);
nand U10004 (N_10004,N_8831,N_9512);
or U10005 (N_10005,N_8625,N_9477);
nand U10006 (N_10006,N_9371,N_9342);
or U10007 (N_10007,N_9510,N_9106);
nand U10008 (N_10008,N_8554,N_8835);
xnor U10009 (N_10009,N_9426,N_9481);
or U10010 (N_10010,N_8430,N_9166);
xnor U10011 (N_10011,N_9467,N_9557);
nand U10012 (N_10012,N_8855,N_8902);
nor U10013 (N_10013,N_8908,N_8778);
or U10014 (N_10014,N_9494,N_9596);
nand U10015 (N_10015,N_8454,N_8732);
xor U10016 (N_10016,N_9313,N_9386);
xnor U10017 (N_10017,N_8457,N_9394);
nand U10018 (N_10018,N_9352,N_9544);
xor U10019 (N_10019,N_8958,N_9530);
xor U10020 (N_10020,N_8901,N_8689);
xor U10021 (N_10021,N_8409,N_9412);
xor U10022 (N_10022,N_9319,N_8994);
or U10023 (N_10023,N_8408,N_9088);
nor U10024 (N_10024,N_9393,N_9037);
nand U10025 (N_10025,N_9340,N_8606);
or U10026 (N_10026,N_9135,N_8757);
and U10027 (N_10027,N_9024,N_9437);
or U10028 (N_10028,N_8477,N_8961);
and U10029 (N_10029,N_9141,N_8674);
and U10030 (N_10030,N_9243,N_8572);
nor U10031 (N_10031,N_8772,N_9086);
and U10032 (N_10032,N_8597,N_9364);
or U10033 (N_10033,N_8885,N_8769);
or U10034 (N_10034,N_8675,N_9378);
nor U10035 (N_10035,N_9456,N_9549);
nand U10036 (N_10036,N_9093,N_9269);
nor U10037 (N_10037,N_9516,N_9079);
nand U10038 (N_10038,N_8783,N_9257);
or U10039 (N_10039,N_9212,N_8832);
or U10040 (N_10040,N_8670,N_8696);
and U10041 (N_10041,N_8488,N_9537);
or U10042 (N_10042,N_9167,N_8414);
and U10043 (N_10043,N_8884,N_9180);
xor U10044 (N_10044,N_8946,N_9347);
nand U10045 (N_10045,N_9188,N_8589);
and U10046 (N_10046,N_9492,N_8543);
xnor U10047 (N_10047,N_8404,N_9545);
xnor U10048 (N_10048,N_8957,N_8863);
nand U10049 (N_10049,N_9231,N_8427);
and U10050 (N_10050,N_8922,N_8449);
or U10051 (N_10051,N_9548,N_9202);
xnor U10052 (N_10052,N_9009,N_9463);
or U10053 (N_10053,N_8476,N_9300);
nand U10054 (N_10054,N_8872,N_9547);
and U10055 (N_10055,N_8578,N_9597);
and U10056 (N_10056,N_9379,N_9230);
nand U10057 (N_10057,N_8710,N_8602);
xor U10058 (N_10058,N_9214,N_9172);
nor U10059 (N_10059,N_9505,N_9028);
and U10060 (N_10060,N_9468,N_9217);
nor U10061 (N_10061,N_8703,N_8460);
and U10062 (N_10062,N_8827,N_9454);
or U10063 (N_10063,N_9108,N_8875);
or U10064 (N_10064,N_8557,N_9483);
nor U10065 (N_10065,N_9185,N_8671);
and U10066 (N_10066,N_8978,N_8599);
xnor U10067 (N_10067,N_8933,N_8800);
nand U10068 (N_10068,N_8605,N_8551);
or U10069 (N_10069,N_8790,N_8981);
nor U10070 (N_10070,N_9348,N_8768);
nand U10071 (N_10071,N_9435,N_9071);
xnor U10072 (N_10072,N_9153,N_8672);
xnor U10073 (N_10073,N_9215,N_8439);
or U10074 (N_10074,N_8502,N_9474);
and U10075 (N_10075,N_8524,N_9409);
nor U10076 (N_10076,N_8781,N_8814);
or U10077 (N_10077,N_9081,N_9066);
or U10078 (N_10078,N_8763,N_8464);
xnor U10079 (N_10079,N_9143,N_9199);
and U10080 (N_10080,N_9256,N_9261);
xor U10081 (N_10081,N_9312,N_8511);
and U10082 (N_10082,N_8708,N_8761);
or U10083 (N_10083,N_8522,N_9198);
nand U10084 (N_10084,N_8940,N_8984);
xnor U10085 (N_10085,N_9452,N_8463);
xnor U10086 (N_10086,N_9539,N_9007);
nor U10087 (N_10087,N_8914,N_9146);
nor U10088 (N_10088,N_9551,N_8916);
nand U10089 (N_10089,N_9148,N_8823);
and U10090 (N_10090,N_8684,N_8799);
and U10091 (N_10091,N_9572,N_9144);
nand U10092 (N_10092,N_9577,N_8423);
nand U10093 (N_10093,N_8809,N_9527);
xor U10094 (N_10094,N_9358,N_9302);
xor U10095 (N_10095,N_9252,N_8764);
xnor U10096 (N_10096,N_9098,N_9359);
or U10097 (N_10097,N_9052,N_8836);
xnor U10098 (N_10098,N_9176,N_8834);
or U10099 (N_10099,N_9042,N_8838);
nand U10100 (N_10100,N_8919,N_8833);
xnor U10101 (N_10101,N_9067,N_8518);
xnor U10102 (N_10102,N_8877,N_9192);
nand U10103 (N_10103,N_8626,N_8742);
xnor U10104 (N_10104,N_9140,N_8942);
nor U10105 (N_10105,N_8654,N_8438);
and U10106 (N_10106,N_8520,N_9470);
or U10107 (N_10107,N_9354,N_9095);
xnor U10108 (N_10108,N_8754,N_8794);
nand U10109 (N_10109,N_9279,N_9432);
xor U10110 (N_10110,N_8528,N_8453);
nor U10111 (N_10111,N_9478,N_9297);
nand U10112 (N_10112,N_9488,N_8820);
nand U10113 (N_10113,N_9034,N_9033);
xor U10114 (N_10114,N_8826,N_9497);
or U10115 (N_10115,N_8779,N_8426);
nor U10116 (N_10116,N_9127,N_9182);
nor U10117 (N_10117,N_8661,N_8693);
nor U10118 (N_10118,N_9012,N_9556);
nand U10119 (N_10119,N_8429,N_8622);
nand U10120 (N_10120,N_9434,N_8907);
nand U10121 (N_10121,N_9104,N_9224);
nor U10122 (N_10122,N_9311,N_9149);
nor U10123 (N_10123,N_8694,N_8731);
nand U10124 (N_10124,N_9447,N_9161);
nand U10125 (N_10125,N_9552,N_9183);
nand U10126 (N_10126,N_9251,N_8571);
or U10127 (N_10127,N_8536,N_8796);
nor U10128 (N_10128,N_9155,N_8458);
xor U10129 (N_10129,N_9484,N_9357);
or U10130 (N_10130,N_9380,N_9107);
xor U10131 (N_10131,N_9555,N_8494);
xnor U10132 (N_10132,N_9245,N_8560);
nor U10133 (N_10133,N_9132,N_8890);
and U10134 (N_10134,N_9250,N_9196);
and U10135 (N_10135,N_9197,N_9325);
nand U10136 (N_10136,N_8635,N_8950);
or U10137 (N_10137,N_8821,N_8455);
or U10138 (N_10138,N_9571,N_9171);
xor U10139 (N_10139,N_8529,N_8864);
and U10140 (N_10140,N_9418,N_9013);
nand U10141 (N_10141,N_9253,N_8743);
nand U10142 (N_10142,N_8471,N_9349);
or U10143 (N_10143,N_8665,N_8889);
xor U10144 (N_10144,N_9258,N_9112);
and U10145 (N_10145,N_9521,N_8545);
xor U10146 (N_10146,N_8588,N_8609);
nand U10147 (N_10147,N_8921,N_8633);
or U10148 (N_10148,N_8766,N_9072);
nor U10149 (N_10149,N_8948,N_8865);
and U10150 (N_10150,N_9421,N_8525);
nor U10151 (N_10151,N_9373,N_8541);
xnor U10152 (N_10152,N_9338,N_9260);
nand U10153 (N_10153,N_8898,N_9296);
nand U10154 (N_10154,N_9309,N_9330);
xnor U10155 (N_10155,N_9462,N_8747);
xor U10156 (N_10156,N_8478,N_8975);
nor U10157 (N_10157,N_8859,N_8923);
and U10158 (N_10158,N_9444,N_8930);
and U10159 (N_10159,N_9267,N_8555);
or U10160 (N_10160,N_8986,N_9411);
nand U10161 (N_10161,N_8699,N_8837);
nor U10162 (N_10162,N_9015,N_9442);
or U10163 (N_10163,N_8744,N_9142);
or U10164 (N_10164,N_8667,N_9353);
or U10165 (N_10165,N_9322,N_9085);
and U10166 (N_10166,N_9194,N_9249);
or U10167 (N_10167,N_9318,N_9567);
nor U10168 (N_10168,N_8717,N_9014);
nand U10169 (N_10169,N_8456,N_8618);
nor U10170 (N_10170,N_8472,N_8929);
nand U10171 (N_10171,N_9561,N_9523);
nor U10172 (N_10172,N_8883,N_8623);
xor U10173 (N_10173,N_8792,N_9216);
xor U10174 (N_10174,N_9356,N_9053);
and U10175 (N_10175,N_8881,N_8896);
or U10176 (N_10176,N_9559,N_8538);
nand U10177 (N_10177,N_9241,N_8736);
and U10178 (N_10178,N_8640,N_9480);
and U10179 (N_10179,N_9138,N_9035);
or U10180 (N_10180,N_8507,N_8542);
nand U10181 (N_10181,N_9455,N_9588);
or U10182 (N_10182,N_8780,N_9489);
nor U10183 (N_10183,N_8552,N_9109);
or U10184 (N_10184,N_9517,N_8753);
or U10185 (N_10185,N_8748,N_8646);
xor U10186 (N_10186,N_9119,N_8668);
nor U10187 (N_10187,N_8756,N_9298);
nor U10188 (N_10188,N_9046,N_9472);
or U10189 (N_10189,N_8591,N_8690);
and U10190 (N_10190,N_9339,N_9465);
or U10191 (N_10191,N_9430,N_8847);
and U10192 (N_10192,N_9294,N_9115);
nand U10193 (N_10193,N_8603,N_8421);
nand U10194 (N_10194,N_8960,N_9568);
xor U10195 (N_10195,N_9101,N_9399);
xor U10196 (N_10196,N_9004,N_8446);
xnor U10197 (N_10197,N_9273,N_9395);
nand U10198 (N_10198,N_8656,N_9291);
xnor U10199 (N_10199,N_8662,N_9292);
nor U10200 (N_10200,N_8850,N_8566);
nor U10201 (N_10201,N_8899,N_9245);
or U10202 (N_10202,N_9524,N_9534);
nor U10203 (N_10203,N_9012,N_9355);
or U10204 (N_10204,N_9004,N_9007);
xnor U10205 (N_10205,N_9229,N_8608);
and U10206 (N_10206,N_9312,N_8870);
nand U10207 (N_10207,N_9385,N_9517);
or U10208 (N_10208,N_8764,N_8620);
nand U10209 (N_10209,N_8966,N_9022);
nand U10210 (N_10210,N_9196,N_9575);
nor U10211 (N_10211,N_9523,N_8972);
nor U10212 (N_10212,N_9248,N_8896);
or U10213 (N_10213,N_8856,N_9145);
xnor U10214 (N_10214,N_8575,N_9573);
or U10215 (N_10215,N_9578,N_8663);
or U10216 (N_10216,N_8870,N_9388);
or U10217 (N_10217,N_9580,N_9040);
nand U10218 (N_10218,N_9112,N_9140);
or U10219 (N_10219,N_9329,N_8919);
nor U10220 (N_10220,N_9427,N_9310);
xor U10221 (N_10221,N_9390,N_9435);
nand U10222 (N_10222,N_9170,N_9283);
and U10223 (N_10223,N_9171,N_8711);
nor U10224 (N_10224,N_8960,N_8646);
and U10225 (N_10225,N_8479,N_8624);
or U10226 (N_10226,N_8439,N_8540);
xor U10227 (N_10227,N_9300,N_8775);
or U10228 (N_10228,N_9079,N_8402);
or U10229 (N_10229,N_8686,N_9395);
or U10230 (N_10230,N_9082,N_9106);
or U10231 (N_10231,N_8923,N_8690);
or U10232 (N_10232,N_9393,N_8888);
or U10233 (N_10233,N_9075,N_8615);
or U10234 (N_10234,N_9412,N_9251);
or U10235 (N_10235,N_9075,N_9132);
nor U10236 (N_10236,N_9007,N_8545);
xnor U10237 (N_10237,N_8721,N_8473);
nand U10238 (N_10238,N_8918,N_8634);
nor U10239 (N_10239,N_9289,N_9273);
and U10240 (N_10240,N_8545,N_9497);
nand U10241 (N_10241,N_8422,N_8830);
or U10242 (N_10242,N_9534,N_8916);
nand U10243 (N_10243,N_8850,N_8545);
and U10244 (N_10244,N_9036,N_8876);
nor U10245 (N_10245,N_9172,N_9410);
nor U10246 (N_10246,N_9211,N_8758);
or U10247 (N_10247,N_9564,N_9501);
and U10248 (N_10248,N_9359,N_8602);
nor U10249 (N_10249,N_9211,N_8828);
and U10250 (N_10250,N_9044,N_9487);
and U10251 (N_10251,N_8700,N_9379);
xor U10252 (N_10252,N_9247,N_8864);
and U10253 (N_10253,N_9524,N_8960);
xor U10254 (N_10254,N_9205,N_9058);
nor U10255 (N_10255,N_9441,N_8889);
or U10256 (N_10256,N_8571,N_8812);
xor U10257 (N_10257,N_8472,N_8941);
nand U10258 (N_10258,N_8985,N_9476);
nand U10259 (N_10259,N_8750,N_9396);
and U10260 (N_10260,N_9268,N_9228);
xor U10261 (N_10261,N_9264,N_9207);
nor U10262 (N_10262,N_8741,N_8545);
or U10263 (N_10263,N_8477,N_9112);
xor U10264 (N_10264,N_9149,N_9476);
or U10265 (N_10265,N_8500,N_8694);
nor U10266 (N_10266,N_8655,N_9027);
nor U10267 (N_10267,N_9502,N_8830);
xor U10268 (N_10268,N_9258,N_8716);
nor U10269 (N_10269,N_8755,N_8486);
and U10270 (N_10270,N_8418,N_9506);
and U10271 (N_10271,N_9357,N_8845);
or U10272 (N_10272,N_9512,N_9367);
and U10273 (N_10273,N_9095,N_9133);
nand U10274 (N_10274,N_8846,N_9227);
or U10275 (N_10275,N_8559,N_9047);
and U10276 (N_10276,N_8836,N_9376);
xnor U10277 (N_10277,N_9445,N_8790);
nor U10278 (N_10278,N_8826,N_9471);
xnor U10279 (N_10279,N_8487,N_9112);
nor U10280 (N_10280,N_9170,N_9164);
nor U10281 (N_10281,N_8712,N_9074);
or U10282 (N_10282,N_9550,N_8886);
xor U10283 (N_10283,N_9210,N_8722);
and U10284 (N_10284,N_8775,N_9256);
xnor U10285 (N_10285,N_9352,N_8773);
and U10286 (N_10286,N_9407,N_8602);
xor U10287 (N_10287,N_8404,N_9396);
or U10288 (N_10288,N_9195,N_9044);
and U10289 (N_10289,N_9274,N_8607);
xor U10290 (N_10290,N_8763,N_9513);
nand U10291 (N_10291,N_9279,N_9191);
nor U10292 (N_10292,N_9375,N_9402);
or U10293 (N_10293,N_9007,N_8821);
or U10294 (N_10294,N_8494,N_9294);
nor U10295 (N_10295,N_8595,N_9129);
nor U10296 (N_10296,N_8570,N_9213);
nand U10297 (N_10297,N_8504,N_9118);
nor U10298 (N_10298,N_8818,N_8563);
nand U10299 (N_10299,N_9398,N_9307);
or U10300 (N_10300,N_8746,N_8571);
xnor U10301 (N_10301,N_8758,N_8600);
and U10302 (N_10302,N_9290,N_8466);
nor U10303 (N_10303,N_8969,N_8988);
or U10304 (N_10304,N_8706,N_9193);
nor U10305 (N_10305,N_9266,N_9573);
nor U10306 (N_10306,N_9382,N_9361);
and U10307 (N_10307,N_9069,N_8636);
or U10308 (N_10308,N_9298,N_8564);
xor U10309 (N_10309,N_8790,N_9084);
or U10310 (N_10310,N_9462,N_9222);
and U10311 (N_10311,N_8810,N_8811);
nor U10312 (N_10312,N_9286,N_8656);
xor U10313 (N_10313,N_8460,N_9302);
or U10314 (N_10314,N_9557,N_9472);
nand U10315 (N_10315,N_8869,N_8645);
xor U10316 (N_10316,N_8881,N_9509);
nor U10317 (N_10317,N_9415,N_9438);
or U10318 (N_10318,N_9064,N_8651);
and U10319 (N_10319,N_8902,N_8541);
xnor U10320 (N_10320,N_8488,N_8684);
xor U10321 (N_10321,N_9234,N_9326);
and U10322 (N_10322,N_9449,N_8730);
nand U10323 (N_10323,N_9043,N_9560);
nand U10324 (N_10324,N_9184,N_9286);
and U10325 (N_10325,N_9354,N_9478);
nor U10326 (N_10326,N_9505,N_8602);
xor U10327 (N_10327,N_8631,N_8409);
nand U10328 (N_10328,N_9439,N_9151);
nand U10329 (N_10329,N_9116,N_8899);
nand U10330 (N_10330,N_8651,N_9560);
xnor U10331 (N_10331,N_8626,N_9441);
nand U10332 (N_10332,N_8634,N_8968);
or U10333 (N_10333,N_9528,N_9036);
nand U10334 (N_10334,N_9134,N_8998);
and U10335 (N_10335,N_9592,N_8731);
xnor U10336 (N_10336,N_8573,N_8781);
nand U10337 (N_10337,N_8410,N_9177);
nor U10338 (N_10338,N_8869,N_8842);
xnor U10339 (N_10339,N_9232,N_9525);
nor U10340 (N_10340,N_8824,N_9030);
nand U10341 (N_10341,N_8472,N_9015);
xor U10342 (N_10342,N_9083,N_8609);
xor U10343 (N_10343,N_9400,N_9543);
nand U10344 (N_10344,N_8793,N_8637);
xor U10345 (N_10345,N_9505,N_9421);
or U10346 (N_10346,N_9577,N_9003);
xnor U10347 (N_10347,N_8998,N_8583);
nand U10348 (N_10348,N_8859,N_8787);
and U10349 (N_10349,N_8916,N_9554);
nor U10350 (N_10350,N_9008,N_9212);
nand U10351 (N_10351,N_8964,N_9268);
or U10352 (N_10352,N_8926,N_8765);
nand U10353 (N_10353,N_8926,N_8402);
nor U10354 (N_10354,N_9471,N_9392);
and U10355 (N_10355,N_9230,N_9304);
or U10356 (N_10356,N_8556,N_9245);
nor U10357 (N_10357,N_9000,N_8475);
and U10358 (N_10358,N_8918,N_9494);
nand U10359 (N_10359,N_8513,N_9350);
or U10360 (N_10360,N_8560,N_8778);
nand U10361 (N_10361,N_8555,N_8661);
and U10362 (N_10362,N_9442,N_8995);
and U10363 (N_10363,N_8522,N_8566);
or U10364 (N_10364,N_8767,N_9405);
xor U10365 (N_10365,N_8505,N_8612);
and U10366 (N_10366,N_9318,N_8722);
or U10367 (N_10367,N_9269,N_9428);
or U10368 (N_10368,N_8755,N_9534);
nand U10369 (N_10369,N_9356,N_8516);
nand U10370 (N_10370,N_9011,N_9266);
nand U10371 (N_10371,N_9096,N_9288);
or U10372 (N_10372,N_8537,N_9145);
nand U10373 (N_10373,N_9323,N_8495);
nor U10374 (N_10374,N_8912,N_8432);
nand U10375 (N_10375,N_9210,N_8526);
or U10376 (N_10376,N_8836,N_9481);
and U10377 (N_10377,N_8800,N_9356);
nor U10378 (N_10378,N_9452,N_8953);
nand U10379 (N_10379,N_8690,N_9139);
nor U10380 (N_10380,N_8666,N_8783);
or U10381 (N_10381,N_8625,N_9002);
nand U10382 (N_10382,N_9461,N_8623);
nor U10383 (N_10383,N_9255,N_8605);
nor U10384 (N_10384,N_8693,N_8778);
nor U10385 (N_10385,N_9175,N_9528);
or U10386 (N_10386,N_8753,N_9100);
nand U10387 (N_10387,N_9215,N_9012);
nor U10388 (N_10388,N_9009,N_8759);
and U10389 (N_10389,N_9322,N_9357);
xor U10390 (N_10390,N_9515,N_9008);
nand U10391 (N_10391,N_8549,N_9082);
nor U10392 (N_10392,N_9547,N_9521);
xor U10393 (N_10393,N_8642,N_9058);
nand U10394 (N_10394,N_8864,N_8534);
or U10395 (N_10395,N_9374,N_9397);
and U10396 (N_10396,N_9304,N_8824);
or U10397 (N_10397,N_8482,N_8670);
and U10398 (N_10398,N_8495,N_8479);
or U10399 (N_10399,N_8897,N_9370);
xor U10400 (N_10400,N_9358,N_8559);
nand U10401 (N_10401,N_9094,N_9023);
xnor U10402 (N_10402,N_8473,N_9032);
nor U10403 (N_10403,N_8882,N_8427);
or U10404 (N_10404,N_8418,N_9206);
and U10405 (N_10405,N_8732,N_8846);
nand U10406 (N_10406,N_8840,N_9223);
nand U10407 (N_10407,N_9333,N_9471);
and U10408 (N_10408,N_8768,N_9417);
xor U10409 (N_10409,N_9501,N_8641);
nor U10410 (N_10410,N_8826,N_9098);
nand U10411 (N_10411,N_8609,N_8430);
nor U10412 (N_10412,N_9364,N_8770);
or U10413 (N_10413,N_8599,N_8585);
or U10414 (N_10414,N_9475,N_8479);
or U10415 (N_10415,N_8561,N_8788);
or U10416 (N_10416,N_8526,N_9438);
nand U10417 (N_10417,N_8887,N_8673);
nor U10418 (N_10418,N_8728,N_9187);
or U10419 (N_10419,N_9262,N_8785);
or U10420 (N_10420,N_8940,N_9544);
nor U10421 (N_10421,N_8865,N_9291);
and U10422 (N_10422,N_9399,N_9492);
nor U10423 (N_10423,N_8760,N_9553);
and U10424 (N_10424,N_8507,N_9254);
nand U10425 (N_10425,N_8887,N_9122);
xnor U10426 (N_10426,N_8947,N_8765);
and U10427 (N_10427,N_9145,N_8405);
nor U10428 (N_10428,N_9591,N_9542);
xor U10429 (N_10429,N_8734,N_8826);
xnor U10430 (N_10430,N_9597,N_8442);
xnor U10431 (N_10431,N_8691,N_9020);
and U10432 (N_10432,N_8774,N_9195);
and U10433 (N_10433,N_8796,N_8730);
nand U10434 (N_10434,N_9013,N_8550);
xnor U10435 (N_10435,N_9318,N_9580);
xor U10436 (N_10436,N_8513,N_8944);
nor U10437 (N_10437,N_9339,N_8997);
nand U10438 (N_10438,N_8666,N_9346);
or U10439 (N_10439,N_8785,N_9010);
xnor U10440 (N_10440,N_8600,N_9465);
and U10441 (N_10441,N_8694,N_8779);
nor U10442 (N_10442,N_9583,N_9214);
and U10443 (N_10443,N_9285,N_8423);
nor U10444 (N_10444,N_8963,N_9493);
xor U10445 (N_10445,N_9508,N_8856);
and U10446 (N_10446,N_8422,N_9408);
xnor U10447 (N_10447,N_9365,N_9335);
nor U10448 (N_10448,N_8940,N_8945);
nand U10449 (N_10449,N_9393,N_8995);
nand U10450 (N_10450,N_8492,N_9203);
nand U10451 (N_10451,N_9071,N_8935);
or U10452 (N_10452,N_8617,N_8963);
nor U10453 (N_10453,N_8738,N_8423);
nor U10454 (N_10454,N_9442,N_8497);
and U10455 (N_10455,N_8811,N_9424);
nor U10456 (N_10456,N_8533,N_9503);
nor U10457 (N_10457,N_9562,N_9142);
and U10458 (N_10458,N_9268,N_9507);
nor U10459 (N_10459,N_9323,N_9447);
and U10460 (N_10460,N_9525,N_9152);
and U10461 (N_10461,N_8685,N_8699);
nor U10462 (N_10462,N_9201,N_9309);
and U10463 (N_10463,N_8822,N_8598);
nor U10464 (N_10464,N_8668,N_8915);
xnor U10465 (N_10465,N_9331,N_8593);
nor U10466 (N_10466,N_9383,N_9576);
xor U10467 (N_10467,N_8947,N_8454);
or U10468 (N_10468,N_8433,N_9237);
xor U10469 (N_10469,N_9542,N_9105);
xnor U10470 (N_10470,N_9335,N_9517);
xnor U10471 (N_10471,N_8489,N_9191);
or U10472 (N_10472,N_9536,N_8710);
nand U10473 (N_10473,N_9554,N_9481);
and U10474 (N_10474,N_8962,N_9342);
and U10475 (N_10475,N_9235,N_9079);
nor U10476 (N_10476,N_8425,N_9267);
or U10477 (N_10477,N_9174,N_8854);
nand U10478 (N_10478,N_8515,N_9115);
and U10479 (N_10479,N_9535,N_8778);
nor U10480 (N_10480,N_8501,N_8504);
or U10481 (N_10481,N_9360,N_8716);
nand U10482 (N_10482,N_8443,N_8756);
and U10483 (N_10483,N_8432,N_9226);
and U10484 (N_10484,N_8870,N_9470);
and U10485 (N_10485,N_8570,N_9067);
nand U10486 (N_10486,N_9052,N_9208);
nand U10487 (N_10487,N_9516,N_9205);
and U10488 (N_10488,N_8681,N_9467);
nand U10489 (N_10489,N_9142,N_9267);
or U10490 (N_10490,N_8826,N_8510);
nor U10491 (N_10491,N_9567,N_9290);
and U10492 (N_10492,N_8412,N_9388);
xnor U10493 (N_10493,N_9565,N_9513);
or U10494 (N_10494,N_9102,N_9399);
xnor U10495 (N_10495,N_8904,N_8569);
and U10496 (N_10496,N_9288,N_8738);
or U10497 (N_10497,N_9467,N_9128);
and U10498 (N_10498,N_8921,N_9513);
nand U10499 (N_10499,N_9319,N_9252);
and U10500 (N_10500,N_9176,N_8979);
xor U10501 (N_10501,N_9390,N_8798);
or U10502 (N_10502,N_8507,N_8991);
nor U10503 (N_10503,N_9108,N_9552);
nand U10504 (N_10504,N_8455,N_9290);
nor U10505 (N_10505,N_8685,N_9036);
xnor U10506 (N_10506,N_8765,N_8404);
and U10507 (N_10507,N_9521,N_8936);
nor U10508 (N_10508,N_9127,N_9273);
xor U10509 (N_10509,N_8731,N_9380);
xnor U10510 (N_10510,N_8815,N_8508);
xor U10511 (N_10511,N_8969,N_9560);
and U10512 (N_10512,N_9382,N_9343);
nor U10513 (N_10513,N_9034,N_9114);
and U10514 (N_10514,N_9195,N_9088);
or U10515 (N_10515,N_8517,N_8773);
and U10516 (N_10516,N_9597,N_9563);
or U10517 (N_10517,N_8601,N_8771);
nor U10518 (N_10518,N_9374,N_9168);
xor U10519 (N_10519,N_8850,N_9124);
or U10520 (N_10520,N_8674,N_9562);
nor U10521 (N_10521,N_9320,N_8626);
xnor U10522 (N_10522,N_8478,N_8607);
or U10523 (N_10523,N_8457,N_8509);
nand U10524 (N_10524,N_9591,N_9279);
and U10525 (N_10525,N_8727,N_8882);
nor U10526 (N_10526,N_8628,N_9424);
nand U10527 (N_10527,N_9219,N_8543);
nand U10528 (N_10528,N_9400,N_8840);
nor U10529 (N_10529,N_8621,N_8866);
xnor U10530 (N_10530,N_8787,N_9482);
nor U10531 (N_10531,N_8837,N_9534);
or U10532 (N_10532,N_8870,N_8850);
or U10533 (N_10533,N_9119,N_9554);
nor U10534 (N_10534,N_8893,N_9312);
xnor U10535 (N_10535,N_8713,N_9326);
nand U10536 (N_10536,N_9565,N_8633);
and U10537 (N_10537,N_8418,N_9463);
and U10538 (N_10538,N_9095,N_9212);
nor U10539 (N_10539,N_9005,N_9546);
or U10540 (N_10540,N_9486,N_8731);
and U10541 (N_10541,N_8773,N_9152);
nor U10542 (N_10542,N_9373,N_8782);
nand U10543 (N_10543,N_8445,N_8997);
nor U10544 (N_10544,N_8740,N_8538);
or U10545 (N_10545,N_9157,N_9115);
nand U10546 (N_10546,N_9019,N_9259);
nor U10547 (N_10547,N_9554,N_8468);
nand U10548 (N_10548,N_8688,N_8963);
and U10549 (N_10549,N_8674,N_8405);
and U10550 (N_10550,N_8533,N_8978);
or U10551 (N_10551,N_9257,N_9503);
nand U10552 (N_10552,N_9209,N_9205);
nor U10553 (N_10553,N_9516,N_9012);
xor U10554 (N_10554,N_8485,N_8940);
nor U10555 (N_10555,N_8878,N_8779);
or U10556 (N_10556,N_8548,N_8513);
nand U10557 (N_10557,N_8633,N_9167);
xnor U10558 (N_10558,N_8428,N_8592);
xor U10559 (N_10559,N_9315,N_8650);
or U10560 (N_10560,N_9258,N_8734);
or U10561 (N_10561,N_9482,N_9038);
nand U10562 (N_10562,N_9022,N_8747);
or U10563 (N_10563,N_9006,N_9425);
or U10564 (N_10564,N_9333,N_8739);
nor U10565 (N_10565,N_8969,N_9304);
nor U10566 (N_10566,N_8491,N_9122);
nor U10567 (N_10567,N_8877,N_8816);
and U10568 (N_10568,N_8701,N_8965);
nor U10569 (N_10569,N_9236,N_8709);
or U10570 (N_10570,N_8626,N_9008);
nand U10571 (N_10571,N_8758,N_8624);
xor U10572 (N_10572,N_9174,N_9572);
nand U10573 (N_10573,N_8991,N_8981);
nand U10574 (N_10574,N_8620,N_8512);
or U10575 (N_10575,N_8528,N_9161);
or U10576 (N_10576,N_9575,N_9324);
nand U10577 (N_10577,N_8725,N_9040);
nor U10578 (N_10578,N_8872,N_9114);
or U10579 (N_10579,N_9275,N_8457);
and U10580 (N_10580,N_8730,N_8885);
or U10581 (N_10581,N_8616,N_9575);
and U10582 (N_10582,N_9154,N_8964);
xor U10583 (N_10583,N_8689,N_9204);
and U10584 (N_10584,N_9061,N_8923);
and U10585 (N_10585,N_9458,N_8843);
nand U10586 (N_10586,N_8973,N_9079);
nor U10587 (N_10587,N_9295,N_9053);
and U10588 (N_10588,N_8548,N_9053);
or U10589 (N_10589,N_8767,N_8493);
nor U10590 (N_10590,N_8717,N_8745);
or U10591 (N_10591,N_9265,N_8629);
or U10592 (N_10592,N_8514,N_9001);
or U10593 (N_10593,N_9038,N_8744);
or U10594 (N_10594,N_9201,N_8783);
and U10595 (N_10595,N_9163,N_8615);
and U10596 (N_10596,N_9391,N_8711);
nand U10597 (N_10597,N_9075,N_9045);
xor U10598 (N_10598,N_9017,N_9544);
and U10599 (N_10599,N_9210,N_9193);
nand U10600 (N_10600,N_9154,N_9181);
or U10601 (N_10601,N_9426,N_8935);
nor U10602 (N_10602,N_9506,N_8422);
or U10603 (N_10603,N_8654,N_9059);
and U10604 (N_10604,N_9599,N_9256);
xor U10605 (N_10605,N_9137,N_9122);
and U10606 (N_10606,N_8483,N_9204);
nor U10607 (N_10607,N_8545,N_9176);
or U10608 (N_10608,N_9425,N_9451);
nor U10609 (N_10609,N_8881,N_8777);
and U10610 (N_10610,N_8858,N_9291);
nor U10611 (N_10611,N_8839,N_9050);
nand U10612 (N_10612,N_8459,N_8751);
and U10613 (N_10613,N_8682,N_8877);
and U10614 (N_10614,N_9008,N_8904);
nor U10615 (N_10615,N_8680,N_9024);
xnor U10616 (N_10616,N_8967,N_9047);
nor U10617 (N_10617,N_9416,N_8623);
xor U10618 (N_10618,N_8916,N_8509);
or U10619 (N_10619,N_8708,N_9103);
nand U10620 (N_10620,N_9039,N_8958);
nand U10621 (N_10621,N_9559,N_9233);
and U10622 (N_10622,N_9250,N_8445);
nand U10623 (N_10623,N_9170,N_9158);
and U10624 (N_10624,N_9567,N_9114);
or U10625 (N_10625,N_8815,N_8931);
or U10626 (N_10626,N_8533,N_8951);
or U10627 (N_10627,N_8553,N_9185);
xnor U10628 (N_10628,N_9023,N_8500);
xnor U10629 (N_10629,N_8902,N_8735);
nor U10630 (N_10630,N_9317,N_8829);
and U10631 (N_10631,N_9310,N_8995);
nor U10632 (N_10632,N_8738,N_8982);
or U10633 (N_10633,N_9270,N_9251);
and U10634 (N_10634,N_8604,N_8432);
and U10635 (N_10635,N_8640,N_8493);
xnor U10636 (N_10636,N_9125,N_9229);
nor U10637 (N_10637,N_9499,N_8988);
or U10638 (N_10638,N_9461,N_9430);
xor U10639 (N_10639,N_8523,N_8951);
nand U10640 (N_10640,N_8848,N_8699);
and U10641 (N_10641,N_9541,N_9557);
and U10642 (N_10642,N_8513,N_8659);
and U10643 (N_10643,N_9069,N_9465);
nand U10644 (N_10644,N_8462,N_8577);
xnor U10645 (N_10645,N_8730,N_9387);
nand U10646 (N_10646,N_9241,N_8964);
nor U10647 (N_10647,N_8871,N_9480);
and U10648 (N_10648,N_8553,N_8671);
nand U10649 (N_10649,N_8991,N_9256);
xnor U10650 (N_10650,N_9335,N_8824);
or U10651 (N_10651,N_8404,N_8945);
or U10652 (N_10652,N_8688,N_8785);
or U10653 (N_10653,N_8636,N_8817);
or U10654 (N_10654,N_9384,N_8663);
or U10655 (N_10655,N_9163,N_8500);
nand U10656 (N_10656,N_8599,N_8478);
nor U10657 (N_10657,N_9509,N_8679);
and U10658 (N_10658,N_8469,N_9262);
and U10659 (N_10659,N_8745,N_8559);
xnor U10660 (N_10660,N_9387,N_8503);
nand U10661 (N_10661,N_8814,N_9449);
or U10662 (N_10662,N_8437,N_9503);
xor U10663 (N_10663,N_8775,N_8917);
xnor U10664 (N_10664,N_9156,N_9491);
nor U10665 (N_10665,N_8636,N_8923);
nor U10666 (N_10666,N_8765,N_9313);
or U10667 (N_10667,N_9032,N_8799);
xor U10668 (N_10668,N_9342,N_9406);
nand U10669 (N_10669,N_8830,N_9352);
nand U10670 (N_10670,N_8874,N_9563);
nor U10671 (N_10671,N_9046,N_8797);
or U10672 (N_10672,N_8567,N_8543);
and U10673 (N_10673,N_9354,N_8404);
or U10674 (N_10674,N_8931,N_8507);
nor U10675 (N_10675,N_8779,N_9045);
or U10676 (N_10676,N_9051,N_8534);
or U10677 (N_10677,N_8469,N_8933);
and U10678 (N_10678,N_8469,N_9546);
and U10679 (N_10679,N_9055,N_8704);
nand U10680 (N_10680,N_9483,N_9019);
nor U10681 (N_10681,N_9428,N_9251);
nand U10682 (N_10682,N_9014,N_9349);
nand U10683 (N_10683,N_8491,N_9567);
and U10684 (N_10684,N_9234,N_8603);
and U10685 (N_10685,N_8455,N_9260);
nand U10686 (N_10686,N_8416,N_8791);
nand U10687 (N_10687,N_8780,N_9440);
or U10688 (N_10688,N_9051,N_8788);
and U10689 (N_10689,N_8766,N_8998);
nor U10690 (N_10690,N_8751,N_9559);
or U10691 (N_10691,N_8938,N_8459);
nand U10692 (N_10692,N_9587,N_9363);
and U10693 (N_10693,N_9337,N_9550);
xor U10694 (N_10694,N_8764,N_8507);
nor U10695 (N_10695,N_8825,N_8848);
or U10696 (N_10696,N_9000,N_9560);
xnor U10697 (N_10697,N_9422,N_9225);
or U10698 (N_10698,N_8741,N_8412);
nor U10699 (N_10699,N_8516,N_9005);
or U10700 (N_10700,N_9558,N_8976);
and U10701 (N_10701,N_8479,N_9064);
xor U10702 (N_10702,N_9285,N_9222);
and U10703 (N_10703,N_9442,N_8455);
nor U10704 (N_10704,N_8672,N_8930);
nor U10705 (N_10705,N_8617,N_8495);
and U10706 (N_10706,N_8817,N_8656);
nand U10707 (N_10707,N_8476,N_9408);
xnor U10708 (N_10708,N_9342,N_8822);
nand U10709 (N_10709,N_9176,N_9533);
xor U10710 (N_10710,N_8752,N_8558);
and U10711 (N_10711,N_8524,N_9513);
or U10712 (N_10712,N_9323,N_8685);
nand U10713 (N_10713,N_8993,N_9591);
nor U10714 (N_10714,N_8874,N_8898);
nand U10715 (N_10715,N_8990,N_8890);
xnor U10716 (N_10716,N_9349,N_9000);
and U10717 (N_10717,N_8509,N_9378);
xor U10718 (N_10718,N_9513,N_9358);
and U10719 (N_10719,N_8516,N_9552);
nor U10720 (N_10720,N_8647,N_9481);
nor U10721 (N_10721,N_8489,N_9035);
xnor U10722 (N_10722,N_8958,N_8617);
nand U10723 (N_10723,N_9446,N_9270);
xnor U10724 (N_10724,N_8791,N_9507);
and U10725 (N_10725,N_8432,N_8507);
xor U10726 (N_10726,N_8825,N_9390);
and U10727 (N_10727,N_8705,N_9289);
nor U10728 (N_10728,N_9525,N_8751);
and U10729 (N_10729,N_9287,N_9084);
xnor U10730 (N_10730,N_9315,N_8845);
xor U10731 (N_10731,N_9415,N_8491);
nand U10732 (N_10732,N_8476,N_8792);
xnor U10733 (N_10733,N_8852,N_9290);
nand U10734 (N_10734,N_8754,N_9491);
nand U10735 (N_10735,N_9043,N_9511);
nand U10736 (N_10736,N_8534,N_8464);
or U10737 (N_10737,N_8944,N_8622);
nor U10738 (N_10738,N_8775,N_8975);
nand U10739 (N_10739,N_8620,N_9092);
or U10740 (N_10740,N_8958,N_9295);
xor U10741 (N_10741,N_8411,N_8555);
xor U10742 (N_10742,N_8412,N_8814);
xor U10743 (N_10743,N_8764,N_9201);
or U10744 (N_10744,N_8815,N_8576);
xor U10745 (N_10745,N_9247,N_9106);
nor U10746 (N_10746,N_8811,N_8868);
xor U10747 (N_10747,N_8933,N_8483);
nand U10748 (N_10748,N_8843,N_9198);
nor U10749 (N_10749,N_9063,N_9103);
nor U10750 (N_10750,N_8996,N_9193);
nor U10751 (N_10751,N_8970,N_8552);
xor U10752 (N_10752,N_9023,N_9171);
and U10753 (N_10753,N_9069,N_9404);
xnor U10754 (N_10754,N_8557,N_8611);
nand U10755 (N_10755,N_9382,N_8562);
nand U10756 (N_10756,N_9554,N_8565);
or U10757 (N_10757,N_9419,N_9064);
nor U10758 (N_10758,N_9284,N_8933);
and U10759 (N_10759,N_9545,N_8491);
xor U10760 (N_10760,N_8696,N_9236);
or U10761 (N_10761,N_9524,N_9269);
nand U10762 (N_10762,N_8550,N_9016);
nand U10763 (N_10763,N_8899,N_9599);
nor U10764 (N_10764,N_9094,N_8595);
nand U10765 (N_10765,N_8893,N_8459);
or U10766 (N_10766,N_9302,N_9225);
and U10767 (N_10767,N_8936,N_8885);
xnor U10768 (N_10768,N_9296,N_9187);
nand U10769 (N_10769,N_8859,N_8948);
nor U10770 (N_10770,N_8907,N_9382);
and U10771 (N_10771,N_8664,N_8760);
nor U10772 (N_10772,N_8857,N_9321);
and U10773 (N_10773,N_8934,N_8520);
or U10774 (N_10774,N_8454,N_9155);
nand U10775 (N_10775,N_9432,N_9399);
xnor U10776 (N_10776,N_9048,N_8519);
and U10777 (N_10777,N_9283,N_9386);
and U10778 (N_10778,N_9110,N_8647);
nor U10779 (N_10779,N_8704,N_8926);
nor U10780 (N_10780,N_8506,N_9457);
or U10781 (N_10781,N_8419,N_8895);
and U10782 (N_10782,N_9577,N_9118);
and U10783 (N_10783,N_8826,N_9424);
or U10784 (N_10784,N_9565,N_9473);
nor U10785 (N_10785,N_9399,N_8834);
xnor U10786 (N_10786,N_9536,N_8627);
nand U10787 (N_10787,N_8520,N_8533);
xnor U10788 (N_10788,N_8702,N_8841);
nand U10789 (N_10789,N_8806,N_9303);
nor U10790 (N_10790,N_8550,N_8440);
xnor U10791 (N_10791,N_8948,N_8755);
nand U10792 (N_10792,N_9406,N_9144);
nor U10793 (N_10793,N_9022,N_8464);
nor U10794 (N_10794,N_8555,N_8982);
or U10795 (N_10795,N_8413,N_8647);
nor U10796 (N_10796,N_8638,N_8935);
xor U10797 (N_10797,N_8459,N_9036);
xor U10798 (N_10798,N_8887,N_9238);
nor U10799 (N_10799,N_8802,N_9530);
or U10800 (N_10800,N_10499,N_9764);
and U10801 (N_10801,N_9690,N_10589);
nand U10802 (N_10802,N_10562,N_10400);
and U10803 (N_10803,N_10471,N_10437);
xor U10804 (N_10804,N_9730,N_9788);
xor U10805 (N_10805,N_10726,N_10584);
nor U10806 (N_10806,N_9945,N_10038);
and U10807 (N_10807,N_9892,N_9819);
and U10808 (N_10808,N_10501,N_10211);
xor U10809 (N_10809,N_10745,N_10637);
or U10810 (N_10810,N_9702,N_10183);
nand U10811 (N_10811,N_10754,N_10326);
xor U10812 (N_10812,N_10480,N_10643);
or U10813 (N_10813,N_10425,N_9697);
and U10814 (N_10814,N_10032,N_9634);
nand U10815 (N_10815,N_10603,N_10468);
nand U10816 (N_10816,N_9709,N_9740);
and U10817 (N_10817,N_10178,N_10129);
nor U10818 (N_10818,N_10460,N_10284);
or U10819 (N_10819,N_9925,N_9761);
and U10820 (N_10820,N_9677,N_10138);
or U10821 (N_10821,N_10370,N_10403);
nor U10822 (N_10822,N_10737,N_10540);
nor U10823 (N_10823,N_9996,N_10538);
nor U10824 (N_10824,N_10219,N_10520);
nand U10825 (N_10825,N_9782,N_9906);
xor U10826 (N_10826,N_10601,N_9679);
nor U10827 (N_10827,N_9937,N_10537);
and U10828 (N_10828,N_9686,N_10733);
or U10829 (N_10829,N_10710,N_10573);
nor U10830 (N_10830,N_10215,N_10026);
and U10831 (N_10831,N_10788,N_9851);
and U10832 (N_10832,N_10122,N_10134);
or U10833 (N_10833,N_10655,N_10670);
and U10834 (N_10834,N_10702,N_9913);
or U10835 (N_10835,N_10181,N_10196);
or U10836 (N_10836,N_10099,N_9883);
or U10837 (N_10837,N_9845,N_9932);
and U10838 (N_10838,N_9768,N_9672);
xor U10839 (N_10839,N_10366,N_10482);
or U10840 (N_10840,N_10447,N_10436);
and U10841 (N_10841,N_10635,N_10160);
and U10842 (N_10842,N_10309,N_10678);
or U10843 (N_10843,N_10582,N_10241);
nand U10844 (N_10844,N_10360,N_10287);
and U10845 (N_10845,N_9715,N_10680);
or U10846 (N_10846,N_10536,N_9678);
nor U10847 (N_10847,N_10387,N_10775);
and U10848 (N_10848,N_10378,N_10469);
xnor U10849 (N_10849,N_10364,N_10263);
or U10850 (N_10850,N_10531,N_9614);
or U10851 (N_10851,N_9814,N_10327);
xor U10852 (N_10852,N_10549,N_9747);
nor U10853 (N_10853,N_10722,N_10596);
nor U10854 (N_10854,N_10345,N_9793);
xor U10855 (N_10855,N_10747,N_10020);
or U10856 (N_10856,N_10590,N_10444);
or U10857 (N_10857,N_9760,N_10258);
or U10858 (N_10858,N_10421,N_10310);
xnor U10859 (N_10859,N_9626,N_10422);
xnor U10860 (N_10860,N_10721,N_9775);
nand U10861 (N_10861,N_10641,N_10332);
and U10862 (N_10862,N_9710,N_10318);
and U10863 (N_10863,N_10336,N_10632);
and U10864 (N_10864,N_10485,N_10218);
nor U10865 (N_10865,N_10517,N_9833);
xnor U10866 (N_10866,N_10015,N_9629);
or U10867 (N_10867,N_10247,N_10095);
or U10868 (N_10868,N_9772,N_10652);
nor U10869 (N_10869,N_10348,N_10797);
nor U10870 (N_10870,N_10342,N_10303);
or U10871 (N_10871,N_10158,N_10101);
nor U10872 (N_10872,N_9783,N_10346);
or U10873 (N_10873,N_10767,N_10225);
and U10874 (N_10874,N_10774,N_10669);
or U10875 (N_10875,N_10073,N_9859);
xnor U10876 (N_10876,N_9687,N_10229);
xor U10877 (N_10877,N_10579,N_10049);
or U10878 (N_10878,N_10314,N_10270);
nor U10879 (N_10879,N_10093,N_9893);
nand U10880 (N_10880,N_9743,N_9790);
nand U10881 (N_10881,N_10081,N_10240);
and U10882 (N_10882,N_10102,N_9928);
and U10883 (N_10883,N_10174,N_10135);
xnor U10884 (N_10884,N_9717,N_9870);
nand U10885 (N_10885,N_10627,N_9974);
xnor U10886 (N_10886,N_10459,N_10242);
and U10887 (N_10887,N_10397,N_10037);
and U10888 (N_10888,N_10454,N_10491);
nor U10889 (N_10889,N_10315,N_10118);
and U10890 (N_10890,N_10018,N_10285);
and U10891 (N_10891,N_10526,N_9750);
nor U10892 (N_10892,N_10202,N_10142);
nand U10893 (N_10893,N_10542,N_10711);
nor U10894 (N_10894,N_10466,N_9746);
or U10895 (N_10895,N_9981,N_9637);
xor U10896 (N_10896,N_10349,N_10365);
nand U10897 (N_10897,N_9770,N_10362);
or U10898 (N_10898,N_10002,N_9899);
or U10899 (N_10899,N_10406,N_9773);
nor U10900 (N_10900,N_10237,N_9795);
nor U10901 (N_10901,N_10671,N_10035);
nor U10902 (N_10902,N_9791,N_9869);
nor U10903 (N_10903,N_9834,N_10781);
or U10904 (N_10904,N_10104,N_9966);
or U10905 (N_10905,N_10250,N_9967);
and U10906 (N_10906,N_9920,N_9780);
and U10907 (N_10907,N_10067,N_9956);
or U10908 (N_10908,N_10773,N_9642);
nor U10909 (N_10909,N_10167,N_9615);
or U10910 (N_10910,N_10273,N_10451);
or U10911 (N_10911,N_10771,N_10173);
xnor U10912 (N_10912,N_10511,N_10690);
xnor U10913 (N_10913,N_10044,N_10199);
xor U10914 (N_10914,N_10098,N_10039);
and U10915 (N_10915,N_10431,N_10324);
and U10916 (N_10916,N_10010,N_10207);
and U10917 (N_10917,N_10008,N_9602);
and U10918 (N_10918,N_9805,N_10291);
nand U10919 (N_10919,N_9989,N_10791);
nor U10920 (N_10920,N_9734,N_10709);
and U10921 (N_10921,N_10137,N_10496);
or U10922 (N_10922,N_10486,N_9821);
or U10923 (N_10923,N_10782,N_9829);
nor U10924 (N_10924,N_10519,N_10625);
xnor U10925 (N_10925,N_10283,N_10047);
nand U10926 (N_10926,N_9613,N_10765);
nor U10927 (N_10927,N_10335,N_10708);
and U10928 (N_10928,N_9900,N_9670);
xnor U10929 (N_10929,N_10379,N_10108);
nand U10930 (N_10930,N_10232,N_9965);
nand U10931 (N_10931,N_9999,N_10017);
and U10932 (N_10932,N_10779,N_9986);
nand U10933 (N_10933,N_9942,N_10739);
or U10934 (N_10934,N_10727,N_9646);
and U10935 (N_10935,N_9929,N_9864);
nor U10936 (N_10936,N_9857,N_10701);
or U10937 (N_10937,N_9603,N_10029);
nor U10938 (N_10938,N_9701,N_10464);
xnor U10939 (N_10939,N_9691,N_9946);
and U10940 (N_10940,N_10186,N_10377);
nand U10941 (N_10941,N_10417,N_9976);
nor U10942 (N_10942,N_10221,N_9838);
xnor U10943 (N_10943,N_9897,N_9902);
xor U10944 (N_10944,N_9910,N_10569);
and U10945 (N_10945,N_10347,N_9604);
nand U10946 (N_10946,N_10510,N_10087);
nand U10947 (N_10947,N_10339,N_10715);
or U10948 (N_10948,N_9718,N_10206);
or U10949 (N_10949,N_10027,N_9875);
nand U10950 (N_10950,N_9964,N_10665);
and U10951 (N_10951,N_9781,N_10021);
xnor U10952 (N_10952,N_10676,N_9837);
and U10953 (N_10953,N_10052,N_10793);
xnor U10954 (N_10954,N_10050,N_9903);
xnor U10955 (N_10955,N_9962,N_10673);
or U10956 (N_10956,N_10629,N_10148);
nor U10957 (N_10957,N_10630,N_9663);
and U10958 (N_10958,N_10649,N_10506);
nand U10959 (N_10959,N_9844,N_9605);
and U10960 (N_10960,N_9777,N_10507);
nand U10961 (N_10961,N_9804,N_10235);
xor U10962 (N_10962,N_9675,N_10505);
nor U10963 (N_10963,N_10109,N_9668);
nor U10964 (N_10964,N_9921,N_9798);
and U10965 (N_10965,N_10341,N_10488);
nand U10966 (N_10966,N_10605,N_10508);
xor U10967 (N_10967,N_10645,N_10063);
nand U10968 (N_10968,N_10518,N_10016);
nor U10969 (N_10969,N_9971,N_9803);
xnor U10970 (N_10970,N_10561,N_9891);
nor U10971 (N_10971,N_10144,N_10415);
xor U10972 (N_10972,N_10139,N_10162);
and U10973 (N_10973,N_10369,N_10180);
nor U10974 (N_10974,N_10043,N_9918);
nor U10975 (N_10975,N_9830,N_10187);
and U10976 (N_10976,N_10545,N_10521);
nand U10977 (N_10977,N_10736,N_10357);
and U10978 (N_10978,N_9968,N_10746);
nand U10979 (N_10979,N_10166,N_10011);
xnor U10980 (N_10980,N_10019,N_9722);
or U10981 (N_10981,N_10295,N_10544);
and U10982 (N_10982,N_10407,N_10145);
nor U10983 (N_10983,N_10654,N_10717);
xnor U10984 (N_10984,N_9708,N_9674);
xnor U10985 (N_10985,N_10317,N_10720);
nor U10986 (N_10986,N_10618,N_10045);
and U10987 (N_10987,N_10621,N_10306);
xor U10988 (N_10988,N_10006,N_9994);
nor U10989 (N_10989,N_10648,N_10344);
xnor U10990 (N_10990,N_10395,N_10410);
xor U10991 (N_10991,N_9737,N_9738);
nand U10992 (N_10992,N_10785,N_10394);
nand U10993 (N_10993,N_10492,N_9990);
nand U10994 (N_10994,N_9970,N_9885);
nand U10995 (N_10995,N_10435,N_10373);
nand U10996 (N_10996,N_10419,N_10132);
or U10997 (N_10997,N_10619,N_10688);
nor U10998 (N_10998,N_10402,N_9610);
or U10999 (N_10999,N_10684,N_10164);
nand U11000 (N_11000,N_9954,N_10522);
or U11001 (N_11001,N_10012,N_9649);
and U11002 (N_11002,N_9880,N_10340);
nand U11003 (N_11003,N_9665,N_10695);
and U11004 (N_11004,N_10732,N_9852);
or U11005 (N_11005,N_10565,N_9939);
or U11006 (N_11006,N_10420,N_10080);
or U11007 (N_11007,N_9930,N_10716);
and U11008 (N_11008,N_9644,N_9822);
and U11009 (N_11009,N_10091,N_9786);
nor U11010 (N_11010,N_9640,N_10128);
nand U11011 (N_11011,N_9895,N_10193);
nor U11012 (N_11012,N_9600,N_10735);
or U11013 (N_11013,N_10659,N_10552);
xnor U11014 (N_11014,N_10581,N_10024);
xor U11015 (N_11015,N_10764,N_9693);
xor U11016 (N_11016,N_10792,N_9630);
nand U11017 (N_11017,N_10473,N_9787);
and U11018 (N_11018,N_10177,N_10616);
nor U11019 (N_11019,N_9769,N_10243);
xor U11020 (N_11020,N_10712,N_10548);
nand U11021 (N_11021,N_9664,N_10493);
nor U11022 (N_11022,N_9694,N_10592);
or U11023 (N_11023,N_10130,N_10083);
and U11024 (N_11024,N_10650,N_10116);
nand U11025 (N_11025,N_9914,N_10543);
and U11026 (N_11026,N_10509,N_10770);
or U11027 (N_11027,N_10343,N_9779);
xnor U11028 (N_11028,N_9641,N_10667);
nand U11029 (N_11029,N_10168,N_9941);
xor U11030 (N_11030,N_10594,N_10430);
or U11031 (N_11031,N_10796,N_10598);
or U11032 (N_11032,N_10337,N_10070);
and U11033 (N_11033,N_10413,N_10481);
or U11034 (N_11034,N_10230,N_10117);
nand U11035 (N_11035,N_10704,N_10386);
xor U11036 (N_11036,N_9959,N_10133);
nand U11037 (N_11037,N_10147,N_10110);
xor U11038 (N_11038,N_10089,N_9661);
nand U11039 (N_11039,N_10401,N_9624);
and U11040 (N_11040,N_10758,N_10533);
and U11041 (N_11041,N_9901,N_10301);
nor U11042 (N_11042,N_9645,N_10191);
or U11043 (N_11043,N_10216,N_9998);
xnor U11044 (N_11044,N_9681,N_10375);
nand U11045 (N_11045,N_10224,N_9993);
and U11046 (N_11046,N_10299,N_10330);
xor U11047 (N_11047,N_10208,N_10361);
and U11048 (N_11048,N_9911,N_10528);
or U11049 (N_11049,N_10749,N_10352);
and U11050 (N_11050,N_10624,N_10723);
or U11051 (N_11051,N_10268,N_9997);
xnor U11052 (N_11052,N_10428,N_10244);
xor U11053 (N_11053,N_10609,N_10790);
nor U11054 (N_11054,N_10612,N_10638);
or U11055 (N_11055,N_10405,N_10563);
or U11056 (N_11056,N_10192,N_9720);
or U11057 (N_11057,N_9935,N_10153);
and U11058 (N_11058,N_9607,N_10575);
nor U11059 (N_11059,N_10307,N_9817);
nor U11060 (N_11060,N_10639,N_10190);
or U11061 (N_11061,N_9673,N_9877);
or U11062 (N_11062,N_9628,N_10033);
nand U11063 (N_11063,N_10560,N_10390);
nand U11064 (N_11064,N_10321,N_10189);
and U11065 (N_11065,N_10408,N_9806);
or U11066 (N_11066,N_10231,N_10429);
xnor U11067 (N_11067,N_10530,N_9625);
and U11068 (N_11068,N_10277,N_10079);
or U11069 (N_11069,N_9618,N_9705);
or U11070 (N_11070,N_9983,N_10280);
nand U11071 (N_11071,N_9872,N_10114);
nor U11072 (N_11072,N_10113,N_9706);
nor U11073 (N_11073,N_10274,N_10691);
xnor U11074 (N_11074,N_10571,N_10040);
and U11075 (N_11075,N_9807,N_9741);
and U11076 (N_11076,N_9889,N_9666);
and U11077 (N_11077,N_9688,N_9888);
nand U11078 (N_11078,N_10457,N_9656);
and U11079 (N_11079,N_10265,N_10127);
nand U11080 (N_11080,N_10768,N_10103);
xnor U11081 (N_11081,N_9862,N_9927);
or U11082 (N_11082,N_10640,N_10312);
and U11083 (N_11083,N_9842,N_10157);
nor U11084 (N_11084,N_10674,N_10185);
and U11085 (N_11085,N_9638,N_10078);
nand U11086 (N_11086,N_9831,N_10069);
xor U11087 (N_11087,N_9977,N_9703);
nor U11088 (N_11088,N_10743,N_10239);
or U11089 (N_11089,N_10220,N_10683);
or U11090 (N_11090,N_9756,N_9643);
or U11091 (N_11091,N_10706,N_10097);
nand U11092 (N_11092,N_10256,N_10411);
xor U11093 (N_11093,N_9723,N_9812);
nand U11094 (N_11094,N_9758,N_10119);
nand U11095 (N_11095,N_9736,N_9878);
nor U11096 (N_11096,N_10703,N_10692);
nor U11097 (N_11097,N_10651,N_10380);
xnor U11098 (N_11098,N_10175,N_10212);
xor U11099 (N_11099,N_10551,N_10246);
xor U11100 (N_11100,N_10574,N_9704);
nor U11101 (N_11101,N_9716,N_10267);
and U11102 (N_11102,N_10586,N_10182);
nor U11103 (N_11103,N_10799,N_9912);
and U11104 (N_11104,N_10595,N_10031);
xor U11105 (N_11105,N_10599,N_10534);
nand U11106 (N_11106,N_9802,N_10497);
nand U11107 (N_11107,N_9909,N_10356);
and U11108 (N_11108,N_10752,N_10210);
xnor U11109 (N_11109,N_9608,N_10353);
and U11110 (N_11110,N_9759,N_10022);
xor U11111 (N_11111,N_10151,N_10014);
xnor U11112 (N_11112,N_9952,N_10448);
nor U11113 (N_11113,N_9809,N_10282);
and U11114 (N_11114,N_10555,N_9898);
xnor U11115 (N_11115,N_9987,N_10311);
and U11116 (N_11116,N_9894,N_10516);
nor U11117 (N_11117,N_10276,N_10278);
or U11118 (N_11118,N_10553,N_10730);
nand U11119 (N_11119,N_10213,N_9606);
nor U11120 (N_11120,N_10440,N_10550);
or U11121 (N_11121,N_10786,N_9823);
nand U11122 (N_11122,N_10759,N_9616);
xnor U11123 (N_11123,N_10539,N_10458);
nand U11124 (N_11124,N_9868,N_9726);
or U11125 (N_11125,N_10580,N_9727);
or U11126 (N_11126,N_10724,N_9774);
or U11127 (N_11127,N_10741,N_10475);
and U11128 (N_11128,N_10060,N_10056);
nand U11129 (N_11129,N_10245,N_9683);
nand U11130 (N_11130,N_10500,N_9982);
xor U11131 (N_11131,N_9978,N_9980);
nand U11132 (N_11132,N_9813,N_9865);
nor U11133 (N_11133,N_10484,N_10359);
xor U11134 (N_11134,N_9733,N_9651);
nor U11135 (N_11135,N_9731,N_10750);
nor U11136 (N_11136,N_9876,N_10131);
nor U11137 (N_11137,N_10642,N_10065);
xor U11138 (N_11138,N_10179,N_9908);
or U11139 (N_11139,N_10381,N_9818);
nand U11140 (N_11140,N_9936,N_9794);
and U11141 (N_11141,N_9922,N_10409);
or U11142 (N_11142,N_10689,N_10628);
nor U11143 (N_11143,N_10476,N_9698);
xnor U11144 (N_11144,N_10698,N_10763);
and U11145 (N_11145,N_10068,N_10439);
nand U11146 (N_11146,N_10198,N_10587);
or U11147 (N_11147,N_10115,N_9655);
nand U11148 (N_11148,N_9695,N_10123);
nand U11149 (N_11149,N_10322,N_10718);
or U11150 (N_11150,N_9662,N_10613);
or U11151 (N_11151,N_10391,N_10610);
xor U11152 (N_11152,N_10634,N_10023);
and U11153 (N_11153,N_10432,N_10383);
or U11154 (N_11154,N_10234,N_10472);
and U11155 (N_11155,N_10470,N_10568);
xnor U11156 (N_11156,N_10748,N_10107);
and U11157 (N_11157,N_10490,N_10668);
nor U11158 (N_11158,N_10254,N_9719);
and U11159 (N_11159,N_9725,N_9826);
nand U11160 (N_11160,N_9755,N_10433);
and U11161 (N_11161,N_10456,N_10384);
and U11162 (N_11162,N_10072,N_9854);
and U11163 (N_11163,N_10152,N_10566);
or U11164 (N_11164,N_9846,N_9824);
xnor U11165 (N_11165,N_9700,N_9848);
xor U11166 (N_11166,N_9948,N_9680);
xnor U11167 (N_11167,N_10719,N_10392);
and U11168 (N_11168,N_9792,N_9947);
xor U11169 (N_11169,N_9940,N_10294);
nand U11170 (N_11170,N_10184,N_10096);
and U11171 (N_11171,N_9754,N_10251);
nor U11172 (N_11172,N_9633,N_9856);
xor U11173 (N_11173,N_9953,N_10092);
or U11174 (N_11174,N_10567,N_10358);
and U11175 (N_11175,N_10591,N_9742);
xnor U11176 (N_11176,N_10662,N_10209);
nor U11177 (N_11177,N_10557,N_10515);
or U11178 (N_11178,N_10535,N_10214);
and U11179 (N_11179,N_10363,N_10653);
nor U11180 (N_11180,N_10661,N_10057);
xor U11181 (N_11181,N_10281,N_10374);
or U11182 (N_11182,N_10351,N_10487);
nand U11183 (N_11183,N_9801,N_9884);
or U11184 (N_11184,N_10141,N_10755);
or U11185 (N_11185,N_10205,N_10685);
or U11186 (N_11186,N_9707,N_10693);
nor U11187 (N_11187,N_10197,N_10611);
xor U11188 (N_11188,N_9796,N_10121);
nor U11189 (N_11189,N_10154,N_9654);
and U11190 (N_11190,N_10279,N_9988);
nor U11191 (N_11191,N_10570,N_10778);
nor U11192 (N_11192,N_10248,N_10477);
and U11193 (N_11193,N_10004,N_9620);
xnor U11194 (N_11194,N_10125,N_9843);
nor U11195 (N_11195,N_9871,N_10094);
and U11196 (N_11196,N_10238,N_10672);
and U11197 (N_11197,N_10172,N_10762);
nor U11198 (N_11198,N_10412,N_10705);
nand U11199 (N_11199,N_9778,N_10228);
or U11200 (N_11200,N_10787,N_10414);
or U11201 (N_11201,N_10264,N_10577);
nor U11202 (N_11202,N_10597,N_10631);
and U11203 (N_11203,N_9647,N_10259);
and U11204 (N_11204,N_10734,N_10679);
xor U11205 (N_11205,N_10156,N_10664);
xor U11206 (N_11206,N_10041,N_10074);
nand U11207 (N_11207,N_10588,N_10200);
nand U11208 (N_11208,N_9890,N_10028);
or U11209 (N_11209,N_10760,N_9745);
nand U11210 (N_11210,N_10687,N_10626);
and U11211 (N_11211,N_10660,N_10169);
or U11212 (N_11212,N_10077,N_10088);
nor U11213 (N_11213,N_10416,N_10443);
xnor U11214 (N_11214,N_10636,N_10696);
and U11215 (N_11215,N_10656,N_10249);
or U11216 (N_11216,N_9631,N_10647);
and U11217 (N_11217,N_10071,N_9721);
nor U11218 (N_11218,N_10498,N_10769);
nor U11219 (N_11219,N_10319,N_10546);
xnor U11220 (N_11220,N_10502,N_10048);
or U11221 (N_11221,N_10742,N_9950);
xor U11222 (N_11222,N_9622,N_9682);
nand U11223 (N_11223,N_9763,N_9799);
nor U11224 (N_11224,N_10009,N_9963);
or U11225 (N_11225,N_10461,N_10170);
or U11226 (N_11226,N_10293,N_9652);
and U11227 (N_11227,N_10325,N_10617);
and U11228 (N_11228,N_9749,N_10001);
or U11229 (N_11229,N_10260,N_10426);
nor U11230 (N_11230,N_9621,N_9619);
or U11231 (N_11231,N_9767,N_10013);
xnor U11232 (N_11232,N_10155,N_10298);
nand U11233 (N_11233,N_9896,N_9827);
and U11234 (N_11234,N_10697,N_10053);
and U11235 (N_11235,N_9797,N_10304);
nand U11236 (N_11236,N_10478,N_10707);
nand U11237 (N_11237,N_10449,N_10075);
or U11238 (N_11238,N_9934,N_9776);
nor U11239 (N_11239,N_9860,N_10261);
and U11240 (N_11240,N_9969,N_10054);
and U11241 (N_11241,N_9808,N_10320);
nand U11242 (N_11242,N_10699,N_9601);
nor U11243 (N_11243,N_10255,N_9951);
and U11244 (N_11244,N_9765,N_10136);
or U11245 (N_11245,N_9992,N_10558);
nand U11246 (N_11246,N_9816,N_9784);
or U11247 (N_11247,N_10290,N_10495);
nand U11248 (N_11248,N_10404,N_10504);
nor U11249 (N_11249,N_10262,N_10140);
or U11250 (N_11250,N_10382,N_9714);
and U11251 (N_11251,N_10376,N_10494);
nand U11252 (N_11252,N_10622,N_9713);
nand U11253 (N_11253,N_10604,N_9917);
and U11254 (N_11254,N_10297,N_10453);
nand U11255 (N_11255,N_10331,N_9825);
nand U11256 (N_11256,N_10794,N_10424);
nand U11257 (N_11257,N_10780,N_10203);
xnor U11258 (N_11258,N_10757,N_9931);
and U11259 (N_11259,N_10713,N_9753);
or U11260 (N_11260,N_10418,N_10201);
or U11261 (N_11261,N_10427,N_9696);
nand U11262 (N_11262,N_10194,N_10666);
and U11263 (N_11263,N_10188,N_10657);
or U11264 (N_11264,N_10030,N_10556);
xnor U11265 (N_11265,N_10620,N_9887);
nand U11266 (N_11266,N_9979,N_10051);
nor U11267 (N_11267,N_10463,N_9752);
xor U11268 (N_11268,N_10305,N_9609);
or U11269 (N_11269,N_10585,N_9915);
or U11270 (N_11270,N_10161,N_9676);
nor U11271 (N_11271,N_10064,N_10350);
or U11272 (N_11272,N_10252,N_9867);
or U11273 (N_11273,N_9995,N_10236);
or U11274 (N_11274,N_10076,N_10465);
xnor U11275 (N_11275,N_9639,N_9669);
and U11276 (N_11276,N_9724,N_10393);
and U11277 (N_11277,N_9832,N_10503);
nand U11278 (N_11278,N_10761,N_10614);
nor U11279 (N_11279,N_10328,N_10288);
or U11280 (N_11280,N_10058,N_10789);
xor U11281 (N_11281,N_9658,N_9650);
or U11282 (N_11282,N_10334,N_9748);
xor U11283 (N_11283,N_10559,N_10036);
or U11284 (N_11284,N_10313,N_10007);
nor U11285 (N_11285,N_9861,N_10195);
nand U11286 (N_11286,N_10323,N_10150);
or U11287 (N_11287,N_10615,N_10005);
or U11288 (N_11288,N_10100,N_9849);
and U11289 (N_11289,N_9938,N_10738);
xnor U11290 (N_11290,N_10663,N_10474);
and U11291 (N_11291,N_10120,N_10514);
xnor U11292 (N_11292,N_10751,N_10554);
and U11293 (N_11293,N_10608,N_10452);
nand U11294 (N_11294,N_9850,N_10222);
nand U11295 (N_11295,N_9958,N_10355);
or U11296 (N_11296,N_9766,N_9635);
and U11297 (N_11297,N_9712,N_10446);
or U11298 (N_11298,N_9657,N_10112);
or U11299 (N_11299,N_10085,N_10633);
or U11300 (N_11300,N_10681,N_10784);
or U11301 (N_11301,N_10798,N_10042);
nor U11302 (N_11302,N_10606,N_10729);
nand U11303 (N_11303,N_10223,N_10385);
xor U11304 (N_11304,N_9728,N_10523);
xor U11305 (N_11305,N_9653,N_10700);
nor U11306 (N_11306,N_9961,N_10149);
xor U11307 (N_11307,N_10547,N_9762);
xnor U11308 (N_11308,N_9943,N_10602);
xnor U11309 (N_11309,N_9836,N_9984);
nand U11310 (N_11310,N_10308,N_10658);
or U11311 (N_11311,N_9711,N_10532);
or U11312 (N_11312,N_10286,N_9879);
and U11313 (N_11313,N_9632,N_9623);
nor U11314 (N_11314,N_10371,N_10677);
xor U11315 (N_11315,N_9847,N_9811);
nand U11316 (N_11316,N_9840,N_10272);
and U11317 (N_11317,N_10034,N_10783);
xnor U11318 (N_11318,N_10171,N_10524);
or U11319 (N_11319,N_10753,N_10644);
xnor U11320 (N_11320,N_9684,N_10576);
nand U11321 (N_11321,N_9771,N_10163);
xnor U11322 (N_11322,N_10725,N_10527);
or U11323 (N_11323,N_9699,N_10269);
nand U11324 (N_11324,N_10003,N_10572);
xor U11325 (N_11325,N_10434,N_10106);
or U11326 (N_11326,N_9835,N_9611);
nand U11327 (N_11327,N_10479,N_10084);
nor U11328 (N_11328,N_9904,N_10300);
or U11329 (N_11329,N_10399,N_10728);
or U11330 (N_11330,N_9973,N_10217);
xor U11331 (N_11331,N_9648,N_10367);
or U11332 (N_11332,N_9858,N_10455);
and U11333 (N_11333,N_10777,N_10489);
and U11334 (N_11334,N_9960,N_10124);
nand U11335 (N_11335,N_10513,N_10289);
or U11336 (N_11336,N_10646,N_10462);
and U11337 (N_11337,N_9785,N_9689);
nor U11338 (N_11338,N_10000,N_9757);
nand U11339 (N_11339,N_10525,N_9744);
nand U11340 (N_11340,N_9617,N_10271);
or U11341 (N_11341,N_10143,N_9685);
xor U11342 (N_11342,N_9916,N_9612);
nand U11343 (N_11343,N_10564,N_10204);
or U11344 (N_11344,N_9991,N_9659);
nand U11345 (N_11345,N_9732,N_9820);
xor U11346 (N_11346,N_10292,N_9873);
or U11347 (N_11347,N_9874,N_10529);
nor U11348 (N_11348,N_10159,N_10766);
or U11349 (N_11349,N_10731,N_9919);
and U11350 (N_11350,N_10483,N_10583);
nand U11351 (N_11351,N_10438,N_9739);
nand U11352 (N_11352,N_10795,N_10253);
nand U11353 (N_11353,N_9671,N_10450);
nand U11354 (N_11354,N_9923,N_10257);
nand U11355 (N_11355,N_10441,N_9955);
or U11356 (N_11356,N_10333,N_10686);
and U11357 (N_11357,N_9924,N_10082);
xnor U11358 (N_11358,N_10066,N_10090);
xor U11359 (N_11359,N_10061,N_9729);
xor U11360 (N_11360,N_9882,N_10302);
nand U11361 (N_11361,N_9815,N_10682);
nand U11362 (N_11362,N_10740,N_10398);
nor U11363 (N_11363,N_9905,N_10233);
and U11364 (N_11364,N_10694,N_10176);
and U11365 (N_11365,N_9692,N_9636);
and U11366 (N_11366,N_9828,N_9907);
xnor U11367 (N_11367,N_10445,N_10055);
or U11368 (N_11368,N_10756,N_10046);
nand U11369 (N_11369,N_10675,N_9972);
xor U11370 (N_11370,N_9855,N_10578);
nand U11371 (N_11371,N_9789,N_9866);
nor U11372 (N_11372,N_10744,N_9660);
and U11373 (N_11373,N_10396,N_9627);
xor U11374 (N_11374,N_10593,N_10600);
nand U11375 (N_11375,N_10772,N_10059);
and U11376 (N_11376,N_10275,N_10329);
xor U11377 (N_11377,N_10086,N_10316);
and U11378 (N_11378,N_9975,N_10105);
and U11379 (N_11379,N_10541,N_9751);
xor U11380 (N_11380,N_10226,N_9957);
and U11381 (N_11381,N_10372,N_10388);
and U11382 (N_11382,N_9667,N_10442);
xor U11383 (N_11383,N_10146,N_10062);
nand U11384 (N_11384,N_10423,N_9949);
nand U11385 (N_11385,N_10165,N_10338);
nor U11386 (N_11386,N_10227,N_10389);
nor U11387 (N_11387,N_9841,N_10296);
nor U11388 (N_11388,N_10714,N_10111);
xor U11389 (N_11389,N_10126,N_9863);
nand U11390 (N_11390,N_10368,N_10776);
nor U11391 (N_11391,N_9839,N_9800);
or U11392 (N_11392,N_10025,N_9881);
and U11393 (N_11393,N_10607,N_10623);
xor U11394 (N_11394,N_9735,N_9985);
or U11395 (N_11395,N_10266,N_9944);
nand U11396 (N_11396,N_9886,N_9853);
or U11397 (N_11397,N_9933,N_9810);
and U11398 (N_11398,N_10354,N_10467);
or U11399 (N_11399,N_10512,N_9926);
and U11400 (N_11400,N_10187,N_9737);
and U11401 (N_11401,N_10746,N_10592);
or U11402 (N_11402,N_10379,N_10439);
nand U11403 (N_11403,N_10449,N_9679);
nor U11404 (N_11404,N_10485,N_10447);
xnor U11405 (N_11405,N_10509,N_9927);
xnor U11406 (N_11406,N_9901,N_10558);
nor U11407 (N_11407,N_10593,N_9942);
and U11408 (N_11408,N_10130,N_10299);
or U11409 (N_11409,N_10670,N_9894);
and U11410 (N_11410,N_10502,N_9720);
or U11411 (N_11411,N_10454,N_10699);
or U11412 (N_11412,N_9897,N_9638);
nand U11413 (N_11413,N_10617,N_10594);
nor U11414 (N_11414,N_10212,N_10596);
and U11415 (N_11415,N_9968,N_10225);
nor U11416 (N_11416,N_9777,N_10636);
xnor U11417 (N_11417,N_10060,N_10782);
nor U11418 (N_11418,N_9933,N_9907);
or U11419 (N_11419,N_10007,N_10336);
xnor U11420 (N_11420,N_10438,N_10123);
xnor U11421 (N_11421,N_10094,N_10251);
or U11422 (N_11422,N_10272,N_10755);
and U11423 (N_11423,N_10219,N_10021);
or U11424 (N_11424,N_10576,N_10252);
nand U11425 (N_11425,N_10096,N_10331);
and U11426 (N_11426,N_9819,N_10039);
nand U11427 (N_11427,N_10109,N_9916);
or U11428 (N_11428,N_9905,N_10586);
nor U11429 (N_11429,N_10272,N_9743);
and U11430 (N_11430,N_9785,N_10604);
or U11431 (N_11431,N_10734,N_10597);
and U11432 (N_11432,N_10187,N_9695);
and U11433 (N_11433,N_10772,N_10475);
nor U11434 (N_11434,N_10715,N_10492);
nand U11435 (N_11435,N_9869,N_9931);
nand U11436 (N_11436,N_10485,N_10026);
nand U11437 (N_11437,N_10596,N_10564);
xor U11438 (N_11438,N_10772,N_10592);
xor U11439 (N_11439,N_10693,N_9744);
xor U11440 (N_11440,N_10269,N_9604);
nor U11441 (N_11441,N_9666,N_9646);
nor U11442 (N_11442,N_9866,N_10301);
or U11443 (N_11443,N_10205,N_10383);
nor U11444 (N_11444,N_10426,N_10733);
nor U11445 (N_11445,N_10770,N_10583);
and U11446 (N_11446,N_10171,N_10481);
xor U11447 (N_11447,N_10358,N_9911);
xor U11448 (N_11448,N_10504,N_9670);
and U11449 (N_11449,N_10483,N_10729);
or U11450 (N_11450,N_9873,N_10002);
xor U11451 (N_11451,N_9797,N_9787);
xor U11452 (N_11452,N_10216,N_9633);
nor U11453 (N_11453,N_9913,N_10498);
nor U11454 (N_11454,N_10497,N_10673);
nor U11455 (N_11455,N_9933,N_9609);
xnor U11456 (N_11456,N_10156,N_9665);
and U11457 (N_11457,N_10554,N_9959);
nand U11458 (N_11458,N_9848,N_9635);
and U11459 (N_11459,N_10612,N_10679);
xnor U11460 (N_11460,N_10273,N_9765);
or U11461 (N_11461,N_9956,N_10038);
or U11462 (N_11462,N_10782,N_9752);
or U11463 (N_11463,N_10158,N_10282);
xor U11464 (N_11464,N_10577,N_10453);
nand U11465 (N_11465,N_10233,N_9772);
nand U11466 (N_11466,N_10745,N_9731);
nor U11467 (N_11467,N_10240,N_10655);
and U11468 (N_11468,N_10358,N_10380);
nor U11469 (N_11469,N_10780,N_10274);
xor U11470 (N_11470,N_10699,N_9822);
and U11471 (N_11471,N_9947,N_10635);
and U11472 (N_11472,N_9946,N_9974);
or U11473 (N_11473,N_9674,N_9775);
nand U11474 (N_11474,N_9650,N_10649);
and U11475 (N_11475,N_10761,N_10771);
and U11476 (N_11476,N_10449,N_10436);
xor U11477 (N_11477,N_10762,N_10223);
xor U11478 (N_11478,N_10362,N_10659);
nor U11479 (N_11479,N_9707,N_10782);
and U11480 (N_11480,N_10088,N_10735);
and U11481 (N_11481,N_10624,N_10513);
nor U11482 (N_11482,N_10292,N_9961);
nand U11483 (N_11483,N_10576,N_10164);
nand U11484 (N_11484,N_10218,N_10082);
or U11485 (N_11485,N_9919,N_10646);
nor U11486 (N_11486,N_10388,N_10649);
or U11487 (N_11487,N_9975,N_10361);
xnor U11488 (N_11488,N_9708,N_10251);
xnor U11489 (N_11489,N_10417,N_10445);
nand U11490 (N_11490,N_10177,N_10473);
xor U11491 (N_11491,N_9657,N_10636);
xor U11492 (N_11492,N_10109,N_10699);
and U11493 (N_11493,N_10451,N_10203);
nor U11494 (N_11494,N_10440,N_9821);
xnor U11495 (N_11495,N_9745,N_9965);
xor U11496 (N_11496,N_9766,N_9897);
nand U11497 (N_11497,N_10596,N_10378);
nand U11498 (N_11498,N_10019,N_9924);
nor U11499 (N_11499,N_10516,N_10289);
and U11500 (N_11500,N_9717,N_10044);
or U11501 (N_11501,N_10468,N_10462);
or U11502 (N_11502,N_9930,N_10770);
nand U11503 (N_11503,N_10334,N_10344);
nor U11504 (N_11504,N_10737,N_10494);
and U11505 (N_11505,N_10389,N_10186);
and U11506 (N_11506,N_9714,N_10663);
nand U11507 (N_11507,N_10443,N_9660);
nor U11508 (N_11508,N_9790,N_10110);
and U11509 (N_11509,N_10090,N_10200);
nor U11510 (N_11510,N_9893,N_10233);
and U11511 (N_11511,N_10759,N_10453);
or U11512 (N_11512,N_9676,N_10570);
nor U11513 (N_11513,N_10175,N_10354);
or U11514 (N_11514,N_10692,N_10155);
or U11515 (N_11515,N_10791,N_10443);
and U11516 (N_11516,N_9749,N_9916);
xor U11517 (N_11517,N_9609,N_10682);
nor U11518 (N_11518,N_10387,N_10293);
nand U11519 (N_11519,N_10137,N_9800);
or U11520 (N_11520,N_10251,N_10111);
and U11521 (N_11521,N_10571,N_10406);
nand U11522 (N_11522,N_10715,N_9604);
and U11523 (N_11523,N_9716,N_10477);
xnor U11524 (N_11524,N_10545,N_9868);
nand U11525 (N_11525,N_10337,N_10216);
nand U11526 (N_11526,N_9960,N_10754);
nor U11527 (N_11527,N_9681,N_9932);
or U11528 (N_11528,N_9687,N_10504);
xor U11529 (N_11529,N_9764,N_10104);
nand U11530 (N_11530,N_10270,N_10437);
nor U11531 (N_11531,N_10733,N_10114);
xnor U11532 (N_11532,N_10745,N_10497);
nor U11533 (N_11533,N_10254,N_9725);
and U11534 (N_11534,N_9655,N_9710);
nor U11535 (N_11535,N_9632,N_10536);
xnor U11536 (N_11536,N_10133,N_10353);
and U11537 (N_11537,N_9616,N_10309);
xnor U11538 (N_11538,N_9968,N_10317);
or U11539 (N_11539,N_9947,N_9662);
nand U11540 (N_11540,N_10284,N_9826);
and U11541 (N_11541,N_10217,N_10286);
and U11542 (N_11542,N_9900,N_10548);
nor U11543 (N_11543,N_10209,N_10248);
xnor U11544 (N_11544,N_9759,N_9801);
xor U11545 (N_11545,N_10673,N_10786);
nor U11546 (N_11546,N_10233,N_9608);
and U11547 (N_11547,N_9772,N_10131);
nand U11548 (N_11548,N_10068,N_9895);
and U11549 (N_11549,N_10276,N_9857);
nand U11550 (N_11550,N_10295,N_10702);
nor U11551 (N_11551,N_9858,N_9784);
or U11552 (N_11552,N_10406,N_9682);
nor U11553 (N_11553,N_10641,N_10420);
xnor U11554 (N_11554,N_10725,N_10243);
nand U11555 (N_11555,N_10367,N_10491);
and U11556 (N_11556,N_10700,N_10013);
xnor U11557 (N_11557,N_10155,N_10426);
or U11558 (N_11558,N_10006,N_10091);
and U11559 (N_11559,N_10099,N_9914);
nand U11560 (N_11560,N_10267,N_10337);
and U11561 (N_11561,N_10290,N_10797);
and U11562 (N_11562,N_10735,N_10164);
or U11563 (N_11563,N_10407,N_9891);
and U11564 (N_11564,N_10799,N_10536);
or U11565 (N_11565,N_10469,N_10323);
and U11566 (N_11566,N_9679,N_9935);
nor U11567 (N_11567,N_10102,N_10224);
nor U11568 (N_11568,N_10683,N_10307);
nand U11569 (N_11569,N_10060,N_9799);
and U11570 (N_11570,N_10487,N_10764);
and U11571 (N_11571,N_10187,N_9759);
and U11572 (N_11572,N_10694,N_10668);
xnor U11573 (N_11573,N_10743,N_10020);
or U11574 (N_11574,N_10179,N_9747);
and U11575 (N_11575,N_9727,N_10306);
nor U11576 (N_11576,N_10473,N_10656);
or U11577 (N_11577,N_9862,N_10682);
or U11578 (N_11578,N_10506,N_10100);
nor U11579 (N_11579,N_9668,N_10338);
nand U11580 (N_11580,N_10621,N_10749);
and U11581 (N_11581,N_10017,N_10021);
and U11582 (N_11582,N_10713,N_10557);
and U11583 (N_11583,N_10239,N_9683);
nor U11584 (N_11584,N_9612,N_10718);
nand U11585 (N_11585,N_9865,N_10330);
and U11586 (N_11586,N_10045,N_10708);
xnor U11587 (N_11587,N_9673,N_10294);
or U11588 (N_11588,N_10509,N_10462);
nor U11589 (N_11589,N_9692,N_9647);
and U11590 (N_11590,N_9870,N_10329);
nand U11591 (N_11591,N_10757,N_9969);
or U11592 (N_11592,N_9609,N_10644);
nand U11593 (N_11593,N_9635,N_10372);
or U11594 (N_11594,N_10527,N_10448);
or U11595 (N_11595,N_10436,N_10332);
nand U11596 (N_11596,N_10241,N_10522);
and U11597 (N_11597,N_9638,N_10722);
or U11598 (N_11598,N_10359,N_10026);
nand U11599 (N_11599,N_10031,N_10225);
xnor U11600 (N_11600,N_9979,N_9666);
or U11601 (N_11601,N_9948,N_10321);
xor U11602 (N_11602,N_9915,N_10020);
xor U11603 (N_11603,N_10319,N_10419);
and U11604 (N_11604,N_10610,N_9890);
and U11605 (N_11605,N_10205,N_10006);
xor U11606 (N_11606,N_10267,N_10557);
xor U11607 (N_11607,N_9643,N_10785);
xor U11608 (N_11608,N_9608,N_10033);
and U11609 (N_11609,N_10634,N_10317);
or U11610 (N_11610,N_10633,N_10581);
or U11611 (N_11611,N_9916,N_10063);
or U11612 (N_11612,N_9965,N_10311);
or U11613 (N_11613,N_9930,N_9637);
xor U11614 (N_11614,N_10700,N_9672);
and U11615 (N_11615,N_10221,N_10642);
and U11616 (N_11616,N_9725,N_10671);
xor U11617 (N_11617,N_9627,N_10346);
nor U11618 (N_11618,N_9663,N_10149);
nand U11619 (N_11619,N_9615,N_10576);
nand U11620 (N_11620,N_10756,N_10410);
nor U11621 (N_11621,N_9894,N_10283);
xnor U11622 (N_11622,N_10670,N_9996);
nor U11623 (N_11623,N_10234,N_9884);
xor U11624 (N_11624,N_10554,N_9962);
or U11625 (N_11625,N_10208,N_10021);
or U11626 (N_11626,N_10771,N_10103);
nand U11627 (N_11627,N_10157,N_10633);
nor U11628 (N_11628,N_9867,N_9749);
nor U11629 (N_11629,N_10103,N_10181);
or U11630 (N_11630,N_9665,N_9992);
nor U11631 (N_11631,N_9865,N_10661);
nor U11632 (N_11632,N_10734,N_10214);
nor U11633 (N_11633,N_10479,N_10232);
xnor U11634 (N_11634,N_9900,N_10405);
or U11635 (N_11635,N_9764,N_10694);
or U11636 (N_11636,N_10351,N_10653);
nor U11637 (N_11637,N_9764,N_10312);
xnor U11638 (N_11638,N_10017,N_10407);
nor U11639 (N_11639,N_10427,N_9927);
or U11640 (N_11640,N_10415,N_9896);
nor U11641 (N_11641,N_9697,N_10223);
and U11642 (N_11642,N_9687,N_9803);
nor U11643 (N_11643,N_10290,N_9663);
nor U11644 (N_11644,N_10705,N_10318);
nand U11645 (N_11645,N_10692,N_9723);
and U11646 (N_11646,N_10321,N_10430);
and U11647 (N_11647,N_9786,N_10020);
or U11648 (N_11648,N_10215,N_10429);
nand U11649 (N_11649,N_10671,N_9941);
and U11650 (N_11650,N_10294,N_9900);
or U11651 (N_11651,N_9970,N_10503);
and U11652 (N_11652,N_10585,N_10357);
and U11653 (N_11653,N_10082,N_9949);
nor U11654 (N_11654,N_9854,N_9858);
or U11655 (N_11655,N_10759,N_9723);
nand U11656 (N_11656,N_10443,N_10588);
or U11657 (N_11657,N_10231,N_10173);
and U11658 (N_11658,N_10304,N_9893);
nor U11659 (N_11659,N_9966,N_9719);
or U11660 (N_11660,N_10570,N_10214);
and U11661 (N_11661,N_10155,N_10591);
nor U11662 (N_11662,N_10194,N_10145);
and U11663 (N_11663,N_10712,N_9836);
nand U11664 (N_11664,N_10458,N_9606);
nand U11665 (N_11665,N_10262,N_9862);
nor U11666 (N_11666,N_9926,N_9925);
nor U11667 (N_11667,N_9756,N_10374);
nor U11668 (N_11668,N_9661,N_10618);
xnor U11669 (N_11669,N_10333,N_10792);
xor U11670 (N_11670,N_9855,N_9605);
or U11671 (N_11671,N_9757,N_10274);
or U11672 (N_11672,N_10394,N_9881);
and U11673 (N_11673,N_9860,N_10131);
or U11674 (N_11674,N_10727,N_9628);
xnor U11675 (N_11675,N_9746,N_9688);
and U11676 (N_11676,N_10730,N_10696);
and U11677 (N_11677,N_10368,N_10160);
xor U11678 (N_11678,N_10485,N_10206);
nor U11679 (N_11679,N_9860,N_10702);
xnor U11680 (N_11680,N_10773,N_10162);
or U11681 (N_11681,N_10142,N_9992);
and U11682 (N_11682,N_10471,N_9714);
nor U11683 (N_11683,N_10663,N_10343);
nand U11684 (N_11684,N_10168,N_9713);
nor U11685 (N_11685,N_10784,N_10471);
nand U11686 (N_11686,N_10017,N_10179);
and U11687 (N_11687,N_9624,N_10264);
xor U11688 (N_11688,N_9695,N_10515);
and U11689 (N_11689,N_10326,N_10627);
nand U11690 (N_11690,N_10261,N_10124);
xnor U11691 (N_11691,N_9907,N_10245);
nor U11692 (N_11692,N_10317,N_10545);
or U11693 (N_11693,N_10473,N_10338);
nand U11694 (N_11694,N_10231,N_9746);
and U11695 (N_11695,N_10011,N_10109);
nor U11696 (N_11696,N_9976,N_10152);
or U11697 (N_11697,N_9828,N_10566);
nor U11698 (N_11698,N_10601,N_9946);
xor U11699 (N_11699,N_10306,N_9848);
and U11700 (N_11700,N_9987,N_10247);
xnor U11701 (N_11701,N_10571,N_10213);
nand U11702 (N_11702,N_9917,N_9840);
or U11703 (N_11703,N_9714,N_10794);
nor U11704 (N_11704,N_10405,N_10582);
or U11705 (N_11705,N_9757,N_9702);
nand U11706 (N_11706,N_10109,N_10088);
nand U11707 (N_11707,N_10225,N_9920);
nor U11708 (N_11708,N_9761,N_9725);
nor U11709 (N_11709,N_10747,N_9745);
nor U11710 (N_11710,N_10494,N_9977);
xnor U11711 (N_11711,N_10168,N_10064);
or U11712 (N_11712,N_9851,N_10625);
nand U11713 (N_11713,N_10595,N_10416);
nand U11714 (N_11714,N_9793,N_9809);
nor U11715 (N_11715,N_10312,N_10379);
nand U11716 (N_11716,N_10007,N_9724);
nor U11717 (N_11717,N_10523,N_10014);
or U11718 (N_11718,N_10250,N_10780);
nand U11719 (N_11719,N_9975,N_10699);
xnor U11720 (N_11720,N_9964,N_9806);
and U11721 (N_11721,N_9677,N_9617);
nand U11722 (N_11722,N_10568,N_10365);
or U11723 (N_11723,N_10401,N_9761);
or U11724 (N_11724,N_10393,N_10012);
and U11725 (N_11725,N_10547,N_10508);
nand U11726 (N_11726,N_9804,N_10632);
nor U11727 (N_11727,N_9650,N_10183);
or U11728 (N_11728,N_10717,N_9788);
and U11729 (N_11729,N_9885,N_10046);
or U11730 (N_11730,N_9602,N_10644);
nand U11731 (N_11731,N_9643,N_9940);
xor U11732 (N_11732,N_10006,N_10103);
or U11733 (N_11733,N_9931,N_10660);
xor U11734 (N_11734,N_10325,N_10188);
and U11735 (N_11735,N_10079,N_9775);
and U11736 (N_11736,N_10727,N_10373);
nand U11737 (N_11737,N_9939,N_10731);
nor U11738 (N_11738,N_10010,N_9877);
and U11739 (N_11739,N_9907,N_10462);
or U11740 (N_11740,N_10614,N_9612);
and U11741 (N_11741,N_10529,N_10521);
and U11742 (N_11742,N_10044,N_10473);
xor U11743 (N_11743,N_9830,N_9653);
xor U11744 (N_11744,N_10768,N_10419);
nand U11745 (N_11745,N_10239,N_10131);
nand U11746 (N_11746,N_9884,N_9921);
nor U11747 (N_11747,N_10185,N_9761);
and U11748 (N_11748,N_9822,N_10722);
nor U11749 (N_11749,N_10620,N_9914);
nor U11750 (N_11750,N_10277,N_10408);
xor U11751 (N_11751,N_9847,N_10226);
nand U11752 (N_11752,N_10431,N_9715);
and U11753 (N_11753,N_10006,N_9680);
nand U11754 (N_11754,N_10100,N_10691);
and U11755 (N_11755,N_10740,N_10479);
nand U11756 (N_11756,N_9918,N_9640);
and U11757 (N_11757,N_10050,N_10777);
or U11758 (N_11758,N_10571,N_10623);
or U11759 (N_11759,N_10717,N_9824);
nand U11760 (N_11760,N_9983,N_9908);
nor U11761 (N_11761,N_9968,N_10545);
and U11762 (N_11762,N_10264,N_10783);
nand U11763 (N_11763,N_9743,N_10016);
and U11764 (N_11764,N_10680,N_10308);
xor U11765 (N_11765,N_10633,N_9705);
nand U11766 (N_11766,N_10313,N_9707);
nand U11767 (N_11767,N_9745,N_9989);
xnor U11768 (N_11768,N_9702,N_10513);
xor U11769 (N_11769,N_9673,N_10101);
nor U11770 (N_11770,N_9788,N_9674);
or U11771 (N_11771,N_9764,N_10235);
or U11772 (N_11772,N_10381,N_9958);
nor U11773 (N_11773,N_10554,N_9684);
xnor U11774 (N_11774,N_9744,N_10400);
and U11775 (N_11775,N_10505,N_10677);
nor U11776 (N_11776,N_10276,N_10661);
nor U11777 (N_11777,N_10082,N_9657);
and U11778 (N_11778,N_10797,N_9637);
or U11779 (N_11779,N_10639,N_9938);
nor U11780 (N_11780,N_10185,N_10723);
or U11781 (N_11781,N_10734,N_9661);
nor U11782 (N_11782,N_9959,N_9932);
nor U11783 (N_11783,N_10610,N_10243);
or U11784 (N_11784,N_10456,N_10117);
nor U11785 (N_11785,N_10093,N_10338);
nor U11786 (N_11786,N_9805,N_9828);
nor U11787 (N_11787,N_10241,N_9762);
or U11788 (N_11788,N_10077,N_9688);
or U11789 (N_11789,N_9604,N_10474);
nand U11790 (N_11790,N_9760,N_9846);
nor U11791 (N_11791,N_10449,N_9622);
or U11792 (N_11792,N_10679,N_10335);
xor U11793 (N_11793,N_10451,N_9628);
nand U11794 (N_11794,N_9867,N_10364);
xnor U11795 (N_11795,N_10419,N_10752);
or U11796 (N_11796,N_10092,N_10315);
xor U11797 (N_11797,N_9843,N_10052);
nand U11798 (N_11798,N_9883,N_10194);
or U11799 (N_11799,N_9823,N_10484);
nand U11800 (N_11800,N_9952,N_10046);
nand U11801 (N_11801,N_10755,N_10576);
or U11802 (N_11802,N_10371,N_10650);
or U11803 (N_11803,N_10524,N_10737);
or U11804 (N_11804,N_9957,N_10284);
and U11805 (N_11805,N_10651,N_10036);
xnor U11806 (N_11806,N_9668,N_10025);
and U11807 (N_11807,N_10345,N_9623);
nor U11808 (N_11808,N_10707,N_9624);
xnor U11809 (N_11809,N_10367,N_10422);
and U11810 (N_11810,N_10772,N_10370);
xnor U11811 (N_11811,N_10674,N_9661);
or U11812 (N_11812,N_9761,N_10561);
and U11813 (N_11813,N_10540,N_10645);
xor U11814 (N_11814,N_10200,N_10539);
nand U11815 (N_11815,N_10142,N_9625);
nor U11816 (N_11816,N_9906,N_10596);
nor U11817 (N_11817,N_10121,N_9698);
and U11818 (N_11818,N_9646,N_10637);
nor U11819 (N_11819,N_9721,N_9606);
nand U11820 (N_11820,N_9947,N_9672);
and U11821 (N_11821,N_9831,N_9888);
and U11822 (N_11822,N_10347,N_10588);
and U11823 (N_11823,N_10790,N_9814);
nor U11824 (N_11824,N_10395,N_10057);
xor U11825 (N_11825,N_10676,N_9826);
xnor U11826 (N_11826,N_10572,N_10758);
and U11827 (N_11827,N_9935,N_9916);
nor U11828 (N_11828,N_10120,N_9615);
and U11829 (N_11829,N_10580,N_9819);
xnor U11830 (N_11830,N_9777,N_10765);
xor U11831 (N_11831,N_10504,N_10792);
xor U11832 (N_11832,N_10288,N_10152);
xnor U11833 (N_11833,N_10033,N_10646);
nor U11834 (N_11834,N_9923,N_10268);
or U11835 (N_11835,N_9765,N_9782);
nor U11836 (N_11836,N_9838,N_10069);
nor U11837 (N_11837,N_10083,N_10599);
xnor U11838 (N_11838,N_10157,N_9987);
and U11839 (N_11839,N_9922,N_10180);
or U11840 (N_11840,N_10569,N_9631);
and U11841 (N_11841,N_10666,N_9687);
nor U11842 (N_11842,N_9636,N_10736);
nor U11843 (N_11843,N_9975,N_9971);
xor U11844 (N_11844,N_9749,N_10415);
or U11845 (N_11845,N_10361,N_9856);
nand U11846 (N_11846,N_10393,N_10578);
nand U11847 (N_11847,N_10740,N_9892);
and U11848 (N_11848,N_9783,N_10438);
xnor U11849 (N_11849,N_9969,N_10402);
nor U11850 (N_11850,N_9763,N_10512);
nor U11851 (N_11851,N_10279,N_10507);
xnor U11852 (N_11852,N_10384,N_9639);
xnor U11853 (N_11853,N_10765,N_9817);
and U11854 (N_11854,N_10471,N_9638);
nor U11855 (N_11855,N_10029,N_9994);
and U11856 (N_11856,N_9970,N_9951);
nor U11857 (N_11857,N_9744,N_9926);
or U11858 (N_11858,N_9988,N_10297);
nor U11859 (N_11859,N_10389,N_9855);
xnor U11860 (N_11860,N_10181,N_10579);
nor U11861 (N_11861,N_10042,N_10465);
and U11862 (N_11862,N_10212,N_10337);
nor U11863 (N_11863,N_10601,N_10768);
xnor U11864 (N_11864,N_10263,N_9846);
xor U11865 (N_11865,N_9890,N_10154);
or U11866 (N_11866,N_10197,N_10078);
nor U11867 (N_11867,N_10159,N_9850);
nor U11868 (N_11868,N_10427,N_10198);
nand U11869 (N_11869,N_10728,N_10589);
or U11870 (N_11870,N_10273,N_9966);
nor U11871 (N_11871,N_10179,N_9613);
nor U11872 (N_11872,N_10167,N_10474);
nand U11873 (N_11873,N_9974,N_10011);
nor U11874 (N_11874,N_9816,N_10501);
xnor U11875 (N_11875,N_10129,N_10322);
and U11876 (N_11876,N_10284,N_10725);
xnor U11877 (N_11877,N_10077,N_9874);
and U11878 (N_11878,N_9920,N_10269);
and U11879 (N_11879,N_9903,N_9712);
or U11880 (N_11880,N_10736,N_10791);
and U11881 (N_11881,N_10681,N_10517);
nand U11882 (N_11882,N_10444,N_10729);
nor U11883 (N_11883,N_9639,N_9971);
or U11884 (N_11884,N_9660,N_10379);
nand U11885 (N_11885,N_9769,N_10200);
nor U11886 (N_11886,N_10570,N_9848);
nor U11887 (N_11887,N_10768,N_10694);
and U11888 (N_11888,N_9979,N_10405);
nand U11889 (N_11889,N_10422,N_9830);
and U11890 (N_11890,N_9678,N_10003);
xnor U11891 (N_11891,N_9747,N_10001);
nor U11892 (N_11892,N_9826,N_10582);
or U11893 (N_11893,N_10005,N_9663);
nor U11894 (N_11894,N_10382,N_9936);
nand U11895 (N_11895,N_9633,N_10145);
nor U11896 (N_11896,N_9870,N_10315);
nor U11897 (N_11897,N_10695,N_9636);
or U11898 (N_11898,N_9949,N_9952);
or U11899 (N_11899,N_10709,N_10728);
nor U11900 (N_11900,N_9637,N_10556);
nor U11901 (N_11901,N_10388,N_10403);
or U11902 (N_11902,N_10320,N_9611);
nand U11903 (N_11903,N_9635,N_10690);
xor U11904 (N_11904,N_10075,N_9865);
and U11905 (N_11905,N_10072,N_9959);
xnor U11906 (N_11906,N_10363,N_10503);
nor U11907 (N_11907,N_10223,N_9857);
nand U11908 (N_11908,N_9630,N_10250);
nor U11909 (N_11909,N_10372,N_10351);
or U11910 (N_11910,N_10719,N_10469);
and U11911 (N_11911,N_10242,N_9752);
or U11912 (N_11912,N_10021,N_10313);
nor U11913 (N_11913,N_10522,N_10436);
nand U11914 (N_11914,N_10309,N_9740);
and U11915 (N_11915,N_10450,N_10395);
and U11916 (N_11916,N_10707,N_10569);
or U11917 (N_11917,N_9804,N_10793);
nand U11918 (N_11918,N_10439,N_10542);
and U11919 (N_11919,N_10082,N_10536);
and U11920 (N_11920,N_10718,N_10043);
and U11921 (N_11921,N_9839,N_10425);
xor U11922 (N_11922,N_10681,N_10385);
nor U11923 (N_11923,N_10690,N_10351);
or U11924 (N_11924,N_9636,N_9972);
nand U11925 (N_11925,N_10286,N_9674);
and U11926 (N_11926,N_9829,N_10127);
nand U11927 (N_11927,N_10664,N_10129);
nand U11928 (N_11928,N_10099,N_9839);
nand U11929 (N_11929,N_10520,N_10442);
xor U11930 (N_11930,N_10787,N_10083);
and U11931 (N_11931,N_9961,N_9714);
nor U11932 (N_11932,N_10495,N_10168);
and U11933 (N_11933,N_9887,N_10288);
or U11934 (N_11934,N_10156,N_10104);
and U11935 (N_11935,N_10173,N_9977);
nand U11936 (N_11936,N_9687,N_10749);
nand U11937 (N_11937,N_10484,N_10441);
and U11938 (N_11938,N_10551,N_10252);
nand U11939 (N_11939,N_9999,N_9678);
or U11940 (N_11940,N_10182,N_10047);
and U11941 (N_11941,N_10634,N_9859);
or U11942 (N_11942,N_9996,N_9754);
and U11943 (N_11943,N_9849,N_9671);
and U11944 (N_11944,N_10625,N_10439);
nor U11945 (N_11945,N_9650,N_9855);
or U11946 (N_11946,N_10316,N_10603);
nor U11947 (N_11947,N_10512,N_10481);
xor U11948 (N_11948,N_10069,N_10552);
xor U11949 (N_11949,N_10530,N_10717);
or U11950 (N_11950,N_10783,N_9917);
nand U11951 (N_11951,N_10781,N_10291);
nand U11952 (N_11952,N_9807,N_10232);
xnor U11953 (N_11953,N_10282,N_10596);
and U11954 (N_11954,N_10525,N_10737);
and U11955 (N_11955,N_10356,N_9933);
and U11956 (N_11956,N_9624,N_9799);
or U11957 (N_11957,N_10240,N_10287);
nor U11958 (N_11958,N_9979,N_9871);
nand U11959 (N_11959,N_9911,N_10254);
or U11960 (N_11960,N_10404,N_10316);
xor U11961 (N_11961,N_10063,N_9778);
or U11962 (N_11962,N_9866,N_9952);
or U11963 (N_11963,N_10190,N_10646);
nand U11964 (N_11964,N_10719,N_10730);
xnor U11965 (N_11965,N_10293,N_10066);
and U11966 (N_11966,N_9975,N_10427);
or U11967 (N_11967,N_10460,N_10666);
nand U11968 (N_11968,N_10243,N_9623);
xor U11969 (N_11969,N_9833,N_10182);
xor U11970 (N_11970,N_9644,N_10199);
or U11971 (N_11971,N_10090,N_9612);
xnor U11972 (N_11972,N_9860,N_9904);
nor U11973 (N_11973,N_10463,N_10700);
nor U11974 (N_11974,N_10170,N_10023);
nand U11975 (N_11975,N_10122,N_10431);
nand U11976 (N_11976,N_10047,N_10272);
nor U11977 (N_11977,N_9960,N_10378);
or U11978 (N_11978,N_10502,N_10580);
nor U11979 (N_11979,N_9610,N_10358);
and U11980 (N_11980,N_10666,N_10602);
and U11981 (N_11981,N_9720,N_10341);
or U11982 (N_11982,N_10632,N_10499);
nor U11983 (N_11983,N_9755,N_10594);
xnor U11984 (N_11984,N_9861,N_10699);
xnor U11985 (N_11985,N_9763,N_10607);
and U11986 (N_11986,N_10058,N_10265);
nor U11987 (N_11987,N_10060,N_10283);
xor U11988 (N_11988,N_9904,N_10563);
xor U11989 (N_11989,N_9954,N_10306);
and U11990 (N_11990,N_9972,N_9652);
and U11991 (N_11991,N_10268,N_9684);
and U11992 (N_11992,N_10766,N_10389);
or U11993 (N_11993,N_9975,N_10350);
or U11994 (N_11994,N_10319,N_9735);
or U11995 (N_11995,N_10323,N_10799);
or U11996 (N_11996,N_10175,N_9907);
and U11997 (N_11997,N_10763,N_10530);
xor U11998 (N_11998,N_10013,N_9782);
nor U11999 (N_11999,N_10223,N_9960);
and U12000 (N_12000,N_11508,N_11310);
nor U12001 (N_12001,N_11984,N_11309);
and U12002 (N_12002,N_11082,N_11979);
nor U12003 (N_12003,N_11431,N_11237);
nor U12004 (N_12004,N_11316,N_11071);
nand U12005 (N_12005,N_10851,N_11534);
nand U12006 (N_12006,N_11946,N_10825);
and U12007 (N_12007,N_10831,N_11335);
xor U12008 (N_12008,N_11696,N_11297);
and U12009 (N_12009,N_11416,N_11328);
or U12010 (N_12010,N_11397,N_11379);
or U12011 (N_12011,N_11306,N_11827);
nand U12012 (N_12012,N_11111,N_10998);
xor U12013 (N_12013,N_11432,N_11807);
xnor U12014 (N_12014,N_11214,N_11831);
nand U12015 (N_12015,N_11065,N_11650);
nand U12016 (N_12016,N_11716,N_10928);
nand U12017 (N_12017,N_11825,N_11002);
or U12018 (N_12018,N_11277,N_10919);
nor U12019 (N_12019,N_11126,N_11725);
and U12020 (N_12020,N_11582,N_11899);
xnor U12021 (N_12021,N_11654,N_11786);
xor U12022 (N_12022,N_10983,N_11143);
nand U12023 (N_12023,N_10884,N_11391);
xor U12024 (N_12024,N_11801,N_11415);
or U12025 (N_12025,N_11729,N_11727);
nand U12026 (N_12026,N_11285,N_11498);
nor U12027 (N_12027,N_11469,N_11988);
or U12028 (N_12028,N_11781,N_11061);
xor U12029 (N_12029,N_11512,N_10853);
nand U12030 (N_12030,N_11934,N_11983);
nor U12031 (N_12031,N_11077,N_11336);
nor U12032 (N_12032,N_11278,N_11630);
and U12033 (N_12033,N_11457,N_11689);
xnor U12034 (N_12034,N_11063,N_11153);
nand U12035 (N_12035,N_11228,N_11000);
and U12036 (N_12036,N_11600,N_11364);
and U12037 (N_12037,N_10860,N_11787);
or U12038 (N_12038,N_11537,N_11872);
xor U12039 (N_12039,N_10913,N_11293);
xor U12040 (N_12040,N_10874,N_10981);
or U12041 (N_12041,N_11034,N_11499);
xor U12042 (N_12042,N_11251,N_10985);
xor U12043 (N_12043,N_10869,N_11514);
and U12044 (N_12044,N_10973,N_11884);
nor U12045 (N_12045,N_11171,N_11996);
nor U12046 (N_12046,N_11642,N_10861);
and U12047 (N_12047,N_11059,N_10866);
xor U12048 (N_12048,N_10976,N_11964);
nand U12049 (N_12049,N_10865,N_11181);
and U12050 (N_12050,N_11715,N_10814);
or U12051 (N_12051,N_11990,N_11795);
nand U12052 (N_12052,N_11957,N_11953);
xnor U12053 (N_12053,N_11064,N_10960);
and U12054 (N_12054,N_10999,N_11039);
nor U12055 (N_12055,N_11058,N_11791);
nand U12056 (N_12056,N_10835,N_11671);
nand U12057 (N_12057,N_11404,N_11012);
nor U12058 (N_12058,N_10822,N_11850);
and U12059 (N_12059,N_11331,N_11510);
nand U12060 (N_12060,N_11521,N_11579);
and U12061 (N_12061,N_11121,N_11652);
nand U12062 (N_12062,N_10809,N_11895);
xnor U12063 (N_12063,N_11806,N_11166);
and U12064 (N_12064,N_10878,N_10944);
nand U12065 (N_12065,N_11625,N_11922);
nor U12066 (N_12066,N_11770,N_11019);
and U12067 (N_12067,N_11322,N_11474);
or U12068 (N_12068,N_11665,N_11615);
or U12069 (N_12069,N_11644,N_11131);
xnor U12070 (N_12070,N_11095,N_11330);
and U12071 (N_12071,N_11461,N_11094);
and U12072 (N_12072,N_10832,N_11647);
nand U12073 (N_12073,N_11837,N_11243);
nor U12074 (N_12074,N_11334,N_11167);
or U12075 (N_12075,N_11805,N_11769);
and U12076 (N_12076,N_10958,N_10974);
nand U12077 (N_12077,N_11235,N_11538);
xor U12078 (N_12078,N_10885,N_11699);
or U12079 (N_12079,N_11317,N_10895);
nor U12080 (N_12080,N_11370,N_10932);
and U12081 (N_12081,N_10833,N_11042);
or U12082 (N_12082,N_11473,N_11023);
xor U12083 (N_12083,N_11004,N_11352);
nor U12084 (N_12084,N_10948,N_11426);
or U12085 (N_12085,N_11568,N_11728);
or U12086 (N_12086,N_11129,N_11950);
or U12087 (N_12087,N_11500,N_11174);
or U12088 (N_12088,N_10980,N_11666);
and U12089 (N_12089,N_11454,N_11680);
nand U12090 (N_12090,N_11467,N_11357);
and U12091 (N_12091,N_11907,N_10888);
or U12092 (N_12092,N_11854,N_11623);
nor U12093 (N_12093,N_11718,N_11157);
xnor U12094 (N_12094,N_10952,N_11810);
or U12095 (N_12095,N_11551,N_11458);
or U12096 (N_12096,N_11637,N_11075);
or U12097 (N_12097,N_11304,N_11993);
nand U12098 (N_12098,N_11120,N_10977);
nand U12099 (N_12099,N_11497,N_11299);
nor U12100 (N_12100,N_11160,N_11511);
or U12101 (N_12101,N_11029,N_11453);
nand U12102 (N_12102,N_11057,N_10996);
nor U12103 (N_12103,N_11970,N_11893);
xnor U12104 (N_12104,N_11954,N_10927);
or U12105 (N_12105,N_11219,N_11536);
nor U12106 (N_12106,N_11282,N_11387);
and U12107 (N_12107,N_11202,N_11267);
nand U12108 (N_12108,N_11502,N_11035);
and U12109 (N_12109,N_11616,N_11212);
nor U12110 (N_12110,N_11083,N_11303);
xnor U12111 (N_12111,N_11274,N_11909);
nand U12112 (N_12112,N_11930,N_11906);
or U12113 (N_12113,N_11005,N_10859);
nor U12114 (N_12114,N_11694,N_11835);
nor U12115 (N_12115,N_11460,N_11741);
and U12116 (N_12116,N_11532,N_11752);
nor U12117 (N_12117,N_11624,N_10921);
nor U12118 (N_12118,N_11130,N_11662);
and U12119 (N_12119,N_11448,N_11385);
nor U12120 (N_12120,N_10947,N_11584);
xnor U12121 (N_12121,N_11679,N_11221);
and U12122 (N_12122,N_11576,N_11485);
xnor U12123 (N_12123,N_11043,N_11503);
nand U12124 (N_12124,N_11258,N_11880);
nand U12125 (N_12125,N_11941,N_11535);
xor U12126 (N_12126,N_11275,N_11320);
or U12127 (N_12127,N_11686,N_11108);
nor U12128 (N_12128,N_11931,N_11505);
nor U12129 (N_12129,N_11692,N_11472);
and U12130 (N_12130,N_11001,N_11691);
and U12131 (N_12131,N_11560,N_11917);
nor U12132 (N_12132,N_10898,N_11719);
or U12133 (N_12133,N_11046,N_11972);
or U12134 (N_12134,N_11969,N_11009);
xor U12135 (N_12135,N_11127,N_11312);
nor U12136 (N_12136,N_11090,N_11627);
and U12137 (N_12137,N_11087,N_11829);
nor U12138 (N_12138,N_11084,N_11868);
and U12139 (N_12139,N_11150,N_10930);
nor U12140 (N_12140,N_11891,N_10810);
xor U12141 (N_12141,N_11247,N_11484);
xor U12142 (N_12142,N_11355,N_11667);
or U12143 (N_12143,N_10965,N_10972);
or U12144 (N_12144,N_11471,N_11832);
or U12145 (N_12145,N_11403,N_11173);
nand U12146 (N_12146,N_11550,N_11928);
and U12147 (N_12147,N_11670,N_11295);
or U12148 (N_12148,N_11981,N_11661);
nand U12149 (N_12149,N_11902,N_10867);
nor U12150 (N_12150,N_11390,N_11105);
nand U12151 (N_12151,N_11700,N_11421);
or U12152 (N_12152,N_10901,N_11062);
or U12153 (N_12153,N_11722,N_11755);
nor U12154 (N_12154,N_11447,N_11300);
and U12155 (N_12155,N_10934,N_11738);
and U12156 (N_12156,N_11554,N_11146);
or U12157 (N_12157,N_11115,N_11269);
xor U12158 (N_12158,N_10883,N_10801);
nor U12159 (N_12159,N_10955,N_11112);
and U12160 (N_12160,N_11091,N_11684);
nor U12161 (N_12161,N_11657,N_11635);
or U12162 (N_12162,N_11053,N_11268);
and U12163 (N_12163,N_11525,N_11669);
xnor U12164 (N_12164,N_10969,N_11271);
nand U12165 (N_12165,N_11855,N_11629);
nand U12166 (N_12166,N_11949,N_10845);
or U12167 (N_12167,N_11775,N_11339);
or U12168 (N_12168,N_11250,N_11375);
and U12169 (N_12169,N_10918,N_11956);
or U12170 (N_12170,N_11798,N_10922);
or U12171 (N_12171,N_11377,N_10802);
xnor U12172 (N_12172,N_11027,N_11528);
or U12173 (N_12173,N_10838,N_11555);
nand U12174 (N_12174,N_11726,N_11744);
and U12175 (N_12175,N_11351,N_11483);
and U12176 (N_12176,N_11276,N_10893);
nor U12177 (N_12177,N_11252,N_11997);
xor U12178 (N_12178,N_11638,N_10982);
and U12179 (N_12179,N_10992,N_11257);
xnor U12180 (N_12180,N_11631,N_11476);
xnor U12181 (N_12181,N_10836,N_10954);
and U12182 (N_12182,N_11601,N_11707);
and U12183 (N_12183,N_11688,N_11260);
or U12184 (N_12184,N_11543,N_11571);
and U12185 (N_12185,N_11305,N_11117);
or U12186 (N_12186,N_11687,N_10873);
nand U12187 (N_12187,N_11480,N_11881);
nor U12188 (N_12188,N_11778,N_11402);
nor U12189 (N_12189,N_11870,N_11583);
or U12190 (N_12190,N_11368,N_11927);
xor U12191 (N_12191,N_10827,N_11517);
or U12192 (N_12192,N_11937,N_11570);
and U12193 (N_12193,N_11055,N_11395);
xor U12194 (N_12194,N_10819,N_11493);
nand U12195 (N_12195,N_11109,N_11819);
nor U12196 (N_12196,N_11991,N_11343);
or U12197 (N_12197,N_10920,N_11459);
and U12198 (N_12198,N_11169,N_11010);
or U12199 (N_12199,N_11710,N_11045);
and U12200 (N_12200,N_10894,N_11158);
nand U12201 (N_12201,N_10896,N_11162);
nand U12202 (N_12202,N_11342,N_11420);
xor U12203 (N_12203,N_11489,N_11292);
or U12204 (N_12204,N_11313,N_10828);
nor U12205 (N_12205,N_11248,N_11749);
nor U12206 (N_12206,N_11877,N_11713);
nor U12207 (N_12207,N_11308,N_11302);
nor U12208 (N_12208,N_11605,N_11656);
xnor U12209 (N_12209,N_10936,N_10800);
xor U12210 (N_12210,N_11541,N_11332);
xnor U12211 (N_12211,N_11581,N_11976);
nand U12212 (N_12212,N_11040,N_11523);
and U12213 (N_12213,N_10905,N_11675);
xor U12214 (N_12214,N_11294,N_11464);
nor U12215 (N_12215,N_11178,N_11279);
nand U12216 (N_12216,N_11620,N_11041);
xnor U12217 (N_12217,N_11951,N_11182);
and U12218 (N_12218,N_11522,N_11333);
nand U12219 (N_12219,N_11712,N_11843);
or U12220 (N_12220,N_11764,N_11736);
or U12221 (N_12221,N_11080,N_11575);
nor U12222 (N_12222,N_11149,N_11967);
xnor U12223 (N_12223,N_11614,N_11735);
xnor U12224 (N_12224,N_11818,N_11871);
or U12225 (N_12225,N_11409,N_11834);
nor U12226 (N_12226,N_11663,N_11486);
xor U12227 (N_12227,N_11878,N_11549);
and U12228 (N_12228,N_11455,N_11353);
nand U12229 (N_12229,N_11233,N_11050);
nand U12230 (N_12230,N_11591,N_10986);
xor U12231 (N_12231,N_11721,N_11345);
or U12232 (N_12232,N_11933,N_11900);
or U12233 (N_12233,N_11873,N_11905);
and U12234 (N_12234,N_11841,N_10988);
and U12235 (N_12235,N_11366,N_10943);
xnor U12236 (N_12236,N_10891,N_11208);
nor U12237 (N_12237,N_11619,N_11446);
nand U12238 (N_12238,N_11093,N_11848);
xnor U12239 (N_12239,N_11589,N_11915);
and U12240 (N_12240,N_11546,N_11414);
xnor U12241 (N_12241,N_10806,N_11860);
and U12242 (N_12242,N_10911,N_11435);
xor U12243 (N_12243,N_11465,N_11626);
or U12244 (N_12244,N_11176,N_11865);
xor U12245 (N_12245,N_11020,N_11482);
and U12246 (N_12246,N_11847,N_11968);
and U12247 (N_12247,N_11759,N_10964);
or U12248 (N_12248,N_11200,N_11114);
nand U12249 (N_12249,N_11539,N_11490);
and U12250 (N_12250,N_11863,N_11923);
nand U12251 (N_12251,N_11265,N_11365);
or U12252 (N_12252,N_11369,N_11411);
nor U12253 (N_12253,N_11466,N_10849);
nor U12254 (N_12254,N_11363,N_10967);
xnor U12255 (N_12255,N_11542,N_11621);
nand U12256 (N_12256,N_10994,N_11596);
nand U12257 (N_12257,N_11098,N_11389);
or U12258 (N_12258,N_11441,N_11586);
nor U12259 (N_12259,N_11945,N_11141);
nor U12260 (N_12260,N_10815,N_10817);
nor U12261 (N_12261,N_11217,N_11659);
nor U12262 (N_12262,N_11226,N_10916);
or U12263 (N_12263,N_11753,N_11036);
nand U12264 (N_12264,N_11006,N_11740);
nor U12265 (N_12265,N_11481,N_11495);
nand U12266 (N_12266,N_11147,N_11188);
nand U12267 (N_12267,N_11883,N_11709);
and U12268 (N_12268,N_10857,N_10938);
nand U12269 (N_12269,N_11393,N_10995);
nor U12270 (N_12270,N_10813,N_11804);
nand U12271 (N_12271,N_11487,N_11745);
xnor U12272 (N_12272,N_11989,N_11030);
and U12273 (N_12273,N_11588,N_11428);
and U12274 (N_12274,N_11677,N_11761);
xnor U12275 (N_12275,N_11164,N_11401);
nor U12276 (N_12276,N_11216,N_11348);
and U12277 (N_12277,N_11919,N_11253);
xnor U12278 (N_12278,N_11693,N_11326);
and U12279 (N_12279,N_11540,N_11565);
xnor U12280 (N_12280,N_11918,N_11732);
nor U12281 (N_12281,N_11698,N_11245);
nor U12282 (N_12282,N_11018,N_11417);
and U12283 (N_12283,N_11144,N_10887);
and U12284 (N_12284,N_10876,N_11910);
nor U12285 (N_12285,N_11220,N_10991);
and U12286 (N_12286,N_11742,N_11594);
or U12287 (N_12287,N_11301,N_11206);
nor U12288 (N_12288,N_11737,N_11177);
or U12289 (N_12289,N_11885,N_11405);
and U12290 (N_12290,N_10931,N_11622);
nor U12291 (N_12291,N_11443,N_11561);
and U12292 (N_12292,N_11604,N_11789);
nand U12293 (N_12293,N_10870,N_11066);
nand U12294 (N_12294,N_11329,N_11307);
nor U12295 (N_12295,N_11232,N_11597);
nor U12296 (N_12296,N_11658,N_11724);
or U12297 (N_12297,N_10803,N_11664);
nand U12298 (N_12298,N_11152,N_11032);
and U12299 (N_12299,N_11985,N_11362);
and U12300 (N_12300,N_11383,N_11705);
nand U12301 (N_12301,N_11003,N_11189);
and U12302 (N_12302,N_10897,N_11122);
xor U12303 (N_12303,N_11739,N_11223);
and U12304 (N_12304,N_11099,N_11840);
nand U12305 (N_12305,N_11572,N_11430);
nand U12306 (N_12306,N_11204,N_11359);
nor U12307 (N_12307,N_10956,N_11506);
xnor U12308 (N_12308,N_11649,N_11168);
nor U12309 (N_12309,N_11321,N_11349);
xor U12310 (N_12310,N_11569,N_11074);
and U12311 (N_12311,N_11777,N_11185);
or U12312 (N_12312,N_11165,N_10879);
and U12313 (N_12313,N_11110,N_11283);
and U12314 (N_12314,N_11350,N_11051);
nand U12315 (N_12315,N_11288,N_11151);
or U12316 (N_12316,N_11504,N_11524);
nor U12317 (N_12317,N_11047,N_11874);
nand U12318 (N_12318,N_11452,N_11995);
nand U12319 (N_12319,N_11780,N_11672);
and U12320 (N_12320,N_11653,N_11270);
nand U12321 (N_12321,N_11125,N_11078);
and U12322 (N_12322,N_11450,N_11943);
xnor U12323 (N_12323,N_11592,N_11184);
nand U12324 (N_12324,N_11785,N_11346);
or U12325 (N_12325,N_11451,N_11824);
nor U12326 (N_12326,N_10997,N_11763);
or U12327 (N_12327,N_11648,N_11861);
or U12328 (N_12328,N_11747,N_10970);
nand U12329 (N_12329,N_11044,N_10963);
and U12330 (N_12330,N_11711,N_11384);
xnor U12331 (N_12331,N_11690,N_11231);
nand U12332 (N_12332,N_11708,N_11695);
nand U12333 (N_12333,N_11180,N_10823);
nand U12334 (N_12334,N_11776,N_10862);
or U12335 (N_12335,N_11932,N_11734);
nand U12336 (N_12336,N_11097,N_11618);
or U12337 (N_12337,N_11319,N_11340);
and U12338 (N_12338,N_11086,N_11449);
nand U12339 (N_12339,N_11903,N_11227);
nor U12340 (N_12340,N_11610,N_10892);
xor U12341 (N_12341,N_10903,N_11757);
and U12342 (N_12342,N_11992,N_11758);
and U12343 (N_12343,N_11136,N_11145);
or U12344 (N_12344,N_10909,N_11314);
nor U12345 (N_12345,N_11028,N_11398);
nand U12346 (N_12346,N_11566,N_10837);
nor U12347 (N_12347,N_11236,N_11007);
xnor U12348 (N_12348,N_11103,N_10826);
or U12349 (N_12349,N_11354,N_11820);
nand U12350 (N_12350,N_11193,N_11702);
or U12351 (N_12351,N_11731,N_11456);
and U12352 (N_12352,N_11636,N_11939);
xnor U12353 (N_12353,N_11286,N_11701);
nor U12354 (N_12354,N_11921,N_11971);
xor U12355 (N_12355,N_10949,N_10807);
nor U12356 (N_12356,N_11142,N_11697);
xnor U12357 (N_12357,N_11808,N_11124);
and U12358 (N_12358,N_10877,N_11423);
or U12359 (N_12359,N_10925,N_11845);
and U12360 (N_12360,N_11811,N_11386);
xor U12361 (N_12361,N_11913,N_11748);
nor U12362 (N_12362,N_11641,N_11017);
nor U12363 (N_12363,N_10914,N_11816);
and U12364 (N_12364,N_11085,N_10904);
nand U12365 (N_12365,N_11682,N_10852);
and U12366 (N_12366,N_11817,N_11215);
xnor U12367 (N_12367,N_10989,N_11526);
or U12368 (N_12368,N_10915,N_11407);
and U12369 (N_12369,N_11060,N_11914);
nand U12370 (N_12370,N_11730,N_11733);
and U12371 (N_12371,N_11205,N_11259);
nand U12372 (N_12372,N_10966,N_11199);
or U12373 (N_12373,N_11815,N_11507);
nor U12374 (N_12374,N_10990,N_10834);
or U12375 (N_12375,N_11519,N_11318);
and U12376 (N_12376,N_11133,N_11706);
or U12377 (N_12377,N_11138,N_11069);
xnor U12378 (N_12378,N_11496,N_11553);
xnor U12379 (N_12379,N_11544,N_11812);
nor U12380 (N_12380,N_11844,N_11024);
nand U12381 (N_12381,N_11961,N_11037);
and U12382 (N_12382,N_11054,N_11955);
and U12383 (N_12383,N_11925,N_11977);
and U12384 (N_12384,N_11929,N_11234);
nor U12385 (N_12385,N_11008,N_11547);
nand U12386 (N_12386,N_11263,N_10929);
and U12387 (N_12387,N_10975,N_11284);
nor U12388 (N_12388,N_10808,N_11170);
xor U12389 (N_12389,N_11876,N_11959);
or U12390 (N_12390,N_11358,N_11557);
nand U12391 (N_12391,N_11225,N_11839);
and U12392 (N_12392,N_11965,N_11272);
xor U12393 (N_12393,N_10900,N_11192);
nor U12394 (N_12394,N_11833,N_11425);
and U12395 (N_12395,N_10899,N_10881);
nand U12396 (N_12396,N_10880,N_11867);
nor U12397 (N_12397,N_11836,N_11823);
or U12398 (N_12398,N_11137,N_11021);
nand U12399 (N_12399,N_10945,N_10993);
nand U12400 (N_12400,N_11509,N_11952);
xor U12401 (N_12401,N_11793,N_11246);
or U12402 (N_12402,N_10939,N_11924);
nand U12403 (N_12403,N_10829,N_11113);
nor U12404 (N_12404,N_10933,N_11296);
xnor U12405 (N_12405,N_11790,N_11378);
nor U12406 (N_12406,N_11862,N_10805);
nor U12407 (N_12407,N_11374,N_11978);
and U12408 (N_12408,N_10910,N_11849);
xor U12409 (N_12409,N_11073,N_11750);
nor U12410 (N_12410,N_11942,N_11559);
nand U12411 (N_12411,N_11797,N_11244);
or U12412 (N_12412,N_11574,N_11545);
and U12413 (N_12413,N_11261,N_11768);
or U12414 (N_12414,N_11118,N_11864);
or U12415 (N_12415,N_11249,N_11645);
and U12416 (N_12416,N_10951,N_11935);
nor U12417 (N_12417,N_10950,N_11372);
and U12418 (N_12418,N_11218,N_11381);
nand U12419 (N_12419,N_11888,N_11894);
nor U12420 (N_12420,N_11119,N_11762);
xor U12421 (N_12421,N_11161,N_11014);
or U12422 (N_12422,N_11760,N_11291);
and U12423 (N_12423,N_11580,N_11940);
or U12424 (N_12424,N_10889,N_11281);
or U12425 (N_12425,N_10912,N_10856);
xnor U12426 (N_12426,N_11606,N_11478);
nand U12427 (N_12427,N_11774,N_11767);
nor U12428 (N_12428,N_10847,N_11194);
nor U12429 (N_12429,N_10987,N_11866);
or U12430 (N_12430,N_11643,N_11814);
and U12431 (N_12431,N_11974,N_11239);
nand U12432 (N_12432,N_11429,N_11016);
xnor U12433 (N_12433,N_10804,N_11463);
or U12434 (N_12434,N_10962,N_11958);
and U12435 (N_12435,N_10818,N_10941);
xor U12436 (N_12436,N_10926,N_10841);
and U12437 (N_12437,N_10882,N_11563);
nor U12438 (N_12438,N_11183,N_11593);
nand U12439 (N_12439,N_11361,N_11765);
and U12440 (N_12440,N_11963,N_10959);
nor U12441 (N_12441,N_11548,N_11821);
nor U12442 (N_12442,N_11025,N_11187);
nor U12443 (N_12443,N_10843,N_11628);
xor U12444 (N_12444,N_11186,N_10961);
and U12445 (N_12445,N_10935,N_11533);
nor U12446 (N_12446,N_11515,N_11324);
nor U12447 (N_12447,N_11201,N_11723);
nor U12448 (N_12448,N_11792,N_11516);
nor U12449 (N_12449,N_11609,N_11338);
xnor U12450 (N_12450,N_10830,N_11678);
nor U12451 (N_12451,N_10984,N_10871);
nor U12452 (N_12452,N_11031,N_11681);
xor U12453 (N_12453,N_10937,N_11373);
xnor U12454 (N_12454,N_11813,N_11879);
or U12455 (N_12455,N_11298,N_11424);
and U12456 (N_12456,N_11238,N_11102);
xor U12457 (N_12457,N_11273,N_11107);
nand U12458 (N_12458,N_10846,N_11155);
and U12459 (N_12459,N_11280,N_11966);
or U12460 (N_12460,N_11809,N_11886);
or U12461 (N_12461,N_10890,N_11327);
nand U12462 (N_12462,N_11056,N_11897);
nor U12463 (N_12463,N_11222,N_10917);
xor U12464 (N_12464,N_11026,N_11756);
xor U12465 (N_12465,N_11049,N_11828);
nor U12466 (N_12466,N_11889,N_11901);
nor U12467 (N_12467,N_11419,N_11088);
or U12468 (N_12468,N_11926,N_11717);
nand U12469 (N_12469,N_11772,N_11987);
or U12470 (N_12470,N_11191,N_11800);
xor U12471 (N_12471,N_11564,N_11360);
and U12472 (N_12472,N_10863,N_11494);
nand U12473 (N_12473,N_11052,N_11773);
and U12474 (N_12474,N_10811,N_11139);
nor U12475 (N_12475,N_11079,N_11676);
nor U12476 (N_12476,N_10858,N_11356);
or U12477 (N_12477,N_11175,N_11822);
xnor U12478 (N_12478,N_11197,N_11148);
nand U12479 (N_12479,N_11788,N_10923);
nor U12480 (N_12480,N_11646,N_11392);
xor U12481 (N_12481,N_11068,N_11096);
or U12482 (N_12482,N_11617,N_10906);
xnor U12483 (N_12483,N_10848,N_11033);
and U12484 (N_12484,N_11936,N_11412);
nor U12485 (N_12485,N_11089,N_11577);
and U12486 (N_12486,N_11999,N_11224);
or U12487 (N_12487,N_11944,N_10946);
and U12488 (N_12488,N_11703,N_11433);
and U12489 (N_12489,N_11887,N_11556);
and U12490 (N_12490,N_11254,N_11771);
or U12491 (N_12491,N_11962,N_10924);
xnor U12492 (N_12492,N_10953,N_11890);
nand U12493 (N_12493,N_11802,N_11266);
nor U12494 (N_12494,N_10816,N_11196);
or U12495 (N_12495,N_10908,N_11070);
xor U12496 (N_12496,N_11852,N_10820);
or U12497 (N_12497,N_11858,N_11229);
or U12498 (N_12498,N_11857,N_10855);
nand U12499 (N_12499,N_11746,N_11916);
xor U12500 (N_12500,N_11264,N_11067);
xor U12501 (N_12501,N_10850,N_11683);
xor U12502 (N_12502,N_11973,N_11599);
nand U12503 (N_12503,N_11492,N_11994);
nor U12504 (N_12504,N_11655,N_11567);
nand U12505 (N_12505,N_11948,N_11896);
and U12506 (N_12506,N_10907,N_10978);
nor U12507 (N_12507,N_11960,N_11634);
and U12508 (N_12508,N_11578,N_11347);
nand U12509 (N_12509,N_11826,N_11529);
and U12510 (N_12510,N_11337,N_10864);
nor U12511 (N_12511,N_11595,N_11437);
nor U12512 (N_12512,N_11408,N_10875);
and U12513 (N_12513,N_10824,N_11190);
nand U12514 (N_12514,N_11904,N_11602);
and U12515 (N_12515,N_11132,N_11444);
and U12516 (N_12516,N_11323,N_11598);
xor U12517 (N_12517,N_11341,N_11530);
nand U12518 (N_12518,N_11325,N_11830);
nand U12519 (N_12519,N_11491,N_11851);
xnor U12520 (N_12520,N_11908,N_11607);
nor U12521 (N_12521,N_11660,N_11195);
and U12522 (N_12522,N_11982,N_11668);
and U12523 (N_12523,N_11633,N_11552);
xor U12524 (N_12524,N_11783,N_11869);
xnor U12525 (N_12525,N_11438,N_11072);
xor U12526 (N_12526,N_11803,N_11673);
or U12527 (N_12527,N_11975,N_11242);
or U12528 (N_12528,N_11399,N_11920);
and U12529 (N_12529,N_10839,N_11048);
nor U12530 (N_12530,N_11856,N_11140);
or U12531 (N_12531,N_11784,N_11290);
nor U12532 (N_12532,N_11163,N_11892);
nor U12533 (N_12533,N_11106,N_11376);
nor U12534 (N_12534,N_11442,N_11766);
xnor U12535 (N_12535,N_11853,N_10840);
nand U12536 (N_12536,N_11603,N_10902);
xnor U12537 (N_12537,N_11198,N_11859);
nand U12538 (N_12538,N_11123,N_11400);
and U12539 (N_12539,N_11846,N_11782);
and U12540 (N_12540,N_11640,N_11685);
or U12541 (N_12541,N_11256,N_11898);
and U12542 (N_12542,N_11380,N_11875);
or U12543 (N_12543,N_11262,N_11531);
or U12544 (N_12544,N_11427,N_11445);
and U12545 (N_12545,N_11468,N_11311);
or U12546 (N_12546,N_11475,N_11720);
nand U12547 (N_12547,N_11612,N_10940);
xnor U12548 (N_12548,N_11394,N_11590);
nor U12549 (N_12549,N_10886,N_11315);
nor U12550 (N_12550,N_11513,N_11396);
nand U12551 (N_12551,N_11172,N_11799);
or U12552 (N_12552,N_10812,N_11092);
nand U12553 (N_12553,N_11573,N_11207);
xnor U12554 (N_12554,N_10872,N_11488);
or U12555 (N_12555,N_11213,N_11128);
and U12556 (N_12556,N_11651,N_11211);
nand U12557 (N_12557,N_11704,N_11585);
xnor U12558 (N_12558,N_11439,N_11639);
xor U12559 (N_12559,N_11527,N_11794);
nor U12560 (N_12560,N_10942,N_10842);
xor U12561 (N_12561,N_11367,N_11100);
nor U12562 (N_12562,N_11101,N_11608);
and U12563 (N_12563,N_11135,N_11611);
nor U12564 (N_12564,N_11912,N_11754);
xnor U12565 (N_12565,N_11134,N_11440);
or U12566 (N_12566,N_11156,N_11240);
nor U12567 (N_12567,N_11081,N_11518);
xnor U12568 (N_12568,N_11422,N_11410);
xor U12569 (N_12569,N_11013,N_11255);
nor U12570 (N_12570,N_11751,N_11674);
xor U12571 (N_12571,N_11159,N_11462);
and U12572 (N_12572,N_11986,N_11938);
xnor U12573 (N_12573,N_11911,N_11076);
xnor U12574 (N_12574,N_11210,N_10844);
nand U12575 (N_12575,N_11838,N_11388);
or U12576 (N_12576,N_11104,N_11479);
xor U12577 (N_12577,N_11413,N_11015);
nor U12578 (N_12578,N_10979,N_11289);
nor U12579 (N_12579,N_11562,N_11022);
xnor U12580 (N_12580,N_11882,N_11434);
xor U12581 (N_12581,N_10821,N_11406);
xor U12582 (N_12582,N_11179,N_11558);
nand U12583 (N_12583,N_10854,N_11241);
nor U12584 (N_12584,N_11371,N_11947);
or U12585 (N_12585,N_11796,N_11980);
and U12586 (N_12586,N_11779,N_10957);
or U12587 (N_12587,N_11714,N_11743);
and U12588 (N_12588,N_11587,N_11436);
nor U12589 (N_12589,N_11209,N_11501);
nand U12590 (N_12590,N_11842,N_11613);
or U12591 (N_12591,N_10968,N_11344);
and U12592 (N_12592,N_11520,N_11477);
xor U12593 (N_12593,N_11230,N_11418);
nand U12594 (N_12594,N_11998,N_10971);
or U12595 (N_12595,N_11470,N_11382);
nand U12596 (N_12596,N_11287,N_11154);
and U12597 (N_12597,N_11011,N_10868);
or U12598 (N_12598,N_11116,N_11632);
xnor U12599 (N_12599,N_11203,N_11038);
nor U12600 (N_12600,N_11357,N_11439);
xnor U12601 (N_12601,N_11648,N_11350);
or U12602 (N_12602,N_10833,N_11669);
xor U12603 (N_12603,N_11020,N_11627);
nand U12604 (N_12604,N_11214,N_11222);
and U12605 (N_12605,N_11181,N_11444);
nor U12606 (N_12606,N_10941,N_11565);
or U12607 (N_12607,N_11584,N_11105);
nand U12608 (N_12608,N_11119,N_10871);
and U12609 (N_12609,N_11704,N_10849);
and U12610 (N_12610,N_10891,N_11074);
nand U12611 (N_12611,N_10805,N_11261);
xor U12612 (N_12612,N_11544,N_11541);
and U12613 (N_12613,N_11905,N_11503);
nor U12614 (N_12614,N_10913,N_11057);
nor U12615 (N_12615,N_11254,N_11018);
xnor U12616 (N_12616,N_11284,N_11959);
nand U12617 (N_12617,N_11763,N_11554);
nand U12618 (N_12618,N_11035,N_11840);
nor U12619 (N_12619,N_11192,N_11047);
and U12620 (N_12620,N_11039,N_11711);
or U12621 (N_12621,N_11773,N_11328);
xor U12622 (N_12622,N_11378,N_11238);
xnor U12623 (N_12623,N_11032,N_11154);
and U12624 (N_12624,N_11233,N_11685);
or U12625 (N_12625,N_11621,N_11650);
nand U12626 (N_12626,N_11869,N_11245);
xor U12627 (N_12627,N_11336,N_11036);
xor U12628 (N_12628,N_10959,N_11406);
or U12629 (N_12629,N_11111,N_11713);
and U12630 (N_12630,N_11274,N_11505);
and U12631 (N_12631,N_11774,N_11501);
nand U12632 (N_12632,N_11613,N_11289);
nor U12633 (N_12633,N_11100,N_11565);
or U12634 (N_12634,N_11331,N_11393);
nand U12635 (N_12635,N_11475,N_11686);
nand U12636 (N_12636,N_11450,N_11980);
and U12637 (N_12637,N_11998,N_11832);
nor U12638 (N_12638,N_10943,N_11406);
nand U12639 (N_12639,N_11153,N_11459);
nand U12640 (N_12640,N_11959,N_11016);
or U12641 (N_12641,N_11818,N_11143);
nor U12642 (N_12642,N_11104,N_11322);
nor U12643 (N_12643,N_11603,N_11342);
and U12644 (N_12644,N_11265,N_11127);
nor U12645 (N_12645,N_11889,N_11609);
nand U12646 (N_12646,N_11448,N_11518);
or U12647 (N_12647,N_11738,N_10810);
nand U12648 (N_12648,N_10946,N_11263);
or U12649 (N_12649,N_11143,N_11454);
or U12650 (N_12650,N_11153,N_11803);
nor U12651 (N_12651,N_11697,N_11736);
and U12652 (N_12652,N_11226,N_11287);
nand U12653 (N_12653,N_11547,N_10904);
and U12654 (N_12654,N_11871,N_11953);
nand U12655 (N_12655,N_11113,N_11875);
nand U12656 (N_12656,N_11183,N_11391);
nor U12657 (N_12657,N_10803,N_11299);
or U12658 (N_12658,N_10971,N_10937);
nor U12659 (N_12659,N_11689,N_11580);
nor U12660 (N_12660,N_11877,N_11946);
or U12661 (N_12661,N_10869,N_11151);
nand U12662 (N_12662,N_10915,N_11869);
nor U12663 (N_12663,N_11165,N_11302);
nand U12664 (N_12664,N_11372,N_11191);
xnor U12665 (N_12665,N_11097,N_11389);
nand U12666 (N_12666,N_10899,N_11660);
xor U12667 (N_12667,N_11632,N_11607);
or U12668 (N_12668,N_11553,N_11677);
nand U12669 (N_12669,N_11929,N_11922);
nand U12670 (N_12670,N_11103,N_11196);
xor U12671 (N_12671,N_11512,N_11236);
xor U12672 (N_12672,N_11299,N_11042);
and U12673 (N_12673,N_11998,N_11592);
nand U12674 (N_12674,N_11956,N_11416);
and U12675 (N_12675,N_11781,N_11021);
xor U12676 (N_12676,N_11631,N_11194);
and U12677 (N_12677,N_11889,N_11430);
xor U12678 (N_12678,N_11127,N_11638);
and U12679 (N_12679,N_11008,N_10829);
nand U12680 (N_12680,N_11599,N_11940);
nor U12681 (N_12681,N_11478,N_11529);
or U12682 (N_12682,N_11264,N_11144);
nor U12683 (N_12683,N_10867,N_10991);
and U12684 (N_12684,N_11775,N_11122);
or U12685 (N_12685,N_11907,N_11068);
nand U12686 (N_12686,N_11212,N_11651);
xor U12687 (N_12687,N_11732,N_11686);
xor U12688 (N_12688,N_10941,N_11806);
nand U12689 (N_12689,N_11038,N_11842);
nor U12690 (N_12690,N_11151,N_10953);
xnor U12691 (N_12691,N_11660,N_11336);
nor U12692 (N_12692,N_11401,N_10841);
or U12693 (N_12693,N_11338,N_11301);
nor U12694 (N_12694,N_11710,N_11320);
xor U12695 (N_12695,N_11952,N_11853);
and U12696 (N_12696,N_11498,N_11525);
nor U12697 (N_12697,N_10995,N_11811);
xnor U12698 (N_12698,N_11575,N_11131);
xnor U12699 (N_12699,N_11545,N_11063);
or U12700 (N_12700,N_11279,N_11373);
nand U12701 (N_12701,N_11343,N_11538);
and U12702 (N_12702,N_11498,N_11299);
or U12703 (N_12703,N_11806,N_11695);
xor U12704 (N_12704,N_11992,N_11988);
nand U12705 (N_12705,N_11627,N_11495);
or U12706 (N_12706,N_11968,N_11362);
xnor U12707 (N_12707,N_10826,N_11761);
nand U12708 (N_12708,N_11027,N_11541);
nand U12709 (N_12709,N_11684,N_11271);
and U12710 (N_12710,N_11331,N_11278);
nand U12711 (N_12711,N_10950,N_11241);
or U12712 (N_12712,N_11265,N_11058);
and U12713 (N_12713,N_11007,N_11064);
nand U12714 (N_12714,N_11219,N_10919);
or U12715 (N_12715,N_11000,N_10923);
and U12716 (N_12716,N_11218,N_11073);
nand U12717 (N_12717,N_11318,N_11819);
xor U12718 (N_12718,N_11506,N_11941);
and U12719 (N_12719,N_11680,N_11823);
xnor U12720 (N_12720,N_11071,N_11474);
or U12721 (N_12721,N_11784,N_11268);
or U12722 (N_12722,N_11265,N_11151);
nor U12723 (N_12723,N_11878,N_10924);
and U12724 (N_12724,N_11383,N_11080);
or U12725 (N_12725,N_10937,N_11797);
nor U12726 (N_12726,N_11006,N_10878);
and U12727 (N_12727,N_11130,N_11445);
or U12728 (N_12728,N_11882,N_10926);
and U12729 (N_12729,N_10866,N_10896);
and U12730 (N_12730,N_11454,N_11893);
or U12731 (N_12731,N_10997,N_11700);
nor U12732 (N_12732,N_11618,N_11977);
or U12733 (N_12733,N_11370,N_11915);
or U12734 (N_12734,N_10886,N_11821);
nand U12735 (N_12735,N_11714,N_11586);
nor U12736 (N_12736,N_11849,N_11691);
nand U12737 (N_12737,N_11558,N_11819);
and U12738 (N_12738,N_11061,N_11368);
nor U12739 (N_12739,N_11926,N_11455);
and U12740 (N_12740,N_10890,N_11029);
or U12741 (N_12741,N_11790,N_11300);
or U12742 (N_12742,N_11160,N_11958);
and U12743 (N_12743,N_11903,N_11184);
or U12744 (N_12744,N_11544,N_11300);
and U12745 (N_12745,N_11490,N_11754);
xor U12746 (N_12746,N_11581,N_11095);
xor U12747 (N_12747,N_11449,N_11891);
nand U12748 (N_12748,N_11789,N_11612);
nor U12749 (N_12749,N_11035,N_11096);
nand U12750 (N_12750,N_11453,N_11277);
nor U12751 (N_12751,N_11306,N_10870);
nor U12752 (N_12752,N_11987,N_11992);
or U12753 (N_12753,N_11128,N_11154);
and U12754 (N_12754,N_11269,N_11587);
xnor U12755 (N_12755,N_10855,N_11450);
nor U12756 (N_12756,N_11642,N_11501);
xnor U12757 (N_12757,N_11545,N_11345);
nand U12758 (N_12758,N_11722,N_11637);
and U12759 (N_12759,N_11583,N_11651);
nor U12760 (N_12760,N_11808,N_10938);
xor U12761 (N_12761,N_10838,N_11946);
nor U12762 (N_12762,N_10907,N_10875);
nor U12763 (N_12763,N_11568,N_11133);
xor U12764 (N_12764,N_11639,N_11919);
xor U12765 (N_12765,N_11622,N_11261);
and U12766 (N_12766,N_11973,N_11453);
and U12767 (N_12767,N_11161,N_10861);
or U12768 (N_12768,N_11522,N_11928);
or U12769 (N_12769,N_11661,N_10941);
and U12770 (N_12770,N_11750,N_11438);
nor U12771 (N_12771,N_10909,N_11882);
and U12772 (N_12772,N_11501,N_11585);
xnor U12773 (N_12773,N_11688,N_11927);
xnor U12774 (N_12774,N_11723,N_11763);
nand U12775 (N_12775,N_11694,N_11902);
nand U12776 (N_12776,N_11356,N_11825);
xnor U12777 (N_12777,N_11585,N_11518);
nor U12778 (N_12778,N_11052,N_11069);
nand U12779 (N_12779,N_11162,N_11240);
xnor U12780 (N_12780,N_11046,N_11871);
nand U12781 (N_12781,N_11868,N_11155);
xnor U12782 (N_12782,N_11528,N_10858);
and U12783 (N_12783,N_11507,N_11782);
or U12784 (N_12784,N_11232,N_11143);
xnor U12785 (N_12785,N_11740,N_11593);
and U12786 (N_12786,N_11768,N_11107);
or U12787 (N_12787,N_11375,N_10956);
xor U12788 (N_12788,N_11558,N_11343);
and U12789 (N_12789,N_11037,N_10902);
nand U12790 (N_12790,N_11448,N_11628);
or U12791 (N_12791,N_11676,N_10812);
or U12792 (N_12792,N_11456,N_10967);
xnor U12793 (N_12793,N_11903,N_11634);
xnor U12794 (N_12794,N_11509,N_10929);
nor U12795 (N_12795,N_11402,N_11924);
xnor U12796 (N_12796,N_11091,N_11125);
and U12797 (N_12797,N_11713,N_11708);
nand U12798 (N_12798,N_10832,N_11112);
xor U12799 (N_12799,N_11475,N_11961);
xnor U12800 (N_12800,N_10959,N_10992);
or U12801 (N_12801,N_10910,N_10890);
nor U12802 (N_12802,N_11423,N_10927);
and U12803 (N_12803,N_10840,N_11440);
or U12804 (N_12804,N_11625,N_11388);
xnor U12805 (N_12805,N_11726,N_10958);
and U12806 (N_12806,N_11509,N_10871);
xnor U12807 (N_12807,N_11111,N_11727);
nand U12808 (N_12808,N_10974,N_10980);
nor U12809 (N_12809,N_10964,N_11970);
and U12810 (N_12810,N_11862,N_11291);
nand U12811 (N_12811,N_11595,N_11646);
or U12812 (N_12812,N_11145,N_11103);
xnor U12813 (N_12813,N_11524,N_11454);
nor U12814 (N_12814,N_10922,N_11671);
nor U12815 (N_12815,N_11468,N_11751);
nand U12816 (N_12816,N_11813,N_11329);
and U12817 (N_12817,N_11299,N_11634);
nand U12818 (N_12818,N_11067,N_11394);
or U12819 (N_12819,N_11897,N_10869);
nand U12820 (N_12820,N_11072,N_11157);
and U12821 (N_12821,N_11754,N_10971);
and U12822 (N_12822,N_10935,N_10930);
nand U12823 (N_12823,N_11216,N_11647);
or U12824 (N_12824,N_11206,N_11077);
nand U12825 (N_12825,N_11776,N_11924);
xnor U12826 (N_12826,N_11515,N_11407);
xor U12827 (N_12827,N_11502,N_11256);
nand U12828 (N_12828,N_11549,N_11718);
and U12829 (N_12829,N_11869,N_10888);
xnor U12830 (N_12830,N_11396,N_11389);
xnor U12831 (N_12831,N_11853,N_11658);
nor U12832 (N_12832,N_11267,N_11206);
and U12833 (N_12833,N_10937,N_11149);
nand U12834 (N_12834,N_11811,N_11114);
nor U12835 (N_12835,N_11022,N_11447);
nor U12836 (N_12836,N_11814,N_11437);
and U12837 (N_12837,N_11337,N_11610);
nor U12838 (N_12838,N_11363,N_11740);
nor U12839 (N_12839,N_11740,N_11132);
and U12840 (N_12840,N_10883,N_10943);
and U12841 (N_12841,N_11511,N_11673);
or U12842 (N_12842,N_11305,N_11721);
or U12843 (N_12843,N_11749,N_11879);
or U12844 (N_12844,N_11107,N_11842);
xor U12845 (N_12845,N_11250,N_10845);
nand U12846 (N_12846,N_11562,N_10800);
or U12847 (N_12847,N_11330,N_11052);
xor U12848 (N_12848,N_11021,N_11657);
or U12849 (N_12849,N_11295,N_11109);
xor U12850 (N_12850,N_11951,N_11430);
nor U12851 (N_12851,N_11052,N_11904);
nor U12852 (N_12852,N_11652,N_10900);
nand U12853 (N_12853,N_11894,N_11976);
or U12854 (N_12854,N_11459,N_11819);
nor U12855 (N_12855,N_11813,N_11061);
or U12856 (N_12856,N_11465,N_11384);
and U12857 (N_12857,N_11778,N_11702);
nor U12858 (N_12858,N_10891,N_11461);
or U12859 (N_12859,N_11187,N_11199);
or U12860 (N_12860,N_11968,N_11397);
or U12861 (N_12861,N_11996,N_11386);
and U12862 (N_12862,N_11066,N_11665);
nor U12863 (N_12863,N_11325,N_11785);
nand U12864 (N_12864,N_11361,N_11912);
and U12865 (N_12865,N_11661,N_11424);
nor U12866 (N_12866,N_11180,N_11946);
nor U12867 (N_12867,N_11233,N_11528);
and U12868 (N_12868,N_11144,N_11063);
and U12869 (N_12869,N_10931,N_11933);
and U12870 (N_12870,N_11752,N_11785);
xnor U12871 (N_12871,N_11542,N_11006);
nor U12872 (N_12872,N_10814,N_11041);
or U12873 (N_12873,N_11611,N_11776);
and U12874 (N_12874,N_11925,N_11097);
xor U12875 (N_12875,N_11953,N_11149);
xor U12876 (N_12876,N_11855,N_11759);
or U12877 (N_12877,N_11243,N_11771);
and U12878 (N_12878,N_11757,N_11514);
or U12879 (N_12879,N_11810,N_11398);
or U12880 (N_12880,N_11158,N_11033);
or U12881 (N_12881,N_11960,N_11948);
nor U12882 (N_12882,N_11381,N_11189);
xnor U12883 (N_12883,N_11333,N_11309);
nor U12884 (N_12884,N_11080,N_11013);
and U12885 (N_12885,N_10903,N_11392);
xnor U12886 (N_12886,N_11095,N_11483);
nor U12887 (N_12887,N_11220,N_11061);
and U12888 (N_12888,N_11667,N_11806);
xnor U12889 (N_12889,N_11170,N_11932);
and U12890 (N_12890,N_10948,N_11019);
or U12891 (N_12891,N_11919,N_11150);
or U12892 (N_12892,N_11339,N_11107);
nor U12893 (N_12893,N_11459,N_11581);
nand U12894 (N_12894,N_11941,N_11676);
nand U12895 (N_12895,N_11523,N_11851);
xor U12896 (N_12896,N_11054,N_11587);
nand U12897 (N_12897,N_10956,N_11577);
nor U12898 (N_12898,N_11887,N_11904);
xor U12899 (N_12899,N_11946,N_11900);
nand U12900 (N_12900,N_11365,N_11284);
nand U12901 (N_12901,N_11192,N_11950);
xor U12902 (N_12902,N_11078,N_10892);
xor U12903 (N_12903,N_11223,N_11874);
xnor U12904 (N_12904,N_11193,N_11345);
nor U12905 (N_12905,N_10924,N_11184);
or U12906 (N_12906,N_11734,N_11852);
nor U12907 (N_12907,N_11156,N_11230);
nand U12908 (N_12908,N_11277,N_10853);
or U12909 (N_12909,N_11133,N_10891);
nor U12910 (N_12910,N_10896,N_11155);
nor U12911 (N_12911,N_10976,N_10979);
nor U12912 (N_12912,N_11863,N_11632);
nor U12913 (N_12913,N_10881,N_11811);
and U12914 (N_12914,N_11629,N_11067);
nand U12915 (N_12915,N_11241,N_10905);
and U12916 (N_12916,N_11110,N_11951);
xnor U12917 (N_12917,N_11097,N_11483);
xnor U12918 (N_12918,N_11949,N_11381);
nand U12919 (N_12919,N_11518,N_11176);
and U12920 (N_12920,N_11519,N_11936);
and U12921 (N_12921,N_11351,N_11420);
or U12922 (N_12922,N_10985,N_11327);
nand U12923 (N_12923,N_11262,N_11809);
nand U12924 (N_12924,N_11805,N_11125);
xnor U12925 (N_12925,N_11860,N_11918);
xor U12926 (N_12926,N_11357,N_11757);
and U12927 (N_12927,N_11405,N_10995);
or U12928 (N_12928,N_11380,N_10807);
nand U12929 (N_12929,N_10930,N_11966);
xnor U12930 (N_12930,N_11469,N_11843);
and U12931 (N_12931,N_11206,N_11070);
nand U12932 (N_12932,N_10919,N_11241);
xor U12933 (N_12933,N_11343,N_11676);
and U12934 (N_12934,N_11642,N_11403);
nand U12935 (N_12935,N_11009,N_11550);
nor U12936 (N_12936,N_11507,N_11264);
nand U12937 (N_12937,N_11747,N_11894);
nand U12938 (N_12938,N_11446,N_11057);
nand U12939 (N_12939,N_11017,N_11524);
xnor U12940 (N_12940,N_11138,N_11384);
nand U12941 (N_12941,N_11180,N_11740);
xnor U12942 (N_12942,N_11281,N_10814);
nor U12943 (N_12943,N_10927,N_10862);
and U12944 (N_12944,N_11442,N_11551);
or U12945 (N_12945,N_11034,N_11025);
or U12946 (N_12946,N_11930,N_11075);
nor U12947 (N_12947,N_11624,N_10923);
xor U12948 (N_12948,N_11189,N_11770);
and U12949 (N_12949,N_10805,N_11591);
xnor U12950 (N_12950,N_11957,N_11294);
and U12951 (N_12951,N_11716,N_11684);
nand U12952 (N_12952,N_11758,N_11778);
xor U12953 (N_12953,N_11255,N_11525);
xnor U12954 (N_12954,N_11380,N_11373);
xnor U12955 (N_12955,N_11491,N_11110);
nor U12956 (N_12956,N_11941,N_11890);
nor U12957 (N_12957,N_11759,N_11715);
nand U12958 (N_12958,N_11205,N_11607);
nand U12959 (N_12959,N_11328,N_11667);
nand U12960 (N_12960,N_10874,N_11818);
nor U12961 (N_12961,N_10988,N_11186);
xnor U12962 (N_12962,N_11560,N_11430);
nor U12963 (N_12963,N_11660,N_11129);
nor U12964 (N_12964,N_11562,N_11901);
xor U12965 (N_12965,N_11630,N_11141);
nand U12966 (N_12966,N_11164,N_11222);
and U12967 (N_12967,N_11772,N_11168);
xnor U12968 (N_12968,N_10943,N_11692);
xnor U12969 (N_12969,N_11493,N_11452);
nor U12970 (N_12970,N_11059,N_11887);
or U12971 (N_12971,N_10954,N_10830);
xnor U12972 (N_12972,N_11219,N_11044);
nor U12973 (N_12973,N_10955,N_11770);
nand U12974 (N_12974,N_11685,N_11841);
xnor U12975 (N_12975,N_11211,N_11353);
or U12976 (N_12976,N_10830,N_11250);
nor U12977 (N_12977,N_11604,N_11070);
or U12978 (N_12978,N_10990,N_11579);
xnor U12979 (N_12979,N_11219,N_11833);
nand U12980 (N_12980,N_11257,N_11047);
or U12981 (N_12981,N_11979,N_11562);
and U12982 (N_12982,N_11881,N_11195);
or U12983 (N_12983,N_11522,N_11060);
nand U12984 (N_12984,N_11398,N_11074);
xor U12985 (N_12985,N_11228,N_11896);
nand U12986 (N_12986,N_11666,N_11547);
xnor U12987 (N_12987,N_11552,N_11786);
and U12988 (N_12988,N_10800,N_11645);
nor U12989 (N_12989,N_11352,N_10942);
nand U12990 (N_12990,N_11408,N_11443);
or U12991 (N_12991,N_11534,N_11522);
nand U12992 (N_12992,N_11934,N_11908);
and U12993 (N_12993,N_11261,N_11919);
nor U12994 (N_12994,N_11514,N_11171);
xor U12995 (N_12995,N_10827,N_11434);
nand U12996 (N_12996,N_11148,N_11145);
nor U12997 (N_12997,N_11842,N_11248);
or U12998 (N_12998,N_11141,N_11772);
xnor U12999 (N_12999,N_11694,N_11831);
and U13000 (N_13000,N_11083,N_11673);
nor U13001 (N_13001,N_11002,N_11925);
nand U13002 (N_13002,N_11695,N_10819);
xnor U13003 (N_13003,N_11414,N_11534);
or U13004 (N_13004,N_11403,N_11896);
nor U13005 (N_13005,N_11312,N_11196);
xnor U13006 (N_13006,N_10880,N_10888);
xnor U13007 (N_13007,N_11422,N_11067);
or U13008 (N_13008,N_11477,N_11130);
or U13009 (N_13009,N_11577,N_11695);
and U13010 (N_13010,N_11514,N_10851);
or U13011 (N_13011,N_11787,N_11950);
xor U13012 (N_13012,N_11587,N_11336);
nand U13013 (N_13013,N_11791,N_11581);
nor U13014 (N_13014,N_11779,N_11900);
and U13015 (N_13015,N_11434,N_10954);
and U13016 (N_13016,N_11699,N_11038);
xor U13017 (N_13017,N_10985,N_11033);
nor U13018 (N_13018,N_11024,N_11163);
nand U13019 (N_13019,N_11977,N_11307);
nand U13020 (N_13020,N_11222,N_11302);
and U13021 (N_13021,N_11763,N_11422);
or U13022 (N_13022,N_11990,N_11582);
xor U13023 (N_13023,N_11482,N_11809);
nor U13024 (N_13024,N_11655,N_11431);
or U13025 (N_13025,N_11813,N_11018);
nand U13026 (N_13026,N_11934,N_11501);
or U13027 (N_13027,N_11698,N_11937);
or U13028 (N_13028,N_10923,N_11155);
and U13029 (N_13029,N_11404,N_11034);
nand U13030 (N_13030,N_11434,N_10978);
and U13031 (N_13031,N_10990,N_10985);
nor U13032 (N_13032,N_11589,N_11856);
nand U13033 (N_13033,N_11738,N_10809);
xor U13034 (N_13034,N_11631,N_10849);
xnor U13035 (N_13035,N_11143,N_11396);
or U13036 (N_13036,N_11001,N_11822);
nor U13037 (N_13037,N_11841,N_10996);
nor U13038 (N_13038,N_11477,N_11678);
and U13039 (N_13039,N_11247,N_11929);
and U13040 (N_13040,N_11761,N_11465);
nor U13041 (N_13041,N_11444,N_11165);
nand U13042 (N_13042,N_11170,N_11630);
xor U13043 (N_13043,N_11284,N_11638);
nand U13044 (N_13044,N_11309,N_10813);
xor U13045 (N_13045,N_11102,N_11318);
xor U13046 (N_13046,N_11973,N_10982);
or U13047 (N_13047,N_11987,N_11588);
and U13048 (N_13048,N_10960,N_11931);
nor U13049 (N_13049,N_11516,N_11714);
and U13050 (N_13050,N_11631,N_11490);
or U13051 (N_13051,N_11787,N_11323);
xor U13052 (N_13052,N_11156,N_11177);
xnor U13053 (N_13053,N_11836,N_11993);
nor U13054 (N_13054,N_11671,N_11775);
or U13055 (N_13055,N_11587,N_11297);
or U13056 (N_13056,N_11599,N_10918);
nor U13057 (N_13057,N_11777,N_11651);
or U13058 (N_13058,N_11638,N_11287);
nor U13059 (N_13059,N_11921,N_10871);
and U13060 (N_13060,N_11091,N_11476);
nor U13061 (N_13061,N_11683,N_11711);
xor U13062 (N_13062,N_11960,N_11489);
nor U13063 (N_13063,N_10898,N_11613);
nor U13064 (N_13064,N_10988,N_11658);
and U13065 (N_13065,N_11440,N_10958);
nand U13066 (N_13066,N_11732,N_11566);
nand U13067 (N_13067,N_11284,N_11933);
or U13068 (N_13068,N_11547,N_11901);
nor U13069 (N_13069,N_11092,N_10801);
and U13070 (N_13070,N_11508,N_11507);
nor U13071 (N_13071,N_11868,N_11091);
and U13072 (N_13072,N_11071,N_11811);
nand U13073 (N_13073,N_11652,N_11859);
and U13074 (N_13074,N_11012,N_11476);
or U13075 (N_13075,N_11933,N_11899);
xnor U13076 (N_13076,N_10810,N_11428);
nor U13077 (N_13077,N_11517,N_11212);
nand U13078 (N_13078,N_11261,N_11993);
nor U13079 (N_13079,N_11383,N_11710);
xnor U13080 (N_13080,N_11955,N_10814);
or U13081 (N_13081,N_11327,N_11781);
and U13082 (N_13082,N_10969,N_11342);
and U13083 (N_13083,N_11228,N_11821);
nor U13084 (N_13084,N_10831,N_11788);
xor U13085 (N_13085,N_11963,N_11046);
and U13086 (N_13086,N_11656,N_11111);
and U13087 (N_13087,N_10828,N_10856);
or U13088 (N_13088,N_11874,N_11845);
nor U13089 (N_13089,N_11256,N_11489);
nand U13090 (N_13090,N_11377,N_11008);
and U13091 (N_13091,N_10840,N_11514);
or U13092 (N_13092,N_11363,N_10894);
or U13093 (N_13093,N_11679,N_11526);
and U13094 (N_13094,N_11724,N_11603);
nor U13095 (N_13095,N_11480,N_11883);
nor U13096 (N_13096,N_11617,N_11730);
nand U13097 (N_13097,N_11985,N_10947);
and U13098 (N_13098,N_11598,N_11586);
and U13099 (N_13099,N_11621,N_11235);
and U13100 (N_13100,N_11317,N_11787);
nor U13101 (N_13101,N_11390,N_10898);
xnor U13102 (N_13102,N_10983,N_11669);
nand U13103 (N_13103,N_11838,N_11273);
nand U13104 (N_13104,N_11813,N_11023);
nand U13105 (N_13105,N_10876,N_11226);
and U13106 (N_13106,N_11317,N_11698);
nand U13107 (N_13107,N_10841,N_10803);
nor U13108 (N_13108,N_11921,N_11272);
and U13109 (N_13109,N_11451,N_11090);
or U13110 (N_13110,N_10832,N_11131);
xor U13111 (N_13111,N_11978,N_11930);
or U13112 (N_13112,N_11496,N_11914);
nand U13113 (N_13113,N_11861,N_11063);
nor U13114 (N_13114,N_10920,N_11116);
nand U13115 (N_13115,N_11496,N_11387);
or U13116 (N_13116,N_11243,N_11689);
and U13117 (N_13117,N_11844,N_11322);
and U13118 (N_13118,N_11487,N_11803);
or U13119 (N_13119,N_11200,N_11731);
nor U13120 (N_13120,N_10901,N_11338);
or U13121 (N_13121,N_11733,N_11398);
and U13122 (N_13122,N_10899,N_11417);
xor U13123 (N_13123,N_11841,N_11715);
nand U13124 (N_13124,N_11550,N_11908);
and U13125 (N_13125,N_11720,N_11255);
nand U13126 (N_13126,N_11644,N_11997);
or U13127 (N_13127,N_11827,N_11857);
or U13128 (N_13128,N_11012,N_11826);
nand U13129 (N_13129,N_11675,N_10855);
nor U13130 (N_13130,N_11151,N_11240);
nor U13131 (N_13131,N_11524,N_10881);
and U13132 (N_13132,N_11416,N_11281);
nand U13133 (N_13133,N_11426,N_11220);
nor U13134 (N_13134,N_11964,N_11510);
nand U13135 (N_13135,N_11946,N_11499);
xnor U13136 (N_13136,N_11741,N_11935);
or U13137 (N_13137,N_10976,N_11671);
or U13138 (N_13138,N_11072,N_11330);
nor U13139 (N_13139,N_11144,N_11196);
xor U13140 (N_13140,N_10851,N_11405);
nor U13141 (N_13141,N_11580,N_10833);
and U13142 (N_13142,N_11675,N_11008);
nand U13143 (N_13143,N_10919,N_11253);
nand U13144 (N_13144,N_11338,N_11221);
and U13145 (N_13145,N_10846,N_11850);
and U13146 (N_13146,N_10844,N_11434);
nand U13147 (N_13147,N_11590,N_10851);
nor U13148 (N_13148,N_11267,N_11713);
xnor U13149 (N_13149,N_11930,N_11253);
nor U13150 (N_13150,N_11585,N_10997);
nand U13151 (N_13151,N_11433,N_11235);
nand U13152 (N_13152,N_11710,N_11762);
or U13153 (N_13153,N_10900,N_11524);
xor U13154 (N_13154,N_11838,N_11610);
xnor U13155 (N_13155,N_11303,N_11352);
xor U13156 (N_13156,N_11208,N_10820);
xor U13157 (N_13157,N_11301,N_11931);
nand U13158 (N_13158,N_11308,N_11640);
xor U13159 (N_13159,N_11959,N_11168);
or U13160 (N_13160,N_10906,N_11999);
xor U13161 (N_13161,N_11401,N_11403);
and U13162 (N_13162,N_11146,N_11914);
nor U13163 (N_13163,N_11455,N_11910);
xnor U13164 (N_13164,N_10825,N_11106);
and U13165 (N_13165,N_11793,N_11783);
xnor U13166 (N_13166,N_11025,N_11365);
or U13167 (N_13167,N_11052,N_11609);
nor U13168 (N_13168,N_11808,N_10813);
nand U13169 (N_13169,N_10886,N_10915);
or U13170 (N_13170,N_11497,N_11275);
and U13171 (N_13171,N_11493,N_11171);
and U13172 (N_13172,N_11424,N_10850);
and U13173 (N_13173,N_11496,N_10983);
or U13174 (N_13174,N_11345,N_11913);
nand U13175 (N_13175,N_11527,N_11528);
nor U13176 (N_13176,N_11962,N_11594);
nand U13177 (N_13177,N_11969,N_11118);
nor U13178 (N_13178,N_11897,N_11703);
xor U13179 (N_13179,N_11235,N_11715);
nor U13180 (N_13180,N_11631,N_11903);
or U13181 (N_13181,N_11551,N_11990);
and U13182 (N_13182,N_10910,N_11734);
nor U13183 (N_13183,N_11963,N_11891);
and U13184 (N_13184,N_11420,N_10989);
nand U13185 (N_13185,N_11480,N_11904);
or U13186 (N_13186,N_10803,N_10840);
xnor U13187 (N_13187,N_11087,N_10812);
xor U13188 (N_13188,N_11779,N_11103);
or U13189 (N_13189,N_11561,N_11385);
nand U13190 (N_13190,N_11458,N_11413);
nor U13191 (N_13191,N_11649,N_11735);
and U13192 (N_13192,N_11755,N_11192);
nor U13193 (N_13193,N_11513,N_11173);
or U13194 (N_13194,N_11460,N_11381);
nand U13195 (N_13195,N_11084,N_11745);
xnor U13196 (N_13196,N_11258,N_11793);
nor U13197 (N_13197,N_11590,N_11863);
or U13198 (N_13198,N_11893,N_11973);
nand U13199 (N_13199,N_10873,N_11219);
and U13200 (N_13200,N_12522,N_12970);
nand U13201 (N_13201,N_12633,N_12246);
nor U13202 (N_13202,N_12704,N_12049);
nand U13203 (N_13203,N_13115,N_12496);
xnor U13204 (N_13204,N_12197,N_12994);
xnor U13205 (N_13205,N_12059,N_12206);
nand U13206 (N_13206,N_13095,N_12914);
xor U13207 (N_13207,N_12763,N_13041);
or U13208 (N_13208,N_12601,N_13002);
nor U13209 (N_13209,N_12649,N_13110);
and U13210 (N_13210,N_13026,N_12379);
or U13211 (N_13211,N_12116,N_12533);
xnor U13212 (N_13212,N_12671,N_13035);
and U13213 (N_13213,N_12385,N_12882);
nor U13214 (N_13214,N_12057,N_12226);
and U13215 (N_13215,N_12802,N_12983);
and U13216 (N_13216,N_12129,N_12718);
or U13217 (N_13217,N_12073,N_12563);
nand U13218 (N_13218,N_12909,N_12866);
and U13219 (N_13219,N_12363,N_12894);
nand U13220 (N_13220,N_13032,N_12027);
nor U13221 (N_13221,N_12176,N_12456);
nand U13222 (N_13222,N_12334,N_12175);
nor U13223 (N_13223,N_12958,N_12579);
and U13224 (N_13224,N_12873,N_12191);
nand U13225 (N_13225,N_12449,N_12309);
nand U13226 (N_13226,N_12636,N_13129);
nand U13227 (N_13227,N_12901,N_12090);
xnor U13228 (N_13228,N_12665,N_12227);
and U13229 (N_13229,N_12211,N_12719);
xor U13230 (N_13230,N_12692,N_12731);
xor U13231 (N_13231,N_12588,N_12083);
or U13232 (N_13232,N_13088,N_13163);
xnor U13233 (N_13233,N_12183,N_12823);
nand U13234 (N_13234,N_12233,N_12615);
nand U13235 (N_13235,N_12479,N_12004);
nor U13236 (N_13236,N_12310,N_13057);
nor U13237 (N_13237,N_12408,N_13093);
xor U13238 (N_13238,N_13109,N_13187);
nand U13239 (N_13239,N_12820,N_12338);
nor U13240 (N_13240,N_12068,N_12656);
or U13241 (N_13241,N_12635,N_12199);
and U13242 (N_13242,N_13039,N_12593);
and U13243 (N_13243,N_12908,N_12660);
nor U13244 (N_13244,N_12691,N_12121);
nor U13245 (N_13245,N_12320,N_12487);
nand U13246 (N_13246,N_12913,N_12888);
xor U13247 (N_13247,N_13104,N_12626);
or U13248 (N_13248,N_12134,N_12260);
nand U13249 (N_13249,N_12082,N_12461);
and U13250 (N_13250,N_12741,N_12160);
nand U13251 (N_13251,N_12587,N_12344);
or U13252 (N_13252,N_13118,N_13178);
or U13253 (N_13253,N_12207,N_12637);
and U13254 (N_13254,N_12960,N_13033);
and U13255 (N_13255,N_12234,N_12333);
or U13256 (N_13256,N_12433,N_12232);
and U13257 (N_13257,N_12291,N_12289);
and U13258 (N_13258,N_12119,N_13185);
and U13259 (N_13259,N_12186,N_12341);
nor U13260 (N_13260,N_12854,N_12906);
nor U13261 (N_13261,N_13006,N_12013);
nor U13262 (N_13262,N_12431,N_12876);
or U13263 (N_13263,N_12747,N_12592);
and U13264 (N_13264,N_12219,N_12564);
nand U13265 (N_13265,N_12323,N_12076);
or U13266 (N_13266,N_12046,N_12272);
or U13267 (N_13267,N_12172,N_12971);
xnor U13268 (N_13268,N_12816,N_12865);
nor U13269 (N_13269,N_12951,N_13116);
nand U13270 (N_13270,N_13122,N_12541);
nand U13271 (N_13271,N_12628,N_12613);
and U13272 (N_13272,N_12723,N_13005);
or U13273 (N_13273,N_13100,N_12275);
and U13274 (N_13274,N_12304,N_12240);
or U13275 (N_13275,N_12209,N_12263);
and U13276 (N_13276,N_12806,N_12834);
nand U13277 (N_13277,N_12403,N_12441);
or U13278 (N_13278,N_12003,N_12221);
nor U13279 (N_13279,N_12993,N_13184);
or U13280 (N_13280,N_12895,N_12949);
nor U13281 (N_13281,N_12627,N_12482);
and U13282 (N_13282,N_12946,N_12915);
and U13283 (N_13283,N_12158,N_12911);
or U13284 (N_13284,N_12574,N_12437);
xnor U13285 (N_13285,N_13091,N_12887);
and U13286 (N_13286,N_12150,N_12714);
and U13287 (N_13287,N_12336,N_12361);
nand U13288 (N_13288,N_13176,N_12066);
nand U13289 (N_13289,N_12780,N_12390);
nand U13290 (N_13290,N_12167,N_12114);
xnor U13291 (N_13291,N_13136,N_12241);
nor U13292 (N_13292,N_12047,N_13098);
xor U13293 (N_13293,N_12280,N_12662);
and U13294 (N_13294,N_12043,N_12460);
nor U13295 (N_13295,N_13105,N_12427);
and U13296 (N_13296,N_12358,N_12113);
nand U13297 (N_13297,N_12598,N_12515);
nand U13298 (N_13298,N_12669,N_12445);
and U13299 (N_13299,N_12870,N_12781);
nor U13300 (N_13300,N_12130,N_12135);
or U13301 (N_13301,N_12967,N_12827);
or U13302 (N_13302,N_13013,N_12954);
or U13303 (N_13303,N_12836,N_12006);
xnor U13304 (N_13304,N_12265,N_12857);
or U13305 (N_13305,N_12596,N_12185);
nor U13306 (N_13306,N_13059,N_12282);
and U13307 (N_13307,N_12171,N_12026);
nor U13308 (N_13308,N_13103,N_12484);
nor U13309 (N_13309,N_12767,N_12143);
nor U13310 (N_13310,N_12752,N_12093);
and U13311 (N_13311,N_12629,N_12568);
nand U13312 (N_13312,N_12115,N_13055);
nand U13313 (N_13313,N_12110,N_12848);
and U13314 (N_13314,N_12589,N_12721);
and U13315 (N_13315,N_12516,N_13155);
or U13316 (N_13316,N_12506,N_12594);
nand U13317 (N_13317,N_12330,N_13124);
nand U13318 (N_13318,N_13101,N_12400);
nor U13319 (N_13319,N_12355,N_13111);
and U13320 (N_13320,N_12772,N_12939);
and U13321 (N_13321,N_12843,N_12771);
and U13322 (N_13322,N_12436,N_12773);
or U13323 (N_13323,N_12508,N_12012);
xor U13324 (N_13324,N_12672,N_12283);
nor U13325 (N_13325,N_12488,N_12092);
nand U13326 (N_13326,N_12060,N_12904);
or U13327 (N_13327,N_13191,N_12069);
nand U13328 (N_13328,N_12019,N_12632);
nand U13329 (N_13329,N_12389,N_12216);
and U13330 (N_13330,N_12335,N_12735);
nand U13331 (N_13331,N_13177,N_12397);
or U13332 (N_13332,N_13148,N_12395);
nand U13333 (N_13333,N_12828,N_12268);
xor U13334 (N_13334,N_12641,N_12029);
nor U13335 (N_13335,N_12365,N_12753);
and U13336 (N_13336,N_12862,N_12236);
and U13337 (N_13337,N_12063,N_12664);
nor U13338 (N_13338,N_12961,N_12988);
nand U13339 (N_13339,N_12301,N_12243);
and U13340 (N_13340,N_12750,N_12164);
nand U13341 (N_13341,N_12072,N_12572);
nand U13342 (N_13342,N_12803,N_13160);
nor U13343 (N_13343,N_12490,N_12276);
and U13344 (N_13344,N_13074,N_12965);
nand U13345 (N_13345,N_12536,N_12432);
and U13346 (N_13346,N_12010,N_13043);
or U13347 (N_13347,N_12316,N_12039);
or U13348 (N_13348,N_12108,N_12486);
xnor U13349 (N_13349,N_12077,N_12071);
or U13350 (N_13350,N_12535,N_13156);
or U13351 (N_13351,N_12148,N_12811);
nand U13352 (N_13352,N_12373,N_12132);
nand U13353 (N_13353,N_12789,N_12693);
and U13354 (N_13354,N_12737,N_12878);
nand U13355 (N_13355,N_12493,N_12896);
or U13356 (N_13356,N_12308,N_12253);
nor U13357 (N_13357,N_12776,N_12630);
nand U13358 (N_13358,N_13068,N_12331);
or U13359 (N_13359,N_12998,N_12306);
or U13360 (N_13360,N_13084,N_12530);
and U13361 (N_13361,N_12645,N_12852);
xor U13362 (N_13362,N_12791,N_12549);
or U13363 (N_13363,N_12290,N_12996);
or U13364 (N_13364,N_12087,N_12782);
and U13365 (N_13365,N_12005,N_12052);
or U13366 (N_13366,N_13120,N_12619);
nand U13367 (N_13367,N_12571,N_12466);
and U13368 (N_13368,N_13114,N_13186);
nand U13369 (N_13369,N_13189,N_13128);
or U13370 (N_13370,N_12295,N_12512);
or U13371 (N_13371,N_12975,N_12138);
nor U13372 (N_13372,N_12864,N_13142);
nor U13373 (N_13373,N_12284,N_12898);
nor U13374 (N_13374,N_12997,N_12473);
nor U13375 (N_13375,N_12956,N_12668);
nor U13376 (N_13376,N_12410,N_12399);
nand U13377 (N_13377,N_13011,N_12156);
or U13378 (N_13378,N_12703,N_12585);
or U13379 (N_13379,N_12281,N_12494);
nor U13380 (N_13380,N_12332,N_12278);
nand U13381 (N_13381,N_12794,N_12270);
nand U13382 (N_13382,N_12959,N_13135);
nor U13383 (N_13383,N_12770,N_12795);
nor U13384 (N_13384,N_12697,N_12980);
or U13385 (N_13385,N_12829,N_12418);
nand U13386 (N_13386,N_12044,N_12098);
and U13387 (N_13387,N_12603,N_12817);
nor U13388 (N_13388,N_12294,N_12972);
xnor U13389 (N_13389,N_13180,N_12107);
and U13390 (N_13390,N_12105,N_12855);
and U13391 (N_13391,N_12402,N_12384);
nand U13392 (N_13392,N_12326,N_12679);
nor U13393 (N_13393,N_12805,N_13067);
or U13394 (N_13394,N_12078,N_12774);
xnor U13395 (N_13395,N_13069,N_13017);
and U13396 (N_13396,N_13112,N_12483);
nor U13397 (N_13397,N_12061,N_13165);
nand U13398 (N_13398,N_12231,N_12392);
xor U13399 (N_13399,N_12351,N_12492);
xor U13400 (N_13400,N_13094,N_12863);
and U13401 (N_13401,N_12256,N_12599);
nor U13402 (N_13402,N_12678,N_12342);
or U13403 (N_13403,N_12801,N_12877);
nand U13404 (N_13404,N_12015,N_13194);
or U13405 (N_13405,N_12048,N_12126);
nor U13406 (N_13406,N_13150,N_12765);
xor U13407 (N_13407,N_12910,N_13056);
xor U13408 (N_13408,N_12080,N_12962);
nand U13409 (N_13409,N_12383,N_13126);
nand U13410 (N_13410,N_12065,N_12396);
and U13411 (N_13411,N_12182,N_12017);
xnor U13412 (N_13412,N_12872,N_12248);
nor U13413 (N_13413,N_12178,N_12354);
and U13414 (N_13414,N_12844,N_12976);
nand U13415 (N_13415,N_13117,N_12732);
nor U13416 (N_13416,N_12239,N_12931);
xor U13417 (N_13417,N_12722,N_12986);
and U13418 (N_13418,N_12858,N_12525);
xnor U13419 (N_13419,N_12454,N_12345);
and U13420 (N_13420,N_13016,N_12462);
or U13421 (N_13421,N_12147,N_12526);
nor U13422 (N_13422,N_13138,N_12458);
or U13423 (N_13423,N_12607,N_12471);
and U13424 (N_13424,N_12808,N_12886);
or U13425 (N_13425,N_12120,N_12101);
and U13426 (N_13426,N_13166,N_12343);
and U13427 (N_13427,N_12356,N_12685);
nand U13428 (N_13428,N_12899,N_13060);
or U13429 (N_13429,N_12277,N_12498);
and U13430 (N_13430,N_13137,N_12838);
or U13431 (N_13431,N_12037,N_12459);
nor U13432 (N_13432,N_13190,N_12028);
xor U13433 (N_13433,N_13167,N_12405);
xnor U13434 (N_13434,N_12969,N_12538);
xor U13435 (N_13435,N_12086,N_12597);
or U13436 (N_13436,N_12885,N_12810);
or U13437 (N_13437,N_13102,N_12742);
or U13438 (N_13438,N_12190,N_12329);
xnor U13439 (N_13439,N_12787,N_12469);
nor U13440 (N_13440,N_12935,N_12897);
xnor U13441 (N_13441,N_12404,N_12255);
or U13442 (N_13442,N_12495,N_13054);
nor U13443 (N_13443,N_13197,N_12944);
nand U13444 (N_13444,N_13097,N_12166);
xnor U13445 (N_13445,N_12875,N_12799);
or U13446 (N_13446,N_12040,N_12520);
nor U13447 (N_13447,N_12687,N_12035);
nor U13448 (N_13448,N_12930,N_12995);
and U13449 (N_13449,N_12020,N_12045);
nand U13450 (N_13450,N_12386,N_12507);
nand U13451 (N_13451,N_13121,N_12570);
or U13452 (N_13452,N_13050,N_12798);
and U13453 (N_13453,N_12837,N_12924);
nor U13454 (N_13454,N_12267,N_12936);
xnor U13455 (N_13455,N_13183,N_12624);
and U13456 (N_13456,N_12832,N_12740);
xnor U13457 (N_13457,N_12973,N_12502);
or U13458 (N_13458,N_12056,N_12686);
nor U13459 (N_13459,N_12409,N_12425);
xor U13460 (N_13460,N_12426,N_12033);
nand U13461 (N_13461,N_13099,N_12102);
or U13462 (N_13462,N_12450,N_12586);
or U13463 (N_13463,N_12874,N_12748);
nor U13464 (N_13464,N_12153,N_12238);
xnor U13465 (N_13465,N_13079,N_12476);
nor U13466 (N_13466,N_13038,N_13131);
nor U13467 (N_13467,N_12474,N_12809);
and U13468 (N_13468,N_13021,N_12123);
xnor U13469 (N_13469,N_12642,N_13080);
nor U13470 (N_13470,N_13020,N_12394);
xor U13471 (N_13471,N_13089,N_12067);
and U13472 (N_13472,N_12555,N_12955);
nand U13473 (N_13473,N_12084,N_12759);
xor U13474 (N_13474,N_12591,N_12764);
nor U13475 (N_13475,N_12407,N_12413);
and U13476 (N_13476,N_13072,N_12918);
or U13477 (N_13477,N_12677,N_12058);
nand U13478 (N_13478,N_12839,N_12938);
nor U13479 (N_13479,N_12707,N_13040);
or U13480 (N_13480,N_12485,N_12546);
nor U13481 (N_13481,N_12325,N_12111);
nand U13482 (N_13482,N_12145,N_12055);
nor U13483 (N_13483,N_13063,N_12783);
xnor U13484 (N_13484,N_12706,N_12177);
and U13485 (N_13485,N_12237,N_12831);
nand U13486 (N_13486,N_12726,N_12163);
nand U13487 (N_13487,N_12941,N_12725);
or U13488 (N_13488,N_12339,N_12419);
or U13489 (N_13489,N_12736,N_12000);
xnor U13490 (N_13490,N_12757,N_13092);
nor U13491 (N_13491,N_12165,N_12286);
and U13492 (N_13492,N_12311,N_12009);
xor U13493 (N_13493,N_13027,N_12879);
and U13494 (N_13494,N_12391,N_12968);
nor U13495 (N_13495,N_13065,N_12928);
xor U13496 (N_13496,N_12925,N_13139);
and U13497 (N_13497,N_13066,N_12435);
and U13498 (N_13498,N_12024,N_12375);
nor U13499 (N_13499,N_12513,N_13044);
xnor U13500 (N_13500,N_12372,N_12845);
or U13501 (N_13501,N_12274,N_12842);
xnor U13502 (N_13502,N_12204,N_13158);
xnor U13503 (N_13503,N_12923,N_12903);
nor U13504 (N_13504,N_12659,N_13173);
and U13505 (N_13505,N_12374,N_12919);
nor U13506 (N_13506,N_13076,N_12141);
xnor U13507 (N_13507,N_12117,N_12880);
nand U13508 (N_13508,N_12766,N_12529);
xor U13509 (N_13509,N_13087,N_13010);
and U13510 (N_13510,N_12985,N_13162);
nand U13511 (N_13511,N_12749,N_13046);
or U13512 (N_13512,N_12189,N_12205);
and U13513 (N_13513,N_12144,N_12595);
xnor U13514 (N_13514,N_12584,N_12245);
or U13515 (N_13515,N_13014,N_12658);
and U13516 (N_13516,N_12833,N_12524);
nor U13517 (N_13517,N_12269,N_12327);
nor U13518 (N_13518,N_13024,N_12464);
nor U13519 (N_13519,N_12540,N_12813);
or U13520 (N_13520,N_12319,N_12670);
nor U13521 (N_13521,N_12312,N_12523);
nor U13522 (N_13522,N_12159,N_12902);
and U13523 (N_13523,N_12088,N_12353);
and U13524 (N_13524,N_12360,N_12195);
or U13525 (N_13525,N_12651,N_12576);
xnor U13526 (N_13526,N_12881,N_12314);
nand U13527 (N_13527,N_12168,N_12511);
nand U13528 (N_13528,N_13003,N_12556);
xor U13529 (N_13529,N_13077,N_12042);
or U13530 (N_13530,N_12974,N_12840);
nor U13531 (N_13531,N_12643,N_12273);
nand U13532 (N_13532,N_12318,N_12822);
and U13533 (N_13533,N_12359,N_12539);
nand U13534 (N_13534,N_12640,N_12398);
nand U13535 (N_13535,N_12279,N_13127);
nand U13536 (N_13536,N_12032,N_12963);
xor U13537 (N_13537,N_12517,N_12094);
or U13538 (N_13538,N_12106,N_12545);
or U13539 (N_13539,N_12440,N_13049);
and U13540 (N_13540,N_12022,N_12883);
nor U13541 (N_13541,N_12202,N_12777);
xor U13542 (N_13542,N_12755,N_12259);
nand U13543 (N_13543,N_13012,N_13195);
nand U13544 (N_13544,N_13147,N_12821);
nand U13545 (N_13545,N_12444,N_12618);
xnor U13546 (N_13546,N_12324,N_12382);
xnor U13547 (N_13547,N_12451,N_12531);
xor U13548 (N_13548,N_12011,N_13085);
and U13549 (N_13549,N_12676,N_12152);
and U13550 (N_13550,N_12992,N_12646);
and U13551 (N_13551,N_12151,N_12537);
nor U13552 (N_13552,N_12711,N_12137);
xnor U13553 (N_13553,N_12868,N_12681);
xnor U13554 (N_13554,N_12743,N_12631);
nand U13555 (N_13555,N_13125,N_13051);
and U13556 (N_13556,N_12565,N_12447);
and U13557 (N_13557,N_12779,N_12023);
nand U13558 (N_13558,N_12554,N_12644);
xor U13559 (N_13559,N_12945,N_13034);
xor U13560 (N_13560,N_12684,N_12465);
nand U13561 (N_13561,N_13001,N_12254);
nand U13562 (N_13562,N_12733,N_13108);
xor U13563 (N_13563,N_12169,N_12491);
xnor U13564 (N_13564,N_12021,N_12620);
nor U13565 (N_13565,N_12103,N_12869);
nor U13566 (N_13566,N_12322,N_13198);
xor U13567 (N_13567,N_12380,N_12340);
nor U13568 (N_13568,N_12235,N_13154);
and U13569 (N_13569,N_12756,N_13090);
nand U13570 (N_13570,N_12184,N_13151);
nand U13571 (N_13571,N_12991,N_12463);
nand U13572 (N_13572,N_12608,N_12890);
xor U13573 (N_13573,N_12790,N_12667);
nand U13574 (N_13574,N_12412,N_13113);
nor U13575 (N_13575,N_12299,N_12188);
or U13576 (N_13576,N_12952,N_12990);
or U13577 (N_13577,N_12746,N_12504);
or U13578 (N_13578,N_12406,N_12503);
nand U13579 (N_13579,N_12162,N_12715);
or U13580 (N_13580,N_12792,N_12287);
nor U13581 (N_13581,N_12293,N_12079);
nand U13582 (N_13582,N_12814,N_12125);
xor U13583 (N_13583,N_13053,N_12943);
and U13584 (N_13584,N_13004,N_12720);
xor U13585 (N_13585,N_12214,N_12929);
nand U13586 (N_13586,N_12109,N_12713);
xnor U13587 (N_13587,N_12758,N_12155);
nand U13588 (N_13588,N_12519,N_12567);
xor U13589 (N_13589,N_12179,N_12621);
nand U13590 (N_13590,N_12610,N_12984);
xor U13591 (N_13591,N_12414,N_13081);
or U13592 (N_13592,N_13052,N_12786);
nand U13593 (N_13593,N_12442,N_12142);
xnor U13594 (N_13594,N_13061,N_12217);
or U13595 (N_13595,N_12215,N_12112);
and U13596 (N_13596,N_12835,N_12614);
or U13597 (N_13597,N_12096,N_12860);
or U13598 (N_13598,N_12377,N_12018);
nor U13599 (N_13599,N_12518,N_13036);
and U13600 (N_13600,N_12648,N_13082);
or U13601 (N_13601,N_12244,N_12229);
and U13602 (N_13602,N_12266,N_12070);
and U13603 (N_13603,N_12712,N_12210);
xor U13604 (N_13604,N_12551,N_13164);
xnor U13605 (N_13605,N_12007,N_12446);
nand U13606 (N_13606,N_12443,N_12934);
xor U13607 (N_13607,N_12455,N_13146);
or U13608 (N_13608,N_12738,N_12761);
and U13609 (N_13609,N_12303,N_12258);
nor U13610 (N_13610,N_12977,N_12578);
or U13611 (N_13611,N_12001,N_12604);
nand U13612 (N_13612,N_12652,N_12501);
or U13613 (N_13613,N_12292,N_12905);
and U13614 (N_13614,N_12136,N_12016);
nor U13615 (N_13615,N_12422,N_12247);
nor U13616 (N_13616,N_13132,N_13083);
or U13617 (N_13617,N_12193,N_12600);
and U13618 (N_13618,N_13071,N_12218);
xor U13619 (N_13619,N_12388,N_12700);
and U13620 (N_13620,N_12804,N_12785);
nand U13621 (N_13621,N_12543,N_13073);
xor U13622 (N_13622,N_13019,N_12118);
nand U13623 (N_13623,N_12989,N_12769);
nand U13624 (N_13624,N_13106,N_12370);
nand U13625 (N_13625,N_12611,N_12940);
xnor U13626 (N_13626,N_12580,N_12417);
or U13627 (N_13627,N_12367,N_12349);
xnor U13628 (N_13628,N_13009,N_12054);
and U13629 (N_13629,N_12411,N_12133);
and U13630 (N_13630,N_12213,N_12357);
or U13631 (N_13631,N_12784,N_12228);
nor U13632 (N_13632,N_12192,N_12350);
xor U13633 (N_13633,N_12696,N_12085);
or U13634 (N_13634,N_12302,N_12583);
nand U13635 (N_13635,N_12760,N_12477);
nand U13636 (N_13636,N_13141,N_12249);
xor U13637 (N_13637,N_12364,N_12856);
nand U13638 (N_13638,N_12500,N_12230);
nor U13639 (N_13639,N_13029,N_12739);
xor U13640 (N_13640,N_12481,N_12181);
nand U13641 (N_13641,N_12051,N_12553);
and U13642 (N_13642,N_13152,N_13174);
nand U13643 (N_13643,N_12730,N_12734);
xor U13644 (N_13644,N_12926,N_12846);
or U13645 (N_13645,N_12222,N_12139);
nor U13646 (N_13646,N_12104,N_12573);
and U13647 (N_13647,N_12457,N_12321);
nand U13648 (N_13648,N_12666,N_12489);
xnor U13649 (N_13649,N_13175,N_12062);
nor U13650 (N_13650,N_12650,N_12948);
or U13651 (N_13651,N_13144,N_13133);
nor U13652 (N_13652,N_12438,N_12499);
nor U13653 (N_13653,N_12220,N_12612);
nand U13654 (N_13654,N_13179,N_12428);
and U13655 (N_13655,N_12429,N_12089);
nand U13656 (N_13656,N_12434,N_12699);
and U13657 (N_13657,N_12964,N_13123);
or U13658 (N_13658,N_12025,N_12654);
xnor U13659 (N_13659,N_13025,N_12548);
and U13660 (N_13660,N_12819,N_12871);
or U13661 (N_13661,N_12053,N_12724);
nor U13662 (N_13662,N_12912,N_12050);
xor U13663 (N_13663,N_12867,N_12097);
nand U13664 (N_13664,N_12847,N_12581);
or U13665 (N_13665,N_12602,N_12250);
and U13666 (N_13666,N_12544,N_12127);
and U13667 (N_13667,N_12550,N_13107);
xor U13668 (N_13668,N_12122,N_12609);
or U13669 (N_13669,N_12762,N_12682);
nor U13670 (N_13670,N_12953,N_12744);
and U13671 (N_13671,N_12095,N_13018);
or U13672 (N_13672,N_12528,N_12448);
and U13673 (N_13673,N_12099,N_12307);
nor U13674 (N_13674,N_12675,N_12261);
nand U13675 (N_13675,N_12634,N_12884);
and U13676 (N_13676,N_12657,N_13000);
and U13677 (N_13677,N_13182,N_12688);
or U13678 (N_13678,N_12701,N_12198);
nor U13679 (N_13679,N_12557,N_13078);
xor U13680 (N_13680,N_12947,N_12663);
or U13681 (N_13681,N_12393,N_12173);
nand U13682 (N_13682,N_12942,N_12212);
or U13683 (N_13683,N_12982,N_12423);
nor U13684 (N_13684,N_13042,N_12074);
xnor U13685 (N_13685,N_12566,N_13145);
nand U13686 (N_13686,N_13171,N_12534);
nor U13687 (N_13687,N_12690,N_12366);
nand U13688 (N_13688,N_12745,N_12920);
nand U13689 (N_13689,N_12552,N_12187);
and U13690 (N_13690,N_12807,N_12348);
or U13691 (N_13691,N_12625,N_12014);
xnor U13692 (N_13692,N_12369,N_12937);
and U13693 (N_13693,N_12420,N_12709);
or U13694 (N_13694,N_12547,N_12978);
and U13695 (N_13695,N_13140,N_12710);
nand U13696 (N_13696,N_12146,N_12100);
nor U13697 (N_13697,N_12957,N_13169);
and U13698 (N_13698,N_12716,N_12661);
or U13699 (N_13699,N_12922,N_12981);
xnor U13700 (N_13700,N_12775,N_12788);
or U13701 (N_13701,N_12157,N_12416);
or U13702 (N_13702,N_13037,N_13143);
nor U13703 (N_13703,N_12623,N_12337);
and U13704 (N_13704,N_12560,N_12475);
or U13705 (N_13705,N_13062,N_12683);
xnor U13706 (N_13706,N_13047,N_12297);
nor U13707 (N_13707,N_12346,N_12196);
nor U13708 (N_13708,N_12892,N_12590);
nand U13709 (N_13709,N_12917,N_12900);
xnor U13710 (N_13710,N_12315,N_13022);
and U13711 (N_13711,N_12242,N_12562);
nand U13712 (N_13712,N_12036,N_12264);
or U13713 (N_13713,N_12430,N_12861);
and U13714 (N_13714,N_12893,N_12569);
nand U13715 (N_13715,N_12616,N_12708);
and U13716 (N_13716,N_12850,N_12223);
nor U13717 (N_13717,N_12439,N_12031);
or U13718 (N_13718,N_12932,N_12296);
and U13719 (N_13719,N_13119,N_12124);
nand U13720 (N_13720,N_13023,N_13161);
nor U13721 (N_13721,N_13064,N_12728);
xnor U13722 (N_13722,N_12575,N_12041);
and U13723 (N_13723,N_12285,N_12288);
xnor U13724 (N_13724,N_13015,N_12131);
or U13725 (N_13725,N_12797,N_12091);
xnor U13726 (N_13726,N_12966,N_12830);
nor U13727 (N_13727,N_12034,N_12768);
nand U13728 (N_13728,N_12891,N_12497);
nor U13729 (N_13729,N_12081,N_12796);
nor U13730 (N_13730,N_12378,N_12347);
nand U13731 (N_13731,N_12841,N_13031);
nand U13732 (N_13732,N_13192,N_12815);
xnor U13733 (N_13733,N_12849,N_12313);
or U13734 (N_13734,N_12532,N_13149);
nor U13735 (N_13735,N_13159,N_13086);
nor U13736 (N_13736,N_13153,N_12251);
nand U13737 (N_13737,N_12328,N_12174);
nand U13738 (N_13738,N_12149,N_12824);
nand U13739 (N_13739,N_12300,N_12702);
or U13740 (N_13740,N_12729,N_12075);
xnor U13741 (N_13741,N_13075,N_13058);
nand U13742 (N_13742,N_12224,N_12727);
nand U13743 (N_13743,N_13157,N_12606);
xor U13744 (N_13744,N_12180,N_12653);
and U13745 (N_13745,N_12208,N_12695);
or U13746 (N_13746,N_12826,N_12825);
and U13747 (N_13747,N_13030,N_12605);
or U13748 (N_13748,N_12298,N_12200);
nand U13749 (N_13749,N_12505,N_12262);
nor U13750 (N_13750,N_12927,N_12201);
or U13751 (N_13751,N_12362,N_12257);
or U13752 (N_13752,N_12271,N_13008);
nor U13753 (N_13753,N_12674,N_12950);
xor U13754 (N_13754,N_12689,N_12851);
nor U13755 (N_13755,N_12478,N_13007);
xnor U13756 (N_13756,N_12510,N_12509);
nor U13757 (N_13757,N_13168,N_12317);
nand U13758 (N_13758,N_12907,N_12800);
nor U13759 (N_13759,N_12559,N_12617);
or U13760 (N_13760,N_12859,N_12527);
nor U13761 (N_13761,N_12638,N_12453);
nor U13762 (N_13762,N_12717,N_12376);
or U13763 (N_13763,N_13096,N_13170);
or U13764 (N_13764,N_12622,N_12514);
or U13765 (N_13765,N_13193,N_13188);
nor U13766 (N_13766,N_12352,N_12170);
nand U13767 (N_13767,N_12577,N_12778);
xnor U13768 (N_13768,N_13181,N_12480);
xnor U13769 (N_13769,N_12751,N_12754);
or U13770 (N_13770,N_12030,N_12401);
or U13771 (N_13771,N_12818,N_12064);
and U13772 (N_13772,N_12381,N_12368);
nand U13773 (N_13773,N_12680,N_12639);
or U13774 (N_13774,N_12252,N_12203);
nand U13775 (N_13775,N_12194,N_12793);
and U13776 (N_13776,N_12305,N_12812);
nand U13777 (N_13777,N_12933,N_12128);
xnor U13778 (N_13778,N_12582,N_13134);
or U13779 (N_13779,N_12154,N_12387);
xnor U13780 (N_13780,N_12853,N_12002);
nor U13781 (N_13781,N_13196,N_13130);
nor U13782 (N_13782,N_12424,N_12470);
nand U13783 (N_13783,N_12521,N_12705);
nand U13784 (N_13784,N_12038,N_12647);
xnor U13785 (N_13785,N_12542,N_12468);
nor U13786 (N_13786,N_12921,N_12415);
nand U13787 (N_13787,N_12889,N_12161);
nor U13788 (N_13788,N_12421,N_12655);
and U13789 (N_13789,N_12673,N_12916);
and U13790 (N_13790,N_12698,N_12999);
nand U13791 (N_13791,N_12467,N_13070);
or U13792 (N_13792,N_12371,N_12558);
and U13793 (N_13793,N_12987,N_12979);
and U13794 (N_13794,N_12008,N_13172);
and U13795 (N_13795,N_13199,N_12225);
xor U13796 (N_13796,N_12140,N_12561);
nand U13797 (N_13797,N_13048,N_13028);
nor U13798 (N_13798,N_12452,N_13045);
nor U13799 (N_13799,N_12472,N_12694);
or U13800 (N_13800,N_12708,N_12894);
or U13801 (N_13801,N_12579,N_12758);
xnor U13802 (N_13802,N_12194,N_12995);
and U13803 (N_13803,N_13126,N_13016);
nand U13804 (N_13804,N_12664,N_12811);
nor U13805 (N_13805,N_13021,N_12219);
and U13806 (N_13806,N_12899,N_12835);
nand U13807 (N_13807,N_12297,N_12352);
nor U13808 (N_13808,N_12292,N_13178);
or U13809 (N_13809,N_12182,N_12918);
nor U13810 (N_13810,N_12294,N_13007);
and U13811 (N_13811,N_13025,N_12678);
and U13812 (N_13812,N_12347,N_13056);
xnor U13813 (N_13813,N_12218,N_12389);
nand U13814 (N_13814,N_12125,N_12981);
nor U13815 (N_13815,N_13167,N_12399);
nor U13816 (N_13816,N_12427,N_12242);
nor U13817 (N_13817,N_12852,N_12700);
xnor U13818 (N_13818,N_13143,N_12992);
and U13819 (N_13819,N_12431,N_12139);
and U13820 (N_13820,N_12318,N_12759);
xor U13821 (N_13821,N_12655,N_12137);
and U13822 (N_13822,N_13053,N_12142);
nand U13823 (N_13823,N_12313,N_12055);
and U13824 (N_13824,N_12388,N_12524);
xor U13825 (N_13825,N_12204,N_12048);
nor U13826 (N_13826,N_12519,N_12293);
and U13827 (N_13827,N_12361,N_12557);
and U13828 (N_13828,N_12939,N_12862);
nor U13829 (N_13829,N_12001,N_12821);
nor U13830 (N_13830,N_12933,N_12810);
and U13831 (N_13831,N_12669,N_12282);
and U13832 (N_13832,N_12915,N_12865);
nand U13833 (N_13833,N_12225,N_12895);
nand U13834 (N_13834,N_12335,N_12465);
nor U13835 (N_13835,N_12357,N_12287);
and U13836 (N_13836,N_13042,N_12016);
xor U13837 (N_13837,N_13086,N_12894);
nand U13838 (N_13838,N_12506,N_13163);
xor U13839 (N_13839,N_13025,N_13164);
nand U13840 (N_13840,N_13115,N_12696);
nor U13841 (N_13841,N_12488,N_12943);
nor U13842 (N_13842,N_12679,N_12296);
xor U13843 (N_13843,N_12594,N_12872);
nand U13844 (N_13844,N_12712,N_12732);
or U13845 (N_13845,N_12000,N_12454);
nand U13846 (N_13846,N_12401,N_12744);
nand U13847 (N_13847,N_12980,N_12359);
or U13848 (N_13848,N_12335,N_12255);
or U13849 (N_13849,N_12197,N_12333);
xnor U13850 (N_13850,N_12978,N_12382);
nand U13851 (N_13851,N_13072,N_12104);
or U13852 (N_13852,N_13067,N_12329);
xor U13853 (N_13853,N_12537,N_12894);
nor U13854 (N_13854,N_13064,N_12664);
nor U13855 (N_13855,N_12161,N_12276);
nand U13856 (N_13856,N_12004,N_12150);
nor U13857 (N_13857,N_13085,N_12537);
and U13858 (N_13858,N_12483,N_12401);
nor U13859 (N_13859,N_13154,N_12089);
or U13860 (N_13860,N_12875,N_12852);
or U13861 (N_13861,N_13192,N_13136);
nor U13862 (N_13862,N_12823,N_12737);
nor U13863 (N_13863,N_12261,N_12280);
nand U13864 (N_13864,N_13193,N_12327);
xnor U13865 (N_13865,N_12119,N_12952);
and U13866 (N_13866,N_12534,N_12196);
nor U13867 (N_13867,N_12049,N_12037);
nand U13868 (N_13868,N_12105,N_13067);
nand U13869 (N_13869,N_13183,N_12774);
or U13870 (N_13870,N_12679,N_12125);
nand U13871 (N_13871,N_13002,N_12642);
or U13872 (N_13872,N_12723,N_12027);
xor U13873 (N_13873,N_12842,N_12469);
xor U13874 (N_13874,N_12545,N_12628);
nand U13875 (N_13875,N_12693,N_12349);
and U13876 (N_13876,N_12797,N_13028);
and U13877 (N_13877,N_12861,N_13045);
and U13878 (N_13878,N_12195,N_13165);
or U13879 (N_13879,N_12256,N_12481);
or U13880 (N_13880,N_12885,N_13033);
or U13881 (N_13881,N_13128,N_12945);
and U13882 (N_13882,N_12207,N_12073);
or U13883 (N_13883,N_12412,N_13095);
and U13884 (N_13884,N_12276,N_12280);
xnor U13885 (N_13885,N_12809,N_12053);
nand U13886 (N_13886,N_12633,N_12928);
and U13887 (N_13887,N_12394,N_12608);
nor U13888 (N_13888,N_12515,N_12979);
nor U13889 (N_13889,N_12260,N_12795);
nand U13890 (N_13890,N_13111,N_12211);
or U13891 (N_13891,N_12736,N_13181);
nor U13892 (N_13892,N_12576,N_12379);
nor U13893 (N_13893,N_12201,N_12030);
nor U13894 (N_13894,N_12483,N_12012);
nor U13895 (N_13895,N_12422,N_12244);
xnor U13896 (N_13896,N_12690,N_12751);
nand U13897 (N_13897,N_12079,N_12464);
nor U13898 (N_13898,N_12255,N_12620);
nand U13899 (N_13899,N_12733,N_12672);
xnor U13900 (N_13900,N_12213,N_12910);
and U13901 (N_13901,N_12451,N_12992);
xor U13902 (N_13902,N_13147,N_12186);
nand U13903 (N_13903,N_12760,N_12381);
or U13904 (N_13904,N_13176,N_12312);
nand U13905 (N_13905,N_12309,N_13139);
nand U13906 (N_13906,N_12360,N_12288);
or U13907 (N_13907,N_12180,N_12980);
and U13908 (N_13908,N_13114,N_12166);
xnor U13909 (N_13909,N_12067,N_12777);
nor U13910 (N_13910,N_12014,N_12645);
xor U13911 (N_13911,N_12265,N_12282);
nor U13912 (N_13912,N_12787,N_12367);
nand U13913 (N_13913,N_12780,N_12729);
nor U13914 (N_13914,N_12927,N_12946);
and U13915 (N_13915,N_12881,N_12709);
xnor U13916 (N_13916,N_12773,N_13086);
or U13917 (N_13917,N_12653,N_12654);
nor U13918 (N_13918,N_12135,N_12926);
and U13919 (N_13919,N_12177,N_12419);
and U13920 (N_13920,N_13081,N_12576);
or U13921 (N_13921,N_12825,N_12963);
and U13922 (N_13922,N_12419,N_12811);
nor U13923 (N_13923,N_13027,N_12802);
xor U13924 (N_13924,N_12601,N_13194);
nor U13925 (N_13925,N_12497,N_12778);
xnor U13926 (N_13926,N_12868,N_12056);
xnor U13927 (N_13927,N_12318,N_12606);
xor U13928 (N_13928,N_12800,N_12594);
nand U13929 (N_13929,N_13117,N_12258);
xnor U13930 (N_13930,N_12617,N_12237);
nor U13931 (N_13931,N_12789,N_12229);
xnor U13932 (N_13932,N_12422,N_12634);
nand U13933 (N_13933,N_12543,N_13182);
xnor U13934 (N_13934,N_12152,N_13088);
xor U13935 (N_13935,N_12180,N_12520);
nand U13936 (N_13936,N_13147,N_12536);
xnor U13937 (N_13937,N_12835,N_13070);
nor U13938 (N_13938,N_12498,N_12094);
nand U13939 (N_13939,N_12614,N_12502);
nor U13940 (N_13940,N_12876,N_12462);
or U13941 (N_13941,N_12622,N_12519);
and U13942 (N_13942,N_12767,N_12992);
nand U13943 (N_13943,N_12394,N_12510);
nor U13944 (N_13944,N_12693,N_12628);
nor U13945 (N_13945,N_12108,N_12046);
nor U13946 (N_13946,N_12655,N_12104);
nand U13947 (N_13947,N_12263,N_13110);
or U13948 (N_13948,N_12962,N_12310);
or U13949 (N_13949,N_12882,N_12346);
nor U13950 (N_13950,N_13150,N_12949);
nand U13951 (N_13951,N_12888,N_12433);
xor U13952 (N_13952,N_12297,N_12387);
nand U13953 (N_13953,N_12685,N_12559);
and U13954 (N_13954,N_12817,N_12443);
or U13955 (N_13955,N_12145,N_13165);
nand U13956 (N_13956,N_12289,N_12317);
nand U13957 (N_13957,N_12364,N_12027);
xor U13958 (N_13958,N_12249,N_12034);
nand U13959 (N_13959,N_12837,N_12792);
xor U13960 (N_13960,N_12484,N_12058);
xor U13961 (N_13961,N_12026,N_12523);
nor U13962 (N_13962,N_12525,N_12979);
and U13963 (N_13963,N_12806,N_12194);
and U13964 (N_13964,N_13099,N_12798);
nor U13965 (N_13965,N_12844,N_12413);
nor U13966 (N_13966,N_13155,N_13105);
xor U13967 (N_13967,N_12553,N_12721);
xor U13968 (N_13968,N_13153,N_12492);
or U13969 (N_13969,N_12765,N_12518);
xor U13970 (N_13970,N_12255,N_12375);
nor U13971 (N_13971,N_12875,N_12847);
and U13972 (N_13972,N_12976,N_12099);
xor U13973 (N_13973,N_12918,N_12405);
nand U13974 (N_13974,N_12185,N_12914);
nor U13975 (N_13975,N_12365,N_13142);
nor U13976 (N_13976,N_12099,N_12510);
nor U13977 (N_13977,N_12087,N_12573);
or U13978 (N_13978,N_12270,N_12689);
nor U13979 (N_13979,N_13152,N_12311);
nor U13980 (N_13980,N_12668,N_13021);
nand U13981 (N_13981,N_12478,N_12037);
nand U13982 (N_13982,N_12271,N_12026);
and U13983 (N_13983,N_13043,N_12794);
nand U13984 (N_13984,N_12860,N_12746);
nor U13985 (N_13985,N_12427,N_12485);
nor U13986 (N_13986,N_13159,N_13059);
nor U13987 (N_13987,N_13165,N_12762);
nor U13988 (N_13988,N_12057,N_12478);
and U13989 (N_13989,N_12591,N_12967);
xor U13990 (N_13990,N_12494,N_12834);
nor U13991 (N_13991,N_12744,N_12557);
or U13992 (N_13992,N_12350,N_12057);
and U13993 (N_13993,N_12014,N_12535);
or U13994 (N_13994,N_12790,N_12587);
and U13995 (N_13995,N_12083,N_12198);
nand U13996 (N_13996,N_12223,N_12048);
xnor U13997 (N_13997,N_12409,N_13014);
and U13998 (N_13998,N_12106,N_12719);
or U13999 (N_13999,N_13162,N_13050);
and U14000 (N_14000,N_12130,N_12054);
or U14001 (N_14001,N_12845,N_12411);
nand U14002 (N_14002,N_12581,N_12320);
nand U14003 (N_14003,N_12501,N_12970);
nor U14004 (N_14004,N_12215,N_12636);
nor U14005 (N_14005,N_12387,N_12246);
nand U14006 (N_14006,N_12025,N_12760);
nand U14007 (N_14007,N_12484,N_12949);
nor U14008 (N_14008,N_12951,N_12016);
xnor U14009 (N_14009,N_12564,N_12452);
or U14010 (N_14010,N_12729,N_12988);
nand U14011 (N_14011,N_12122,N_12557);
and U14012 (N_14012,N_13004,N_12102);
nand U14013 (N_14013,N_13144,N_12859);
nand U14014 (N_14014,N_12796,N_12566);
nor U14015 (N_14015,N_12030,N_12564);
nor U14016 (N_14016,N_12249,N_12240);
nor U14017 (N_14017,N_12627,N_12915);
nand U14018 (N_14018,N_13032,N_12910);
xor U14019 (N_14019,N_12049,N_12325);
nor U14020 (N_14020,N_12302,N_12341);
nand U14021 (N_14021,N_12645,N_12911);
or U14022 (N_14022,N_12778,N_12114);
xnor U14023 (N_14023,N_13063,N_12513);
or U14024 (N_14024,N_12283,N_12676);
or U14025 (N_14025,N_12091,N_12389);
nor U14026 (N_14026,N_12942,N_13095);
nand U14027 (N_14027,N_12531,N_12721);
and U14028 (N_14028,N_12653,N_12099);
and U14029 (N_14029,N_12989,N_12151);
xnor U14030 (N_14030,N_12887,N_12750);
nor U14031 (N_14031,N_12372,N_12062);
and U14032 (N_14032,N_12310,N_12989);
xnor U14033 (N_14033,N_12493,N_12172);
xnor U14034 (N_14034,N_12571,N_12256);
or U14035 (N_14035,N_12615,N_13105);
nor U14036 (N_14036,N_12509,N_12628);
and U14037 (N_14037,N_12889,N_13187);
xor U14038 (N_14038,N_12098,N_12485);
or U14039 (N_14039,N_12365,N_12422);
nor U14040 (N_14040,N_12576,N_12765);
xnor U14041 (N_14041,N_12439,N_12344);
or U14042 (N_14042,N_12870,N_12946);
nand U14043 (N_14043,N_12655,N_12418);
and U14044 (N_14044,N_13020,N_12274);
or U14045 (N_14045,N_12842,N_13145);
xnor U14046 (N_14046,N_12888,N_12292);
nand U14047 (N_14047,N_13165,N_12256);
xor U14048 (N_14048,N_12289,N_12374);
and U14049 (N_14049,N_12481,N_12791);
nand U14050 (N_14050,N_12726,N_12579);
nand U14051 (N_14051,N_13036,N_12354);
xnor U14052 (N_14052,N_12637,N_12551);
or U14053 (N_14053,N_12019,N_12405);
and U14054 (N_14054,N_12129,N_12560);
nor U14055 (N_14055,N_12804,N_12492);
or U14056 (N_14056,N_12967,N_12387);
xor U14057 (N_14057,N_12263,N_13121);
or U14058 (N_14058,N_12243,N_12490);
or U14059 (N_14059,N_12755,N_12586);
or U14060 (N_14060,N_12037,N_12701);
or U14061 (N_14061,N_12473,N_13167);
or U14062 (N_14062,N_13092,N_12667);
xor U14063 (N_14063,N_12020,N_12236);
xor U14064 (N_14064,N_12729,N_12921);
and U14065 (N_14065,N_12393,N_12009);
nor U14066 (N_14066,N_13036,N_12065);
nor U14067 (N_14067,N_12622,N_13034);
and U14068 (N_14068,N_12940,N_13193);
xnor U14069 (N_14069,N_13048,N_12761);
xnor U14070 (N_14070,N_12850,N_12578);
or U14071 (N_14071,N_12464,N_12433);
nand U14072 (N_14072,N_12242,N_13067);
and U14073 (N_14073,N_12565,N_13150);
nor U14074 (N_14074,N_12568,N_12107);
or U14075 (N_14075,N_12048,N_12264);
nor U14076 (N_14076,N_12902,N_12745);
xnor U14077 (N_14077,N_12547,N_13190);
xnor U14078 (N_14078,N_12884,N_12019);
or U14079 (N_14079,N_12087,N_12973);
and U14080 (N_14080,N_12129,N_12075);
nor U14081 (N_14081,N_13078,N_12232);
xnor U14082 (N_14082,N_12801,N_12268);
nand U14083 (N_14083,N_13006,N_12199);
nor U14084 (N_14084,N_12795,N_12959);
nand U14085 (N_14085,N_12674,N_12561);
nor U14086 (N_14086,N_12252,N_12404);
nand U14087 (N_14087,N_12973,N_13086);
nand U14088 (N_14088,N_12784,N_12562);
or U14089 (N_14089,N_12929,N_12972);
and U14090 (N_14090,N_13163,N_12502);
nand U14091 (N_14091,N_12160,N_12146);
nor U14092 (N_14092,N_12878,N_12211);
nor U14093 (N_14093,N_13130,N_12890);
and U14094 (N_14094,N_12737,N_12158);
nor U14095 (N_14095,N_12234,N_12564);
xnor U14096 (N_14096,N_12887,N_13146);
xnor U14097 (N_14097,N_12187,N_12683);
nor U14098 (N_14098,N_12088,N_12880);
and U14099 (N_14099,N_12405,N_12681);
nor U14100 (N_14100,N_13037,N_12553);
and U14101 (N_14101,N_12758,N_12388);
or U14102 (N_14102,N_12176,N_12024);
or U14103 (N_14103,N_12564,N_13068);
xor U14104 (N_14104,N_12815,N_12973);
or U14105 (N_14105,N_12647,N_13168);
nand U14106 (N_14106,N_13118,N_13188);
and U14107 (N_14107,N_12860,N_13072);
nand U14108 (N_14108,N_12664,N_12410);
xor U14109 (N_14109,N_12823,N_12810);
or U14110 (N_14110,N_12132,N_12316);
and U14111 (N_14111,N_12170,N_12790);
and U14112 (N_14112,N_12250,N_13049);
xor U14113 (N_14113,N_13154,N_13125);
or U14114 (N_14114,N_12380,N_13052);
or U14115 (N_14115,N_12026,N_13154);
nor U14116 (N_14116,N_12149,N_12390);
xnor U14117 (N_14117,N_12314,N_12555);
nor U14118 (N_14118,N_12347,N_12772);
nor U14119 (N_14119,N_12415,N_12793);
xor U14120 (N_14120,N_12283,N_12979);
or U14121 (N_14121,N_13095,N_13144);
or U14122 (N_14122,N_12487,N_12400);
nor U14123 (N_14123,N_12874,N_12005);
nor U14124 (N_14124,N_12853,N_12280);
xor U14125 (N_14125,N_12608,N_13166);
nand U14126 (N_14126,N_12531,N_12412);
nor U14127 (N_14127,N_13095,N_12513);
nor U14128 (N_14128,N_12644,N_12095);
nor U14129 (N_14129,N_13197,N_12168);
nand U14130 (N_14130,N_12278,N_12536);
or U14131 (N_14131,N_12498,N_12660);
or U14132 (N_14132,N_13167,N_12691);
nor U14133 (N_14133,N_12067,N_13008);
nand U14134 (N_14134,N_12923,N_13125);
or U14135 (N_14135,N_12935,N_12283);
nor U14136 (N_14136,N_12349,N_12375);
nor U14137 (N_14137,N_12558,N_12990);
nor U14138 (N_14138,N_12710,N_12976);
or U14139 (N_14139,N_12825,N_12609);
and U14140 (N_14140,N_12557,N_12784);
or U14141 (N_14141,N_12017,N_13154);
nor U14142 (N_14142,N_12483,N_12980);
nand U14143 (N_14143,N_12686,N_12430);
xor U14144 (N_14144,N_12602,N_12561);
nand U14145 (N_14145,N_12687,N_12539);
xnor U14146 (N_14146,N_12645,N_12667);
nand U14147 (N_14147,N_12153,N_12179);
and U14148 (N_14148,N_12495,N_12932);
and U14149 (N_14149,N_12196,N_12491);
nand U14150 (N_14150,N_12923,N_12372);
xor U14151 (N_14151,N_12900,N_12766);
and U14152 (N_14152,N_12202,N_12618);
nand U14153 (N_14153,N_12157,N_12109);
and U14154 (N_14154,N_13000,N_12914);
nand U14155 (N_14155,N_12992,N_12713);
nand U14156 (N_14156,N_12755,N_12039);
and U14157 (N_14157,N_12912,N_12637);
and U14158 (N_14158,N_12194,N_12661);
xor U14159 (N_14159,N_12741,N_12131);
and U14160 (N_14160,N_12163,N_12167);
and U14161 (N_14161,N_12886,N_12009);
or U14162 (N_14162,N_13151,N_12897);
xnor U14163 (N_14163,N_12779,N_12731);
nand U14164 (N_14164,N_12188,N_13054);
xor U14165 (N_14165,N_12626,N_12905);
or U14166 (N_14166,N_12811,N_12899);
and U14167 (N_14167,N_12991,N_12236);
xnor U14168 (N_14168,N_12899,N_12231);
nand U14169 (N_14169,N_12707,N_12797);
nor U14170 (N_14170,N_12621,N_12047);
or U14171 (N_14171,N_12206,N_12458);
nor U14172 (N_14172,N_12524,N_12403);
nand U14173 (N_14173,N_12847,N_12190);
and U14174 (N_14174,N_12185,N_12024);
and U14175 (N_14175,N_13128,N_12179);
nand U14176 (N_14176,N_12662,N_13030);
or U14177 (N_14177,N_12138,N_12158);
nand U14178 (N_14178,N_12183,N_12505);
xor U14179 (N_14179,N_12839,N_12108);
xnor U14180 (N_14180,N_12562,N_12093);
nand U14181 (N_14181,N_12093,N_12490);
or U14182 (N_14182,N_12256,N_12390);
xor U14183 (N_14183,N_12712,N_12897);
xnor U14184 (N_14184,N_13146,N_12557);
xor U14185 (N_14185,N_12889,N_12742);
nand U14186 (N_14186,N_12098,N_12964);
nor U14187 (N_14187,N_12349,N_12333);
or U14188 (N_14188,N_12849,N_12868);
xor U14189 (N_14189,N_12795,N_13129);
nor U14190 (N_14190,N_12235,N_12194);
xor U14191 (N_14191,N_12274,N_12462);
or U14192 (N_14192,N_12524,N_12851);
nand U14193 (N_14193,N_12403,N_12390);
nor U14194 (N_14194,N_12660,N_12481);
nand U14195 (N_14195,N_12537,N_12675);
nand U14196 (N_14196,N_12168,N_12403);
nand U14197 (N_14197,N_12247,N_12508);
nand U14198 (N_14198,N_12310,N_12936);
and U14199 (N_14199,N_12564,N_12749);
or U14200 (N_14200,N_12191,N_12563);
and U14201 (N_14201,N_12358,N_13004);
or U14202 (N_14202,N_12005,N_12327);
and U14203 (N_14203,N_12698,N_12991);
or U14204 (N_14204,N_12865,N_12952);
or U14205 (N_14205,N_12108,N_12241);
and U14206 (N_14206,N_12089,N_12912);
nand U14207 (N_14207,N_12262,N_12961);
nor U14208 (N_14208,N_12393,N_12333);
nand U14209 (N_14209,N_12245,N_12820);
or U14210 (N_14210,N_12259,N_12879);
and U14211 (N_14211,N_12371,N_12853);
nor U14212 (N_14212,N_12173,N_12888);
and U14213 (N_14213,N_12840,N_12182);
and U14214 (N_14214,N_12496,N_12787);
xor U14215 (N_14215,N_12190,N_13046);
nor U14216 (N_14216,N_12883,N_12156);
and U14217 (N_14217,N_12264,N_12552);
or U14218 (N_14218,N_12508,N_13133);
and U14219 (N_14219,N_12457,N_12910);
nor U14220 (N_14220,N_12982,N_12197);
nor U14221 (N_14221,N_12541,N_12511);
or U14222 (N_14222,N_12069,N_12117);
xor U14223 (N_14223,N_12486,N_12781);
nand U14224 (N_14224,N_12894,N_13161);
nor U14225 (N_14225,N_12066,N_13050);
or U14226 (N_14226,N_13146,N_12664);
nor U14227 (N_14227,N_12830,N_12550);
and U14228 (N_14228,N_13052,N_12246);
or U14229 (N_14229,N_12897,N_12469);
nand U14230 (N_14230,N_12255,N_12102);
and U14231 (N_14231,N_12817,N_13141);
and U14232 (N_14232,N_12414,N_12503);
nand U14233 (N_14233,N_12970,N_13077);
nor U14234 (N_14234,N_12971,N_12897);
nor U14235 (N_14235,N_13147,N_12014);
and U14236 (N_14236,N_12342,N_12451);
and U14237 (N_14237,N_12995,N_12017);
or U14238 (N_14238,N_12522,N_12015);
nor U14239 (N_14239,N_13110,N_12977);
and U14240 (N_14240,N_12290,N_13119);
or U14241 (N_14241,N_12495,N_12394);
nand U14242 (N_14242,N_12740,N_13080);
and U14243 (N_14243,N_12237,N_12375);
or U14244 (N_14244,N_13196,N_12699);
xnor U14245 (N_14245,N_13011,N_12380);
xnor U14246 (N_14246,N_13094,N_12377);
or U14247 (N_14247,N_12980,N_12036);
nand U14248 (N_14248,N_12846,N_12261);
or U14249 (N_14249,N_12567,N_13077);
and U14250 (N_14250,N_13199,N_12499);
xnor U14251 (N_14251,N_12221,N_12914);
and U14252 (N_14252,N_12922,N_13063);
xor U14253 (N_14253,N_12459,N_12293);
or U14254 (N_14254,N_12044,N_13123);
xor U14255 (N_14255,N_12923,N_12726);
and U14256 (N_14256,N_12374,N_12954);
xnor U14257 (N_14257,N_12236,N_12329);
xor U14258 (N_14258,N_12681,N_12317);
nand U14259 (N_14259,N_12696,N_12370);
nor U14260 (N_14260,N_12272,N_12692);
and U14261 (N_14261,N_12652,N_12903);
nor U14262 (N_14262,N_12647,N_12664);
nand U14263 (N_14263,N_12517,N_12221);
nor U14264 (N_14264,N_12006,N_12279);
xor U14265 (N_14265,N_12858,N_12791);
and U14266 (N_14266,N_12277,N_12650);
nand U14267 (N_14267,N_12067,N_12123);
xnor U14268 (N_14268,N_12010,N_12793);
and U14269 (N_14269,N_12171,N_12462);
nand U14270 (N_14270,N_13023,N_12190);
xnor U14271 (N_14271,N_12964,N_12725);
nor U14272 (N_14272,N_12069,N_13118);
and U14273 (N_14273,N_12185,N_12111);
nor U14274 (N_14274,N_12501,N_12018);
or U14275 (N_14275,N_12804,N_13077);
xor U14276 (N_14276,N_12520,N_12391);
and U14277 (N_14277,N_12851,N_12839);
nor U14278 (N_14278,N_12110,N_12646);
nand U14279 (N_14279,N_12032,N_12074);
and U14280 (N_14280,N_12414,N_12159);
nand U14281 (N_14281,N_12250,N_13121);
and U14282 (N_14282,N_12670,N_12660);
and U14283 (N_14283,N_13045,N_13074);
nor U14284 (N_14284,N_12764,N_13197);
or U14285 (N_14285,N_13129,N_12646);
and U14286 (N_14286,N_12754,N_13005);
and U14287 (N_14287,N_12467,N_12546);
nor U14288 (N_14288,N_12454,N_12614);
nand U14289 (N_14289,N_12837,N_12523);
nor U14290 (N_14290,N_12952,N_12737);
nor U14291 (N_14291,N_13132,N_12412);
and U14292 (N_14292,N_13053,N_12707);
and U14293 (N_14293,N_13172,N_12345);
or U14294 (N_14294,N_12943,N_12098);
and U14295 (N_14295,N_12276,N_12720);
xor U14296 (N_14296,N_13040,N_12515);
xor U14297 (N_14297,N_12100,N_13036);
nand U14298 (N_14298,N_12735,N_13164);
and U14299 (N_14299,N_12083,N_12692);
xnor U14300 (N_14300,N_12221,N_12366);
xor U14301 (N_14301,N_12466,N_12228);
and U14302 (N_14302,N_12512,N_12114);
and U14303 (N_14303,N_12514,N_12742);
xor U14304 (N_14304,N_12861,N_12669);
and U14305 (N_14305,N_12166,N_12077);
nor U14306 (N_14306,N_12272,N_12690);
xor U14307 (N_14307,N_12579,N_12301);
nand U14308 (N_14308,N_12766,N_12132);
and U14309 (N_14309,N_13157,N_13099);
xor U14310 (N_14310,N_13035,N_12296);
nand U14311 (N_14311,N_12455,N_12731);
and U14312 (N_14312,N_12799,N_12623);
and U14313 (N_14313,N_13038,N_12211);
nand U14314 (N_14314,N_12277,N_12198);
xnor U14315 (N_14315,N_13058,N_12268);
nand U14316 (N_14316,N_12701,N_12915);
xnor U14317 (N_14317,N_12178,N_12301);
or U14318 (N_14318,N_12452,N_12572);
xnor U14319 (N_14319,N_12796,N_12286);
nor U14320 (N_14320,N_12516,N_12039);
or U14321 (N_14321,N_12589,N_12800);
and U14322 (N_14322,N_12928,N_12382);
nand U14323 (N_14323,N_12187,N_13141);
nor U14324 (N_14324,N_12687,N_12233);
xnor U14325 (N_14325,N_12174,N_12095);
nor U14326 (N_14326,N_12638,N_13185);
nand U14327 (N_14327,N_12910,N_12158);
nand U14328 (N_14328,N_12364,N_12426);
xor U14329 (N_14329,N_12289,N_12666);
and U14330 (N_14330,N_12025,N_13017);
xor U14331 (N_14331,N_12267,N_12216);
nand U14332 (N_14332,N_12172,N_12897);
and U14333 (N_14333,N_12736,N_13028);
nor U14334 (N_14334,N_12516,N_12062);
and U14335 (N_14335,N_12811,N_12838);
and U14336 (N_14336,N_12746,N_12464);
and U14337 (N_14337,N_12295,N_13137);
or U14338 (N_14338,N_13174,N_12222);
xor U14339 (N_14339,N_12687,N_12088);
and U14340 (N_14340,N_12967,N_12672);
and U14341 (N_14341,N_12234,N_12448);
xor U14342 (N_14342,N_12618,N_12888);
nand U14343 (N_14343,N_12438,N_12943);
or U14344 (N_14344,N_13115,N_13087);
or U14345 (N_14345,N_12739,N_12493);
nor U14346 (N_14346,N_12103,N_12671);
or U14347 (N_14347,N_12358,N_12460);
xnor U14348 (N_14348,N_12476,N_13091);
nor U14349 (N_14349,N_12696,N_12536);
and U14350 (N_14350,N_13136,N_12923);
or U14351 (N_14351,N_12635,N_12181);
xor U14352 (N_14352,N_12905,N_12556);
nor U14353 (N_14353,N_13137,N_12040);
or U14354 (N_14354,N_12283,N_12777);
nand U14355 (N_14355,N_12560,N_13176);
or U14356 (N_14356,N_12541,N_12810);
xnor U14357 (N_14357,N_12995,N_12202);
or U14358 (N_14358,N_12606,N_12906);
xor U14359 (N_14359,N_12697,N_12462);
xnor U14360 (N_14360,N_12656,N_12022);
and U14361 (N_14361,N_12468,N_12166);
and U14362 (N_14362,N_12109,N_12939);
and U14363 (N_14363,N_12146,N_12385);
and U14364 (N_14364,N_12316,N_12493);
nand U14365 (N_14365,N_12074,N_13179);
nand U14366 (N_14366,N_12932,N_12510);
xnor U14367 (N_14367,N_12806,N_12638);
nor U14368 (N_14368,N_12936,N_12050);
and U14369 (N_14369,N_12200,N_13061);
nor U14370 (N_14370,N_12927,N_12158);
nand U14371 (N_14371,N_12379,N_12206);
nor U14372 (N_14372,N_12546,N_12155);
or U14373 (N_14373,N_12894,N_13000);
nand U14374 (N_14374,N_12724,N_12691);
nand U14375 (N_14375,N_12580,N_12119);
and U14376 (N_14376,N_12640,N_12365);
nor U14377 (N_14377,N_12264,N_12371);
nand U14378 (N_14378,N_13163,N_12362);
xnor U14379 (N_14379,N_12082,N_12711);
xnor U14380 (N_14380,N_13069,N_12029);
nand U14381 (N_14381,N_12122,N_12763);
nor U14382 (N_14382,N_13174,N_12074);
xor U14383 (N_14383,N_12840,N_13029);
or U14384 (N_14384,N_12374,N_12940);
or U14385 (N_14385,N_13084,N_12863);
nor U14386 (N_14386,N_12368,N_12029);
nand U14387 (N_14387,N_12069,N_12441);
xnor U14388 (N_14388,N_12395,N_12722);
or U14389 (N_14389,N_12020,N_12533);
nand U14390 (N_14390,N_12164,N_12132);
xnor U14391 (N_14391,N_12520,N_12628);
nor U14392 (N_14392,N_12441,N_13167);
xor U14393 (N_14393,N_12487,N_12122);
nand U14394 (N_14394,N_12069,N_12185);
xnor U14395 (N_14395,N_12584,N_13011);
nor U14396 (N_14396,N_12015,N_12526);
nand U14397 (N_14397,N_12115,N_12575);
or U14398 (N_14398,N_12801,N_12540);
or U14399 (N_14399,N_12707,N_12309);
nor U14400 (N_14400,N_14203,N_13929);
nor U14401 (N_14401,N_13787,N_14193);
and U14402 (N_14402,N_14140,N_13873);
xor U14403 (N_14403,N_13515,N_13745);
and U14404 (N_14404,N_13721,N_13453);
and U14405 (N_14405,N_14122,N_14345);
nor U14406 (N_14406,N_13661,N_13848);
nand U14407 (N_14407,N_13459,N_14190);
nor U14408 (N_14408,N_14396,N_13240);
and U14409 (N_14409,N_14314,N_14337);
nand U14410 (N_14410,N_13755,N_14038);
and U14411 (N_14411,N_13920,N_14353);
nor U14412 (N_14412,N_13671,N_13539);
xnor U14413 (N_14413,N_14305,N_13563);
or U14414 (N_14414,N_13783,N_14044);
and U14415 (N_14415,N_14136,N_13485);
or U14416 (N_14416,N_13341,N_14301);
or U14417 (N_14417,N_13296,N_13207);
nor U14418 (N_14418,N_13514,N_13319);
xnor U14419 (N_14419,N_13982,N_13821);
and U14420 (N_14420,N_13407,N_13952);
nor U14421 (N_14421,N_13224,N_14178);
nor U14422 (N_14422,N_13217,N_13531);
nor U14423 (N_14423,N_13849,N_13827);
xnor U14424 (N_14424,N_14053,N_13942);
nor U14425 (N_14425,N_13964,N_13494);
nand U14426 (N_14426,N_13340,N_13447);
nor U14427 (N_14427,N_13321,N_13985);
and U14428 (N_14428,N_13512,N_13616);
or U14429 (N_14429,N_13290,N_13245);
xnor U14430 (N_14430,N_14105,N_13715);
or U14431 (N_14431,N_13639,N_13660);
xor U14432 (N_14432,N_13590,N_13579);
nand U14433 (N_14433,N_13792,N_14196);
or U14434 (N_14434,N_14008,N_13901);
nand U14435 (N_14435,N_13853,N_13753);
and U14436 (N_14436,N_13936,N_13550);
xor U14437 (N_14437,N_13423,N_13835);
or U14438 (N_14438,N_13683,N_13606);
xnor U14439 (N_14439,N_13306,N_13438);
nand U14440 (N_14440,N_13836,N_13642);
and U14441 (N_14441,N_14232,N_13749);
or U14442 (N_14442,N_13713,N_14030);
and U14443 (N_14443,N_14321,N_14060);
xor U14444 (N_14444,N_13347,N_13211);
xnor U14445 (N_14445,N_14253,N_13264);
nand U14446 (N_14446,N_14341,N_13335);
xor U14447 (N_14447,N_14137,N_14179);
xnor U14448 (N_14448,N_14094,N_13561);
nand U14449 (N_14449,N_13786,N_13497);
nand U14450 (N_14450,N_14183,N_14120);
nor U14451 (N_14451,N_13720,N_13948);
xnor U14452 (N_14452,N_14207,N_14151);
xor U14453 (N_14453,N_14174,N_14262);
xor U14454 (N_14454,N_14263,N_13719);
xnor U14455 (N_14455,N_13578,N_13268);
xor U14456 (N_14456,N_13300,N_14258);
and U14457 (N_14457,N_13338,N_13957);
nor U14458 (N_14458,N_14343,N_14319);
nor U14459 (N_14459,N_13656,N_14168);
nand U14460 (N_14460,N_13443,N_13595);
or U14461 (N_14461,N_13962,N_13331);
nand U14462 (N_14462,N_13665,N_13612);
and U14463 (N_14463,N_14013,N_14288);
and U14464 (N_14464,N_14330,N_14074);
nor U14465 (N_14465,N_13591,N_14054);
and U14466 (N_14466,N_13686,N_13261);
xor U14467 (N_14467,N_14176,N_13898);
nor U14468 (N_14468,N_14004,N_14336);
nor U14469 (N_14469,N_14089,N_14049);
or U14470 (N_14470,N_14302,N_14043);
nor U14471 (N_14471,N_13712,N_13470);
nor U14472 (N_14472,N_13634,N_14028);
and U14473 (N_14473,N_14270,N_13846);
or U14474 (N_14474,N_13343,N_14068);
or U14475 (N_14475,N_13249,N_13458);
and U14476 (N_14476,N_14208,N_14329);
xor U14477 (N_14477,N_13894,N_14058);
nor U14478 (N_14478,N_14388,N_13482);
nor U14479 (N_14479,N_13337,N_13789);
and U14480 (N_14480,N_13259,N_14006);
and U14481 (N_14481,N_13492,N_13609);
or U14482 (N_14482,N_14128,N_13658);
and U14483 (N_14483,N_14078,N_13980);
or U14484 (N_14484,N_14310,N_13698);
and U14485 (N_14485,N_14211,N_13927);
nand U14486 (N_14486,N_13554,N_13843);
nor U14487 (N_14487,N_14047,N_13450);
xor U14488 (N_14488,N_14346,N_14217);
nor U14489 (N_14489,N_13205,N_13733);
xnor U14490 (N_14490,N_14248,N_13823);
or U14491 (N_14491,N_13604,N_13750);
and U14492 (N_14492,N_14086,N_14278);
nand U14493 (N_14493,N_14342,N_14308);
or U14494 (N_14494,N_13232,N_14260);
xor U14495 (N_14495,N_13722,N_13299);
nand U14496 (N_14496,N_13857,N_13670);
nand U14497 (N_14497,N_13687,N_13707);
or U14498 (N_14498,N_13781,N_14103);
nand U14499 (N_14499,N_14095,N_14204);
and U14500 (N_14500,N_13778,N_14017);
and U14501 (N_14501,N_13363,N_13852);
and U14502 (N_14502,N_13969,N_13931);
xor U14503 (N_14503,N_13914,N_14261);
xnor U14504 (N_14504,N_14134,N_13371);
and U14505 (N_14505,N_13882,N_13999);
nand U14506 (N_14506,N_13412,N_13283);
nand U14507 (N_14507,N_14188,N_13418);
xnor U14508 (N_14508,N_13565,N_13355);
nand U14509 (N_14509,N_13206,N_14218);
xnor U14510 (N_14510,N_13972,N_13735);
or U14511 (N_14511,N_13488,N_14340);
or U14512 (N_14512,N_13904,N_13717);
xnor U14513 (N_14513,N_13394,N_14173);
xnor U14514 (N_14514,N_13677,N_13788);
and U14515 (N_14515,N_14275,N_14266);
and U14516 (N_14516,N_13699,N_14376);
nand U14517 (N_14517,N_14399,N_14177);
nor U14518 (N_14518,N_13732,N_13923);
or U14519 (N_14519,N_13430,N_14077);
nand U14520 (N_14520,N_13681,N_14228);
xnor U14521 (N_14521,N_13480,N_14117);
or U14522 (N_14522,N_14011,N_14156);
and U14523 (N_14523,N_13820,N_14000);
and U14524 (N_14524,N_13771,N_13489);
nor U14525 (N_14525,N_13758,N_13344);
nand U14526 (N_14526,N_13888,N_13332);
nor U14527 (N_14527,N_14127,N_14390);
nor U14528 (N_14528,N_14363,N_13596);
nand U14529 (N_14529,N_14045,N_13621);
or U14530 (N_14530,N_13404,N_13708);
xor U14531 (N_14531,N_14227,N_13932);
and U14532 (N_14532,N_13504,N_13210);
nand U14533 (N_14533,N_14322,N_14056);
xor U14534 (N_14534,N_14298,N_13669);
xor U14535 (N_14535,N_13776,N_13653);
and U14536 (N_14536,N_13968,N_14306);
or U14537 (N_14537,N_13560,N_13441);
nor U14538 (N_14538,N_13916,N_14025);
or U14539 (N_14539,N_13826,N_13572);
and U14540 (N_14540,N_14237,N_13599);
nand U14541 (N_14541,N_14328,N_13295);
nor U14542 (N_14542,N_13602,N_13314);
or U14543 (N_14543,N_13472,N_13231);
nand U14544 (N_14544,N_14316,N_13463);
and U14545 (N_14545,N_14130,N_13933);
and U14546 (N_14546,N_13950,N_13945);
nor U14547 (N_14547,N_13524,N_13905);
nand U14548 (N_14548,N_13954,N_13203);
nor U14549 (N_14549,N_13416,N_14032);
xor U14550 (N_14550,N_13958,N_14338);
nor U14551 (N_14551,N_13659,N_14398);
nor U14552 (N_14552,N_13695,N_13348);
nand U14553 (N_14553,N_13705,N_13824);
nand U14554 (N_14554,N_13608,N_13375);
nand U14555 (N_14555,N_13626,N_13651);
nor U14556 (N_14556,N_13493,N_14065);
and U14557 (N_14557,N_13637,N_13541);
nand U14558 (N_14558,N_14239,N_13468);
or U14559 (N_14559,N_14285,N_14313);
xor U14560 (N_14560,N_13487,N_13839);
nand U14561 (N_14561,N_14093,N_13770);
and U14562 (N_14562,N_14022,N_14215);
or U14563 (N_14563,N_13513,N_13614);
nor U14564 (N_14564,N_13395,N_14225);
and U14565 (N_14565,N_14115,N_13924);
xnor U14566 (N_14566,N_14146,N_14231);
and U14567 (N_14567,N_13522,N_14100);
xnor U14568 (N_14568,N_13235,N_14080);
nor U14569 (N_14569,N_13528,N_13877);
or U14570 (N_14570,N_13293,N_13833);
nor U14571 (N_14571,N_14297,N_14166);
and U14572 (N_14572,N_14354,N_14244);
nand U14573 (N_14573,N_13435,N_14073);
nand U14574 (N_14574,N_13403,N_13361);
or U14575 (N_14575,N_13704,N_13456);
xnor U14576 (N_14576,N_14057,N_14165);
xnor U14577 (N_14577,N_13775,N_14023);
nor U14578 (N_14578,N_13501,N_13349);
xnor U14579 (N_14579,N_13584,N_13803);
xor U14580 (N_14580,N_13992,N_14265);
nor U14581 (N_14581,N_13908,N_13483);
nor U14582 (N_14582,N_13866,N_13861);
nor U14583 (N_14583,N_13844,N_13411);
nand U14584 (N_14584,N_13391,N_13318);
and U14585 (N_14585,N_13938,N_14251);
nor U14586 (N_14586,N_13542,N_13213);
or U14587 (N_14587,N_13397,N_13367);
nor U14588 (N_14588,N_13219,N_14087);
xor U14589 (N_14589,N_13913,N_13376);
xnor U14590 (N_14590,N_14175,N_13613);
xor U14591 (N_14591,N_14169,N_14163);
nor U14592 (N_14592,N_14090,N_13657);
nand U14593 (N_14593,N_13362,N_13855);
and U14594 (N_14594,N_13706,N_13620);
nor U14595 (N_14595,N_13947,N_13520);
nor U14596 (N_14596,N_13988,N_14294);
or U14597 (N_14597,N_13473,N_13436);
xor U14598 (N_14598,N_13280,N_14061);
nor U14599 (N_14599,N_13762,N_13703);
xnor U14600 (N_14600,N_13214,N_13648);
and U14601 (N_14601,N_13736,N_13433);
nor U14602 (N_14602,N_13727,N_14132);
nand U14603 (N_14603,N_13384,N_14250);
or U14604 (N_14604,N_13804,N_13327);
nor U14605 (N_14605,N_13500,N_14158);
or U14606 (N_14606,N_14256,N_14172);
nor U14607 (N_14607,N_14002,N_14113);
or U14608 (N_14608,N_13242,N_13491);
xnor U14609 (N_14609,N_13334,N_13558);
or U14610 (N_14610,N_14167,N_14198);
nand U14611 (N_14611,N_13955,N_13495);
nand U14612 (N_14612,N_13576,N_14069);
xnor U14613 (N_14613,N_13258,N_13734);
and U14614 (N_14614,N_14299,N_13464);
nor U14615 (N_14615,N_13311,N_14318);
nand U14616 (N_14616,N_14397,N_14352);
nand U14617 (N_14617,N_14282,N_13260);
and U14618 (N_14618,N_14213,N_14331);
and U14619 (N_14619,N_13477,N_13265);
nand U14620 (N_14620,N_13586,N_14351);
xnor U14621 (N_14621,N_13409,N_14223);
xnor U14622 (N_14622,N_13352,N_14064);
nor U14623 (N_14623,N_14361,N_13233);
xnor U14624 (N_14624,N_14212,N_14037);
or U14625 (N_14625,N_14210,N_13697);
nor U14626 (N_14626,N_13215,N_13401);
and U14627 (N_14627,N_14154,N_13377);
nor U14628 (N_14628,N_13806,N_13588);
or U14629 (N_14629,N_13809,N_14186);
nor U14630 (N_14630,N_14255,N_13617);
or U14631 (N_14631,N_13997,N_14320);
nor U14632 (N_14632,N_13868,N_14300);
or U14633 (N_14633,N_14234,N_13593);
nor U14634 (N_14634,N_13346,N_13990);
and U14635 (N_14635,N_13742,N_13538);
nor U14636 (N_14636,N_14076,N_13519);
nor U14637 (N_14637,N_13752,N_13413);
or U14638 (N_14638,N_14135,N_13396);
nand U14639 (N_14639,N_14161,N_13850);
xor U14640 (N_14640,N_14194,N_13312);
or U14641 (N_14641,N_13802,N_13622);
or U14642 (N_14642,N_13829,N_13269);
nor U14643 (N_14643,N_13801,N_13452);
or U14644 (N_14644,N_13336,N_13284);
or U14645 (N_14645,N_13582,N_13879);
nand U14646 (N_14646,N_13815,N_14171);
nor U14647 (N_14647,N_14139,N_14170);
xor U14648 (N_14648,N_14291,N_14119);
or U14649 (N_14649,N_14111,N_14019);
and U14650 (N_14650,N_13667,N_13603);
or U14651 (N_14651,N_13814,N_13981);
or U14652 (N_14652,N_13429,N_13949);
nand U14653 (N_14653,N_13390,N_13325);
and U14654 (N_14654,N_13222,N_13445);
nand U14655 (N_14655,N_13887,N_14041);
nand U14656 (N_14656,N_13666,N_13816);
nor U14657 (N_14657,N_13310,N_14238);
xor U14658 (N_14658,N_13819,N_13454);
nand U14659 (N_14659,N_14355,N_13571);
and U14660 (N_14660,N_13966,N_14051);
nor U14661 (N_14661,N_13448,N_13257);
xnor U14662 (N_14662,N_14245,N_13529);
and U14663 (N_14663,N_13961,N_14254);
nor U14664 (N_14664,N_13886,N_13973);
and U14665 (N_14665,N_13370,N_13818);
nand U14666 (N_14666,N_13368,N_14380);
or U14667 (N_14667,N_14145,N_14116);
or U14668 (N_14668,N_13523,N_13763);
or U14669 (N_14669,N_14372,N_13568);
nand U14670 (N_14670,N_13323,N_14205);
nor U14671 (N_14671,N_13339,N_13974);
or U14672 (N_14672,N_13526,N_13518);
or U14673 (N_14673,N_13746,N_13780);
and U14674 (N_14674,N_14233,N_13891);
xor U14675 (N_14675,N_13379,N_13530);
nand U14676 (N_14676,N_14366,N_13684);
nor U14677 (N_14677,N_14121,N_14379);
or U14678 (N_14678,N_13393,N_14187);
or U14679 (N_14679,N_13625,N_14085);
and U14680 (N_14680,N_13897,N_13747);
or U14681 (N_14681,N_13305,N_14184);
nor U14682 (N_14682,N_13592,N_13793);
xnor U14683 (N_14683,N_13825,N_13466);
or U14684 (N_14684,N_14209,N_13986);
nand U14685 (N_14685,N_13896,N_14035);
or U14686 (N_14686,N_13354,N_13641);
nand U14687 (N_14687,N_13226,N_14277);
nand U14688 (N_14688,N_13469,N_14036);
xnor U14689 (N_14689,N_13587,N_14375);
nor U14690 (N_14690,N_13883,N_13556);
or U14691 (N_14691,N_14200,N_13859);
and U14692 (N_14692,N_13930,N_13303);
nor U14693 (N_14693,N_13615,N_13724);
and U14694 (N_14694,N_13505,N_13381);
xnor U14695 (N_14695,N_13508,N_14382);
and U14696 (N_14696,N_14142,N_13860);
xor U14697 (N_14697,N_13817,N_14040);
nand U14698 (N_14698,N_13643,N_13243);
and U14699 (N_14699,N_13629,N_13754);
and U14700 (N_14700,N_13449,N_13864);
and U14701 (N_14701,N_13800,N_13646);
or U14702 (N_14702,N_14129,N_13989);
or U14703 (N_14703,N_13543,N_14155);
nand U14704 (N_14704,N_13330,N_13967);
nand U14705 (N_14705,N_13907,N_14222);
xor U14706 (N_14706,N_13479,N_13941);
xnor U14707 (N_14707,N_14109,N_13333);
xor U14708 (N_14708,N_13872,N_13509);
nand U14709 (N_14709,N_14348,N_13751);
or U14710 (N_14710,N_13632,N_13238);
xnor U14711 (N_14711,N_14349,N_13965);
nand U14712 (N_14712,N_14162,N_13840);
xor U14713 (N_14713,N_13970,N_13672);
or U14714 (N_14714,N_13380,N_14104);
xor U14715 (N_14715,N_13553,N_14384);
xnor U14716 (N_14716,N_13583,N_13200);
nor U14717 (N_14717,N_14050,N_14125);
nor U14718 (N_14718,N_13378,N_13790);
nor U14719 (N_14719,N_13507,N_13741);
nand U14720 (N_14720,N_13977,N_13884);
xor U14721 (N_14721,N_14191,N_13607);
or U14722 (N_14722,N_14098,N_14026);
or U14723 (N_14723,N_14383,N_13533);
and U14724 (N_14724,N_14071,N_14229);
nor U14725 (N_14725,N_13984,N_14257);
and U14726 (N_14726,N_13534,N_13995);
nor U14727 (N_14727,N_14230,N_14206);
xor U14728 (N_14728,N_13517,N_13960);
nand U14729 (N_14729,N_14048,N_13419);
or U14730 (N_14730,N_13208,N_14333);
and U14731 (N_14731,N_13421,N_13701);
nand U14732 (N_14732,N_13716,N_13976);
xnor U14733 (N_14733,N_14020,N_13502);
nand U14734 (N_14734,N_14377,N_14003);
and U14735 (N_14735,N_14042,N_13385);
xor U14736 (N_14736,N_13481,N_14079);
and U14737 (N_14737,N_14276,N_13212);
nor U14738 (N_14738,N_13313,N_13324);
and U14739 (N_14739,N_13241,N_14101);
nand U14740 (N_14740,N_14016,N_14339);
nand U14741 (N_14741,N_13405,N_13460);
nand U14742 (N_14742,N_14034,N_13434);
xor U14743 (N_14743,N_14367,N_13221);
or U14744 (N_14744,N_13702,N_14327);
and U14745 (N_14745,N_13983,N_13766);
or U14746 (N_14746,N_14334,N_14009);
xnor U14747 (N_14747,N_13725,N_14392);
or U14748 (N_14748,N_13700,N_14235);
nand U14749 (N_14749,N_13834,N_14293);
nand U14750 (N_14750,N_13428,N_14387);
or U14751 (N_14751,N_14356,N_14062);
nand U14752 (N_14752,N_13871,N_13906);
nor U14753 (N_14753,N_14102,N_13810);
xor U14754 (N_14754,N_13777,N_14148);
and U14755 (N_14755,N_14046,N_13358);
nor U14756 (N_14756,N_13227,N_13490);
and U14757 (N_14757,N_14014,N_14133);
nand U14758 (N_14758,N_13228,N_13889);
nand U14759 (N_14759,N_13425,N_13427);
xor U14760 (N_14760,N_13546,N_14052);
nand U14761 (N_14761,N_13544,N_13611);
nand U14762 (N_14762,N_13636,N_14099);
and U14763 (N_14763,N_13691,N_13710);
nor U14764 (N_14764,N_13287,N_13255);
or U14765 (N_14765,N_13917,N_13773);
xnor U14766 (N_14766,N_13743,N_13581);
nand U14767 (N_14767,N_13663,N_14389);
xor U14768 (N_14768,N_13253,N_13890);
xnor U14769 (N_14769,N_14202,N_13784);
nor U14770 (N_14770,N_13444,N_13442);
and U14771 (N_14771,N_14005,N_13838);
nand U14772 (N_14772,N_13645,N_13457);
and U14773 (N_14773,N_13322,N_13365);
xor U14774 (N_14774,N_13426,N_14157);
xor U14775 (N_14775,N_14272,N_13878);
nor U14776 (N_14776,N_13910,N_13748);
nor U14777 (N_14777,N_13628,N_13431);
nor U14778 (N_14778,N_14055,N_13963);
and U14779 (N_14779,N_13939,N_14224);
nor U14780 (N_14780,N_13580,N_13461);
xor U14781 (N_14781,N_13439,N_13286);
and U14782 (N_14782,N_13369,N_14106);
or U14783 (N_14783,N_13373,N_14324);
nand U14784 (N_14784,N_14214,N_13402);
nand U14785 (N_14785,N_13366,N_14373);
and U14786 (N_14786,N_13919,N_13711);
nor U14787 (N_14787,N_13756,N_13351);
xor U14788 (N_14788,N_14118,N_13830);
nand U14789 (N_14789,N_13797,N_14259);
nor U14790 (N_14790,N_14083,N_14236);
xor U14791 (N_14791,N_14311,N_13547);
nor U14792 (N_14792,N_13408,N_13357);
nor U14793 (N_14793,N_13761,N_13652);
nand U14794 (N_14794,N_13577,N_13765);
xor U14795 (N_14795,N_13304,N_13946);
xor U14796 (N_14796,N_13399,N_13417);
nand U14797 (N_14797,N_14273,N_13574);
or U14798 (N_14798,N_13297,N_13881);
or U14799 (N_14799,N_13218,N_14290);
and U14800 (N_14800,N_13918,N_14201);
xnor U14801 (N_14801,N_14072,N_13486);
nand U14802 (N_14802,N_13739,N_13635);
and U14803 (N_14803,N_13548,N_13799);
nand U14804 (N_14804,N_14182,N_13272);
nor U14805 (N_14805,N_13309,N_13638);
nand U14806 (N_14806,N_13266,N_13812);
or U14807 (N_14807,N_13610,N_14114);
or U14808 (N_14808,N_14199,N_13899);
nand U14809 (N_14809,N_13476,N_14216);
nand U14810 (N_14810,N_13682,N_14015);
nor U14811 (N_14811,N_13909,N_13555);
or U14812 (N_14812,N_14394,N_13204);
and U14813 (N_14813,N_14091,N_13308);
and U14814 (N_14814,N_13307,N_14385);
and U14815 (N_14815,N_14284,N_13842);
and U14816 (N_14816,N_13422,N_13624);
xnor U14817 (N_14817,N_13410,N_14247);
nand U14818 (N_14818,N_13654,N_14364);
or U14819 (N_14819,N_13630,N_14082);
or U14820 (N_14820,N_14393,N_13282);
and U14821 (N_14821,N_13991,N_13594);
nand U14822 (N_14822,N_13386,N_13225);
or U14823 (N_14823,N_13317,N_14181);
xnor U14824 (N_14824,N_13549,N_14303);
nand U14825 (N_14825,N_13854,N_14197);
nor U14826 (N_14826,N_13270,N_14143);
nor U14827 (N_14827,N_14281,N_13302);
or U14828 (N_14828,N_13769,N_13811);
nand U14829 (N_14829,N_13726,N_13521);
xor U14830 (N_14830,N_13237,N_13679);
xnor U14831 (N_14831,N_14066,N_13274);
or U14832 (N_14832,N_13230,N_14279);
nor U14833 (N_14833,N_14033,N_14280);
and U14834 (N_14834,N_13372,N_13794);
xnor U14835 (N_14835,N_14075,N_14362);
and U14836 (N_14836,N_14195,N_13598);
xor U14837 (N_14837,N_13993,N_13278);
nor U14838 (N_14838,N_14024,N_13564);
and U14839 (N_14839,N_13360,N_14192);
xor U14840 (N_14840,N_14021,N_13688);
or U14841 (N_14841,N_13767,N_13696);
xor U14842 (N_14842,N_13432,N_13858);
nand U14843 (N_14843,N_14189,N_13315);
nand U14844 (N_14844,N_13292,N_13953);
or U14845 (N_14845,N_14012,N_13757);
nor U14846 (N_14846,N_14152,N_13951);
and U14847 (N_14847,N_13664,N_13281);
xor U14848 (N_14848,N_13503,N_14360);
xor U14849 (N_14849,N_13680,N_13345);
nand U14850 (N_14850,N_13813,N_13223);
nor U14851 (N_14851,N_13692,N_14110);
xnor U14852 (N_14852,N_14381,N_13647);
and U14853 (N_14853,N_13779,N_13471);
and U14854 (N_14854,N_13465,N_13911);
and U14855 (N_14855,N_13935,N_13841);
or U14856 (N_14856,N_13398,N_14007);
nor U14857 (N_14857,N_13285,N_14325);
and U14858 (N_14858,N_14365,N_14160);
and U14859 (N_14859,N_14039,N_13869);
nor U14860 (N_14860,N_14287,N_13414);
nand U14861 (N_14861,N_13847,N_14144);
xor U14862 (N_14862,N_13236,N_14219);
or U14863 (N_14863,N_14370,N_14063);
and U14864 (N_14864,N_14368,N_14031);
and U14865 (N_14865,N_14267,N_13928);
or U14866 (N_14866,N_13856,N_13808);
xnor U14867 (N_14867,N_13619,N_13209);
or U14868 (N_14868,N_14138,N_13248);
nand U14869 (N_14869,N_13496,N_14108);
or U14870 (N_14870,N_14344,N_13902);
nand U14871 (N_14871,N_13987,N_14164);
xnor U14872 (N_14872,N_13718,N_13244);
or U14873 (N_14873,N_13903,N_13600);
or U14874 (N_14874,N_13895,N_13301);
nand U14875 (N_14875,N_13685,N_13251);
and U14876 (N_14876,N_13668,N_13536);
nand U14877 (N_14877,N_13252,N_14112);
and U14878 (N_14878,N_13552,N_14374);
xor U14879 (N_14879,N_13467,N_13356);
and U14880 (N_14880,N_13807,N_13831);
xor U14881 (N_14881,N_13420,N_13785);
xor U14882 (N_14882,N_13880,N_14070);
or U14883 (N_14883,N_13239,N_13744);
or U14884 (N_14884,N_13511,N_13925);
and U14885 (N_14885,N_13723,N_14147);
nand U14886 (N_14886,N_13537,N_14221);
nand U14887 (N_14887,N_13627,N_14326);
xnor U14888 (N_14888,N_13689,N_13474);
or U14889 (N_14889,N_13760,N_14335);
nand U14890 (N_14890,N_13737,N_14357);
and U14891 (N_14891,N_13455,N_14295);
and U14892 (N_14892,N_13498,N_13714);
xor U14893 (N_14893,N_13575,N_13730);
nor U14894 (N_14894,N_13862,N_14180);
or U14895 (N_14895,N_13912,N_13557);
nand U14896 (N_14896,N_13527,N_13921);
nand U14897 (N_14897,N_13832,N_14371);
nand U14898 (N_14898,N_13220,N_13937);
nand U14899 (N_14899,N_13956,N_14317);
nand U14900 (N_14900,N_14131,N_13383);
nor U14901 (N_14901,N_14141,N_14378);
and U14902 (N_14902,N_14312,N_13247);
xor U14903 (N_14903,N_13262,N_13900);
or U14904 (N_14904,N_13545,N_13201);
xor U14905 (N_14905,N_13516,N_13690);
nor U14906 (N_14906,N_13738,N_13374);
xor U14907 (N_14907,N_14067,N_13288);
or U14908 (N_14908,N_13675,N_13996);
or U14909 (N_14909,N_13328,N_14391);
or U14910 (N_14910,N_13915,N_13229);
or U14911 (N_14911,N_13540,N_13400);
and U14912 (N_14912,N_13440,N_13851);
nor U14913 (N_14913,N_13876,N_13475);
nor U14914 (N_14914,N_13926,N_14092);
nand U14915 (N_14915,N_13795,N_14350);
or U14916 (N_14916,N_13676,N_13650);
or U14917 (N_14917,N_13693,N_13353);
xor U14918 (N_14918,N_13618,N_14010);
nor U14919 (N_14919,N_13277,N_13451);
nor U14920 (N_14920,N_13216,N_14264);
xor U14921 (N_14921,N_14084,N_14123);
nor U14922 (N_14922,N_13674,N_14126);
or U14923 (N_14923,N_13316,N_14029);
or U14924 (N_14924,N_14088,N_13535);
xor U14925 (N_14925,N_14185,N_13863);
nand U14926 (N_14926,N_13275,N_13709);
xnor U14927 (N_14927,N_13246,N_13959);
and U14928 (N_14928,N_13298,N_13267);
or U14929 (N_14929,N_13633,N_13655);
nor U14930 (N_14930,N_13796,N_14107);
nand U14931 (N_14931,N_14359,N_13202);
nand U14932 (N_14932,N_13729,N_13273);
or U14933 (N_14933,N_13279,N_13623);
nand U14934 (N_14934,N_13822,N_13874);
or U14935 (N_14935,N_14243,N_13350);
or U14936 (N_14936,N_14242,N_14309);
xnor U14937 (N_14937,N_14252,N_14159);
xnor U14938 (N_14938,N_13845,N_13551);
xor U14939 (N_14939,N_13276,N_14386);
nor U14940 (N_14940,N_13759,N_14274);
and U14941 (N_14941,N_13828,N_13764);
nor U14942 (N_14942,N_13731,N_13446);
xnor U14943 (N_14943,N_13994,N_14323);
nor U14944 (N_14944,N_13662,N_14220);
xnor U14945 (N_14945,N_13573,N_13559);
xor U14946 (N_14946,N_14296,N_13234);
or U14947 (N_14947,N_13478,N_13678);
xor U14948 (N_14948,N_14149,N_14240);
nor U14949 (N_14949,N_14286,N_13649);
nand U14950 (N_14950,N_13774,N_13597);
nor U14951 (N_14951,N_13589,N_13805);
and U14952 (N_14952,N_14358,N_13342);
nor U14953 (N_14953,N_13865,N_13837);
nand U14954 (N_14954,N_13892,N_14292);
nor U14955 (N_14955,N_13605,N_13740);
or U14956 (N_14956,N_14018,N_14150);
and U14957 (N_14957,N_13971,N_13263);
nand U14958 (N_14958,N_13254,N_13424);
or U14959 (N_14959,N_13978,N_13437);
and U14960 (N_14960,N_13943,N_14124);
nand U14961 (N_14961,N_14283,N_13388);
nor U14962 (N_14962,N_14027,N_13506);
nor U14963 (N_14963,N_13631,N_14315);
or U14964 (N_14964,N_14268,N_14226);
xor U14965 (N_14965,N_13359,N_13934);
xor U14966 (N_14966,N_13294,N_14096);
or U14967 (N_14967,N_14271,N_13289);
and U14968 (N_14968,N_13499,N_13772);
nand U14969 (N_14969,N_13462,N_13975);
nor U14970 (N_14970,N_14289,N_13406);
and U14971 (N_14971,N_13329,N_13532);
xor U14972 (N_14972,N_13694,N_13798);
nor U14973 (N_14973,N_14249,N_13601);
nor U14974 (N_14974,N_13364,N_13392);
or U14975 (N_14975,N_13673,N_14097);
nor U14976 (N_14976,N_13566,N_13940);
or U14977 (N_14977,N_13867,N_13728);
nor U14978 (N_14978,N_14153,N_13870);
xor U14979 (N_14979,N_13944,N_13271);
nand U14980 (N_14980,N_14241,N_13415);
nor U14981 (N_14981,N_13768,N_13640);
or U14982 (N_14982,N_13875,N_13256);
nand U14983 (N_14983,N_13525,N_14347);
nor U14984 (N_14984,N_14269,N_13644);
and U14985 (N_14985,N_13567,N_13979);
xor U14986 (N_14986,N_13510,N_13998);
and U14987 (N_14987,N_14332,N_13791);
or U14988 (N_14988,N_14001,N_13382);
nand U14989 (N_14989,N_14059,N_13389);
and U14990 (N_14990,N_13922,N_13250);
nor U14991 (N_14991,N_13326,N_13782);
or U14992 (N_14992,N_14304,N_13484);
and U14993 (N_14993,N_13893,N_13320);
nor U14994 (N_14994,N_13885,N_14369);
or U14995 (N_14995,N_14395,N_13291);
nor U14996 (N_14996,N_14246,N_13562);
and U14997 (N_14997,N_13570,N_13585);
nand U14998 (N_14998,N_13569,N_14307);
or U14999 (N_14999,N_13387,N_14081);
and U15000 (N_15000,N_14089,N_13982);
xnor U15001 (N_15001,N_13405,N_13351);
and U15002 (N_15002,N_13785,N_13888);
and U15003 (N_15003,N_14112,N_13583);
nor U15004 (N_15004,N_13712,N_14050);
xnor U15005 (N_15005,N_13290,N_14035);
or U15006 (N_15006,N_13475,N_14310);
nor U15007 (N_15007,N_13301,N_13869);
or U15008 (N_15008,N_14264,N_13940);
or U15009 (N_15009,N_13437,N_14168);
nor U15010 (N_15010,N_13550,N_13813);
or U15011 (N_15011,N_14377,N_14116);
nor U15012 (N_15012,N_13382,N_14356);
xnor U15013 (N_15013,N_14209,N_13317);
and U15014 (N_15014,N_14165,N_14004);
nand U15015 (N_15015,N_13620,N_13780);
xnor U15016 (N_15016,N_14247,N_13997);
xnor U15017 (N_15017,N_14246,N_14323);
nor U15018 (N_15018,N_13530,N_13290);
xor U15019 (N_15019,N_13497,N_13347);
and U15020 (N_15020,N_14063,N_14243);
and U15021 (N_15021,N_13861,N_13646);
and U15022 (N_15022,N_14018,N_13844);
nand U15023 (N_15023,N_13726,N_14193);
xor U15024 (N_15024,N_13660,N_13950);
nor U15025 (N_15025,N_13940,N_14043);
nand U15026 (N_15026,N_13279,N_14329);
or U15027 (N_15027,N_13387,N_13530);
and U15028 (N_15028,N_13590,N_13405);
xor U15029 (N_15029,N_13657,N_13533);
nor U15030 (N_15030,N_13519,N_13733);
nand U15031 (N_15031,N_13537,N_14066);
nor U15032 (N_15032,N_14014,N_13478);
or U15033 (N_15033,N_13486,N_13942);
nor U15034 (N_15034,N_13891,N_14057);
xnor U15035 (N_15035,N_14091,N_13546);
nand U15036 (N_15036,N_13295,N_14175);
xor U15037 (N_15037,N_14110,N_13372);
nand U15038 (N_15038,N_14284,N_13569);
or U15039 (N_15039,N_13230,N_13450);
and U15040 (N_15040,N_13983,N_13843);
or U15041 (N_15041,N_13607,N_13216);
or U15042 (N_15042,N_14032,N_14331);
and U15043 (N_15043,N_13307,N_14015);
xor U15044 (N_15044,N_13293,N_13688);
or U15045 (N_15045,N_13583,N_13554);
nor U15046 (N_15046,N_13576,N_13569);
xor U15047 (N_15047,N_13837,N_14362);
nand U15048 (N_15048,N_14058,N_13416);
nand U15049 (N_15049,N_14105,N_13897);
xnor U15050 (N_15050,N_13216,N_13217);
and U15051 (N_15051,N_13690,N_14142);
nor U15052 (N_15052,N_13492,N_14170);
xnor U15053 (N_15053,N_14050,N_13410);
and U15054 (N_15054,N_13331,N_14335);
or U15055 (N_15055,N_14375,N_13963);
xor U15056 (N_15056,N_14075,N_13834);
and U15057 (N_15057,N_13532,N_13829);
nand U15058 (N_15058,N_13384,N_13606);
xor U15059 (N_15059,N_14324,N_13526);
nand U15060 (N_15060,N_14218,N_13400);
nor U15061 (N_15061,N_14088,N_14379);
xor U15062 (N_15062,N_13776,N_14205);
nand U15063 (N_15063,N_14280,N_13665);
or U15064 (N_15064,N_13558,N_13499);
or U15065 (N_15065,N_14245,N_13236);
or U15066 (N_15066,N_13297,N_13845);
nor U15067 (N_15067,N_13638,N_13352);
nor U15068 (N_15068,N_13676,N_14018);
nor U15069 (N_15069,N_14217,N_13945);
nand U15070 (N_15070,N_13991,N_14371);
nand U15071 (N_15071,N_13672,N_13836);
nand U15072 (N_15072,N_13606,N_13633);
and U15073 (N_15073,N_14369,N_13309);
or U15074 (N_15074,N_14281,N_13647);
nor U15075 (N_15075,N_14061,N_13747);
nand U15076 (N_15076,N_14005,N_13295);
xor U15077 (N_15077,N_13680,N_14350);
and U15078 (N_15078,N_13831,N_13229);
or U15079 (N_15079,N_13428,N_14188);
or U15080 (N_15080,N_14288,N_13706);
nand U15081 (N_15081,N_14229,N_13421);
or U15082 (N_15082,N_13556,N_14237);
xor U15083 (N_15083,N_13578,N_14291);
nor U15084 (N_15084,N_13786,N_14363);
xor U15085 (N_15085,N_13325,N_13573);
and U15086 (N_15086,N_14006,N_13329);
nand U15087 (N_15087,N_13837,N_13925);
xnor U15088 (N_15088,N_14022,N_14246);
or U15089 (N_15089,N_14206,N_13545);
nor U15090 (N_15090,N_13415,N_13949);
nand U15091 (N_15091,N_14041,N_13893);
nor U15092 (N_15092,N_14146,N_13570);
xor U15093 (N_15093,N_13917,N_13568);
xnor U15094 (N_15094,N_13703,N_14219);
nand U15095 (N_15095,N_13696,N_13229);
and U15096 (N_15096,N_13442,N_13230);
and U15097 (N_15097,N_13900,N_14231);
xnor U15098 (N_15098,N_14023,N_13307);
nor U15099 (N_15099,N_13608,N_13364);
nand U15100 (N_15100,N_13850,N_14064);
xor U15101 (N_15101,N_14078,N_13417);
and U15102 (N_15102,N_14010,N_13759);
xor U15103 (N_15103,N_13421,N_13371);
nand U15104 (N_15104,N_14331,N_13604);
nand U15105 (N_15105,N_13716,N_14151);
nor U15106 (N_15106,N_13876,N_13286);
nor U15107 (N_15107,N_14388,N_13262);
xor U15108 (N_15108,N_14241,N_13522);
or U15109 (N_15109,N_13314,N_13418);
xnor U15110 (N_15110,N_14249,N_13883);
nand U15111 (N_15111,N_14023,N_13218);
xor U15112 (N_15112,N_13723,N_14273);
xor U15113 (N_15113,N_13299,N_13717);
and U15114 (N_15114,N_13890,N_13589);
or U15115 (N_15115,N_13211,N_13898);
or U15116 (N_15116,N_13874,N_13447);
or U15117 (N_15117,N_13676,N_13276);
or U15118 (N_15118,N_14395,N_14070);
nor U15119 (N_15119,N_14182,N_14206);
or U15120 (N_15120,N_13793,N_13943);
nor U15121 (N_15121,N_13698,N_14009);
nor U15122 (N_15122,N_13920,N_13312);
xnor U15123 (N_15123,N_13756,N_13692);
xor U15124 (N_15124,N_13746,N_13835);
nor U15125 (N_15125,N_14328,N_13243);
and U15126 (N_15126,N_13641,N_13760);
xnor U15127 (N_15127,N_14390,N_14225);
and U15128 (N_15128,N_14214,N_13417);
xor U15129 (N_15129,N_13761,N_13798);
nand U15130 (N_15130,N_13685,N_14169);
and U15131 (N_15131,N_13418,N_14071);
nor U15132 (N_15132,N_13831,N_13861);
or U15133 (N_15133,N_13307,N_13252);
nor U15134 (N_15134,N_13551,N_13704);
and U15135 (N_15135,N_13890,N_13278);
or U15136 (N_15136,N_14117,N_13675);
or U15137 (N_15137,N_13548,N_13327);
nand U15138 (N_15138,N_13751,N_13855);
nand U15139 (N_15139,N_14287,N_13745);
or U15140 (N_15140,N_13590,N_14188);
or U15141 (N_15141,N_13258,N_13793);
and U15142 (N_15142,N_13425,N_13478);
xnor U15143 (N_15143,N_13636,N_14047);
nor U15144 (N_15144,N_13486,N_13638);
or U15145 (N_15145,N_13303,N_13825);
nor U15146 (N_15146,N_14139,N_13977);
xnor U15147 (N_15147,N_13718,N_13851);
xor U15148 (N_15148,N_13374,N_14297);
xnor U15149 (N_15149,N_13530,N_13631);
xor U15150 (N_15150,N_14030,N_13822);
nand U15151 (N_15151,N_13795,N_13518);
xnor U15152 (N_15152,N_13442,N_14079);
xnor U15153 (N_15153,N_13996,N_13624);
and U15154 (N_15154,N_14279,N_13811);
nor U15155 (N_15155,N_13819,N_13994);
and U15156 (N_15156,N_14213,N_13775);
or U15157 (N_15157,N_13918,N_14365);
xnor U15158 (N_15158,N_13525,N_13763);
nor U15159 (N_15159,N_14304,N_13631);
and U15160 (N_15160,N_13388,N_14293);
nor U15161 (N_15161,N_13504,N_14295);
nor U15162 (N_15162,N_13758,N_13696);
xor U15163 (N_15163,N_13262,N_13919);
or U15164 (N_15164,N_13389,N_13520);
xnor U15165 (N_15165,N_13254,N_13793);
and U15166 (N_15166,N_13284,N_13452);
or U15167 (N_15167,N_13785,N_13679);
xor U15168 (N_15168,N_13806,N_14170);
xor U15169 (N_15169,N_14269,N_13972);
or U15170 (N_15170,N_14069,N_13266);
nand U15171 (N_15171,N_13954,N_13431);
or U15172 (N_15172,N_13720,N_13326);
nor U15173 (N_15173,N_13736,N_13978);
and U15174 (N_15174,N_13673,N_13864);
or U15175 (N_15175,N_14073,N_13954);
nor U15176 (N_15176,N_13982,N_13210);
or U15177 (N_15177,N_13510,N_13562);
and U15178 (N_15178,N_13633,N_13208);
and U15179 (N_15179,N_13806,N_13394);
xnor U15180 (N_15180,N_13286,N_13446);
nand U15181 (N_15181,N_13540,N_14375);
and U15182 (N_15182,N_14219,N_13233);
nor U15183 (N_15183,N_14273,N_14162);
or U15184 (N_15184,N_14019,N_13758);
nand U15185 (N_15185,N_14086,N_13424);
or U15186 (N_15186,N_14031,N_14077);
or U15187 (N_15187,N_13905,N_13782);
nor U15188 (N_15188,N_14192,N_13271);
nand U15189 (N_15189,N_13297,N_14046);
xor U15190 (N_15190,N_14137,N_13703);
or U15191 (N_15191,N_13323,N_13506);
and U15192 (N_15192,N_14039,N_13296);
xor U15193 (N_15193,N_14064,N_14266);
and U15194 (N_15194,N_14312,N_14130);
nand U15195 (N_15195,N_14298,N_13795);
nand U15196 (N_15196,N_13347,N_13858);
xor U15197 (N_15197,N_13275,N_14329);
nor U15198 (N_15198,N_13676,N_13353);
nor U15199 (N_15199,N_14318,N_13698);
xnor U15200 (N_15200,N_13513,N_13624);
nand U15201 (N_15201,N_13246,N_14300);
or U15202 (N_15202,N_13757,N_14254);
and U15203 (N_15203,N_13883,N_13924);
and U15204 (N_15204,N_13408,N_14009);
nor U15205 (N_15205,N_14197,N_13451);
or U15206 (N_15206,N_14361,N_13598);
or U15207 (N_15207,N_13538,N_14153);
or U15208 (N_15208,N_14304,N_13997);
and U15209 (N_15209,N_14371,N_13967);
nand U15210 (N_15210,N_13955,N_13840);
xor U15211 (N_15211,N_14398,N_13582);
or U15212 (N_15212,N_13724,N_13366);
and U15213 (N_15213,N_14016,N_14380);
or U15214 (N_15214,N_14116,N_13308);
or U15215 (N_15215,N_13326,N_13393);
and U15216 (N_15216,N_13656,N_14017);
or U15217 (N_15217,N_13702,N_13215);
and U15218 (N_15218,N_13861,N_13407);
nor U15219 (N_15219,N_13525,N_13245);
nor U15220 (N_15220,N_14039,N_14098);
nor U15221 (N_15221,N_13875,N_14306);
or U15222 (N_15222,N_13665,N_13261);
or U15223 (N_15223,N_14192,N_13973);
or U15224 (N_15224,N_13623,N_14357);
and U15225 (N_15225,N_13462,N_14080);
nand U15226 (N_15226,N_13230,N_13214);
xnor U15227 (N_15227,N_13399,N_13878);
nand U15228 (N_15228,N_14117,N_13315);
nor U15229 (N_15229,N_13283,N_13618);
xor U15230 (N_15230,N_13821,N_13534);
nand U15231 (N_15231,N_14024,N_13994);
xor U15232 (N_15232,N_13581,N_13535);
nand U15233 (N_15233,N_14308,N_13596);
or U15234 (N_15234,N_14264,N_13879);
or U15235 (N_15235,N_13883,N_14018);
nand U15236 (N_15236,N_13429,N_13242);
xnor U15237 (N_15237,N_13864,N_14300);
nand U15238 (N_15238,N_13301,N_13605);
nor U15239 (N_15239,N_13803,N_14357);
xor U15240 (N_15240,N_14117,N_14007);
and U15241 (N_15241,N_13569,N_13691);
xnor U15242 (N_15242,N_13887,N_14032);
nor U15243 (N_15243,N_13976,N_14010);
xor U15244 (N_15244,N_14247,N_13352);
xor U15245 (N_15245,N_13773,N_13344);
nor U15246 (N_15246,N_13835,N_13217);
nor U15247 (N_15247,N_13660,N_14236);
or U15248 (N_15248,N_13661,N_13419);
or U15249 (N_15249,N_13961,N_13560);
nand U15250 (N_15250,N_13533,N_13371);
nand U15251 (N_15251,N_13924,N_13771);
nand U15252 (N_15252,N_13558,N_14082);
or U15253 (N_15253,N_13859,N_14346);
nand U15254 (N_15254,N_13521,N_13371);
or U15255 (N_15255,N_13770,N_13708);
and U15256 (N_15256,N_14327,N_13811);
and U15257 (N_15257,N_13638,N_13772);
nor U15258 (N_15258,N_13363,N_13350);
xor U15259 (N_15259,N_14206,N_14040);
nor U15260 (N_15260,N_13755,N_13909);
and U15261 (N_15261,N_14247,N_13989);
xor U15262 (N_15262,N_13213,N_13263);
and U15263 (N_15263,N_13744,N_13352);
and U15264 (N_15264,N_14207,N_13979);
or U15265 (N_15265,N_13870,N_13368);
xnor U15266 (N_15266,N_13549,N_13830);
nor U15267 (N_15267,N_13315,N_13286);
nor U15268 (N_15268,N_13954,N_14212);
xor U15269 (N_15269,N_13938,N_14239);
and U15270 (N_15270,N_13759,N_13753);
nor U15271 (N_15271,N_13485,N_13567);
or U15272 (N_15272,N_13318,N_13299);
or U15273 (N_15273,N_14304,N_13723);
nand U15274 (N_15274,N_13602,N_13546);
nand U15275 (N_15275,N_13708,N_14085);
xnor U15276 (N_15276,N_14341,N_13307);
or U15277 (N_15277,N_13748,N_13432);
or U15278 (N_15278,N_14050,N_13784);
nand U15279 (N_15279,N_13376,N_14130);
xor U15280 (N_15280,N_13242,N_13316);
and U15281 (N_15281,N_13895,N_14394);
nand U15282 (N_15282,N_13472,N_13303);
or U15283 (N_15283,N_13316,N_13569);
or U15284 (N_15284,N_13604,N_13727);
and U15285 (N_15285,N_13359,N_14269);
or U15286 (N_15286,N_13200,N_14070);
nor U15287 (N_15287,N_13653,N_14057);
or U15288 (N_15288,N_13478,N_13842);
xor U15289 (N_15289,N_13794,N_14097);
nor U15290 (N_15290,N_13944,N_13410);
or U15291 (N_15291,N_13348,N_14084);
nor U15292 (N_15292,N_14115,N_13485);
and U15293 (N_15293,N_13370,N_13316);
nor U15294 (N_15294,N_14075,N_13939);
and U15295 (N_15295,N_14390,N_13593);
or U15296 (N_15296,N_13790,N_13400);
nand U15297 (N_15297,N_14350,N_13219);
nor U15298 (N_15298,N_14037,N_14150);
nor U15299 (N_15299,N_14184,N_13699);
or U15300 (N_15300,N_13247,N_13384);
nor U15301 (N_15301,N_13956,N_13585);
nand U15302 (N_15302,N_13418,N_14232);
nand U15303 (N_15303,N_13988,N_13911);
and U15304 (N_15304,N_14268,N_13961);
xor U15305 (N_15305,N_13360,N_14131);
xor U15306 (N_15306,N_13671,N_13817);
nor U15307 (N_15307,N_13622,N_13401);
xnor U15308 (N_15308,N_14341,N_13431);
and U15309 (N_15309,N_14158,N_13430);
nor U15310 (N_15310,N_14037,N_14044);
and U15311 (N_15311,N_13776,N_13346);
nand U15312 (N_15312,N_14310,N_13579);
or U15313 (N_15313,N_13833,N_14237);
nand U15314 (N_15314,N_13401,N_13254);
xnor U15315 (N_15315,N_13937,N_13668);
or U15316 (N_15316,N_13847,N_14182);
nor U15317 (N_15317,N_14001,N_13798);
and U15318 (N_15318,N_13899,N_13261);
nand U15319 (N_15319,N_13464,N_13981);
xor U15320 (N_15320,N_14171,N_14187);
xnor U15321 (N_15321,N_13253,N_13767);
nand U15322 (N_15322,N_13477,N_13231);
and U15323 (N_15323,N_14319,N_14168);
xor U15324 (N_15324,N_13217,N_14189);
nand U15325 (N_15325,N_14126,N_13913);
nor U15326 (N_15326,N_13844,N_13575);
xnor U15327 (N_15327,N_13513,N_13570);
xor U15328 (N_15328,N_13959,N_13996);
xnor U15329 (N_15329,N_14236,N_14027);
xnor U15330 (N_15330,N_13417,N_13477);
nor U15331 (N_15331,N_13628,N_14045);
nor U15332 (N_15332,N_13733,N_13420);
xor U15333 (N_15333,N_13953,N_14263);
and U15334 (N_15334,N_13999,N_13970);
or U15335 (N_15335,N_14385,N_13516);
nor U15336 (N_15336,N_13898,N_13382);
nor U15337 (N_15337,N_13327,N_13590);
nor U15338 (N_15338,N_14150,N_13302);
xor U15339 (N_15339,N_13689,N_13366);
nor U15340 (N_15340,N_13784,N_13262);
and U15341 (N_15341,N_14180,N_13762);
and U15342 (N_15342,N_13766,N_14039);
xor U15343 (N_15343,N_13420,N_13457);
and U15344 (N_15344,N_14211,N_13361);
xnor U15345 (N_15345,N_14128,N_13824);
nand U15346 (N_15346,N_13538,N_13805);
nand U15347 (N_15347,N_13483,N_14279);
and U15348 (N_15348,N_13753,N_13345);
or U15349 (N_15349,N_14154,N_14179);
nor U15350 (N_15350,N_14227,N_13290);
nand U15351 (N_15351,N_14351,N_14136);
nor U15352 (N_15352,N_13309,N_14262);
and U15353 (N_15353,N_13890,N_13938);
and U15354 (N_15354,N_13802,N_13321);
and U15355 (N_15355,N_14206,N_14289);
nor U15356 (N_15356,N_14320,N_14358);
nor U15357 (N_15357,N_13441,N_14235);
or U15358 (N_15358,N_13689,N_13218);
xor U15359 (N_15359,N_13555,N_13414);
xnor U15360 (N_15360,N_14070,N_14306);
xor U15361 (N_15361,N_14154,N_13796);
nor U15362 (N_15362,N_13293,N_13457);
nor U15363 (N_15363,N_14307,N_13627);
nand U15364 (N_15364,N_13489,N_14050);
nor U15365 (N_15365,N_13527,N_13996);
and U15366 (N_15366,N_13530,N_13678);
xnor U15367 (N_15367,N_13504,N_13858);
nor U15368 (N_15368,N_13876,N_13854);
or U15369 (N_15369,N_13225,N_13369);
xnor U15370 (N_15370,N_14224,N_14219);
xnor U15371 (N_15371,N_14343,N_14147);
or U15372 (N_15372,N_13940,N_14327);
and U15373 (N_15373,N_13955,N_13279);
nand U15374 (N_15374,N_14222,N_13886);
or U15375 (N_15375,N_13330,N_14110);
xor U15376 (N_15376,N_13502,N_14047);
nand U15377 (N_15377,N_14064,N_13436);
nor U15378 (N_15378,N_13271,N_13779);
nand U15379 (N_15379,N_13221,N_14156);
xor U15380 (N_15380,N_13275,N_14044);
xor U15381 (N_15381,N_13725,N_13653);
xnor U15382 (N_15382,N_13549,N_14275);
nand U15383 (N_15383,N_14285,N_14080);
xnor U15384 (N_15384,N_14012,N_13423);
xnor U15385 (N_15385,N_14285,N_13850);
nand U15386 (N_15386,N_14384,N_14231);
nor U15387 (N_15387,N_14339,N_13958);
xor U15388 (N_15388,N_14336,N_13476);
nand U15389 (N_15389,N_14069,N_13602);
nor U15390 (N_15390,N_13229,N_13493);
nor U15391 (N_15391,N_13494,N_13205);
and U15392 (N_15392,N_13516,N_13877);
or U15393 (N_15393,N_13611,N_13573);
nand U15394 (N_15394,N_13653,N_14181);
or U15395 (N_15395,N_13337,N_13233);
and U15396 (N_15396,N_13993,N_13464);
xnor U15397 (N_15397,N_13234,N_13856);
nand U15398 (N_15398,N_13547,N_13828);
and U15399 (N_15399,N_13379,N_14218);
or U15400 (N_15400,N_14226,N_14335);
and U15401 (N_15401,N_13611,N_13218);
xor U15402 (N_15402,N_13966,N_13772);
nand U15403 (N_15403,N_13544,N_14306);
and U15404 (N_15404,N_14299,N_14046);
and U15405 (N_15405,N_13575,N_14002);
xor U15406 (N_15406,N_13890,N_14238);
or U15407 (N_15407,N_13884,N_13917);
or U15408 (N_15408,N_13776,N_13737);
or U15409 (N_15409,N_13910,N_14238);
nor U15410 (N_15410,N_13407,N_13419);
xor U15411 (N_15411,N_14121,N_14345);
or U15412 (N_15412,N_13264,N_13218);
nand U15413 (N_15413,N_13233,N_13333);
xor U15414 (N_15414,N_13727,N_13728);
nand U15415 (N_15415,N_14258,N_13899);
and U15416 (N_15416,N_13560,N_14010);
xnor U15417 (N_15417,N_14141,N_13508);
and U15418 (N_15418,N_13813,N_13486);
and U15419 (N_15419,N_13590,N_13308);
nand U15420 (N_15420,N_14240,N_14363);
xor U15421 (N_15421,N_14091,N_13600);
or U15422 (N_15422,N_14177,N_14168);
nor U15423 (N_15423,N_13392,N_13546);
or U15424 (N_15424,N_13956,N_13338);
or U15425 (N_15425,N_14154,N_13938);
nand U15426 (N_15426,N_14067,N_13222);
and U15427 (N_15427,N_13707,N_13743);
or U15428 (N_15428,N_13480,N_14044);
nor U15429 (N_15429,N_14064,N_13387);
or U15430 (N_15430,N_13426,N_13316);
nand U15431 (N_15431,N_14222,N_13922);
nand U15432 (N_15432,N_13925,N_14213);
and U15433 (N_15433,N_13523,N_13508);
nand U15434 (N_15434,N_13644,N_13509);
nand U15435 (N_15435,N_13454,N_14242);
or U15436 (N_15436,N_13625,N_14257);
nor U15437 (N_15437,N_13393,N_14141);
nor U15438 (N_15438,N_14049,N_13610);
and U15439 (N_15439,N_14111,N_13750);
or U15440 (N_15440,N_13287,N_13311);
and U15441 (N_15441,N_14180,N_13619);
nor U15442 (N_15442,N_14354,N_13679);
nor U15443 (N_15443,N_13743,N_13660);
or U15444 (N_15444,N_13794,N_13371);
xnor U15445 (N_15445,N_13405,N_13338);
nor U15446 (N_15446,N_13723,N_13540);
xor U15447 (N_15447,N_13523,N_13565);
or U15448 (N_15448,N_14294,N_13804);
and U15449 (N_15449,N_13693,N_14185);
or U15450 (N_15450,N_13276,N_13513);
or U15451 (N_15451,N_13901,N_13458);
and U15452 (N_15452,N_13251,N_14055);
nor U15453 (N_15453,N_14070,N_13717);
nor U15454 (N_15454,N_13494,N_13920);
or U15455 (N_15455,N_14289,N_13477);
nor U15456 (N_15456,N_14084,N_14194);
xor U15457 (N_15457,N_13806,N_13396);
nor U15458 (N_15458,N_13835,N_13873);
or U15459 (N_15459,N_14311,N_14194);
and U15460 (N_15460,N_14332,N_13571);
or U15461 (N_15461,N_14285,N_13456);
and U15462 (N_15462,N_13258,N_13700);
nor U15463 (N_15463,N_14384,N_13886);
xnor U15464 (N_15464,N_13583,N_13931);
and U15465 (N_15465,N_13250,N_13213);
nor U15466 (N_15466,N_13411,N_14016);
xor U15467 (N_15467,N_14212,N_14152);
and U15468 (N_15468,N_13224,N_14001);
nor U15469 (N_15469,N_13712,N_14094);
xnor U15470 (N_15470,N_13917,N_14050);
nor U15471 (N_15471,N_14329,N_13819);
xor U15472 (N_15472,N_13615,N_13431);
and U15473 (N_15473,N_14170,N_13947);
xnor U15474 (N_15474,N_14339,N_14159);
or U15475 (N_15475,N_14086,N_13251);
nand U15476 (N_15476,N_14366,N_14089);
nand U15477 (N_15477,N_14140,N_13634);
xnor U15478 (N_15478,N_13556,N_14140);
or U15479 (N_15479,N_13633,N_14234);
xnor U15480 (N_15480,N_13626,N_14196);
nor U15481 (N_15481,N_14125,N_13759);
xnor U15482 (N_15482,N_13373,N_13492);
and U15483 (N_15483,N_13607,N_14290);
or U15484 (N_15484,N_13847,N_13357);
nor U15485 (N_15485,N_14248,N_13483);
xnor U15486 (N_15486,N_14105,N_13958);
or U15487 (N_15487,N_13923,N_13618);
and U15488 (N_15488,N_13954,N_14082);
and U15489 (N_15489,N_14375,N_13553);
or U15490 (N_15490,N_13964,N_13757);
or U15491 (N_15491,N_13781,N_13227);
xnor U15492 (N_15492,N_14297,N_14028);
and U15493 (N_15493,N_13802,N_13528);
and U15494 (N_15494,N_13985,N_14194);
and U15495 (N_15495,N_14160,N_13443);
or U15496 (N_15496,N_13963,N_14127);
xnor U15497 (N_15497,N_13711,N_13818);
and U15498 (N_15498,N_14209,N_13674);
nand U15499 (N_15499,N_13657,N_14017);
or U15500 (N_15500,N_14280,N_14099);
or U15501 (N_15501,N_14206,N_13609);
nor U15502 (N_15502,N_13953,N_13411);
nand U15503 (N_15503,N_13591,N_13685);
nand U15504 (N_15504,N_14146,N_13760);
or U15505 (N_15505,N_13482,N_14031);
or U15506 (N_15506,N_13283,N_13973);
xor U15507 (N_15507,N_14377,N_13334);
nand U15508 (N_15508,N_14142,N_13723);
and U15509 (N_15509,N_13364,N_13930);
or U15510 (N_15510,N_13493,N_14314);
nor U15511 (N_15511,N_13832,N_14318);
and U15512 (N_15512,N_13363,N_13532);
nand U15513 (N_15513,N_13668,N_13815);
and U15514 (N_15514,N_14137,N_14381);
xor U15515 (N_15515,N_13502,N_13681);
xnor U15516 (N_15516,N_13247,N_14330);
nor U15517 (N_15517,N_13811,N_13374);
or U15518 (N_15518,N_13336,N_14360);
nor U15519 (N_15519,N_13509,N_13259);
nand U15520 (N_15520,N_13546,N_14305);
nand U15521 (N_15521,N_14245,N_13379);
and U15522 (N_15522,N_13895,N_13844);
and U15523 (N_15523,N_13804,N_13769);
or U15524 (N_15524,N_14061,N_13611);
or U15525 (N_15525,N_14198,N_13550);
xnor U15526 (N_15526,N_13306,N_14011);
nand U15527 (N_15527,N_13957,N_13205);
and U15528 (N_15528,N_14111,N_13499);
and U15529 (N_15529,N_13987,N_14186);
xor U15530 (N_15530,N_13402,N_13369);
nand U15531 (N_15531,N_14050,N_14046);
and U15532 (N_15532,N_13557,N_14147);
nor U15533 (N_15533,N_13319,N_13536);
or U15534 (N_15534,N_13707,N_13428);
xnor U15535 (N_15535,N_14314,N_13736);
and U15536 (N_15536,N_13977,N_13753);
nor U15537 (N_15537,N_13272,N_13679);
nand U15538 (N_15538,N_14233,N_13406);
nand U15539 (N_15539,N_14376,N_14397);
or U15540 (N_15540,N_13800,N_13231);
and U15541 (N_15541,N_14247,N_13883);
or U15542 (N_15542,N_13618,N_13216);
nor U15543 (N_15543,N_13753,N_13878);
xor U15544 (N_15544,N_14334,N_14066);
nor U15545 (N_15545,N_13877,N_13490);
and U15546 (N_15546,N_13282,N_13672);
and U15547 (N_15547,N_14205,N_13931);
xor U15548 (N_15548,N_13526,N_14199);
and U15549 (N_15549,N_13486,N_13714);
nand U15550 (N_15550,N_14276,N_14050);
and U15551 (N_15551,N_14339,N_14288);
xnor U15552 (N_15552,N_13220,N_14306);
nand U15553 (N_15553,N_13849,N_13577);
nand U15554 (N_15554,N_13689,N_13370);
xnor U15555 (N_15555,N_13359,N_14037);
nand U15556 (N_15556,N_14222,N_13637);
or U15557 (N_15557,N_14316,N_14373);
or U15558 (N_15558,N_14052,N_13739);
or U15559 (N_15559,N_14327,N_13725);
nand U15560 (N_15560,N_13769,N_14270);
xnor U15561 (N_15561,N_13280,N_14278);
nand U15562 (N_15562,N_14129,N_14146);
nor U15563 (N_15563,N_13901,N_13648);
xor U15564 (N_15564,N_13775,N_14211);
or U15565 (N_15565,N_13606,N_14188);
nand U15566 (N_15566,N_13437,N_13449);
nor U15567 (N_15567,N_13824,N_13588);
or U15568 (N_15568,N_13594,N_14348);
xor U15569 (N_15569,N_14388,N_13650);
or U15570 (N_15570,N_14268,N_13697);
nor U15571 (N_15571,N_13445,N_13810);
nor U15572 (N_15572,N_13763,N_13655);
nor U15573 (N_15573,N_14358,N_13417);
xnor U15574 (N_15574,N_13200,N_13715);
xor U15575 (N_15575,N_14216,N_13480);
nor U15576 (N_15576,N_13751,N_13248);
and U15577 (N_15577,N_13377,N_13469);
or U15578 (N_15578,N_14373,N_13779);
or U15579 (N_15579,N_14054,N_13646);
nor U15580 (N_15580,N_13588,N_13497);
and U15581 (N_15581,N_13798,N_14346);
or U15582 (N_15582,N_13507,N_14181);
nand U15583 (N_15583,N_13761,N_13363);
and U15584 (N_15584,N_14025,N_13448);
xor U15585 (N_15585,N_14359,N_13776);
or U15586 (N_15586,N_13601,N_13965);
or U15587 (N_15587,N_13866,N_13971);
nor U15588 (N_15588,N_13513,N_13798);
nor U15589 (N_15589,N_14093,N_13438);
or U15590 (N_15590,N_14370,N_14231);
xnor U15591 (N_15591,N_14293,N_13825);
xor U15592 (N_15592,N_13239,N_14387);
nand U15593 (N_15593,N_13322,N_13664);
xnor U15594 (N_15594,N_14230,N_13759);
nor U15595 (N_15595,N_13768,N_13928);
xor U15596 (N_15596,N_13903,N_13635);
nand U15597 (N_15597,N_13888,N_13913);
or U15598 (N_15598,N_13932,N_13499);
xor U15599 (N_15599,N_14374,N_14324);
xnor U15600 (N_15600,N_14820,N_15460);
and U15601 (N_15601,N_14884,N_14644);
xnor U15602 (N_15602,N_15191,N_14710);
nand U15603 (N_15603,N_15379,N_14615);
or U15604 (N_15604,N_15344,N_15522);
xnor U15605 (N_15605,N_14446,N_14769);
and U15606 (N_15606,N_14704,N_14471);
or U15607 (N_15607,N_14583,N_14547);
xnor U15608 (N_15608,N_15197,N_14738);
and U15609 (N_15609,N_14431,N_15442);
nand U15610 (N_15610,N_14756,N_15001);
xor U15611 (N_15611,N_14826,N_15220);
or U15612 (N_15612,N_14876,N_14485);
nor U15613 (N_15613,N_15129,N_15260);
and U15614 (N_15614,N_15428,N_15541);
or U15615 (N_15615,N_14669,N_15340);
xor U15616 (N_15616,N_14605,N_15421);
and U15617 (N_15617,N_14722,N_14847);
nor U15618 (N_15618,N_14478,N_15560);
nor U15619 (N_15619,N_14652,N_15301);
nor U15620 (N_15620,N_14590,N_14842);
xor U15621 (N_15621,N_14527,N_14479);
nand U15622 (N_15622,N_14401,N_15273);
and U15623 (N_15623,N_15293,N_14683);
xor U15624 (N_15624,N_14767,N_15278);
xnor U15625 (N_15625,N_14708,N_15140);
or U15626 (N_15626,N_14855,N_15246);
or U15627 (N_15627,N_15350,N_15235);
or U15628 (N_15628,N_14544,N_15099);
or U15629 (N_15629,N_15586,N_14865);
and U15630 (N_15630,N_15389,N_15103);
nand U15631 (N_15631,N_15267,N_15020);
and U15632 (N_15632,N_14740,N_14895);
nand U15633 (N_15633,N_15162,N_15217);
nand U15634 (N_15634,N_14733,N_14435);
or U15635 (N_15635,N_15331,N_15531);
and U15636 (N_15636,N_14588,N_15381);
nand U15637 (N_15637,N_14966,N_15375);
xnor U15638 (N_15638,N_15582,N_14961);
nor U15639 (N_15639,N_15223,N_14405);
and U15640 (N_15640,N_14823,N_15313);
and U15641 (N_15641,N_15324,N_14506);
or U15642 (N_15642,N_15334,N_14711);
xor U15643 (N_15643,N_14635,N_15112);
and U15644 (N_15644,N_14808,N_14724);
nand U15645 (N_15645,N_15537,N_14627);
nand U15646 (N_15646,N_14452,N_15005);
xor U15647 (N_15647,N_15154,N_14620);
nor U15648 (N_15648,N_15006,N_14905);
and U15649 (N_15649,N_15370,N_14600);
or U15650 (N_15650,N_14940,N_14429);
nand U15651 (N_15651,N_14987,N_14534);
or U15652 (N_15652,N_14508,N_15115);
and U15653 (N_15653,N_14893,N_14954);
nand U15654 (N_15654,N_14480,N_15357);
nor U15655 (N_15655,N_15404,N_15050);
xor U15656 (N_15656,N_15161,N_15205);
xnor U15657 (N_15657,N_15319,N_15489);
nand U15658 (N_15658,N_15427,N_15320);
or U15659 (N_15659,N_15414,N_15349);
and U15660 (N_15660,N_14903,N_15144);
or U15661 (N_15661,N_15296,N_14696);
nand U15662 (N_15662,N_14771,N_14721);
nand U15663 (N_15663,N_14490,N_15336);
xnor U15664 (N_15664,N_14580,N_14688);
and U15665 (N_15665,N_14720,N_15596);
nand U15666 (N_15666,N_15086,N_14602);
nor U15667 (N_15667,N_15171,N_15533);
xor U15668 (N_15668,N_15432,N_14734);
xnor U15669 (N_15669,N_14542,N_15431);
nor U15670 (N_15670,N_15092,N_14586);
or U15671 (N_15671,N_14593,N_15568);
nand U15672 (N_15672,N_14845,N_15405);
and U15673 (N_15673,N_15031,N_15282);
or U15674 (N_15674,N_15277,N_14426);
or U15675 (N_15675,N_15315,N_14818);
xnor U15676 (N_15676,N_15048,N_15231);
and U15677 (N_15677,N_14984,N_14629);
xnor U15678 (N_15678,N_14568,N_14481);
xor U15679 (N_15679,N_14877,N_14653);
and U15680 (N_15680,N_14904,N_14607);
xor U15681 (N_15681,N_15089,N_15206);
nor U15682 (N_15682,N_15594,N_14929);
nor U15683 (N_15683,N_14703,N_15169);
xor U15684 (N_15684,N_15581,N_14496);
xor U15685 (N_15685,N_15043,N_15034);
nand U15686 (N_15686,N_15555,N_15054);
xnor U15687 (N_15687,N_15148,N_15430);
xor U15688 (N_15688,N_15107,N_15532);
nand U15689 (N_15689,N_15036,N_14690);
or U15690 (N_15690,N_15438,N_14456);
nand U15691 (N_15691,N_14493,N_15348);
and U15692 (N_15692,N_15083,N_15425);
xor U15693 (N_15693,N_14817,N_15091);
nand U15694 (N_15694,N_15362,N_14854);
and U15695 (N_15695,N_15500,N_14535);
and U15696 (N_15696,N_15012,N_15396);
or U15697 (N_15697,N_14764,N_14870);
nor U15698 (N_15698,N_15367,N_14606);
nor U15699 (N_15699,N_14512,N_14744);
nor U15700 (N_15700,N_15024,N_14555);
or U15701 (N_15701,N_14746,N_15587);
and U15702 (N_15702,N_14623,N_14851);
nand U15703 (N_15703,N_15070,N_15076);
nand U15704 (N_15704,N_15519,N_14666);
and U15705 (N_15705,N_14751,N_14622);
and U15706 (N_15706,N_15420,N_15286);
nand U15707 (N_15707,N_15041,N_14505);
xnor U15708 (N_15708,N_15477,N_15482);
nor U15709 (N_15709,N_15047,N_14835);
nand U15710 (N_15710,N_15072,N_15310);
and U15711 (N_15711,N_14773,N_15157);
nor U15712 (N_15712,N_14483,N_15517);
xor U15713 (N_15713,N_15287,N_14799);
xor U15714 (N_15714,N_15548,N_15455);
xor U15715 (N_15715,N_14444,N_15291);
nor U15716 (N_15716,N_14858,N_15534);
xnor U15717 (N_15717,N_14420,N_15366);
or U15718 (N_15718,N_15285,N_14702);
nand U15719 (N_15719,N_15028,N_15377);
or U15720 (N_15720,N_15535,N_14766);
xor U15721 (N_15721,N_15272,N_15547);
or U15722 (N_15722,N_14924,N_14868);
or U15723 (N_15723,N_15074,N_15289);
or U15724 (N_15724,N_14960,N_15158);
or U15725 (N_15725,N_15569,N_15242);
nor U15726 (N_15726,N_15382,N_14783);
nand U15727 (N_15727,N_15193,N_14942);
and U15728 (N_15728,N_14457,N_14592);
or U15729 (N_15729,N_15199,N_14561);
nor U15730 (N_15730,N_15204,N_15451);
and U15731 (N_15731,N_15557,N_14890);
nand U15732 (N_15732,N_15003,N_15390);
xnor U15733 (N_15733,N_14927,N_15021);
or U15734 (N_15734,N_15599,N_15508);
nor U15735 (N_15735,N_15056,N_14828);
nor U15736 (N_15736,N_15338,N_14470);
xor U15737 (N_15737,N_14819,N_15280);
nor U15738 (N_15738,N_14687,N_15225);
nand U15739 (N_15739,N_15149,N_14413);
nor U15740 (N_15740,N_14665,N_14533);
xor U15741 (N_15741,N_15543,N_14912);
xor U15742 (N_15742,N_14827,N_15450);
and U15743 (N_15743,N_14609,N_15327);
or U15744 (N_15744,N_15514,N_15049);
nand U15745 (N_15745,N_15307,N_15393);
nor U15746 (N_15746,N_15251,N_14415);
xor U15747 (N_15747,N_15419,N_14936);
nor U15748 (N_15748,N_14680,N_14403);
xnor U15749 (N_15749,N_15398,N_14894);
nor U15750 (N_15750,N_15330,N_14944);
nand U15751 (N_15751,N_14811,N_14971);
and U15752 (N_15752,N_15440,N_14735);
nor U15753 (N_15753,N_14423,N_15448);
nor U15754 (N_15754,N_14500,N_14739);
nor U15755 (N_15755,N_15247,N_14888);
and U15756 (N_15756,N_14805,N_15067);
or U15757 (N_15757,N_15332,N_14613);
and U15758 (N_15758,N_14775,N_14408);
nor U15759 (N_15759,N_14852,N_14539);
and U15760 (N_15760,N_14624,N_15170);
nor U15761 (N_15761,N_15088,N_14715);
or U15762 (N_15762,N_15011,N_15152);
nand U15763 (N_15763,N_14731,N_15406);
nand U15764 (N_15764,N_14474,N_15407);
nor U15765 (N_15765,N_15224,N_15521);
xor U15766 (N_15766,N_14917,N_15399);
nand U15767 (N_15767,N_15198,N_14673);
nor U15768 (N_15768,N_14667,N_15476);
nor U15769 (N_15769,N_14645,N_15556);
xnor U15770 (N_15770,N_14797,N_15059);
nand U15771 (N_15771,N_14430,N_15464);
or U15772 (N_15772,N_14492,N_15134);
nand U15773 (N_15773,N_14909,N_14840);
and U15774 (N_15774,N_15490,N_14445);
or U15775 (N_15775,N_15025,N_15459);
or U15776 (N_15776,N_14642,N_15417);
nor U15777 (N_15777,N_15497,N_15493);
or U15778 (N_15778,N_15068,N_15004);
nor U15779 (N_15779,N_14567,N_14857);
or U15780 (N_15780,N_15243,N_15228);
and U15781 (N_15781,N_15507,N_15387);
and U15782 (N_15782,N_15471,N_14685);
xnor U15783 (N_15783,N_14737,N_15110);
nand U15784 (N_15784,N_15567,N_14460);
nor U15785 (N_15785,N_14648,N_14689);
and U15786 (N_15786,N_14860,N_15299);
nand U15787 (N_15787,N_14869,N_14730);
or U15788 (N_15788,N_15312,N_14906);
nor U15789 (N_15789,N_14822,N_14639);
xnor U15790 (N_15790,N_15325,N_15426);
nor U15791 (N_15791,N_14864,N_15133);
or U15792 (N_15792,N_15055,N_15274);
and U15793 (N_15793,N_14617,N_14713);
nor U15794 (N_15794,N_14521,N_14848);
xnor U15795 (N_15795,N_14575,N_15119);
and U15796 (N_15796,N_14914,N_14548);
or U15797 (N_15797,N_14462,N_15027);
nand U15798 (N_15798,N_15187,N_14981);
nand U15799 (N_15799,N_15141,N_14947);
nand U15800 (N_15800,N_14650,N_15167);
or U15801 (N_15801,N_15098,N_14564);
or U15802 (N_15802,N_15104,N_14712);
nand U15803 (N_15803,N_14992,N_14990);
and U15804 (N_15804,N_15314,N_15499);
xor U15805 (N_15805,N_15253,N_14502);
nor U15806 (N_15806,N_14499,N_14755);
or U15807 (N_15807,N_15335,N_15178);
and U15808 (N_15808,N_15550,N_14861);
and U15809 (N_15809,N_15576,N_14867);
or U15810 (N_15810,N_14532,N_14576);
and U15811 (N_15811,N_14682,N_15589);
and U15812 (N_15812,N_15485,N_15265);
nand U15813 (N_15813,N_14886,N_14849);
or U15814 (N_15814,N_15392,N_14853);
and U15815 (N_15815,N_14803,N_15094);
and U15816 (N_15816,N_15565,N_14986);
and U15817 (N_15817,N_14824,N_15135);
and U15818 (N_15818,N_14946,N_14509);
and U15819 (N_15819,N_15013,N_14911);
nor U15820 (N_15820,N_14816,N_15216);
or U15821 (N_15821,N_15062,N_14427);
and U15822 (N_15822,N_15524,N_15174);
nor U15823 (N_15823,N_14786,N_14630);
nand U15824 (N_15824,N_15308,N_14638);
nor U15825 (N_15825,N_15269,N_15435);
xnor U15826 (N_15826,N_15413,N_15010);
and U15827 (N_15827,N_14441,N_15394);
nand U15828 (N_15828,N_14691,N_14809);
nand U15829 (N_15829,N_15304,N_14530);
nor U15830 (N_15830,N_15380,N_14464);
and U15831 (N_15831,N_14898,N_14443);
nand U15832 (N_15832,N_14684,N_15443);
xor U15833 (N_15833,N_14791,N_14418);
or U15834 (N_15834,N_15495,N_14804);
xor U15835 (N_15835,N_15343,N_15039);
and U15836 (N_15836,N_14616,N_14782);
or U15837 (N_15837,N_14973,N_14465);
or U15838 (N_15838,N_15040,N_15029);
and U15839 (N_15839,N_15258,N_15529);
nand U15840 (N_15840,N_14422,N_14697);
or U15841 (N_15841,N_14979,N_15468);
xor U15842 (N_15842,N_14969,N_15552);
nor U15843 (N_15843,N_14553,N_15172);
or U15844 (N_15844,N_14436,N_15069);
nand U15845 (N_15845,N_15237,N_15329);
or U15846 (N_15846,N_14473,N_14439);
or U15847 (N_15847,N_15182,N_15361);
and U15848 (N_15848,N_14748,N_14656);
nor U15849 (N_15849,N_14993,N_15470);
or U15850 (N_15850,N_15026,N_14813);
nand U15851 (N_15851,N_15369,N_15570);
xor U15852 (N_15852,N_15118,N_14424);
or U15853 (N_15853,N_15147,N_15573);
nor U15854 (N_15854,N_15143,N_15388);
nand U15855 (N_15855,N_15395,N_15288);
and U15856 (N_15856,N_14798,N_15322);
and U15857 (N_15857,N_14806,N_15108);
xnor U15858 (N_15858,N_15252,N_15064);
and U15859 (N_15859,N_15057,N_15527);
nor U15860 (N_15860,N_14700,N_15590);
and U15861 (N_15861,N_14599,N_14821);
or U15862 (N_15862,N_14698,N_15592);
nor U15863 (N_15863,N_14693,N_14515);
nand U15864 (N_15864,N_15202,N_15544);
or U15865 (N_15865,N_14559,N_14589);
nor U15866 (N_15866,N_14566,N_15058);
nor U15867 (N_15867,N_15297,N_15512);
nor U15868 (N_15868,N_14922,N_14726);
or U15869 (N_15869,N_15101,N_14603);
nor U15870 (N_15870,N_14651,N_15368);
nand U15871 (N_15871,N_14701,N_14511);
nand U15872 (N_15872,N_15422,N_14625);
nand U15873 (N_15873,N_14777,N_15408);
nand U15874 (N_15874,N_15444,N_14663);
and U15875 (N_15875,N_14763,N_14438);
or U15876 (N_15876,N_14972,N_15106);
nand U15877 (N_15877,N_14707,N_14582);
xor U15878 (N_15878,N_14692,N_15096);
xnor U15879 (N_15879,N_14646,N_15015);
nand U15880 (N_15880,N_14794,N_14581);
nor U15881 (N_15881,N_14482,N_14531);
and U15882 (N_15882,N_14846,N_14409);
and U15883 (N_15883,N_15479,N_14432);
and U15884 (N_15884,N_14999,N_14779);
nor U15885 (N_15885,N_14611,N_14448);
or U15886 (N_15886,N_14621,N_15097);
nand U15887 (N_15887,N_15341,N_15233);
nor U15888 (N_15888,N_14519,N_15211);
xor U15889 (N_15889,N_15276,N_14983);
or U15890 (N_15890,N_14654,N_14404);
nor U15891 (N_15891,N_14612,N_15415);
or U15892 (N_15892,N_15542,N_14836);
xnor U15893 (N_15893,N_15100,N_14543);
or U15894 (N_15894,N_14610,N_15510);
or U15895 (N_15895,N_14565,N_14887);
nor U15896 (N_15896,N_15078,N_14699);
nand U15897 (N_15897,N_15401,N_15077);
nor U15898 (N_15898,N_14552,N_15292);
or U15899 (N_15899,N_15463,N_15084);
nand U15900 (N_15900,N_15126,N_15595);
nor U15901 (N_15901,N_14557,N_15591);
and U15902 (N_15902,N_14489,N_14503);
or U15903 (N_15903,N_15538,N_15436);
or U15904 (N_15904,N_14709,N_14976);
nor U15905 (N_15905,N_15472,N_15458);
xor U15906 (N_15906,N_14844,N_15462);
and U15907 (N_15907,N_14814,N_14501);
nor U15908 (N_15908,N_14469,N_14837);
and U15909 (N_15909,N_15188,N_14977);
nor U15910 (N_15910,N_14859,N_14545);
xor U15911 (N_15911,N_14714,N_14965);
nor U15912 (N_15912,N_14810,N_15222);
xnor U15913 (N_15913,N_14668,N_15017);
nand U15914 (N_15914,N_15245,N_14863);
xor U15915 (N_15915,N_14466,N_15186);
and U15916 (N_15916,N_14742,N_15121);
or U15917 (N_15917,N_15238,N_14494);
or U15918 (N_15918,N_15264,N_14945);
nand U15919 (N_15919,N_15345,N_15053);
nand U15920 (N_15920,N_14451,N_15411);
or U15921 (N_15921,N_14476,N_15457);
xor U15922 (N_15922,N_15081,N_14881);
nand U15923 (N_15923,N_14885,N_14829);
or U15924 (N_15924,N_15351,N_14467);
nand U15925 (N_15925,N_15305,N_14866);
nor U15926 (N_15926,N_14455,N_14765);
xnor U15927 (N_15927,N_14760,N_15481);
and U15928 (N_15928,N_14729,N_15266);
and U15929 (N_15929,N_15232,N_14664);
nand U15930 (N_15930,N_14923,N_14419);
and U15931 (N_15931,N_14571,N_15111);
nand U15932 (N_15932,N_15488,N_15032);
xnor U15933 (N_15933,N_15469,N_14749);
or U15934 (N_15934,N_15539,N_15545);
or U15935 (N_15935,N_15494,N_14628);
and U15936 (N_15936,N_15478,N_15528);
xnor U15937 (N_15937,N_14908,N_15262);
nand U15938 (N_15938,N_14781,N_15023);
and U15939 (N_15939,N_15270,N_14416);
nand U15940 (N_15940,N_14510,N_14995);
or U15941 (N_15941,N_14491,N_14784);
xor U15942 (N_15942,N_14449,N_14934);
or U15943 (N_15943,N_14524,N_14572);
and U15944 (N_15944,N_14728,N_14634);
or U15945 (N_15945,N_15434,N_14495);
and U15946 (N_15946,N_14716,N_14930);
xor U15947 (N_15947,N_14618,N_15423);
nand U15948 (N_15948,N_15201,N_15208);
or U15949 (N_15949,N_14516,N_14772);
nand U15950 (N_15950,N_15146,N_14897);
nor U15951 (N_15951,N_14770,N_15530);
nor U15952 (N_15952,N_14768,N_15139);
or U15953 (N_15953,N_15066,N_14498);
or U15954 (N_15954,N_15160,N_15060);
or U15955 (N_15955,N_15333,N_15095);
xnor U15956 (N_15956,N_14434,N_15079);
and U15957 (N_15957,N_14891,N_14796);
nor U15958 (N_15958,N_15281,N_15184);
nor U15959 (N_15959,N_15227,N_15487);
nor U15960 (N_15960,N_14695,N_14525);
or U15961 (N_15961,N_15486,N_15356);
nand U15962 (N_15962,N_15386,N_14591);
or U15963 (N_15963,N_15580,N_14998);
xnor U15964 (N_15964,N_14608,N_15412);
nor U15965 (N_15965,N_15009,N_14631);
nor U15966 (N_15966,N_15339,N_14717);
nand U15967 (N_15967,N_15298,N_14518);
and U15968 (N_15968,N_15249,N_14486);
and U15969 (N_15969,N_15558,N_15513);
or U15970 (N_15970,N_15168,N_14901);
and U15971 (N_15971,N_14758,N_15194);
and U15972 (N_15972,N_15502,N_15503);
xor U15973 (N_15973,N_14800,N_14595);
nand U15974 (N_15974,N_15128,N_14745);
or U15975 (N_15975,N_14838,N_15234);
xor U15976 (N_15976,N_15321,N_14678);
nor U15977 (N_15977,N_15153,N_15452);
nor U15978 (N_15978,N_14787,N_15372);
and U15979 (N_15979,N_14454,N_14513);
and U15980 (N_15980,N_14632,N_15230);
nor U15981 (N_15981,N_15213,N_15566);
nand U15982 (N_15982,N_15584,N_15433);
nand U15983 (N_15983,N_14921,N_15473);
nor U15984 (N_15984,N_15200,N_15446);
or U15985 (N_15985,N_15373,N_14659);
xnor U15986 (N_15986,N_14604,N_14974);
xor U15987 (N_15987,N_15145,N_15065);
and U15988 (N_15988,N_14596,N_15116);
nand U15989 (N_15989,N_15183,N_14585);
or U15990 (N_15990,N_14407,N_15203);
nor U15991 (N_15991,N_14879,N_15165);
or U15992 (N_15992,N_15579,N_14959);
nor U15993 (N_15993,N_15042,N_14450);
and U15994 (N_15994,N_15082,N_15352);
nor U15995 (N_15995,N_14425,N_15302);
nor U15996 (N_15996,N_14793,N_14962);
nor U15997 (N_15997,N_15306,N_14896);
and U15998 (N_15998,N_15113,N_15456);
nor U15999 (N_15999,N_15244,N_14830);
or U16000 (N_16000,N_14957,N_14967);
nor U16001 (N_16001,N_14932,N_15504);
nand U16002 (N_16002,N_14633,N_15105);
nand U16003 (N_16003,N_14414,N_14761);
nand U16004 (N_16004,N_14952,N_14935);
nand U16005 (N_16005,N_15181,N_15391);
and U16006 (N_16006,N_14440,N_15207);
and U16007 (N_16007,N_14902,N_14458);
xnor U16008 (N_16008,N_14637,N_15439);
xnor U16009 (N_16009,N_15030,N_15303);
nor U16010 (N_16010,N_15080,N_14640);
or U16011 (N_16011,N_14538,N_15035);
nor U16012 (N_16012,N_14743,N_15526);
nand U16013 (N_16013,N_14694,N_15124);
xnor U16014 (N_16014,N_14558,N_14862);
nor U16015 (N_16015,N_15290,N_14719);
and U16016 (N_16016,N_14958,N_14661);
nand U16017 (N_16017,N_15323,N_14956);
nor U16018 (N_16018,N_15492,N_15598);
and U16019 (N_16019,N_14675,N_14562);
nor U16020 (N_16020,N_14926,N_14941);
and U16021 (N_16021,N_15416,N_14718);
and U16022 (N_16022,N_15196,N_15424);
xor U16023 (N_16023,N_14918,N_14874);
nor U16024 (N_16024,N_14402,N_15525);
xnor U16025 (N_16025,N_14801,N_15175);
nand U16026 (N_16026,N_15061,N_14910);
xor U16027 (N_16027,N_15014,N_15179);
nor U16028 (N_16028,N_14517,N_15268);
nor U16029 (N_16029,N_15051,N_15554);
or U16030 (N_16030,N_15018,N_15418);
xor U16031 (N_16031,N_14825,N_15505);
xor U16032 (N_16032,N_15360,N_14815);
xor U16033 (N_16033,N_15483,N_15071);
xnor U16034 (N_16034,N_14614,N_15397);
nand U16035 (N_16035,N_14577,N_15073);
or U16036 (N_16036,N_15256,N_14889);
or U16037 (N_16037,N_15559,N_15410);
nand U16038 (N_16038,N_15046,N_15221);
nor U16039 (N_16039,N_15597,N_15248);
or U16040 (N_16040,N_14802,N_15536);
nand U16041 (N_16041,N_14400,N_15271);
xnor U16042 (N_16042,N_14980,N_15441);
nor U16043 (N_16043,N_15523,N_14437);
or U16044 (N_16044,N_15342,N_15593);
or U16045 (N_16045,N_15498,N_15259);
nor U16046 (N_16046,N_14412,N_14850);
and U16047 (N_16047,N_15163,N_15016);
xor U16048 (N_16048,N_14832,N_15358);
nand U16049 (N_16049,N_15137,N_14875);
and U16050 (N_16050,N_14727,N_14563);
xnor U16051 (N_16051,N_15019,N_14556);
or U16052 (N_16052,N_15384,N_14529);
and U16053 (N_16053,N_14507,N_14985);
nor U16054 (N_16054,N_14523,N_15402);
xor U16055 (N_16055,N_15177,N_15037);
and U16056 (N_16056,N_14453,N_15453);
xor U16057 (N_16057,N_15214,N_14560);
or U16058 (N_16058,N_15093,N_14994);
nor U16059 (N_16059,N_15583,N_14780);
or U16060 (N_16060,N_15318,N_15326);
or U16061 (N_16061,N_15131,N_15239);
nor U16062 (N_16062,N_14671,N_14569);
xor U16063 (N_16063,N_14933,N_15008);
and U16064 (N_16064,N_15575,N_15577);
nand U16065 (N_16065,N_14900,N_15354);
or U16066 (N_16066,N_14514,N_15540);
and U16067 (N_16067,N_14892,N_15561);
or U16068 (N_16068,N_15585,N_14792);
and U16069 (N_16069,N_14475,N_15190);
or U16070 (N_16070,N_15142,N_15491);
nor U16071 (N_16071,N_14574,N_14597);
nor U16072 (N_16072,N_15374,N_15506);
nand U16073 (N_16073,N_14578,N_15275);
xnor U16074 (N_16074,N_15002,N_15363);
and U16075 (N_16075,N_15378,N_14754);
or U16076 (N_16076,N_15496,N_15300);
nand U16077 (N_16077,N_14497,N_14641);
xnor U16078 (N_16078,N_14883,N_14598);
and U16079 (N_16079,N_14939,N_14551);
or U16080 (N_16080,N_15549,N_14488);
nor U16081 (N_16081,N_14706,N_15461);
and U16082 (N_16082,N_14920,N_15516);
xor U16083 (N_16083,N_15117,N_15546);
or U16084 (N_16084,N_14536,N_14522);
and U16085 (N_16085,N_15123,N_15518);
nor U16086 (N_16086,N_14601,N_15130);
xnor U16087 (N_16087,N_15236,N_15572);
nor U16088 (N_16088,N_14410,N_15090);
or U16089 (N_16089,N_14487,N_15127);
nor U16090 (N_16090,N_14636,N_14988);
xor U16091 (N_16091,N_15311,N_15000);
or U16092 (N_16092,N_14677,N_15209);
nand U16093 (N_16093,N_15044,N_14579);
xnor U16094 (N_16094,N_14406,N_14747);
xor U16095 (N_16095,N_15578,N_15562);
and U16096 (N_16096,N_15063,N_15337);
nor U16097 (N_16097,N_15075,N_14540);
xnor U16098 (N_16098,N_14789,N_15226);
nor U16099 (N_16099,N_14778,N_15520);
nor U16100 (N_16100,N_15588,N_14417);
nor U16101 (N_16101,N_15365,N_14871);
and U16102 (N_16102,N_15409,N_14899);
xnor U16103 (N_16103,N_15255,N_14785);
or U16104 (N_16104,N_14681,N_14975);
xnor U16105 (N_16105,N_15295,N_15007);
nand U16106 (N_16106,N_15195,N_15574);
nand U16107 (N_16107,N_15501,N_15263);
nor U16108 (N_16108,N_14584,N_15102);
nand U16109 (N_16109,N_14968,N_14472);
or U16110 (N_16110,N_14949,N_15316);
and U16111 (N_16111,N_15371,N_15156);
and U16112 (N_16112,N_15215,N_14741);
or U16113 (N_16113,N_15317,N_15564);
or U16114 (N_16114,N_15180,N_15257);
or U16115 (N_16115,N_15449,N_15445);
nor U16116 (N_16116,N_14776,N_15114);
or U16117 (N_16117,N_14953,N_14878);
xor U16118 (N_16118,N_14686,N_15571);
nand U16119 (N_16119,N_14428,N_15467);
xnor U16120 (N_16120,N_15176,N_14872);
or U16121 (N_16121,N_15551,N_14541);
nand U16122 (N_16122,N_15553,N_14626);
nor U16123 (N_16123,N_15284,N_14916);
xnor U16124 (N_16124,N_15240,N_15480);
and U16125 (N_16125,N_14520,N_14991);
xnor U16126 (N_16126,N_14963,N_14970);
nor U16127 (N_16127,N_14619,N_15085);
and U16128 (N_16128,N_15437,N_15038);
and U16129 (N_16129,N_14411,N_15563);
and U16130 (N_16130,N_15138,N_14676);
or U16131 (N_16131,N_15022,N_14978);
nor U16132 (N_16132,N_15385,N_14907);
nand U16133 (N_16133,N_14831,N_14759);
nor U16134 (N_16134,N_15210,N_14753);
nor U16135 (N_16135,N_14554,N_15447);
xnor U16136 (N_16136,N_15403,N_14421);
xnor U16137 (N_16137,N_14468,N_15353);
and U16138 (N_16138,N_14856,N_14587);
nor U16139 (N_16139,N_14790,N_14657);
or U16140 (N_16140,N_15045,N_14672);
or U16141 (N_16141,N_14459,N_14833);
xnor U16142 (N_16142,N_14913,N_14807);
nor U16143 (N_16143,N_14925,N_14982);
nor U16144 (N_16144,N_14723,N_14950);
xnor U16145 (N_16145,N_14660,N_14752);
xor U16146 (N_16146,N_14750,N_15466);
nand U16147 (N_16147,N_15087,N_14997);
or U16148 (N_16148,N_14880,N_14573);
nor U16149 (N_16149,N_15279,N_14774);
nand U16150 (N_16150,N_15511,N_15309);
xnor U16151 (N_16151,N_15400,N_14662);
nor U16152 (N_16152,N_15328,N_15122);
and U16153 (N_16153,N_14915,N_14736);
xnor U16154 (N_16154,N_15429,N_15484);
nand U16155 (N_16155,N_15185,N_15376);
and U16156 (N_16156,N_15294,N_14928);
or U16157 (N_16157,N_14461,N_15150);
xnor U16158 (N_16158,N_15254,N_14643);
xnor U16159 (N_16159,N_15474,N_15189);
and U16160 (N_16160,N_14549,N_14537);
nor U16161 (N_16161,N_14843,N_14732);
or U16162 (N_16162,N_15241,N_15515);
nor U16163 (N_16163,N_15283,N_15192);
nor U16164 (N_16164,N_15109,N_15151);
xor U16165 (N_16165,N_14964,N_14841);
or U16166 (N_16166,N_14834,N_15132);
nor U16167 (N_16167,N_14679,N_15033);
and U16168 (N_16168,N_14463,N_14550);
xnor U16169 (N_16169,N_14442,N_14931);
nand U16170 (N_16170,N_14937,N_14938);
xnor U16171 (N_16171,N_14655,N_14484);
and U16172 (N_16172,N_15355,N_14762);
xor U16173 (N_16173,N_15347,N_14570);
and U16174 (N_16174,N_15125,N_15159);
and U16175 (N_16175,N_14526,N_15136);
xnor U16176 (N_16176,N_14839,N_14658);
and U16177 (N_16177,N_14943,N_15454);
and U16178 (N_16178,N_15218,N_14528);
xor U16179 (N_16179,N_14989,N_14674);
nor U16180 (N_16180,N_14948,N_15261);
or U16181 (N_16181,N_15475,N_14705);
and U16182 (N_16182,N_14757,N_15120);
xor U16183 (N_16183,N_14594,N_15465);
or U16184 (N_16184,N_15250,N_14788);
nand U16185 (N_16185,N_15229,N_15219);
or U16186 (N_16186,N_14504,N_14812);
nand U16187 (N_16187,N_15346,N_14873);
nor U16188 (N_16188,N_14951,N_14546);
or U16189 (N_16189,N_14647,N_14433);
xnor U16190 (N_16190,N_15212,N_15509);
nor U16191 (N_16191,N_14447,N_15052);
nor U16192 (N_16192,N_15155,N_14670);
nand U16193 (N_16193,N_14955,N_14882);
and U16194 (N_16194,N_15173,N_15166);
nor U16195 (N_16195,N_14795,N_14996);
nand U16196 (N_16196,N_15364,N_14919);
or U16197 (N_16197,N_14649,N_15359);
nand U16198 (N_16198,N_15383,N_14725);
or U16199 (N_16199,N_15164,N_14477);
nor U16200 (N_16200,N_14890,N_14476);
or U16201 (N_16201,N_14810,N_15136);
or U16202 (N_16202,N_14732,N_14556);
and U16203 (N_16203,N_14672,N_14460);
nor U16204 (N_16204,N_15447,N_14823);
nor U16205 (N_16205,N_14681,N_15391);
nand U16206 (N_16206,N_14401,N_14534);
nor U16207 (N_16207,N_15285,N_14453);
and U16208 (N_16208,N_15595,N_14644);
nor U16209 (N_16209,N_15450,N_15460);
or U16210 (N_16210,N_14809,N_14877);
and U16211 (N_16211,N_15066,N_14506);
xor U16212 (N_16212,N_15166,N_14636);
and U16213 (N_16213,N_15166,N_14524);
and U16214 (N_16214,N_14417,N_15123);
or U16215 (N_16215,N_14567,N_15012);
and U16216 (N_16216,N_15211,N_15275);
nor U16217 (N_16217,N_15154,N_14545);
and U16218 (N_16218,N_14423,N_15093);
xnor U16219 (N_16219,N_14412,N_14804);
or U16220 (N_16220,N_15592,N_15217);
or U16221 (N_16221,N_14638,N_14893);
or U16222 (N_16222,N_14647,N_15527);
nor U16223 (N_16223,N_14783,N_15231);
or U16224 (N_16224,N_15530,N_15235);
and U16225 (N_16225,N_15038,N_14719);
xor U16226 (N_16226,N_14613,N_14659);
and U16227 (N_16227,N_15078,N_14807);
or U16228 (N_16228,N_14680,N_14538);
nand U16229 (N_16229,N_14867,N_14793);
or U16230 (N_16230,N_15012,N_15207);
nand U16231 (N_16231,N_14558,N_15114);
nand U16232 (N_16232,N_15042,N_15008);
nand U16233 (N_16233,N_14834,N_14864);
and U16234 (N_16234,N_14534,N_14484);
nand U16235 (N_16235,N_15052,N_15319);
xor U16236 (N_16236,N_14548,N_15038);
or U16237 (N_16237,N_14676,N_14800);
or U16238 (N_16238,N_14558,N_15174);
nand U16239 (N_16239,N_14826,N_14473);
xor U16240 (N_16240,N_14780,N_14976);
nor U16241 (N_16241,N_14866,N_14481);
nor U16242 (N_16242,N_14799,N_15342);
nand U16243 (N_16243,N_15257,N_15299);
nand U16244 (N_16244,N_14829,N_15087);
nor U16245 (N_16245,N_15268,N_15150);
nor U16246 (N_16246,N_14430,N_14670);
nand U16247 (N_16247,N_15283,N_14891);
xnor U16248 (N_16248,N_15438,N_15496);
nor U16249 (N_16249,N_15310,N_14422);
nand U16250 (N_16250,N_15336,N_14968);
and U16251 (N_16251,N_14837,N_14513);
and U16252 (N_16252,N_15296,N_14843);
xor U16253 (N_16253,N_14826,N_15461);
xnor U16254 (N_16254,N_14973,N_15537);
nor U16255 (N_16255,N_15487,N_15486);
nand U16256 (N_16256,N_15338,N_14488);
or U16257 (N_16257,N_15244,N_15302);
nand U16258 (N_16258,N_14839,N_15315);
nand U16259 (N_16259,N_14430,N_14489);
nand U16260 (N_16260,N_15357,N_14482);
nor U16261 (N_16261,N_15044,N_14989);
nand U16262 (N_16262,N_15356,N_15364);
or U16263 (N_16263,N_15489,N_14775);
or U16264 (N_16264,N_14619,N_15519);
and U16265 (N_16265,N_14536,N_15087);
and U16266 (N_16266,N_14443,N_14918);
nor U16267 (N_16267,N_15507,N_14546);
xnor U16268 (N_16268,N_14692,N_15351);
nand U16269 (N_16269,N_15468,N_14635);
and U16270 (N_16270,N_14767,N_14631);
or U16271 (N_16271,N_15272,N_15247);
nand U16272 (N_16272,N_14704,N_15455);
nor U16273 (N_16273,N_14634,N_15306);
nand U16274 (N_16274,N_14712,N_15066);
or U16275 (N_16275,N_14937,N_15244);
xnor U16276 (N_16276,N_15045,N_15554);
and U16277 (N_16277,N_14931,N_15451);
xor U16278 (N_16278,N_14987,N_14696);
nor U16279 (N_16279,N_15567,N_14667);
nand U16280 (N_16280,N_14595,N_14514);
xor U16281 (N_16281,N_15096,N_14579);
and U16282 (N_16282,N_14795,N_14624);
nor U16283 (N_16283,N_14572,N_14531);
and U16284 (N_16284,N_15495,N_15133);
and U16285 (N_16285,N_14420,N_14459);
and U16286 (N_16286,N_15530,N_15046);
nand U16287 (N_16287,N_14656,N_14446);
nor U16288 (N_16288,N_14974,N_15409);
nand U16289 (N_16289,N_14748,N_14466);
or U16290 (N_16290,N_15572,N_15339);
nand U16291 (N_16291,N_15120,N_14546);
nor U16292 (N_16292,N_15280,N_14715);
nor U16293 (N_16293,N_15159,N_14584);
and U16294 (N_16294,N_15555,N_14453);
or U16295 (N_16295,N_14818,N_14865);
nor U16296 (N_16296,N_14571,N_15086);
nand U16297 (N_16297,N_15334,N_14953);
or U16298 (N_16298,N_14510,N_15363);
and U16299 (N_16299,N_15332,N_14869);
and U16300 (N_16300,N_15279,N_15295);
and U16301 (N_16301,N_14745,N_15317);
xor U16302 (N_16302,N_15587,N_15035);
or U16303 (N_16303,N_15449,N_14403);
xor U16304 (N_16304,N_14848,N_15008);
and U16305 (N_16305,N_15304,N_14404);
nor U16306 (N_16306,N_15482,N_15558);
xnor U16307 (N_16307,N_15155,N_14621);
or U16308 (N_16308,N_14626,N_14948);
or U16309 (N_16309,N_15280,N_14711);
xor U16310 (N_16310,N_15129,N_15590);
nand U16311 (N_16311,N_14933,N_14632);
or U16312 (N_16312,N_14860,N_15075);
nor U16313 (N_16313,N_15121,N_14444);
and U16314 (N_16314,N_15201,N_15558);
nor U16315 (N_16315,N_15233,N_14854);
nor U16316 (N_16316,N_14797,N_15419);
nor U16317 (N_16317,N_15260,N_14919);
xnor U16318 (N_16318,N_15311,N_15336);
xor U16319 (N_16319,N_14510,N_14696);
or U16320 (N_16320,N_14810,N_15545);
or U16321 (N_16321,N_14965,N_14809);
or U16322 (N_16322,N_14683,N_15363);
nor U16323 (N_16323,N_15414,N_14524);
nor U16324 (N_16324,N_15425,N_14507);
xor U16325 (N_16325,N_15160,N_14516);
nor U16326 (N_16326,N_14909,N_15152);
xor U16327 (N_16327,N_15412,N_14702);
or U16328 (N_16328,N_14451,N_14817);
xnor U16329 (N_16329,N_14758,N_14918);
xnor U16330 (N_16330,N_15280,N_14619);
and U16331 (N_16331,N_15155,N_14931);
nor U16332 (N_16332,N_14584,N_14751);
and U16333 (N_16333,N_14936,N_15059);
nor U16334 (N_16334,N_15560,N_15454);
xor U16335 (N_16335,N_15351,N_15342);
nand U16336 (N_16336,N_15428,N_14526);
nand U16337 (N_16337,N_14529,N_14767);
nand U16338 (N_16338,N_14471,N_15422);
nand U16339 (N_16339,N_14696,N_14663);
nor U16340 (N_16340,N_14759,N_14774);
nand U16341 (N_16341,N_15463,N_15272);
xor U16342 (N_16342,N_14527,N_14665);
xnor U16343 (N_16343,N_14775,N_14607);
nor U16344 (N_16344,N_14877,N_14550);
nand U16345 (N_16345,N_15594,N_15308);
xnor U16346 (N_16346,N_15412,N_15546);
or U16347 (N_16347,N_14906,N_14708);
or U16348 (N_16348,N_15128,N_14955);
nand U16349 (N_16349,N_15307,N_14648);
or U16350 (N_16350,N_14924,N_14903);
xnor U16351 (N_16351,N_14560,N_15159);
or U16352 (N_16352,N_14761,N_14912);
or U16353 (N_16353,N_15031,N_15544);
xor U16354 (N_16354,N_14880,N_15261);
or U16355 (N_16355,N_15187,N_15040);
xnor U16356 (N_16356,N_15117,N_14912);
or U16357 (N_16357,N_15427,N_15244);
nand U16358 (N_16358,N_15341,N_14459);
and U16359 (N_16359,N_14946,N_15533);
nand U16360 (N_16360,N_15065,N_15204);
xnor U16361 (N_16361,N_14946,N_15296);
and U16362 (N_16362,N_15050,N_15568);
nand U16363 (N_16363,N_15413,N_15377);
xor U16364 (N_16364,N_15277,N_15279);
nand U16365 (N_16365,N_14604,N_15571);
and U16366 (N_16366,N_15091,N_15027);
xor U16367 (N_16367,N_14737,N_15106);
nand U16368 (N_16368,N_14480,N_14519);
and U16369 (N_16369,N_14706,N_14413);
xnor U16370 (N_16370,N_14753,N_15318);
and U16371 (N_16371,N_14934,N_15436);
and U16372 (N_16372,N_14727,N_15347);
xnor U16373 (N_16373,N_14766,N_15312);
nor U16374 (N_16374,N_14887,N_15109);
or U16375 (N_16375,N_14760,N_15571);
xnor U16376 (N_16376,N_14605,N_14994);
and U16377 (N_16377,N_15039,N_14659);
nor U16378 (N_16378,N_15442,N_15237);
or U16379 (N_16379,N_14529,N_15400);
xor U16380 (N_16380,N_15485,N_14755);
and U16381 (N_16381,N_14586,N_15279);
and U16382 (N_16382,N_15309,N_14444);
and U16383 (N_16383,N_15170,N_15465);
xnor U16384 (N_16384,N_14676,N_15029);
or U16385 (N_16385,N_14648,N_14424);
nand U16386 (N_16386,N_15306,N_14916);
and U16387 (N_16387,N_14605,N_14747);
and U16388 (N_16388,N_14682,N_14618);
or U16389 (N_16389,N_15109,N_15411);
and U16390 (N_16390,N_15467,N_14906);
xnor U16391 (N_16391,N_15381,N_15148);
nor U16392 (N_16392,N_14865,N_15338);
nor U16393 (N_16393,N_14957,N_15187);
xnor U16394 (N_16394,N_14723,N_14932);
or U16395 (N_16395,N_14501,N_15284);
nand U16396 (N_16396,N_15214,N_14688);
xor U16397 (N_16397,N_15423,N_14717);
xor U16398 (N_16398,N_14902,N_15404);
nor U16399 (N_16399,N_14539,N_15330);
or U16400 (N_16400,N_14468,N_14780);
xnor U16401 (N_16401,N_14963,N_15098);
nor U16402 (N_16402,N_15392,N_14438);
or U16403 (N_16403,N_14922,N_14925);
or U16404 (N_16404,N_14990,N_14837);
xnor U16405 (N_16405,N_14804,N_14561);
and U16406 (N_16406,N_14717,N_15193);
or U16407 (N_16407,N_15113,N_14746);
or U16408 (N_16408,N_15514,N_14492);
xor U16409 (N_16409,N_15047,N_15051);
nor U16410 (N_16410,N_15417,N_14981);
xnor U16411 (N_16411,N_15009,N_15292);
or U16412 (N_16412,N_14916,N_14686);
nor U16413 (N_16413,N_14883,N_15244);
nand U16414 (N_16414,N_14444,N_15299);
nor U16415 (N_16415,N_15124,N_14969);
or U16416 (N_16416,N_15282,N_14956);
nand U16417 (N_16417,N_15446,N_14989);
nor U16418 (N_16418,N_14665,N_14646);
nand U16419 (N_16419,N_14473,N_14601);
xor U16420 (N_16420,N_14632,N_14509);
nand U16421 (N_16421,N_15416,N_15238);
nand U16422 (N_16422,N_15527,N_15504);
nor U16423 (N_16423,N_14708,N_15533);
xnor U16424 (N_16424,N_14908,N_15361);
nand U16425 (N_16425,N_14435,N_15462);
and U16426 (N_16426,N_14587,N_14883);
or U16427 (N_16427,N_14570,N_14705);
nor U16428 (N_16428,N_14468,N_15437);
or U16429 (N_16429,N_14795,N_15579);
or U16430 (N_16430,N_15517,N_14759);
or U16431 (N_16431,N_14810,N_15396);
and U16432 (N_16432,N_15252,N_14542);
xnor U16433 (N_16433,N_14559,N_15302);
nand U16434 (N_16434,N_14412,N_14456);
or U16435 (N_16435,N_14967,N_15427);
nand U16436 (N_16436,N_14808,N_15001);
and U16437 (N_16437,N_14836,N_14817);
xnor U16438 (N_16438,N_15003,N_15462);
xnor U16439 (N_16439,N_15573,N_14526);
xnor U16440 (N_16440,N_15116,N_15206);
or U16441 (N_16441,N_15050,N_15586);
or U16442 (N_16442,N_14540,N_14530);
or U16443 (N_16443,N_14691,N_15280);
nor U16444 (N_16444,N_15179,N_15073);
nor U16445 (N_16445,N_15171,N_14499);
nand U16446 (N_16446,N_15484,N_15027);
and U16447 (N_16447,N_15327,N_15467);
nor U16448 (N_16448,N_14684,N_14756);
or U16449 (N_16449,N_15095,N_14673);
nand U16450 (N_16450,N_15372,N_15435);
nand U16451 (N_16451,N_15018,N_15295);
nand U16452 (N_16452,N_15157,N_14459);
xnor U16453 (N_16453,N_15179,N_14622);
nor U16454 (N_16454,N_15260,N_15172);
nand U16455 (N_16455,N_15544,N_14773);
xnor U16456 (N_16456,N_15236,N_14577);
nor U16457 (N_16457,N_15531,N_15505);
xor U16458 (N_16458,N_14611,N_15287);
xor U16459 (N_16459,N_14792,N_15493);
and U16460 (N_16460,N_14833,N_15329);
or U16461 (N_16461,N_14709,N_14563);
nor U16462 (N_16462,N_14962,N_14942);
nand U16463 (N_16463,N_14673,N_15544);
and U16464 (N_16464,N_14425,N_15480);
or U16465 (N_16465,N_14515,N_14595);
or U16466 (N_16466,N_15181,N_15422);
xnor U16467 (N_16467,N_14908,N_14559);
nand U16468 (N_16468,N_14618,N_14565);
nor U16469 (N_16469,N_14475,N_15304);
and U16470 (N_16470,N_14505,N_15064);
xnor U16471 (N_16471,N_15121,N_14473);
or U16472 (N_16472,N_15559,N_15578);
and U16473 (N_16473,N_15204,N_14943);
xnor U16474 (N_16474,N_14616,N_15202);
nor U16475 (N_16475,N_15132,N_14540);
xnor U16476 (N_16476,N_14659,N_15388);
nand U16477 (N_16477,N_15049,N_14466);
nor U16478 (N_16478,N_14880,N_15155);
nand U16479 (N_16479,N_15014,N_14628);
or U16480 (N_16480,N_15208,N_15258);
or U16481 (N_16481,N_15407,N_15231);
xor U16482 (N_16482,N_15301,N_14767);
xnor U16483 (N_16483,N_14928,N_15511);
and U16484 (N_16484,N_14533,N_15259);
or U16485 (N_16485,N_15111,N_14836);
and U16486 (N_16486,N_14836,N_15543);
and U16487 (N_16487,N_14531,N_15022);
xnor U16488 (N_16488,N_14674,N_15062);
or U16489 (N_16489,N_14696,N_15096);
and U16490 (N_16490,N_15451,N_14802);
or U16491 (N_16491,N_14631,N_15095);
or U16492 (N_16492,N_15278,N_15355);
or U16493 (N_16493,N_14830,N_15328);
and U16494 (N_16494,N_15265,N_14632);
and U16495 (N_16495,N_14844,N_14964);
nand U16496 (N_16496,N_15423,N_14829);
nor U16497 (N_16497,N_14587,N_14745);
xor U16498 (N_16498,N_14729,N_15530);
nor U16499 (N_16499,N_14426,N_15317);
nand U16500 (N_16500,N_14434,N_14591);
xnor U16501 (N_16501,N_15277,N_14873);
or U16502 (N_16502,N_15189,N_15393);
and U16503 (N_16503,N_15537,N_14950);
or U16504 (N_16504,N_14469,N_14682);
xor U16505 (N_16505,N_15119,N_14920);
nand U16506 (N_16506,N_15563,N_15072);
nor U16507 (N_16507,N_15181,N_14973);
nor U16508 (N_16508,N_14993,N_14471);
or U16509 (N_16509,N_14767,N_14541);
nor U16510 (N_16510,N_14671,N_14755);
nor U16511 (N_16511,N_15521,N_15250);
and U16512 (N_16512,N_14947,N_15183);
xor U16513 (N_16513,N_15541,N_14918);
nand U16514 (N_16514,N_15394,N_14902);
nor U16515 (N_16515,N_15516,N_14728);
xor U16516 (N_16516,N_15025,N_15437);
xnor U16517 (N_16517,N_15165,N_14501);
xor U16518 (N_16518,N_14971,N_15047);
and U16519 (N_16519,N_14693,N_14619);
nor U16520 (N_16520,N_14549,N_14541);
nand U16521 (N_16521,N_14511,N_14745);
nor U16522 (N_16522,N_15268,N_14452);
or U16523 (N_16523,N_14996,N_15543);
xor U16524 (N_16524,N_15167,N_14681);
nand U16525 (N_16525,N_14702,N_15030);
and U16526 (N_16526,N_15076,N_15314);
or U16527 (N_16527,N_14681,N_15471);
xor U16528 (N_16528,N_15354,N_15356);
and U16529 (N_16529,N_15327,N_15284);
and U16530 (N_16530,N_15043,N_14998);
nand U16531 (N_16531,N_14430,N_15472);
xnor U16532 (N_16532,N_15226,N_15053);
and U16533 (N_16533,N_14969,N_14419);
nand U16534 (N_16534,N_15529,N_14975);
and U16535 (N_16535,N_15373,N_14750);
nand U16536 (N_16536,N_14848,N_14462);
nand U16537 (N_16537,N_14679,N_15220);
or U16538 (N_16538,N_14825,N_15447);
xor U16539 (N_16539,N_15323,N_15411);
or U16540 (N_16540,N_14705,N_14942);
nor U16541 (N_16541,N_15401,N_15306);
or U16542 (N_16542,N_15557,N_15189);
or U16543 (N_16543,N_15236,N_15301);
and U16544 (N_16544,N_14564,N_14724);
or U16545 (N_16545,N_15296,N_15548);
and U16546 (N_16546,N_14435,N_15375);
and U16547 (N_16547,N_15140,N_14707);
nand U16548 (N_16548,N_14484,N_14838);
nor U16549 (N_16549,N_15567,N_14822);
nand U16550 (N_16550,N_15328,N_14999);
nand U16551 (N_16551,N_15134,N_14461);
nor U16552 (N_16552,N_14507,N_14972);
and U16553 (N_16553,N_14518,N_14811);
or U16554 (N_16554,N_14490,N_14574);
or U16555 (N_16555,N_14618,N_14459);
and U16556 (N_16556,N_15304,N_15542);
or U16557 (N_16557,N_14998,N_15268);
nand U16558 (N_16558,N_15320,N_14678);
nand U16559 (N_16559,N_14493,N_15516);
and U16560 (N_16560,N_15290,N_15433);
or U16561 (N_16561,N_14468,N_15540);
nor U16562 (N_16562,N_14418,N_15227);
nor U16563 (N_16563,N_15076,N_14479);
nor U16564 (N_16564,N_14897,N_14846);
nand U16565 (N_16565,N_14758,N_14459);
and U16566 (N_16566,N_14514,N_14539);
nand U16567 (N_16567,N_15369,N_14621);
and U16568 (N_16568,N_15232,N_15144);
nor U16569 (N_16569,N_14446,N_14442);
or U16570 (N_16570,N_14886,N_15447);
nor U16571 (N_16571,N_15185,N_14947);
xnor U16572 (N_16572,N_15042,N_14451);
xor U16573 (N_16573,N_14990,N_15108);
nor U16574 (N_16574,N_15368,N_14604);
or U16575 (N_16575,N_15536,N_15197);
or U16576 (N_16576,N_15044,N_15157);
and U16577 (N_16577,N_15092,N_14741);
and U16578 (N_16578,N_15202,N_15035);
and U16579 (N_16579,N_14573,N_15406);
nand U16580 (N_16580,N_14556,N_14847);
nor U16581 (N_16581,N_15048,N_15391);
nor U16582 (N_16582,N_14928,N_14685);
or U16583 (N_16583,N_15289,N_15495);
nor U16584 (N_16584,N_15111,N_15528);
nor U16585 (N_16585,N_15351,N_14918);
nand U16586 (N_16586,N_15318,N_14546);
or U16587 (N_16587,N_14748,N_14850);
or U16588 (N_16588,N_14695,N_14547);
or U16589 (N_16589,N_14528,N_14816);
nand U16590 (N_16590,N_14822,N_14827);
xor U16591 (N_16591,N_15352,N_14777);
and U16592 (N_16592,N_14518,N_14656);
xnor U16593 (N_16593,N_14538,N_14699);
nor U16594 (N_16594,N_15268,N_15496);
nor U16595 (N_16595,N_14799,N_14419);
nand U16596 (N_16596,N_15243,N_15558);
and U16597 (N_16597,N_14949,N_14437);
or U16598 (N_16598,N_15410,N_14782);
nand U16599 (N_16599,N_15257,N_14493);
xnor U16600 (N_16600,N_14701,N_14870);
and U16601 (N_16601,N_14952,N_15407);
nand U16602 (N_16602,N_15105,N_15011);
xor U16603 (N_16603,N_14872,N_15562);
or U16604 (N_16604,N_15024,N_15508);
or U16605 (N_16605,N_15011,N_15538);
or U16606 (N_16606,N_14742,N_15004);
and U16607 (N_16607,N_15119,N_15504);
nand U16608 (N_16608,N_15317,N_15350);
xor U16609 (N_16609,N_14863,N_14509);
or U16610 (N_16610,N_14644,N_14936);
and U16611 (N_16611,N_14605,N_14522);
or U16612 (N_16612,N_15330,N_14469);
or U16613 (N_16613,N_14575,N_15264);
xnor U16614 (N_16614,N_14507,N_15146);
xor U16615 (N_16615,N_15145,N_14817);
and U16616 (N_16616,N_14619,N_14575);
nor U16617 (N_16617,N_15190,N_14490);
nor U16618 (N_16618,N_15354,N_15363);
nor U16619 (N_16619,N_14923,N_14583);
and U16620 (N_16620,N_14545,N_14795);
nand U16621 (N_16621,N_15038,N_14871);
xor U16622 (N_16622,N_14726,N_15591);
xnor U16623 (N_16623,N_15084,N_15521);
xor U16624 (N_16624,N_14472,N_15450);
xor U16625 (N_16625,N_14866,N_15532);
nand U16626 (N_16626,N_15361,N_15062);
nor U16627 (N_16627,N_14991,N_14837);
xnor U16628 (N_16628,N_15390,N_15510);
xnor U16629 (N_16629,N_14414,N_14980);
nand U16630 (N_16630,N_14881,N_15218);
nand U16631 (N_16631,N_14917,N_15117);
nand U16632 (N_16632,N_15326,N_14576);
and U16633 (N_16633,N_14423,N_14738);
xor U16634 (N_16634,N_15120,N_14732);
xor U16635 (N_16635,N_15009,N_15527);
or U16636 (N_16636,N_14806,N_14474);
nand U16637 (N_16637,N_14639,N_14515);
and U16638 (N_16638,N_15148,N_15326);
nor U16639 (N_16639,N_14994,N_15009);
and U16640 (N_16640,N_15311,N_15257);
nor U16641 (N_16641,N_14851,N_14594);
nor U16642 (N_16642,N_15129,N_14707);
and U16643 (N_16643,N_14766,N_14570);
xor U16644 (N_16644,N_14742,N_15390);
nor U16645 (N_16645,N_15168,N_14447);
nor U16646 (N_16646,N_15003,N_14769);
and U16647 (N_16647,N_14624,N_14709);
and U16648 (N_16648,N_15523,N_14503);
and U16649 (N_16649,N_15348,N_14496);
nand U16650 (N_16650,N_14921,N_15340);
or U16651 (N_16651,N_15419,N_14714);
or U16652 (N_16652,N_14617,N_15109);
xor U16653 (N_16653,N_15435,N_14468);
nand U16654 (N_16654,N_14896,N_14406);
or U16655 (N_16655,N_14466,N_14452);
or U16656 (N_16656,N_15162,N_14845);
and U16657 (N_16657,N_14994,N_15333);
and U16658 (N_16658,N_14689,N_15599);
xor U16659 (N_16659,N_15322,N_15036);
xor U16660 (N_16660,N_14945,N_14479);
nor U16661 (N_16661,N_14463,N_15583);
nand U16662 (N_16662,N_14851,N_15114);
and U16663 (N_16663,N_15009,N_15080);
and U16664 (N_16664,N_15150,N_15247);
and U16665 (N_16665,N_14915,N_15232);
xnor U16666 (N_16666,N_14735,N_14862);
nand U16667 (N_16667,N_15064,N_14478);
xnor U16668 (N_16668,N_15258,N_15030);
xor U16669 (N_16669,N_15446,N_15455);
nor U16670 (N_16670,N_15292,N_14845);
xor U16671 (N_16671,N_15315,N_15346);
and U16672 (N_16672,N_14680,N_15309);
nand U16673 (N_16673,N_14611,N_14891);
nor U16674 (N_16674,N_14551,N_15110);
and U16675 (N_16675,N_14568,N_15507);
nor U16676 (N_16676,N_15273,N_15066);
nand U16677 (N_16677,N_15220,N_14953);
nor U16678 (N_16678,N_15153,N_15161);
nand U16679 (N_16679,N_14853,N_14429);
nor U16680 (N_16680,N_14932,N_14588);
nand U16681 (N_16681,N_14499,N_14400);
and U16682 (N_16682,N_14654,N_14518);
or U16683 (N_16683,N_15082,N_15170);
xor U16684 (N_16684,N_14589,N_15099);
nand U16685 (N_16685,N_14462,N_14449);
and U16686 (N_16686,N_15488,N_15260);
nand U16687 (N_16687,N_15571,N_15585);
and U16688 (N_16688,N_14698,N_15558);
or U16689 (N_16689,N_14888,N_14722);
xnor U16690 (N_16690,N_14855,N_14630);
or U16691 (N_16691,N_15419,N_14840);
nor U16692 (N_16692,N_14799,N_15067);
nand U16693 (N_16693,N_14944,N_14877);
nand U16694 (N_16694,N_15536,N_14467);
or U16695 (N_16695,N_14966,N_15088);
and U16696 (N_16696,N_15511,N_15590);
xnor U16697 (N_16697,N_14848,N_15014);
nor U16698 (N_16698,N_14612,N_14699);
or U16699 (N_16699,N_14900,N_15504);
nor U16700 (N_16700,N_15078,N_15461);
xnor U16701 (N_16701,N_14770,N_14835);
or U16702 (N_16702,N_15155,N_15058);
nor U16703 (N_16703,N_14647,N_15400);
xor U16704 (N_16704,N_14446,N_15127);
nor U16705 (N_16705,N_14603,N_14554);
xnor U16706 (N_16706,N_14755,N_15170);
nor U16707 (N_16707,N_15087,N_15111);
nor U16708 (N_16708,N_15307,N_15215);
nand U16709 (N_16709,N_14516,N_14905);
or U16710 (N_16710,N_15535,N_14702);
or U16711 (N_16711,N_15425,N_15327);
nor U16712 (N_16712,N_15370,N_14554);
nand U16713 (N_16713,N_15586,N_15026);
nor U16714 (N_16714,N_14590,N_14488);
xnor U16715 (N_16715,N_15184,N_15158);
nand U16716 (N_16716,N_15403,N_15322);
and U16717 (N_16717,N_14458,N_15152);
or U16718 (N_16718,N_15078,N_14770);
nand U16719 (N_16719,N_15252,N_15100);
nor U16720 (N_16720,N_14755,N_15578);
xor U16721 (N_16721,N_15566,N_15378);
and U16722 (N_16722,N_15548,N_15181);
or U16723 (N_16723,N_15088,N_15025);
or U16724 (N_16724,N_15570,N_14487);
and U16725 (N_16725,N_15194,N_14704);
xor U16726 (N_16726,N_15319,N_14442);
or U16727 (N_16727,N_15329,N_15121);
and U16728 (N_16728,N_14695,N_14512);
or U16729 (N_16729,N_15399,N_15432);
and U16730 (N_16730,N_14808,N_14630);
and U16731 (N_16731,N_14918,N_14536);
nand U16732 (N_16732,N_15251,N_15182);
xnor U16733 (N_16733,N_15481,N_15528);
xnor U16734 (N_16734,N_14687,N_14683);
and U16735 (N_16735,N_14965,N_15124);
nor U16736 (N_16736,N_15560,N_14408);
nand U16737 (N_16737,N_14945,N_15563);
or U16738 (N_16738,N_15091,N_15051);
nand U16739 (N_16739,N_15053,N_14520);
nand U16740 (N_16740,N_14966,N_14735);
xnor U16741 (N_16741,N_15564,N_14882);
or U16742 (N_16742,N_15356,N_14417);
xor U16743 (N_16743,N_14866,N_14520);
nor U16744 (N_16744,N_15045,N_14905);
and U16745 (N_16745,N_15256,N_15396);
and U16746 (N_16746,N_14814,N_14634);
nand U16747 (N_16747,N_15413,N_15339);
nand U16748 (N_16748,N_14878,N_15112);
xnor U16749 (N_16749,N_15517,N_15179);
nor U16750 (N_16750,N_15490,N_15011);
xnor U16751 (N_16751,N_14779,N_15499);
xnor U16752 (N_16752,N_14756,N_15072);
nor U16753 (N_16753,N_15501,N_15050);
nor U16754 (N_16754,N_15514,N_15556);
nand U16755 (N_16755,N_14584,N_14844);
or U16756 (N_16756,N_15291,N_14761);
and U16757 (N_16757,N_14483,N_15518);
or U16758 (N_16758,N_14554,N_15008);
or U16759 (N_16759,N_15425,N_14553);
nor U16760 (N_16760,N_14736,N_14588);
nand U16761 (N_16761,N_15451,N_14433);
nor U16762 (N_16762,N_14640,N_15557);
and U16763 (N_16763,N_15552,N_15497);
nand U16764 (N_16764,N_15530,N_15531);
nor U16765 (N_16765,N_14693,N_15280);
nor U16766 (N_16766,N_14450,N_15001);
nand U16767 (N_16767,N_15562,N_14645);
xnor U16768 (N_16768,N_14640,N_14549);
xor U16769 (N_16769,N_15479,N_15355);
nor U16770 (N_16770,N_14476,N_14688);
xor U16771 (N_16771,N_15068,N_15531);
nor U16772 (N_16772,N_14815,N_14693);
nor U16773 (N_16773,N_14452,N_14922);
nor U16774 (N_16774,N_14487,N_14418);
nand U16775 (N_16775,N_14592,N_15526);
xnor U16776 (N_16776,N_15380,N_14880);
nand U16777 (N_16777,N_15477,N_14463);
xnor U16778 (N_16778,N_14618,N_15304);
and U16779 (N_16779,N_15546,N_14683);
nand U16780 (N_16780,N_15076,N_15147);
and U16781 (N_16781,N_14495,N_15275);
nand U16782 (N_16782,N_15187,N_14438);
or U16783 (N_16783,N_14732,N_14532);
nor U16784 (N_16784,N_15459,N_15223);
and U16785 (N_16785,N_14511,N_14577);
or U16786 (N_16786,N_14909,N_14967);
nand U16787 (N_16787,N_15154,N_15040);
nand U16788 (N_16788,N_15534,N_15473);
nand U16789 (N_16789,N_15454,N_15095);
nor U16790 (N_16790,N_14923,N_14983);
nand U16791 (N_16791,N_15308,N_15239);
or U16792 (N_16792,N_15056,N_15563);
nand U16793 (N_16793,N_14802,N_14538);
nand U16794 (N_16794,N_14757,N_15296);
xor U16795 (N_16795,N_15265,N_14793);
xnor U16796 (N_16796,N_14567,N_15152);
nor U16797 (N_16797,N_14550,N_15339);
nand U16798 (N_16798,N_14631,N_14552);
nor U16799 (N_16799,N_14956,N_15283);
or U16800 (N_16800,N_16243,N_16615);
nor U16801 (N_16801,N_15837,N_15891);
or U16802 (N_16802,N_15870,N_16616);
xnor U16803 (N_16803,N_16575,N_15928);
nand U16804 (N_16804,N_16671,N_15844);
nand U16805 (N_16805,N_16069,N_15936);
or U16806 (N_16806,N_16656,N_16597);
or U16807 (N_16807,N_16689,N_16638);
and U16808 (N_16808,N_15974,N_16274);
xor U16809 (N_16809,N_15739,N_16114);
nand U16810 (N_16810,N_16008,N_15795);
xnor U16811 (N_16811,N_16448,N_16709);
nor U16812 (N_16812,N_16633,N_16596);
or U16813 (N_16813,N_16494,N_15742);
or U16814 (N_16814,N_16515,N_15694);
nand U16815 (N_16815,N_16681,N_15665);
and U16816 (N_16816,N_16737,N_15965);
nor U16817 (N_16817,N_15863,N_15849);
xnor U16818 (N_16818,N_15894,N_16761);
nand U16819 (N_16819,N_16343,N_16792);
nor U16820 (N_16820,N_16099,N_16520);
xnor U16821 (N_16821,N_15733,N_16079);
or U16822 (N_16822,N_16407,N_16493);
nand U16823 (N_16823,N_16036,N_16693);
or U16824 (N_16824,N_16351,N_15935);
nor U16825 (N_16825,N_15772,N_16798);
nor U16826 (N_16826,N_16478,N_16499);
nand U16827 (N_16827,N_16553,N_16053);
and U16828 (N_16828,N_15982,N_16423);
nor U16829 (N_16829,N_16608,N_16454);
or U16830 (N_16830,N_16348,N_16316);
nand U16831 (N_16831,N_15846,N_15930);
or U16832 (N_16832,N_16362,N_15612);
and U16833 (N_16833,N_16531,N_16613);
and U16834 (N_16834,N_16367,N_16406);
nor U16835 (N_16835,N_16731,N_15831);
xnor U16836 (N_16836,N_16146,N_16264);
nand U16837 (N_16837,N_15686,N_16547);
nor U16838 (N_16838,N_16320,N_16503);
or U16839 (N_16839,N_15964,N_16746);
nand U16840 (N_16840,N_16758,N_16391);
nand U16841 (N_16841,N_16446,N_16463);
or U16842 (N_16842,N_16513,N_15720);
nand U16843 (N_16843,N_16542,N_16117);
and U16844 (N_16844,N_16738,N_15829);
and U16845 (N_16845,N_16369,N_16701);
or U16846 (N_16846,N_16696,N_16509);
nand U16847 (N_16847,N_16620,N_16471);
nand U16848 (N_16848,N_16037,N_16310);
nor U16849 (N_16849,N_15864,N_16632);
nor U16850 (N_16850,N_16570,N_15826);
nand U16851 (N_16851,N_16532,N_16357);
or U16852 (N_16852,N_16516,N_15745);
nor U16853 (N_16853,N_16569,N_16375);
xor U16854 (N_16854,N_16094,N_16276);
and U16855 (N_16855,N_16497,N_15911);
nor U16856 (N_16856,N_15721,N_15832);
and U16857 (N_16857,N_16285,N_16724);
xor U16858 (N_16858,N_15661,N_16031);
and U16859 (N_16859,N_16694,N_16534);
and U16860 (N_16860,N_16245,N_16476);
and U16861 (N_16861,N_15933,N_16562);
and U16862 (N_16862,N_16517,N_15938);
xnor U16863 (N_16863,N_16759,N_16734);
or U16864 (N_16864,N_16281,N_16279);
nand U16865 (N_16865,N_15646,N_15635);
and U16866 (N_16866,N_16490,N_15610);
nand U16867 (N_16867,N_16480,N_15613);
nor U16868 (N_16868,N_16544,N_15840);
or U16869 (N_16869,N_16048,N_16530);
and U16870 (N_16870,N_16664,N_15991);
nand U16871 (N_16871,N_16300,N_16609);
nor U16872 (N_16872,N_16441,N_16359);
nand U16873 (N_16873,N_15885,N_16271);
xor U16874 (N_16874,N_16226,N_16392);
nor U16875 (N_16875,N_16102,N_15709);
nor U16876 (N_16876,N_15784,N_15898);
and U16877 (N_16877,N_16697,N_16501);
nor U16878 (N_16878,N_16019,N_16539);
and U16879 (N_16879,N_16447,N_16555);
nand U16880 (N_16880,N_15619,N_16091);
or U16881 (N_16881,N_16443,N_16202);
nand U16882 (N_16882,N_16421,N_15980);
or U16883 (N_16883,N_16365,N_16280);
nor U16884 (N_16884,N_15710,N_16009);
nand U16885 (N_16885,N_15778,N_16698);
or U16886 (N_16886,N_15960,N_15645);
or U16887 (N_16887,N_15887,N_16690);
or U16888 (N_16888,N_15999,N_16084);
nor U16889 (N_16889,N_15948,N_16751);
nand U16890 (N_16890,N_15804,N_16433);
xor U16891 (N_16891,N_15757,N_16042);
or U16892 (N_16892,N_16686,N_15644);
nand U16893 (N_16893,N_15724,N_15970);
nand U16894 (N_16894,N_16060,N_16435);
or U16895 (N_16895,N_16722,N_16248);
xor U16896 (N_16896,N_15701,N_16641);
nor U16897 (N_16897,N_15748,N_16670);
nor U16898 (N_16898,N_16651,N_16304);
nand U16899 (N_16899,N_16715,N_16049);
or U16900 (N_16900,N_15608,N_15663);
xor U16901 (N_16901,N_16229,N_16201);
xnor U16902 (N_16902,N_15954,N_16629);
nor U16903 (N_16903,N_16762,N_16788);
xnor U16904 (N_16904,N_16186,N_15637);
or U16905 (N_16905,N_16345,N_15725);
or U16906 (N_16906,N_16429,N_16437);
nor U16907 (N_16907,N_16073,N_16370);
nand U16908 (N_16908,N_16470,N_16381);
nand U16909 (N_16909,N_16288,N_15830);
nor U16910 (N_16910,N_16126,N_16234);
xor U16911 (N_16911,N_16712,N_16156);
and U16912 (N_16912,N_16169,N_15897);
xor U16913 (N_16913,N_16753,N_16572);
nand U16914 (N_16914,N_16247,N_16554);
nand U16915 (N_16915,N_16536,N_16538);
xnor U16916 (N_16916,N_16233,N_16332);
and U16917 (N_16917,N_15975,N_16395);
nand U16918 (N_16918,N_16356,N_16565);
xor U16919 (N_16919,N_16765,N_15681);
nor U16920 (N_16920,N_16790,N_15769);
nor U16921 (N_16921,N_16595,N_16654);
nand U16922 (N_16922,N_16377,N_16373);
or U16923 (N_16923,N_15951,N_15882);
or U16924 (N_16924,N_16504,N_16016);
nand U16925 (N_16925,N_15825,N_16294);
xor U16926 (N_16926,N_16462,N_15865);
nand U16927 (N_16927,N_16030,N_16749);
or U16928 (N_16928,N_16071,N_16723);
or U16929 (N_16929,N_15861,N_16191);
nand U16930 (N_16930,N_15672,N_16623);
and U16931 (N_16931,N_15845,N_16695);
and U16932 (N_16932,N_15767,N_16218);
nand U16933 (N_16933,N_16023,N_16334);
and U16934 (N_16934,N_16107,N_16702);
xor U16935 (N_16935,N_15766,N_15969);
nor U16936 (N_16936,N_15943,N_16321);
nor U16937 (N_16937,N_16436,N_16237);
xnor U16938 (N_16938,N_16183,N_16479);
xnor U16939 (N_16939,N_16070,N_16127);
nor U16940 (N_16940,N_15787,N_15746);
and U16941 (N_16941,N_16333,N_16590);
nand U16942 (N_16942,N_16747,N_16648);
nand U16943 (N_16943,N_16363,N_16543);
and U16944 (N_16944,N_16610,N_15878);
nand U16945 (N_16945,N_16401,N_15922);
nor U16946 (N_16946,N_15723,N_16272);
xnor U16947 (N_16947,N_16510,N_15881);
xnor U16948 (N_16948,N_16215,N_16013);
xnor U16949 (N_16949,N_16062,N_16038);
and U16950 (N_16950,N_16061,N_16305);
nor U16951 (N_16951,N_16262,N_16151);
xnor U16952 (N_16952,N_15817,N_15913);
xnor U16953 (N_16953,N_15989,N_16598);
nor U16954 (N_16954,N_16768,N_15850);
and U16955 (N_16955,N_15696,N_16467);
and U16956 (N_16956,N_15744,N_16647);
or U16957 (N_16957,N_15920,N_16740);
nand U16958 (N_16958,N_16054,N_15666);
xor U16959 (N_16959,N_16133,N_16637);
nor U16960 (N_16960,N_16491,N_15628);
and U16961 (N_16961,N_15947,N_15973);
or U16962 (N_16962,N_16605,N_16385);
or U16963 (N_16963,N_16529,N_15717);
or U16964 (N_16964,N_16707,N_15722);
or U16965 (N_16965,N_16082,N_16779);
and U16966 (N_16966,N_16258,N_15629);
nor U16967 (N_16967,N_16228,N_15956);
xor U16968 (N_16968,N_16167,N_16742);
nand U16969 (N_16969,N_16594,N_16130);
nand U16970 (N_16970,N_15994,N_15893);
nand U16971 (N_16971,N_16604,N_15877);
xor U16972 (N_16972,N_16044,N_16175);
nor U16973 (N_16973,N_16064,N_15702);
and U16974 (N_16974,N_16001,N_16549);
and U16975 (N_16975,N_15823,N_15713);
or U16976 (N_16976,N_16018,N_15946);
xor U16977 (N_16977,N_15961,N_16282);
nor U16978 (N_16978,N_16662,N_16685);
or U16979 (N_16979,N_15821,N_16705);
nand U16980 (N_16980,N_15729,N_16521);
xnor U16981 (N_16981,N_16780,N_16118);
or U16982 (N_16982,N_16209,N_16242);
nand U16983 (N_16983,N_16492,N_16726);
or U16984 (N_16984,N_16511,N_15662);
xor U16985 (N_16985,N_15670,N_16618);
or U16986 (N_16986,N_15914,N_16227);
or U16987 (N_16987,N_16100,N_16564);
and U16988 (N_16988,N_16177,N_15602);
or U16989 (N_16989,N_15750,N_16464);
and U16990 (N_16990,N_16525,N_15658);
xnor U16991 (N_16991,N_16125,N_16307);
and U16992 (N_16992,N_16302,N_16550);
or U16993 (N_16993,N_15867,N_16646);
nor U16994 (N_16994,N_15698,N_15976);
nand U16995 (N_16995,N_15799,N_16643);
nand U16996 (N_16996,N_16568,N_16354);
nand U16997 (N_16997,N_16444,N_16092);
and U16998 (N_16998,N_16195,N_16355);
and U16999 (N_16999,N_15945,N_16541);
xor U17000 (N_17000,N_16663,N_15689);
nor U17001 (N_17001,N_16261,N_16022);
or U17002 (N_17002,N_16291,N_16159);
or U17003 (N_17003,N_16330,N_15952);
xor U17004 (N_17004,N_15773,N_16396);
xor U17005 (N_17005,N_15622,N_15874);
nor U17006 (N_17006,N_16170,N_16010);
nor U17007 (N_17007,N_15718,N_15939);
xnor U17008 (N_17008,N_15692,N_15909);
nor U17009 (N_17009,N_16344,N_15653);
xor U17010 (N_17010,N_16434,N_16526);
or U17011 (N_17011,N_15794,N_15866);
nand U17012 (N_17012,N_15682,N_16412);
nor U17013 (N_17013,N_16556,N_16376);
xor U17014 (N_17014,N_15782,N_16413);
nor U17015 (N_17015,N_16393,N_16756);
or U17016 (N_17016,N_16131,N_16484);
nand U17017 (N_17017,N_15899,N_15621);
nand U17018 (N_17018,N_16257,N_16505);
xnor U17019 (N_17019,N_15932,N_16074);
or U17020 (N_17020,N_15798,N_16210);
xnor U17021 (N_17021,N_16140,N_15906);
nand U17022 (N_17022,N_16661,N_15754);
xnor U17023 (N_17023,N_16457,N_16194);
and U17024 (N_17024,N_16003,N_16224);
nand U17025 (N_17025,N_16111,N_16507);
nor U17026 (N_17026,N_15732,N_15719);
or U17027 (N_17027,N_16253,N_16522);
nand U17028 (N_17028,N_16653,N_15679);
nor U17029 (N_17029,N_15786,N_16329);
or U17030 (N_17030,N_15998,N_15925);
and U17031 (N_17031,N_15983,N_16587);
nor U17032 (N_17032,N_16736,N_16750);
and U17033 (N_17033,N_15796,N_16383);
nand U17034 (N_17034,N_15923,N_15981);
nand U17035 (N_17035,N_15634,N_16056);
nor U17036 (N_17036,N_15985,N_16277);
nand U17037 (N_17037,N_15751,N_16297);
or U17038 (N_17038,N_16573,N_16085);
nor U17039 (N_17039,N_15901,N_16136);
or U17040 (N_17040,N_15953,N_15736);
nand U17041 (N_17041,N_16639,N_15731);
nor U17042 (N_17042,N_16113,N_16523);
xor U17043 (N_17043,N_16625,N_15756);
or U17044 (N_17044,N_15673,N_16551);
or U17045 (N_17045,N_16442,N_16265);
xor U17046 (N_17046,N_15706,N_15912);
nor U17047 (N_17047,N_16399,N_15802);
or U17048 (N_17048,N_16287,N_16578);
or U17049 (N_17049,N_15684,N_16745);
nand U17050 (N_17050,N_16027,N_16179);
or U17051 (N_17051,N_16496,N_16152);
nor U17052 (N_17052,N_15889,N_16489);
and U17053 (N_17053,N_15620,N_16764);
nor U17054 (N_17054,N_16181,N_15810);
xnor U17055 (N_17055,N_16459,N_15765);
nand U17056 (N_17056,N_16577,N_16090);
xor U17057 (N_17057,N_16097,N_15781);
xnor U17058 (N_17058,N_16767,N_16290);
and U17059 (N_17059,N_16314,N_16386);
nor U17060 (N_17060,N_15824,N_16600);
nor U17061 (N_17061,N_16431,N_15971);
xor U17062 (N_17062,N_16089,N_16350);
and U17063 (N_17063,N_16483,N_16217);
nor U17064 (N_17064,N_16164,N_15926);
and U17065 (N_17065,N_16711,N_15642);
nand U17066 (N_17066,N_16340,N_15842);
or U17067 (N_17067,N_16408,N_16752);
nor U17068 (N_17068,N_16174,N_15915);
xor U17069 (N_17069,N_15903,N_15785);
and U17070 (N_17070,N_15779,N_15838);
and U17071 (N_17071,N_16046,N_16624);
nand U17072 (N_17072,N_16098,N_15836);
nor U17073 (N_17073,N_16360,N_15605);
nor U17074 (N_17074,N_16667,N_16755);
nor U17075 (N_17075,N_15603,N_15737);
nor U17076 (N_17076,N_15942,N_16109);
nand U17077 (N_17077,N_16093,N_15807);
nor U17078 (N_17078,N_16727,N_16256);
or U17079 (N_17079,N_16208,N_16405);
or U17080 (N_17080,N_16675,N_16692);
xor U17081 (N_17081,N_15630,N_16419);
or U17082 (N_17082,N_16766,N_16087);
nor U17083 (N_17083,N_16137,N_16791);
nand U17084 (N_17084,N_16628,N_15918);
nor U17085 (N_17085,N_16239,N_15996);
or U17086 (N_17086,N_15879,N_16485);
nand U17087 (N_17087,N_16083,N_16477);
xor U17088 (N_17088,N_16771,N_16558);
xor U17089 (N_17089,N_16424,N_16672);
xnor U17090 (N_17090,N_15789,N_16487);
nand U17091 (N_17091,N_15927,N_16458);
nor U17092 (N_17092,N_15966,N_16583);
nor U17093 (N_17093,N_16728,N_16785);
and U17094 (N_17094,N_16591,N_15660);
xnor U17095 (N_17095,N_15924,N_16077);
or U17096 (N_17096,N_16739,N_16472);
xor U17097 (N_17097,N_15809,N_15631);
and U17098 (N_17098,N_16200,N_16295);
nor U17099 (N_17099,N_15822,N_16537);
nand U17100 (N_17100,N_16041,N_16409);
or U17101 (N_17101,N_16335,N_16799);
and U17102 (N_17102,N_15959,N_16754);
xor U17103 (N_17103,N_16189,N_16361);
nor U17104 (N_17104,N_16222,N_16216);
or U17105 (N_17105,N_16518,N_16270);
xor U17106 (N_17106,N_16602,N_16576);
nor U17107 (N_17107,N_16006,N_15955);
and U17108 (N_17108,N_16708,N_16328);
and U17109 (N_17109,N_15931,N_16076);
and U17110 (N_17110,N_16427,N_15664);
nand U17111 (N_17111,N_15636,N_15868);
and U17112 (N_17112,N_16473,N_16631);
and U17113 (N_17113,N_15690,N_16124);
nand U17114 (N_17114,N_15848,N_15856);
nand U17115 (N_17115,N_16184,N_15738);
or U17116 (N_17116,N_16545,N_15900);
nand U17117 (N_17117,N_16422,N_15820);
or U17118 (N_17118,N_16153,N_15740);
or U17119 (N_17119,N_15654,N_16327);
or U17120 (N_17120,N_15873,N_16450);
nand U17121 (N_17121,N_15668,N_16508);
or U17122 (N_17122,N_16668,N_16081);
or U17123 (N_17123,N_16225,N_15703);
or U17124 (N_17124,N_15680,N_16410);
or U17125 (N_17125,N_15940,N_15678);
and U17126 (N_17126,N_15806,N_15683);
nor U17127 (N_17127,N_16095,N_15919);
and U17128 (N_17128,N_16634,N_16086);
or U17129 (N_17129,N_16246,N_15651);
or U17130 (N_17130,N_16353,N_16260);
and U17131 (N_17131,N_16561,N_16772);
nor U17132 (N_17132,N_16687,N_15855);
nor U17133 (N_17133,N_16255,N_15614);
or U17134 (N_17134,N_16787,N_15640);
nand U17135 (N_17135,N_16283,N_16559);
nand U17136 (N_17136,N_16254,N_16389);
and U17137 (N_17137,N_15803,N_16718);
nand U17138 (N_17138,N_16371,N_16721);
xnor U17139 (N_17139,N_16683,N_16557);
xnor U17140 (N_17140,N_16730,N_15854);
nor U17141 (N_17141,N_16002,N_15761);
xor U17142 (N_17142,N_15852,N_16415);
and U17143 (N_17143,N_15984,N_16123);
and U17144 (N_17144,N_15958,N_16778);
nor U17145 (N_17145,N_16364,N_16252);
nor U17146 (N_17146,N_16051,N_16552);
nor U17147 (N_17147,N_16158,N_16691);
xor U17148 (N_17148,N_16223,N_16374);
nand U17149 (N_17149,N_16417,N_16299);
xnor U17150 (N_17150,N_16420,N_15601);
nand U17151 (N_17151,N_15941,N_16005);
and U17152 (N_17152,N_15699,N_16045);
and U17153 (N_17153,N_15727,N_16703);
nand U17154 (N_17154,N_16599,N_16238);
nor U17155 (N_17155,N_15929,N_16744);
nand U17156 (N_17156,N_16055,N_16678);
xnor U17157 (N_17157,N_15711,N_16533);
xor U17158 (N_17158,N_15650,N_16676);
xnor U17159 (N_17159,N_15657,N_16432);
nand U17160 (N_17160,N_16400,N_16372);
nand U17161 (N_17161,N_15775,N_16068);
nor U17162 (N_17162,N_16700,N_15977);
nand U17163 (N_17163,N_15851,N_16581);
and U17164 (N_17164,N_16250,N_15624);
or U17165 (N_17165,N_16358,N_16622);
nor U17166 (N_17166,N_15997,N_16197);
or U17167 (N_17167,N_16148,N_16313);
nand U17168 (N_17168,N_16154,N_16449);
nor U17169 (N_17169,N_16007,N_16112);
xor U17170 (N_17170,N_15978,N_15808);
nand U17171 (N_17171,N_16560,N_15895);
and U17172 (N_17172,N_15655,N_16176);
nand U17173 (N_17173,N_16713,N_15693);
and U17174 (N_17174,N_16677,N_16161);
and U17175 (N_17175,N_16021,N_15675);
xor U17176 (N_17176,N_16000,N_15712);
xor U17177 (N_17177,N_15801,N_15749);
xnor U17178 (N_17178,N_16714,N_15758);
or U17179 (N_17179,N_16786,N_15780);
and U17180 (N_17180,N_16269,N_16394);
nor U17181 (N_17181,N_16387,N_16655);
and U17182 (N_17182,N_16162,N_16193);
nor U17183 (N_17183,N_16075,N_16579);
and U17184 (N_17184,N_15735,N_16289);
xor U17185 (N_17185,N_15704,N_16585);
nor U17186 (N_17186,N_16035,N_16214);
and U17187 (N_17187,N_16199,N_15627);
xnor U17188 (N_17188,N_16660,N_16249);
xor U17189 (N_17189,N_15990,N_16292);
nor U17190 (N_17190,N_15728,N_16757);
nor U17191 (N_17191,N_16352,N_16286);
nor U17192 (N_17192,N_15859,N_16466);
xnor U17193 (N_17193,N_16612,N_15659);
and U17194 (N_17194,N_15726,N_16104);
nand U17195 (N_17195,N_15714,N_16145);
nand U17196 (N_17196,N_16339,N_15949);
and U17197 (N_17197,N_16635,N_16735);
nor U17198 (N_17198,N_16567,N_16318);
xnor U17199 (N_17199,N_16777,N_16157);
and U17200 (N_17200,N_16182,N_16627);
or U17201 (N_17201,N_15858,N_16582);
nor U17202 (N_17202,N_16284,N_15774);
or U17203 (N_17203,N_16793,N_15857);
nor U17204 (N_17204,N_15812,N_16106);
and U17205 (N_17205,N_16101,N_15791);
and U17206 (N_17206,N_16719,N_16207);
nor U17207 (N_17207,N_16213,N_16240);
nor U17208 (N_17208,N_16425,N_16155);
or U17209 (N_17209,N_15884,N_16451);
or U17210 (N_17210,N_16263,N_16129);
xnor U17211 (N_17211,N_16122,N_16760);
xor U17212 (N_17212,N_16273,N_15697);
nand U17213 (N_17213,N_16047,N_15609);
or U17214 (N_17214,N_16528,N_15793);
xnor U17215 (N_17215,N_16043,N_15705);
and U17216 (N_17216,N_16192,N_15649);
nand U17217 (N_17217,N_16398,N_15768);
nor U17218 (N_17218,N_16034,N_16614);
and U17219 (N_17219,N_16445,N_16236);
nor U17220 (N_17220,N_16020,N_15910);
or U17221 (N_17221,N_15988,N_16346);
nand U17222 (N_17222,N_15875,N_15993);
nand U17223 (N_17223,N_15888,N_15695);
nor U17224 (N_17224,N_16187,N_15730);
nand U17225 (N_17225,N_16774,N_16453);
nor U17226 (N_17226,N_15600,N_15734);
or U17227 (N_17227,N_15760,N_16789);
and U17228 (N_17228,N_16776,N_16134);
or U17229 (N_17229,N_16584,N_16657);
and U17230 (N_17230,N_15834,N_16601);
or U17231 (N_17231,N_15896,N_15916);
nand U17232 (N_17232,N_15671,N_16278);
and U17233 (N_17233,N_15853,N_16172);
or U17234 (N_17234,N_16232,N_15677);
or U17235 (N_17235,N_15676,N_16315);
nor U17236 (N_17236,N_16666,N_15921);
and U17237 (N_17237,N_15687,N_16688);
and U17238 (N_17238,N_16468,N_15752);
or U17239 (N_17239,N_15776,N_15816);
nor U17240 (N_17240,N_16729,N_16241);
or U17241 (N_17241,N_16308,N_16326);
and U17242 (N_17242,N_16275,N_16781);
and U17243 (N_17243,N_15771,N_16379);
xor U17244 (N_17244,N_16546,N_16469);
xnor U17245 (N_17245,N_15759,N_16580);
and U17246 (N_17246,N_15652,N_15905);
and U17247 (N_17247,N_16004,N_16717);
nand U17248 (N_17248,N_15643,N_16141);
xnor U17249 (N_17249,N_16519,N_15691);
nand U17250 (N_17250,N_15638,N_16196);
or U17251 (N_17251,N_15962,N_16115);
and U17252 (N_17252,N_16699,N_16050);
nand U17253 (N_17253,N_16486,N_15950);
nand U17254 (N_17254,N_16474,N_15869);
and U17255 (N_17255,N_16630,N_16312);
and U17256 (N_17256,N_16748,N_16325);
and U17257 (N_17257,N_16796,N_16150);
or U17258 (N_17258,N_16650,N_16619);
xor U17259 (N_17259,N_16535,N_16725);
nand U17260 (N_17260,N_16482,N_15633);
and U17261 (N_17261,N_16072,N_16642);
or U17262 (N_17262,N_16163,N_16014);
nand U17263 (N_17263,N_16058,N_16430);
xnor U17264 (N_17264,N_16524,N_15763);
nor U17265 (N_17265,N_15783,N_16397);
nor U17266 (N_17266,N_16204,N_16571);
nand U17267 (N_17267,N_16040,N_16682);
nand U17268 (N_17268,N_16171,N_16033);
xnor U17269 (N_17269,N_15790,N_16180);
xor U17270 (N_17270,N_16652,N_16121);
and U17271 (N_17271,N_16795,N_16012);
xnor U17272 (N_17272,N_16311,N_15847);
nor U17273 (N_17273,N_16319,N_16331);
xor U17274 (N_17274,N_16298,N_16024);
xor U17275 (N_17275,N_15908,N_15615);
nand U17276 (N_17276,N_16783,N_16211);
and U17277 (N_17277,N_16540,N_15907);
and U17278 (N_17278,N_15688,N_16065);
or U17279 (N_17279,N_16710,N_15986);
xor U17280 (N_17280,N_15862,N_16452);
nand U17281 (N_17281,N_16132,N_16382);
or U17282 (N_17282,N_15741,N_16784);
nand U17283 (N_17283,N_15937,N_16669);
or U17284 (N_17284,N_15639,N_16704);
nor U17285 (N_17285,N_16078,N_16640);
or U17286 (N_17286,N_16566,N_15707);
or U17287 (N_17287,N_16110,N_16165);
xnor U17288 (N_17288,N_16028,N_16388);
and U17289 (N_17289,N_15813,N_16680);
xnor U17290 (N_17290,N_16105,N_16498);
or U17291 (N_17291,N_16716,N_16782);
and U17292 (N_17292,N_16178,N_15828);
nor U17293 (N_17293,N_16293,N_15604);
nor U17294 (N_17294,N_16029,N_15987);
and U17295 (N_17295,N_15700,N_16720);
nand U17296 (N_17296,N_15883,N_16166);
xor U17297 (N_17297,N_16512,N_16366);
and U17298 (N_17298,N_15968,N_16411);
xnor U17299 (N_17299,N_16770,N_16135);
and U17300 (N_17300,N_15979,N_15995);
xnor U17301 (N_17301,N_16506,N_16743);
nor U17302 (N_17302,N_16015,N_16120);
or U17303 (N_17303,N_16244,N_15934);
xor U17304 (N_17304,N_16475,N_16636);
nor U17305 (N_17305,N_16188,N_16142);
and U17306 (N_17306,N_16052,N_16378);
and U17307 (N_17307,N_16741,N_15972);
xor U17308 (N_17308,N_15770,N_15835);
and U17309 (N_17309,N_15814,N_15872);
and U17310 (N_17310,N_15685,N_15792);
nand U17311 (N_17311,N_16426,N_16527);
nand U17312 (N_17312,N_15818,N_16205);
or U17313 (N_17313,N_15611,N_16323);
xor U17314 (N_17314,N_16347,N_15647);
xnor U17315 (N_17315,N_16548,N_16732);
nand U17316 (N_17316,N_16349,N_16108);
and U17317 (N_17317,N_16198,N_15777);
nor U17318 (N_17318,N_16221,N_16251);
nor U17319 (N_17319,N_15764,N_16185);
nand U17320 (N_17320,N_16059,N_15944);
nand U17321 (N_17321,N_16147,N_16593);
or U17322 (N_17322,N_15833,N_16231);
nor U17323 (N_17323,N_16465,N_16139);
nand U17324 (N_17324,N_16168,N_15886);
xor U17325 (N_17325,N_15607,N_16266);
nand U17326 (N_17326,N_16220,N_15674);
xor U17327 (N_17327,N_16402,N_16067);
or U17328 (N_17328,N_16495,N_16460);
xnor U17329 (N_17329,N_15967,N_16645);
and U17330 (N_17330,N_16665,N_15963);
xnor U17331 (N_17331,N_16025,N_15747);
or U17332 (N_17332,N_15669,N_16502);
nor U17333 (N_17333,N_16586,N_16611);
nor U17334 (N_17334,N_16679,N_16368);
and U17335 (N_17335,N_16455,N_16384);
or U17336 (N_17336,N_16428,N_16440);
xnor U17337 (N_17337,N_16439,N_16138);
and U17338 (N_17338,N_15617,N_16337);
nor U17339 (N_17339,N_15648,N_16606);
xnor U17340 (N_17340,N_16119,N_16589);
nor U17341 (N_17341,N_16342,N_16309);
and U17342 (N_17342,N_16659,N_16322);
or U17343 (N_17343,N_16267,N_15616);
xnor U17344 (N_17344,N_16303,N_15860);
nor U17345 (N_17345,N_16160,N_16797);
nand U17346 (N_17346,N_16514,N_16203);
or U17347 (N_17347,N_15827,N_16626);
and U17348 (N_17348,N_15715,N_16341);
or U17349 (N_17349,N_15815,N_15892);
xnor U17350 (N_17350,N_16649,N_15904);
nor U17351 (N_17351,N_16621,N_16414);
or U17352 (N_17352,N_16456,N_15788);
xnor U17353 (N_17353,N_16438,N_15762);
xor U17354 (N_17354,N_16461,N_16173);
or U17355 (N_17355,N_16011,N_16219);
xnor U17356 (N_17356,N_16775,N_16066);
or U17357 (N_17357,N_16390,N_15902);
or U17358 (N_17358,N_15716,N_16088);
or U17359 (N_17359,N_16773,N_16674);
or U17360 (N_17360,N_16603,N_16206);
xor U17361 (N_17361,N_16481,N_15606);
xnor U17362 (N_17362,N_15708,N_15819);
or U17363 (N_17363,N_16644,N_16306);
and U17364 (N_17364,N_16080,N_16794);
and U17365 (N_17365,N_15890,N_15957);
nand U17366 (N_17366,N_16296,N_16403);
nand U17367 (N_17367,N_16488,N_16763);
nand U17368 (N_17368,N_15641,N_16144);
and U17369 (N_17369,N_16574,N_16128);
nor U17370 (N_17370,N_16039,N_16380);
xnor U17371 (N_17371,N_15626,N_16684);
nand U17372 (N_17372,N_16658,N_15753);
and U17373 (N_17373,N_16026,N_16230);
nand U17374 (N_17374,N_16032,N_16317);
xor U17375 (N_17375,N_16063,N_15805);
and U17376 (N_17376,N_16336,N_15618);
and U17377 (N_17377,N_15667,N_16404);
or U17378 (N_17378,N_16143,N_16617);
nor U17379 (N_17379,N_16673,N_15743);
nand U17380 (N_17380,N_16017,N_16338);
nor U17381 (N_17381,N_15841,N_16149);
and U17382 (N_17382,N_16769,N_15880);
xnor U17383 (N_17383,N_15843,N_16324);
and U17384 (N_17384,N_16190,N_16418);
and U17385 (N_17385,N_16592,N_15755);
or U17386 (N_17386,N_15797,N_15625);
nor U17387 (N_17387,N_16733,N_16500);
nand U17388 (N_17388,N_16563,N_16268);
or U17389 (N_17389,N_15917,N_16706);
nor U17390 (N_17390,N_15992,N_16116);
nand U17391 (N_17391,N_16235,N_16212);
or U17392 (N_17392,N_15623,N_16607);
nor U17393 (N_17393,N_16259,N_16057);
nor U17394 (N_17394,N_15839,N_16301);
and U17395 (N_17395,N_15800,N_16103);
nor U17396 (N_17396,N_16416,N_16588);
and U17397 (N_17397,N_15811,N_15632);
and U17398 (N_17398,N_15656,N_16096);
nand U17399 (N_17399,N_15871,N_15876);
xnor U17400 (N_17400,N_16214,N_15665);
and U17401 (N_17401,N_16718,N_16700);
nand U17402 (N_17402,N_15898,N_16428);
nor U17403 (N_17403,N_16160,N_15717);
xor U17404 (N_17404,N_16427,N_16755);
and U17405 (N_17405,N_16290,N_16581);
xor U17406 (N_17406,N_16046,N_16747);
nor U17407 (N_17407,N_15765,N_15629);
nand U17408 (N_17408,N_15754,N_16188);
nand U17409 (N_17409,N_16473,N_15604);
xnor U17410 (N_17410,N_15943,N_15661);
nor U17411 (N_17411,N_15919,N_16689);
nand U17412 (N_17412,N_16723,N_16019);
and U17413 (N_17413,N_15671,N_16233);
nor U17414 (N_17414,N_15934,N_16278);
nand U17415 (N_17415,N_16215,N_16388);
xnor U17416 (N_17416,N_16268,N_16544);
and U17417 (N_17417,N_15805,N_15849);
nor U17418 (N_17418,N_16174,N_15749);
nor U17419 (N_17419,N_16367,N_15811);
nor U17420 (N_17420,N_15985,N_16790);
and U17421 (N_17421,N_15989,N_16086);
nor U17422 (N_17422,N_16687,N_16342);
nor U17423 (N_17423,N_16586,N_16457);
or U17424 (N_17424,N_16776,N_15631);
or U17425 (N_17425,N_15706,N_16296);
nand U17426 (N_17426,N_16666,N_15674);
and U17427 (N_17427,N_16628,N_16078);
xor U17428 (N_17428,N_16198,N_16133);
xor U17429 (N_17429,N_15802,N_15618);
nor U17430 (N_17430,N_16079,N_15714);
and U17431 (N_17431,N_15956,N_16384);
nor U17432 (N_17432,N_16549,N_15624);
nand U17433 (N_17433,N_16053,N_16321);
xnor U17434 (N_17434,N_15795,N_16719);
xor U17435 (N_17435,N_15923,N_16605);
xor U17436 (N_17436,N_16237,N_15772);
xnor U17437 (N_17437,N_16634,N_15762);
nor U17438 (N_17438,N_16445,N_16618);
nor U17439 (N_17439,N_15921,N_16304);
and U17440 (N_17440,N_16127,N_15677);
xor U17441 (N_17441,N_16231,N_15888);
and U17442 (N_17442,N_16793,N_15994);
nand U17443 (N_17443,N_16073,N_16150);
nor U17444 (N_17444,N_15674,N_16696);
nand U17445 (N_17445,N_16601,N_16040);
or U17446 (N_17446,N_16331,N_16714);
nor U17447 (N_17447,N_16283,N_16634);
nor U17448 (N_17448,N_16207,N_16026);
nor U17449 (N_17449,N_15726,N_15801);
and U17450 (N_17450,N_15651,N_15741);
nand U17451 (N_17451,N_16394,N_16785);
nor U17452 (N_17452,N_16340,N_15962);
nand U17453 (N_17453,N_16210,N_16266);
nand U17454 (N_17454,N_15972,N_16377);
nor U17455 (N_17455,N_16113,N_16546);
nand U17456 (N_17456,N_16379,N_16414);
or U17457 (N_17457,N_16232,N_16473);
or U17458 (N_17458,N_16383,N_16080);
or U17459 (N_17459,N_16059,N_15963);
and U17460 (N_17460,N_16361,N_16496);
or U17461 (N_17461,N_16604,N_16388);
xor U17462 (N_17462,N_15909,N_16763);
and U17463 (N_17463,N_15901,N_15603);
and U17464 (N_17464,N_16390,N_15808);
and U17465 (N_17465,N_16127,N_15804);
nor U17466 (N_17466,N_15830,N_16778);
nand U17467 (N_17467,N_15801,N_16058);
nor U17468 (N_17468,N_16023,N_16256);
or U17469 (N_17469,N_15600,N_16789);
and U17470 (N_17470,N_15682,N_15822);
and U17471 (N_17471,N_15899,N_16347);
xnor U17472 (N_17472,N_16579,N_16180);
xor U17473 (N_17473,N_16544,N_16267);
nand U17474 (N_17474,N_16048,N_16437);
nand U17475 (N_17475,N_16576,N_16048);
and U17476 (N_17476,N_16213,N_16214);
nor U17477 (N_17477,N_15669,N_16220);
or U17478 (N_17478,N_16514,N_15620);
nor U17479 (N_17479,N_16773,N_16519);
xor U17480 (N_17480,N_16443,N_15811);
or U17481 (N_17481,N_16099,N_15627);
and U17482 (N_17482,N_16735,N_16310);
xnor U17483 (N_17483,N_16510,N_15665);
xor U17484 (N_17484,N_16093,N_16322);
nor U17485 (N_17485,N_15742,N_16339);
and U17486 (N_17486,N_16023,N_15944);
xor U17487 (N_17487,N_15681,N_16528);
or U17488 (N_17488,N_16158,N_16299);
nand U17489 (N_17489,N_15843,N_16774);
and U17490 (N_17490,N_15790,N_16636);
nor U17491 (N_17491,N_15952,N_16463);
xor U17492 (N_17492,N_16180,N_16707);
and U17493 (N_17493,N_16707,N_16659);
nor U17494 (N_17494,N_15843,N_16112);
nor U17495 (N_17495,N_16350,N_16614);
nor U17496 (N_17496,N_15638,N_16673);
xnor U17497 (N_17497,N_16184,N_15622);
xor U17498 (N_17498,N_16596,N_15814);
nor U17499 (N_17499,N_16084,N_16320);
nor U17500 (N_17500,N_15779,N_15660);
xor U17501 (N_17501,N_15918,N_16346);
or U17502 (N_17502,N_15858,N_15987);
nor U17503 (N_17503,N_16597,N_16418);
nand U17504 (N_17504,N_16485,N_15655);
nor U17505 (N_17505,N_15700,N_15627);
or U17506 (N_17506,N_16264,N_16451);
nor U17507 (N_17507,N_16465,N_16694);
xor U17508 (N_17508,N_15634,N_16181);
or U17509 (N_17509,N_16626,N_16351);
nand U17510 (N_17510,N_16307,N_16475);
and U17511 (N_17511,N_15613,N_16134);
or U17512 (N_17512,N_16289,N_16124);
or U17513 (N_17513,N_15862,N_16100);
or U17514 (N_17514,N_15955,N_16147);
or U17515 (N_17515,N_16552,N_16547);
nand U17516 (N_17516,N_15811,N_16454);
and U17517 (N_17517,N_16433,N_15884);
or U17518 (N_17518,N_15796,N_16474);
nor U17519 (N_17519,N_16160,N_16616);
xor U17520 (N_17520,N_16249,N_15954);
xor U17521 (N_17521,N_16178,N_15689);
and U17522 (N_17522,N_16447,N_16330);
nor U17523 (N_17523,N_16377,N_16507);
and U17524 (N_17524,N_16417,N_16322);
xor U17525 (N_17525,N_16721,N_16775);
xor U17526 (N_17526,N_15642,N_16052);
xor U17527 (N_17527,N_16798,N_16532);
nor U17528 (N_17528,N_16649,N_15842);
nor U17529 (N_17529,N_16003,N_16187);
xnor U17530 (N_17530,N_15839,N_16348);
or U17531 (N_17531,N_16205,N_16301);
nand U17532 (N_17532,N_15661,N_16470);
nand U17533 (N_17533,N_15759,N_15793);
and U17534 (N_17534,N_16258,N_16341);
and U17535 (N_17535,N_15600,N_16102);
nor U17536 (N_17536,N_15765,N_16763);
nand U17537 (N_17537,N_16074,N_15877);
nand U17538 (N_17538,N_16649,N_16424);
or U17539 (N_17539,N_15802,N_16619);
nor U17540 (N_17540,N_16611,N_16107);
and U17541 (N_17541,N_15710,N_16092);
xor U17542 (N_17542,N_15702,N_15829);
nor U17543 (N_17543,N_15687,N_16024);
nand U17544 (N_17544,N_15685,N_15622);
xor U17545 (N_17545,N_16434,N_15895);
and U17546 (N_17546,N_16161,N_15802);
and U17547 (N_17547,N_15779,N_16585);
nor U17548 (N_17548,N_16021,N_16705);
xnor U17549 (N_17549,N_16697,N_16111);
nand U17550 (N_17550,N_15980,N_15747);
nor U17551 (N_17551,N_15971,N_16265);
or U17552 (N_17552,N_16048,N_15607);
xor U17553 (N_17553,N_15896,N_16162);
nor U17554 (N_17554,N_16387,N_16762);
or U17555 (N_17555,N_16086,N_15948);
nand U17556 (N_17556,N_16194,N_15715);
nand U17557 (N_17557,N_16461,N_16722);
and U17558 (N_17558,N_15953,N_15983);
nand U17559 (N_17559,N_16740,N_16391);
and U17560 (N_17560,N_16209,N_16681);
nand U17561 (N_17561,N_15650,N_16099);
or U17562 (N_17562,N_15767,N_16145);
or U17563 (N_17563,N_15823,N_16042);
or U17564 (N_17564,N_16290,N_16591);
and U17565 (N_17565,N_16681,N_16581);
or U17566 (N_17566,N_15802,N_15774);
nor U17567 (N_17567,N_16093,N_16669);
and U17568 (N_17568,N_16360,N_16579);
xnor U17569 (N_17569,N_15665,N_15750);
xor U17570 (N_17570,N_15955,N_16796);
or U17571 (N_17571,N_15835,N_16439);
nand U17572 (N_17572,N_16459,N_15789);
nand U17573 (N_17573,N_16092,N_15934);
xnor U17574 (N_17574,N_16027,N_15669);
nor U17575 (N_17575,N_15740,N_15950);
nor U17576 (N_17576,N_16602,N_16543);
nor U17577 (N_17577,N_16058,N_16246);
and U17578 (N_17578,N_16086,N_15691);
and U17579 (N_17579,N_16095,N_16364);
xor U17580 (N_17580,N_15857,N_15759);
xnor U17581 (N_17581,N_15916,N_15716);
nand U17582 (N_17582,N_16045,N_15854);
xnor U17583 (N_17583,N_15672,N_16650);
xnor U17584 (N_17584,N_16699,N_15902);
nand U17585 (N_17585,N_16230,N_15658);
nand U17586 (N_17586,N_16043,N_16272);
nor U17587 (N_17587,N_15959,N_16412);
nor U17588 (N_17588,N_16485,N_16362);
xnor U17589 (N_17589,N_15778,N_16463);
or U17590 (N_17590,N_15922,N_16265);
or U17591 (N_17591,N_16413,N_16362);
nor U17592 (N_17592,N_16516,N_16578);
nand U17593 (N_17593,N_16681,N_16247);
nand U17594 (N_17594,N_15849,N_15709);
xor U17595 (N_17595,N_16795,N_16496);
or U17596 (N_17596,N_15601,N_16144);
nor U17597 (N_17597,N_16283,N_16488);
xnor U17598 (N_17598,N_15751,N_16517);
nand U17599 (N_17599,N_16239,N_16651);
and U17600 (N_17600,N_16573,N_15952);
and U17601 (N_17601,N_16594,N_15804);
nand U17602 (N_17602,N_16175,N_16660);
or U17603 (N_17603,N_16007,N_16126);
nor U17604 (N_17604,N_15644,N_16470);
and U17605 (N_17605,N_16022,N_16794);
or U17606 (N_17606,N_15952,N_16092);
or U17607 (N_17607,N_16583,N_16215);
or U17608 (N_17608,N_15617,N_15717);
nor U17609 (N_17609,N_16232,N_16013);
or U17610 (N_17610,N_16423,N_16322);
and U17611 (N_17611,N_16374,N_16496);
nor U17612 (N_17612,N_16215,N_16705);
and U17613 (N_17613,N_15821,N_15845);
xor U17614 (N_17614,N_16034,N_15890);
or U17615 (N_17615,N_15764,N_16331);
nor U17616 (N_17616,N_15838,N_16285);
xnor U17617 (N_17617,N_15841,N_16701);
xor U17618 (N_17618,N_16091,N_16172);
xor U17619 (N_17619,N_15813,N_16411);
nand U17620 (N_17620,N_15656,N_16059);
and U17621 (N_17621,N_15632,N_16087);
and U17622 (N_17622,N_15912,N_16492);
nor U17623 (N_17623,N_16573,N_16799);
xnor U17624 (N_17624,N_16693,N_16262);
nand U17625 (N_17625,N_15953,N_16344);
nand U17626 (N_17626,N_16082,N_16099);
or U17627 (N_17627,N_15842,N_16431);
nor U17628 (N_17628,N_16019,N_15801);
nor U17629 (N_17629,N_15692,N_15740);
and U17630 (N_17630,N_15866,N_15930);
or U17631 (N_17631,N_15893,N_16216);
xnor U17632 (N_17632,N_15804,N_15685);
and U17633 (N_17633,N_16309,N_16053);
nor U17634 (N_17634,N_16265,N_16214);
or U17635 (N_17635,N_16377,N_15665);
nor U17636 (N_17636,N_15724,N_16314);
xnor U17637 (N_17637,N_16263,N_15892);
nor U17638 (N_17638,N_16025,N_16111);
and U17639 (N_17639,N_16419,N_16498);
nand U17640 (N_17640,N_16364,N_15675);
and U17641 (N_17641,N_15692,N_16119);
nand U17642 (N_17642,N_15656,N_16126);
or U17643 (N_17643,N_16598,N_16596);
nand U17644 (N_17644,N_16088,N_15930);
and U17645 (N_17645,N_16359,N_15855);
and U17646 (N_17646,N_15879,N_16291);
or U17647 (N_17647,N_16697,N_16736);
or U17648 (N_17648,N_16575,N_16411);
nor U17649 (N_17649,N_16049,N_16733);
or U17650 (N_17650,N_16095,N_16405);
or U17651 (N_17651,N_16167,N_15801);
or U17652 (N_17652,N_16655,N_16609);
or U17653 (N_17653,N_16141,N_15871);
nand U17654 (N_17654,N_16254,N_16686);
and U17655 (N_17655,N_16400,N_15979);
xnor U17656 (N_17656,N_16159,N_15991);
xor U17657 (N_17657,N_16167,N_16310);
and U17658 (N_17658,N_16291,N_15953);
or U17659 (N_17659,N_16159,N_16138);
nand U17660 (N_17660,N_16234,N_16557);
nor U17661 (N_17661,N_16453,N_15788);
nor U17662 (N_17662,N_16784,N_16598);
nor U17663 (N_17663,N_16426,N_16794);
and U17664 (N_17664,N_16402,N_15798);
nand U17665 (N_17665,N_16017,N_15683);
nor U17666 (N_17666,N_16790,N_15852);
nor U17667 (N_17667,N_16284,N_15831);
nand U17668 (N_17668,N_16799,N_15999);
and U17669 (N_17669,N_16710,N_16032);
nand U17670 (N_17670,N_16478,N_15721);
nor U17671 (N_17671,N_16092,N_15928);
or U17672 (N_17672,N_15755,N_15891);
or U17673 (N_17673,N_15866,N_16637);
nand U17674 (N_17674,N_15834,N_16172);
and U17675 (N_17675,N_16550,N_16119);
or U17676 (N_17676,N_16453,N_16163);
xor U17677 (N_17677,N_16530,N_15736);
or U17678 (N_17678,N_16464,N_16101);
or U17679 (N_17679,N_15896,N_15990);
nor U17680 (N_17680,N_16310,N_16791);
nor U17681 (N_17681,N_16217,N_16380);
nor U17682 (N_17682,N_16712,N_15654);
nand U17683 (N_17683,N_16224,N_16018);
and U17684 (N_17684,N_15849,N_16642);
nor U17685 (N_17685,N_16286,N_16345);
nand U17686 (N_17686,N_15617,N_16290);
xor U17687 (N_17687,N_15602,N_15909);
and U17688 (N_17688,N_16003,N_16430);
and U17689 (N_17689,N_16532,N_16171);
nand U17690 (N_17690,N_15869,N_15630);
xor U17691 (N_17691,N_16463,N_16784);
nand U17692 (N_17692,N_15916,N_16393);
nor U17693 (N_17693,N_15987,N_16630);
or U17694 (N_17694,N_16049,N_16657);
nor U17695 (N_17695,N_16023,N_15755);
nand U17696 (N_17696,N_16266,N_16698);
nand U17697 (N_17697,N_15767,N_15968);
or U17698 (N_17698,N_16488,N_15755);
nor U17699 (N_17699,N_15971,N_16449);
or U17700 (N_17700,N_16796,N_16516);
or U17701 (N_17701,N_16605,N_16759);
and U17702 (N_17702,N_15911,N_16106);
xnor U17703 (N_17703,N_16543,N_16463);
nor U17704 (N_17704,N_16283,N_16722);
xnor U17705 (N_17705,N_16772,N_16446);
xnor U17706 (N_17706,N_15749,N_16562);
and U17707 (N_17707,N_16194,N_16477);
nor U17708 (N_17708,N_15923,N_16450);
xor U17709 (N_17709,N_16532,N_16693);
nand U17710 (N_17710,N_16356,N_16649);
and U17711 (N_17711,N_16335,N_16219);
and U17712 (N_17712,N_16324,N_16678);
xor U17713 (N_17713,N_16295,N_16033);
nand U17714 (N_17714,N_15728,N_16358);
and U17715 (N_17715,N_16311,N_16331);
or U17716 (N_17716,N_16003,N_15789);
and U17717 (N_17717,N_15705,N_16047);
xnor U17718 (N_17718,N_16390,N_16596);
nor U17719 (N_17719,N_15962,N_16469);
nor U17720 (N_17720,N_16284,N_15770);
nor U17721 (N_17721,N_16532,N_16170);
nand U17722 (N_17722,N_15921,N_16297);
nand U17723 (N_17723,N_16289,N_16294);
and U17724 (N_17724,N_15953,N_15891);
or U17725 (N_17725,N_16673,N_16357);
or U17726 (N_17726,N_15692,N_16444);
or U17727 (N_17727,N_16622,N_16531);
and U17728 (N_17728,N_16671,N_16236);
and U17729 (N_17729,N_15739,N_16119);
nor U17730 (N_17730,N_15627,N_16583);
and U17731 (N_17731,N_16164,N_15608);
xnor U17732 (N_17732,N_15637,N_15819);
and U17733 (N_17733,N_15931,N_15750);
nor U17734 (N_17734,N_16084,N_16471);
nand U17735 (N_17735,N_16539,N_16023);
nand U17736 (N_17736,N_15612,N_16393);
nand U17737 (N_17737,N_16617,N_15629);
nand U17738 (N_17738,N_16439,N_15906);
xnor U17739 (N_17739,N_16584,N_16024);
and U17740 (N_17740,N_16150,N_15719);
nand U17741 (N_17741,N_15981,N_16347);
nand U17742 (N_17742,N_16225,N_16586);
xor U17743 (N_17743,N_15774,N_16533);
xnor U17744 (N_17744,N_15751,N_16129);
xnor U17745 (N_17745,N_16205,N_16402);
and U17746 (N_17746,N_16084,N_16260);
and U17747 (N_17747,N_16259,N_16085);
xor U17748 (N_17748,N_16072,N_15642);
nand U17749 (N_17749,N_16293,N_16531);
nand U17750 (N_17750,N_16658,N_16640);
or U17751 (N_17751,N_16334,N_16647);
and U17752 (N_17752,N_16230,N_15676);
nand U17753 (N_17753,N_16186,N_16400);
nor U17754 (N_17754,N_16256,N_16429);
nand U17755 (N_17755,N_16114,N_15852);
xnor U17756 (N_17756,N_16161,N_16135);
nand U17757 (N_17757,N_16109,N_16224);
and U17758 (N_17758,N_16148,N_16044);
or U17759 (N_17759,N_16363,N_16516);
or U17760 (N_17760,N_16234,N_16764);
and U17761 (N_17761,N_15908,N_16270);
and U17762 (N_17762,N_16538,N_16217);
nor U17763 (N_17763,N_15628,N_15804);
and U17764 (N_17764,N_15758,N_16109);
or U17765 (N_17765,N_16014,N_16618);
and U17766 (N_17766,N_15912,N_15657);
and U17767 (N_17767,N_16331,N_16405);
or U17768 (N_17768,N_15673,N_16309);
xnor U17769 (N_17769,N_16006,N_15697);
or U17770 (N_17770,N_15774,N_16787);
or U17771 (N_17771,N_16370,N_15778);
and U17772 (N_17772,N_15990,N_16743);
and U17773 (N_17773,N_15939,N_16472);
or U17774 (N_17774,N_16198,N_16361);
and U17775 (N_17775,N_15688,N_16386);
nor U17776 (N_17776,N_16710,N_16261);
or U17777 (N_17777,N_16155,N_16009);
nand U17778 (N_17778,N_16140,N_16031);
and U17779 (N_17779,N_16768,N_16023);
and U17780 (N_17780,N_15662,N_16631);
xor U17781 (N_17781,N_16612,N_16569);
or U17782 (N_17782,N_16078,N_16737);
nand U17783 (N_17783,N_16014,N_16612);
nand U17784 (N_17784,N_16582,N_16589);
and U17785 (N_17785,N_16033,N_16443);
nand U17786 (N_17786,N_16422,N_16794);
and U17787 (N_17787,N_16657,N_16678);
nor U17788 (N_17788,N_15882,N_16516);
xor U17789 (N_17789,N_16310,N_16688);
nor U17790 (N_17790,N_16266,N_16582);
and U17791 (N_17791,N_16353,N_16020);
or U17792 (N_17792,N_16489,N_16618);
nor U17793 (N_17793,N_16675,N_16743);
nand U17794 (N_17794,N_16279,N_16280);
nor U17795 (N_17795,N_15618,N_16078);
and U17796 (N_17796,N_16477,N_16473);
xnor U17797 (N_17797,N_15727,N_15928);
and U17798 (N_17798,N_16407,N_16451);
or U17799 (N_17799,N_16509,N_16425);
nor U17800 (N_17800,N_16274,N_16419);
and U17801 (N_17801,N_15751,N_16651);
nor U17802 (N_17802,N_16232,N_16726);
and U17803 (N_17803,N_16358,N_16642);
nor U17804 (N_17804,N_16171,N_15910);
or U17805 (N_17805,N_15871,N_16065);
or U17806 (N_17806,N_16647,N_15765);
and U17807 (N_17807,N_16310,N_15692);
and U17808 (N_17808,N_16787,N_16715);
xnor U17809 (N_17809,N_15683,N_16322);
or U17810 (N_17810,N_16633,N_15816);
nand U17811 (N_17811,N_16559,N_15970);
and U17812 (N_17812,N_16256,N_15980);
nor U17813 (N_17813,N_15759,N_15680);
and U17814 (N_17814,N_16336,N_16030);
xor U17815 (N_17815,N_16728,N_15794);
and U17816 (N_17816,N_16330,N_16035);
or U17817 (N_17817,N_16478,N_16138);
nor U17818 (N_17818,N_16796,N_16404);
xnor U17819 (N_17819,N_16653,N_16028);
or U17820 (N_17820,N_16701,N_16024);
nor U17821 (N_17821,N_16036,N_16429);
and U17822 (N_17822,N_16391,N_15607);
or U17823 (N_17823,N_15907,N_15958);
xor U17824 (N_17824,N_16085,N_16003);
and U17825 (N_17825,N_15614,N_16139);
or U17826 (N_17826,N_16209,N_16530);
nand U17827 (N_17827,N_16287,N_15684);
nand U17828 (N_17828,N_16645,N_16522);
xor U17829 (N_17829,N_16698,N_16085);
xor U17830 (N_17830,N_16642,N_16025);
and U17831 (N_17831,N_16442,N_16552);
xor U17832 (N_17832,N_15877,N_15893);
xor U17833 (N_17833,N_16051,N_16782);
nand U17834 (N_17834,N_16081,N_16109);
and U17835 (N_17835,N_16513,N_16572);
nor U17836 (N_17836,N_16549,N_15691);
xnor U17837 (N_17837,N_15970,N_16206);
and U17838 (N_17838,N_15985,N_16782);
xnor U17839 (N_17839,N_15761,N_16604);
nor U17840 (N_17840,N_15805,N_15934);
and U17841 (N_17841,N_16615,N_15717);
nand U17842 (N_17842,N_15671,N_16041);
nor U17843 (N_17843,N_16681,N_16396);
xor U17844 (N_17844,N_16581,N_16454);
or U17845 (N_17845,N_16559,N_16122);
nand U17846 (N_17846,N_16155,N_16052);
and U17847 (N_17847,N_15996,N_16166);
nand U17848 (N_17848,N_15835,N_16079);
or U17849 (N_17849,N_15952,N_15990);
or U17850 (N_17850,N_16699,N_15836);
xor U17851 (N_17851,N_15865,N_16488);
nand U17852 (N_17852,N_16132,N_15684);
or U17853 (N_17853,N_15696,N_16212);
nand U17854 (N_17854,N_15728,N_15940);
xnor U17855 (N_17855,N_16272,N_16117);
and U17856 (N_17856,N_16171,N_16245);
and U17857 (N_17857,N_16219,N_16126);
xor U17858 (N_17858,N_15923,N_16205);
xnor U17859 (N_17859,N_15963,N_16453);
and U17860 (N_17860,N_16270,N_16568);
nand U17861 (N_17861,N_16436,N_16576);
xnor U17862 (N_17862,N_16579,N_15950);
nand U17863 (N_17863,N_16258,N_16093);
xnor U17864 (N_17864,N_15809,N_16079);
xor U17865 (N_17865,N_15899,N_16538);
xnor U17866 (N_17866,N_16616,N_16442);
xnor U17867 (N_17867,N_16155,N_16363);
or U17868 (N_17868,N_16767,N_15613);
xor U17869 (N_17869,N_15883,N_16239);
or U17870 (N_17870,N_16262,N_16645);
nor U17871 (N_17871,N_16452,N_15631);
or U17872 (N_17872,N_16093,N_16440);
nor U17873 (N_17873,N_15972,N_16062);
and U17874 (N_17874,N_16374,N_15650);
xor U17875 (N_17875,N_16029,N_16471);
nor U17876 (N_17876,N_16498,N_15840);
xor U17877 (N_17877,N_16399,N_15978);
xnor U17878 (N_17878,N_15952,N_15987);
or U17879 (N_17879,N_16654,N_15719);
and U17880 (N_17880,N_16525,N_16523);
xnor U17881 (N_17881,N_16538,N_15716);
nand U17882 (N_17882,N_16198,N_16286);
nor U17883 (N_17883,N_16299,N_16196);
xor U17884 (N_17884,N_15911,N_16443);
xor U17885 (N_17885,N_16352,N_16710);
or U17886 (N_17886,N_16721,N_16422);
nand U17887 (N_17887,N_15600,N_16226);
nand U17888 (N_17888,N_16547,N_16714);
and U17889 (N_17889,N_16273,N_15966);
and U17890 (N_17890,N_15933,N_16634);
and U17891 (N_17891,N_15696,N_15700);
xnor U17892 (N_17892,N_16291,N_16177);
nand U17893 (N_17893,N_16657,N_15720);
and U17894 (N_17894,N_16137,N_16120);
nor U17895 (N_17895,N_16461,N_15771);
nor U17896 (N_17896,N_15684,N_15863);
nor U17897 (N_17897,N_16279,N_16532);
xnor U17898 (N_17898,N_15668,N_16748);
nor U17899 (N_17899,N_16078,N_16367);
nor U17900 (N_17900,N_16769,N_15861);
and U17901 (N_17901,N_16791,N_16017);
or U17902 (N_17902,N_15883,N_16558);
xnor U17903 (N_17903,N_16010,N_16434);
nor U17904 (N_17904,N_16778,N_15842);
or U17905 (N_17905,N_16421,N_16530);
and U17906 (N_17906,N_15825,N_16237);
or U17907 (N_17907,N_16488,N_15741);
and U17908 (N_17908,N_16590,N_16023);
or U17909 (N_17909,N_16380,N_16791);
and U17910 (N_17910,N_15940,N_16260);
and U17911 (N_17911,N_16335,N_16024);
xor U17912 (N_17912,N_16103,N_16263);
and U17913 (N_17913,N_16069,N_15780);
xnor U17914 (N_17914,N_16123,N_16549);
xnor U17915 (N_17915,N_15764,N_16548);
nor U17916 (N_17916,N_16362,N_15632);
nand U17917 (N_17917,N_16392,N_16319);
nand U17918 (N_17918,N_16636,N_16538);
nand U17919 (N_17919,N_16628,N_16496);
nand U17920 (N_17920,N_15783,N_15864);
and U17921 (N_17921,N_16518,N_15720);
and U17922 (N_17922,N_16744,N_16374);
nor U17923 (N_17923,N_16781,N_16386);
nand U17924 (N_17924,N_15974,N_15882);
nor U17925 (N_17925,N_16538,N_15959);
or U17926 (N_17926,N_16578,N_16571);
xor U17927 (N_17927,N_16011,N_16049);
nor U17928 (N_17928,N_16759,N_16670);
and U17929 (N_17929,N_15750,N_15823);
and U17930 (N_17930,N_16749,N_16440);
or U17931 (N_17931,N_15737,N_15640);
or U17932 (N_17932,N_16447,N_16250);
nand U17933 (N_17933,N_16723,N_15918);
xnor U17934 (N_17934,N_15656,N_16169);
and U17935 (N_17935,N_15972,N_16096);
nor U17936 (N_17936,N_16616,N_16756);
nor U17937 (N_17937,N_16135,N_16175);
and U17938 (N_17938,N_16098,N_16218);
nand U17939 (N_17939,N_15735,N_15630);
nor U17940 (N_17940,N_16059,N_15897);
nor U17941 (N_17941,N_15721,N_15868);
xnor U17942 (N_17942,N_16729,N_16350);
or U17943 (N_17943,N_16555,N_16087);
nor U17944 (N_17944,N_15848,N_16606);
xor U17945 (N_17945,N_15819,N_16586);
nand U17946 (N_17946,N_16289,N_16135);
or U17947 (N_17947,N_15847,N_15889);
nand U17948 (N_17948,N_15896,N_16011);
and U17949 (N_17949,N_16098,N_16434);
or U17950 (N_17950,N_16433,N_15866);
and U17951 (N_17951,N_16289,N_16334);
and U17952 (N_17952,N_16179,N_16258);
or U17953 (N_17953,N_15792,N_15788);
xor U17954 (N_17954,N_16787,N_16611);
nor U17955 (N_17955,N_16541,N_16679);
and U17956 (N_17956,N_15975,N_16444);
nor U17957 (N_17957,N_16239,N_16786);
xnor U17958 (N_17958,N_15828,N_15857);
xnor U17959 (N_17959,N_16687,N_16127);
or U17960 (N_17960,N_16400,N_15810);
nand U17961 (N_17961,N_15696,N_16665);
and U17962 (N_17962,N_16005,N_16267);
nand U17963 (N_17963,N_15724,N_16500);
and U17964 (N_17964,N_16132,N_16794);
and U17965 (N_17965,N_16647,N_15673);
and U17966 (N_17966,N_16130,N_15932);
and U17967 (N_17967,N_15823,N_16581);
and U17968 (N_17968,N_16278,N_15814);
or U17969 (N_17969,N_15949,N_16374);
nand U17970 (N_17970,N_16713,N_15711);
or U17971 (N_17971,N_15675,N_16699);
or U17972 (N_17972,N_16682,N_16372);
and U17973 (N_17973,N_16472,N_15746);
nor U17974 (N_17974,N_16263,N_16528);
nand U17975 (N_17975,N_16380,N_16004);
nor U17976 (N_17976,N_16661,N_16523);
or U17977 (N_17977,N_15957,N_15655);
and U17978 (N_17978,N_15617,N_16714);
or U17979 (N_17979,N_16654,N_15785);
and U17980 (N_17980,N_16000,N_15909);
xor U17981 (N_17981,N_16681,N_16608);
and U17982 (N_17982,N_16044,N_16430);
nor U17983 (N_17983,N_16633,N_16726);
nand U17984 (N_17984,N_16586,N_16269);
xor U17985 (N_17985,N_15706,N_16316);
nor U17986 (N_17986,N_16546,N_16221);
nor U17987 (N_17987,N_16439,N_16293);
nand U17988 (N_17988,N_16388,N_16518);
or U17989 (N_17989,N_15718,N_16180);
nand U17990 (N_17990,N_16247,N_15900);
nand U17991 (N_17991,N_16727,N_16665);
xor U17992 (N_17992,N_16220,N_16168);
nor U17993 (N_17993,N_15611,N_16411);
and U17994 (N_17994,N_16017,N_16295);
nand U17995 (N_17995,N_16331,N_16477);
nor U17996 (N_17996,N_16053,N_16364);
xnor U17997 (N_17997,N_16772,N_15826);
nand U17998 (N_17998,N_15759,N_16065);
or U17999 (N_17999,N_16422,N_16286);
and U18000 (N_18000,N_17052,N_17902);
nor U18001 (N_18001,N_17203,N_17268);
xor U18002 (N_18002,N_16826,N_17973);
nor U18003 (N_18003,N_17633,N_17719);
xor U18004 (N_18004,N_17798,N_17486);
and U18005 (N_18005,N_17690,N_17082);
nor U18006 (N_18006,N_16912,N_17684);
or U18007 (N_18007,N_17861,N_17614);
nand U18008 (N_18008,N_16831,N_16889);
nor U18009 (N_18009,N_17780,N_17514);
or U18010 (N_18010,N_17980,N_17771);
and U18011 (N_18011,N_17083,N_17863);
and U18012 (N_18012,N_17033,N_17160);
nand U18013 (N_18013,N_17939,N_16983);
nand U18014 (N_18014,N_17652,N_17742);
xnor U18015 (N_18015,N_17169,N_16813);
xnor U18016 (N_18016,N_17774,N_17316);
nand U18017 (N_18017,N_17458,N_17537);
and U18018 (N_18018,N_17376,N_17923);
nor U18019 (N_18019,N_17872,N_17635);
or U18020 (N_18020,N_17870,N_16802);
nand U18021 (N_18021,N_17163,N_17740);
nand U18022 (N_18022,N_17747,N_17851);
nor U18023 (N_18023,N_16943,N_17200);
xnor U18024 (N_18024,N_17871,N_17366);
or U18025 (N_18025,N_17425,N_17415);
and U18026 (N_18026,N_17062,N_17648);
and U18027 (N_18027,N_17734,N_16921);
nand U18028 (N_18028,N_17258,N_17249);
xor U18029 (N_18029,N_17176,N_17718);
nand U18030 (N_18030,N_17839,N_17960);
nand U18031 (N_18031,N_17977,N_17264);
xnor U18032 (N_18032,N_17476,N_17009);
or U18033 (N_18033,N_17398,N_17876);
nand U18034 (N_18034,N_17976,N_17820);
nand U18035 (N_18035,N_17613,N_17595);
and U18036 (N_18036,N_17515,N_17253);
or U18037 (N_18037,N_17324,N_17859);
xor U18038 (N_18038,N_17528,N_17015);
and U18039 (N_18039,N_17619,N_17251);
and U18040 (N_18040,N_17165,N_17498);
xor U18041 (N_18041,N_17322,N_17461);
xor U18042 (N_18042,N_17447,N_17215);
or U18043 (N_18043,N_17523,N_16890);
and U18044 (N_18044,N_16982,N_17815);
and U18045 (N_18045,N_17315,N_17529);
and U18046 (N_18046,N_17847,N_17267);
and U18047 (N_18047,N_16884,N_17683);
or U18048 (N_18048,N_17762,N_17812);
xor U18049 (N_18049,N_17763,N_17544);
xnor U18050 (N_18050,N_17339,N_17494);
xnor U18051 (N_18051,N_17412,N_17705);
or U18052 (N_18052,N_17834,N_17618);
nor U18053 (N_18053,N_17724,N_17021);
xor U18054 (N_18054,N_17752,N_17416);
nor U18055 (N_18055,N_17707,N_17354);
or U18056 (N_18056,N_16855,N_17346);
nand U18057 (N_18057,N_17569,N_17842);
xnor U18058 (N_18058,N_17521,N_17301);
and U18059 (N_18059,N_17908,N_17749);
xor U18060 (N_18060,N_16990,N_17290);
xnor U18061 (N_18061,N_17916,N_17556);
and U18062 (N_18062,N_17188,N_17917);
or U18063 (N_18063,N_16951,N_17548);
nand U18064 (N_18064,N_17000,N_17985);
xnor U18065 (N_18065,N_16887,N_17883);
and U18066 (N_18066,N_16876,N_17199);
nor U18067 (N_18067,N_17138,N_17185);
nor U18068 (N_18068,N_17887,N_17371);
or U18069 (N_18069,N_17961,N_17038);
xnor U18070 (N_18070,N_17472,N_17586);
nand U18071 (N_18071,N_17091,N_17475);
nand U18072 (N_18072,N_17443,N_17426);
nand U18073 (N_18073,N_17095,N_17533);
or U18074 (N_18074,N_17775,N_16851);
and U18075 (N_18075,N_17671,N_16965);
nor U18076 (N_18076,N_17123,N_17404);
nor U18077 (N_18077,N_17993,N_17010);
nor U18078 (N_18078,N_17103,N_17596);
and U18079 (N_18079,N_17470,N_17209);
xor U18080 (N_18080,N_17625,N_17406);
xnor U18081 (N_18081,N_17144,N_17356);
nor U18082 (N_18082,N_17282,N_16918);
and U18083 (N_18083,N_17706,N_17841);
or U18084 (N_18084,N_17727,N_17177);
nor U18085 (N_18085,N_17609,N_17604);
or U18086 (N_18086,N_17431,N_17304);
nor U18087 (N_18087,N_16994,N_17658);
and U18088 (N_18088,N_16872,N_17807);
xnor U18089 (N_18089,N_17418,N_17410);
and U18090 (N_18090,N_17168,N_17195);
xnor U18091 (N_18091,N_17142,N_16961);
or U18092 (N_18092,N_17938,N_16938);
nor U18093 (N_18093,N_17270,N_16853);
xor U18094 (N_18094,N_17137,N_17906);
xor U18095 (N_18095,N_17636,N_17140);
and U18096 (N_18096,N_16863,N_17161);
or U18097 (N_18097,N_17744,N_17483);
nor U18098 (N_18098,N_17532,N_17988);
nor U18099 (N_18099,N_17827,N_17293);
or U18100 (N_18100,N_17881,N_16870);
or U18101 (N_18101,N_17034,N_16922);
xnor U18102 (N_18102,N_16968,N_17351);
nand U18103 (N_18103,N_17682,N_17286);
nor U18104 (N_18104,N_17440,N_17929);
and U18105 (N_18105,N_17184,N_17835);
or U18106 (N_18106,N_17904,N_17287);
and U18107 (N_18107,N_17480,N_17983);
or U18108 (N_18108,N_17358,N_17954);
or U18109 (N_18109,N_17273,N_17477);
xnor U18110 (N_18110,N_17232,N_17832);
and U18111 (N_18111,N_17814,N_17893);
and U18112 (N_18112,N_17868,N_16899);
and U18113 (N_18113,N_17387,N_17784);
nor U18114 (N_18114,N_17029,N_17673);
or U18115 (N_18115,N_17074,N_17712);
or U18116 (N_18116,N_17298,N_17219);
nand U18117 (N_18117,N_16935,N_17332);
nor U18118 (N_18118,N_17539,N_17182);
nand U18119 (N_18119,N_17550,N_17720);
xnor U18120 (N_18120,N_17114,N_17023);
nand U18121 (N_18121,N_16842,N_16984);
or U18122 (N_18122,N_17221,N_17765);
nor U18123 (N_18123,N_17922,N_17989);
and U18124 (N_18124,N_16864,N_17849);
nor U18125 (N_18125,N_17069,N_17901);
nand U18126 (N_18126,N_17124,N_17650);
nand U18127 (N_18127,N_17030,N_17357);
nor U18128 (N_18128,N_17723,N_17998);
and U18129 (N_18129,N_16907,N_17466);
nor U18130 (N_18130,N_17921,N_17198);
nor U18131 (N_18131,N_17288,N_17846);
and U18132 (N_18132,N_17259,N_17111);
xor U18133 (N_18133,N_17255,N_17878);
nor U18134 (N_18134,N_16931,N_17601);
or U18135 (N_18135,N_17855,N_17150);
nor U18136 (N_18136,N_17152,N_17996);
and U18137 (N_18137,N_17552,N_17745);
nand U18138 (N_18138,N_17924,N_16875);
nand U18139 (N_18139,N_16999,N_16911);
and U18140 (N_18140,N_17218,N_17369);
nor U18141 (N_18141,N_17585,N_17553);
and U18142 (N_18142,N_17167,N_17858);
and U18143 (N_18143,N_16959,N_17299);
or U18144 (N_18144,N_17736,N_17520);
xnor U18145 (N_18145,N_17640,N_17795);
or U18146 (N_18146,N_16878,N_17309);
xor U18147 (N_18147,N_17330,N_17790);
nor U18148 (N_18148,N_16972,N_17700);
and U18149 (N_18149,N_17244,N_16824);
nor U18150 (N_18150,N_17231,N_16850);
nand U18151 (N_18151,N_17056,N_17670);
and U18152 (N_18152,N_17321,N_17016);
xor U18153 (N_18153,N_17263,N_17992);
nor U18154 (N_18154,N_17860,N_17078);
and U18155 (N_18155,N_16955,N_17968);
xnor U18156 (N_18156,N_16900,N_17323);
and U18157 (N_18157,N_17930,N_17757);
and U18158 (N_18158,N_16975,N_17493);
nor U18159 (N_18159,N_17452,N_17420);
nand U18160 (N_18160,N_17344,N_17879);
or U18161 (N_18161,N_16954,N_17910);
nand U18162 (N_18162,N_17730,N_17469);
and U18163 (N_18163,N_17037,N_16926);
and U18164 (N_18164,N_17385,N_17606);
xnor U18165 (N_18165,N_17106,N_16814);
xor U18166 (N_18166,N_16810,N_17283);
xnor U18167 (N_18167,N_17829,N_17157);
nand U18168 (N_18168,N_17984,N_17822);
and U18169 (N_18169,N_17627,N_16945);
or U18170 (N_18170,N_16881,N_17068);
and U18171 (N_18171,N_17838,N_17400);
and U18172 (N_18172,N_17485,N_16962);
and U18173 (N_18173,N_17554,N_17001);
and U18174 (N_18174,N_17972,N_17665);
or U18175 (N_18175,N_17672,N_16976);
and U18176 (N_18176,N_17402,N_17396);
or U18177 (N_18177,N_17125,N_17383);
or U18178 (N_18178,N_17927,N_17252);
xnor U18179 (N_18179,N_17239,N_17227);
nand U18180 (N_18180,N_17122,N_17438);
xnor U18181 (N_18181,N_17139,N_17307);
xnor U18182 (N_18182,N_16829,N_16997);
or U18183 (N_18183,N_16981,N_17563);
or U18184 (N_18184,N_17126,N_17173);
or U18185 (N_18185,N_17560,N_17629);
nor U18186 (N_18186,N_17667,N_17269);
and U18187 (N_18187,N_17555,N_17053);
nand U18188 (N_18188,N_16904,N_17940);
nand U18189 (N_18189,N_17660,N_17534);
or U18190 (N_18190,N_17495,N_17326);
xnor U18191 (N_18191,N_17217,N_16821);
or U18192 (N_18192,N_17701,N_17492);
xor U18193 (N_18193,N_17329,N_16839);
nand U18194 (N_18194,N_17561,N_16923);
xor U18195 (N_18195,N_17733,N_16948);
xor U18196 (N_18196,N_16992,N_17689);
xor U18197 (N_18197,N_17786,N_16800);
nand U18198 (N_18198,N_16919,N_16995);
nand U18199 (N_18199,N_17424,N_17147);
or U18200 (N_18200,N_17362,N_17957);
and U18201 (N_18201,N_16828,N_16905);
or U18202 (N_18202,N_16822,N_17454);
nand U18203 (N_18203,N_17955,N_17007);
and U18204 (N_18204,N_17739,N_17926);
xor U18205 (N_18205,N_17436,N_16836);
nand U18206 (N_18206,N_17496,N_17190);
nor U18207 (N_18207,N_16966,N_17228);
nand U18208 (N_18208,N_16940,N_17025);
nor U18209 (N_18209,N_17119,N_16862);
or U18210 (N_18210,N_16957,N_17570);
and U18211 (N_18211,N_16874,N_17313);
nor U18212 (N_18212,N_17112,N_17393);
and U18213 (N_18213,N_17800,N_17422);
nor U18214 (N_18214,N_17072,N_17035);
xor U18215 (N_18215,N_17811,N_17071);
and U18216 (N_18216,N_17265,N_17368);
and U18217 (N_18217,N_17004,N_17519);
xnor U18218 (N_18218,N_16952,N_17272);
or U18219 (N_18219,N_17699,N_17610);
nor U18220 (N_18220,N_17349,N_17711);
and U18221 (N_18221,N_17801,N_17238);
nor U18222 (N_18222,N_17233,N_17732);
nor U18223 (N_18223,N_17319,N_17064);
nand U18224 (N_18224,N_17802,N_17120);
nand U18225 (N_18225,N_17628,N_17389);
xnor U18226 (N_18226,N_17918,N_17174);
nor U18227 (N_18227,N_16902,N_16989);
and U18228 (N_18228,N_16861,N_17380);
and U18229 (N_18229,N_17503,N_17830);
nand U18230 (N_18230,N_17070,N_17128);
nand U18231 (N_18231,N_17455,N_17220);
or U18232 (N_18232,N_17194,N_17085);
nor U18233 (N_18233,N_17278,N_17943);
xnor U18234 (N_18234,N_16933,N_17409);
nand U18235 (N_18235,N_17237,N_16838);
nand U18236 (N_18236,N_16979,N_17819);
xnor U18237 (N_18237,N_17865,N_16819);
nand U18238 (N_18238,N_17753,N_17783);
nor U18239 (N_18239,N_17439,N_17243);
xor U18240 (N_18240,N_17340,N_16941);
and U18241 (N_18241,N_17006,N_17271);
xnor U18242 (N_18242,N_17372,N_17407);
nor U18243 (N_18243,N_17912,N_17364);
nand U18244 (N_18244,N_16844,N_17262);
xnor U18245 (N_18245,N_17118,N_17970);
or U18246 (N_18246,N_17365,N_17240);
nand U18247 (N_18247,N_17427,N_17448);
xor U18248 (N_18248,N_17662,N_17698);
nor U18249 (N_18249,N_17964,N_17593);
or U18250 (N_18250,N_17442,N_16882);
and U18251 (N_18251,N_17444,N_17709);
nor U18252 (N_18252,N_17417,N_16883);
nand U18253 (N_18253,N_17113,N_17017);
nand U18254 (N_18254,N_17688,N_17681);
xnor U18255 (N_18255,N_17058,N_17279);
and U18256 (N_18256,N_17430,N_17236);
and U18257 (N_18257,N_17411,N_17840);
or U18258 (N_18258,N_17451,N_17668);
xnor U18259 (N_18259,N_17211,N_17919);
and U18260 (N_18260,N_17674,N_17159);
or U18261 (N_18261,N_17145,N_17620);
nand U18262 (N_18262,N_16987,N_17951);
or U18263 (N_18263,N_17837,N_16841);
nor U18264 (N_18264,N_16924,N_17192);
xor U18265 (N_18265,N_16950,N_17027);
nor U18266 (N_18266,N_17026,N_17543);
and U18267 (N_18267,N_17931,N_17474);
and U18268 (N_18268,N_17615,N_17403);
and U18269 (N_18269,N_16980,N_17894);
xor U18270 (N_18270,N_17591,N_17327);
xnor U18271 (N_18271,N_17116,N_17805);
nand U18272 (N_18272,N_17969,N_17468);
xor U18273 (N_18273,N_16996,N_16986);
xor U18274 (N_18274,N_17647,N_17012);
and U18275 (N_18275,N_17680,N_17501);
xor U18276 (N_18276,N_17051,N_16973);
xnor U18277 (N_18277,N_17275,N_17981);
nand U18278 (N_18278,N_17731,N_17024);
nor U18279 (N_18279,N_16934,N_16910);
nand U18280 (N_18280,N_17579,N_17391);
nor U18281 (N_18281,N_17696,N_17948);
nand U18282 (N_18282,N_17577,N_16937);
or U18283 (N_18283,N_17877,N_17979);
nor U18284 (N_18284,N_17453,N_17959);
xor U18285 (N_18285,N_17080,N_17077);
xnor U18286 (N_18286,N_16960,N_17562);
and U18287 (N_18287,N_17090,N_16942);
or U18288 (N_18288,N_16978,N_17445);
nand U18289 (N_18289,N_17675,N_17994);
xnor U18290 (N_18290,N_17896,N_17942);
nor U18291 (N_18291,N_17484,N_17588);
or U18292 (N_18292,N_17646,N_17589);
or U18293 (N_18293,N_17768,N_16837);
or U18294 (N_18294,N_16913,N_17225);
and U18295 (N_18295,N_17508,N_17792);
nand U18296 (N_18296,N_17638,N_16928);
nand U18297 (N_18297,N_17512,N_17121);
or U18298 (N_18298,N_17055,N_17760);
nand U18299 (N_18299,N_17644,N_17204);
nand U18300 (N_18300,N_17289,N_17280);
xnor U18301 (N_18301,N_16991,N_17401);
or U18302 (N_18302,N_17828,N_17623);
nand U18303 (N_18303,N_17018,N_16880);
or U18304 (N_18304,N_17808,N_17716);
nand U18305 (N_18305,N_17833,N_17797);
nand U18306 (N_18306,N_17207,N_17076);
xnor U18307 (N_18307,N_16929,N_17156);
nor U18308 (N_18308,N_17617,N_17110);
or U18309 (N_18309,N_17907,N_17518);
nand U18310 (N_18310,N_17886,N_17054);
xor U18311 (N_18311,N_17748,N_16915);
or U18312 (N_18312,N_17459,N_17936);
nand U18313 (N_18313,N_17148,N_17285);
xnor U18314 (N_18314,N_17934,N_16885);
and U18315 (N_18315,N_17962,N_17245);
xor U18316 (N_18316,N_17965,N_16858);
or U18317 (N_18317,N_16847,N_17506);
xor U18318 (N_18318,N_17261,N_17210);
nand U18319 (N_18319,N_17005,N_17094);
xnor U18320 (N_18320,N_17639,N_17889);
nor U18321 (N_18321,N_17626,N_17041);
nand U18322 (N_18322,N_17487,N_16871);
or U18323 (N_18323,N_17178,N_17414);
nor U18324 (N_18324,N_16804,N_17097);
and U18325 (N_18325,N_16891,N_16849);
xor U18326 (N_18326,N_17325,N_17890);
nor U18327 (N_18327,N_17153,N_17158);
nand U18328 (N_18328,N_17810,N_17900);
nand U18329 (N_18329,N_17587,N_17999);
and U18330 (N_18330,N_17713,N_16843);
nor U18331 (N_18331,N_17741,N_16888);
xor U18332 (N_18332,N_16820,N_17641);
xnor U18333 (N_18333,N_16816,N_17063);
nor U18334 (N_18334,N_17777,N_17995);
or U18335 (N_18335,N_17465,N_17963);
nor U18336 (N_18336,N_16877,N_17405);
nand U18337 (N_18337,N_17205,N_16927);
nand U18338 (N_18338,N_16845,N_17036);
and U18339 (N_18339,N_17428,N_16856);
nand U18340 (N_18340,N_17758,N_17637);
nor U18341 (N_18341,N_17598,N_17818);
nor U18342 (N_18342,N_17394,N_17502);
and U18343 (N_18343,N_17086,N_17597);
nand U18344 (N_18344,N_17093,N_16998);
xor U18345 (N_18345,N_17216,N_17920);
nor U18346 (N_18346,N_17578,N_17778);
nand U18347 (N_18347,N_17911,N_17341);
nand U18348 (N_18348,N_17104,N_17717);
xor U18349 (N_18349,N_17621,N_17379);
or U18350 (N_18350,N_17363,N_17605);
and U18351 (N_18351,N_17117,N_17296);
nand U18352 (N_18352,N_16906,N_17949);
xnor U18353 (N_18353,N_17971,N_17175);
nand U18354 (N_18354,N_17183,N_17915);
or U18355 (N_18355,N_17928,N_17726);
nand U18356 (N_18356,N_17429,N_17488);
xnor U18357 (N_18357,N_16917,N_17862);
xor U18358 (N_18358,N_17320,N_17541);
xnor U18359 (N_18359,N_17791,N_16857);
nor U18360 (N_18360,N_17135,N_17276);
xnor U18361 (N_18361,N_17694,N_17974);
or U18362 (N_18362,N_17105,N_17504);
or U18363 (N_18363,N_17347,N_17663);
xnor U18364 (N_18364,N_17715,N_17317);
and U18365 (N_18365,N_17845,N_17946);
or U18366 (N_18366,N_17743,N_17446);
nor U18367 (N_18367,N_17399,N_16925);
or U18368 (N_18368,N_17599,N_17134);
nand U18369 (N_18369,N_17982,N_17678);
or U18370 (N_18370,N_17754,N_16949);
nor U18371 (N_18371,N_17222,N_17008);
or U18372 (N_18372,N_17978,N_17722);
nand U18373 (N_18373,N_17456,N_17359);
or U18374 (N_18374,N_17513,N_16914);
nor U18375 (N_18375,N_17292,N_17067);
or U18376 (N_18376,N_17108,N_17566);
nand U18377 (N_18377,N_17099,N_17014);
xor U18378 (N_18378,N_17704,N_16835);
or U18379 (N_18379,N_17821,N_17735);
xnor U18380 (N_18380,N_17857,N_17728);
nor U18381 (N_18381,N_17129,N_16834);
and U18382 (N_18382,N_17952,N_16825);
xor U18383 (N_18383,N_17869,N_17300);
nand U18384 (N_18384,N_17558,N_16809);
xnor U18385 (N_18385,N_17079,N_17306);
xnor U18386 (N_18386,N_17831,N_17434);
or U18387 (N_18387,N_17527,N_17181);
xnor U18388 (N_18388,N_16896,N_16854);
nor U18389 (N_18389,N_17019,N_17944);
and U18390 (N_18390,N_16958,N_17266);
and U18391 (N_18391,N_17098,N_17043);
nand U18392 (N_18392,N_17193,N_17274);
nor U18393 (N_18393,N_17549,N_17729);
xor U18394 (N_18394,N_17305,N_17464);
or U18395 (N_18395,N_17028,N_17151);
nand U18396 (N_18396,N_17499,N_17524);
or U18397 (N_18397,N_17224,N_16893);
or U18398 (N_18398,N_16969,N_17676);
xor U18399 (N_18399,N_17413,N_17785);
or U18400 (N_18400,N_17953,N_17651);
and U18401 (N_18401,N_17467,N_17213);
nand U18402 (N_18402,N_17809,N_16967);
nor U18403 (N_18403,N_16956,N_17941);
or U18404 (N_18404,N_17866,N_17350);
and U18405 (N_18405,N_16868,N_17049);
nor U18406 (N_18406,N_17109,N_17505);
xor U18407 (N_18407,N_17950,N_17816);
nor U18408 (N_18408,N_17208,N_17759);
nand U18409 (N_18409,N_17914,N_17769);
nor U18410 (N_18410,N_17656,N_16970);
nand U18411 (N_18411,N_17526,N_17423);
xor U18412 (N_18412,N_17891,N_17721);
or U18413 (N_18413,N_17612,N_17884);
xnor U18414 (N_18414,N_16846,N_16860);
nand U18415 (N_18415,N_17202,N_17382);
xnor U18416 (N_18416,N_17449,N_16898);
xnor U18417 (N_18417,N_17378,N_17066);
nor U18418 (N_18418,N_16964,N_17525);
or U18419 (N_18419,N_17260,N_17880);
xor U18420 (N_18420,N_17582,N_17281);
and U18421 (N_18421,N_17065,N_17302);
nor U18422 (N_18422,N_17856,N_17328);
nor U18423 (N_18423,N_17115,N_17888);
nor U18424 (N_18424,N_17482,N_17473);
xnor U18425 (N_18425,N_17565,N_17530);
or U18426 (N_18426,N_16897,N_17042);
or U18427 (N_18427,N_17654,N_17574);
nor U18428 (N_18428,N_17966,N_17229);
nor U18429 (N_18429,N_17048,N_17642);
and U18430 (N_18430,N_17360,N_17779);
nor U18431 (N_18431,N_17746,N_17864);
nor U18432 (N_18432,N_17295,N_17457);
or U18433 (N_18433,N_17710,N_17045);
nor U18434 (N_18434,N_16985,N_17975);
nor U18435 (N_18435,N_16953,N_17516);
nor U18436 (N_18436,N_16805,N_17803);
xor U18437 (N_18437,N_17102,N_17510);
xnor U18438 (N_18438,N_16873,N_16879);
and U18439 (N_18439,N_17162,N_17107);
xnor U18440 (N_18440,N_17352,N_17047);
nand U18441 (N_18441,N_16974,N_17538);
nor U18442 (N_18442,N_17463,N_17419);
or U18443 (N_18443,N_17789,N_17767);
nand U18444 (N_18444,N_17248,N_17899);
nor U18445 (N_18445,N_17377,N_17630);
and U18446 (N_18446,N_17491,N_17435);
xor U18447 (N_18447,N_16892,N_16848);
nor U18448 (N_18448,N_17214,N_17146);
and U18449 (N_18449,N_17310,N_16811);
or U18450 (N_18450,N_16852,N_17003);
nand U18451 (N_18451,N_17693,N_17686);
and U18452 (N_18452,N_17772,N_17172);
nor U18453 (N_18453,N_17885,N_17294);
xor U18454 (N_18454,N_17817,N_17632);
nand U18455 (N_18455,N_17397,N_17154);
nand U18456 (N_18456,N_17559,N_17594);
or U18457 (N_18457,N_17571,N_17254);
xor U18458 (N_18458,N_17206,N_17450);
nand U18459 (N_18459,N_17046,N_17853);
xnor U18460 (N_18460,N_17823,N_17836);
nand U18461 (N_18461,N_17040,N_17246);
and U18462 (N_18462,N_17787,N_17002);
or U18463 (N_18463,N_17471,N_17657);
nor U18464 (N_18464,N_17337,N_17186);
or U18465 (N_18465,N_17522,N_17773);
nor U18466 (N_18466,N_17250,N_17164);
nand U18467 (N_18467,N_17958,N_17584);
nor U18468 (N_18468,N_17875,N_17575);
nor U18469 (N_18469,N_17611,N_17750);
nor U18470 (N_18470,N_16895,N_17564);
or U18471 (N_18471,N_17603,N_17130);
nor U18472 (N_18472,N_17655,N_17854);
nor U18473 (N_18473,N_17687,N_17607);
nor U18474 (N_18474,N_16867,N_17898);
nor U18475 (N_18475,N_17334,N_17551);
or U18476 (N_18476,N_17697,N_17702);
or U18477 (N_18477,N_17945,N_17087);
or U18478 (N_18478,N_17247,N_17421);
nor U18479 (N_18479,N_16977,N_17256);
nand U18480 (N_18480,N_17634,N_17196);
nand U18481 (N_18481,N_17441,N_17373);
nand U18482 (N_18482,N_17133,N_17489);
nand U18483 (N_18483,N_17677,N_17545);
nor U18484 (N_18484,N_17355,N_17991);
or U18485 (N_18485,N_17437,N_16830);
and U18486 (N_18486,N_16807,N_16808);
or U18487 (N_18487,N_17013,N_17131);
xnor U18488 (N_18488,N_17084,N_17061);
and U18489 (N_18489,N_17297,N_17235);
nor U18490 (N_18490,N_17990,N_17039);
nor U18491 (N_18491,N_17166,N_17947);
nor U18492 (N_18492,N_17191,N_16866);
xor U18493 (N_18493,N_16946,N_17500);
nor U18494 (N_18494,N_17799,N_17059);
xor U18495 (N_18495,N_17873,N_17781);
nand U18496 (N_18496,N_17653,N_17725);
nor U18497 (N_18497,N_17141,N_17882);
nor U18498 (N_18498,N_17011,N_17764);
or U18499 (N_18499,N_17590,N_16832);
nor U18500 (N_18500,N_17685,N_17649);
and U18501 (N_18501,N_17874,N_17987);
or U18502 (N_18502,N_17179,N_17170);
nand U18503 (N_18503,N_17032,N_17291);
nor U18504 (N_18504,N_17659,N_17348);
nand U18505 (N_18505,N_16936,N_17092);
nand U18506 (N_18506,N_17737,N_17101);
nor U18507 (N_18507,N_17751,N_17096);
xnor U18508 (N_18508,N_17234,N_17223);
xor U18509 (N_18509,N_17331,N_17661);
nand U18510 (N_18510,N_16930,N_17284);
xor U18511 (N_18511,N_17242,N_17189);
or U18512 (N_18512,N_17536,N_16840);
xnor U18513 (N_18513,N_16817,N_16963);
or U18514 (N_18514,N_17390,N_17738);
or U18515 (N_18515,N_17517,N_17692);
nand U18516 (N_18516,N_17695,N_17031);
nand U18517 (N_18517,N_16801,N_17903);
and U18518 (N_18518,N_17967,N_17583);
nor U18519 (N_18519,N_17187,N_17540);
and U18520 (N_18520,N_17666,N_17277);
or U18521 (N_18521,N_17643,N_17714);
xor U18522 (N_18522,N_17075,N_17535);
xor U18523 (N_18523,N_17844,N_17497);
or U18524 (N_18524,N_17825,N_17308);
xor U18525 (N_18525,N_16827,N_17892);
nor U18526 (N_18526,N_17804,N_17608);
and U18527 (N_18527,N_17333,N_17703);
xor U18528 (N_18528,N_16803,N_17462);
nand U18529 (N_18529,N_17057,N_17171);
and U18530 (N_18530,N_16939,N_17073);
nand U18531 (N_18531,N_17622,N_17576);
nand U18532 (N_18532,N_17794,N_17766);
xor U18533 (N_18533,N_17132,N_17572);
and U18534 (N_18534,N_17370,N_17852);
nor U18535 (N_18535,N_17511,N_17088);
and U18536 (N_18536,N_17581,N_17312);
nor U18537 (N_18537,N_17843,N_16894);
or U18538 (N_18538,N_16833,N_17303);
nor U18539 (N_18539,N_17933,N_17782);
and U18540 (N_18540,N_17460,N_17761);
and U18541 (N_18541,N_17212,N_17592);
or U18542 (N_18542,N_17568,N_17616);
nor U18543 (N_18543,N_17897,N_17342);
and U18544 (N_18544,N_16947,N_17909);
and U18545 (N_18545,N_17600,N_17509);
xor U18546 (N_18546,N_17756,N_17478);
nor U18547 (N_18547,N_17127,N_16909);
or U18548 (N_18548,N_17180,N_17230);
xnor U18549 (N_18549,N_17826,N_16865);
and U18550 (N_18550,N_17573,N_16901);
and U18551 (N_18551,N_17567,N_17314);
and U18552 (N_18552,N_17089,N_16818);
or U18553 (N_18553,N_17679,N_17793);
xnor U18554 (N_18554,N_16988,N_17956);
and U18555 (N_18555,N_17507,N_17813);
nor U18556 (N_18556,N_17155,N_17669);
xnor U18557 (N_18557,N_16971,N_17050);
and U18558 (N_18558,N_17776,N_17691);
xor U18559 (N_18559,N_17986,N_17353);
nor U18560 (N_18560,N_16944,N_17631);
and U18561 (N_18561,N_17481,N_17136);
xnor U18562 (N_18562,N_17770,N_17143);
xor U18563 (N_18563,N_17081,N_17020);
or U18564 (N_18564,N_17645,N_16869);
nand U18565 (N_18565,N_17624,N_17335);
and U18566 (N_18566,N_17343,N_17531);
nand U18567 (N_18567,N_17580,N_16932);
xor U18568 (N_18568,N_17937,N_17338);
or U18569 (N_18569,N_17345,N_17044);
xor U18570 (N_18570,N_16903,N_17408);
xor U18571 (N_18571,N_17336,N_17433);
or U18572 (N_18572,N_16908,N_17388);
or U18573 (N_18573,N_16859,N_17381);
xnor U18574 (N_18574,N_17395,N_17318);
nand U18575 (N_18575,N_17547,N_17060);
nor U18576 (N_18576,N_17788,N_17602);
xnor U18577 (N_18577,N_17490,N_17546);
and U18578 (N_18578,N_17100,N_16815);
and U18579 (N_18579,N_17557,N_17374);
nand U18580 (N_18580,N_17708,N_17542);
or U18581 (N_18581,N_17241,N_17913);
and U18582 (N_18582,N_17895,N_16806);
or U18583 (N_18583,N_17848,N_17997);
nor U18584 (N_18584,N_16993,N_17479);
nor U18585 (N_18585,N_16886,N_17022);
or U18586 (N_18586,N_16812,N_17755);
xor U18587 (N_18587,N_17905,N_17149);
or U18588 (N_18588,N_17384,N_17806);
xor U18589 (N_18589,N_17257,N_17850);
nor U18590 (N_18590,N_16920,N_17311);
nand U18591 (N_18591,N_17935,N_17796);
xor U18592 (N_18592,N_17361,N_17932);
or U18593 (N_18593,N_16823,N_17367);
xnor U18594 (N_18594,N_17201,N_17226);
xnor U18595 (N_18595,N_17824,N_17432);
xnor U18596 (N_18596,N_17867,N_17664);
nand U18597 (N_18597,N_17386,N_17392);
nand U18598 (N_18598,N_16916,N_17375);
nand U18599 (N_18599,N_17925,N_17197);
xnor U18600 (N_18600,N_17315,N_17989);
and U18601 (N_18601,N_17046,N_17160);
or U18602 (N_18602,N_17211,N_17175);
nand U18603 (N_18603,N_17393,N_17763);
and U18604 (N_18604,N_17067,N_17529);
or U18605 (N_18605,N_17784,N_17994);
nor U18606 (N_18606,N_16842,N_17377);
nand U18607 (N_18607,N_17369,N_17138);
nand U18608 (N_18608,N_17612,N_16953);
or U18609 (N_18609,N_17836,N_17630);
or U18610 (N_18610,N_16982,N_17126);
and U18611 (N_18611,N_17945,N_17289);
nor U18612 (N_18612,N_17507,N_17207);
or U18613 (N_18613,N_17441,N_17528);
xor U18614 (N_18614,N_17201,N_17878);
and U18615 (N_18615,N_17964,N_17161);
nand U18616 (N_18616,N_17386,N_17468);
and U18617 (N_18617,N_17693,N_16800);
nor U18618 (N_18618,N_17759,N_17951);
nand U18619 (N_18619,N_17821,N_17653);
xnor U18620 (N_18620,N_17178,N_17183);
nand U18621 (N_18621,N_17831,N_17758);
or U18622 (N_18622,N_17605,N_17531);
xor U18623 (N_18623,N_16989,N_17749);
xor U18624 (N_18624,N_17911,N_16902);
and U18625 (N_18625,N_16861,N_16874);
and U18626 (N_18626,N_16820,N_17972);
or U18627 (N_18627,N_17087,N_17450);
nand U18628 (N_18628,N_17613,N_17253);
or U18629 (N_18629,N_17169,N_17101);
nand U18630 (N_18630,N_17355,N_17319);
nand U18631 (N_18631,N_16990,N_17868);
xor U18632 (N_18632,N_17964,N_17134);
nand U18633 (N_18633,N_17475,N_17669);
nand U18634 (N_18634,N_17068,N_16899);
xor U18635 (N_18635,N_16837,N_17558);
xor U18636 (N_18636,N_17327,N_17366);
xnor U18637 (N_18637,N_16955,N_17570);
or U18638 (N_18638,N_17453,N_17390);
nand U18639 (N_18639,N_17067,N_17696);
and U18640 (N_18640,N_17278,N_17668);
nor U18641 (N_18641,N_17979,N_17968);
nand U18642 (N_18642,N_17810,N_16883);
or U18643 (N_18643,N_17899,N_17905);
or U18644 (N_18644,N_17192,N_17211);
and U18645 (N_18645,N_17482,N_17375);
and U18646 (N_18646,N_17195,N_17727);
or U18647 (N_18647,N_17368,N_16836);
nand U18648 (N_18648,N_17103,N_17936);
and U18649 (N_18649,N_17895,N_17788);
xor U18650 (N_18650,N_16972,N_17486);
and U18651 (N_18651,N_17573,N_17564);
or U18652 (N_18652,N_17802,N_17037);
or U18653 (N_18653,N_16920,N_17981);
or U18654 (N_18654,N_17591,N_17246);
xor U18655 (N_18655,N_17373,N_17561);
or U18656 (N_18656,N_16994,N_17957);
nand U18657 (N_18657,N_17755,N_16825);
nand U18658 (N_18658,N_17752,N_17433);
nor U18659 (N_18659,N_17929,N_16806);
or U18660 (N_18660,N_17218,N_17803);
and U18661 (N_18661,N_16956,N_17012);
nor U18662 (N_18662,N_17833,N_17608);
nor U18663 (N_18663,N_17448,N_17458);
and U18664 (N_18664,N_16872,N_17598);
xnor U18665 (N_18665,N_17792,N_17454);
and U18666 (N_18666,N_16827,N_17329);
nand U18667 (N_18667,N_17109,N_17078);
xnor U18668 (N_18668,N_16941,N_17396);
nor U18669 (N_18669,N_17885,N_17711);
xor U18670 (N_18670,N_17012,N_17216);
nand U18671 (N_18671,N_17284,N_17133);
xnor U18672 (N_18672,N_17053,N_17985);
nor U18673 (N_18673,N_16848,N_17377);
nor U18674 (N_18674,N_17034,N_17544);
nor U18675 (N_18675,N_17820,N_17209);
xnor U18676 (N_18676,N_17380,N_17141);
and U18677 (N_18677,N_17456,N_17387);
nand U18678 (N_18678,N_16916,N_17847);
or U18679 (N_18679,N_17027,N_17402);
nand U18680 (N_18680,N_17949,N_17490);
nor U18681 (N_18681,N_17414,N_16946);
nand U18682 (N_18682,N_17709,N_17920);
nor U18683 (N_18683,N_17320,N_17082);
xnor U18684 (N_18684,N_16827,N_17726);
nor U18685 (N_18685,N_17015,N_17636);
xor U18686 (N_18686,N_16944,N_17418);
or U18687 (N_18687,N_17245,N_17866);
or U18688 (N_18688,N_17723,N_17220);
and U18689 (N_18689,N_16899,N_16866);
and U18690 (N_18690,N_17477,N_17767);
nor U18691 (N_18691,N_16822,N_17426);
xor U18692 (N_18692,N_17297,N_17762);
and U18693 (N_18693,N_17283,N_17515);
and U18694 (N_18694,N_16921,N_17267);
or U18695 (N_18695,N_17518,N_17066);
nand U18696 (N_18696,N_17277,N_17289);
or U18697 (N_18697,N_17415,N_16866);
xnor U18698 (N_18698,N_16810,N_16968);
nand U18699 (N_18699,N_17865,N_17912);
and U18700 (N_18700,N_17030,N_17633);
xor U18701 (N_18701,N_17454,N_17060);
and U18702 (N_18702,N_17914,N_17372);
nand U18703 (N_18703,N_17564,N_17045);
nand U18704 (N_18704,N_17646,N_17360);
nor U18705 (N_18705,N_17761,N_17163);
nand U18706 (N_18706,N_17796,N_17759);
or U18707 (N_18707,N_17013,N_16943);
and U18708 (N_18708,N_17029,N_17293);
nand U18709 (N_18709,N_17855,N_17021);
or U18710 (N_18710,N_17074,N_17839);
nor U18711 (N_18711,N_17213,N_17453);
nor U18712 (N_18712,N_17246,N_17740);
xnor U18713 (N_18713,N_17698,N_17997);
nand U18714 (N_18714,N_17630,N_17776);
nand U18715 (N_18715,N_17890,N_17637);
nor U18716 (N_18716,N_17194,N_17230);
nand U18717 (N_18717,N_17848,N_16969);
nor U18718 (N_18718,N_17127,N_17837);
nor U18719 (N_18719,N_16852,N_16841);
or U18720 (N_18720,N_17178,N_17319);
nand U18721 (N_18721,N_17564,N_17625);
and U18722 (N_18722,N_17980,N_17393);
and U18723 (N_18723,N_17667,N_16936);
nor U18724 (N_18724,N_17010,N_17658);
and U18725 (N_18725,N_16932,N_17953);
or U18726 (N_18726,N_17453,N_17633);
or U18727 (N_18727,N_17471,N_17445);
or U18728 (N_18728,N_17736,N_17584);
xnor U18729 (N_18729,N_16903,N_17251);
nand U18730 (N_18730,N_16990,N_17482);
xor U18731 (N_18731,N_17459,N_17918);
xnor U18732 (N_18732,N_17246,N_16852);
and U18733 (N_18733,N_17744,N_16831);
xnor U18734 (N_18734,N_17230,N_17415);
nand U18735 (N_18735,N_16853,N_17652);
or U18736 (N_18736,N_17199,N_16928);
xor U18737 (N_18737,N_17787,N_17902);
nand U18738 (N_18738,N_17463,N_17563);
nor U18739 (N_18739,N_17079,N_17918);
nor U18740 (N_18740,N_17762,N_16939);
xor U18741 (N_18741,N_17972,N_17322);
nand U18742 (N_18742,N_17793,N_17922);
xor U18743 (N_18743,N_17224,N_17463);
nor U18744 (N_18744,N_16890,N_17123);
nor U18745 (N_18745,N_17681,N_17834);
and U18746 (N_18746,N_16883,N_16820);
nor U18747 (N_18747,N_17958,N_17557);
nor U18748 (N_18748,N_17992,N_17129);
xor U18749 (N_18749,N_16836,N_17987);
nor U18750 (N_18750,N_17001,N_17699);
or U18751 (N_18751,N_17309,N_17844);
nand U18752 (N_18752,N_17121,N_17454);
nand U18753 (N_18753,N_17043,N_17877);
or U18754 (N_18754,N_17394,N_17693);
and U18755 (N_18755,N_17989,N_17118);
nor U18756 (N_18756,N_16965,N_17626);
and U18757 (N_18757,N_17001,N_17300);
xnor U18758 (N_18758,N_17964,N_17096);
and U18759 (N_18759,N_16889,N_17849);
and U18760 (N_18760,N_17808,N_17066);
nand U18761 (N_18761,N_17348,N_17673);
and U18762 (N_18762,N_17327,N_16837);
nand U18763 (N_18763,N_16810,N_17156);
xor U18764 (N_18764,N_17704,N_17006);
xor U18765 (N_18765,N_17619,N_17165);
xor U18766 (N_18766,N_17967,N_17881);
nor U18767 (N_18767,N_17396,N_17074);
nand U18768 (N_18768,N_17144,N_17474);
nor U18769 (N_18769,N_16880,N_17562);
or U18770 (N_18770,N_16821,N_17587);
and U18771 (N_18771,N_17809,N_16851);
or U18772 (N_18772,N_17930,N_17740);
xnor U18773 (N_18773,N_16893,N_17480);
nand U18774 (N_18774,N_17599,N_16907);
and U18775 (N_18775,N_16822,N_17548);
xnor U18776 (N_18776,N_16877,N_16881);
and U18777 (N_18777,N_17001,N_16916);
xor U18778 (N_18778,N_17556,N_17294);
or U18779 (N_18779,N_17301,N_17180);
and U18780 (N_18780,N_17830,N_16960);
or U18781 (N_18781,N_16825,N_17547);
or U18782 (N_18782,N_17967,N_17659);
nor U18783 (N_18783,N_17277,N_17578);
or U18784 (N_18784,N_17745,N_17915);
and U18785 (N_18785,N_17376,N_17306);
xor U18786 (N_18786,N_16920,N_17717);
or U18787 (N_18787,N_17888,N_17372);
nand U18788 (N_18788,N_17406,N_17637);
nor U18789 (N_18789,N_16884,N_17954);
nand U18790 (N_18790,N_16881,N_17203);
xnor U18791 (N_18791,N_17923,N_17591);
and U18792 (N_18792,N_17282,N_17139);
or U18793 (N_18793,N_16964,N_17673);
xnor U18794 (N_18794,N_17312,N_17572);
and U18795 (N_18795,N_16904,N_17458);
nor U18796 (N_18796,N_17924,N_17649);
and U18797 (N_18797,N_17996,N_17302);
nor U18798 (N_18798,N_17950,N_17229);
xor U18799 (N_18799,N_17516,N_17102);
nand U18800 (N_18800,N_17951,N_17429);
or U18801 (N_18801,N_17822,N_17134);
nand U18802 (N_18802,N_17757,N_17608);
nand U18803 (N_18803,N_17038,N_17309);
nand U18804 (N_18804,N_17632,N_17182);
or U18805 (N_18805,N_17114,N_16924);
or U18806 (N_18806,N_17381,N_17777);
nand U18807 (N_18807,N_17186,N_16956);
nor U18808 (N_18808,N_17732,N_16849);
nor U18809 (N_18809,N_17443,N_16968);
and U18810 (N_18810,N_17137,N_17616);
and U18811 (N_18811,N_17520,N_17500);
xor U18812 (N_18812,N_17120,N_17721);
and U18813 (N_18813,N_17892,N_17186);
nand U18814 (N_18814,N_16970,N_17539);
nor U18815 (N_18815,N_17454,N_17103);
nand U18816 (N_18816,N_17916,N_17460);
nand U18817 (N_18817,N_17972,N_17131);
or U18818 (N_18818,N_17036,N_16894);
nand U18819 (N_18819,N_17746,N_17597);
xor U18820 (N_18820,N_17075,N_17111);
and U18821 (N_18821,N_17729,N_17042);
or U18822 (N_18822,N_16943,N_17309);
xnor U18823 (N_18823,N_17575,N_17764);
nand U18824 (N_18824,N_17465,N_16928);
xnor U18825 (N_18825,N_17743,N_16871);
nor U18826 (N_18826,N_17410,N_17183);
and U18827 (N_18827,N_17002,N_17883);
xnor U18828 (N_18828,N_17418,N_17877);
and U18829 (N_18829,N_17203,N_17663);
or U18830 (N_18830,N_17454,N_16987);
xor U18831 (N_18831,N_17012,N_17265);
nor U18832 (N_18832,N_17083,N_17133);
and U18833 (N_18833,N_17145,N_17894);
nor U18834 (N_18834,N_17362,N_16809);
xnor U18835 (N_18835,N_17437,N_17461);
or U18836 (N_18836,N_17931,N_17634);
nor U18837 (N_18837,N_17766,N_17425);
nor U18838 (N_18838,N_17776,N_17010);
nor U18839 (N_18839,N_17866,N_17022);
and U18840 (N_18840,N_17159,N_17661);
nand U18841 (N_18841,N_17265,N_17707);
nand U18842 (N_18842,N_17640,N_17619);
and U18843 (N_18843,N_17004,N_16994);
xnor U18844 (N_18844,N_17466,N_17396);
nor U18845 (N_18845,N_17032,N_17893);
xor U18846 (N_18846,N_17743,N_17430);
xnor U18847 (N_18847,N_17549,N_17416);
and U18848 (N_18848,N_16937,N_17094);
nor U18849 (N_18849,N_17137,N_17649);
nand U18850 (N_18850,N_17898,N_17932);
or U18851 (N_18851,N_17594,N_17244);
or U18852 (N_18852,N_17112,N_17548);
xor U18853 (N_18853,N_17532,N_17758);
xnor U18854 (N_18854,N_17951,N_17140);
xor U18855 (N_18855,N_17808,N_17593);
and U18856 (N_18856,N_17852,N_16992);
nand U18857 (N_18857,N_17001,N_17574);
xnor U18858 (N_18858,N_17794,N_17476);
xnor U18859 (N_18859,N_17986,N_17434);
or U18860 (N_18860,N_16815,N_17084);
or U18861 (N_18861,N_17624,N_17102);
xor U18862 (N_18862,N_17706,N_17847);
xnor U18863 (N_18863,N_17816,N_17209);
or U18864 (N_18864,N_17456,N_17706);
and U18865 (N_18865,N_17132,N_17227);
or U18866 (N_18866,N_16819,N_17112);
nand U18867 (N_18867,N_17462,N_16860);
or U18868 (N_18868,N_17987,N_16922);
or U18869 (N_18869,N_17129,N_17080);
or U18870 (N_18870,N_17595,N_17101);
xor U18871 (N_18871,N_17984,N_17314);
xor U18872 (N_18872,N_16903,N_17469);
nand U18873 (N_18873,N_17280,N_16991);
or U18874 (N_18874,N_17076,N_17613);
nand U18875 (N_18875,N_17369,N_17557);
nand U18876 (N_18876,N_17293,N_17460);
xnor U18877 (N_18877,N_17624,N_16807);
xnor U18878 (N_18878,N_17863,N_16810);
or U18879 (N_18879,N_16985,N_16948);
nand U18880 (N_18880,N_16949,N_17988);
or U18881 (N_18881,N_17274,N_16981);
xor U18882 (N_18882,N_17731,N_16808);
and U18883 (N_18883,N_17261,N_17974);
xor U18884 (N_18884,N_17051,N_17132);
and U18885 (N_18885,N_17059,N_16968);
or U18886 (N_18886,N_17388,N_17179);
and U18887 (N_18887,N_17200,N_17408);
xnor U18888 (N_18888,N_17904,N_17087);
xnor U18889 (N_18889,N_17380,N_16957);
and U18890 (N_18890,N_17509,N_17463);
xnor U18891 (N_18891,N_17375,N_17080);
xnor U18892 (N_18892,N_17335,N_16822);
nand U18893 (N_18893,N_17623,N_17949);
and U18894 (N_18894,N_17469,N_17696);
or U18895 (N_18895,N_16941,N_17309);
nand U18896 (N_18896,N_17953,N_17229);
nand U18897 (N_18897,N_17410,N_17195);
nand U18898 (N_18898,N_16983,N_16978);
or U18899 (N_18899,N_16937,N_17312);
or U18900 (N_18900,N_17562,N_17732);
nor U18901 (N_18901,N_17455,N_17023);
or U18902 (N_18902,N_17127,N_17171);
or U18903 (N_18903,N_17235,N_17606);
and U18904 (N_18904,N_17174,N_17466);
xnor U18905 (N_18905,N_17161,N_17960);
nand U18906 (N_18906,N_17599,N_17192);
or U18907 (N_18907,N_16919,N_17020);
nor U18908 (N_18908,N_16840,N_16924);
and U18909 (N_18909,N_17967,N_17537);
and U18910 (N_18910,N_17126,N_17593);
xor U18911 (N_18911,N_17402,N_17386);
or U18912 (N_18912,N_16849,N_17295);
nor U18913 (N_18913,N_17707,N_16938);
nor U18914 (N_18914,N_16931,N_16873);
nor U18915 (N_18915,N_17812,N_17180);
xor U18916 (N_18916,N_17977,N_17598);
or U18917 (N_18917,N_17889,N_17043);
xor U18918 (N_18918,N_17728,N_17138);
nand U18919 (N_18919,N_17031,N_17084);
nor U18920 (N_18920,N_17910,N_17803);
and U18921 (N_18921,N_17330,N_16859);
and U18922 (N_18922,N_17244,N_17490);
xnor U18923 (N_18923,N_17344,N_17793);
xor U18924 (N_18924,N_17242,N_17869);
nor U18925 (N_18925,N_16996,N_17053);
and U18926 (N_18926,N_17951,N_17431);
nand U18927 (N_18927,N_17080,N_17703);
or U18928 (N_18928,N_17642,N_17327);
and U18929 (N_18929,N_17801,N_17200);
nand U18930 (N_18930,N_17695,N_17365);
nand U18931 (N_18931,N_17089,N_17809);
and U18932 (N_18932,N_17613,N_17140);
nand U18933 (N_18933,N_17847,N_17368);
nand U18934 (N_18934,N_17439,N_17826);
and U18935 (N_18935,N_17018,N_17307);
xor U18936 (N_18936,N_17088,N_17134);
nand U18937 (N_18937,N_17390,N_17876);
or U18938 (N_18938,N_17960,N_17049);
nor U18939 (N_18939,N_17708,N_16960);
xnor U18940 (N_18940,N_17425,N_17629);
xor U18941 (N_18941,N_17407,N_16877);
nor U18942 (N_18942,N_17785,N_17013);
nor U18943 (N_18943,N_16983,N_16856);
or U18944 (N_18944,N_17580,N_17071);
or U18945 (N_18945,N_17664,N_17331);
xnor U18946 (N_18946,N_17102,N_17740);
nor U18947 (N_18947,N_17488,N_17330);
xor U18948 (N_18948,N_17604,N_17244);
nor U18949 (N_18949,N_17236,N_17888);
nand U18950 (N_18950,N_17002,N_17842);
or U18951 (N_18951,N_17056,N_16921);
nor U18952 (N_18952,N_16980,N_17339);
nand U18953 (N_18953,N_17624,N_17056);
nand U18954 (N_18954,N_17422,N_17315);
or U18955 (N_18955,N_17066,N_17210);
nand U18956 (N_18956,N_17153,N_17971);
and U18957 (N_18957,N_17735,N_17538);
and U18958 (N_18958,N_16823,N_17456);
or U18959 (N_18959,N_17164,N_16853);
nor U18960 (N_18960,N_17393,N_17849);
or U18961 (N_18961,N_17903,N_17961);
nor U18962 (N_18962,N_17521,N_17516);
nor U18963 (N_18963,N_17655,N_17680);
or U18964 (N_18964,N_17108,N_17488);
and U18965 (N_18965,N_17644,N_17046);
or U18966 (N_18966,N_17766,N_17405);
or U18967 (N_18967,N_17116,N_17959);
nor U18968 (N_18968,N_17443,N_17380);
nor U18969 (N_18969,N_17603,N_17374);
and U18970 (N_18970,N_17962,N_17071);
or U18971 (N_18971,N_16854,N_17306);
or U18972 (N_18972,N_16866,N_17313);
and U18973 (N_18973,N_17486,N_17505);
or U18974 (N_18974,N_17240,N_16923);
xor U18975 (N_18975,N_17528,N_17103);
or U18976 (N_18976,N_17891,N_17424);
or U18977 (N_18977,N_17704,N_17035);
xnor U18978 (N_18978,N_17516,N_17392);
xor U18979 (N_18979,N_17317,N_17508);
nor U18980 (N_18980,N_17157,N_17204);
nor U18981 (N_18981,N_17601,N_17967);
and U18982 (N_18982,N_17217,N_17852);
xnor U18983 (N_18983,N_17154,N_17563);
xnor U18984 (N_18984,N_17883,N_17737);
or U18985 (N_18985,N_17839,N_17102);
xor U18986 (N_18986,N_17097,N_17727);
and U18987 (N_18987,N_17071,N_17849);
or U18988 (N_18988,N_16889,N_16806);
and U18989 (N_18989,N_16834,N_17096);
and U18990 (N_18990,N_17223,N_17633);
nand U18991 (N_18991,N_17487,N_17503);
and U18992 (N_18992,N_17742,N_16973);
nand U18993 (N_18993,N_16885,N_16817);
or U18994 (N_18994,N_17841,N_17118);
nor U18995 (N_18995,N_17487,N_17979);
or U18996 (N_18996,N_17479,N_17530);
nor U18997 (N_18997,N_16812,N_17163);
nand U18998 (N_18998,N_17224,N_17281);
nor U18999 (N_18999,N_17464,N_17869);
nor U19000 (N_19000,N_17000,N_17972);
nor U19001 (N_19001,N_17962,N_17078);
or U19002 (N_19002,N_17046,N_17563);
xor U19003 (N_19003,N_17495,N_17558);
nor U19004 (N_19004,N_17706,N_17499);
or U19005 (N_19005,N_17825,N_17673);
and U19006 (N_19006,N_17810,N_17049);
nor U19007 (N_19007,N_16982,N_17249);
nand U19008 (N_19008,N_17356,N_17408);
and U19009 (N_19009,N_17888,N_17946);
and U19010 (N_19010,N_17859,N_17415);
xnor U19011 (N_19011,N_17959,N_17756);
or U19012 (N_19012,N_16924,N_17386);
and U19013 (N_19013,N_17744,N_16874);
nor U19014 (N_19014,N_17298,N_17823);
or U19015 (N_19015,N_17865,N_17591);
nor U19016 (N_19016,N_17992,N_17202);
xor U19017 (N_19017,N_17435,N_17515);
nor U19018 (N_19018,N_17267,N_17987);
xor U19019 (N_19019,N_17681,N_17769);
xnor U19020 (N_19020,N_17898,N_17722);
nand U19021 (N_19021,N_17047,N_16874);
and U19022 (N_19022,N_17633,N_17628);
nor U19023 (N_19023,N_17604,N_17785);
nand U19024 (N_19024,N_17235,N_16813);
or U19025 (N_19025,N_17497,N_17270);
xnor U19026 (N_19026,N_17838,N_17751);
and U19027 (N_19027,N_17603,N_16841);
or U19028 (N_19028,N_17645,N_17572);
xnor U19029 (N_19029,N_17326,N_17746);
nand U19030 (N_19030,N_17243,N_17959);
nand U19031 (N_19031,N_17455,N_16960);
or U19032 (N_19032,N_17850,N_17337);
xnor U19033 (N_19033,N_17107,N_17374);
xnor U19034 (N_19034,N_16854,N_17060);
nor U19035 (N_19035,N_16802,N_17762);
or U19036 (N_19036,N_17983,N_17510);
nor U19037 (N_19037,N_17291,N_17871);
or U19038 (N_19038,N_16860,N_17458);
or U19039 (N_19039,N_17757,N_17214);
nand U19040 (N_19040,N_17611,N_17541);
xnor U19041 (N_19041,N_17511,N_17718);
nand U19042 (N_19042,N_17675,N_17179);
xor U19043 (N_19043,N_17708,N_17121);
xor U19044 (N_19044,N_16806,N_17489);
nor U19045 (N_19045,N_17297,N_17253);
xnor U19046 (N_19046,N_16915,N_17980);
nor U19047 (N_19047,N_17800,N_16866);
and U19048 (N_19048,N_17348,N_17431);
nor U19049 (N_19049,N_17379,N_17774);
xor U19050 (N_19050,N_17221,N_16912);
and U19051 (N_19051,N_17185,N_17979);
nand U19052 (N_19052,N_17842,N_17297);
xnor U19053 (N_19053,N_17537,N_17652);
and U19054 (N_19054,N_16918,N_17912);
nor U19055 (N_19055,N_17116,N_16939);
xor U19056 (N_19056,N_17867,N_17841);
nor U19057 (N_19057,N_17954,N_17361);
xnor U19058 (N_19058,N_16817,N_17678);
nor U19059 (N_19059,N_17783,N_17524);
or U19060 (N_19060,N_17192,N_17513);
and U19061 (N_19061,N_17992,N_16871);
nor U19062 (N_19062,N_17303,N_17890);
and U19063 (N_19063,N_17363,N_17610);
and U19064 (N_19064,N_17271,N_17260);
or U19065 (N_19065,N_17664,N_17469);
xor U19066 (N_19066,N_17812,N_17055);
xor U19067 (N_19067,N_17968,N_17854);
xnor U19068 (N_19068,N_17093,N_17319);
and U19069 (N_19069,N_16915,N_17767);
and U19070 (N_19070,N_17659,N_17251);
or U19071 (N_19071,N_17568,N_17988);
or U19072 (N_19072,N_17435,N_16835);
nor U19073 (N_19073,N_17531,N_17259);
and U19074 (N_19074,N_17918,N_17488);
xnor U19075 (N_19075,N_17757,N_17341);
and U19076 (N_19076,N_16981,N_17130);
or U19077 (N_19077,N_17333,N_17406);
nor U19078 (N_19078,N_17329,N_17126);
xor U19079 (N_19079,N_17644,N_17126);
xnor U19080 (N_19080,N_17533,N_17615);
or U19081 (N_19081,N_17315,N_17416);
or U19082 (N_19082,N_17031,N_17524);
or U19083 (N_19083,N_17579,N_16936);
nor U19084 (N_19084,N_16935,N_17503);
nor U19085 (N_19085,N_17499,N_16857);
nor U19086 (N_19086,N_17221,N_17958);
or U19087 (N_19087,N_17871,N_17360);
nand U19088 (N_19088,N_17420,N_16956);
nor U19089 (N_19089,N_17605,N_17656);
nor U19090 (N_19090,N_17906,N_17474);
xnor U19091 (N_19091,N_17897,N_17842);
and U19092 (N_19092,N_17114,N_17459);
nand U19093 (N_19093,N_17984,N_16931);
and U19094 (N_19094,N_17576,N_17470);
and U19095 (N_19095,N_17442,N_17462);
or U19096 (N_19096,N_17602,N_17985);
nor U19097 (N_19097,N_17383,N_17584);
nand U19098 (N_19098,N_17871,N_17044);
or U19099 (N_19099,N_17459,N_17250);
and U19100 (N_19100,N_17217,N_17474);
nor U19101 (N_19101,N_17712,N_17388);
nor U19102 (N_19102,N_17752,N_16967);
nor U19103 (N_19103,N_17849,N_17930);
nand U19104 (N_19104,N_17660,N_17524);
and U19105 (N_19105,N_17456,N_17507);
nand U19106 (N_19106,N_16992,N_16904);
nor U19107 (N_19107,N_17739,N_17368);
xor U19108 (N_19108,N_17974,N_17304);
or U19109 (N_19109,N_17413,N_17628);
or U19110 (N_19110,N_17830,N_17009);
or U19111 (N_19111,N_17048,N_17434);
and U19112 (N_19112,N_16954,N_17928);
xnor U19113 (N_19113,N_17617,N_17513);
or U19114 (N_19114,N_17646,N_16892);
xor U19115 (N_19115,N_16896,N_17379);
nand U19116 (N_19116,N_17990,N_17905);
xor U19117 (N_19117,N_17248,N_17091);
xnor U19118 (N_19118,N_17915,N_17576);
or U19119 (N_19119,N_16893,N_17363);
xor U19120 (N_19120,N_17934,N_17907);
nand U19121 (N_19121,N_17971,N_17680);
or U19122 (N_19122,N_16940,N_17678);
and U19123 (N_19123,N_17788,N_17702);
and U19124 (N_19124,N_16825,N_17943);
or U19125 (N_19125,N_17762,N_17264);
xnor U19126 (N_19126,N_16820,N_17611);
or U19127 (N_19127,N_17031,N_17184);
xnor U19128 (N_19128,N_17193,N_17385);
nor U19129 (N_19129,N_17639,N_17303);
and U19130 (N_19130,N_17862,N_17420);
or U19131 (N_19131,N_17654,N_17450);
or U19132 (N_19132,N_17870,N_17687);
or U19133 (N_19133,N_17657,N_17630);
or U19134 (N_19134,N_17505,N_17871);
or U19135 (N_19135,N_17053,N_17074);
nand U19136 (N_19136,N_17533,N_17086);
or U19137 (N_19137,N_17198,N_16879);
nor U19138 (N_19138,N_16913,N_17312);
nor U19139 (N_19139,N_17629,N_17743);
or U19140 (N_19140,N_17187,N_17483);
or U19141 (N_19141,N_17916,N_17061);
xnor U19142 (N_19142,N_17177,N_17893);
or U19143 (N_19143,N_17817,N_17239);
nor U19144 (N_19144,N_16883,N_17487);
xor U19145 (N_19145,N_17013,N_17169);
xor U19146 (N_19146,N_17995,N_17974);
and U19147 (N_19147,N_17965,N_17508);
xor U19148 (N_19148,N_17202,N_17606);
nor U19149 (N_19149,N_17849,N_17990);
or U19150 (N_19150,N_16898,N_17775);
and U19151 (N_19151,N_17454,N_16821);
or U19152 (N_19152,N_17321,N_17019);
nand U19153 (N_19153,N_17046,N_17211);
or U19154 (N_19154,N_17007,N_17052);
nand U19155 (N_19155,N_17058,N_17792);
nor U19156 (N_19156,N_16955,N_17622);
or U19157 (N_19157,N_16907,N_17759);
or U19158 (N_19158,N_17589,N_17186);
or U19159 (N_19159,N_16843,N_16818);
or U19160 (N_19160,N_17117,N_17504);
nand U19161 (N_19161,N_17337,N_17446);
nand U19162 (N_19162,N_16865,N_17043);
and U19163 (N_19163,N_17990,N_17630);
or U19164 (N_19164,N_16970,N_17447);
nor U19165 (N_19165,N_16836,N_17155);
or U19166 (N_19166,N_17225,N_17376);
and U19167 (N_19167,N_16927,N_17025);
and U19168 (N_19168,N_16958,N_17594);
nor U19169 (N_19169,N_16851,N_17094);
nor U19170 (N_19170,N_17300,N_17667);
nand U19171 (N_19171,N_17713,N_17167);
nand U19172 (N_19172,N_16975,N_17428);
nor U19173 (N_19173,N_17260,N_16974);
xor U19174 (N_19174,N_16943,N_17312);
nor U19175 (N_19175,N_17509,N_17860);
nor U19176 (N_19176,N_17699,N_17616);
nand U19177 (N_19177,N_17749,N_17171);
xor U19178 (N_19178,N_17771,N_17757);
or U19179 (N_19179,N_16864,N_17549);
and U19180 (N_19180,N_17371,N_16940);
or U19181 (N_19181,N_17735,N_17396);
xnor U19182 (N_19182,N_16864,N_16874);
nand U19183 (N_19183,N_17343,N_17338);
and U19184 (N_19184,N_17150,N_17892);
or U19185 (N_19185,N_16963,N_17534);
nor U19186 (N_19186,N_17650,N_17289);
nand U19187 (N_19187,N_17277,N_16841);
xnor U19188 (N_19188,N_17266,N_17599);
nor U19189 (N_19189,N_17742,N_16836);
and U19190 (N_19190,N_17724,N_17307);
xor U19191 (N_19191,N_17430,N_17365);
or U19192 (N_19192,N_17096,N_17924);
and U19193 (N_19193,N_17151,N_17736);
nand U19194 (N_19194,N_17224,N_17320);
nand U19195 (N_19195,N_17607,N_17767);
or U19196 (N_19196,N_17830,N_17271);
and U19197 (N_19197,N_17361,N_17049);
and U19198 (N_19198,N_17540,N_17103);
or U19199 (N_19199,N_16821,N_17545);
or U19200 (N_19200,N_18268,N_18117);
nand U19201 (N_19201,N_19037,N_18493);
nor U19202 (N_19202,N_18567,N_18911);
nand U19203 (N_19203,N_19128,N_18201);
nand U19204 (N_19204,N_18831,N_18052);
xnor U19205 (N_19205,N_18637,N_19182);
and U19206 (N_19206,N_19160,N_18149);
xnor U19207 (N_19207,N_18711,N_18286);
and U19208 (N_19208,N_18144,N_18293);
or U19209 (N_19209,N_18501,N_18071);
nand U19210 (N_19210,N_19167,N_19046);
nor U19211 (N_19211,N_18464,N_18307);
nand U19212 (N_19212,N_18992,N_18685);
nor U19213 (N_19213,N_18826,N_19100);
xnor U19214 (N_19214,N_18323,N_18243);
nor U19215 (N_19215,N_18388,N_19047);
or U19216 (N_19216,N_18748,N_19003);
xor U19217 (N_19217,N_18446,N_18219);
nor U19218 (N_19218,N_18866,N_18542);
nor U19219 (N_19219,N_18533,N_18861);
and U19220 (N_19220,N_18937,N_18130);
and U19221 (N_19221,N_19148,N_18284);
nand U19222 (N_19222,N_18447,N_18562);
xnor U19223 (N_19223,N_18109,N_18234);
or U19224 (N_19224,N_19051,N_18101);
nand U19225 (N_19225,N_18420,N_19087);
nand U19226 (N_19226,N_19183,N_18348);
and U19227 (N_19227,N_19112,N_18032);
and U19228 (N_19228,N_19159,N_18322);
nand U19229 (N_19229,N_18521,N_18356);
or U19230 (N_19230,N_18191,N_18702);
xnor U19231 (N_19231,N_18865,N_18821);
nand U19232 (N_19232,N_18553,N_19166);
nor U19233 (N_19233,N_19065,N_18504);
and U19234 (N_19234,N_19172,N_18855);
and U19235 (N_19235,N_18918,N_18329);
or U19236 (N_19236,N_18262,N_18183);
nand U19237 (N_19237,N_18700,N_18409);
nor U19238 (N_19238,N_18291,N_19060);
and U19239 (N_19239,N_19009,N_18424);
nand U19240 (N_19240,N_18445,N_18078);
xnor U19241 (N_19241,N_18554,N_18742);
or U19242 (N_19242,N_18058,N_18684);
or U19243 (N_19243,N_18298,N_18867);
xor U19244 (N_19244,N_18245,N_18378);
xnor U19245 (N_19245,N_18210,N_18308);
xnor U19246 (N_19246,N_18043,N_18285);
and U19247 (N_19247,N_19106,N_18580);
or U19248 (N_19248,N_18393,N_19143);
nand U19249 (N_19249,N_18668,N_18946);
or U19250 (N_19250,N_18523,N_19028);
nand U19251 (N_19251,N_18033,N_18749);
or U19252 (N_19252,N_19080,N_18551);
nand U19253 (N_19253,N_19135,N_18640);
nand U19254 (N_19254,N_19178,N_18670);
or U19255 (N_19255,N_18190,N_18386);
xor U19256 (N_19256,N_18251,N_18380);
and U19257 (N_19257,N_19125,N_18539);
or U19258 (N_19258,N_18652,N_18878);
nand U19259 (N_19259,N_18026,N_18951);
or U19260 (N_19260,N_19042,N_18087);
nand U19261 (N_19261,N_18544,N_19108);
nand U19262 (N_19262,N_19161,N_18028);
nor U19263 (N_19263,N_18153,N_18686);
nor U19264 (N_19264,N_18770,N_18324);
or U19265 (N_19265,N_19070,N_18633);
and U19266 (N_19266,N_18828,N_19038);
and U19267 (N_19267,N_18563,N_18723);
and U19268 (N_19268,N_18766,N_18140);
or U19269 (N_19269,N_18823,N_18790);
or U19270 (N_19270,N_19000,N_18600);
xor U19271 (N_19271,N_18269,N_18736);
xnor U19272 (N_19272,N_18949,N_18247);
xor U19273 (N_19273,N_18564,N_18205);
and U19274 (N_19274,N_18891,N_19036);
or U19275 (N_19275,N_18660,N_18977);
and U19276 (N_19276,N_18494,N_18240);
xnor U19277 (N_19277,N_18187,N_18296);
or U19278 (N_19278,N_18721,N_18787);
or U19279 (N_19279,N_18089,N_18925);
and U19280 (N_19280,N_18436,N_18344);
nand U19281 (N_19281,N_18485,N_19029);
nor U19282 (N_19282,N_18777,N_19123);
or U19283 (N_19283,N_19071,N_19191);
or U19284 (N_19284,N_18304,N_18801);
xor U19285 (N_19285,N_18145,N_19120);
nor U19286 (N_19286,N_18569,N_18159);
or U19287 (N_19287,N_18055,N_18710);
xor U19288 (N_19288,N_19156,N_18706);
xor U19289 (N_19289,N_18889,N_18317);
and U19290 (N_19290,N_18080,N_18856);
nor U19291 (N_19291,N_18060,N_18953);
nand U19292 (N_19292,N_19077,N_18178);
xor U19293 (N_19293,N_18428,N_18834);
xnor U19294 (N_19294,N_18372,N_18273);
xor U19295 (N_19295,N_18110,N_18796);
nand U19296 (N_19296,N_18797,N_18756);
or U19297 (N_19297,N_19119,N_18241);
nand U19298 (N_19298,N_18361,N_18687);
nand U19299 (N_19299,N_18235,N_18371);
or U19300 (N_19300,N_19078,N_18500);
and U19301 (N_19301,N_18387,N_18582);
or U19302 (N_19302,N_19084,N_18068);
nor U19303 (N_19303,N_18715,N_18041);
nand U19304 (N_19304,N_18595,N_19032);
nand U19305 (N_19305,N_18261,N_18738);
nand U19306 (N_19306,N_18963,N_18490);
nand U19307 (N_19307,N_19139,N_18905);
nor U19308 (N_19308,N_18276,N_18990);
nand U19309 (N_19309,N_18817,N_19059);
nor U19310 (N_19310,N_18466,N_18627);
or U19311 (N_19311,N_18568,N_18746);
nor U19312 (N_19312,N_18753,N_18368);
nand U19313 (N_19313,N_18793,N_18351);
and U19314 (N_19314,N_18666,N_18152);
nor U19315 (N_19315,N_18642,N_18000);
nor U19316 (N_19316,N_19013,N_18852);
or U19317 (N_19317,N_18989,N_19014);
or U19318 (N_19318,N_18385,N_18237);
nand U19319 (N_19319,N_18007,N_18907);
or U19320 (N_19320,N_18585,N_18292);
xnor U19321 (N_19321,N_19027,N_18807);
xor U19322 (N_19322,N_19010,N_18921);
xor U19323 (N_19323,N_18195,N_18476);
nor U19324 (N_19324,N_18935,N_18279);
and U19325 (N_19325,N_18957,N_18054);
and U19326 (N_19326,N_18625,N_18440);
or U19327 (N_19327,N_18875,N_18389);
xor U19328 (N_19328,N_18454,N_19099);
xnor U19329 (N_19329,N_19169,N_18531);
xnor U19330 (N_19330,N_18690,N_18184);
and U19331 (N_19331,N_18948,N_18325);
nor U19332 (N_19332,N_18981,N_18773);
nand U19333 (N_19333,N_18207,N_18526);
nand U19334 (N_19334,N_18091,N_18776);
nand U19335 (N_19335,N_18837,N_18747);
nand U19336 (N_19336,N_18806,N_18864);
or U19337 (N_19337,N_18758,N_18976);
or U19338 (N_19338,N_19041,N_19045);
nor U19339 (N_19339,N_18212,N_18919);
or U19340 (N_19340,N_18941,N_18970);
xor U19341 (N_19341,N_18106,N_18674);
nand U19342 (N_19342,N_18509,N_18172);
nand U19343 (N_19343,N_18426,N_18636);
or U19344 (N_19344,N_18162,N_18347);
or U19345 (N_19345,N_18359,N_19083);
nand U19346 (N_19346,N_18743,N_18546);
nor U19347 (N_19347,N_18651,N_19104);
nand U19348 (N_19348,N_19016,N_19069);
nor U19349 (N_19349,N_18714,N_18363);
nand U19350 (N_19350,N_18175,N_18137);
or U19351 (N_19351,N_18857,N_18073);
and U19352 (N_19352,N_18006,N_18362);
nor U19353 (N_19353,N_19068,N_19035);
nand U19354 (N_19354,N_18759,N_18350);
nor U19355 (N_19355,N_19179,N_18044);
xnor U19356 (N_19356,N_18467,N_18489);
xnor U19357 (N_19357,N_18532,N_18181);
xnor U19358 (N_19358,N_19199,N_19103);
or U19359 (N_19359,N_18377,N_18617);
xor U19360 (N_19360,N_18631,N_19102);
nor U19361 (N_19361,N_19170,N_18571);
and U19362 (N_19362,N_19015,N_18938);
nor U19363 (N_19363,N_18601,N_19131);
nand U19364 (N_19364,N_18832,N_18517);
or U19365 (N_19365,N_19105,N_18735);
nand U19366 (N_19366,N_18973,N_18682);
nand U19367 (N_19367,N_19192,N_18148);
or U19368 (N_19368,N_18885,N_18062);
and U19369 (N_19369,N_18451,N_18200);
and U19370 (N_19370,N_19053,N_18186);
xnor U19371 (N_19371,N_18960,N_18716);
xor U19372 (N_19372,N_18752,N_18053);
or U19373 (N_19373,N_18482,N_18590);
or U19374 (N_19374,N_18473,N_18672);
xnor U19375 (N_19375,N_18411,N_19140);
nor U19376 (N_19376,N_18098,N_18203);
or U19377 (N_19377,N_18854,N_18146);
or U19378 (N_19378,N_18846,N_18892);
and U19379 (N_19379,N_18441,N_18722);
xor U19380 (N_19380,N_18404,N_18903);
nor U19381 (N_19381,N_18683,N_18463);
xnor U19382 (N_19382,N_19186,N_18619);
xor U19383 (N_19383,N_18802,N_18461);
or U19384 (N_19384,N_18699,N_19006);
xor U19385 (N_19385,N_18077,N_18530);
and U19386 (N_19386,N_18868,N_18750);
xnor U19387 (N_19387,N_18986,N_18248);
and U19388 (N_19388,N_18782,N_18114);
nor U19389 (N_19389,N_18193,N_18405);
and U19390 (N_19390,N_19110,N_18495);
nand U19391 (N_19391,N_18199,N_18084);
nand U19392 (N_19392,N_18609,N_18290);
and U19393 (N_19393,N_18851,N_18592);
xnor U19394 (N_19394,N_18720,N_19141);
xor U19395 (N_19395,N_18624,N_19194);
or U19396 (N_19396,N_18520,N_18815);
and U19397 (N_19397,N_18578,N_18616);
xnor U19398 (N_19398,N_18769,N_18877);
or U19399 (N_19399,N_18206,N_18825);
nand U19400 (N_19400,N_18671,N_18943);
nand U19401 (N_19401,N_19153,N_18416);
xnor U19402 (N_19402,N_18842,N_18566);
xnor U19403 (N_19403,N_18128,N_18635);
and U19404 (N_19404,N_18653,N_18418);
nand U19405 (N_19405,N_18040,N_18099);
xor U19406 (N_19406,N_18713,N_18956);
and U19407 (N_19407,N_18522,N_18994);
xnor U19408 (N_19408,N_18102,N_19109);
or U19409 (N_19409,N_19039,N_19033);
xor U19410 (N_19410,N_18880,N_19176);
nor U19411 (N_19411,N_18050,N_18845);
nand U19412 (N_19412,N_18545,N_18719);
nand U19413 (N_19413,N_18228,N_18518);
xnor U19414 (N_19414,N_18391,N_19132);
or U19415 (N_19415,N_18883,N_19012);
nand U19416 (N_19416,N_18584,N_18650);
or U19417 (N_19417,N_18468,N_18384);
nor U19418 (N_19418,N_19081,N_18122);
nor U19419 (N_19419,N_18641,N_18449);
or U19420 (N_19420,N_19061,N_18931);
xor U19421 (N_19421,N_19017,N_18264);
or U19422 (N_19422,N_18390,N_18983);
nand U19423 (N_19423,N_18302,N_18222);
nor U19424 (N_19424,N_18620,N_18496);
nor U19425 (N_19425,N_19076,N_18955);
nand U19426 (N_19426,N_18991,N_19184);
or U19427 (N_19427,N_18312,N_18987);
or U19428 (N_19428,N_18392,N_18486);
and U19429 (N_19429,N_18768,N_18734);
and U19430 (N_19430,N_18180,N_18019);
nor U19431 (N_19431,N_18059,N_18427);
or U19432 (N_19432,N_19001,N_19113);
and U19433 (N_19433,N_19040,N_18330);
nand U19434 (N_19434,N_18460,N_18737);
nand U19435 (N_19435,N_18929,N_18621);
and U19436 (N_19436,N_18176,N_18096);
or U19437 (N_19437,N_18039,N_18015);
or U19438 (N_19438,N_18063,N_18311);
and U19439 (N_19439,N_18125,N_18622);
nor U19440 (N_19440,N_18579,N_18353);
xnor U19441 (N_19441,N_18197,N_19115);
nor U19442 (N_19442,N_18689,N_18278);
nand U19443 (N_19443,N_18541,N_18744);
nor U19444 (N_19444,N_18728,N_19150);
xor U19445 (N_19445,N_18357,N_18004);
nor U19446 (N_19446,N_18663,N_18367);
xnor U19447 (N_19447,N_18602,N_18288);
and U19448 (N_19448,N_19181,N_18785);
or U19449 (N_19449,N_18263,N_19050);
nand U19450 (N_19450,N_18643,N_18408);
nand U19451 (N_19451,N_18189,N_18656);
and U19452 (N_19452,N_18613,N_18901);
nand U19453 (N_19453,N_18423,N_18001);
xnor U19454 (N_19454,N_18419,N_18606);
nand U19455 (N_19455,N_18853,N_18092);
xor U19456 (N_19456,N_19151,N_18373);
and U19457 (N_19457,N_18629,N_18154);
and U19458 (N_19458,N_18338,N_18487);
nor U19459 (N_19459,N_18213,N_18993);
xor U19460 (N_19460,N_18480,N_19018);
and U19461 (N_19461,N_18431,N_18086);
nand U19462 (N_19462,N_18303,N_18471);
nor U19463 (N_19463,N_18300,N_18131);
nand U19464 (N_19464,N_18394,N_18442);
or U19465 (N_19465,N_19152,N_18025);
xor U19466 (N_19466,N_18381,N_18761);
nand U19467 (N_19467,N_18610,N_18100);
nor U19468 (N_19468,N_18794,N_18751);
nor U19469 (N_19469,N_18847,N_18873);
and U19470 (N_19470,N_18034,N_19067);
or U19471 (N_19471,N_18863,N_18297);
nor U19472 (N_19472,N_18401,N_18022);
nor U19473 (N_19473,N_18558,N_18915);
nand U19474 (N_19474,N_19142,N_18150);
or U19475 (N_19475,N_18588,N_18133);
nand U19476 (N_19476,N_18654,N_18049);
xnor U19477 (N_19477,N_18603,N_18811);
xor U19478 (N_19478,N_18141,N_18575);
or U19479 (N_19479,N_18491,N_18065);
or U19480 (N_19480,N_19082,N_18255);
and U19481 (N_19481,N_19093,N_18018);
xor U19482 (N_19482,N_18927,N_18574);
or U19483 (N_19483,N_18524,N_18549);
nand U19484 (N_19484,N_18374,N_18573);
xor U19485 (N_19485,N_18267,N_18910);
or U19486 (N_19486,N_19096,N_19049);
and U19487 (N_19487,N_19187,N_18031);
nor U19488 (N_19488,N_18085,N_18223);
and U19489 (N_19489,N_18540,N_18754);
nand U19490 (N_19490,N_18792,N_18890);
nor U19491 (N_19491,N_18341,N_18326);
xnor U19492 (N_19492,N_19021,N_18398);
xnor U19493 (N_19493,N_19129,N_18536);
xnor U19494 (N_19494,N_18820,N_19146);
nor U19495 (N_19495,N_18366,N_18155);
or U19496 (N_19496,N_18923,N_18996);
and U19497 (N_19497,N_18694,N_18259);
and U19498 (N_19498,N_19101,N_18701);
nor U19499 (N_19499,N_19063,N_18772);
nor U19500 (N_19500,N_19144,N_18462);
nand U19501 (N_19501,N_19055,N_18111);
nor U19502 (N_19502,N_18333,N_18978);
nor U19503 (N_19503,N_19121,N_19145);
nor U19504 (N_19504,N_18979,N_18547);
or U19505 (N_19505,N_18589,N_19097);
xnor U19506 (N_19506,N_18529,N_18882);
or U19507 (N_19507,N_18599,N_18104);
nor U19508 (N_19508,N_18675,N_18475);
and U19509 (N_19509,N_19133,N_18012);
and U19510 (N_19510,N_18254,N_18107);
nand U19511 (N_19511,N_18434,N_19025);
nor U19512 (N_19512,N_18453,N_18321);
nand U19513 (N_19513,N_18778,N_18849);
nand U19514 (N_19514,N_18294,N_18337);
and U19515 (N_19515,N_19072,N_18410);
and U19516 (N_19516,N_18048,N_18593);
or U19517 (N_19517,N_18733,N_18543);
nand U19518 (N_19518,N_18075,N_18587);
nand U19519 (N_19519,N_18315,N_18972);
and U19520 (N_19520,N_18225,N_19019);
and U19521 (N_19521,N_18841,N_19173);
nand U19522 (N_19522,N_18681,N_18667);
nand U19523 (N_19523,N_18375,N_18679);
nand U19524 (N_19524,N_18334,N_18809);
and U19525 (N_19525,N_18604,N_18764);
or U19526 (N_19526,N_18899,N_18975);
nor U19527 (N_19527,N_18724,N_18605);
xnor U19528 (N_19528,N_18934,N_18512);
nor U19529 (N_19529,N_18661,N_19197);
xor U19530 (N_19530,N_18800,N_18655);
nor U19531 (N_19531,N_18669,N_18355);
nor U19532 (N_19532,N_18011,N_18008);
nand U19533 (N_19533,N_18340,N_19118);
and U19534 (N_19534,N_18450,N_18510);
xnor U19535 (N_19535,N_18396,N_18204);
and U19536 (N_19536,N_18014,N_18379);
nor U19537 (N_19537,N_18763,N_18893);
nor U19538 (N_19538,N_18271,N_18328);
xor U19539 (N_19539,N_18572,N_18550);
nand U19540 (N_19540,N_18795,N_18402);
nor U19541 (N_19541,N_18704,N_19030);
xor U19542 (N_19542,N_19024,N_18707);
or U19543 (N_19543,N_18274,N_18969);
xnor U19544 (N_19544,N_18157,N_18912);
nor U19545 (N_19545,N_18229,N_18708);
nor U19546 (N_19546,N_19008,N_18739);
or U19547 (N_19547,N_18933,N_18677);
or U19548 (N_19548,N_18083,N_18697);
nor U19549 (N_19549,N_18009,N_18499);
nand U19550 (N_19550,N_18607,N_18665);
nand U19551 (N_19551,N_18557,N_18581);
and U19552 (N_19552,N_18914,N_19175);
nand U19553 (N_19553,N_18535,N_18177);
nand U19554 (N_19554,N_18432,N_18185);
or U19555 (N_19555,N_18780,N_19079);
nand U19556 (N_19556,N_18134,N_18027);
and U19557 (N_19557,N_18030,N_18791);
nand U19558 (N_19558,N_18139,N_18103);
xnor U19559 (N_19559,N_18999,N_18064);
or U19560 (N_19560,N_18349,N_18095);
xor U19561 (N_19561,N_18252,N_18896);
nand U19562 (N_19562,N_18437,N_19091);
or U19563 (N_19563,N_18997,N_18505);
and U19564 (N_19564,N_18819,N_18774);
xnor U19565 (N_19565,N_18630,N_18940);
nor U19566 (N_19566,N_18198,N_18513);
xnor U19567 (N_19567,N_19180,N_18354);
or U19568 (N_19568,N_19185,N_18097);
xor U19569 (N_19569,N_18673,N_18647);
nor U19570 (N_19570,N_18013,N_18998);
nand U19571 (N_19571,N_18844,N_19154);
nand U19572 (N_19572,N_18968,N_19107);
xnor U19573 (N_19573,N_18320,N_18082);
or U19574 (N_19574,N_18478,N_18771);
or U19575 (N_19575,N_18784,N_18555);
nand U19576 (N_19576,N_18634,N_18803);
and U19577 (N_19577,N_18638,N_18980);
xor U19578 (N_19578,N_19163,N_18249);
nor U19579 (N_19579,N_18061,N_18429);
xnor U19580 (N_19580,N_18345,N_18074);
and U19581 (N_19581,N_18215,N_18138);
nor U19582 (N_19582,N_18121,N_18649);
nor U19583 (N_19583,N_18364,N_18182);
or U19584 (N_19584,N_19137,N_18755);
and U19585 (N_19585,N_18257,N_18488);
and U19586 (N_19586,N_18214,N_18151);
and U19587 (N_19587,N_18370,N_18691);
nor U19588 (N_19588,N_18692,N_18789);
nand U19589 (N_19589,N_18648,N_18950);
nand U19590 (N_19590,N_18397,N_18066);
or U19591 (N_19591,N_18173,N_18051);
nor U19592 (N_19592,N_18962,N_18280);
and U19593 (N_19593,N_18369,N_18258);
and U19594 (N_19594,N_18360,N_18289);
nor U19595 (N_19595,N_18021,N_18430);
nor U19596 (N_19596,N_18120,N_18209);
xor U19597 (N_19597,N_18515,N_18042);
and U19598 (N_19598,N_19147,N_18244);
and U19599 (N_19599,N_19155,N_19126);
or U19600 (N_19600,N_18870,N_18732);
and U19601 (N_19601,N_18818,N_18952);
xnor U19602 (N_19602,N_18788,N_19052);
and U19603 (N_19603,N_18498,N_19138);
nand U19604 (N_19604,N_18452,N_18835);
or U19605 (N_19605,N_18067,N_18448);
or U19606 (N_19606,N_18167,N_18399);
or U19607 (N_19607,N_18343,N_18422);
and U19608 (N_19608,N_18570,N_19085);
nand U19609 (N_19609,N_18417,N_19048);
xnor U19610 (N_19610,N_18887,N_18023);
nor U19611 (N_19611,N_18238,N_18614);
xor U19612 (N_19612,N_18838,N_18586);
or U19613 (N_19613,N_18160,N_18848);
or U19614 (N_19614,N_18712,N_18046);
nor U19615 (N_19615,N_18594,N_18232);
and U19616 (N_19616,N_18045,N_18805);
xnor U19617 (N_19617,N_18696,N_19026);
or U19618 (N_19618,N_18628,N_18779);
xor U19619 (N_19619,N_18319,N_19165);
or U19620 (N_19620,N_18310,N_19190);
and U19621 (N_19621,N_18525,N_18383);
nand U19622 (N_19622,N_19124,N_18862);
xnor U19623 (N_19623,N_19056,N_18400);
nand U19624 (N_19624,N_18306,N_18860);
and U19625 (N_19625,N_18678,N_18967);
and U19626 (N_19626,N_18226,N_18703);
and U19627 (N_19627,N_18886,N_18472);
xor U19628 (N_19628,N_18982,N_18560);
xnor U19629 (N_19629,N_18900,N_18124);
xnor U19630 (N_19630,N_18810,N_18469);
nand U19631 (N_19631,N_19020,N_18726);
nor U19632 (N_19632,N_18029,N_18514);
or U19633 (N_19633,N_18984,N_18680);
nand U19634 (N_19634,N_18781,N_18403);
nor U19635 (N_19635,N_19011,N_18171);
and U19636 (N_19636,N_18644,N_18830);
xor U19637 (N_19637,N_18455,N_18236);
nand U19638 (N_19638,N_19090,N_19168);
nor U19639 (N_19639,N_18947,N_18657);
and U19640 (N_19640,N_18413,N_18301);
and U19641 (N_19641,N_18164,N_18129);
and U19642 (N_19642,N_18211,N_18037);
nor U19643 (N_19643,N_18908,N_18618);
xor U19644 (N_19644,N_18843,N_18088);
xor U19645 (N_19645,N_18503,N_18725);
and U19646 (N_19646,N_18108,N_19054);
or U19647 (N_19647,N_18163,N_18352);
and U19648 (N_19648,N_18395,N_18729);
or U19649 (N_19649,N_18762,N_18143);
nand U19650 (N_19650,N_18477,N_18559);
or U19651 (N_19651,N_18827,N_19130);
and U19652 (N_19652,N_18816,N_18507);
and U19653 (N_19653,N_18016,N_18327);
and U19654 (N_19654,N_18528,N_18208);
and U19655 (N_19655,N_19086,N_18556);
xnor U19656 (N_19656,N_18342,N_18458);
nor U19657 (N_19657,N_18688,N_18740);
and U19658 (N_19658,N_18822,N_19188);
xor U19659 (N_19659,N_18727,N_18483);
nand U19660 (N_19660,N_19134,N_18767);
nor U19661 (N_19661,N_18295,N_18010);
nor U19662 (N_19662,N_18433,N_19114);
and U19663 (N_19663,N_18537,N_18765);
and U19664 (N_19664,N_18115,N_18804);
or U19665 (N_19665,N_18305,N_18233);
or U19666 (N_19666,N_18272,N_18147);
and U19667 (N_19667,N_19074,N_18709);
xor U19668 (N_19668,N_18474,N_18093);
xor U19669 (N_19669,N_18920,N_18116);
nand U19670 (N_19670,N_18484,N_18850);
xor U19671 (N_19671,N_18365,N_18336);
nand U19672 (N_19672,N_18783,N_18597);
and U19673 (N_19673,N_18662,N_18425);
nor U19674 (N_19674,N_18718,N_18407);
and U19675 (N_19675,N_18839,N_18971);
xnor U19676 (N_19676,N_18005,N_18869);
nand U19677 (N_19677,N_18479,N_18456);
nor U19678 (N_19678,N_18443,N_19162);
nor U19679 (N_19679,N_18611,N_19189);
nand U19680 (N_19680,N_18283,N_18906);
xor U19681 (N_19681,N_18090,N_18135);
nand U19682 (N_19682,N_19136,N_18916);
xor U19683 (N_19683,N_18118,N_18511);
and U19684 (N_19684,N_18928,N_18775);
xor U19685 (N_19685,N_18961,N_18985);
nand U19686 (N_19686,N_18057,N_18814);
or U19687 (N_19687,N_18612,N_18224);
nor U19688 (N_19688,N_18376,N_19164);
and U19689 (N_19689,N_18829,N_18904);
xor U19690 (N_19690,N_18898,N_18412);
xor U19691 (N_19691,N_18858,N_18888);
nor U19692 (N_19692,N_18196,N_18192);
and U19693 (N_19693,N_18260,N_18036);
or U19694 (N_19694,N_18909,N_19177);
nand U19695 (N_19695,N_18127,N_18548);
nor U19696 (N_19696,N_18565,N_18119);
nand U19697 (N_19697,N_18786,N_18256);
xnor U19698 (N_19698,N_18757,N_18250);
or U19699 (N_19699,N_18126,N_18246);
xnor U19700 (N_19700,N_18265,N_18438);
or U19701 (N_19701,N_18335,N_18465);
xnor U19702 (N_19702,N_18132,N_18658);
or U19703 (N_19703,N_18174,N_18299);
nand U19704 (N_19704,N_18492,N_18936);
and U19705 (N_19705,N_18958,N_19196);
nor U19706 (N_19706,N_18506,N_18113);
and U19707 (N_19707,N_18623,N_19171);
and U19708 (N_19708,N_18038,N_18339);
nand U19709 (N_19709,N_19043,N_19158);
xnor U19710 (N_19710,N_18871,N_18798);
and U19711 (N_19711,N_18406,N_18481);
nor U19712 (N_19712,N_18332,N_18717);
or U19713 (N_19713,N_18932,N_18897);
nor U19714 (N_19714,N_19088,N_18596);
and U19715 (N_19715,N_18470,N_18874);
xnor U19716 (N_19716,N_18824,N_19022);
nor U19717 (N_19717,N_19098,N_18230);
nand U19718 (N_19718,N_18188,N_18318);
nor U19719 (N_19719,N_18281,N_19066);
nor U19720 (N_19720,N_18421,N_18161);
xor U19721 (N_19721,N_19031,N_18414);
or U19722 (N_19722,N_18698,N_18277);
or U19723 (N_19723,N_18105,N_18168);
and U19724 (N_19724,N_18194,N_18591);
xnor U19725 (N_19725,N_18502,N_18995);
xnor U19726 (N_19726,N_18812,N_19117);
and U19727 (N_19727,N_19149,N_18072);
nand U19728 (N_19728,N_18382,N_18913);
xnor U19729 (N_19729,N_19062,N_18730);
nor U19730 (N_19730,N_18459,N_19092);
xor U19731 (N_19731,N_19064,N_18287);
nand U19732 (N_19732,N_18024,N_18926);
and U19733 (N_19733,N_18954,N_18583);
nor U19734 (N_19734,N_18220,N_18645);
or U19735 (N_19735,N_18964,N_19127);
nor U19736 (N_19736,N_18415,N_18136);
or U19737 (N_19737,N_19058,N_18227);
or U19738 (N_19738,N_18538,N_18840);
nor U19739 (N_19739,N_19195,N_18693);
nor U19740 (N_19740,N_18942,N_18218);
nand U19741 (N_19741,N_18179,N_19073);
nor U19742 (N_19742,N_18282,N_18202);
xor U19743 (N_19743,N_18930,N_18444);
nor U19744 (N_19744,N_18094,N_19034);
nand U19745 (N_19745,N_18519,N_18165);
or U19746 (N_19746,N_19095,N_18457);
and U19747 (N_19747,N_18216,N_18156);
nor U19748 (N_19748,N_18358,N_18945);
or U19749 (N_19749,N_18598,N_19057);
nor U19750 (N_19750,N_18056,N_18516);
nor U19751 (N_19751,N_18166,N_19075);
xnor U19752 (N_19752,N_19116,N_18615);
or U19753 (N_19753,N_18876,N_18070);
nor U19754 (N_19754,N_18239,N_18988);
nor U19755 (N_19755,N_18859,N_18435);
xnor U19756 (N_19756,N_18576,N_18959);
xor U19757 (N_19757,N_18309,N_18902);
xnor U19758 (N_19758,N_19023,N_18266);
xnor U19759 (N_19759,N_18017,N_18695);
and U19760 (N_19760,N_18316,N_18924);
and U19761 (N_19761,N_18331,N_18664);
nor U19762 (N_19762,N_18047,N_18799);
nor U19763 (N_19763,N_18577,N_18081);
and U19764 (N_19764,N_18242,N_18170);
and U19765 (N_19765,N_18561,N_18922);
nand U19766 (N_19766,N_18270,N_18895);
or U19767 (N_19767,N_18076,N_18069);
or U19768 (N_19768,N_18508,N_18253);
xor U19769 (N_19769,N_18169,N_18439);
xnor U19770 (N_19770,N_18002,N_18608);
nor U19771 (N_19771,N_18275,N_18966);
nor U19772 (N_19772,N_18813,N_18231);
and U19773 (N_19773,N_19002,N_18639);
nor U19774 (N_19774,N_18079,N_18760);
or U19775 (N_19775,N_18879,N_18112);
xnor U19776 (N_19776,N_18534,N_19005);
nand U19777 (N_19777,N_18881,N_18314);
nand U19778 (N_19778,N_18142,N_19044);
nor U19779 (N_19779,N_18944,N_19198);
or U19780 (N_19780,N_18632,N_18872);
or U19781 (N_19781,N_18221,N_18003);
or U19782 (N_19782,N_18020,N_18741);
xor U19783 (N_19783,N_19157,N_18123);
xnor U19784 (N_19784,N_18497,N_18965);
nor U19785 (N_19785,N_18158,N_18626);
nor U19786 (N_19786,N_18974,N_18917);
nand U19787 (N_19787,N_19111,N_18833);
or U19788 (N_19788,N_18552,N_19094);
and U19789 (N_19789,N_18731,N_18313);
nand U19790 (N_19790,N_18939,N_19174);
nor U19791 (N_19791,N_18745,N_18527);
or U19792 (N_19792,N_18884,N_18217);
and U19793 (N_19793,N_19007,N_18705);
xor U19794 (N_19794,N_18676,N_18894);
nand U19795 (N_19795,N_19122,N_19004);
and U19796 (N_19796,N_18035,N_18346);
nand U19797 (N_19797,N_19193,N_18646);
nand U19798 (N_19798,N_19089,N_18659);
xor U19799 (N_19799,N_18836,N_18808);
or U19800 (N_19800,N_19104,N_18641);
xnor U19801 (N_19801,N_18260,N_18966);
and U19802 (N_19802,N_18267,N_18294);
nand U19803 (N_19803,N_18059,N_18018);
nand U19804 (N_19804,N_18389,N_18136);
and U19805 (N_19805,N_18434,N_19175);
or U19806 (N_19806,N_18293,N_18298);
or U19807 (N_19807,N_19141,N_18277);
or U19808 (N_19808,N_19024,N_18391);
or U19809 (N_19809,N_18651,N_18444);
xor U19810 (N_19810,N_19148,N_19023);
nand U19811 (N_19811,N_18829,N_18050);
xor U19812 (N_19812,N_18213,N_18064);
and U19813 (N_19813,N_18495,N_18369);
nor U19814 (N_19814,N_18303,N_18159);
nor U19815 (N_19815,N_18063,N_18514);
nor U19816 (N_19816,N_18011,N_19113);
nand U19817 (N_19817,N_18630,N_18872);
xnor U19818 (N_19818,N_19184,N_18828);
nor U19819 (N_19819,N_18019,N_18093);
or U19820 (N_19820,N_18268,N_18389);
and U19821 (N_19821,N_18459,N_18739);
nand U19822 (N_19822,N_18374,N_18137);
nor U19823 (N_19823,N_19148,N_18346);
nand U19824 (N_19824,N_18022,N_18670);
nor U19825 (N_19825,N_18710,N_18987);
nand U19826 (N_19826,N_18692,N_18002);
nor U19827 (N_19827,N_18139,N_19056);
nor U19828 (N_19828,N_19033,N_18252);
and U19829 (N_19829,N_18093,N_18251);
nor U19830 (N_19830,N_18883,N_18716);
or U19831 (N_19831,N_18316,N_18953);
and U19832 (N_19832,N_18247,N_18419);
nand U19833 (N_19833,N_19110,N_19012);
nand U19834 (N_19834,N_18120,N_18548);
nand U19835 (N_19835,N_18202,N_18064);
or U19836 (N_19836,N_19026,N_18344);
xor U19837 (N_19837,N_18701,N_18481);
and U19838 (N_19838,N_18186,N_18303);
xnor U19839 (N_19839,N_18203,N_18286);
or U19840 (N_19840,N_18813,N_18499);
nand U19841 (N_19841,N_18421,N_18837);
nor U19842 (N_19842,N_18773,N_19143);
nand U19843 (N_19843,N_18712,N_18449);
nor U19844 (N_19844,N_18485,N_18948);
and U19845 (N_19845,N_18582,N_19037);
nand U19846 (N_19846,N_18637,N_18512);
nand U19847 (N_19847,N_18061,N_19003);
xor U19848 (N_19848,N_18274,N_18688);
and U19849 (N_19849,N_18487,N_18455);
nor U19850 (N_19850,N_18356,N_19157);
and U19851 (N_19851,N_19059,N_18533);
xnor U19852 (N_19852,N_18778,N_18954);
xor U19853 (N_19853,N_18740,N_19092);
nor U19854 (N_19854,N_19064,N_18007);
nor U19855 (N_19855,N_18469,N_18930);
xor U19856 (N_19856,N_18887,N_18383);
and U19857 (N_19857,N_18181,N_19160);
and U19858 (N_19858,N_19003,N_18443);
nand U19859 (N_19859,N_18187,N_18166);
nor U19860 (N_19860,N_18977,N_18870);
xnor U19861 (N_19861,N_18627,N_18512);
xor U19862 (N_19862,N_18233,N_18610);
or U19863 (N_19863,N_18832,N_18977);
and U19864 (N_19864,N_18085,N_18504);
and U19865 (N_19865,N_18540,N_18156);
and U19866 (N_19866,N_19010,N_19112);
and U19867 (N_19867,N_18775,N_19106);
xnor U19868 (N_19868,N_18183,N_18312);
nand U19869 (N_19869,N_18969,N_18818);
nor U19870 (N_19870,N_18758,N_18785);
nor U19871 (N_19871,N_18531,N_18018);
or U19872 (N_19872,N_18211,N_18803);
or U19873 (N_19873,N_18238,N_18654);
xnor U19874 (N_19874,N_18648,N_18135);
or U19875 (N_19875,N_18068,N_19143);
and U19876 (N_19876,N_18782,N_18343);
or U19877 (N_19877,N_18532,N_18380);
or U19878 (N_19878,N_19121,N_19067);
nand U19879 (N_19879,N_18196,N_18655);
nand U19880 (N_19880,N_18253,N_18069);
or U19881 (N_19881,N_19129,N_18546);
nor U19882 (N_19882,N_19091,N_18754);
or U19883 (N_19883,N_19026,N_18362);
nand U19884 (N_19884,N_18142,N_19108);
nor U19885 (N_19885,N_18338,N_18388);
or U19886 (N_19886,N_19040,N_18923);
xor U19887 (N_19887,N_19001,N_18058);
and U19888 (N_19888,N_18857,N_18958);
nor U19889 (N_19889,N_18560,N_18672);
and U19890 (N_19890,N_18683,N_18296);
or U19891 (N_19891,N_18456,N_18641);
nor U19892 (N_19892,N_18442,N_18050);
xnor U19893 (N_19893,N_18509,N_18298);
nor U19894 (N_19894,N_18049,N_18688);
or U19895 (N_19895,N_18054,N_18302);
xnor U19896 (N_19896,N_18885,N_18227);
xor U19897 (N_19897,N_18841,N_19106);
xor U19898 (N_19898,N_18457,N_18942);
or U19899 (N_19899,N_18653,N_18677);
and U19900 (N_19900,N_18688,N_18988);
and U19901 (N_19901,N_18318,N_18975);
xor U19902 (N_19902,N_18737,N_18959);
xnor U19903 (N_19903,N_18689,N_18647);
nor U19904 (N_19904,N_18245,N_18064);
and U19905 (N_19905,N_18155,N_18589);
or U19906 (N_19906,N_18565,N_18741);
xnor U19907 (N_19907,N_18453,N_18815);
and U19908 (N_19908,N_18471,N_18830);
xnor U19909 (N_19909,N_18885,N_18728);
and U19910 (N_19910,N_18231,N_18173);
and U19911 (N_19911,N_18940,N_18612);
nor U19912 (N_19912,N_18198,N_19180);
xnor U19913 (N_19913,N_18538,N_18317);
nor U19914 (N_19914,N_18245,N_18382);
nand U19915 (N_19915,N_18744,N_19126);
and U19916 (N_19916,N_18774,N_19008);
and U19917 (N_19917,N_18021,N_19120);
nor U19918 (N_19918,N_18937,N_18082);
and U19919 (N_19919,N_18820,N_18246);
nand U19920 (N_19920,N_18480,N_19038);
and U19921 (N_19921,N_18891,N_19154);
nand U19922 (N_19922,N_18783,N_18364);
xor U19923 (N_19923,N_18241,N_18798);
nand U19924 (N_19924,N_18821,N_18369);
or U19925 (N_19925,N_18791,N_18787);
and U19926 (N_19926,N_19170,N_18209);
and U19927 (N_19927,N_18915,N_18312);
nand U19928 (N_19928,N_19155,N_18424);
and U19929 (N_19929,N_18377,N_18108);
nand U19930 (N_19930,N_18511,N_18137);
xnor U19931 (N_19931,N_19199,N_18569);
nand U19932 (N_19932,N_18006,N_19181);
and U19933 (N_19933,N_18602,N_19047);
or U19934 (N_19934,N_18833,N_19188);
or U19935 (N_19935,N_18492,N_19086);
and U19936 (N_19936,N_18419,N_18218);
nand U19937 (N_19937,N_18894,N_19080);
nand U19938 (N_19938,N_18585,N_18064);
xnor U19939 (N_19939,N_18036,N_18577);
and U19940 (N_19940,N_18952,N_19041);
xor U19941 (N_19941,N_19144,N_19080);
or U19942 (N_19942,N_18903,N_18559);
nor U19943 (N_19943,N_18091,N_18082);
nor U19944 (N_19944,N_18411,N_18585);
nand U19945 (N_19945,N_18013,N_18312);
xnor U19946 (N_19946,N_19162,N_18205);
xor U19947 (N_19947,N_18938,N_18373);
nand U19948 (N_19948,N_18294,N_18042);
xnor U19949 (N_19949,N_18590,N_18170);
nor U19950 (N_19950,N_18380,N_18715);
and U19951 (N_19951,N_18741,N_18171);
nor U19952 (N_19952,N_18721,N_18016);
xnor U19953 (N_19953,N_18096,N_18539);
and U19954 (N_19954,N_18796,N_18371);
nor U19955 (N_19955,N_18209,N_18980);
and U19956 (N_19956,N_18739,N_18723);
nor U19957 (N_19957,N_19054,N_18045);
or U19958 (N_19958,N_18157,N_18777);
and U19959 (N_19959,N_18130,N_18469);
nor U19960 (N_19960,N_18334,N_18548);
or U19961 (N_19961,N_18777,N_18384);
and U19962 (N_19962,N_18515,N_18914);
and U19963 (N_19963,N_18263,N_19013);
or U19964 (N_19964,N_18518,N_19162);
nand U19965 (N_19965,N_18347,N_18252);
xor U19966 (N_19966,N_18975,N_18419);
and U19967 (N_19967,N_19093,N_18159);
or U19968 (N_19968,N_18344,N_18715);
nor U19969 (N_19969,N_18907,N_19028);
xor U19970 (N_19970,N_18284,N_18191);
and U19971 (N_19971,N_18186,N_18865);
and U19972 (N_19972,N_18664,N_18989);
or U19973 (N_19973,N_18192,N_18839);
xnor U19974 (N_19974,N_18667,N_18724);
or U19975 (N_19975,N_18270,N_18928);
xnor U19976 (N_19976,N_18334,N_18423);
or U19977 (N_19977,N_18895,N_18999);
nor U19978 (N_19978,N_18968,N_18920);
xnor U19979 (N_19979,N_18182,N_19172);
and U19980 (N_19980,N_18027,N_18453);
or U19981 (N_19981,N_18505,N_18199);
nand U19982 (N_19982,N_18920,N_18222);
and U19983 (N_19983,N_18120,N_18861);
or U19984 (N_19984,N_18317,N_18986);
nand U19985 (N_19985,N_19089,N_18244);
nand U19986 (N_19986,N_18620,N_18789);
and U19987 (N_19987,N_18857,N_18147);
nor U19988 (N_19988,N_19016,N_18576);
nand U19989 (N_19989,N_18052,N_18919);
xor U19990 (N_19990,N_19096,N_18490);
xnor U19991 (N_19991,N_19151,N_18506);
nand U19992 (N_19992,N_18494,N_19069);
nand U19993 (N_19993,N_19198,N_18211);
and U19994 (N_19994,N_19070,N_18716);
xor U19995 (N_19995,N_19009,N_18653);
and U19996 (N_19996,N_18835,N_18265);
xnor U19997 (N_19997,N_18571,N_18568);
nor U19998 (N_19998,N_18542,N_18371);
or U19999 (N_19999,N_18355,N_18918);
or U20000 (N_20000,N_18799,N_19051);
xnor U20001 (N_20001,N_18705,N_18866);
and U20002 (N_20002,N_18849,N_18131);
or U20003 (N_20003,N_18466,N_18279);
nand U20004 (N_20004,N_18467,N_18687);
xnor U20005 (N_20005,N_18279,N_18958);
nor U20006 (N_20006,N_19153,N_18751);
xor U20007 (N_20007,N_18297,N_18312);
nor U20008 (N_20008,N_18319,N_18603);
nand U20009 (N_20009,N_18406,N_18649);
nand U20010 (N_20010,N_19074,N_18138);
and U20011 (N_20011,N_19050,N_18929);
and U20012 (N_20012,N_18201,N_18451);
nand U20013 (N_20013,N_18556,N_18992);
nor U20014 (N_20014,N_18680,N_19133);
nand U20015 (N_20015,N_18613,N_18263);
or U20016 (N_20016,N_18625,N_18174);
xor U20017 (N_20017,N_18143,N_18531);
nand U20018 (N_20018,N_18306,N_18708);
xor U20019 (N_20019,N_18550,N_18848);
and U20020 (N_20020,N_18796,N_18735);
xnor U20021 (N_20021,N_18094,N_18305);
and U20022 (N_20022,N_18377,N_18567);
and U20023 (N_20023,N_18180,N_18435);
nor U20024 (N_20024,N_19169,N_19117);
nor U20025 (N_20025,N_18025,N_18073);
xnor U20026 (N_20026,N_19174,N_18705);
nor U20027 (N_20027,N_18433,N_18336);
or U20028 (N_20028,N_18961,N_18296);
xnor U20029 (N_20029,N_19092,N_18431);
xnor U20030 (N_20030,N_18667,N_18379);
xor U20031 (N_20031,N_18250,N_18663);
nand U20032 (N_20032,N_18047,N_18927);
or U20033 (N_20033,N_18594,N_19045);
or U20034 (N_20034,N_18259,N_19130);
or U20035 (N_20035,N_18091,N_19074);
or U20036 (N_20036,N_19080,N_18882);
and U20037 (N_20037,N_18168,N_18028);
xnor U20038 (N_20038,N_18007,N_18186);
and U20039 (N_20039,N_18371,N_18640);
and U20040 (N_20040,N_18298,N_18765);
xnor U20041 (N_20041,N_18594,N_18905);
and U20042 (N_20042,N_18756,N_18912);
and U20043 (N_20043,N_18605,N_18488);
and U20044 (N_20044,N_19138,N_18147);
and U20045 (N_20045,N_18830,N_18278);
nand U20046 (N_20046,N_18646,N_19055);
and U20047 (N_20047,N_18215,N_18471);
or U20048 (N_20048,N_18609,N_18558);
or U20049 (N_20049,N_18446,N_18580);
or U20050 (N_20050,N_18687,N_18078);
or U20051 (N_20051,N_18613,N_18704);
or U20052 (N_20052,N_18371,N_18604);
nand U20053 (N_20053,N_18707,N_18477);
xor U20054 (N_20054,N_18008,N_18864);
nor U20055 (N_20055,N_18494,N_18421);
nand U20056 (N_20056,N_19155,N_18309);
and U20057 (N_20057,N_18984,N_18223);
nand U20058 (N_20058,N_18625,N_18871);
nor U20059 (N_20059,N_18131,N_18714);
or U20060 (N_20060,N_18838,N_18105);
or U20061 (N_20061,N_18188,N_18863);
nand U20062 (N_20062,N_18446,N_18776);
xor U20063 (N_20063,N_18581,N_18896);
and U20064 (N_20064,N_18072,N_18050);
nand U20065 (N_20065,N_19199,N_18124);
and U20066 (N_20066,N_18131,N_19010);
and U20067 (N_20067,N_18404,N_19086);
or U20068 (N_20068,N_19047,N_18993);
xnor U20069 (N_20069,N_18367,N_18412);
nor U20070 (N_20070,N_18589,N_18085);
and U20071 (N_20071,N_19085,N_18531);
nor U20072 (N_20072,N_18504,N_19090);
and U20073 (N_20073,N_19199,N_18452);
nand U20074 (N_20074,N_19023,N_18798);
xnor U20075 (N_20075,N_19088,N_18009);
nand U20076 (N_20076,N_18621,N_18521);
or U20077 (N_20077,N_18061,N_19094);
nand U20078 (N_20078,N_18886,N_18161);
and U20079 (N_20079,N_18187,N_18819);
nor U20080 (N_20080,N_18999,N_19179);
nand U20081 (N_20081,N_19001,N_18690);
nor U20082 (N_20082,N_18821,N_18768);
xor U20083 (N_20083,N_18040,N_18383);
and U20084 (N_20084,N_18370,N_18597);
xor U20085 (N_20085,N_18847,N_19065);
and U20086 (N_20086,N_19091,N_18941);
nor U20087 (N_20087,N_18271,N_18497);
and U20088 (N_20088,N_18690,N_18003);
or U20089 (N_20089,N_19163,N_18981);
xor U20090 (N_20090,N_18032,N_18876);
xor U20091 (N_20091,N_18510,N_18039);
xnor U20092 (N_20092,N_18590,N_18576);
nand U20093 (N_20093,N_18498,N_18790);
nor U20094 (N_20094,N_19171,N_18987);
nor U20095 (N_20095,N_18119,N_18826);
and U20096 (N_20096,N_19000,N_18364);
xor U20097 (N_20097,N_18502,N_19070);
and U20098 (N_20098,N_18264,N_18240);
and U20099 (N_20099,N_18937,N_18605);
xnor U20100 (N_20100,N_18709,N_18954);
nor U20101 (N_20101,N_18424,N_18917);
xor U20102 (N_20102,N_19017,N_18332);
and U20103 (N_20103,N_18537,N_18138);
or U20104 (N_20104,N_18206,N_18048);
nor U20105 (N_20105,N_18233,N_18633);
xnor U20106 (N_20106,N_18982,N_18521);
nor U20107 (N_20107,N_18959,N_19146);
nand U20108 (N_20108,N_18477,N_18724);
xnor U20109 (N_20109,N_18458,N_18388);
nand U20110 (N_20110,N_18201,N_19008);
and U20111 (N_20111,N_18533,N_18484);
xnor U20112 (N_20112,N_18553,N_19189);
nor U20113 (N_20113,N_18012,N_18067);
nor U20114 (N_20114,N_18964,N_18524);
nor U20115 (N_20115,N_18469,N_18187);
nand U20116 (N_20116,N_18187,N_18860);
xor U20117 (N_20117,N_18939,N_18278);
nand U20118 (N_20118,N_18056,N_18566);
xor U20119 (N_20119,N_18587,N_18447);
and U20120 (N_20120,N_18251,N_18879);
nor U20121 (N_20121,N_18775,N_18836);
xor U20122 (N_20122,N_18337,N_18795);
and U20123 (N_20123,N_18800,N_19058);
or U20124 (N_20124,N_18712,N_18107);
and U20125 (N_20125,N_18135,N_18781);
nand U20126 (N_20126,N_18899,N_18252);
xnor U20127 (N_20127,N_18375,N_18865);
nor U20128 (N_20128,N_18871,N_18531);
nand U20129 (N_20129,N_18516,N_18897);
nor U20130 (N_20130,N_18850,N_18359);
nor U20131 (N_20131,N_19141,N_18689);
xor U20132 (N_20132,N_18387,N_18658);
or U20133 (N_20133,N_18447,N_18079);
nand U20134 (N_20134,N_18502,N_18264);
or U20135 (N_20135,N_18413,N_18667);
xnor U20136 (N_20136,N_18124,N_18508);
xnor U20137 (N_20137,N_18485,N_18271);
and U20138 (N_20138,N_19078,N_18977);
nand U20139 (N_20139,N_18960,N_18390);
or U20140 (N_20140,N_18247,N_19067);
and U20141 (N_20141,N_18103,N_18630);
or U20142 (N_20142,N_18188,N_18041);
xor U20143 (N_20143,N_18618,N_19157);
xor U20144 (N_20144,N_18665,N_18774);
nor U20145 (N_20145,N_18135,N_18946);
nor U20146 (N_20146,N_18567,N_18004);
or U20147 (N_20147,N_18575,N_18564);
nand U20148 (N_20148,N_19080,N_18173);
and U20149 (N_20149,N_18415,N_18539);
or U20150 (N_20150,N_18908,N_19167);
xnor U20151 (N_20151,N_18703,N_18517);
and U20152 (N_20152,N_18800,N_19059);
nor U20153 (N_20153,N_19076,N_18431);
nand U20154 (N_20154,N_18162,N_19104);
xnor U20155 (N_20155,N_18626,N_18358);
and U20156 (N_20156,N_18705,N_19134);
nor U20157 (N_20157,N_19032,N_18030);
nor U20158 (N_20158,N_18171,N_18920);
xnor U20159 (N_20159,N_18629,N_18704);
or U20160 (N_20160,N_18431,N_18851);
or U20161 (N_20161,N_18105,N_18868);
xor U20162 (N_20162,N_18860,N_18178);
xor U20163 (N_20163,N_18078,N_18523);
xor U20164 (N_20164,N_18158,N_18714);
nor U20165 (N_20165,N_18667,N_18283);
and U20166 (N_20166,N_19129,N_18543);
nor U20167 (N_20167,N_18233,N_18811);
nor U20168 (N_20168,N_18025,N_18956);
or U20169 (N_20169,N_19136,N_18778);
xnor U20170 (N_20170,N_18430,N_18304);
xor U20171 (N_20171,N_18558,N_18153);
or U20172 (N_20172,N_18338,N_18838);
nand U20173 (N_20173,N_18851,N_19049);
nor U20174 (N_20174,N_18124,N_18819);
nand U20175 (N_20175,N_18649,N_18859);
nor U20176 (N_20176,N_18428,N_18783);
xor U20177 (N_20177,N_18258,N_19033);
and U20178 (N_20178,N_18760,N_18023);
and U20179 (N_20179,N_19070,N_18138);
xor U20180 (N_20180,N_18067,N_18799);
xor U20181 (N_20181,N_18379,N_18491);
or U20182 (N_20182,N_18586,N_18170);
xor U20183 (N_20183,N_18545,N_18710);
and U20184 (N_20184,N_18936,N_18486);
nand U20185 (N_20185,N_18814,N_18046);
nand U20186 (N_20186,N_19175,N_18068);
and U20187 (N_20187,N_18232,N_18507);
nand U20188 (N_20188,N_18201,N_18517);
and U20189 (N_20189,N_18133,N_19101);
or U20190 (N_20190,N_18378,N_18989);
xnor U20191 (N_20191,N_19175,N_18335);
and U20192 (N_20192,N_19057,N_18145);
nor U20193 (N_20193,N_18958,N_18375);
and U20194 (N_20194,N_19079,N_18651);
or U20195 (N_20195,N_18463,N_18187);
xnor U20196 (N_20196,N_18607,N_18531);
nor U20197 (N_20197,N_18674,N_19070);
nand U20198 (N_20198,N_18545,N_18028);
or U20199 (N_20199,N_19033,N_18476);
xnor U20200 (N_20200,N_18897,N_18922);
xor U20201 (N_20201,N_19037,N_18766);
xor U20202 (N_20202,N_18266,N_18224);
nand U20203 (N_20203,N_18640,N_18136);
nand U20204 (N_20204,N_18643,N_18456);
nor U20205 (N_20205,N_19134,N_18682);
xnor U20206 (N_20206,N_18498,N_18431);
or U20207 (N_20207,N_18270,N_18346);
or U20208 (N_20208,N_18846,N_19192);
or U20209 (N_20209,N_18899,N_18375);
or U20210 (N_20210,N_18174,N_18866);
nor U20211 (N_20211,N_19170,N_18689);
nand U20212 (N_20212,N_18339,N_19131);
or U20213 (N_20213,N_18523,N_18896);
xnor U20214 (N_20214,N_18838,N_18470);
nand U20215 (N_20215,N_19112,N_18859);
nor U20216 (N_20216,N_18445,N_18810);
nor U20217 (N_20217,N_18103,N_18216);
nor U20218 (N_20218,N_19113,N_19141);
or U20219 (N_20219,N_18654,N_18461);
nand U20220 (N_20220,N_18723,N_18614);
or U20221 (N_20221,N_18127,N_19152);
nand U20222 (N_20222,N_18204,N_18389);
or U20223 (N_20223,N_18056,N_18382);
or U20224 (N_20224,N_18418,N_19168);
or U20225 (N_20225,N_18176,N_18235);
nor U20226 (N_20226,N_18042,N_18056);
nand U20227 (N_20227,N_18143,N_18701);
or U20228 (N_20228,N_18356,N_18825);
and U20229 (N_20229,N_18747,N_18834);
or U20230 (N_20230,N_18981,N_18073);
nor U20231 (N_20231,N_18881,N_18153);
nand U20232 (N_20232,N_18234,N_18735);
xor U20233 (N_20233,N_18170,N_18427);
xnor U20234 (N_20234,N_18411,N_18595);
and U20235 (N_20235,N_18617,N_18212);
xnor U20236 (N_20236,N_18337,N_18537);
xor U20237 (N_20237,N_18644,N_18827);
xnor U20238 (N_20238,N_18021,N_18728);
or U20239 (N_20239,N_18911,N_18500);
nand U20240 (N_20240,N_18934,N_18101);
or U20241 (N_20241,N_18383,N_18695);
or U20242 (N_20242,N_18316,N_18403);
or U20243 (N_20243,N_18958,N_18294);
nor U20244 (N_20244,N_18932,N_18310);
nand U20245 (N_20245,N_18264,N_18587);
nand U20246 (N_20246,N_18626,N_18595);
and U20247 (N_20247,N_18017,N_18971);
or U20248 (N_20248,N_18060,N_19112);
or U20249 (N_20249,N_18750,N_18754);
or U20250 (N_20250,N_18307,N_18965);
and U20251 (N_20251,N_19151,N_18054);
xor U20252 (N_20252,N_18770,N_18638);
and U20253 (N_20253,N_18087,N_18412);
nand U20254 (N_20254,N_19122,N_18308);
nor U20255 (N_20255,N_18917,N_18925);
xor U20256 (N_20256,N_18468,N_18287);
or U20257 (N_20257,N_18987,N_19193);
xnor U20258 (N_20258,N_18059,N_18920);
nand U20259 (N_20259,N_18674,N_19001);
or U20260 (N_20260,N_18208,N_18976);
nor U20261 (N_20261,N_18254,N_18668);
nand U20262 (N_20262,N_18086,N_18909);
nand U20263 (N_20263,N_18997,N_18618);
or U20264 (N_20264,N_19119,N_18152);
xor U20265 (N_20265,N_18242,N_18810);
xor U20266 (N_20266,N_18112,N_18017);
xnor U20267 (N_20267,N_19115,N_18639);
or U20268 (N_20268,N_18436,N_18587);
nand U20269 (N_20269,N_19022,N_18375);
or U20270 (N_20270,N_18672,N_19190);
nor U20271 (N_20271,N_18824,N_18730);
xnor U20272 (N_20272,N_18529,N_18168);
or U20273 (N_20273,N_19138,N_18282);
and U20274 (N_20274,N_18072,N_19140);
nor U20275 (N_20275,N_18111,N_18178);
nand U20276 (N_20276,N_18437,N_18544);
and U20277 (N_20277,N_18494,N_18917);
and U20278 (N_20278,N_18244,N_18405);
nand U20279 (N_20279,N_18324,N_19173);
xnor U20280 (N_20280,N_18416,N_19049);
or U20281 (N_20281,N_18193,N_18749);
and U20282 (N_20282,N_18109,N_18395);
nor U20283 (N_20283,N_18960,N_18194);
nor U20284 (N_20284,N_18367,N_18584);
or U20285 (N_20285,N_18353,N_18912);
nor U20286 (N_20286,N_18112,N_18087);
nor U20287 (N_20287,N_18917,N_18789);
and U20288 (N_20288,N_18914,N_18585);
nand U20289 (N_20289,N_18625,N_18496);
or U20290 (N_20290,N_18249,N_18712);
nand U20291 (N_20291,N_18225,N_18979);
xnor U20292 (N_20292,N_18807,N_18512);
xnor U20293 (N_20293,N_18458,N_19091);
nor U20294 (N_20294,N_18590,N_18448);
nor U20295 (N_20295,N_18557,N_18971);
nand U20296 (N_20296,N_18319,N_19044);
and U20297 (N_20297,N_18443,N_18225);
nor U20298 (N_20298,N_18035,N_18058);
or U20299 (N_20299,N_18956,N_18076);
xor U20300 (N_20300,N_19046,N_18018);
and U20301 (N_20301,N_18289,N_19065);
xnor U20302 (N_20302,N_18030,N_18268);
nand U20303 (N_20303,N_19195,N_18554);
or U20304 (N_20304,N_18737,N_18834);
xnor U20305 (N_20305,N_18517,N_18519);
and U20306 (N_20306,N_19136,N_18867);
nor U20307 (N_20307,N_18944,N_18041);
nor U20308 (N_20308,N_18768,N_18616);
and U20309 (N_20309,N_19144,N_18614);
and U20310 (N_20310,N_19198,N_18449);
or U20311 (N_20311,N_19100,N_18641);
nor U20312 (N_20312,N_18012,N_19048);
nor U20313 (N_20313,N_19065,N_18714);
nor U20314 (N_20314,N_18418,N_18249);
and U20315 (N_20315,N_18526,N_19141);
xnor U20316 (N_20316,N_19109,N_18326);
or U20317 (N_20317,N_18952,N_18520);
nor U20318 (N_20318,N_18240,N_19090);
or U20319 (N_20319,N_19187,N_19097);
nor U20320 (N_20320,N_18547,N_18862);
or U20321 (N_20321,N_18183,N_18566);
nor U20322 (N_20322,N_18133,N_18715);
and U20323 (N_20323,N_18905,N_18447);
nor U20324 (N_20324,N_18017,N_18637);
nand U20325 (N_20325,N_18098,N_18622);
nand U20326 (N_20326,N_18879,N_18917);
nor U20327 (N_20327,N_18872,N_19085);
or U20328 (N_20328,N_19092,N_18005);
xnor U20329 (N_20329,N_18827,N_18873);
or U20330 (N_20330,N_19006,N_18214);
nand U20331 (N_20331,N_19102,N_18037);
or U20332 (N_20332,N_18529,N_18002);
nand U20333 (N_20333,N_18288,N_18645);
xor U20334 (N_20334,N_18975,N_18259);
nand U20335 (N_20335,N_18897,N_18215);
nand U20336 (N_20336,N_18848,N_18206);
nor U20337 (N_20337,N_18621,N_18372);
nor U20338 (N_20338,N_18039,N_18114);
xor U20339 (N_20339,N_18192,N_19138);
or U20340 (N_20340,N_18952,N_18308);
nand U20341 (N_20341,N_18820,N_19125);
xor U20342 (N_20342,N_18792,N_18729);
nor U20343 (N_20343,N_18744,N_18030);
and U20344 (N_20344,N_19091,N_18691);
xor U20345 (N_20345,N_18333,N_18930);
or U20346 (N_20346,N_18667,N_18884);
xor U20347 (N_20347,N_18884,N_18188);
and U20348 (N_20348,N_18713,N_18841);
or U20349 (N_20349,N_18995,N_19124);
and U20350 (N_20350,N_18649,N_18009);
xnor U20351 (N_20351,N_18148,N_18340);
or U20352 (N_20352,N_18602,N_18229);
and U20353 (N_20353,N_18409,N_19121);
nand U20354 (N_20354,N_19130,N_18617);
nor U20355 (N_20355,N_18503,N_18264);
nor U20356 (N_20356,N_18064,N_18068);
xnor U20357 (N_20357,N_18186,N_18961);
nand U20358 (N_20358,N_18506,N_18203);
or U20359 (N_20359,N_18929,N_19150);
nor U20360 (N_20360,N_18538,N_18350);
nand U20361 (N_20361,N_18297,N_18652);
xor U20362 (N_20362,N_19102,N_18164);
or U20363 (N_20363,N_18970,N_18601);
or U20364 (N_20364,N_18385,N_18196);
and U20365 (N_20365,N_18713,N_18577);
or U20366 (N_20366,N_18776,N_19084);
nand U20367 (N_20367,N_18015,N_18042);
and U20368 (N_20368,N_18454,N_18974);
nand U20369 (N_20369,N_18185,N_19054);
or U20370 (N_20370,N_18579,N_18464);
or U20371 (N_20371,N_19046,N_18659);
xor U20372 (N_20372,N_18458,N_18301);
nand U20373 (N_20373,N_18229,N_19199);
xnor U20374 (N_20374,N_18289,N_18506);
or U20375 (N_20375,N_18006,N_18269);
nor U20376 (N_20376,N_19041,N_18042);
xor U20377 (N_20377,N_18253,N_18734);
or U20378 (N_20378,N_18768,N_18917);
nand U20379 (N_20379,N_19034,N_18119);
and U20380 (N_20380,N_18749,N_18686);
xnor U20381 (N_20381,N_18726,N_19130);
xnor U20382 (N_20382,N_18384,N_18906);
xor U20383 (N_20383,N_19174,N_18582);
or U20384 (N_20384,N_18630,N_18657);
and U20385 (N_20385,N_18219,N_18018);
nor U20386 (N_20386,N_18615,N_18563);
or U20387 (N_20387,N_18515,N_18301);
and U20388 (N_20388,N_18996,N_19140);
nand U20389 (N_20389,N_18636,N_18012);
xnor U20390 (N_20390,N_18714,N_18870);
nand U20391 (N_20391,N_18516,N_18805);
and U20392 (N_20392,N_19157,N_18663);
nand U20393 (N_20393,N_18243,N_18542);
xnor U20394 (N_20394,N_18940,N_18149);
nor U20395 (N_20395,N_18684,N_18735);
or U20396 (N_20396,N_18266,N_18373);
or U20397 (N_20397,N_18882,N_18462);
or U20398 (N_20398,N_18248,N_18944);
nand U20399 (N_20399,N_18070,N_18002);
xor U20400 (N_20400,N_19998,N_19364);
nand U20401 (N_20401,N_19965,N_20053);
xnor U20402 (N_20402,N_19784,N_19827);
xnor U20403 (N_20403,N_19456,N_20078);
or U20404 (N_20404,N_20373,N_19297);
nor U20405 (N_20405,N_20188,N_19569);
and U20406 (N_20406,N_19306,N_20204);
or U20407 (N_20407,N_20353,N_19481);
nor U20408 (N_20408,N_19863,N_20161);
nor U20409 (N_20409,N_20362,N_20144);
nand U20410 (N_20410,N_19338,N_19346);
and U20411 (N_20411,N_19415,N_19752);
nor U20412 (N_20412,N_19988,N_19514);
nand U20413 (N_20413,N_19851,N_19220);
nand U20414 (N_20414,N_20192,N_20147);
nor U20415 (N_20415,N_19386,N_19910);
xor U20416 (N_20416,N_19465,N_19337);
xor U20417 (N_20417,N_20396,N_20319);
xor U20418 (N_20418,N_19219,N_19410);
nand U20419 (N_20419,N_19906,N_20110);
nand U20420 (N_20420,N_19258,N_19432);
nor U20421 (N_20421,N_20339,N_19886);
or U20422 (N_20422,N_19589,N_20072);
nor U20423 (N_20423,N_19417,N_19896);
nand U20424 (N_20424,N_20342,N_20334);
or U20425 (N_20425,N_19250,N_19796);
nor U20426 (N_20426,N_19881,N_19763);
nor U20427 (N_20427,N_19257,N_19530);
xnor U20428 (N_20428,N_19603,N_19550);
nand U20429 (N_20429,N_19421,N_20018);
and U20430 (N_20430,N_19332,N_20357);
nor U20431 (N_20431,N_19807,N_20379);
xnor U20432 (N_20432,N_19838,N_19620);
and U20433 (N_20433,N_19503,N_19388);
nor U20434 (N_20434,N_19290,N_19591);
or U20435 (N_20435,N_20366,N_20142);
nor U20436 (N_20436,N_19358,N_19643);
and U20437 (N_20437,N_20191,N_19246);
or U20438 (N_20438,N_20386,N_19624);
and U20439 (N_20439,N_20063,N_19307);
xnor U20440 (N_20440,N_19675,N_20257);
and U20441 (N_20441,N_19314,N_19983);
nor U20442 (N_20442,N_20202,N_19995);
nand U20443 (N_20443,N_20069,N_20076);
or U20444 (N_20444,N_19333,N_19535);
and U20445 (N_20445,N_19966,N_19962);
and U20446 (N_20446,N_19731,N_19518);
nand U20447 (N_20447,N_19210,N_19800);
nand U20448 (N_20448,N_20274,N_19485);
and U20449 (N_20449,N_19335,N_20114);
nor U20450 (N_20450,N_20228,N_19799);
xor U20451 (N_20451,N_20197,N_20231);
nor U20452 (N_20452,N_19859,N_20208);
nor U20453 (N_20453,N_19522,N_20020);
xnor U20454 (N_20454,N_19814,N_19304);
and U20455 (N_20455,N_20329,N_19952);
nand U20456 (N_20456,N_20042,N_19967);
nand U20457 (N_20457,N_19590,N_20187);
nor U20458 (N_20458,N_20303,N_19991);
nor U20459 (N_20459,N_20037,N_19561);
nand U20460 (N_20460,N_19607,N_19657);
nor U20461 (N_20461,N_19272,N_20252);
xnor U20462 (N_20462,N_20213,N_19493);
and U20463 (N_20463,N_20256,N_19549);
xnor U20464 (N_20464,N_19292,N_19982);
nand U20465 (N_20465,N_19804,N_19371);
and U20466 (N_20466,N_19733,N_19725);
nor U20467 (N_20467,N_19336,N_19226);
nand U20468 (N_20468,N_19263,N_20012);
xor U20469 (N_20469,N_19266,N_19626);
and U20470 (N_20470,N_20101,N_19638);
xor U20471 (N_20471,N_19958,N_20013);
xor U20472 (N_20472,N_19444,N_19699);
nor U20473 (N_20473,N_19204,N_20295);
nand U20474 (N_20474,N_19259,N_20064);
xnor U20475 (N_20475,N_19368,N_20368);
xnor U20476 (N_20476,N_19283,N_19565);
nor U20477 (N_20477,N_20333,N_19779);
nor U20478 (N_20478,N_19564,N_19761);
and U20479 (N_20479,N_19217,N_20314);
or U20480 (N_20480,N_19667,N_19331);
or U20481 (N_20481,N_19370,N_19671);
nor U20482 (N_20482,N_20091,N_19883);
nor U20483 (N_20483,N_19319,N_20022);
and U20484 (N_20484,N_19653,N_19941);
nor U20485 (N_20485,N_19512,N_20381);
nand U20486 (N_20486,N_19918,N_19323);
and U20487 (N_20487,N_19679,N_20394);
xnor U20488 (N_20488,N_20308,N_19367);
xnor U20489 (N_20489,N_20145,N_19401);
and U20490 (N_20490,N_19477,N_19637);
nor U20491 (N_20491,N_20121,N_20002);
and U20492 (N_20492,N_20137,N_20027);
nor U20493 (N_20493,N_20341,N_19762);
xor U20494 (N_20494,N_20085,N_20289);
xnor U20495 (N_20495,N_20277,N_19207);
nand U20496 (N_20496,N_19377,N_19789);
and U20497 (N_20497,N_19553,N_19347);
nor U20498 (N_20498,N_20209,N_20116);
nor U20499 (N_20499,N_19686,N_19802);
and U20500 (N_20500,N_19909,N_19855);
and U20501 (N_20501,N_19341,N_19900);
nand U20502 (N_20502,N_20105,N_20235);
nor U20503 (N_20503,N_19632,N_20302);
and U20504 (N_20504,N_19580,N_19531);
nor U20505 (N_20505,N_19869,N_19466);
nor U20506 (N_20506,N_19646,N_19280);
or U20507 (N_20507,N_19354,N_20138);
nand U20508 (N_20508,N_19443,N_20071);
nor U20509 (N_20509,N_19539,N_19633);
and U20510 (N_20510,N_19769,N_19957);
nor U20511 (N_20511,N_19935,N_20151);
nand U20512 (N_20512,N_19943,N_19911);
or U20513 (N_20513,N_19684,N_19422);
nor U20514 (N_20514,N_19730,N_19760);
nand U20515 (N_20515,N_19495,N_19841);
nor U20516 (N_20516,N_20221,N_20107);
nand U20517 (N_20517,N_19451,N_19666);
and U20518 (N_20518,N_20306,N_19287);
nor U20519 (N_20519,N_19221,N_19641);
nor U20520 (N_20520,N_20016,N_19857);
and U20521 (N_20521,N_19703,N_19599);
nor U20522 (N_20522,N_20359,N_19571);
or U20523 (N_20523,N_20172,N_19772);
nor U20524 (N_20524,N_19406,N_19889);
xor U20525 (N_20525,N_20031,N_19892);
or U20526 (N_20526,N_19449,N_20040);
nor U20527 (N_20527,N_19606,N_20011);
and U20528 (N_20528,N_19714,N_19588);
or U20529 (N_20529,N_19527,N_19473);
xnor U20530 (N_20530,N_19985,N_20205);
or U20531 (N_20531,N_19915,N_19541);
xor U20532 (N_20532,N_19515,N_19426);
or U20533 (N_20533,N_20021,N_20177);
and U20534 (N_20534,N_19200,N_19349);
and U20535 (N_20535,N_20301,N_20203);
nand U20536 (N_20536,N_20033,N_20247);
nor U20537 (N_20537,N_19999,N_20025);
xnor U20538 (N_20538,N_19291,N_19668);
or U20539 (N_20539,N_19865,N_19794);
and U20540 (N_20540,N_20195,N_19931);
or U20541 (N_20541,N_19930,N_20146);
and U20542 (N_20542,N_19510,N_19391);
nor U20543 (N_20543,N_19871,N_19395);
or U20544 (N_20544,N_20350,N_19617);
and U20545 (N_20545,N_19592,N_19954);
or U20546 (N_20546,N_19317,N_19236);
xor U20547 (N_20547,N_19662,N_19526);
or U20548 (N_20548,N_20399,N_19251);
or U20549 (N_20549,N_19487,N_19720);
nand U20550 (N_20550,N_19390,N_20060);
or U20551 (N_20551,N_20181,N_19939);
nand U20552 (N_20552,N_19665,N_19570);
nand U20553 (N_20553,N_19458,N_19436);
nor U20554 (N_20554,N_19254,N_19212);
and U20555 (N_20555,N_19608,N_19300);
and U20556 (N_20556,N_19551,N_19833);
nor U20557 (N_20557,N_20307,N_20113);
xnor U20558 (N_20558,N_19489,N_19741);
xnor U20559 (N_20559,N_19384,N_19398);
or U20560 (N_20560,N_19378,N_19205);
or U20561 (N_20561,N_20226,N_20075);
or U20562 (N_20562,N_19735,N_20123);
or U20563 (N_20563,N_20248,N_19506);
and U20564 (N_20564,N_19424,N_19659);
xor U20565 (N_20565,N_19284,N_19381);
xnor U20566 (N_20566,N_19340,N_19225);
xnor U20567 (N_20567,N_20038,N_19791);
nand U20568 (N_20568,N_19834,N_20236);
xnor U20569 (N_20569,N_19955,N_19989);
or U20570 (N_20570,N_20304,N_19276);
or U20571 (N_20571,N_19427,N_19308);
nand U20572 (N_20572,N_20288,N_19673);
and U20573 (N_20573,N_19650,N_19818);
nor U20574 (N_20574,N_19598,N_19343);
nand U20575 (N_20575,N_20019,N_20239);
and U20576 (N_20576,N_20176,N_20264);
and U20577 (N_20577,N_20153,N_19862);
xnor U20578 (N_20578,N_19704,N_19285);
xor U20579 (N_20579,N_20154,N_20265);
nor U20580 (N_20580,N_19959,N_19969);
nor U20581 (N_20581,N_19584,N_19694);
or U20582 (N_20582,N_20272,N_20152);
and U20583 (N_20583,N_20266,N_20215);
nor U20584 (N_20584,N_19867,N_20238);
nand U20585 (N_20585,N_19743,N_19594);
nand U20586 (N_20586,N_19600,N_19680);
nor U20587 (N_20587,N_19609,N_20294);
nor U20588 (N_20588,N_19475,N_19375);
nand U20589 (N_20589,N_19396,N_19310);
nor U20590 (N_20590,N_19759,N_20321);
or U20591 (N_20591,N_19929,N_19687);
nand U20592 (N_20592,N_19562,N_19322);
nor U20593 (N_20593,N_19233,N_20185);
xor U20594 (N_20594,N_19293,N_19718);
nor U20595 (N_20595,N_19739,N_19576);
nor U20596 (N_20596,N_19279,N_20035);
nand U20597 (N_20597,N_20249,N_19414);
or U20598 (N_20598,N_20349,N_19655);
or U20599 (N_20599,N_19615,N_20131);
or U20600 (N_20600,N_20008,N_19438);
nor U20601 (N_20601,N_19925,N_19628);
and U20602 (N_20602,N_20062,N_19275);
nor U20603 (N_20603,N_19877,N_19708);
or U20604 (N_20604,N_19873,N_19234);
or U20605 (N_20605,N_19843,N_20074);
nand U20606 (N_20606,N_20026,N_20229);
xnor U20607 (N_20607,N_19819,N_19298);
nand U20608 (N_20608,N_19810,N_19996);
or U20609 (N_20609,N_19492,N_20164);
and U20610 (N_20610,N_19932,N_19472);
nand U20611 (N_20611,N_19888,N_20029);
nor U20612 (N_20612,N_19854,N_20007);
or U20613 (N_20613,N_20331,N_20099);
xor U20614 (N_20614,N_20365,N_20190);
or U20615 (N_20615,N_19927,N_20001);
nand U20616 (N_20616,N_20242,N_20118);
nand U20617 (N_20617,N_19719,N_19216);
and U20618 (N_20618,N_19578,N_19705);
xor U20619 (N_20619,N_20270,N_20380);
nor U20620 (N_20620,N_19602,N_20312);
and U20621 (N_20621,N_19270,N_19747);
or U20622 (N_20622,N_20047,N_20360);
xnor U20623 (N_20623,N_19328,N_19664);
or U20624 (N_20624,N_19920,N_20377);
or U20625 (N_20625,N_19788,N_19245);
and U20626 (N_20626,N_20096,N_20382);
nand U20627 (N_20627,N_19459,N_19677);
or U20628 (N_20628,N_19893,N_19875);
nand U20629 (N_20629,N_19946,N_19907);
or U20630 (N_20630,N_20230,N_20286);
nor U20631 (N_20631,N_19716,N_19866);
nor U20632 (N_20632,N_19479,N_19711);
nor U20633 (N_20633,N_19261,N_19764);
nand U20634 (N_20634,N_19621,N_20196);
nand U20635 (N_20635,N_19474,N_20034);
nand U20636 (N_20636,N_19636,N_20119);
or U20637 (N_20637,N_19555,N_19848);
nand U20638 (N_20638,N_19498,N_19385);
and U20639 (N_20639,N_20067,N_19790);
xor U20640 (N_20640,N_19501,N_19237);
nand U20641 (N_20641,N_19548,N_20348);
or U20642 (N_20642,N_20262,N_20059);
or U20643 (N_20643,N_20251,N_20108);
nor U20644 (N_20644,N_19256,N_19729);
nor U20645 (N_20645,N_20030,N_19691);
nor U20646 (N_20646,N_19547,N_19454);
xnor U20647 (N_20647,N_19360,N_20343);
xnor U20648 (N_20648,N_19441,N_20255);
nand U20649 (N_20649,N_19698,N_19742);
and U20650 (N_20650,N_19230,N_19971);
or U20651 (N_20651,N_19658,N_20175);
xnor U20652 (N_20652,N_19861,N_19945);
or U20653 (N_20653,N_19605,N_19960);
xnor U20654 (N_20654,N_19901,N_19654);
and U20655 (N_20655,N_19619,N_19339);
or U20656 (N_20656,N_19575,N_19774);
and U20657 (N_20657,N_19899,N_20148);
nand U20658 (N_20658,N_20328,N_19728);
nand U20659 (N_20659,N_20160,N_19469);
xnor U20660 (N_20660,N_19423,N_20070);
or U20661 (N_20661,N_19844,N_19651);
nand U20662 (N_20662,N_19648,N_19849);
xnor U20663 (N_20663,N_20309,N_20345);
xor U20664 (N_20664,N_19815,N_20244);
nand U20665 (N_20665,N_19478,N_19404);
or U20666 (N_20666,N_20092,N_19924);
nor U20667 (N_20667,N_19897,N_19228);
nor U20668 (N_20668,N_19649,N_20170);
or U20669 (N_20669,N_19921,N_20158);
nor U20670 (N_20670,N_20254,N_20102);
or U20671 (N_20671,N_19975,N_19842);
or U20672 (N_20672,N_19509,N_19235);
nand U20673 (N_20673,N_19483,N_20260);
nor U20674 (N_20674,N_20135,N_19350);
nand U20675 (N_20675,N_19357,N_20003);
nor U20676 (N_20676,N_19533,N_19832);
nor U20677 (N_20677,N_19579,N_19723);
xor U20678 (N_20678,N_20206,N_20337);
nor U20679 (N_20679,N_19745,N_19542);
and U20680 (N_20680,N_19872,N_20278);
or U20681 (N_20681,N_19273,N_20237);
nor U20682 (N_20682,N_19271,N_20287);
or U20683 (N_20683,N_19614,N_19734);
and U20684 (N_20684,N_19712,N_19903);
or U20685 (N_20685,N_19977,N_19302);
nand U20686 (N_20686,N_19964,N_20139);
nor U20687 (N_20687,N_20155,N_19211);
xor U20688 (N_20688,N_19811,N_19693);
or U20689 (N_20689,N_19644,N_19778);
nor U20690 (N_20690,N_19963,N_19242);
nand U20691 (N_20691,N_20182,N_20245);
nor U20692 (N_20692,N_20082,N_19738);
and U20693 (N_20693,N_19351,N_19768);
nor U20694 (N_20694,N_19968,N_20088);
and U20695 (N_20695,N_19688,N_20372);
nand U20696 (N_20696,N_19560,N_19356);
xor U20697 (N_20697,N_20388,N_20010);
nor U20698 (N_20698,N_19353,N_20103);
and U20699 (N_20699,N_19222,N_19631);
and U20700 (N_20700,N_19853,N_20117);
xnor U20701 (N_20701,N_19919,N_19532);
nor U20702 (N_20702,N_20065,N_19203);
xnor U20703 (N_20703,N_20178,N_20327);
nand U20704 (N_20704,N_19468,N_19467);
and U20705 (N_20705,N_20391,N_19826);
or U20706 (N_20706,N_20273,N_19365);
xor U20707 (N_20707,N_19201,N_19403);
nor U20708 (N_20708,N_20212,N_19647);
xor U20709 (N_20709,N_19836,N_19260);
and U20710 (N_20710,N_19215,N_19326);
and U20711 (N_20711,N_19462,N_19990);
and U20712 (N_20712,N_19816,N_20214);
or U20713 (N_20713,N_19808,N_19223);
nor U20714 (N_20714,N_20057,N_20336);
or U20715 (N_20715,N_19218,N_19597);
or U20716 (N_20716,N_19978,N_20315);
nand U20717 (N_20717,N_19858,N_19979);
nand U20718 (N_20718,N_19253,N_19616);
xor U20719 (N_20719,N_19786,N_19255);
or U20720 (N_20720,N_19572,N_20090);
xnor U20721 (N_20721,N_19405,N_19635);
xor U20722 (N_20722,N_20267,N_19268);
nor U20723 (N_20723,N_19721,N_19566);
nor U20724 (N_20724,N_20384,N_19757);
nand U20725 (N_20725,N_20055,N_20173);
and U20726 (N_20726,N_19613,N_20130);
and U20727 (N_20727,N_20335,N_19824);
nor U20728 (N_20728,N_19244,N_20028);
and U20729 (N_20729,N_19868,N_20004);
xor U20730 (N_20730,N_19431,N_19981);
or U20731 (N_20731,N_19448,N_20169);
xnor U20732 (N_20732,N_19435,N_19724);
xor U20733 (N_20733,N_20310,N_19828);
nand U20734 (N_20734,N_19545,N_19685);
xor U20735 (N_20735,N_19612,N_19519);
nand U20736 (N_20736,N_19732,N_19296);
xnor U20737 (N_20737,N_20299,N_19315);
xnor U20738 (N_20738,N_19372,N_20198);
xor U20739 (N_20739,N_19793,N_19722);
or U20740 (N_20740,N_19209,N_19581);
or U20741 (N_20741,N_19318,N_19894);
nand U20742 (N_20742,N_19249,N_19394);
xor U20743 (N_20743,N_19656,N_19277);
xor U20744 (N_20744,N_20324,N_20376);
and U20745 (N_20745,N_19683,N_20189);
nor U20746 (N_20746,N_20149,N_20290);
nor U20747 (N_20747,N_19311,N_19864);
nand U20748 (N_20748,N_20036,N_19773);
nand U20749 (N_20749,N_19880,N_20320);
and U20750 (N_20750,N_19563,N_20271);
or U20751 (N_20751,N_19830,N_20375);
nand U20752 (N_20752,N_19574,N_20106);
nand U20753 (N_20753,N_20371,N_19630);
or U20754 (N_20754,N_19480,N_19709);
xnor U20755 (N_20755,N_19587,N_19885);
and U20756 (N_20756,N_19697,N_19812);
nand U20757 (N_20757,N_19846,N_19765);
and U20758 (N_20758,N_19392,N_19442);
nor U20759 (N_20759,N_19744,N_20332);
xor U20760 (N_20760,N_20369,N_19992);
xor U20761 (N_20761,N_19727,N_19274);
nor U20762 (N_20762,N_19402,N_20005);
nand U20763 (N_20763,N_19879,N_19439);
and U20764 (N_20764,N_19922,N_20387);
xnor U20765 (N_20765,N_19513,N_19416);
nor U20766 (N_20766,N_20300,N_20136);
or U20767 (N_20767,N_20279,N_19663);
nor U20768 (N_20768,N_19625,N_20241);
nand U20769 (N_20769,N_19269,N_19970);
xnor U20770 (N_20770,N_19681,N_19520);
nor U20771 (N_20771,N_19248,N_19383);
xnor U20772 (N_20772,N_19238,N_20133);
xnor U20773 (N_20773,N_19289,N_19330);
and U20774 (N_20774,N_20186,N_20081);
nor U20775 (N_20775,N_19652,N_20087);
nor U20776 (N_20776,N_19455,N_19379);
or U20777 (N_20777,N_19460,N_19433);
or U20778 (N_20778,N_19767,N_19419);
xnor U20779 (N_20779,N_20363,N_19239);
nand U20780 (N_20780,N_19316,N_19912);
nor U20781 (N_20781,N_19334,N_20084);
nor U20782 (N_20782,N_20323,N_20068);
nand U20783 (N_20783,N_19825,N_19882);
and U20784 (N_20784,N_19707,N_20017);
xnor U20785 (N_20785,N_19345,N_19627);
xor U20786 (N_20786,N_19953,N_19453);
or U20787 (N_20787,N_19700,N_20268);
and U20788 (N_20788,N_19782,N_19874);
nor U20789 (N_20789,N_19488,N_19890);
xnor U20790 (N_20790,N_19408,N_20162);
or U20791 (N_20791,N_19552,N_20127);
nand U20792 (N_20792,N_20109,N_20397);
nand U20793 (N_20793,N_20043,N_19247);
xnor U20794 (N_20794,N_19511,N_20165);
nor U20795 (N_20795,N_20233,N_19822);
and U20796 (N_20796,N_20398,N_20234);
xnor U20797 (N_20797,N_20193,N_20222);
nor U20798 (N_20798,N_19938,N_19944);
xnor U20799 (N_20799,N_19777,N_20132);
nor U20800 (N_20800,N_19710,N_19813);
nand U20801 (N_20801,N_20352,N_20141);
nand U20802 (N_20802,N_19984,N_20383);
nor U20803 (N_20803,N_19393,N_19523);
or U20804 (N_20804,N_19771,N_19286);
nand U20805 (N_20805,N_20200,N_19583);
xor U20806 (N_20806,N_19715,N_19775);
nand U20807 (N_20807,N_19781,N_19840);
or U20808 (N_20808,N_20066,N_19536);
xor U20809 (N_20809,N_19876,N_19736);
xor U20810 (N_20810,N_19726,N_19471);
nand U20811 (N_20811,N_19327,N_20305);
nor U20812 (N_20812,N_19766,N_20325);
xnor U20813 (N_20813,N_19792,N_20318);
xor U20814 (N_20814,N_19281,N_19577);
nor U20815 (N_20815,N_19947,N_20166);
and U20816 (N_20816,N_19837,N_19803);
nand U20817 (N_20817,N_19546,N_19342);
or U20818 (N_20818,N_20095,N_20243);
xnor U20819 (N_20819,N_19457,N_19329);
nand U20820 (N_20820,N_19692,N_19490);
and U20821 (N_20821,N_19785,N_20171);
and U20822 (N_20822,N_20183,N_20098);
xnor U20823 (N_20823,N_19937,N_19312);
nand U20824 (N_20824,N_19213,N_20207);
nand U20825 (N_20825,N_20385,N_19387);
or U20826 (N_20826,N_19748,N_19887);
nor U20827 (N_20827,N_19642,N_19908);
nor U20828 (N_20828,N_19610,N_19231);
nand U20829 (N_20829,N_20389,N_20216);
or U20830 (N_20830,N_19676,N_20378);
nor U20831 (N_20831,N_20199,N_19904);
nand U20832 (N_20832,N_20015,N_19753);
xor U20833 (N_20833,N_19740,N_19267);
xor U20834 (N_20834,N_19325,N_20126);
or U20835 (N_20835,N_19986,N_19770);
nand U20836 (N_20836,N_19505,N_19850);
xor U20837 (N_20837,N_19993,N_19623);
xor U20838 (N_20838,N_20326,N_19362);
and U20839 (N_20839,N_19634,N_20048);
nand U20840 (N_20840,N_20293,N_20250);
or U20841 (N_20841,N_19973,N_19829);
nor U20842 (N_20842,N_19913,N_19695);
or U20843 (N_20843,N_19409,N_19412);
and U20844 (N_20844,N_19847,N_19240);
nor U20845 (N_20845,N_19278,N_19702);
nor U20846 (N_20846,N_20393,N_20058);
and U20847 (N_20847,N_19507,N_19497);
and U20848 (N_20848,N_19557,N_19593);
nor U20849 (N_20849,N_20317,N_19949);
xor U20850 (N_20850,N_20044,N_19554);
nand U20851 (N_20851,N_19573,N_19437);
nand U20852 (N_20852,N_19420,N_19852);
xnor U20853 (N_20853,N_20184,N_20258);
nand U20854 (N_20854,N_20282,N_20280);
nand U20855 (N_20855,N_20049,N_19309);
nand U20856 (N_20856,N_19363,N_19916);
nand U20857 (N_20857,N_20129,N_19696);
nand U20858 (N_20858,N_20023,N_20358);
nand U20859 (N_20859,N_19482,N_19756);
nand U20860 (N_20860,N_20051,N_19529);
and U20861 (N_20861,N_19817,N_19987);
nand U20862 (N_20862,N_19359,N_19713);
nor U20863 (N_20863,N_19224,N_19678);
xnor U20864 (N_20864,N_19798,N_19596);
xor U20865 (N_20865,N_19961,N_19208);
nor U20866 (N_20866,N_20240,N_19556);
and U20867 (N_20867,N_19568,N_19229);
nand U20868 (N_20868,N_19202,N_20291);
and U20869 (N_20869,N_19926,N_20374);
xnor U20870 (N_20870,N_19936,N_19543);
nor U20871 (N_20871,N_20159,N_19461);
nand U20872 (N_20872,N_19355,N_20163);
or U20873 (N_20873,N_20330,N_20297);
and U20874 (N_20874,N_19538,N_20218);
xnor U20875 (N_20875,N_19486,N_20322);
nand U20876 (N_20876,N_20150,N_19418);
and U20877 (N_20877,N_20125,N_20024);
nor U20878 (N_20878,N_19674,N_19504);
nor U20879 (N_20879,N_19750,N_19682);
or U20880 (N_20880,N_19629,N_19942);
nor U20881 (N_20881,N_19352,N_20263);
nand U20882 (N_20882,N_20006,N_19878);
and U20883 (N_20883,N_20367,N_19524);
nor U20884 (N_20884,N_19265,N_20281);
or U20885 (N_20885,N_19320,N_19809);
nor U20886 (N_20886,N_19321,N_19956);
and U20887 (N_20887,N_20219,N_19407);
nand U20888 (N_20888,N_20351,N_19494);
xor U20889 (N_20889,N_20168,N_19950);
nand U20890 (N_20890,N_19373,N_19934);
nand U20891 (N_20891,N_19380,N_19434);
nor U20892 (N_20892,N_19399,N_19400);
nand U20893 (N_20893,N_20354,N_19951);
and U20894 (N_20894,N_19749,N_19301);
nand U20895 (N_20895,N_19540,N_20009);
nor U20896 (N_20896,N_20283,N_19940);
and U20897 (N_20897,N_19476,N_19997);
xnor U20898 (N_20898,N_20223,N_20045);
nor U20899 (N_20899,N_19496,N_19502);
xnor U20900 (N_20900,N_19559,N_20225);
or U20901 (N_20901,N_19411,N_19820);
nor U20902 (N_20902,N_19348,N_19517);
or U20903 (N_20903,N_20211,N_20284);
or U20904 (N_20904,N_20000,N_19758);
nand U20905 (N_20905,N_19528,N_19839);
nor U20906 (N_20906,N_20346,N_19914);
nand U20907 (N_20907,N_19464,N_19537);
or U20908 (N_20908,N_19282,N_19689);
xor U20909 (N_20909,N_20157,N_20167);
and U20910 (N_20910,N_19660,N_19382);
or U20911 (N_20911,N_19463,N_20086);
nand U20912 (N_20912,N_20054,N_19611);
and U20913 (N_20913,N_20298,N_19622);
xnor U20914 (N_20914,N_19717,N_20120);
nor U20915 (N_20915,N_19917,N_19928);
nand U20916 (N_20916,N_19484,N_19369);
nand U20917 (N_20917,N_19980,N_20128);
or U20918 (N_20918,N_19706,N_20039);
nand U20919 (N_20919,N_19823,N_20246);
xor U20920 (N_20920,N_19366,N_19835);
nand U20921 (N_20921,N_19534,N_19783);
xnor U20922 (N_20922,N_19299,N_19303);
and U20923 (N_20923,N_20080,N_20210);
and U20924 (N_20924,N_20041,N_20052);
and U20925 (N_20925,N_20104,N_19214);
nor U20926 (N_20926,N_19445,N_20392);
or U20927 (N_20927,N_20180,N_19845);
or U20928 (N_20928,N_20338,N_19521);
nand U20929 (N_20929,N_20276,N_20390);
or U20930 (N_20930,N_20364,N_19670);
xor U20931 (N_20931,N_19801,N_19787);
nor U20932 (N_20932,N_19586,N_20083);
nand U20933 (N_20933,N_20077,N_20269);
nand U20934 (N_20934,N_19313,N_20032);
nand U20935 (N_20935,N_19544,N_19884);
xor U20936 (N_20936,N_19923,N_19595);
nor U20937 (N_20937,N_20046,N_20356);
or U20938 (N_20938,N_19232,N_19821);
and U20939 (N_20939,N_19206,N_20232);
xnor U20940 (N_20940,N_20311,N_20340);
xor U20941 (N_20941,N_20347,N_19585);
xor U20942 (N_20942,N_19499,N_19933);
and U20943 (N_20943,N_20224,N_20292);
and U20944 (N_20944,N_20355,N_20134);
nor U20945 (N_20945,N_19264,N_19905);
nor U20946 (N_20946,N_20259,N_19754);
xor U20947 (N_20947,N_20261,N_20112);
nand U20948 (N_20948,N_19500,N_20285);
and U20949 (N_20949,N_19860,N_20094);
nor U20950 (N_20950,N_19639,N_19994);
nor U20951 (N_20951,N_19376,N_20111);
nor U20952 (N_20952,N_19305,N_19948);
xor U20953 (N_20953,N_20316,N_19344);
and U20954 (N_20954,N_19601,N_20089);
nand U20955 (N_20955,N_19295,N_19425);
xor U20956 (N_20956,N_20201,N_19440);
or U20957 (N_20957,N_19525,N_20061);
xor U20958 (N_20958,N_19361,N_20073);
xnor U20959 (N_20959,N_19508,N_20097);
xor U20960 (N_20960,N_19661,N_19640);
nor U20961 (N_20961,N_19972,N_20174);
or U20962 (N_20962,N_19582,N_19294);
xnor U20963 (N_20963,N_20296,N_20140);
and U20964 (N_20964,N_19870,N_19516);
or U20965 (N_20965,N_19491,N_19902);
xor U20966 (N_20966,N_20313,N_19252);
and U20967 (N_20967,N_19746,N_19428);
xnor U20968 (N_20968,N_19262,N_20122);
and U20969 (N_20969,N_20124,N_19288);
nand U20970 (N_20970,N_19805,N_19450);
nand U20971 (N_20971,N_20093,N_20156);
nand U20972 (N_20972,N_19446,N_19751);
and U20973 (N_20973,N_19737,N_19776);
and U20974 (N_20974,N_19976,N_19452);
xnor U20975 (N_20975,N_19470,N_19701);
or U20976 (N_20976,N_19227,N_19690);
nor U20977 (N_20977,N_20143,N_19898);
and U20978 (N_20978,N_19324,N_20014);
nor U20979 (N_20979,N_19856,N_19558);
nor U20980 (N_20980,N_20115,N_20344);
nor U20981 (N_20981,N_19974,N_19604);
nor U20982 (N_20982,N_20395,N_20056);
and U20983 (N_20983,N_19430,N_19397);
nand U20984 (N_20984,N_20227,N_19672);
nor U20985 (N_20985,N_20361,N_19645);
nor U20986 (N_20986,N_20050,N_19241);
xor U20987 (N_20987,N_19389,N_19447);
or U20988 (N_20988,N_19891,N_20194);
xor U20989 (N_20989,N_19243,N_19413);
nor U20990 (N_20990,N_20370,N_19374);
nor U20991 (N_20991,N_19806,N_19831);
and U20992 (N_20992,N_19895,N_19669);
nor U20993 (N_20993,N_20275,N_20100);
xor U20994 (N_20994,N_20079,N_19429);
nor U20995 (N_20995,N_19780,N_19618);
xor U20996 (N_20996,N_19755,N_19567);
xor U20997 (N_20997,N_20220,N_20253);
nor U20998 (N_20998,N_19795,N_20217);
or U20999 (N_20999,N_20179,N_19797);
and U21000 (N_21000,N_20019,N_19373);
xnor U21001 (N_21001,N_20039,N_19505);
and U21002 (N_21002,N_19818,N_19506);
nor U21003 (N_21003,N_19413,N_19570);
nand U21004 (N_21004,N_20375,N_19630);
or U21005 (N_21005,N_19242,N_19857);
and U21006 (N_21006,N_19369,N_19998);
nand U21007 (N_21007,N_20029,N_19336);
nand U21008 (N_21008,N_19484,N_19200);
nor U21009 (N_21009,N_19275,N_19734);
and U21010 (N_21010,N_19359,N_19211);
nand U21011 (N_21011,N_19216,N_19765);
or U21012 (N_21012,N_19600,N_20347);
and U21013 (N_21013,N_20027,N_19730);
or U21014 (N_21014,N_19512,N_19479);
xnor U21015 (N_21015,N_19998,N_19910);
and U21016 (N_21016,N_20015,N_19268);
and U21017 (N_21017,N_19383,N_19297);
or U21018 (N_21018,N_20281,N_19856);
xnor U21019 (N_21019,N_19903,N_19560);
nor U21020 (N_21020,N_20303,N_20304);
or U21021 (N_21021,N_19443,N_19407);
nor U21022 (N_21022,N_20087,N_19213);
or U21023 (N_21023,N_20037,N_20063);
and U21024 (N_21024,N_20162,N_19768);
or U21025 (N_21025,N_19911,N_19611);
nand U21026 (N_21026,N_19903,N_20132);
nand U21027 (N_21027,N_19262,N_19623);
and U21028 (N_21028,N_20172,N_19731);
and U21029 (N_21029,N_19891,N_19223);
or U21030 (N_21030,N_20378,N_19817);
nand U21031 (N_21031,N_19360,N_20385);
nand U21032 (N_21032,N_19437,N_19312);
nor U21033 (N_21033,N_19460,N_19760);
or U21034 (N_21034,N_19201,N_19987);
or U21035 (N_21035,N_20285,N_19206);
and U21036 (N_21036,N_19838,N_19527);
xor U21037 (N_21037,N_20176,N_19619);
and U21038 (N_21038,N_19815,N_20348);
xnor U21039 (N_21039,N_19955,N_20258);
and U21040 (N_21040,N_19763,N_19898);
or U21041 (N_21041,N_20161,N_19387);
xor U21042 (N_21042,N_19394,N_20188);
nand U21043 (N_21043,N_19228,N_19529);
and U21044 (N_21044,N_19744,N_19596);
and U21045 (N_21045,N_19704,N_19991);
or U21046 (N_21046,N_19559,N_19737);
and U21047 (N_21047,N_19991,N_19441);
and U21048 (N_21048,N_19954,N_20139);
and U21049 (N_21049,N_20230,N_19250);
nor U21050 (N_21050,N_19878,N_19362);
xnor U21051 (N_21051,N_19640,N_19767);
nand U21052 (N_21052,N_19730,N_19340);
xor U21053 (N_21053,N_19494,N_19758);
and U21054 (N_21054,N_19859,N_20213);
and U21055 (N_21055,N_19209,N_20319);
or U21056 (N_21056,N_20151,N_19880);
nor U21057 (N_21057,N_19259,N_20296);
xnor U21058 (N_21058,N_19617,N_20018);
xor U21059 (N_21059,N_19462,N_19719);
or U21060 (N_21060,N_19993,N_19204);
or U21061 (N_21061,N_20241,N_19485);
and U21062 (N_21062,N_19670,N_20300);
and U21063 (N_21063,N_19473,N_20067);
xor U21064 (N_21064,N_20030,N_19574);
nand U21065 (N_21065,N_20299,N_19847);
nor U21066 (N_21066,N_19514,N_19921);
nor U21067 (N_21067,N_19242,N_20341);
or U21068 (N_21068,N_19550,N_20217);
xnor U21069 (N_21069,N_19823,N_19973);
nand U21070 (N_21070,N_19350,N_20064);
nor U21071 (N_21071,N_19268,N_19884);
nand U21072 (N_21072,N_19669,N_19255);
or U21073 (N_21073,N_20232,N_19568);
nor U21074 (N_21074,N_19726,N_19735);
nand U21075 (N_21075,N_20399,N_19203);
xnor U21076 (N_21076,N_19832,N_20283);
and U21077 (N_21077,N_19337,N_19768);
nand U21078 (N_21078,N_19260,N_19285);
xor U21079 (N_21079,N_20158,N_19892);
or U21080 (N_21080,N_20072,N_20387);
nand U21081 (N_21081,N_19830,N_19460);
xnor U21082 (N_21082,N_19910,N_19844);
nor U21083 (N_21083,N_20031,N_19795);
and U21084 (N_21084,N_19461,N_20069);
xor U21085 (N_21085,N_19989,N_20344);
xor U21086 (N_21086,N_19555,N_20071);
and U21087 (N_21087,N_19704,N_19529);
nand U21088 (N_21088,N_19685,N_19320);
nor U21089 (N_21089,N_20250,N_19338);
nand U21090 (N_21090,N_19684,N_19674);
or U21091 (N_21091,N_20067,N_19427);
or U21092 (N_21092,N_19614,N_20079);
or U21093 (N_21093,N_19321,N_20171);
and U21094 (N_21094,N_19247,N_20050);
or U21095 (N_21095,N_19292,N_19420);
nand U21096 (N_21096,N_19888,N_19553);
xnor U21097 (N_21097,N_20003,N_19402);
and U21098 (N_21098,N_19305,N_20211);
xnor U21099 (N_21099,N_19303,N_19420);
nand U21100 (N_21100,N_19344,N_19789);
nand U21101 (N_21101,N_19844,N_19820);
and U21102 (N_21102,N_19563,N_20384);
and U21103 (N_21103,N_19498,N_19216);
nand U21104 (N_21104,N_20178,N_19711);
nand U21105 (N_21105,N_19399,N_20187);
xnor U21106 (N_21106,N_19990,N_19488);
and U21107 (N_21107,N_19246,N_19631);
nor U21108 (N_21108,N_19696,N_19936);
or U21109 (N_21109,N_19242,N_19470);
nor U21110 (N_21110,N_19949,N_19617);
nand U21111 (N_21111,N_20330,N_19904);
xor U21112 (N_21112,N_20145,N_20148);
xor U21113 (N_21113,N_20296,N_19349);
xnor U21114 (N_21114,N_20253,N_20385);
or U21115 (N_21115,N_20129,N_19598);
or U21116 (N_21116,N_20205,N_20003);
nor U21117 (N_21117,N_19730,N_19873);
nor U21118 (N_21118,N_20102,N_20201);
nor U21119 (N_21119,N_20219,N_19612);
nand U21120 (N_21120,N_19428,N_19650);
nand U21121 (N_21121,N_20352,N_19636);
nand U21122 (N_21122,N_19685,N_19267);
and U21123 (N_21123,N_20059,N_20221);
and U21124 (N_21124,N_20378,N_20320);
or U21125 (N_21125,N_19826,N_20323);
and U21126 (N_21126,N_19695,N_19588);
or U21127 (N_21127,N_19479,N_19870);
nand U21128 (N_21128,N_19581,N_20019);
or U21129 (N_21129,N_20257,N_20314);
nand U21130 (N_21130,N_20240,N_19600);
xnor U21131 (N_21131,N_19927,N_19438);
xor U21132 (N_21132,N_20164,N_19869);
and U21133 (N_21133,N_19202,N_20140);
xnor U21134 (N_21134,N_19952,N_19475);
or U21135 (N_21135,N_19722,N_19514);
xor U21136 (N_21136,N_19937,N_20093);
or U21137 (N_21137,N_20026,N_19928);
nand U21138 (N_21138,N_19994,N_20396);
nor U21139 (N_21139,N_19336,N_19499);
nand U21140 (N_21140,N_20186,N_19581);
and U21141 (N_21141,N_20363,N_19224);
and U21142 (N_21142,N_19950,N_19278);
nor U21143 (N_21143,N_20206,N_19889);
nand U21144 (N_21144,N_19393,N_20284);
xor U21145 (N_21145,N_19518,N_20127);
or U21146 (N_21146,N_20218,N_20224);
or U21147 (N_21147,N_20299,N_19316);
or U21148 (N_21148,N_19906,N_20013);
or U21149 (N_21149,N_19506,N_19232);
xnor U21150 (N_21150,N_19535,N_20114);
nor U21151 (N_21151,N_19445,N_20099);
nor U21152 (N_21152,N_19896,N_19256);
and U21153 (N_21153,N_20032,N_19775);
xor U21154 (N_21154,N_19539,N_19640);
nor U21155 (N_21155,N_19496,N_19962);
nand U21156 (N_21156,N_20214,N_20273);
xnor U21157 (N_21157,N_20381,N_19927);
nor U21158 (N_21158,N_19808,N_20123);
nor U21159 (N_21159,N_20267,N_19966);
nand U21160 (N_21160,N_19500,N_19676);
or U21161 (N_21161,N_19204,N_19665);
or U21162 (N_21162,N_19395,N_19685);
or U21163 (N_21163,N_19916,N_19540);
nor U21164 (N_21164,N_20190,N_19531);
nor U21165 (N_21165,N_19514,N_19533);
or U21166 (N_21166,N_20148,N_20321);
and U21167 (N_21167,N_20023,N_19993);
and U21168 (N_21168,N_20325,N_19888);
and U21169 (N_21169,N_20275,N_19720);
or U21170 (N_21170,N_19896,N_20179);
nor U21171 (N_21171,N_20197,N_19959);
or U21172 (N_21172,N_20006,N_19778);
xnor U21173 (N_21173,N_20121,N_20198);
nor U21174 (N_21174,N_19393,N_19951);
xnor U21175 (N_21175,N_20245,N_19667);
nor U21176 (N_21176,N_20232,N_19704);
or U21177 (N_21177,N_20058,N_20104);
nor U21178 (N_21178,N_20041,N_20045);
or U21179 (N_21179,N_19239,N_19961);
nor U21180 (N_21180,N_20341,N_19507);
nor U21181 (N_21181,N_20235,N_19545);
nor U21182 (N_21182,N_20022,N_19523);
and U21183 (N_21183,N_19249,N_19379);
and U21184 (N_21184,N_20350,N_20353);
nor U21185 (N_21185,N_20047,N_20072);
nand U21186 (N_21186,N_20015,N_20098);
and U21187 (N_21187,N_19659,N_20019);
nor U21188 (N_21188,N_19958,N_19538);
xor U21189 (N_21189,N_19908,N_20170);
or U21190 (N_21190,N_19897,N_19497);
nor U21191 (N_21191,N_20074,N_19855);
nand U21192 (N_21192,N_19676,N_19264);
and U21193 (N_21193,N_20145,N_19527);
or U21194 (N_21194,N_19206,N_20221);
and U21195 (N_21195,N_20049,N_19215);
xor U21196 (N_21196,N_20383,N_19746);
or U21197 (N_21197,N_19798,N_20202);
xor U21198 (N_21198,N_20212,N_19693);
or U21199 (N_21199,N_19202,N_19543);
and U21200 (N_21200,N_20345,N_20178);
nor U21201 (N_21201,N_19502,N_19521);
or U21202 (N_21202,N_20219,N_20387);
nor U21203 (N_21203,N_19632,N_20206);
nand U21204 (N_21204,N_19436,N_20140);
or U21205 (N_21205,N_19214,N_19524);
or U21206 (N_21206,N_19773,N_20360);
or U21207 (N_21207,N_20221,N_19654);
nand U21208 (N_21208,N_19255,N_19991);
nor U21209 (N_21209,N_19864,N_20146);
or U21210 (N_21210,N_19576,N_19797);
or U21211 (N_21211,N_19465,N_20148);
or U21212 (N_21212,N_20187,N_20176);
nand U21213 (N_21213,N_19269,N_19747);
xnor U21214 (N_21214,N_19268,N_20198);
nor U21215 (N_21215,N_20177,N_19913);
or U21216 (N_21216,N_20060,N_20202);
or U21217 (N_21217,N_19675,N_20348);
nand U21218 (N_21218,N_19240,N_20293);
nand U21219 (N_21219,N_19986,N_19358);
xnor U21220 (N_21220,N_20084,N_20129);
xnor U21221 (N_21221,N_20140,N_20345);
nand U21222 (N_21222,N_20028,N_19514);
nor U21223 (N_21223,N_20039,N_19248);
nand U21224 (N_21224,N_19773,N_19516);
or U21225 (N_21225,N_20286,N_20399);
or U21226 (N_21226,N_20275,N_19321);
or U21227 (N_21227,N_20194,N_19450);
nand U21228 (N_21228,N_19514,N_20366);
nor U21229 (N_21229,N_20220,N_20334);
or U21230 (N_21230,N_19227,N_19527);
or U21231 (N_21231,N_19929,N_19234);
and U21232 (N_21232,N_19290,N_19873);
and U21233 (N_21233,N_19313,N_20046);
nor U21234 (N_21234,N_19286,N_19916);
xor U21235 (N_21235,N_19351,N_19480);
nor U21236 (N_21236,N_19792,N_19265);
nor U21237 (N_21237,N_19422,N_19425);
nor U21238 (N_21238,N_20389,N_19878);
nand U21239 (N_21239,N_20125,N_20203);
nor U21240 (N_21240,N_19462,N_20073);
nor U21241 (N_21241,N_19462,N_20281);
xor U21242 (N_21242,N_20277,N_19292);
xnor U21243 (N_21243,N_19436,N_19325);
xor U21244 (N_21244,N_19736,N_19372);
or U21245 (N_21245,N_20226,N_19702);
xor U21246 (N_21246,N_20120,N_19586);
nand U21247 (N_21247,N_19602,N_19759);
nor U21248 (N_21248,N_19400,N_19434);
xnor U21249 (N_21249,N_20189,N_19219);
and U21250 (N_21250,N_19487,N_20346);
nor U21251 (N_21251,N_19212,N_20058);
xnor U21252 (N_21252,N_19748,N_19552);
xnor U21253 (N_21253,N_19788,N_20145);
xor U21254 (N_21254,N_20382,N_19968);
xor U21255 (N_21255,N_19654,N_19680);
or U21256 (N_21256,N_19248,N_19933);
nand U21257 (N_21257,N_20190,N_19694);
nor U21258 (N_21258,N_20215,N_20311);
nand U21259 (N_21259,N_20294,N_19588);
nand U21260 (N_21260,N_19479,N_19966);
or U21261 (N_21261,N_20380,N_20048);
or U21262 (N_21262,N_20275,N_20155);
xor U21263 (N_21263,N_19590,N_19390);
xor U21264 (N_21264,N_19601,N_19692);
and U21265 (N_21265,N_20330,N_20395);
or U21266 (N_21266,N_19397,N_19411);
nand U21267 (N_21267,N_19929,N_19439);
and U21268 (N_21268,N_20155,N_19324);
xnor U21269 (N_21269,N_19200,N_19803);
and U21270 (N_21270,N_19276,N_19795);
xor U21271 (N_21271,N_19838,N_19730);
nand U21272 (N_21272,N_19750,N_20247);
nor U21273 (N_21273,N_19380,N_20226);
or U21274 (N_21274,N_20332,N_20013);
nor U21275 (N_21275,N_20133,N_19543);
or U21276 (N_21276,N_20331,N_19309);
nor U21277 (N_21277,N_19556,N_19580);
nand U21278 (N_21278,N_19877,N_19903);
or U21279 (N_21279,N_20361,N_20026);
xnor U21280 (N_21280,N_19812,N_20307);
nand U21281 (N_21281,N_20080,N_19424);
and U21282 (N_21282,N_19726,N_19927);
xnor U21283 (N_21283,N_19510,N_19520);
nand U21284 (N_21284,N_20128,N_19535);
or U21285 (N_21285,N_19960,N_20075);
or U21286 (N_21286,N_20308,N_19409);
nand U21287 (N_21287,N_19486,N_20333);
nand U21288 (N_21288,N_19840,N_20000);
nand U21289 (N_21289,N_19816,N_19389);
nand U21290 (N_21290,N_19831,N_20030);
xnor U21291 (N_21291,N_19442,N_19971);
nor U21292 (N_21292,N_20051,N_19567);
xor U21293 (N_21293,N_20276,N_19377);
nand U21294 (N_21294,N_20356,N_20336);
nand U21295 (N_21295,N_20330,N_20028);
xnor U21296 (N_21296,N_20150,N_20149);
and U21297 (N_21297,N_19501,N_20008);
xnor U21298 (N_21298,N_20035,N_19844);
and U21299 (N_21299,N_19720,N_20137);
xor U21300 (N_21300,N_19361,N_19912);
nand U21301 (N_21301,N_19617,N_19754);
xor U21302 (N_21302,N_19444,N_19265);
nor U21303 (N_21303,N_20254,N_19447);
nor U21304 (N_21304,N_19886,N_19862);
nand U21305 (N_21305,N_19605,N_19731);
and U21306 (N_21306,N_19219,N_19498);
nand U21307 (N_21307,N_20315,N_19693);
and U21308 (N_21308,N_19711,N_19426);
xnor U21309 (N_21309,N_19311,N_19489);
and U21310 (N_21310,N_19964,N_19240);
nor U21311 (N_21311,N_19394,N_20172);
or U21312 (N_21312,N_20244,N_20001);
nand U21313 (N_21313,N_20373,N_19969);
or U21314 (N_21314,N_19677,N_20338);
or U21315 (N_21315,N_19213,N_20120);
xor U21316 (N_21316,N_19919,N_19482);
or U21317 (N_21317,N_19612,N_20184);
or U21318 (N_21318,N_20350,N_19534);
nand U21319 (N_21319,N_19235,N_19918);
or U21320 (N_21320,N_19314,N_19341);
or U21321 (N_21321,N_19476,N_20356);
nor U21322 (N_21322,N_20332,N_20186);
and U21323 (N_21323,N_19765,N_20261);
and U21324 (N_21324,N_19977,N_19992);
xor U21325 (N_21325,N_19356,N_20228);
and U21326 (N_21326,N_20367,N_19218);
or U21327 (N_21327,N_20308,N_20270);
and U21328 (N_21328,N_19783,N_19867);
or U21329 (N_21329,N_19797,N_20119);
nor U21330 (N_21330,N_19477,N_20137);
or U21331 (N_21331,N_20301,N_20121);
nor U21332 (N_21332,N_19229,N_20395);
nand U21333 (N_21333,N_19232,N_19828);
or U21334 (N_21334,N_19665,N_20328);
nor U21335 (N_21335,N_20063,N_19805);
nor U21336 (N_21336,N_19714,N_20059);
nand U21337 (N_21337,N_20156,N_20025);
nor U21338 (N_21338,N_19416,N_20208);
and U21339 (N_21339,N_19691,N_19372);
or U21340 (N_21340,N_19398,N_19713);
nand U21341 (N_21341,N_19616,N_19700);
nor U21342 (N_21342,N_19412,N_19598);
and U21343 (N_21343,N_19280,N_20278);
xor U21344 (N_21344,N_20256,N_20049);
or U21345 (N_21345,N_20229,N_19266);
and U21346 (N_21346,N_19942,N_20240);
nor U21347 (N_21347,N_19776,N_19249);
nand U21348 (N_21348,N_19599,N_19236);
xor U21349 (N_21349,N_19639,N_19721);
nor U21350 (N_21350,N_19528,N_19678);
or U21351 (N_21351,N_19875,N_19975);
nor U21352 (N_21352,N_19248,N_19307);
xnor U21353 (N_21353,N_19361,N_19698);
xnor U21354 (N_21354,N_19245,N_19864);
nand U21355 (N_21355,N_19313,N_20103);
or U21356 (N_21356,N_19444,N_19388);
nor U21357 (N_21357,N_19551,N_19544);
or U21358 (N_21358,N_20190,N_20359);
nor U21359 (N_21359,N_20374,N_20301);
xor U21360 (N_21360,N_20363,N_19517);
and U21361 (N_21361,N_20071,N_19257);
or U21362 (N_21362,N_19300,N_19239);
and U21363 (N_21363,N_19212,N_19262);
nand U21364 (N_21364,N_19860,N_19893);
nor U21365 (N_21365,N_19855,N_19544);
or U21366 (N_21366,N_20122,N_20263);
and U21367 (N_21367,N_19674,N_20188);
xnor U21368 (N_21368,N_19310,N_19252);
or U21369 (N_21369,N_20319,N_20378);
or U21370 (N_21370,N_19953,N_19758);
nand U21371 (N_21371,N_20015,N_20170);
xor U21372 (N_21372,N_19741,N_20095);
and U21373 (N_21373,N_19654,N_19690);
and U21374 (N_21374,N_19512,N_19909);
and U21375 (N_21375,N_19515,N_19583);
and U21376 (N_21376,N_19817,N_20095);
and U21377 (N_21377,N_19327,N_19924);
nor U21378 (N_21378,N_19352,N_19895);
nor U21379 (N_21379,N_20348,N_19838);
or U21380 (N_21380,N_20147,N_19804);
or U21381 (N_21381,N_19331,N_19287);
or U21382 (N_21382,N_19863,N_20094);
and U21383 (N_21383,N_19662,N_19632);
xor U21384 (N_21384,N_20109,N_20272);
or U21385 (N_21385,N_19447,N_19535);
and U21386 (N_21386,N_20344,N_19747);
or U21387 (N_21387,N_19977,N_19638);
nand U21388 (N_21388,N_20099,N_20003);
nor U21389 (N_21389,N_19799,N_19938);
nand U21390 (N_21390,N_19995,N_19723);
or U21391 (N_21391,N_20042,N_19991);
xor U21392 (N_21392,N_20331,N_19447);
or U21393 (N_21393,N_19819,N_19270);
nand U21394 (N_21394,N_20380,N_20298);
nand U21395 (N_21395,N_19242,N_19517);
nor U21396 (N_21396,N_19772,N_20002);
and U21397 (N_21397,N_19913,N_20346);
or U21398 (N_21398,N_19830,N_19569);
and U21399 (N_21399,N_19488,N_20145);
or U21400 (N_21400,N_19687,N_19585);
nand U21401 (N_21401,N_20334,N_19593);
nor U21402 (N_21402,N_19750,N_19448);
xnor U21403 (N_21403,N_19391,N_19279);
and U21404 (N_21404,N_20170,N_19559);
nand U21405 (N_21405,N_20229,N_19800);
or U21406 (N_21406,N_20380,N_19726);
and U21407 (N_21407,N_19231,N_19427);
nand U21408 (N_21408,N_19372,N_20149);
xnor U21409 (N_21409,N_19870,N_19589);
xnor U21410 (N_21410,N_20290,N_20006);
and U21411 (N_21411,N_19999,N_19649);
and U21412 (N_21412,N_19571,N_19727);
and U21413 (N_21413,N_20022,N_20035);
nand U21414 (N_21414,N_19423,N_19739);
or U21415 (N_21415,N_19233,N_20124);
and U21416 (N_21416,N_19662,N_19804);
xnor U21417 (N_21417,N_19410,N_19396);
and U21418 (N_21418,N_19361,N_20366);
or U21419 (N_21419,N_19540,N_20195);
nor U21420 (N_21420,N_19719,N_20167);
nand U21421 (N_21421,N_19315,N_19327);
or U21422 (N_21422,N_19658,N_19425);
nor U21423 (N_21423,N_19302,N_19475);
or U21424 (N_21424,N_19810,N_19297);
nand U21425 (N_21425,N_20160,N_19974);
and U21426 (N_21426,N_19430,N_20098);
and U21427 (N_21427,N_20247,N_20252);
nand U21428 (N_21428,N_20339,N_19696);
or U21429 (N_21429,N_20055,N_19898);
nand U21430 (N_21430,N_19303,N_19432);
nand U21431 (N_21431,N_20180,N_19563);
xnor U21432 (N_21432,N_20368,N_19573);
xor U21433 (N_21433,N_19828,N_19978);
and U21434 (N_21434,N_19579,N_20283);
and U21435 (N_21435,N_19758,N_19858);
xor U21436 (N_21436,N_19735,N_19324);
or U21437 (N_21437,N_19961,N_19959);
nor U21438 (N_21438,N_19406,N_20086);
nor U21439 (N_21439,N_19817,N_19220);
xor U21440 (N_21440,N_19644,N_19468);
or U21441 (N_21441,N_20216,N_19630);
nor U21442 (N_21442,N_20287,N_19299);
xnor U21443 (N_21443,N_19522,N_19349);
and U21444 (N_21444,N_20066,N_19696);
xnor U21445 (N_21445,N_19922,N_19343);
nor U21446 (N_21446,N_19390,N_20259);
and U21447 (N_21447,N_19688,N_20204);
or U21448 (N_21448,N_19846,N_19278);
and U21449 (N_21449,N_19891,N_19570);
nor U21450 (N_21450,N_20254,N_19211);
or U21451 (N_21451,N_19315,N_19819);
nand U21452 (N_21452,N_19657,N_19845);
and U21453 (N_21453,N_20228,N_19636);
or U21454 (N_21454,N_20186,N_20052);
xor U21455 (N_21455,N_20211,N_20060);
nor U21456 (N_21456,N_19386,N_19358);
or U21457 (N_21457,N_19839,N_20334);
nand U21458 (N_21458,N_20321,N_19330);
or U21459 (N_21459,N_19975,N_19216);
or U21460 (N_21460,N_19882,N_19411);
xor U21461 (N_21461,N_19402,N_19333);
xor U21462 (N_21462,N_19830,N_20232);
and U21463 (N_21463,N_19856,N_20377);
and U21464 (N_21464,N_19731,N_19849);
or U21465 (N_21465,N_19381,N_19683);
and U21466 (N_21466,N_19721,N_19288);
nand U21467 (N_21467,N_20060,N_19416);
nor U21468 (N_21468,N_19661,N_20140);
nor U21469 (N_21469,N_19378,N_20161);
xnor U21470 (N_21470,N_19302,N_19978);
nand U21471 (N_21471,N_19598,N_19943);
xor U21472 (N_21472,N_20352,N_19806);
nand U21473 (N_21473,N_19948,N_19989);
and U21474 (N_21474,N_19898,N_20029);
xnor U21475 (N_21475,N_19595,N_19542);
or U21476 (N_21476,N_19844,N_19240);
nand U21477 (N_21477,N_20315,N_20349);
or U21478 (N_21478,N_19479,N_20038);
or U21479 (N_21479,N_20369,N_19370);
xnor U21480 (N_21480,N_19520,N_19421);
or U21481 (N_21481,N_20148,N_20091);
or U21482 (N_21482,N_19889,N_20338);
or U21483 (N_21483,N_20346,N_19300);
or U21484 (N_21484,N_19438,N_19808);
and U21485 (N_21485,N_19690,N_19691);
nor U21486 (N_21486,N_19468,N_20365);
xnor U21487 (N_21487,N_19347,N_19307);
and U21488 (N_21488,N_19902,N_19835);
xnor U21489 (N_21489,N_19521,N_20075);
nor U21490 (N_21490,N_19726,N_19628);
nor U21491 (N_21491,N_19996,N_19407);
nor U21492 (N_21492,N_19465,N_19582);
nand U21493 (N_21493,N_19818,N_20393);
nor U21494 (N_21494,N_19407,N_19529);
nor U21495 (N_21495,N_19680,N_19293);
xor U21496 (N_21496,N_19557,N_20305);
xnor U21497 (N_21497,N_19901,N_19557);
nor U21498 (N_21498,N_19472,N_20314);
xnor U21499 (N_21499,N_20082,N_19757);
and U21500 (N_21500,N_19922,N_19848);
xor U21501 (N_21501,N_19231,N_19235);
nor U21502 (N_21502,N_20207,N_20079);
nor U21503 (N_21503,N_20081,N_19565);
or U21504 (N_21504,N_19632,N_20298);
and U21505 (N_21505,N_19843,N_19933);
and U21506 (N_21506,N_20203,N_19566);
nor U21507 (N_21507,N_19737,N_19789);
and U21508 (N_21508,N_19639,N_20070);
nor U21509 (N_21509,N_19529,N_20254);
nand U21510 (N_21510,N_19560,N_20171);
xor U21511 (N_21511,N_19756,N_20171);
xor U21512 (N_21512,N_20122,N_19852);
nor U21513 (N_21513,N_19621,N_19805);
nand U21514 (N_21514,N_19213,N_20105);
xor U21515 (N_21515,N_19806,N_20387);
nand U21516 (N_21516,N_20210,N_19229);
or U21517 (N_21517,N_19565,N_19929);
nor U21518 (N_21518,N_20259,N_19876);
and U21519 (N_21519,N_19444,N_19571);
nand U21520 (N_21520,N_19596,N_19813);
nor U21521 (N_21521,N_19546,N_19817);
xor U21522 (N_21522,N_19475,N_19851);
nor U21523 (N_21523,N_19333,N_20217);
or U21524 (N_21524,N_20160,N_19366);
nand U21525 (N_21525,N_20065,N_20152);
xnor U21526 (N_21526,N_19219,N_19669);
nand U21527 (N_21527,N_19719,N_19286);
or U21528 (N_21528,N_19699,N_19911);
nor U21529 (N_21529,N_20332,N_20248);
nand U21530 (N_21530,N_19881,N_20298);
and U21531 (N_21531,N_20137,N_19701);
nand U21532 (N_21532,N_19285,N_20099);
nor U21533 (N_21533,N_19725,N_20258);
nor U21534 (N_21534,N_19706,N_19817);
xor U21535 (N_21535,N_20117,N_19668);
nand U21536 (N_21536,N_19460,N_19487);
nand U21537 (N_21537,N_19294,N_19518);
or U21538 (N_21538,N_19489,N_20059);
xnor U21539 (N_21539,N_19673,N_19757);
xnor U21540 (N_21540,N_20338,N_20255);
nand U21541 (N_21541,N_19634,N_19505);
nand U21542 (N_21542,N_19501,N_20183);
nand U21543 (N_21543,N_19482,N_19684);
and U21544 (N_21544,N_19734,N_19252);
and U21545 (N_21545,N_19589,N_19541);
or U21546 (N_21546,N_20190,N_19875);
nand U21547 (N_21547,N_19795,N_20206);
and U21548 (N_21548,N_19944,N_19863);
and U21549 (N_21549,N_19457,N_20132);
nand U21550 (N_21550,N_19810,N_19427);
nand U21551 (N_21551,N_19612,N_20369);
xnor U21552 (N_21552,N_19262,N_20332);
and U21553 (N_21553,N_19548,N_19460);
nor U21554 (N_21554,N_19490,N_20083);
or U21555 (N_21555,N_20309,N_20366);
nand U21556 (N_21556,N_19435,N_20131);
and U21557 (N_21557,N_19360,N_19609);
and U21558 (N_21558,N_19697,N_19787);
and U21559 (N_21559,N_20312,N_19726);
and U21560 (N_21560,N_19779,N_19571);
and U21561 (N_21561,N_19410,N_19789);
nor U21562 (N_21562,N_20011,N_19983);
or U21563 (N_21563,N_19705,N_20177);
nor U21564 (N_21564,N_19523,N_19422);
or U21565 (N_21565,N_20323,N_19976);
or U21566 (N_21566,N_19575,N_19296);
nand U21567 (N_21567,N_19815,N_19759);
xnor U21568 (N_21568,N_19652,N_20352);
or U21569 (N_21569,N_19359,N_19769);
and U21570 (N_21570,N_19871,N_19541);
and U21571 (N_21571,N_19406,N_19521);
nand U21572 (N_21572,N_20140,N_20126);
nor U21573 (N_21573,N_20230,N_19215);
and U21574 (N_21574,N_19584,N_19232);
or U21575 (N_21575,N_20162,N_19729);
nand U21576 (N_21576,N_19673,N_19638);
or U21577 (N_21577,N_20226,N_19622);
nor U21578 (N_21578,N_19820,N_19681);
nor U21579 (N_21579,N_20152,N_20031);
nand U21580 (N_21580,N_19342,N_19519);
xor U21581 (N_21581,N_19987,N_20065);
nand U21582 (N_21582,N_20005,N_20216);
or U21583 (N_21583,N_19472,N_19527);
nor U21584 (N_21584,N_19969,N_19830);
nand U21585 (N_21585,N_19808,N_20186);
or U21586 (N_21586,N_19801,N_20250);
and U21587 (N_21587,N_19682,N_20345);
and U21588 (N_21588,N_20005,N_19467);
nand U21589 (N_21589,N_19263,N_19264);
nor U21590 (N_21590,N_20398,N_20372);
nor U21591 (N_21591,N_19454,N_19437);
and U21592 (N_21592,N_19970,N_19266);
or U21593 (N_21593,N_19437,N_19421);
nor U21594 (N_21594,N_19432,N_19403);
or U21595 (N_21595,N_19739,N_20037);
or U21596 (N_21596,N_19866,N_19735);
and U21597 (N_21597,N_19739,N_19940);
or U21598 (N_21598,N_19921,N_19360);
and U21599 (N_21599,N_19427,N_20142);
nor U21600 (N_21600,N_20924,N_20507);
nor U21601 (N_21601,N_20447,N_21583);
or U21602 (N_21602,N_21344,N_20598);
nor U21603 (N_21603,N_21129,N_21315);
and U21604 (N_21604,N_21537,N_21377);
nor U21605 (N_21605,N_20783,N_21272);
or U21606 (N_21606,N_20891,N_20990);
nand U21607 (N_21607,N_21380,N_21440);
and U21608 (N_21608,N_20982,N_20492);
and U21609 (N_21609,N_21200,N_21280);
nand U21610 (N_21610,N_21423,N_21420);
or U21611 (N_21611,N_20499,N_20880);
xnor U21612 (N_21612,N_21564,N_20996);
and U21613 (N_21613,N_21114,N_21293);
and U21614 (N_21614,N_20861,N_20953);
xnor U21615 (N_21615,N_20585,N_21356);
nand U21616 (N_21616,N_20890,N_20976);
and U21617 (N_21617,N_21333,N_21290);
nand U21618 (N_21618,N_21439,N_21268);
nor U21619 (N_21619,N_20883,N_21163);
xnor U21620 (N_21620,N_21015,N_20548);
nor U21621 (N_21621,N_21234,N_20804);
or U21622 (N_21622,N_21236,N_21563);
xor U21623 (N_21623,N_21229,N_20592);
xnor U21624 (N_21624,N_20416,N_21257);
and U21625 (N_21625,N_20852,N_20858);
and U21626 (N_21626,N_21567,N_20420);
or U21627 (N_21627,N_21018,N_21365);
xor U21628 (N_21628,N_21287,N_21297);
and U21629 (N_21629,N_21566,N_21156);
or U21630 (N_21630,N_21582,N_20840);
nand U21631 (N_21631,N_21039,N_20938);
nand U21632 (N_21632,N_20910,N_21006);
nor U21633 (N_21633,N_20856,N_21128);
xor U21634 (N_21634,N_20793,N_20828);
xnor U21635 (N_21635,N_20564,N_20954);
nand U21636 (N_21636,N_20699,N_20668);
xnor U21637 (N_21637,N_20784,N_20693);
nor U21638 (N_21638,N_21349,N_20791);
nor U21639 (N_21639,N_21430,N_20407);
nand U21640 (N_21640,N_21573,N_20415);
nor U21641 (N_21641,N_20503,N_21581);
nand U21642 (N_21642,N_20696,N_20824);
and U21643 (N_21643,N_20772,N_21598);
and U21644 (N_21644,N_21165,N_20899);
nand U21645 (N_21645,N_20554,N_20452);
and U21646 (N_21646,N_21000,N_20808);
nor U21647 (N_21647,N_21080,N_20849);
xnor U21648 (N_21648,N_20848,N_21134);
xor U21649 (N_21649,N_20871,N_21035);
and U21650 (N_21650,N_21104,N_21081);
or U21651 (N_21651,N_21556,N_21189);
xor U21652 (N_21652,N_20587,N_21231);
or U21653 (N_21653,N_20786,N_21249);
xnor U21654 (N_21654,N_21584,N_20866);
nor U21655 (N_21655,N_21352,N_20992);
nand U21656 (N_21656,N_21414,N_21314);
or U21657 (N_21657,N_20664,N_20843);
or U21658 (N_21658,N_20835,N_20624);
nand U21659 (N_21659,N_20588,N_21585);
nand U21660 (N_21660,N_21071,N_21417);
nand U21661 (N_21661,N_21144,N_20497);
nand U21662 (N_21662,N_20544,N_20937);
and U21663 (N_21663,N_20448,N_21111);
nor U21664 (N_21664,N_20568,N_21458);
nor U21665 (N_21665,N_21174,N_21248);
and U21666 (N_21666,N_21456,N_21025);
nor U21667 (N_21667,N_20483,N_21316);
nand U21668 (N_21668,N_21321,N_21118);
nor U21669 (N_21669,N_20961,N_20545);
xnor U21670 (N_21670,N_21577,N_21510);
xor U21671 (N_21671,N_21554,N_21301);
xor U21672 (N_21672,N_20658,N_21469);
nor U21673 (N_21673,N_20977,N_21481);
xor U21674 (N_21674,N_21305,N_20831);
or U21675 (N_21675,N_20517,N_21310);
and U21676 (N_21676,N_20642,N_20667);
or U21677 (N_21677,N_20472,N_20680);
or U21678 (N_21678,N_20757,N_20596);
and U21679 (N_21679,N_21482,N_20951);
or U21680 (N_21680,N_20643,N_20557);
xor U21681 (N_21681,N_20782,N_20901);
and U21682 (N_21682,N_20916,N_21507);
xor U21683 (N_21683,N_21485,N_20809);
or U21684 (N_21684,N_21531,N_21191);
xnor U21685 (N_21685,N_20906,N_20582);
nor U21686 (N_21686,N_20607,N_21056);
and U21687 (N_21687,N_20788,N_21106);
nand U21688 (N_21688,N_21141,N_20747);
and U21689 (N_21689,N_21394,N_21124);
and U21690 (N_21690,N_20688,N_21411);
xor U21691 (N_21691,N_20986,N_20662);
and U21692 (N_21692,N_21100,N_21176);
or U21693 (N_21693,N_20762,N_21175);
xor U21694 (N_21694,N_20549,N_21395);
nor U21695 (N_21695,N_20579,N_21426);
or U21696 (N_21696,N_21451,N_20623);
nand U21697 (N_21697,N_20413,N_20820);
and U21698 (N_21698,N_20745,N_20956);
nor U21699 (N_21699,N_20758,N_20781);
nand U21700 (N_21700,N_20601,N_21233);
nand U21701 (N_21701,N_21361,N_21286);
nor U21702 (N_21702,N_20653,N_21568);
xor U21703 (N_21703,N_21433,N_20690);
nand U21704 (N_21704,N_21328,N_20525);
and U21705 (N_21705,N_20462,N_20622);
nor U21706 (N_21706,N_21218,N_20473);
xnor U21707 (N_21707,N_20754,N_20520);
xnor U21708 (N_21708,N_20755,N_21126);
or U21709 (N_21709,N_20508,N_20519);
nand U21710 (N_21710,N_20586,N_21196);
nor U21711 (N_21711,N_20775,N_21224);
nor U21712 (N_21712,N_20812,N_20567);
or U21713 (N_21713,N_20842,N_20742);
nor U21714 (N_21714,N_21495,N_20423);
nand U21715 (N_21715,N_20947,N_20444);
xor U21716 (N_21716,N_21214,N_21169);
xnor U21717 (N_21717,N_21159,N_21192);
and U21718 (N_21718,N_21232,N_20457);
or U21719 (N_21719,N_20862,N_20735);
and U21720 (N_21720,N_21278,N_21235);
and U21721 (N_21721,N_21487,N_21279);
nor U21722 (N_21722,N_21535,N_21382);
or U21723 (N_21723,N_20608,N_21548);
or U21724 (N_21724,N_20709,N_20576);
xor U21725 (N_21725,N_20966,N_20649);
xor U21726 (N_21726,N_21143,N_20569);
xnor U21727 (N_21727,N_20562,N_20753);
xor U21728 (N_21728,N_21166,N_20454);
or U21729 (N_21729,N_20614,N_20633);
nor U21730 (N_21730,N_21557,N_20750);
or U21731 (N_21731,N_21358,N_21504);
xor U21732 (N_21732,N_20737,N_20510);
and U21733 (N_21733,N_21521,N_20615);
and U21734 (N_21734,N_20634,N_20641);
and U21735 (N_21735,N_20559,N_21202);
xnor U21736 (N_21736,N_20723,N_21449);
xor U21737 (N_21737,N_20540,N_20619);
or U21738 (N_21738,N_20532,N_21139);
xnor U21739 (N_21739,N_20773,N_20401);
nand U21740 (N_21740,N_21147,N_21092);
xnor U21741 (N_21741,N_20629,N_21405);
nor U21742 (N_21742,N_21309,N_21273);
nand U21743 (N_21743,N_20713,N_20731);
nand U21744 (N_21744,N_20580,N_21101);
nor U21745 (N_21745,N_20893,N_21313);
nor U21746 (N_21746,N_20656,N_21589);
and U21747 (N_21747,N_20402,N_21421);
nand U21748 (N_21748,N_20612,N_20962);
or U21749 (N_21749,N_20975,N_20743);
xnor U21750 (N_21750,N_20868,N_21161);
xor U21751 (N_21751,N_21371,N_20513);
nand U21752 (N_21752,N_20518,N_20541);
and U21753 (N_21753,N_20985,N_20853);
nor U21754 (N_21754,N_21325,N_20787);
nor U21755 (N_21755,N_21401,N_21150);
nor U21756 (N_21756,N_21067,N_21076);
and U21757 (N_21757,N_20543,N_21447);
nand U21758 (N_21758,N_21523,N_21289);
and U21759 (N_21759,N_20646,N_20964);
nand U21760 (N_21760,N_20974,N_21070);
or U21761 (N_21761,N_20669,N_21024);
and U21762 (N_21762,N_20878,N_21354);
or U21763 (N_21763,N_21491,N_20636);
xnor U21764 (N_21764,N_20570,N_21442);
xnor U21765 (N_21765,N_20529,N_21259);
or U21766 (N_21766,N_20896,N_20488);
nand U21767 (N_21767,N_20480,N_21553);
or U21768 (N_21768,N_20660,N_21501);
nor U21769 (N_21769,N_21308,N_21167);
or U21770 (N_21770,N_20770,N_20800);
nand U21771 (N_21771,N_21274,N_21351);
and U21772 (N_21772,N_21069,N_21335);
xor U21773 (N_21773,N_21240,N_20704);
and U21774 (N_21774,N_20494,N_21342);
and U21775 (N_21775,N_20616,N_20918);
nor U21776 (N_21776,N_20412,N_21043);
nand U21777 (N_21777,N_20957,N_21580);
nand U21778 (N_21778,N_20493,N_20771);
nor U21779 (N_21779,N_21061,N_20744);
nor U21780 (N_21780,N_20600,N_21552);
xnor U21781 (N_21781,N_21270,N_20888);
nand U21782 (N_21782,N_20522,N_21016);
nor U21783 (N_21783,N_21304,N_21120);
and U21784 (N_21784,N_20434,N_21110);
xor U21785 (N_21785,N_21475,N_20620);
nor U21786 (N_21786,N_21441,N_21045);
nor U21787 (N_21787,N_20955,N_20645);
xor U21788 (N_21788,N_21511,N_20748);
and U21789 (N_21789,N_21152,N_21164);
nor U21790 (N_21790,N_21532,N_21222);
xnor U21791 (N_21791,N_21393,N_21296);
and U21792 (N_21792,N_21539,N_21370);
and U21793 (N_21793,N_21346,N_21422);
xor U21794 (N_21794,N_20897,N_21484);
nand U21795 (N_21795,N_21415,N_21538);
nor U21796 (N_21796,N_20941,N_20952);
nor U21797 (N_21797,N_21123,N_21571);
xnor U21798 (N_21798,N_21561,N_21022);
nor U21799 (N_21799,N_20714,N_21020);
nand U21800 (N_21800,N_20971,N_20440);
xor U21801 (N_21801,N_20767,N_21528);
nor U21802 (N_21802,N_21054,N_20829);
nand U21803 (N_21803,N_21284,N_20983);
or U21804 (N_21804,N_21107,N_21464);
and U21805 (N_21805,N_20637,N_20822);
or U21806 (N_21806,N_21466,N_21432);
and U21807 (N_21807,N_20882,N_20761);
nor U21808 (N_21808,N_20606,N_20987);
or U21809 (N_21809,N_21059,N_20441);
nor U21810 (N_21810,N_20575,N_20591);
nand U21811 (N_21811,N_21350,N_20546);
nor U21812 (N_21812,N_20769,N_20451);
xnor U21813 (N_21813,N_20823,N_20836);
nor U21814 (N_21814,N_21385,N_20915);
nor U21815 (N_21815,N_20491,N_21399);
xor U21816 (N_21816,N_20967,N_20886);
xor U21817 (N_21817,N_20721,N_20655);
nand U21818 (N_21818,N_21245,N_20610);
nor U21819 (N_21819,N_21319,N_21148);
or U21820 (N_21820,N_20832,N_20703);
and U21821 (N_21821,N_20722,N_20930);
xnor U21822 (N_21822,N_21149,N_20602);
nand U21823 (N_21823,N_21033,N_20551);
nor U21824 (N_21824,N_21513,N_20411);
nand U21825 (N_21825,N_21404,N_21254);
nand U21826 (N_21826,N_20706,N_21190);
and U21827 (N_21827,N_21265,N_20902);
nor U21828 (N_21828,N_21586,N_21434);
xor U21829 (N_21829,N_21095,N_20613);
nand U21830 (N_21830,N_20926,N_20827);
xnor U21831 (N_21831,N_21560,N_20617);
nand U21832 (N_21832,N_21140,N_20741);
xor U21833 (N_21833,N_21355,N_21001);
and U21834 (N_21834,N_21221,N_20657);
or U21835 (N_21835,N_20443,N_21443);
and U21836 (N_21836,N_20611,N_20702);
xor U21837 (N_21837,N_21238,N_21195);
and U21838 (N_21838,N_20864,N_20467);
nor U21839 (N_21839,N_20521,N_20959);
nand U21840 (N_21840,N_21072,N_21386);
xnor U21841 (N_21841,N_21010,N_20675);
or U21842 (N_21842,N_21406,N_20919);
nor U21843 (N_21843,N_21089,N_20571);
and U21844 (N_21844,N_21299,N_20536);
xnor U21845 (N_21845,N_21223,N_21294);
xnor U21846 (N_21846,N_20523,N_21283);
or U21847 (N_21847,N_21051,N_20663);
nand U21848 (N_21848,N_20738,N_20449);
and U21849 (N_21849,N_21127,N_20765);
nor U21850 (N_21850,N_20464,N_20875);
or U21851 (N_21851,N_21593,N_21468);
xnor U21852 (N_21852,N_21208,N_20635);
xnor U21853 (N_21853,N_21306,N_21211);
xnor U21854 (N_21854,N_20945,N_21457);
or U21855 (N_21855,N_21239,N_20739);
nand U21856 (N_21856,N_21569,N_20695);
xor U21857 (N_21857,N_21478,N_21063);
nor U21858 (N_21858,N_20980,N_21210);
xor U21859 (N_21859,N_21558,N_20505);
or U21860 (N_21860,N_21392,N_21594);
nor U21861 (N_21861,N_21038,N_21027);
xor U21862 (N_21862,N_21098,N_20685);
xnor U21863 (N_21863,N_21499,N_20700);
xor U21864 (N_21864,N_21138,N_20826);
and U21865 (N_21865,N_21336,N_21271);
nand U21866 (N_21866,N_21282,N_21121);
nand U21867 (N_21867,N_20806,N_20870);
and U21868 (N_21868,N_21023,N_20736);
xnor U21869 (N_21869,N_21550,N_21137);
nor U21870 (N_21870,N_21261,N_21146);
or U21871 (N_21871,N_21360,N_20979);
and U21872 (N_21872,N_21509,N_20430);
nand U21873 (N_21873,N_21402,N_20710);
and U21874 (N_21874,N_20830,N_20504);
and U21875 (N_21875,N_21040,N_21494);
and U21876 (N_21876,N_21409,N_20970);
or U21877 (N_21877,N_21498,N_21267);
nor U21878 (N_21878,N_21389,N_21186);
and U21879 (N_21879,N_20889,N_20458);
xor U21880 (N_21880,N_21122,N_20652);
nor U21881 (N_21881,N_21135,N_21307);
xor U21882 (N_21882,N_21256,N_20450);
xnor U21883 (N_21883,N_20950,N_21330);
and U21884 (N_21884,N_21591,N_20644);
and U21885 (N_21885,N_21005,N_21543);
nand U21886 (N_21886,N_21317,N_21332);
nor U21887 (N_21887,N_21046,N_20500);
or U21888 (N_21888,N_20751,N_20526);
nor U21889 (N_21889,N_20679,N_21034);
or U21890 (N_21890,N_21452,N_21064);
and U21891 (N_21891,N_21388,N_21130);
nand U21892 (N_21892,N_20838,N_21347);
nor U21893 (N_21893,N_21206,N_21028);
nand U21894 (N_21894,N_21207,N_21002);
nor U21895 (N_21895,N_20405,N_21396);
nor U21896 (N_21896,N_20716,N_20417);
and U21897 (N_21897,N_21368,N_20419);
or U21898 (N_21898,N_21445,N_21255);
nand U21899 (N_21899,N_21219,N_20999);
xor U21900 (N_21900,N_21158,N_20844);
nor U21901 (N_21901,N_20816,N_21486);
xor U21902 (N_21902,N_20469,N_21082);
and U21903 (N_21903,N_20989,N_20968);
or U21904 (N_21904,N_20475,N_21112);
or U21905 (N_21905,N_20421,N_21201);
nand U21906 (N_21906,N_20682,N_21077);
or U21907 (N_21907,N_21463,N_21269);
and U21908 (N_21908,N_20903,N_20729);
and U21909 (N_21909,N_20426,N_21518);
or U21910 (N_21910,N_21253,N_21400);
xor U21911 (N_21911,N_21467,N_21363);
xnor U21912 (N_21912,N_20509,N_21182);
or U21913 (N_21913,N_21113,N_20776);
and U21914 (N_21914,N_20673,N_20892);
or U21915 (N_21915,N_21508,N_21424);
or U21916 (N_21916,N_21048,N_20931);
xnor U21917 (N_21917,N_20604,N_21057);
and U21918 (N_21918,N_21145,N_21004);
xnor U21919 (N_21919,N_21230,N_20471);
or U21920 (N_21920,N_21226,N_21108);
nand U21921 (N_21921,N_20553,N_21096);
nand U21922 (N_21922,N_21074,N_20609);
or U21923 (N_21923,N_20640,N_20550);
nand U21924 (N_21924,N_21181,N_21185);
or U21925 (N_21925,N_21084,N_20725);
or U21926 (N_21926,N_21212,N_21533);
xnor U21927 (N_21927,N_20466,N_20501);
xnor U21928 (N_21928,N_21073,N_21418);
or U21929 (N_21929,N_21474,N_21055);
or U21930 (N_21930,N_21331,N_20715);
xnor U21931 (N_21931,N_20797,N_20654);
xor U21932 (N_21932,N_20859,N_21320);
or U21933 (N_21933,N_20631,N_20863);
xor U21934 (N_21934,N_21324,N_20468);
and U21935 (N_21935,N_20907,N_21116);
xnor U21936 (N_21936,N_21407,N_21188);
and U21937 (N_21937,N_20678,N_20885);
nor U21938 (N_21938,N_21217,N_20728);
xor U21939 (N_21939,N_20879,N_20825);
or U21940 (N_21940,N_21042,N_20895);
nor U21941 (N_21941,N_20694,N_20445);
or U21942 (N_21942,N_20565,N_20597);
or U21943 (N_21943,N_20939,N_21381);
and U21944 (N_21944,N_21303,N_20860);
nand U21945 (N_21945,N_20911,N_20594);
nor U21946 (N_21946,N_20484,N_20727);
xnor U21947 (N_21947,N_21031,N_21472);
nor U21948 (N_21948,N_21572,N_21369);
and U21949 (N_21949,N_20436,N_20589);
or U21950 (N_21950,N_20406,N_20867);
nand U21951 (N_21951,N_21437,N_21343);
xor U21952 (N_21952,N_21250,N_20659);
nand U21953 (N_21953,N_21258,N_20900);
xnor U21954 (N_21954,N_21285,N_21479);
xor U21955 (N_21955,N_21170,N_21544);
or U21956 (N_21956,N_21011,N_20626);
nor U21957 (N_21957,N_20805,N_20403);
xnor U21958 (N_21958,N_20778,N_20857);
and U21959 (N_21959,N_20763,N_20799);
nor U21960 (N_21960,N_20628,N_21383);
nand U21961 (N_21961,N_20524,N_20512);
xor U21962 (N_21962,N_21471,N_21157);
xnor U21963 (N_21963,N_20946,N_21109);
xnor U21964 (N_21964,N_21075,N_20681);
or U21965 (N_21965,N_20515,N_20921);
xnor U21966 (N_21966,N_21036,N_21446);
nor U21967 (N_21967,N_20834,N_20795);
nand U21968 (N_21968,N_20936,N_20618);
nor U21969 (N_21969,N_20819,N_20650);
xnor U21970 (N_21970,N_21133,N_20697);
xor U21971 (N_21971,N_21246,N_21168);
xnor U21972 (N_21972,N_21247,N_21288);
nand U21973 (N_21973,N_21085,N_21574);
xor U21974 (N_21974,N_21078,N_21505);
or U21975 (N_21975,N_20780,N_20766);
nor U21976 (N_21976,N_21462,N_20807);
or U21977 (N_21977,N_21547,N_20638);
and U21978 (N_21978,N_20677,N_20969);
and U21979 (N_21979,N_21524,N_21416);
or U21980 (N_21980,N_21291,N_21058);
nand U21981 (N_21981,N_21436,N_20574);
xor U21982 (N_21982,N_20691,N_20539);
and U21983 (N_21983,N_21559,N_20425);
xnor U21984 (N_21984,N_21244,N_21052);
and U21985 (N_21985,N_21529,N_20674);
nor U21986 (N_21986,N_21378,N_20942);
or U21987 (N_21987,N_21488,N_21154);
xnor U21988 (N_21988,N_21008,N_21435);
nor U21989 (N_21989,N_20400,N_21493);
xor U21990 (N_21990,N_21527,N_21012);
nor U21991 (N_21991,N_20884,N_21540);
or U21992 (N_21992,N_20414,N_20833);
nand U21993 (N_21993,N_21341,N_20732);
nand U21994 (N_21994,N_20672,N_20726);
and U21995 (N_21995,N_20877,N_20514);
or U21996 (N_21996,N_21490,N_21251);
nor U21997 (N_21997,N_20427,N_20887);
and U21998 (N_21998,N_21007,N_21515);
and U21999 (N_21999,N_20802,N_21546);
and U22000 (N_22000,N_20839,N_21049);
nand U22001 (N_22001,N_21032,N_21391);
nor U22002 (N_22002,N_20639,N_21180);
xor U22003 (N_22003,N_20692,N_20801);
nor U22004 (N_22004,N_20949,N_21506);
and U22005 (N_22005,N_21171,N_20530);
xor U22006 (N_22006,N_21136,N_21298);
nor U22007 (N_22007,N_21119,N_20790);
or U22008 (N_22008,N_20477,N_21534);
nand U22009 (N_22009,N_20837,N_21536);
or U22010 (N_22010,N_21470,N_21013);
nand U22011 (N_22011,N_21337,N_21530);
and U22012 (N_22012,N_20595,N_20984);
nand U22013 (N_22013,N_21338,N_21281);
nand U22014 (N_22014,N_20913,N_20991);
and U22015 (N_22015,N_21520,N_21311);
nand U22016 (N_22016,N_20707,N_20993);
nor U22017 (N_22017,N_21021,N_20978);
xor U22018 (N_22018,N_20577,N_21172);
nor U22019 (N_22019,N_20846,N_21177);
or U22020 (N_22020,N_21359,N_21353);
nand U22021 (N_22021,N_20908,N_21364);
and U22022 (N_22022,N_20470,N_21565);
nor U22023 (N_22023,N_20408,N_21260);
and U22024 (N_22024,N_20433,N_20798);
nand U22025 (N_22025,N_21194,N_20943);
and U22026 (N_22026,N_21179,N_21105);
or U22027 (N_22027,N_20547,N_20777);
xnor U22028 (N_22028,N_21497,N_20581);
nor U22029 (N_22029,N_20914,N_21228);
nor U22030 (N_22030,N_20528,N_21199);
xor U22031 (N_22031,N_20917,N_20905);
nor U22032 (N_22032,N_20719,N_21275);
or U22033 (N_22033,N_21477,N_20404);
nand U22034 (N_22034,N_21215,N_20810);
nand U22035 (N_22035,N_21326,N_20774);
xnor U22036 (N_22036,N_21438,N_20909);
nor U22037 (N_22037,N_20869,N_20817);
nand U22038 (N_22038,N_21576,N_21086);
nor U22039 (N_22039,N_20482,N_20442);
or U22040 (N_22040,N_20734,N_20498);
xor U22041 (N_22041,N_20851,N_20583);
nor U22042 (N_22042,N_20718,N_20534);
xor U22043 (N_22043,N_20760,N_20872);
and U22044 (N_22044,N_21178,N_21397);
nor U22045 (N_22045,N_20409,N_20803);
xor U22046 (N_22046,N_20671,N_21083);
and U22047 (N_22047,N_21184,N_20698);
xor U22048 (N_22048,N_21483,N_20429);
or U22049 (N_22049,N_20684,N_20847);
or U22050 (N_22050,N_20792,N_21318);
and U22051 (N_22051,N_21264,N_21151);
and U22052 (N_22052,N_20927,N_20687);
xor U22053 (N_22053,N_20489,N_20561);
nor U22054 (N_22054,N_20573,N_21429);
nor U22055 (N_22055,N_20537,N_21339);
nor U22056 (N_22056,N_21068,N_21454);
or U22057 (N_22057,N_21496,N_21329);
nand U22058 (N_22058,N_21091,N_20476);
or U22059 (N_22059,N_20527,N_21242);
nand U22060 (N_22060,N_20733,N_21367);
xnor U22061 (N_22061,N_21384,N_21295);
xnor U22062 (N_22062,N_21312,N_21465);
or U22063 (N_22063,N_20593,N_20994);
or U22064 (N_22064,N_21461,N_20932);
nor U22065 (N_22065,N_21448,N_20661);
xnor U22066 (N_22066,N_20486,N_20625);
or U22067 (N_22067,N_21160,N_21183);
nor U22068 (N_22068,N_21262,N_20683);
and U22069 (N_22069,N_20898,N_21103);
or U22070 (N_22070,N_21162,N_21578);
nor U22071 (N_22071,N_20632,N_21348);
or U22072 (N_22072,N_20873,N_20665);
nand U22073 (N_22073,N_21588,N_20648);
and U22074 (N_22074,N_20818,N_20438);
nor U22075 (N_22075,N_20944,N_21227);
nand U22076 (N_22076,N_21480,N_21590);
and U22077 (N_22077,N_21090,N_20479);
or U22078 (N_22078,N_20965,N_21102);
nand U22079 (N_22079,N_20676,N_21197);
and U22080 (N_22080,N_21019,N_20418);
nor U22081 (N_22081,N_21263,N_21502);
nand U22082 (N_22082,N_21541,N_21060);
nor U22083 (N_22083,N_21017,N_20431);
xor U22084 (N_22084,N_20535,N_20850);
xnor U22085 (N_22085,N_20689,N_20542);
xnor U22086 (N_22086,N_21579,N_21425);
nand U22087 (N_22087,N_20605,N_21216);
xor U22088 (N_22088,N_21087,N_20670);
and U22089 (N_22089,N_20845,N_21357);
xnor U22090 (N_22090,N_21340,N_20578);
xor U22091 (N_22091,N_21398,N_20759);
nor U22092 (N_22092,N_20934,N_20925);
and U22093 (N_22093,N_20563,N_20730);
nor U22094 (N_22094,N_21053,N_20756);
nand U22095 (N_22095,N_20651,N_21555);
nand U22096 (N_22096,N_20740,N_20928);
nor U22097 (N_22097,N_21549,N_20538);
nand U22098 (N_22098,N_20785,N_20894);
and U22099 (N_22099,N_21323,N_21225);
xnor U22100 (N_22100,N_21292,N_20666);
or U22101 (N_22101,N_21431,N_20531);
nor U22102 (N_22102,N_20463,N_21302);
xnor U22103 (N_22103,N_20474,N_21050);
xor U22104 (N_22104,N_20821,N_21209);
nor U22105 (N_22105,N_20584,N_21115);
xnor U22106 (N_22106,N_21009,N_21376);
and U22107 (N_22107,N_20439,N_20768);
nor U22108 (N_22108,N_20920,N_21237);
or U22109 (N_22109,N_20929,N_20566);
or U22110 (N_22110,N_20456,N_20764);
or U22111 (N_22111,N_21276,N_21198);
or U22112 (N_22112,N_21387,N_20621);
nand U22113 (N_22113,N_21519,N_21088);
nand U22114 (N_22114,N_20424,N_21047);
or U22115 (N_22115,N_20705,N_21413);
nor U22116 (N_22116,N_20627,N_20495);
nand U22117 (N_22117,N_21492,N_20854);
nand U22118 (N_22118,N_21444,N_21575);
nand U22119 (N_22119,N_21587,N_20746);
nand U22120 (N_22120,N_20552,N_20437);
or U22121 (N_22121,N_20590,N_21345);
or U22122 (N_22122,N_21412,N_20465);
xor U22123 (N_22123,N_20752,N_20923);
or U22124 (N_22124,N_21522,N_21597);
xnor U22125 (N_22125,N_21117,N_20865);
nand U22126 (N_22126,N_20490,N_21132);
nor U22127 (N_22127,N_20940,N_21503);
nor U22128 (N_22128,N_21373,N_21455);
and U22129 (N_22129,N_20972,N_20904);
and U22130 (N_22130,N_20560,N_21460);
xnor U22131 (N_22131,N_21125,N_20813);
nor U22132 (N_22132,N_21187,N_20701);
nor U22133 (N_22133,N_21453,N_20960);
and U22134 (N_22134,N_21514,N_21419);
nand U22135 (N_22135,N_20481,N_20485);
and U22136 (N_22136,N_21094,N_20446);
or U22137 (N_22137,N_20811,N_21026);
nor U22138 (N_22138,N_20459,N_20555);
or U22139 (N_22139,N_20708,N_20487);
or U22140 (N_22140,N_20997,N_21277);
nor U22141 (N_22141,N_21512,N_20922);
or U22142 (N_22142,N_21450,N_21205);
nand U22143 (N_22143,N_20815,N_20533);
and U22144 (N_22144,N_21097,N_21220);
nor U22145 (N_22145,N_20749,N_20794);
and U22146 (N_22146,N_20963,N_21596);
nand U22147 (N_22147,N_21476,N_21410);
and U22148 (N_22148,N_20460,N_21542);
nand U22149 (N_22149,N_21375,N_20881);
or U22150 (N_22150,N_21334,N_21473);
and U22151 (N_22151,N_21327,N_20516);
or U22152 (N_22152,N_21041,N_21403);
nor U22153 (N_22153,N_21155,N_20599);
nand U22154 (N_22154,N_21459,N_20958);
or U22155 (N_22155,N_21570,N_21300);
nor U22156 (N_22156,N_21517,N_21173);
or U22157 (N_22157,N_20789,N_21029);
nand U22158 (N_22158,N_21243,N_21562);
xor U22159 (N_22159,N_20461,N_21079);
or U22160 (N_22160,N_20948,N_21030);
nand U22161 (N_22161,N_21379,N_20686);
and U22162 (N_22162,N_21044,N_21037);
nor U22163 (N_22163,N_20455,N_21153);
and U22164 (N_22164,N_21500,N_20874);
nor U22165 (N_22165,N_20973,N_21595);
nand U22166 (N_22166,N_20453,N_21489);
xnor U22167 (N_22167,N_20711,N_21203);
or U22168 (N_22168,N_20502,N_21252);
or U22169 (N_22169,N_21099,N_20717);
nor U22170 (N_22170,N_20496,N_21525);
and U22171 (N_22171,N_20814,N_20998);
nor U22172 (N_22172,N_21526,N_21551);
or U22173 (N_22173,N_21408,N_21428);
nor U22174 (N_22174,N_20988,N_20435);
and U22175 (N_22175,N_21390,N_21545);
xnor U22176 (N_22176,N_20556,N_21066);
or U22177 (N_22177,N_20855,N_21062);
nor U22178 (N_22178,N_21322,N_20410);
and U22179 (N_22179,N_21093,N_20647);
and U22180 (N_22180,N_20712,N_20912);
or U22181 (N_22181,N_21014,N_21131);
nand U22182 (N_22182,N_20572,N_21372);
xnor U22183 (N_22183,N_20779,N_21266);
or U22184 (N_22184,N_21599,N_20506);
or U22185 (N_22185,N_20724,N_21065);
or U22186 (N_22186,N_21592,N_20558);
and U22187 (N_22187,N_20720,N_21003);
and U22188 (N_22188,N_20478,N_20933);
xnor U22189 (N_22189,N_21241,N_21516);
nor U22190 (N_22190,N_20796,N_21193);
or U22191 (N_22191,N_21142,N_20511);
and U22192 (N_22192,N_20630,N_21213);
xor U22193 (N_22193,N_20603,N_20935);
nand U22194 (N_22194,N_20432,N_20841);
and U22195 (N_22195,N_20995,N_20422);
nand U22196 (N_22196,N_21362,N_20876);
and U22197 (N_22197,N_21427,N_21374);
nor U22198 (N_22198,N_21366,N_20428);
or U22199 (N_22199,N_20981,N_21204);
nand U22200 (N_22200,N_21579,N_21026);
nor U22201 (N_22201,N_21447,N_21009);
nand U22202 (N_22202,N_21039,N_21431);
xnor U22203 (N_22203,N_20897,N_21051);
nand U22204 (N_22204,N_20973,N_21305);
and U22205 (N_22205,N_21432,N_21539);
xnor U22206 (N_22206,N_21571,N_20425);
nor U22207 (N_22207,N_20546,N_21035);
nand U22208 (N_22208,N_20727,N_20693);
nor U22209 (N_22209,N_20852,N_20533);
nor U22210 (N_22210,N_21327,N_21134);
and U22211 (N_22211,N_21033,N_20688);
nand U22212 (N_22212,N_21457,N_21522);
nand U22213 (N_22213,N_21170,N_20976);
xor U22214 (N_22214,N_21284,N_20440);
xor U22215 (N_22215,N_20551,N_20851);
and U22216 (N_22216,N_20674,N_21025);
nor U22217 (N_22217,N_20685,N_21085);
or U22218 (N_22218,N_21002,N_20620);
and U22219 (N_22219,N_20497,N_21453);
nor U22220 (N_22220,N_20685,N_21543);
xor U22221 (N_22221,N_21169,N_21276);
nand U22222 (N_22222,N_21136,N_20419);
and U22223 (N_22223,N_20690,N_21297);
nand U22224 (N_22224,N_21291,N_20455);
xnor U22225 (N_22225,N_21316,N_20751);
xnor U22226 (N_22226,N_20776,N_21076);
nor U22227 (N_22227,N_21020,N_20401);
or U22228 (N_22228,N_21517,N_21082);
xnor U22229 (N_22229,N_21467,N_21127);
nand U22230 (N_22230,N_20770,N_21509);
and U22231 (N_22231,N_21070,N_21522);
nand U22232 (N_22232,N_21026,N_20731);
and U22233 (N_22233,N_20572,N_21314);
xnor U22234 (N_22234,N_21381,N_21144);
nor U22235 (N_22235,N_20649,N_20598);
nor U22236 (N_22236,N_21552,N_21560);
or U22237 (N_22237,N_20802,N_21056);
nor U22238 (N_22238,N_20491,N_20725);
or U22239 (N_22239,N_20770,N_20528);
or U22240 (N_22240,N_20659,N_21319);
and U22241 (N_22241,N_20782,N_21247);
nand U22242 (N_22242,N_21200,N_21512);
nand U22243 (N_22243,N_20907,N_21439);
xnor U22244 (N_22244,N_20696,N_20685);
or U22245 (N_22245,N_20435,N_20541);
nand U22246 (N_22246,N_21411,N_21127);
nand U22247 (N_22247,N_21328,N_21554);
or U22248 (N_22248,N_20400,N_20431);
or U22249 (N_22249,N_20594,N_20649);
xnor U22250 (N_22250,N_21517,N_20669);
nor U22251 (N_22251,N_21444,N_20665);
xor U22252 (N_22252,N_21019,N_21551);
and U22253 (N_22253,N_20473,N_20840);
and U22254 (N_22254,N_20411,N_20633);
nand U22255 (N_22255,N_21198,N_20779);
nand U22256 (N_22256,N_21114,N_21139);
xor U22257 (N_22257,N_21288,N_20882);
and U22258 (N_22258,N_21304,N_20620);
xnor U22259 (N_22259,N_21042,N_21285);
xnor U22260 (N_22260,N_21429,N_20590);
nand U22261 (N_22261,N_20432,N_20661);
nor U22262 (N_22262,N_20471,N_21352);
nor U22263 (N_22263,N_21419,N_21428);
or U22264 (N_22264,N_20819,N_20957);
and U22265 (N_22265,N_20535,N_21377);
xor U22266 (N_22266,N_21079,N_21182);
nor U22267 (N_22267,N_21007,N_21483);
xor U22268 (N_22268,N_21139,N_21551);
xor U22269 (N_22269,N_20786,N_21473);
or U22270 (N_22270,N_20832,N_20607);
xnor U22271 (N_22271,N_21318,N_21104);
or U22272 (N_22272,N_21530,N_20699);
or U22273 (N_22273,N_21574,N_20545);
and U22274 (N_22274,N_20493,N_21552);
and U22275 (N_22275,N_20518,N_20460);
and U22276 (N_22276,N_20663,N_20434);
or U22277 (N_22277,N_20792,N_20742);
or U22278 (N_22278,N_21086,N_21462);
and U22279 (N_22279,N_21433,N_20455);
nor U22280 (N_22280,N_21149,N_20857);
or U22281 (N_22281,N_21163,N_20625);
nor U22282 (N_22282,N_20658,N_21005);
or U22283 (N_22283,N_20566,N_20956);
nor U22284 (N_22284,N_21526,N_21099);
nand U22285 (N_22285,N_20510,N_20497);
xor U22286 (N_22286,N_21572,N_20573);
nor U22287 (N_22287,N_20941,N_20428);
or U22288 (N_22288,N_20937,N_20943);
xnor U22289 (N_22289,N_21456,N_21472);
or U22290 (N_22290,N_21468,N_20588);
xor U22291 (N_22291,N_20425,N_21230);
nand U22292 (N_22292,N_20717,N_21170);
and U22293 (N_22293,N_21333,N_20707);
xnor U22294 (N_22294,N_20479,N_21255);
nand U22295 (N_22295,N_20921,N_21459);
or U22296 (N_22296,N_20692,N_21033);
or U22297 (N_22297,N_20981,N_21058);
and U22298 (N_22298,N_20946,N_21131);
xnor U22299 (N_22299,N_20439,N_20717);
nand U22300 (N_22300,N_21329,N_21575);
and U22301 (N_22301,N_20781,N_21197);
nor U22302 (N_22302,N_21202,N_20656);
nor U22303 (N_22303,N_21418,N_20430);
nor U22304 (N_22304,N_20635,N_21387);
nand U22305 (N_22305,N_21180,N_20583);
or U22306 (N_22306,N_20753,N_21246);
xnor U22307 (N_22307,N_21406,N_20789);
nor U22308 (N_22308,N_21035,N_21013);
xnor U22309 (N_22309,N_21251,N_20957);
nand U22310 (N_22310,N_21335,N_21005);
xnor U22311 (N_22311,N_20898,N_21180);
xor U22312 (N_22312,N_21003,N_21149);
or U22313 (N_22313,N_20793,N_21328);
xnor U22314 (N_22314,N_20979,N_20606);
or U22315 (N_22315,N_20921,N_21436);
and U22316 (N_22316,N_21171,N_20974);
nor U22317 (N_22317,N_20677,N_21421);
nor U22318 (N_22318,N_20763,N_20549);
nor U22319 (N_22319,N_21087,N_21506);
or U22320 (N_22320,N_20557,N_21478);
nand U22321 (N_22321,N_21462,N_20601);
nand U22322 (N_22322,N_21340,N_20855);
and U22323 (N_22323,N_21001,N_21362);
and U22324 (N_22324,N_20883,N_21478);
xnor U22325 (N_22325,N_20757,N_20736);
xor U22326 (N_22326,N_21434,N_21118);
or U22327 (N_22327,N_21290,N_21246);
nor U22328 (N_22328,N_20789,N_21011);
nand U22329 (N_22329,N_21172,N_20999);
xnor U22330 (N_22330,N_20935,N_20441);
xnor U22331 (N_22331,N_20681,N_21540);
nor U22332 (N_22332,N_21598,N_20844);
or U22333 (N_22333,N_20684,N_21054);
nor U22334 (N_22334,N_21233,N_21473);
or U22335 (N_22335,N_20678,N_21573);
nand U22336 (N_22336,N_20513,N_21413);
nor U22337 (N_22337,N_20944,N_20418);
xnor U22338 (N_22338,N_21354,N_21280);
xnor U22339 (N_22339,N_20881,N_21068);
nor U22340 (N_22340,N_20913,N_20652);
nand U22341 (N_22341,N_21362,N_20955);
nand U22342 (N_22342,N_20681,N_20651);
or U22343 (N_22343,N_20917,N_21248);
or U22344 (N_22344,N_20733,N_20846);
or U22345 (N_22345,N_20897,N_20646);
or U22346 (N_22346,N_21395,N_20508);
xor U22347 (N_22347,N_21375,N_20529);
or U22348 (N_22348,N_21589,N_21121);
nand U22349 (N_22349,N_21326,N_21050);
nor U22350 (N_22350,N_20514,N_21479);
or U22351 (N_22351,N_20743,N_21263);
xnor U22352 (N_22352,N_20519,N_20406);
or U22353 (N_22353,N_20400,N_20837);
nand U22354 (N_22354,N_20694,N_21080);
nor U22355 (N_22355,N_20617,N_20960);
xor U22356 (N_22356,N_21110,N_21073);
nand U22357 (N_22357,N_20694,N_20617);
nor U22358 (N_22358,N_20900,N_21538);
nand U22359 (N_22359,N_20933,N_20920);
nand U22360 (N_22360,N_21220,N_20860);
nand U22361 (N_22361,N_20754,N_21293);
or U22362 (N_22362,N_20462,N_21117);
and U22363 (N_22363,N_20400,N_21199);
and U22364 (N_22364,N_20761,N_20989);
nor U22365 (N_22365,N_20941,N_21109);
or U22366 (N_22366,N_21417,N_20793);
or U22367 (N_22367,N_20627,N_20837);
xnor U22368 (N_22368,N_21038,N_21082);
nand U22369 (N_22369,N_21411,N_21425);
nor U22370 (N_22370,N_20752,N_20472);
or U22371 (N_22371,N_20853,N_21054);
nand U22372 (N_22372,N_20920,N_20877);
nor U22373 (N_22373,N_21533,N_21376);
nand U22374 (N_22374,N_20766,N_20509);
nand U22375 (N_22375,N_21398,N_20968);
xor U22376 (N_22376,N_21465,N_20913);
xnor U22377 (N_22377,N_21461,N_20698);
or U22378 (N_22378,N_20846,N_20577);
nand U22379 (N_22379,N_21387,N_20508);
xnor U22380 (N_22380,N_20412,N_21587);
and U22381 (N_22381,N_21079,N_21024);
nand U22382 (N_22382,N_21027,N_21515);
nand U22383 (N_22383,N_20679,N_20482);
nor U22384 (N_22384,N_21324,N_20526);
and U22385 (N_22385,N_20690,N_21104);
xnor U22386 (N_22386,N_21227,N_21130);
or U22387 (N_22387,N_20920,N_21510);
and U22388 (N_22388,N_20414,N_21097);
nor U22389 (N_22389,N_20872,N_20821);
nand U22390 (N_22390,N_21389,N_21414);
xnor U22391 (N_22391,N_21039,N_20797);
nor U22392 (N_22392,N_20889,N_20893);
nor U22393 (N_22393,N_20551,N_21124);
xnor U22394 (N_22394,N_20965,N_21579);
and U22395 (N_22395,N_20994,N_20692);
nand U22396 (N_22396,N_20939,N_20618);
or U22397 (N_22397,N_20662,N_20877);
xor U22398 (N_22398,N_20672,N_21383);
xor U22399 (N_22399,N_20670,N_20422);
xnor U22400 (N_22400,N_20413,N_21332);
nor U22401 (N_22401,N_20825,N_21483);
xor U22402 (N_22402,N_21437,N_20536);
or U22403 (N_22403,N_21494,N_20710);
xnor U22404 (N_22404,N_21197,N_20744);
nor U22405 (N_22405,N_21134,N_21168);
xor U22406 (N_22406,N_20914,N_21424);
nand U22407 (N_22407,N_20525,N_21406);
nand U22408 (N_22408,N_21026,N_21553);
or U22409 (N_22409,N_20791,N_20476);
or U22410 (N_22410,N_21083,N_20977);
and U22411 (N_22411,N_21016,N_21433);
nand U22412 (N_22412,N_20676,N_20894);
nor U22413 (N_22413,N_21534,N_20841);
nand U22414 (N_22414,N_20588,N_21178);
nor U22415 (N_22415,N_21334,N_20556);
nor U22416 (N_22416,N_20509,N_21114);
nand U22417 (N_22417,N_21351,N_20908);
nand U22418 (N_22418,N_21122,N_21199);
xnor U22419 (N_22419,N_20444,N_20442);
and U22420 (N_22420,N_20868,N_21113);
nor U22421 (N_22421,N_20766,N_20755);
nand U22422 (N_22422,N_20841,N_21387);
nand U22423 (N_22423,N_20624,N_20911);
nand U22424 (N_22424,N_21142,N_21366);
and U22425 (N_22425,N_21087,N_20663);
xor U22426 (N_22426,N_20561,N_20919);
or U22427 (N_22427,N_20915,N_21490);
and U22428 (N_22428,N_20844,N_21137);
nor U22429 (N_22429,N_21542,N_21018);
xor U22430 (N_22430,N_20862,N_20868);
xor U22431 (N_22431,N_20809,N_20863);
and U22432 (N_22432,N_21014,N_20827);
nand U22433 (N_22433,N_20529,N_21533);
nand U22434 (N_22434,N_21050,N_20672);
or U22435 (N_22435,N_20925,N_20600);
xor U22436 (N_22436,N_20883,N_20435);
nand U22437 (N_22437,N_21179,N_20892);
xor U22438 (N_22438,N_20760,N_21266);
nand U22439 (N_22439,N_20760,N_20410);
and U22440 (N_22440,N_21193,N_20554);
and U22441 (N_22441,N_20577,N_21353);
and U22442 (N_22442,N_20459,N_21488);
or U22443 (N_22443,N_20407,N_20670);
and U22444 (N_22444,N_21061,N_20949);
nor U22445 (N_22445,N_20761,N_21112);
nor U22446 (N_22446,N_21159,N_21065);
or U22447 (N_22447,N_20595,N_21188);
nand U22448 (N_22448,N_21079,N_20974);
or U22449 (N_22449,N_21504,N_21392);
nand U22450 (N_22450,N_20523,N_20416);
xor U22451 (N_22451,N_20645,N_21595);
nand U22452 (N_22452,N_20431,N_20895);
xor U22453 (N_22453,N_21572,N_20606);
xnor U22454 (N_22454,N_20942,N_20528);
and U22455 (N_22455,N_21470,N_20795);
nand U22456 (N_22456,N_20684,N_20649);
nand U22457 (N_22457,N_21277,N_21423);
nor U22458 (N_22458,N_21300,N_21535);
nand U22459 (N_22459,N_21395,N_20985);
xor U22460 (N_22460,N_20607,N_21511);
or U22461 (N_22461,N_20957,N_21250);
or U22462 (N_22462,N_21409,N_20630);
and U22463 (N_22463,N_21386,N_20672);
and U22464 (N_22464,N_20661,N_20690);
or U22465 (N_22465,N_21543,N_21083);
and U22466 (N_22466,N_21188,N_20718);
and U22467 (N_22467,N_20817,N_20597);
nand U22468 (N_22468,N_20787,N_21336);
and U22469 (N_22469,N_21353,N_21480);
or U22470 (N_22470,N_21089,N_20971);
and U22471 (N_22471,N_21021,N_21118);
or U22472 (N_22472,N_21490,N_21472);
nor U22473 (N_22473,N_21507,N_21485);
xnor U22474 (N_22474,N_21036,N_20973);
or U22475 (N_22475,N_20647,N_20697);
or U22476 (N_22476,N_20987,N_20524);
or U22477 (N_22477,N_21158,N_21572);
or U22478 (N_22478,N_21360,N_21280);
and U22479 (N_22479,N_21276,N_20482);
nor U22480 (N_22480,N_21213,N_20647);
xor U22481 (N_22481,N_21411,N_21073);
xnor U22482 (N_22482,N_20874,N_20798);
xor U22483 (N_22483,N_21042,N_21391);
and U22484 (N_22484,N_21002,N_21068);
xnor U22485 (N_22485,N_20673,N_21040);
nor U22486 (N_22486,N_21051,N_21594);
xnor U22487 (N_22487,N_21191,N_21017);
or U22488 (N_22488,N_20733,N_21175);
xnor U22489 (N_22489,N_20935,N_20806);
or U22490 (N_22490,N_20877,N_21399);
or U22491 (N_22491,N_21161,N_21101);
xor U22492 (N_22492,N_20535,N_20885);
xnor U22493 (N_22493,N_21036,N_20440);
or U22494 (N_22494,N_20548,N_21350);
nand U22495 (N_22495,N_20948,N_21269);
xor U22496 (N_22496,N_21220,N_20901);
and U22497 (N_22497,N_20503,N_20668);
and U22498 (N_22498,N_20659,N_20737);
or U22499 (N_22499,N_21406,N_20541);
or U22500 (N_22500,N_20535,N_20970);
nand U22501 (N_22501,N_20598,N_21350);
or U22502 (N_22502,N_21448,N_21210);
nor U22503 (N_22503,N_20492,N_21482);
or U22504 (N_22504,N_21112,N_20538);
nor U22505 (N_22505,N_21456,N_20547);
xnor U22506 (N_22506,N_21060,N_20976);
nand U22507 (N_22507,N_20953,N_20562);
nand U22508 (N_22508,N_21583,N_20922);
nor U22509 (N_22509,N_21209,N_20515);
nand U22510 (N_22510,N_21494,N_20484);
xor U22511 (N_22511,N_20729,N_20530);
nor U22512 (N_22512,N_20988,N_21249);
or U22513 (N_22513,N_20754,N_20845);
or U22514 (N_22514,N_21471,N_20734);
and U22515 (N_22515,N_20795,N_20786);
nand U22516 (N_22516,N_21417,N_20662);
nor U22517 (N_22517,N_20997,N_20746);
nor U22518 (N_22518,N_20927,N_21234);
nand U22519 (N_22519,N_21503,N_20637);
or U22520 (N_22520,N_21019,N_21108);
or U22521 (N_22521,N_20591,N_20645);
nor U22522 (N_22522,N_21566,N_21216);
and U22523 (N_22523,N_21467,N_21334);
or U22524 (N_22524,N_20956,N_20879);
or U22525 (N_22525,N_21488,N_20915);
nor U22526 (N_22526,N_21264,N_21009);
or U22527 (N_22527,N_20611,N_20886);
nand U22528 (N_22528,N_21243,N_21402);
or U22529 (N_22529,N_20918,N_21384);
xor U22530 (N_22530,N_20836,N_20854);
nor U22531 (N_22531,N_21597,N_21269);
nor U22532 (N_22532,N_21432,N_21168);
nor U22533 (N_22533,N_20612,N_21534);
nor U22534 (N_22534,N_20513,N_21304);
xor U22535 (N_22535,N_20494,N_20989);
nand U22536 (N_22536,N_20551,N_20645);
nor U22537 (N_22537,N_20997,N_20917);
xnor U22538 (N_22538,N_21555,N_21512);
xnor U22539 (N_22539,N_21088,N_20625);
and U22540 (N_22540,N_21241,N_20736);
and U22541 (N_22541,N_20648,N_20467);
nand U22542 (N_22542,N_20569,N_20691);
xor U22543 (N_22543,N_20705,N_20730);
or U22544 (N_22544,N_21408,N_21076);
and U22545 (N_22545,N_21051,N_20528);
xor U22546 (N_22546,N_20902,N_20777);
nor U22547 (N_22547,N_21420,N_20593);
nor U22548 (N_22548,N_21538,N_21160);
xor U22549 (N_22549,N_20588,N_21296);
or U22550 (N_22550,N_21017,N_21238);
nand U22551 (N_22551,N_21300,N_20641);
nor U22552 (N_22552,N_20468,N_21241);
nor U22553 (N_22553,N_21599,N_20424);
xnor U22554 (N_22554,N_21379,N_20952);
or U22555 (N_22555,N_20486,N_20633);
or U22556 (N_22556,N_20943,N_20779);
nor U22557 (N_22557,N_21234,N_20800);
xor U22558 (N_22558,N_21320,N_20956);
or U22559 (N_22559,N_20658,N_20929);
or U22560 (N_22560,N_21060,N_20790);
nor U22561 (N_22561,N_21252,N_21416);
nor U22562 (N_22562,N_21366,N_21260);
nor U22563 (N_22563,N_20646,N_20899);
or U22564 (N_22564,N_20500,N_20955);
and U22565 (N_22565,N_21253,N_21294);
and U22566 (N_22566,N_20621,N_20646);
and U22567 (N_22567,N_20544,N_20973);
or U22568 (N_22568,N_21562,N_20565);
xnor U22569 (N_22569,N_20755,N_21559);
nand U22570 (N_22570,N_20669,N_21187);
xor U22571 (N_22571,N_21351,N_20560);
and U22572 (N_22572,N_21569,N_21223);
nand U22573 (N_22573,N_20903,N_20858);
nand U22574 (N_22574,N_20695,N_20785);
nor U22575 (N_22575,N_20554,N_21381);
and U22576 (N_22576,N_21408,N_20932);
nor U22577 (N_22577,N_20707,N_20949);
nor U22578 (N_22578,N_21030,N_20755);
nand U22579 (N_22579,N_21551,N_20998);
and U22580 (N_22580,N_20782,N_21103);
nand U22581 (N_22581,N_21546,N_20472);
or U22582 (N_22582,N_21427,N_20946);
nor U22583 (N_22583,N_21189,N_20620);
nand U22584 (N_22584,N_21213,N_20540);
and U22585 (N_22585,N_21001,N_20783);
and U22586 (N_22586,N_21416,N_21023);
and U22587 (N_22587,N_20919,N_21144);
xnor U22588 (N_22588,N_21147,N_21350);
or U22589 (N_22589,N_21126,N_21099);
and U22590 (N_22590,N_20847,N_20968);
or U22591 (N_22591,N_21495,N_21005);
and U22592 (N_22592,N_21513,N_21518);
or U22593 (N_22593,N_20725,N_20659);
or U22594 (N_22594,N_21438,N_21545);
or U22595 (N_22595,N_21191,N_20513);
nor U22596 (N_22596,N_21267,N_20972);
and U22597 (N_22597,N_21451,N_20700);
or U22598 (N_22598,N_20440,N_20425);
nand U22599 (N_22599,N_21484,N_21170);
nand U22600 (N_22600,N_20946,N_21471);
xnor U22601 (N_22601,N_20404,N_20748);
nand U22602 (N_22602,N_20640,N_20616);
nor U22603 (N_22603,N_21520,N_20664);
or U22604 (N_22604,N_21355,N_20446);
nand U22605 (N_22605,N_20842,N_20823);
nor U22606 (N_22606,N_20411,N_20871);
and U22607 (N_22607,N_21115,N_20793);
or U22608 (N_22608,N_21545,N_20464);
and U22609 (N_22609,N_20812,N_21557);
xnor U22610 (N_22610,N_21050,N_20464);
xor U22611 (N_22611,N_21176,N_20842);
nand U22612 (N_22612,N_20492,N_21365);
nand U22613 (N_22613,N_20768,N_21020);
or U22614 (N_22614,N_21134,N_20605);
nor U22615 (N_22615,N_21085,N_21435);
nor U22616 (N_22616,N_21077,N_20689);
and U22617 (N_22617,N_21030,N_21246);
xor U22618 (N_22618,N_21299,N_21518);
or U22619 (N_22619,N_20517,N_20852);
xor U22620 (N_22620,N_20489,N_20837);
nand U22621 (N_22621,N_20472,N_20859);
nor U22622 (N_22622,N_21394,N_21596);
or U22623 (N_22623,N_21246,N_20756);
or U22624 (N_22624,N_21026,N_20691);
nand U22625 (N_22625,N_21191,N_21565);
nor U22626 (N_22626,N_20441,N_21567);
and U22627 (N_22627,N_20594,N_20897);
xnor U22628 (N_22628,N_21260,N_21511);
nor U22629 (N_22629,N_21039,N_20867);
nand U22630 (N_22630,N_20744,N_20875);
or U22631 (N_22631,N_20762,N_21010);
nand U22632 (N_22632,N_21361,N_21354);
nor U22633 (N_22633,N_20700,N_21241);
xnor U22634 (N_22634,N_20674,N_20470);
or U22635 (N_22635,N_21584,N_20491);
nor U22636 (N_22636,N_20810,N_21459);
nor U22637 (N_22637,N_21161,N_20454);
and U22638 (N_22638,N_20664,N_20526);
and U22639 (N_22639,N_21203,N_21388);
nand U22640 (N_22640,N_20787,N_21549);
and U22641 (N_22641,N_20997,N_20914);
or U22642 (N_22642,N_21450,N_20890);
nor U22643 (N_22643,N_21341,N_21253);
xor U22644 (N_22644,N_20896,N_21418);
xor U22645 (N_22645,N_21472,N_20663);
or U22646 (N_22646,N_21076,N_21020);
or U22647 (N_22647,N_21145,N_20638);
xnor U22648 (N_22648,N_20415,N_20705);
nor U22649 (N_22649,N_20688,N_21458);
or U22650 (N_22650,N_21016,N_20920);
or U22651 (N_22651,N_20876,N_21325);
nor U22652 (N_22652,N_20573,N_21096);
nor U22653 (N_22653,N_21315,N_20909);
xnor U22654 (N_22654,N_20569,N_20547);
nor U22655 (N_22655,N_21136,N_20551);
nor U22656 (N_22656,N_21438,N_21239);
nand U22657 (N_22657,N_21494,N_20899);
xor U22658 (N_22658,N_21119,N_20818);
or U22659 (N_22659,N_20797,N_20588);
and U22660 (N_22660,N_21292,N_21402);
xor U22661 (N_22661,N_20805,N_20881);
nor U22662 (N_22662,N_20818,N_20776);
nand U22663 (N_22663,N_20485,N_21095);
xnor U22664 (N_22664,N_21432,N_21511);
nand U22665 (N_22665,N_20641,N_20962);
nor U22666 (N_22666,N_21242,N_21178);
or U22667 (N_22667,N_20743,N_21066);
nor U22668 (N_22668,N_21493,N_20799);
or U22669 (N_22669,N_20857,N_20978);
or U22670 (N_22670,N_21072,N_21042);
and U22671 (N_22671,N_21224,N_20558);
or U22672 (N_22672,N_21431,N_20970);
and U22673 (N_22673,N_21224,N_20976);
and U22674 (N_22674,N_20936,N_20816);
nor U22675 (N_22675,N_20545,N_21586);
and U22676 (N_22676,N_21122,N_21159);
nor U22677 (N_22677,N_21058,N_21286);
and U22678 (N_22678,N_20922,N_20888);
or U22679 (N_22679,N_21233,N_21109);
xor U22680 (N_22680,N_20503,N_20621);
nor U22681 (N_22681,N_21026,N_21567);
and U22682 (N_22682,N_20696,N_21422);
nor U22683 (N_22683,N_21051,N_21020);
xnor U22684 (N_22684,N_20453,N_21272);
and U22685 (N_22685,N_21148,N_21493);
nand U22686 (N_22686,N_21378,N_20629);
or U22687 (N_22687,N_20825,N_21511);
nand U22688 (N_22688,N_20725,N_21200);
and U22689 (N_22689,N_20657,N_20754);
xnor U22690 (N_22690,N_21318,N_21510);
nand U22691 (N_22691,N_21054,N_21389);
nor U22692 (N_22692,N_21416,N_20985);
xnor U22693 (N_22693,N_21469,N_20729);
nor U22694 (N_22694,N_20521,N_21302);
or U22695 (N_22695,N_21230,N_20848);
xor U22696 (N_22696,N_21564,N_20781);
nor U22697 (N_22697,N_21058,N_20471);
or U22698 (N_22698,N_20606,N_20834);
nor U22699 (N_22699,N_20588,N_21090);
or U22700 (N_22700,N_21021,N_21130);
nor U22701 (N_22701,N_21054,N_20915);
nand U22702 (N_22702,N_20751,N_20489);
nor U22703 (N_22703,N_21074,N_21194);
or U22704 (N_22704,N_21086,N_20794);
nand U22705 (N_22705,N_21127,N_21575);
nor U22706 (N_22706,N_20925,N_21519);
nand U22707 (N_22707,N_21397,N_21440);
xnor U22708 (N_22708,N_21498,N_21597);
xnor U22709 (N_22709,N_21132,N_20896);
xor U22710 (N_22710,N_20920,N_20873);
nor U22711 (N_22711,N_20987,N_21469);
and U22712 (N_22712,N_20692,N_20588);
nor U22713 (N_22713,N_20414,N_21491);
xor U22714 (N_22714,N_20664,N_21125);
or U22715 (N_22715,N_20408,N_20712);
or U22716 (N_22716,N_21070,N_21353);
or U22717 (N_22717,N_20970,N_20973);
and U22718 (N_22718,N_21025,N_21117);
xnor U22719 (N_22719,N_21110,N_20542);
nand U22720 (N_22720,N_21448,N_21200);
nand U22721 (N_22721,N_21070,N_20652);
nor U22722 (N_22722,N_20602,N_21079);
or U22723 (N_22723,N_20484,N_20602);
nand U22724 (N_22724,N_20754,N_20848);
or U22725 (N_22725,N_21258,N_20563);
or U22726 (N_22726,N_21551,N_21051);
and U22727 (N_22727,N_20475,N_20546);
or U22728 (N_22728,N_20487,N_21470);
nor U22729 (N_22729,N_20467,N_21338);
xor U22730 (N_22730,N_21426,N_20546);
nand U22731 (N_22731,N_21572,N_21272);
nor U22732 (N_22732,N_21429,N_20414);
xor U22733 (N_22733,N_21164,N_20927);
xor U22734 (N_22734,N_20941,N_21271);
and U22735 (N_22735,N_20954,N_20875);
nor U22736 (N_22736,N_20947,N_20879);
and U22737 (N_22737,N_20978,N_20719);
xor U22738 (N_22738,N_20634,N_20804);
nor U22739 (N_22739,N_20801,N_20793);
nand U22740 (N_22740,N_21281,N_21543);
or U22741 (N_22741,N_21489,N_21236);
and U22742 (N_22742,N_21263,N_21011);
nand U22743 (N_22743,N_20935,N_21127);
xor U22744 (N_22744,N_20689,N_20634);
nand U22745 (N_22745,N_20597,N_20435);
nor U22746 (N_22746,N_20592,N_21334);
or U22747 (N_22747,N_20628,N_21106);
xnor U22748 (N_22748,N_20437,N_21315);
nor U22749 (N_22749,N_20640,N_21475);
or U22750 (N_22750,N_21540,N_20904);
xnor U22751 (N_22751,N_20641,N_21095);
xor U22752 (N_22752,N_20810,N_20537);
nand U22753 (N_22753,N_21302,N_20831);
xor U22754 (N_22754,N_21265,N_21351);
nor U22755 (N_22755,N_21452,N_21137);
and U22756 (N_22756,N_20597,N_21317);
or U22757 (N_22757,N_21149,N_21166);
and U22758 (N_22758,N_20658,N_21482);
nor U22759 (N_22759,N_20734,N_20923);
nand U22760 (N_22760,N_20424,N_21265);
xor U22761 (N_22761,N_20400,N_20907);
xor U22762 (N_22762,N_21135,N_20767);
and U22763 (N_22763,N_20788,N_21381);
nor U22764 (N_22764,N_21271,N_21420);
nor U22765 (N_22765,N_21308,N_20592);
nand U22766 (N_22766,N_20500,N_21518);
or U22767 (N_22767,N_20998,N_21149);
nor U22768 (N_22768,N_21466,N_21113);
or U22769 (N_22769,N_21175,N_21578);
xor U22770 (N_22770,N_21420,N_21171);
and U22771 (N_22771,N_20641,N_21323);
xor U22772 (N_22772,N_20624,N_21378);
xor U22773 (N_22773,N_20970,N_21334);
nor U22774 (N_22774,N_20672,N_21286);
nor U22775 (N_22775,N_21042,N_20419);
nor U22776 (N_22776,N_21332,N_20596);
nor U22777 (N_22777,N_20925,N_20620);
or U22778 (N_22778,N_21180,N_21375);
nor U22779 (N_22779,N_21020,N_21044);
or U22780 (N_22780,N_21146,N_20470);
nand U22781 (N_22781,N_21490,N_21367);
xnor U22782 (N_22782,N_21268,N_20905);
nand U22783 (N_22783,N_20893,N_21095);
or U22784 (N_22784,N_21533,N_20928);
nand U22785 (N_22785,N_21037,N_20849);
xnor U22786 (N_22786,N_20874,N_21377);
and U22787 (N_22787,N_20980,N_20788);
nor U22788 (N_22788,N_20585,N_21551);
xor U22789 (N_22789,N_20802,N_21161);
xor U22790 (N_22790,N_20936,N_21596);
and U22791 (N_22791,N_21467,N_20797);
xnor U22792 (N_22792,N_20835,N_20537);
or U22793 (N_22793,N_21480,N_20690);
and U22794 (N_22794,N_20579,N_20714);
xor U22795 (N_22795,N_20441,N_20429);
and U22796 (N_22796,N_20911,N_20422);
or U22797 (N_22797,N_21056,N_21017);
xnor U22798 (N_22798,N_21427,N_20958);
or U22799 (N_22799,N_21413,N_21213);
or U22800 (N_22800,N_22505,N_22317);
or U22801 (N_22801,N_22154,N_22216);
and U22802 (N_22802,N_21830,N_22601);
and U22803 (N_22803,N_22581,N_21909);
and U22804 (N_22804,N_22611,N_21681);
nor U22805 (N_22805,N_22402,N_22178);
and U22806 (N_22806,N_22684,N_22331);
xor U22807 (N_22807,N_22602,N_22352);
and U22808 (N_22808,N_22788,N_22112);
and U22809 (N_22809,N_22038,N_22255);
or U22810 (N_22810,N_21730,N_22768);
and U22811 (N_22811,N_22660,N_22456);
nor U22812 (N_22812,N_21892,N_22508);
xor U22813 (N_22813,N_22403,N_21929);
and U22814 (N_22814,N_22321,N_21619);
nor U22815 (N_22815,N_22375,N_21974);
nor U22816 (N_22816,N_21947,N_21691);
nand U22817 (N_22817,N_21941,N_21756);
and U22818 (N_22818,N_22503,N_22097);
and U22819 (N_22819,N_22516,N_22401);
nand U22820 (N_22820,N_22442,N_22621);
or U22821 (N_22821,N_21978,N_22268);
nand U22822 (N_22822,N_21684,N_22741);
nand U22823 (N_22823,N_22540,N_21663);
nand U22824 (N_22824,N_22361,N_22098);
and U22825 (N_22825,N_22042,N_22333);
nand U22826 (N_22826,N_22658,N_22431);
nor U22827 (N_22827,N_21608,N_22672);
and U22828 (N_22828,N_22374,N_21823);
or U22829 (N_22829,N_22465,N_22522);
or U22830 (N_22830,N_22613,N_22449);
xnor U22831 (N_22831,N_22765,N_21788);
nor U22832 (N_22832,N_21853,N_22344);
or U22833 (N_22833,N_21808,N_21783);
and U22834 (N_22834,N_22359,N_21751);
nand U22835 (N_22835,N_22118,N_22033);
and U22836 (N_22836,N_22063,N_21686);
nand U22837 (N_22837,N_21656,N_22100);
and U22838 (N_22838,N_22451,N_21948);
nand U22839 (N_22839,N_22500,N_21956);
xnor U22840 (N_22840,N_22019,N_22297);
nand U22841 (N_22841,N_21760,N_22328);
and U22842 (N_22842,N_22641,N_22243);
and U22843 (N_22843,N_21845,N_22134);
nor U22844 (N_22844,N_22723,N_22167);
nand U22845 (N_22845,N_22092,N_22701);
or U22846 (N_22846,N_21786,N_22405);
nor U22847 (N_22847,N_21769,N_21846);
nand U22848 (N_22848,N_22358,N_22687);
and U22849 (N_22849,N_21774,N_22586);
xnor U22850 (N_22850,N_21669,N_22190);
xnor U22851 (N_22851,N_21888,N_22133);
xnor U22852 (N_22852,N_21639,N_22346);
and U22853 (N_22853,N_21922,N_21644);
or U22854 (N_22854,N_22282,N_21942);
nand U22855 (N_22855,N_21838,N_21865);
xor U22856 (N_22856,N_22138,N_21984);
xor U22857 (N_22857,N_22023,N_21805);
and U22858 (N_22858,N_22021,N_21637);
nand U22859 (N_22859,N_22523,N_22096);
or U22860 (N_22860,N_22058,N_22709);
nor U22861 (N_22861,N_22084,N_22683);
or U22862 (N_22862,N_21896,N_21802);
nor U22863 (N_22863,N_22559,N_21626);
nand U22864 (N_22864,N_22435,N_21700);
and U22865 (N_22865,N_21825,N_22079);
or U22866 (N_22866,N_22620,N_22335);
and U22867 (N_22867,N_22647,N_22484);
and U22868 (N_22868,N_22164,N_21718);
nand U22869 (N_22869,N_21621,N_22014);
and U22870 (N_22870,N_21685,N_22357);
nor U22871 (N_22871,N_22764,N_21884);
xor U22872 (N_22872,N_22618,N_21795);
and U22873 (N_22873,N_22201,N_22544);
nand U22874 (N_22874,N_22426,N_22674);
nor U22875 (N_22875,N_22369,N_21631);
or U22876 (N_22876,N_21868,N_22666);
or U22877 (N_22877,N_21812,N_21652);
nor U22878 (N_22878,N_21857,N_22372);
and U22879 (N_22879,N_22156,N_22554);
nor U22880 (N_22880,N_21649,N_21706);
xor U22881 (N_22881,N_21765,N_21910);
nor U22882 (N_22882,N_21728,N_21672);
or U22883 (N_22883,N_22205,N_22490);
xor U22884 (N_22884,N_21657,N_22262);
xor U22885 (N_22885,N_21745,N_22560);
or U22886 (N_22886,N_22434,N_21740);
or U22887 (N_22887,N_22228,N_21891);
xnor U22888 (N_22888,N_22087,N_22527);
nand U22889 (N_22889,N_21806,N_21666);
or U22890 (N_22890,N_21906,N_22147);
nor U22891 (N_22891,N_21655,N_21869);
nand U22892 (N_22892,N_21736,N_21878);
and U22893 (N_22893,N_22475,N_22324);
or U22894 (N_22894,N_22071,N_22771);
xnor U22895 (N_22895,N_22729,N_21612);
nor U22896 (N_22896,N_22746,N_22584);
or U22897 (N_22897,N_22137,N_22142);
nor U22898 (N_22898,N_22782,N_21780);
nor U22899 (N_22899,N_21634,N_22759);
nor U22900 (N_22900,N_21982,N_21750);
nor U22901 (N_22901,N_21659,N_22474);
xor U22902 (N_22902,N_21600,N_22325);
or U22903 (N_22903,N_21933,N_22069);
or U22904 (N_22904,N_21983,N_22495);
and U22905 (N_22905,N_21874,N_21969);
and U22906 (N_22906,N_21628,N_22633);
or U22907 (N_22907,N_21955,N_22141);
or U22908 (N_22908,N_22577,N_22727);
or U22909 (N_22909,N_22747,N_22557);
xnor U22910 (N_22910,N_22790,N_21790);
nor U22911 (N_22911,N_22740,N_22541);
xor U22912 (N_22912,N_21796,N_22341);
and U22913 (N_22913,N_22758,N_22389);
nand U22914 (N_22914,N_22444,N_21986);
and U22915 (N_22915,N_22423,N_22140);
nor U22916 (N_22916,N_21994,N_22238);
or U22917 (N_22917,N_22735,N_21839);
nor U22918 (N_22918,N_21815,N_22607);
nor U22919 (N_22919,N_22281,N_22796);
nand U22920 (N_22920,N_21723,N_21690);
nor U22921 (N_22921,N_22531,N_22309);
xnor U22922 (N_22922,N_22638,N_21602);
nand U22923 (N_22923,N_21988,N_22194);
nor U22924 (N_22924,N_21925,N_22717);
nor U22925 (N_22925,N_22253,N_21957);
or U22926 (N_22926,N_22744,N_22212);
nand U22927 (N_22927,N_22223,N_22061);
nand U22928 (N_22928,N_22240,N_22619);
nand U22929 (N_22929,N_22174,N_22578);
or U22930 (N_22930,N_21981,N_21694);
nor U22931 (N_22931,N_21716,N_21887);
and U22932 (N_22932,N_22215,N_21604);
nor U22933 (N_22933,N_22121,N_21636);
nand U22934 (N_22934,N_22158,N_22318);
or U22935 (N_22935,N_22511,N_22575);
xor U22936 (N_22936,N_22264,N_22404);
or U22937 (N_22937,N_22088,N_21813);
nand U22938 (N_22938,N_22161,N_22032);
xnor U22939 (N_22939,N_21938,N_22193);
xor U22940 (N_22940,N_22573,N_22101);
and U22941 (N_22941,N_21759,N_21829);
and U22942 (N_22942,N_22246,N_22629);
xor U22943 (N_22943,N_22691,N_22363);
and U22944 (N_22944,N_22391,N_21799);
nand U22945 (N_22945,N_21658,N_21989);
and U22946 (N_22946,N_21886,N_22200);
or U22947 (N_22947,N_22606,N_21693);
and U22948 (N_22948,N_22186,N_22794);
nand U22949 (N_22949,N_22080,N_21776);
nand U22950 (N_22950,N_22644,N_22707);
xnor U22951 (N_22951,N_22693,N_22183);
and U22952 (N_22952,N_22168,N_22549);
nand U22953 (N_22953,N_22536,N_22424);
nor U22954 (N_22954,N_21601,N_22676);
nor U22955 (N_22955,N_22416,N_22517);
nor U22956 (N_22956,N_21625,N_22292);
and U22957 (N_22957,N_21703,N_22436);
or U22958 (N_22958,N_22179,N_22177);
nand U22959 (N_22959,N_22387,N_21931);
nor U22960 (N_22960,N_22289,N_22284);
or U22961 (N_22961,N_22148,N_22204);
xnor U22962 (N_22962,N_22635,N_22515);
or U22963 (N_22963,N_21960,N_22129);
nand U22964 (N_22964,N_22585,N_22534);
nor U22965 (N_22965,N_22411,N_22276);
nor U22966 (N_22966,N_22236,N_22713);
or U22967 (N_22967,N_22786,N_21661);
nor U22968 (N_22968,N_21856,N_22132);
nand U22969 (N_22969,N_21827,N_22738);
or U22970 (N_22970,N_22187,N_22422);
nor U22971 (N_22971,N_22766,N_22172);
or U22972 (N_22972,N_22330,N_22224);
nor U22973 (N_22973,N_22085,N_22316);
xnor U22974 (N_22974,N_22260,N_22419);
nor U22975 (N_22975,N_22654,N_21711);
nor U22976 (N_22976,N_22463,N_22157);
or U22977 (N_22977,N_22528,N_22526);
nor U22978 (N_22978,N_21821,N_21905);
nor U22979 (N_22979,N_21735,N_22412);
or U22980 (N_22980,N_22628,N_22365);
and U22981 (N_22981,N_22235,N_21819);
and U22982 (N_22982,N_22181,N_22064);
xnor U22983 (N_22983,N_22645,N_22206);
or U22984 (N_22984,N_22234,N_22327);
and U22985 (N_22985,N_21950,N_22694);
or U22986 (N_22986,N_21822,N_22169);
nor U22987 (N_22987,N_22438,N_21784);
or U22988 (N_22988,N_22524,N_21734);
nand U22989 (N_22989,N_22348,N_22288);
or U22990 (N_22990,N_22565,N_21970);
xnor U22991 (N_22991,N_22093,N_22513);
or U22992 (N_22992,N_22624,N_22450);
and U22993 (N_22993,N_21920,N_22469);
nor U22994 (N_22994,N_21847,N_21698);
nand U22995 (N_22995,N_22399,N_21616);
xnor U22996 (N_22996,N_22115,N_22781);
or U22997 (N_22997,N_22409,N_22433);
nand U22998 (N_22998,N_21951,N_22793);
nand U22999 (N_22999,N_22550,N_21976);
and U23000 (N_23000,N_22538,N_22593);
nor U23001 (N_23001,N_22232,N_22499);
nand U23002 (N_23002,N_22609,N_21773);
nand U23003 (N_23003,N_21864,N_22486);
xnor U23004 (N_23004,N_22108,N_21850);
and U23005 (N_23005,N_21739,N_22407);
nor U23006 (N_23006,N_22126,N_21766);
xor U23007 (N_23007,N_22207,N_22245);
xnor U23008 (N_23008,N_22150,N_21715);
and U23009 (N_23009,N_22686,N_22227);
and U23010 (N_23010,N_21630,N_21605);
xnor U23011 (N_23011,N_22489,N_22339);
xor U23012 (N_23012,N_21966,N_22173);
and U23013 (N_23013,N_22762,N_22350);
nor U23014 (N_23014,N_22259,N_22231);
nand U23015 (N_23015,N_22220,N_22296);
nand U23016 (N_23016,N_22250,N_22663);
nor U23017 (N_23017,N_22198,N_22443);
and U23018 (N_23018,N_22700,N_21676);
and U23019 (N_23019,N_22385,N_22072);
or U23020 (N_23020,N_22082,N_22371);
and U23021 (N_23021,N_22089,N_22616);
nand U23022 (N_23022,N_22267,N_22688);
nor U23023 (N_23023,N_22721,N_22447);
nand U23024 (N_23024,N_22176,N_22300);
xnor U23025 (N_23025,N_22057,N_22046);
or U23026 (N_23026,N_22290,N_21832);
and U23027 (N_23027,N_22308,N_22326);
nor U23028 (N_23028,N_22596,N_22345);
or U23029 (N_23029,N_21871,N_22650);
nor U23030 (N_23030,N_22053,N_22018);
and U23031 (N_23031,N_21623,N_22279);
nor U23032 (N_23032,N_22060,N_22787);
or U23033 (N_23033,N_22780,N_22388);
and U23034 (N_23034,N_21814,N_22591);
nand U23035 (N_23035,N_21963,N_21641);
or U23036 (N_23036,N_22068,N_22214);
xor U23037 (N_23037,N_21949,N_21771);
or U23038 (N_23038,N_21939,N_21744);
nor U23039 (N_23039,N_22697,N_21782);
or U23040 (N_23040,N_22623,N_22144);
xnor U23041 (N_23041,N_21737,N_22661);
or U23042 (N_23042,N_21987,N_22307);
xnor U23043 (N_23043,N_21785,N_22512);
nand U23044 (N_23044,N_22191,N_22714);
nor U23045 (N_23045,N_22073,N_22799);
nor U23046 (N_23046,N_21629,N_21717);
or U23047 (N_23047,N_22689,N_22303);
nand U23048 (N_23048,N_22592,N_21992);
or U23049 (N_23049,N_21862,N_22485);
xor U23050 (N_23050,N_21650,N_22340);
xor U23051 (N_23051,N_22562,N_22553);
xnor U23052 (N_23052,N_22256,N_21617);
and U23053 (N_23053,N_22648,N_21724);
nand U23054 (N_23054,N_22679,N_22272);
nor U23055 (N_23055,N_21654,N_21696);
nand U23056 (N_23056,N_22530,N_22506);
and U23057 (N_23057,N_22580,N_22393);
nand U23058 (N_23058,N_22767,N_22170);
xnor U23059 (N_23059,N_22237,N_22597);
nand U23060 (N_23060,N_21894,N_21917);
nand U23061 (N_23061,N_22772,N_22617);
nand U23062 (N_23062,N_21643,N_21993);
xnor U23063 (N_23063,N_22251,N_22233);
nor U23064 (N_23064,N_22149,N_22519);
nor U23065 (N_23065,N_22478,N_22090);
nand U23066 (N_23066,N_21999,N_22152);
and U23067 (N_23067,N_22384,N_21885);
or U23068 (N_23068,N_21678,N_22702);
and U23069 (N_23069,N_21898,N_22320);
and U23070 (N_23070,N_21818,N_21729);
nor U23071 (N_23071,N_21935,N_22564);
or U23072 (N_23072,N_21985,N_21844);
nand U23073 (N_23073,N_21665,N_22576);
or U23074 (N_23074,N_22130,N_22210);
nor U23075 (N_23075,N_22471,N_22632);
nor U23076 (N_23076,N_22483,N_21901);
xor U23077 (N_23077,N_22381,N_22099);
nand U23078 (N_23078,N_22504,N_22603);
nor U23079 (N_23079,N_21908,N_22081);
nor U23080 (N_23080,N_21775,N_22730);
and U23081 (N_23081,N_22337,N_21882);
and U23082 (N_23082,N_21689,N_22188);
and U23083 (N_23083,N_22479,N_22010);
and U23084 (N_23084,N_22263,N_22291);
or U23085 (N_23085,N_22247,N_22030);
or U23086 (N_23086,N_21996,N_22066);
or U23087 (N_23087,N_21881,N_21803);
xnor U23088 (N_23088,N_22273,N_21633);
nor U23089 (N_23089,N_22171,N_21903);
nand U23090 (N_23090,N_21918,N_21936);
nor U23091 (N_23091,N_21607,N_22464);
or U23092 (N_23092,N_21726,N_22695);
and U23093 (N_23093,N_22421,N_22026);
nand U23094 (N_23094,N_22779,N_22677);
or U23095 (N_23095,N_21889,N_22432);
xnor U23096 (N_23096,N_22347,N_21895);
nand U23097 (N_23097,N_22163,N_22131);
nand U23098 (N_23098,N_21793,N_22248);
nand U23099 (N_23099,N_22151,N_21872);
and U23100 (N_23100,N_22588,N_21642);
or U23101 (N_23101,N_22213,N_22392);
or U23102 (N_23102,N_21753,N_22354);
nand U23103 (N_23103,N_22007,N_21674);
nand U23104 (N_23104,N_22025,N_22703);
nor U23105 (N_23105,N_22008,N_22319);
and U23106 (N_23106,N_22221,N_22783);
or U23107 (N_23107,N_22396,N_22310);
nand U23108 (N_23108,N_22229,N_22301);
and U23109 (N_23109,N_22750,N_22005);
or U23110 (N_23110,N_21851,N_22241);
nor U23111 (N_23111,N_22520,N_21797);
nand U23112 (N_23112,N_22636,N_22052);
xnor U23113 (N_23113,N_22242,N_22751);
and U23114 (N_23114,N_22725,N_21747);
nor U23115 (N_23115,N_22160,N_22468);
nand U23116 (N_23116,N_22535,N_21940);
xor U23117 (N_23117,N_21915,N_22067);
nor U23118 (N_23118,N_22733,N_21849);
xor U23119 (N_23119,N_22095,N_22041);
nor U23120 (N_23120,N_22458,N_22634);
and U23121 (N_23121,N_22383,N_22642);
nor U23122 (N_23122,N_22143,N_22773);
and U23123 (N_23123,N_21748,N_22323);
nor U23124 (N_23124,N_22047,N_21876);
xor U23125 (N_23125,N_22343,N_22366);
and U23126 (N_23126,N_22349,N_21772);
nor U23127 (N_23127,N_22566,N_21660);
nor U23128 (N_23128,N_22031,N_22532);
or U23129 (N_23129,N_22219,N_22257);
nand U23130 (N_23130,N_21725,N_22056);
and U23131 (N_23131,N_22548,N_21880);
xor U23132 (N_23132,N_22120,N_21801);
nand U23133 (N_23133,N_22668,N_22395);
nand U23134 (N_23134,N_22711,N_22441);
xnor U23135 (N_23135,N_22561,N_22502);
xnor U23136 (N_23136,N_22039,N_22208);
nor U23137 (N_23137,N_22054,N_22035);
nor U23138 (N_23138,N_22110,N_21810);
nor U23139 (N_23139,N_22275,N_22077);
or U23140 (N_23140,N_22302,N_22760);
xor U23141 (N_23141,N_22044,N_21677);
xnor U23142 (N_23142,N_21877,N_21977);
xor U23143 (N_23143,N_22690,N_21835);
or U23144 (N_23144,N_22254,N_22552);
or U23145 (N_23145,N_22626,N_21611);
and U23146 (N_23146,N_21638,N_22051);
or U23147 (N_23147,N_22091,N_22153);
nand U23148 (N_23148,N_21778,N_21668);
nor U23149 (N_23149,N_22615,N_21720);
and U23150 (N_23150,N_21704,N_22712);
nor U23151 (N_23151,N_22048,N_21907);
nand U23152 (N_23152,N_21719,N_22545);
and U23153 (N_23153,N_21632,N_22753);
nor U23154 (N_23154,N_21695,N_21912);
nor U23155 (N_23155,N_22128,N_21781);
xnor U23156 (N_23156,N_21916,N_22139);
nor U23157 (N_23157,N_22049,N_21757);
or U23158 (N_23158,N_21767,N_22547);
and U23159 (N_23159,N_22737,N_21904);
and U23160 (N_23160,N_22604,N_22277);
and U23161 (N_23161,N_21727,N_22437);
xor U23162 (N_23162,N_22184,N_21741);
and U23163 (N_23163,N_22332,N_22425);
xnor U23164 (N_23164,N_22571,N_22643);
xnor U23165 (N_23165,N_21651,N_22752);
nand U23166 (N_23166,N_22034,N_22258);
nand U23167 (N_23167,N_22667,N_22590);
and U23168 (N_23168,N_22742,N_22086);
and U23169 (N_23169,N_22127,N_22078);
or U23170 (N_23170,N_21702,N_22718);
nand U23171 (N_23171,N_22106,N_21914);
or U23172 (N_23172,N_22496,N_22798);
xor U23173 (N_23173,N_21615,N_21687);
nor U23174 (N_23174,N_21837,N_22670);
or U23175 (N_23175,N_22651,N_22756);
xor U23176 (N_23176,N_22022,N_21640);
xor U23177 (N_23177,N_21610,N_22795);
nand U23178 (N_23178,N_21959,N_21620);
and U23179 (N_23179,N_22286,N_21701);
nor U23180 (N_23180,N_22665,N_22514);
nor U23181 (N_23181,N_21671,N_22197);
xor U23182 (N_23182,N_22551,N_22518);
or U23183 (N_23183,N_22278,N_21762);
xnor U23184 (N_23184,N_22631,N_21834);
nor U23185 (N_23185,N_22509,N_22311);
nor U23186 (N_23186,N_22065,N_22572);
xnor U23187 (N_23187,N_22608,N_22477);
nand U23188 (N_23188,N_22390,N_22640);
or U23189 (N_23189,N_21928,N_21645);
and U23190 (N_23190,N_22004,N_22778);
xor U23191 (N_23191,N_22037,N_22195);
xnor U23192 (N_23192,N_22589,N_22732);
nor U23193 (N_23193,N_22708,N_22775);
xnor U23194 (N_23194,N_21953,N_22462);
nor U23195 (N_23195,N_21890,N_21975);
nand U23196 (N_23196,N_21964,N_22582);
nand U23197 (N_23197,N_22304,N_22599);
or U23198 (N_23198,N_22016,N_22704);
nand U23199 (N_23199,N_22397,N_21731);
nor U23200 (N_23200,N_22461,N_21768);
and U23201 (N_23201,N_21858,N_21682);
xor U23202 (N_23202,N_21926,N_21683);
and U23203 (N_23203,N_21673,N_22252);
nor U23204 (N_23204,N_21913,N_21763);
nand U23205 (N_23205,N_21680,N_22306);
xnor U23206 (N_23206,N_22415,N_22657);
and U23207 (N_23207,N_21861,N_22298);
xnor U23208 (N_23208,N_21752,N_22420);
and U23209 (N_23209,N_22543,N_22457);
or U23210 (N_23210,N_22622,N_22546);
nand U23211 (N_23211,N_22467,N_22487);
and U23212 (N_23212,N_22230,N_22315);
or U23213 (N_23213,N_21972,N_22002);
nand U23214 (N_23214,N_21944,N_21732);
or U23215 (N_23215,N_21811,N_22028);
xnor U23216 (N_23216,N_22570,N_22413);
and U23217 (N_23217,N_21824,N_22001);
nand U23218 (N_23218,N_21873,N_21746);
nand U23219 (N_23219,N_21709,N_22338);
and U23220 (N_23220,N_22012,N_21800);
or U23221 (N_23221,N_22417,N_22312);
nor U23222 (N_23222,N_22715,N_21770);
nand U23223 (N_23223,N_22013,N_22630);
nor U23224 (N_23224,N_22314,N_22287);
and U23225 (N_23225,N_22470,N_22146);
and U23226 (N_23226,N_21792,N_22239);
xnor U23227 (N_23227,N_22567,N_22710);
and U23228 (N_23228,N_22755,N_21848);
or U23229 (N_23229,N_21902,N_22649);
nor U23230 (N_23230,N_22669,N_22454);
or U23231 (N_23231,N_22777,N_22180);
and U23232 (N_23232,N_21712,N_22192);
and U23233 (N_23233,N_21614,N_22351);
nor U23234 (N_23234,N_22406,N_21624);
and U23235 (N_23235,N_21979,N_22610);
and U23236 (N_23236,N_21946,N_22501);
and U23237 (N_23237,N_22113,N_21749);
or U23238 (N_23238,N_21967,N_22480);
nor U23239 (N_23239,N_21833,N_21860);
xnor U23240 (N_23240,N_22299,N_21613);
nand U23241 (N_23241,N_22070,N_22380);
or U23242 (N_23242,N_21973,N_21883);
and U23243 (N_23243,N_22059,N_21836);
and U23244 (N_23244,N_22598,N_21789);
xor U23245 (N_23245,N_21990,N_22382);
nor U23246 (N_23246,N_22342,N_22083);
nand U23247 (N_23247,N_21688,N_22671);
or U23248 (N_23248,N_21606,N_22776);
and U23249 (N_23249,N_22249,N_22473);
xor U23250 (N_23250,N_22446,N_22125);
nand U23251 (N_23251,N_22116,N_21958);
or U23252 (N_23252,N_21930,N_22364);
nor U23253 (N_23253,N_22024,N_22430);
nand U23254 (N_23254,N_22367,N_21699);
xnor U23255 (N_23255,N_22731,N_22274);
or U23256 (N_23256,N_22020,N_22040);
and U23257 (N_23257,N_21787,N_21662);
nor U23258 (N_23258,N_22785,N_22720);
nand U23259 (N_23259,N_22492,N_22295);
or U23260 (N_23260,N_22199,N_22736);
and U23261 (N_23261,N_22763,N_22211);
or U23262 (N_23262,N_22459,N_22368);
nand U23263 (N_23263,N_22408,N_22105);
nor U23264 (N_23264,N_22739,N_22355);
nor U23265 (N_23265,N_22579,N_22203);
nor U23266 (N_23266,N_21952,N_22466);
or U23267 (N_23267,N_21945,N_22159);
xnor U23268 (N_23268,N_22583,N_22568);
and U23269 (N_23269,N_22659,N_21932);
xnor U23270 (N_23270,N_22353,N_22293);
or U23271 (N_23271,N_22498,N_22507);
or U23272 (N_23272,N_21998,N_22745);
nand U23273 (N_23273,N_22165,N_22218);
xnor U23274 (N_23274,N_22418,N_22334);
and U23275 (N_23275,N_22370,N_21859);
xnor U23276 (N_23276,N_22563,N_21679);
nand U23277 (N_23277,N_22414,N_22225);
and U23278 (N_23278,N_22724,N_21899);
and U23279 (N_23279,N_22135,N_22270);
and U23280 (N_23280,N_22117,N_22185);
nor U23281 (N_23281,N_22043,N_21764);
xnor U23282 (N_23282,N_22662,N_22155);
nand U23283 (N_23283,N_22356,N_22680);
or U23284 (N_23284,N_22094,N_21826);
nor U23285 (N_23285,N_21708,N_22394);
or U23286 (N_23286,N_22761,N_22637);
and U23287 (N_23287,N_22136,N_22558);
and U23288 (N_23288,N_22664,N_21893);
and U23289 (N_23289,N_21761,N_22027);
nor U23290 (N_23290,N_22410,N_21934);
or U23291 (N_23291,N_22050,N_22525);
xor U23292 (N_23292,N_21618,N_22202);
nand U23293 (N_23293,N_21995,N_21900);
xnor U23294 (N_23294,N_21603,N_22734);
nor U23295 (N_23295,N_22009,N_22533);
or U23296 (N_23296,N_22109,N_22556);
nand U23297 (N_23297,N_22594,N_22600);
xnor U23298 (N_23298,N_21675,N_21779);
or U23299 (N_23299,N_21697,N_21991);
or U23300 (N_23300,N_22377,N_22103);
and U23301 (N_23301,N_21820,N_22265);
or U23302 (N_23302,N_21653,N_21670);
nor U23303 (N_23303,N_22445,N_21733);
and U23304 (N_23304,N_22373,N_21648);
nand U23305 (N_23305,N_21705,N_22625);
nand U23306 (N_23306,N_21743,N_22757);
and U23307 (N_23307,N_21924,N_22784);
nor U23308 (N_23308,N_22269,N_21831);
and U23309 (N_23309,N_21867,N_22003);
xnor U23310 (N_23310,N_22271,N_22102);
and U23311 (N_23311,N_21721,N_22015);
and U23312 (N_23312,N_22612,N_21841);
and U23313 (N_23313,N_21897,N_21962);
nor U23314 (N_23314,N_22379,N_22104);
xor U23315 (N_23315,N_22398,N_22652);
nor U23316 (N_23316,N_22614,N_22313);
nand U23317 (N_23317,N_22754,N_22029);
or U23318 (N_23318,N_22675,N_22521);
nor U23319 (N_23319,N_22074,N_22716);
and U23320 (N_23320,N_22111,N_22145);
and U23321 (N_23321,N_22681,N_22743);
nand U23322 (N_23322,N_22482,N_22574);
xnor U23323 (N_23323,N_22011,N_21943);
and U23324 (N_23324,N_21798,N_22653);
or U23325 (N_23325,N_22539,N_22542);
xor U23326 (N_23326,N_22427,N_21911);
nor U23327 (N_23327,N_22075,N_22452);
nor U23328 (N_23328,N_22386,N_22673);
nor U23329 (N_23329,N_22706,N_22209);
nor U23330 (N_23330,N_21997,N_22656);
xor U23331 (N_23331,N_22698,N_22329);
nor U23332 (N_23332,N_22114,N_21954);
or U23333 (N_23333,N_22196,N_22453);
and U23334 (N_23334,N_22123,N_22769);
nor U23335 (N_23335,N_21722,N_21809);
nor U23336 (N_23336,N_21965,N_21777);
and U23337 (N_23337,N_22789,N_22770);
nor U23338 (N_23338,N_21923,N_22189);
and U23339 (N_23339,N_22175,N_22497);
xnor U23340 (N_23340,N_21842,N_22322);
or U23341 (N_23341,N_22266,N_22488);
and U23342 (N_23342,N_21817,N_21714);
xor U23343 (N_23343,N_22494,N_22376);
nand U23344 (N_23344,N_22722,N_22476);
or U23345 (N_23345,N_21710,N_21664);
xor U23346 (N_23346,N_21866,N_22749);
nor U23347 (N_23347,N_22429,N_21875);
xnor U23348 (N_23348,N_22006,N_22455);
and U23349 (N_23349,N_22646,N_22791);
and U23350 (N_23350,N_22107,N_22569);
nor U23351 (N_23351,N_22362,N_21840);
nor U23352 (N_23352,N_21980,N_21758);
xnor U23353 (N_23353,N_21937,N_21742);
and U23354 (N_23354,N_21754,N_22726);
xnor U23355 (N_23355,N_22699,N_21738);
and U23356 (N_23356,N_22555,N_22719);
or U23357 (N_23357,N_22605,N_22124);
nand U23358 (N_23358,N_21794,N_22587);
nor U23359 (N_23359,N_21692,N_22162);
nor U23360 (N_23360,N_21807,N_22378);
or U23361 (N_23361,N_21627,N_21843);
and U23362 (N_23362,N_21879,N_22439);
and U23363 (N_23363,N_22537,N_22055);
or U23364 (N_23364,N_21921,N_21855);
nand U23365 (N_23365,N_22529,N_22797);
nor U23366 (N_23366,N_22222,N_22682);
nand U23367 (N_23367,N_22481,N_21622);
or U23368 (N_23368,N_22122,N_21713);
nand U23369 (N_23369,N_22627,N_22491);
xnor U23370 (N_23370,N_22595,N_22774);
xnor U23371 (N_23371,N_21927,N_22045);
or U23372 (N_23372,N_21852,N_22017);
or U23373 (N_23373,N_21635,N_22472);
and U23374 (N_23374,N_22493,N_22182);
nor U23375 (N_23375,N_22748,N_22360);
or U23376 (N_23376,N_22226,N_22692);
nand U23377 (N_23377,N_22336,N_22460);
nor U23378 (N_23378,N_22217,N_22261);
xor U23379 (N_23379,N_21647,N_21961);
nand U23380 (N_23380,N_22639,N_22678);
xor U23381 (N_23381,N_22285,N_22036);
nand U23382 (N_23382,N_22280,N_21609);
nor U23383 (N_23383,N_21791,N_22400);
or U23384 (N_23384,N_22166,N_22510);
and U23385 (N_23385,N_21971,N_22685);
xor U23386 (N_23386,N_22792,N_22448);
nor U23387 (N_23387,N_22244,N_21854);
or U23388 (N_23388,N_21804,N_21919);
nor U23389 (N_23389,N_22696,N_22305);
or U23390 (N_23390,N_22428,N_22119);
nor U23391 (N_23391,N_22294,N_22283);
or U23392 (N_23392,N_21863,N_21667);
or U23393 (N_23393,N_22062,N_22705);
xor U23394 (N_23394,N_22000,N_21870);
nand U23395 (N_23395,N_22655,N_21755);
nor U23396 (N_23396,N_21646,N_22440);
nor U23397 (N_23397,N_21968,N_22076);
nand U23398 (N_23398,N_21707,N_21828);
nor U23399 (N_23399,N_22728,N_21816);
or U23400 (N_23400,N_21630,N_21844);
nor U23401 (N_23401,N_22603,N_22019);
xnor U23402 (N_23402,N_21605,N_22007);
nand U23403 (N_23403,N_22369,N_22445);
or U23404 (N_23404,N_21640,N_22379);
nor U23405 (N_23405,N_21836,N_22183);
and U23406 (N_23406,N_21924,N_22204);
nand U23407 (N_23407,N_21793,N_22578);
or U23408 (N_23408,N_21752,N_21958);
and U23409 (N_23409,N_22588,N_21635);
nor U23410 (N_23410,N_21650,N_22404);
and U23411 (N_23411,N_22706,N_22088);
nor U23412 (N_23412,N_22592,N_21668);
nor U23413 (N_23413,N_22356,N_21776);
nor U23414 (N_23414,N_22024,N_21891);
xnor U23415 (N_23415,N_22257,N_22721);
xnor U23416 (N_23416,N_21970,N_21945);
nor U23417 (N_23417,N_22780,N_21656);
and U23418 (N_23418,N_21874,N_21638);
xnor U23419 (N_23419,N_22379,N_22497);
nand U23420 (N_23420,N_22477,N_22483);
nand U23421 (N_23421,N_22648,N_22465);
xor U23422 (N_23422,N_22313,N_21690);
nor U23423 (N_23423,N_22653,N_22269);
xnor U23424 (N_23424,N_21918,N_22179);
nor U23425 (N_23425,N_21935,N_21676);
xnor U23426 (N_23426,N_21786,N_21615);
nor U23427 (N_23427,N_21940,N_21958);
or U23428 (N_23428,N_22383,N_22016);
nor U23429 (N_23429,N_22168,N_21740);
nor U23430 (N_23430,N_22254,N_21897);
nor U23431 (N_23431,N_22747,N_22254);
and U23432 (N_23432,N_22144,N_22265);
nor U23433 (N_23433,N_22086,N_21870);
nor U23434 (N_23434,N_21795,N_22265);
xor U23435 (N_23435,N_22631,N_22423);
nand U23436 (N_23436,N_22020,N_22326);
or U23437 (N_23437,N_21738,N_21611);
xnor U23438 (N_23438,N_22653,N_21838);
nand U23439 (N_23439,N_21678,N_22021);
nor U23440 (N_23440,N_22210,N_21790);
or U23441 (N_23441,N_22756,N_22213);
nor U23442 (N_23442,N_22107,N_22080);
and U23443 (N_23443,N_22762,N_22298);
nand U23444 (N_23444,N_22043,N_22300);
and U23445 (N_23445,N_21810,N_22190);
nand U23446 (N_23446,N_22090,N_21615);
nor U23447 (N_23447,N_22719,N_21633);
xnor U23448 (N_23448,N_22667,N_21645);
or U23449 (N_23449,N_22748,N_22714);
or U23450 (N_23450,N_22096,N_21792);
nand U23451 (N_23451,N_22380,N_21984);
xnor U23452 (N_23452,N_22291,N_22698);
nand U23453 (N_23453,N_22329,N_21836);
xnor U23454 (N_23454,N_22094,N_22533);
or U23455 (N_23455,N_22138,N_22231);
or U23456 (N_23456,N_22320,N_21648);
and U23457 (N_23457,N_22026,N_22073);
nand U23458 (N_23458,N_21751,N_22286);
xnor U23459 (N_23459,N_22777,N_22320);
or U23460 (N_23460,N_22342,N_22343);
or U23461 (N_23461,N_22208,N_22259);
and U23462 (N_23462,N_21667,N_21932);
and U23463 (N_23463,N_22421,N_22139);
nor U23464 (N_23464,N_22260,N_22741);
xor U23465 (N_23465,N_22299,N_21863);
nand U23466 (N_23466,N_22711,N_22274);
nand U23467 (N_23467,N_21810,N_22459);
and U23468 (N_23468,N_21897,N_22356);
nor U23469 (N_23469,N_22792,N_22020);
xnor U23470 (N_23470,N_22307,N_21690);
or U23471 (N_23471,N_22058,N_22633);
and U23472 (N_23472,N_21965,N_22255);
or U23473 (N_23473,N_22208,N_21652);
or U23474 (N_23474,N_22649,N_21904);
and U23475 (N_23475,N_22032,N_22064);
and U23476 (N_23476,N_22543,N_22327);
and U23477 (N_23477,N_22214,N_22247);
nand U23478 (N_23478,N_22204,N_22056);
nand U23479 (N_23479,N_22672,N_22232);
nor U23480 (N_23480,N_21617,N_21700);
nor U23481 (N_23481,N_21604,N_21848);
xnor U23482 (N_23482,N_21882,N_22236);
or U23483 (N_23483,N_22462,N_22348);
or U23484 (N_23484,N_22336,N_22724);
and U23485 (N_23485,N_22226,N_21714);
and U23486 (N_23486,N_21743,N_22436);
nand U23487 (N_23487,N_22138,N_22056);
xor U23488 (N_23488,N_21918,N_22197);
nor U23489 (N_23489,N_22357,N_21878);
nand U23490 (N_23490,N_21801,N_21850);
nor U23491 (N_23491,N_22227,N_22484);
or U23492 (N_23492,N_22041,N_22234);
or U23493 (N_23493,N_22702,N_21863);
xor U23494 (N_23494,N_21897,N_22240);
nor U23495 (N_23495,N_21646,N_21871);
or U23496 (N_23496,N_22659,N_22363);
nor U23497 (N_23497,N_22325,N_22406);
nand U23498 (N_23498,N_22503,N_21836);
nand U23499 (N_23499,N_21731,N_22610);
or U23500 (N_23500,N_22519,N_22386);
xor U23501 (N_23501,N_21997,N_21693);
or U23502 (N_23502,N_22550,N_22560);
nor U23503 (N_23503,N_22493,N_22445);
nor U23504 (N_23504,N_22741,N_22701);
and U23505 (N_23505,N_21915,N_21669);
nor U23506 (N_23506,N_22521,N_22345);
xnor U23507 (N_23507,N_22172,N_21960);
nand U23508 (N_23508,N_22235,N_21741);
or U23509 (N_23509,N_21708,N_21610);
nand U23510 (N_23510,N_22703,N_22595);
and U23511 (N_23511,N_22699,N_21999);
or U23512 (N_23512,N_22512,N_21605);
nor U23513 (N_23513,N_22759,N_22271);
and U23514 (N_23514,N_21734,N_22233);
nand U23515 (N_23515,N_22773,N_22505);
nor U23516 (N_23516,N_22056,N_22454);
nor U23517 (N_23517,N_22451,N_22458);
or U23518 (N_23518,N_21914,N_22005);
xnor U23519 (N_23519,N_22170,N_21972);
xor U23520 (N_23520,N_21612,N_22619);
and U23521 (N_23521,N_21943,N_22289);
or U23522 (N_23522,N_22420,N_21716);
xnor U23523 (N_23523,N_22551,N_22633);
nand U23524 (N_23524,N_22477,N_22542);
nand U23525 (N_23525,N_22699,N_21776);
nand U23526 (N_23526,N_22021,N_22460);
and U23527 (N_23527,N_22045,N_21630);
nand U23528 (N_23528,N_21958,N_22144);
and U23529 (N_23529,N_22194,N_22090);
nor U23530 (N_23530,N_22084,N_22598);
nand U23531 (N_23531,N_22295,N_21646);
or U23532 (N_23532,N_21789,N_22455);
nand U23533 (N_23533,N_22680,N_22127);
or U23534 (N_23534,N_22469,N_21647);
or U23535 (N_23535,N_22256,N_22340);
xor U23536 (N_23536,N_22206,N_22541);
nor U23537 (N_23537,N_21959,N_21904);
xor U23538 (N_23538,N_21759,N_21988);
xnor U23539 (N_23539,N_22040,N_22013);
or U23540 (N_23540,N_22737,N_22341);
nand U23541 (N_23541,N_22039,N_22711);
nand U23542 (N_23542,N_22196,N_22058);
and U23543 (N_23543,N_22595,N_21989);
and U23544 (N_23544,N_21995,N_21750);
and U23545 (N_23545,N_21718,N_22602);
xnor U23546 (N_23546,N_22355,N_22383);
or U23547 (N_23547,N_21936,N_22307);
xnor U23548 (N_23548,N_21868,N_22507);
xor U23549 (N_23549,N_22709,N_22686);
nand U23550 (N_23550,N_22413,N_22303);
and U23551 (N_23551,N_21792,N_22234);
nor U23552 (N_23552,N_22550,N_22216);
or U23553 (N_23553,N_22515,N_22431);
nor U23554 (N_23554,N_22784,N_22786);
xor U23555 (N_23555,N_21938,N_22090);
and U23556 (N_23556,N_22218,N_21899);
nand U23557 (N_23557,N_22350,N_21926);
and U23558 (N_23558,N_21978,N_22564);
and U23559 (N_23559,N_22216,N_22042);
nand U23560 (N_23560,N_22690,N_22495);
xor U23561 (N_23561,N_22497,N_21770);
xnor U23562 (N_23562,N_22780,N_22061);
xnor U23563 (N_23563,N_22097,N_21860);
nor U23564 (N_23564,N_21669,N_22294);
nand U23565 (N_23565,N_22691,N_22438);
nand U23566 (N_23566,N_22023,N_22181);
nor U23567 (N_23567,N_22122,N_22072);
or U23568 (N_23568,N_22387,N_21800);
xor U23569 (N_23569,N_22488,N_22714);
or U23570 (N_23570,N_22271,N_22502);
xnor U23571 (N_23571,N_22352,N_22193);
or U23572 (N_23572,N_22496,N_21919);
xnor U23573 (N_23573,N_22765,N_22563);
and U23574 (N_23574,N_22337,N_22136);
nand U23575 (N_23575,N_22693,N_22372);
xnor U23576 (N_23576,N_22056,N_22575);
or U23577 (N_23577,N_22152,N_22070);
xor U23578 (N_23578,N_22794,N_22775);
nand U23579 (N_23579,N_21732,N_22076);
xor U23580 (N_23580,N_21738,N_22308);
and U23581 (N_23581,N_21776,N_21886);
xor U23582 (N_23582,N_22590,N_22009);
or U23583 (N_23583,N_22387,N_22676);
xor U23584 (N_23584,N_21997,N_22519);
nor U23585 (N_23585,N_21873,N_21789);
xnor U23586 (N_23586,N_21917,N_22326);
xnor U23587 (N_23587,N_22221,N_21749);
and U23588 (N_23588,N_22228,N_22243);
xor U23589 (N_23589,N_22115,N_22420);
and U23590 (N_23590,N_21709,N_21650);
and U23591 (N_23591,N_22783,N_22692);
and U23592 (N_23592,N_21758,N_22223);
or U23593 (N_23593,N_22460,N_22500);
or U23594 (N_23594,N_21700,N_22347);
nor U23595 (N_23595,N_21871,N_21866);
and U23596 (N_23596,N_21929,N_22686);
nor U23597 (N_23597,N_22182,N_22301);
xnor U23598 (N_23598,N_22552,N_21778);
nand U23599 (N_23599,N_22256,N_22073);
xor U23600 (N_23600,N_22670,N_22621);
and U23601 (N_23601,N_22308,N_22376);
or U23602 (N_23602,N_22272,N_22435);
or U23603 (N_23603,N_21752,N_22529);
nor U23604 (N_23604,N_22314,N_22026);
and U23605 (N_23605,N_22111,N_21715);
xor U23606 (N_23606,N_22109,N_22010);
nand U23607 (N_23607,N_22575,N_21909);
xor U23608 (N_23608,N_22164,N_22041);
xnor U23609 (N_23609,N_22376,N_22200);
or U23610 (N_23610,N_21939,N_21630);
nand U23611 (N_23611,N_22631,N_22171);
or U23612 (N_23612,N_21743,N_21696);
xor U23613 (N_23613,N_22536,N_22144);
and U23614 (N_23614,N_22733,N_22524);
and U23615 (N_23615,N_22605,N_22138);
xnor U23616 (N_23616,N_22689,N_22080);
or U23617 (N_23617,N_21846,N_22361);
or U23618 (N_23618,N_21981,N_22127);
nor U23619 (N_23619,N_22547,N_22063);
or U23620 (N_23620,N_22008,N_22068);
xnor U23621 (N_23621,N_21857,N_22472);
nand U23622 (N_23622,N_22355,N_21933);
nor U23623 (N_23623,N_22651,N_22699);
nor U23624 (N_23624,N_22318,N_22110);
or U23625 (N_23625,N_22541,N_22363);
nand U23626 (N_23626,N_21937,N_22421);
nand U23627 (N_23627,N_21777,N_22161);
or U23628 (N_23628,N_22601,N_21791);
nand U23629 (N_23629,N_21688,N_22609);
or U23630 (N_23630,N_22325,N_21906);
or U23631 (N_23631,N_22264,N_22080);
or U23632 (N_23632,N_22695,N_22443);
and U23633 (N_23633,N_21760,N_21658);
nor U23634 (N_23634,N_22586,N_22472);
nor U23635 (N_23635,N_21797,N_22335);
xnor U23636 (N_23636,N_22587,N_22248);
and U23637 (N_23637,N_21971,N_22399);
or U23638 (N_23638,N_22581,N_21954);
and U23639 (N_23639,N_21833,N_21756);
xor U23640 (N_23640,N_22621,N_21935);
or U23641 (N_23641,N_22264,N_21767);
xnor U23642 (N_23642,N_22005,N_22568);
or U23643 (N_23643,N_22314,N_22703);
xnor U23644 (N_23644,N_22218,N_22201);
xor U23645 (N_23645,N_22260,N_22189);
and U23646 (N_23646,N_22325,N_21979);
and U23647 (N_23647,N_22206,N_22621);
and U23648 (N_23648,N_21816,N_22090);
nor U23649 (N_23649,N_22385,N_22774);
xnor U23650 (N_23650,N_21996,N_21884);
nand U23651 (N_23651,N_21857,N_22310);
nand U23652 (N_23652,N_22613,N_22021);
nand U23653 (N_23653,N_22068,N_22760);
nand U23654 (N_23654,N_22079,N_21713);
or U23655 (N_23655,N_22685,N_21648);
xnor U23656 (N_23656,N_22003,N_22074);
and U23657 (N_23657,N_22145,N_22203);
nor U23658 (N_23658,N_22617,N_21808);
and U23659 (N_23659,N_22239,N_22156);
or U23660 (N_23660,N_21811,N_21721);
nor U23661 (N_23661,N_21634,N_22744);
or U23662 (N_23662,N_21689,N_21862);
or U23663 (N_23663,N_21705,N_22353);
nand U23664 (N_23664,N_21658,N_21939);
xnor U23665 (N_23665,N_21814,N_22332);
and U23666 (N_23666,N_21778,N_22398);
nor U23667 (N_23667,N_22138,N_22069);
and U23668 (N_23668,N_21745,N_22074);
nor U23669 (N_23669,N_22697,N_22087);
or U23670 (N_23670,N_21674,N_22620);
nand U23671 (N_23671,N_22763,N_22366);
nand U23672 (N_23672,N_22302,N_22309);
nand U23673 (N_23673,N_22115,N_22059);
or U23674 (N_23674,N_21824,N_21889);
or U23675 (N_23675,N_21827,N_22156);
and U23676 (N_23676,N_22043,N_22457);
xor U23677 (N_23677,N_22416,N_22295);
xnor U23678 (N_23678,N_21825,N_21963);
nor U23679 (N_23679,N_22307,N_21663);
or U23680 (N_23680,N_22757,N_22288);
and U23681 (N_23681,N_22448,N_22281);
nor U23682 (N_23682,N_22513,N_21703);
xor U23683 (N_23683,N_22368,N_21752);
or U23684 (N_23684,N_22486,N_21808);
xor U23685 (N_23685,N_21913,N_22042);
xnor U23686 (N_23686,N_22644,N_22512);
xor U23687 (N_23687,N_22668,N_22522);
or U23688 (N_23688,N_22757,N_22583);
and U23689 (N_23689,N_22149,N_22567);
or U23690 (N_23690,N_21654,N_22771);
and U23691 (N_23691,N_22219,N_21742);
xor U23692 (N_23692,N_22425,N_21851);
and U23693 (N_23693,N_21992,N_21812);
and U23694 (N_23694,N_22351,N_22799);
and U23695 (N_23695,N_22627,N_22496);
and U23696 (N_23696,N_22312,N_22797);
or U23697 (N_23697,N_21644,N_22281);
xnor U23698 (N_23698,N_21630,N_22009);
or U23699 (N_23699,N_22285,N_22130);
and U23700 (N_23700,N_21927,N_21758);
and U23701 (N_23701,N_22110,N_21745);
nand U23702 (N_23702,N_22643,N_21736);
nor U23703 (N_23703,N_22652,N_22661);
and U23704 (N_23704,N_22368,N_21929);
nor U23705 (N_23705,N_21929,N_21946);
nand U23706 (N_23706,N_21612,N_22337);
nor U23707 (N_23707,N_21873,N_22636);
or U23708 (N_23708,N_22513,N_22275);
or U23709 (N_23709,N_22374,N_22158);
or U23710 (N_23710,N_22613,N_22081);
nand U23711 (N_23711,N_22263,N_21954);
and U23712 (N_23712,N_22677,N_22489);
nor U23713 (N_23713,N_21895,N_22469);
and U23714 (N_23714,N_21892,N_22523);
nor U23715 (N_23715,N_22746,N_21666);
nor U23716 (N_23716,N_22798,N_22211);
nor U23717 (N_23717,N_21773,N_22404);
xor U23718 (N_23718,N_21846,N_21758);
xor U23719 (N_23719,N_21913,N_22785);
nor U23720 (N_23720,N_21961,N_21608);
nand U23721 (N_23721,N_22688,N_22371);
nor U23722 (N_23722,N_22340,N_22143);
nand U23723 (N_23723,N_21717,N_21898);
or U23724 (N_23724,N_22552,N_22483);
nand U23725 (N_23725,N_21761,N_21777);
and U23726 (N_23726,N_21612,N_22300);
or U23727 (N_23727,N_21828,N_22394);
and U23728 (N_23728,N_22509,N_22736);
and U23729 (N_23729,N_22334,N_22601);
or U23730 (N_23730,N_21733,N_22301);
or U23731 (N_23731,N_22739,N_21767);
or U23732 (N_23732,N_22552,N_22398);
nor U23733 (N_23733,N_21912,N_22115);
nor U23734 (N_23734,N_22445,N_21916);
nor U23735 (N_23735,N_22176,N_22197);
or U23736 (N_23736,N_22661,N_21675);
xor U23737 (N_23737,N_21893,N_22236);
xor U23738 (N_23738,N_21724,N_22300);
nor U23739 (N_23739,N_21711,N_22356);
or U23740 (N_23740,N_21851,N_22305);
nor U23741 (N_23741,N_21865,N_22384);
xnor U23742 (N_23742,N_21868,N_21846);
xnor U23743 (N_23743,N_21773,N_22009);
nor U23744 (N_23744,N_21853,N_22171);
nor U23745 (N_23745,N_22261,N_21884);
and U23746 (N_23746,N_22343,N_22540);
xor U23747 (N_23747,N_21773,N_22050);
nand U23748 (N_23748,N_21977,N_22465);
nand U23749 (N_23749,N_22084,N_21981);
nand U23750 (N_23750,N_21806,N_22206);
nand U23751 (N_23751,N_22650,N_21699);
nor U23752 (N_23752,N_22233,N_21760);
xnor U23753 (N_23753,N_21634,N_21809);
nor U23754 (N_23754,N_22630,N_22221);
and U23755 (N_23755,N_22687,N_21948);
and U23756 (N_23756,N_21671,N_22114);
nor U23757 (N_23757,N_22553,N_22773);
and U23758 (N_23758,N_22022,N_21849);
nor U23759 (N_23759,N_21772,N_22411);
xnor U23760 (N_23760,N_22277,N_22761);
nand U23761 (N_23761,N_21708,N_21738);
nand U23762 (N_23762,N_22328,N_22191);
nor U23763 (N_23763,N_22321,N_21908);
nand U23764 (N_23764,N_21658,N_21978);
and U23765 (N_23765,N_22585,N_21744);
and U23766 (N_23766,N_22396,N_21825);
xnor U23767 (N_23767,N_22406,N_22541);
xor U23768 (N_23768,N_22353,N_21911);
nand U23769 (N_23769,N_22653,N_22790);
and U23770 (N_23770,N_21776,N_22578);
xor U23771 (N_23771,N_22302,N_22471);
nor U23772 (N_23772,N_22296,N_22176);
and U23773 (N_23773,N_22120,N_22433);
nand U23774 (N_23774,N_22773,N_21766);
or U23775 (N_23775,N_22141,N_21635);
or U23776 (N_23776,N_21652,N_22557);
or U23777 (N_23777,N_22340,N_22122);
or U23778 (N_23778,N_22156,N_21931);
nand U23779 (N_23779,N_22558,N_22373);
and U23780 (N_23780,N_22729,N_22084);
or U23781 (N_23781,N_22604,N_22054);
or U23782 (N_23782,N_22774,N_22534);
or U23783 (N_23783,N_22232,N_22019);
nand U23784 (N_23784,N_22720,N_22228);
xnor U23785 (N_23785,N_22140,N_22077);
nand U23786 (N_23786,N_22536,N_21670);
nand U23787 (N_23787,N_22184,N_21747);
nor U23788 (N_23788,N_22199,N_22658);
and U23789 (N_23789,N_21829,N_22155);
nor U23790 (N_23790,N_22623,N_22551);
nand U23791 (N_23791,N_22548,N_21981);
nand U23792 (N_23792,N_22184,N_21841);
nand U23793 (N_23793,N_22685,N_22142);
and U23794 (N_23794,N_22117,N_22133);
nor U23795 (N_23795,N_22797,N_21774);
nor U23796 (N_23796,N_22740,N_21894);
nor U23797 (N_23797,N_21836,N_22709);
nor U23798 (N_23798,N_22537,N_21851);
nor U23799 (N_23799,N_22242,N_21872);
or U23800 (N_23800,N_21990,N_22578);
nor U23801 (N_23801,N_21740,N_22123);
xnor U23802 (N_23802,N_21882,N_22389);
nor U23803 (N_23803,N_22284,N_22144);
and U23804 (N_23804,N_22239,N_22226);
xnor U23805 (N_23805,N_21957,N_22508);
nand U23806 (N_23806,N_22649,N_21676);
and U23807 (N_23807,N_22149,N_22658);
nand U23808 (N_23808,N_22175,N_22659);
nand U23809 (N_23809,N_22432,N_22787);
xnor U23810 (N_23810,N_22718,N_21798);
xor U23811 (N_23811,N_22467,N_21673);
xor U23812 (N_23812,N_22032,N_22471);
xnor U23813 (N_23813,N_22199,N_22165);
nor U23814 (N_23814,N_22323,N_21860);
nand U23815 (N_23815,N_22484,N_22440);
xor U23816 (N_23816,N_21720,N_21917);
xor U23817 (N_23817,N_21816,N_22777);
nand U23818 (N_23818,N_21741,N_22751);
and U23819 (N_23819,N_22516,N_22496);
nor U23820 (N_23820,N_22088,N_22652);
or U23821 (N_23821,N_21942,N_22361);
xnor U23822 (N_23822,N_22100,N_21991);
xnor U23823 (N_23823,N_22249,N_22653);
nor U23824 (N_23824,N_22428,N_22776);
or U23825 (N_23825,N_22586,N_22520);
nor U23826 (N_23826,N_22195,N_21946);
nand U23827 (N_23827,N_22580,N_21998);
xnor U23828 (N_23828,N_22301,N_22003);
or U23829 (N_23829,N_22581,N_21811);
or U23830 (N_23830,N_22128,N_22552);
or U23831 (N_23831,N_22202,N_21989);
nand U23832 (N_23832,N_22157,N_22132);
and U23833 (N_23833,N_21744,N_22399);
nand U23834 (N_23834,N_21847,N_22214);
nor U23835 (N_23835,N_22177,N_22030);
and U23836 (N_23836,N_22276,N_22732);
xnor U23837 (N_23837,N_21989,N_21967);
or U23838 (N_23838,N_22436,N_22200);
nor U23839 (N_23839,N_22672,N_22493);
or U23840 (N_23840,N_22337,N_22295);
or U23841 (N_23841,N_21723,N_22316);
and U23842 (N_23842,N_21900,N_22253);
or U23843 (N_23843,N_21921,N_22248);
xor U23844 (N_23844,N_22364,N_22353);
and U23845 (N_23845,N_21753,N_21749);
and U23846 (N_23846,N_22795,N_21818);
nor U23847 (N_23847,N_22272,N_21891);
nor U23848 (N_23848,N_21972,N_22641);
or U23849 (N_23849,N_22317,N_21678);
or U23850 (N_23850,N_21939,N_22044);
nand U23851 (N_23851,N_22171,N_21636);
xnor U23852 (N_23852,N_21760,N_21834);
nor U23853 (N_23853,N_22565,N_22323);
and U23854 (N_23854,N_22769,N_21966);
nor U23855 (N_23855,N_21964,N_21912);
nand U23856 (N_23856,N_22103,N_22319);
xnor U23857 (N_23857,N_21810,N_22194);
xor U23858 (N_23858,N_22795,N_22548);
xnor U23859 (N_23859,N_21918,N_21691);
nor U23860 (N_23860,N_22448,N_22240);
xnor U23861 (N_23861,N_22320,N_21798);
nand U23862 (N_23862,N_22591,N_21822);
and U23863 (N_23863,N_22582,N_22267);
or U23864 (N_23864,N_22720,N_21621);
or U23865 (N_23865,N_21791,N_21835);
xor U23866 (N_23866,N_21781,N_21740);
nand U23867 (N_23867,N_22560,N_22473);
xor U23868 (N_23868,N_22282,N_22445);
xnor U23869 (N_23869,N_21971,N_22064);
and U23870 (N_23870,N_22298,N_22745);
or U23871 (N_23871,N_21658,N_22705);
or U23872 (N_23872,N_22116,N_22508);
xnor U23873 (N_23873,N_22511,N_22299);
or U23874 (N_23874,N_22110,N_22578);
or U23875 (N_23875,N_22667,N_21986);
and U23876 (N_23876,N_22451,N_21678);
xnor U23877 (N_23877,N_22089,N_22790);
or U23878 (N_23878,N_21856,N_22731);
nor U23879 (N_23879,N_22347,N_22621);
xor U23880 (N_23880,N_22485,N_22420);
nor U23881 (N_23881,N_21665,N_21767);
nand U23882 (N_23882,N_22695,N_22405);
and U23883 (N_23883,N_22040,N_22411);
nor U23884 (N_23884,N_22601,N_22645);
nand U23885 (N_23885,N_22465,N_22012);
nand U23886 (N_23886,N_22536,N_21967);
nor U23887 (N_23887,N_22015,N_22056);
xnor U23888 (N_23888,N_22318,N_22377);
xnor U23889 (N_23889,N_22544,N_21728);
nor U23890 (N_23890,N_22109,N_22773);
xnor U23891 (N_23891,N_21797,N_21629);
nand U23892 (N_23892,N_22003,N_22288);
or U23893 (N_23893,N_21773,N_22787);
nand U23894 (N_23894,N_22662,N_21702);
xor U23895 (N_23895,N_22287,N_22711);
and U23896 (N_23896,N_21770,N_22705);
nor U23897 (N_23897,N_21914,N_22277);
nor U23898 (N_23898,N_22034,N_22576);
nor U23899 (N_23899,N_22303,N_22655);
nand U23900 (N_23900,N_22313,N_22182);
and U23901 (N_23901,N_21772,N_21909);
nor U23902 (N_23902,N_21825,N_21822);
nor U23903 (N_23903,N_21641,N_22354);
and U23904 (N_23904,N_22359,N_21651);
xnor U23905 (N_23905,N_22778,N_21659);
xor U23906 (N_23906,N_21727,N_22591);
nor U23907 (N_23907,N_22469,N_22235);
nor U23908 (N_23908,N_21658,N_22683);
nand U23909 (N_23909,N_21673,N_22736);
nand U23910 (N_23910,N_21685,N_21785);
xor U23911 (N_23911,N_22537,N_21718);
and U23912 (N_23912,N_21946,N_22639);
and U23913 (N_23913,N_21616,N_22419);
xor U23914 (N_23914,N_22761,N_22149);
xnor U23915 (N_23915,N_22207,N_22368);
xor U23916 (N_23916,N_21734,N_22236);
nand U23917 (N_23917,N_22422,N_22108);
nand U23918 (N_23918,N_21640,N_21651);
or U23919 (N_23919,N_22124,N_22649);
or U23920 (N_23920,N_22117,N_22423);
and U23921 (N_23921,N_22605,N_22797);
nor U23922 (N_23922,N_21754,N_22126);
xor U23923 (N_23923,N_22008,N_21755);
xor U23924 (N_23924,N_22573,N_22447);
and U23925 (N_23925,N_22376,N_21894);
xnor U23926 (N_23926,N_22156,N_22247);
nor U23927 (N_23927,N_21747,N_22600);
nand U23928 (N_23928,N_21827,N_21714);
or U23929 (N_23929,N_22786,N_22112);
nor U23930 (N_23930,N_22570,N_22546);
and U23931 (N_23931,N_22669,N_22420);
nand U23932 (N_23932,N_21839,N_22390);
and U23933 (N_23933,N_22391,N_22609);
or U23934 (N_23934,N_22116,N_21910);
nor U23935 (N_23935,N_21968,N_22019);
nor U23936 (N_23936,N_22400,N_22188);
or U23937 (N_23937,N_22178,N_22353);
nand U23938 (N_23938,N_22404,N_22139);
nor U23939 (N_23939,N_22161,N_21845);
nor U23940 (N_23940,N_22715,N_22653);
or U23941 (N_23941,N_22047,N_22100);
or U23942 (N_23942,N_22110,N_22236);
nand U23943 (N_23943,N_22712,N_21835);
nand U23944 (N_23944,N_22388,N_22778);
nor U23945 (N_23945,N_22122,N_22674);
nor U23946 (N_23946,N_22613,N_22031);
nor U23947 (N_23947,N_22431,N_22248);
nand U23948 (N_23948,N_22715,N_22633);
nand U23949 (N_23949,N_22594,N_22714);
xor U23950 (N_23950,N_21957,N_21968);
nor U23951 (N_23951,N_22552,N_21803);
or U23952 (N_23952,N_21881,N_22585);
nand U23953 (N_23953,N_22434,N_22751);
and U23954 (N_23954,N_22738,N_21799);
nor U23955 (N_23955,N_21736,N_21698);
nor U23956 (N_23956,N_22273,N_21889);
nor U23957 (N_23957,N_22578,N_21804);
xnor U23958 (N_23958,N_21667,N_21707);
nand U23959 (N_23959,N_22632,N_22642);
nand U23960 (N_23960,N_22628,N_21850);
nor U23961 (N_23961,N_22168,N_21711);
nor U23962 (N_23962,N_22271,N_22562);
nand U23963 (N_23963,N_21843,N_21774);
xnor U23964 (N_23964,N_22650,N_22716);
or U23965 (N_23965,N_22300,N_22531);
and U23966 (N_23966,N_22512,N_21864);
nand U23967 (N_23967,N_21707,N_22176);
and U23968 (N_23968,N_21825,N_22111);
nand U23969 (N_23969,N_22457,N_22083);
nor U23970 (N_23970,N_21959,N_22610);
and U23971 (N_23971,N_22477,N_22350);
nand U23972 (N_23972,N_22355,N_22127);
or U23973 (N_23973,N_22338,N_21720);
and U23974 (N_23974,N_22186,N_22637);
and U23975 (N_23975,N_22766,N_21952);
or U23976 (N_23976,N_21956,N_22637);
xor U23977 (N_23977,N_22566,N_21869);
xor U23978 (N_23978,N_22111,N_21886);
and U23979 (N_23979,N_22057,N_22326);
nand U23980 (N_23980,N_22242,N_22069);
nand U23981 (N_23981,N_21683,N_22625);
or U23982 (N_23982,N_21659,N_22135);
and U23983 (N_23983,N_22554,N_21730);
xor U23984 (N_23984,N_22673,N_22183);
nand U23985 (N_23985,N_22329,N_22552);
xor U23986 (N_23986,N_22036,N_22031);
nand U23987 (N_23987,N_22497,N_21851);
nor U23988 (N_23988,N_22320,N_22483);
or U23989 (N_23989,N_22266,N_22502);
nand U23990 (N_23990,N_21891,N_22160);
nor U23991 (N_23991,N_21949,N_22356);
xor U23992 (N_23992,N_22736,N_22240);
nor U23993 (N_23993,N_21763,N_22058);
nand U23994 (N_23994,N_22694,N_21935);
nor U23995 (N_23995,N_21978,N_22194);
nor U23996 (N_23996,N_21619,N_22493);
and U23997 (N_23997,N_22187,N_22565);
or U23998 (N_23998,N_21771,N_22360);
or U23999 (N_23999,N_22174,N_22167);
nor U24000 (N_24000,N_23328,N_23582);
nor U24001 (N_24001,N_22898,N_23021);
xor U24002 (N_24002,N_23144,N_23827);
xnor U24003 (N_24003,N_23624,N_22839);
nand U24004 (N_24004,N_23033,N_23937);
nand U24005 (N_24005,N_23704,N_23526);
nand U24006 (N_24006,N_23335,N_23226);
and U24007 (N_24007,N_23185,N_23364);
xnor U24008 (N_24008,N_23622,N_22862);
nand U24009 (N_24009,N_23732,N_23849);
xnor U24010 (N_24010,N_23797,N_23778);
or U24011 (N_24011,N_23087,N_23259);
and U24012 (N_24012,N_23352,N_23479);
or U24013 (N_24013,N_23942,N_23320);
or U24014 (N_24014,N_23971,N_23260);
nor U24015 (N_24015,N_22879,N_22903);
or U24016 (N_24016,N_22918,N_22951);
or U24017 (N_24017,N_23857,N_23264);
or U24018 (N_24018,N_23903,N_23905);
xor U24019 (N_24019,N_23672,N_23785);
nor U24020 (N_24020,N_22856,N_23366);
nor U24021 (N_24021,N_22958,N_23899);
nor U24022 (N_24022,N_23691,N_23040);
xnor U24023 (N_24023,N_23728,N_23554);
nor U24024 (N_24024,N_23338,N_23140);
nor U24025 (N_24025,N_23263,N_23161);
nand U24026 (N_24026,N_23451,N_23434);
and U24027 (N_24027,N_23463,N_23080);
and U24028 (N_24028,N_23841,N_23870);
nand U24029 (N_24029,N_23314,N_23201);
nand U24030 (N_24030,N_23074,N_22847);
and U24031 (N_24031,N_23138,N_22866);
nor U24032 (N_24032,N_23085,N_23294);
nand U24033 (N_24033,N_23025,N_23030);
or U24034 (N_24034,N_23362,N_23258);
or U24035 (N_24035,N_23315,N_23938);
nand U24036 (N_24036,N_23754,N_23324);
xor U24037 (N_24037,N_23823,N_23141);
and U24038 (N_24038,N_23219,N_23643);
nand U24039 (N_24039,N_23867,N_22973);
nor U24040 (N_24040,N_23255,N_23012);
nor U24041 (N_24041,N_23218,N_23664);
or U24042 (N_24042,N_23380,N_23117);
nor U24043 (N_24043,N_23828,N_23336);
or U24044 (N_24044,N_23099,N_22960);
or U24045 (N_24045,N_22977,N_23344);
or U24046 (N_24046,N_22886,N_23330);
xor U24047 (N_24047,N_23319,N_23019);
nand U24048 (N_24048,N_23415,N_23641);
and U24049 (N_24049,N_22873,N_23859);
nand U24050 (N_24050,N_23091,N_23714);
nor U24051 (N_24051,N_23274,N_23240);
or U24052 (N_24052,N_23963,N_23855);
xor U24053 (N_24053,N_23733,N_23498);
and U24054 (N_24054,N_23084,N_23716);
or U24055 (N_24055,N_23408,N_23375);
and U24056 (N_24056,N_23273,N_23097);
and U24057 (N_24057,N_23003,N_23900);
nand U24058 (N_24058,N_23647,N_23172);
nor U24059 (N_24059,N_23946,N_23383);
and U24060 (N_24060,N_23460,N_23416);
or U24061 (N_24061,N_23165,N_23835);
nand U24062 (N_24062,N_23029,N_22806);
xor U24063 (N_24063,N_23960,N_22831);
or U24064 (N_24064,N_23514,N_23974);
and U24065 (N_24065,N_23384,N_23035);
nand U24066 (N_24066,N_22822,N_23904);
or U24067 (N_24067,N_23048,N_23548);
and U24068 (N_24068,N_23277,N_23500);
or U24069 (N_24069,N_23764,N_23881);
nand U24070 (N_24070,N_23478,N_22966);
and U24071 (N_24071,N_23129,N_23148);
nand U24072 (N_24072,N_23822,N_23678);
nand U24073 (N_24073,N_22825,N_23627);
nand U24074 (N_24074,N_23155,N_23568);
nand U24075 (N_24075,N_23300,N_23756);
nand U24076 (N_24076,N_23312,N_23353);
or U24077 (N_24077,N_22957,N_23707);
nor U24078 (N_24078,N_23605,N_23923);
xor U24079 (N_24079,N_23351,N_23819);
xnor U24080 (N_24080,N_23020,N_23565);
nand U24081 (N_24081,N_23360,N_23102);
and U24082 (N_24082,N_22816,N_22889);
and U24083 (N_24083,N_22930,N_23875);
nor U24084 (N_24084,N_23382,N_23788);
nor U24085 (N_24085,N_23598,N_23023);
and U24086 (N_24086,N_22990,N_23028);
and U24087 (N_24087,N_23958,N_23615);
and U24088 (N_24088,N_23735,N_23246);
nor U24089 (N_24089,N_23537,N_23008);
nor U24090 (N_24090,N_23729,N_23781);
nor U24091 (N_24091,N_23722,N_22875);
nor U24092 (N_24092,N_23513,N_22907);
xnor U24093 (N_24093,N_22902,N_23724);
or U24094 (N_24094,N_23913,N_23053);
or U24095 (N_24095,N_23430,N_23474);
xnor U24096 (N_24096,N_23492,N_23060);
or U24097 (N_24097,N_23531,N_23342);
nor U24098 (N_24098,N_23317,N_23614);
and U24099 (N_24099,N_23794,N_23107);
and U24100 (N_24100,N_23517,N_23066);
or U24101 (N_24101,N_23313,N_22858);
and U24102 (N_24102,N_23755,N_23578);
or U24103 (N_24103,N_23447,N_22919);
or U24104 (N_24104,N_22987,N_23136);
and U24105 (N_24105,N_23972,N_23295);
and U24106 (N_24106,N_23638,N_22859);
xor U24107 (N_24107,N_23297,N_23431);
and U24108 (N_24108,N_23372,N_23907);
or U24109 (N_24109,N_23697,N_23190);
xor U24110 (N_24110,N_23385,N_23202);
and U24111 (N_24111,N_22827,N_23376);
nor U24112 (N_24112,N_23403,N_23483);
xnor U24113 (N_24113,N_23316,N_23949);
or U24114 (N_24114,N_23977,N_23442);
and U24115 (N_24115,N_23848,N_23734);
and U24116 (N_24116,N_23522,N_23292);
nor U24117 (N_24117,N_23773,N_23104);
nor U24118 (N_24118,N_23301,N_23878);
or U24119 (N_24119,N_23405,N_23092);
nand U24120 (N_24120,N_23983,N_23753);
and U24121 (N_24121,N_23518,N_23976);
or U24122 (N_24122,N_22956,N_23922);
nand U24123 (N_24123,N_23992,N_23234);
nand U24124 (N_24124,N_23731,N_22833);
and U24125 (N_24125,N_23547,N_23632);
xnor U24126 (N_24126,N_22949,N_23469);
and U24127 (N_24127,N_22830,N_22983);
nor U24128 (N_24128,N_23279,N_23365);
and U24129 (N_24129,N_22985,N_23546);
nor U24130 (N_24130,N_22835,N_23874);
and U24131 (N_24131,N_23445,N_23560);
nand U24132 (N_24132,N_23188,N_23212);
xnor U24133 (N_24133,N_23061,N_23891);
nand U24134 (N_24134,N_23723,N_22942);
nor U24135 (N_24135,N_23127,N_23629);
nand U24136 (N_24136,N_23933,N_23078);
nor U24137 (N_24137,N_23536,N_23304);
nor U24138 (N_24138,N_23062,N_23676);
and U24139 (N_24139,N_23989,N_23285);
and U24140 (N_24140,N_23196,N_23644);
nand U24141 (N_24141,N_23556,N_23490);
nor U24142 (N_24142,N_23860,N_23527);
or U24143 (N_24143,N_23950,N_23007);
and U24144 (N_24144,N_23801,N_23419);
nand U24145 (N_24145,N_23094,N_23966);
xnor U24146 (N_24146,N_22984,N_23786);
xor U24147 (N_24147,N_23250,N_23705);
and U24148 (N_24148,N_23122,N_23610);
nand U24149 (N_24149,N_23191,N_23909);
nand U24150 (N_24150,N_23863,N_23709);
or U24151 (N_24151,N_23215,N_23799);
and U24152 (N_24152,N_23450,N_23597);
and U24153 (N_24153,N_23776,N_23746);
and U24154 (N_24154,N_23955,N_23884);
xor U24155 (N_24155,N_23402,N_22874);
nor U24156 (N_24156,N_23011,N_23484);
or U24157 (N_24157,N_23532,N_23157);
and U24158 (N_24158,N_23350,N_23043);
nor U24159 (N_24159,N_23412,N_23700);
and U24160 (N_24160,N_23692,N_23608);
xor U24161 (N_24161,N_22811,N_23256);
xor U24162 (N_24162,N_23687,N_23908);
or U24163 (N_24163,N_22932,N_23941);
or U24164 (N_24164,N_23952,N_23868);
nand U24165 (N_24165,N_23004,N_22894);
xor U24166 (N_24166,N_23984,N_23843);
or U24167 (N_24167,N_23679,N_23675);
and U24168 (N_24168,N_23920,N_23036);
xnor U24169 (N_24169,N_23747,N_23824);
or U24170 (N_24170,N_22884,N_23184);
and U24171 (N_24171,N_23559,N_22895);
or U24172 (N_24172,N_23276,N_22878);
xnor U24173 (N_24173,N_23210,N_23990);
or U24174 (N_24174,N_22861,N_23363);
or U24175 (N_24175,N_23683,N_23354);
or U24176 (N_24176,N_22967,N_23349);
or U24177 (N_24177,N_23507,N_23648);
and U24178 (N_24178,N_23804,N_23454);
nand U24179 (N_24179,N_23051,N_22869);
and U24180 (N_24180,N_23703,N_23699);
xnor U24181 (N_24181,N_23334,N_23713);
xor U24182 (N_24182,N_23540,N_23805);
and U24183 (N_24183,N_23082,N_23842);
or U24184 (N_24184,N_23592,N_23951);
xor U24185 (N_24185,N_23488,N_23956);
or U24186 (N_24186,N_23180,N_22880);
or U24187 (N_24187,N_23481,N_23195);
and U24188 (N_24188,N_23331,N_22908);
and U24189 (N_24189,N_23470,N_23927);
or U24190 (N_24190,N_23525,N_23248);
xnor U24191 (N_24191,N_23310,N_23437);
nand U24192 (N_24192,N_23052,N_23257);
nand U24193 (N_24193,N_22804,N_22963);
nand U24194 (N_24194,N_23070,N_23772);
nor U24195 (N_24195,N_23817,N_23885);
or U24196 (N_24196,N_23561,N_22909);
and U24197 (N_24197,N_23549,N_22913);
nor U24198 (N_24198,N_22937,N_23591);
xor U24199 (N_24199,N_23642,N_23010);
xnor U24200 (N_24200,N_23777,N_23550);
or U24201 (N_24201,N_22948,N_23737);
and U24202 (N_24202,N_23996,N_22991);
nor U24203 (N_24203,N_22953,N_23580);
and U24204 (N_24204,N_23742,N_23586);
and U24205 (N_24205,N_23836,N_23613);
nor U24206 (N_24206,N_23281,N_23398);
or U24207 (N_24207,N_23182,N_23611);
or U24208 (N_24208,N_23137,N_22964);
or U24209 (N_24209,N_23837,N_22802);
xor U24210 (N_24210,N_23649,N_23037);
nand U24211 (N_24211,N_23109,N_23111);
nor U24212 (N_24212,N_23853,N_23539);
nand U24213 (N_24213,N_22851,N_23032);
xor U24214 (N_24214,N_23476,N_23243);
xor U24215 (N_24215,N_23551,N_23286);
and U24216 (N_24216,N_22999,N_23229);
or U24217 (N_24217,N_23465,N_22935);
or U24218 (N_24218,N_23523,N_23736);
and U24219 (N_24219,N_23046,N_23417);
and U24220 (N_24220,N_23216,N_23738);
and U24221 (N_24221,N_23410,N_23861);
or U24222 (N_24222,N_23566,N_23386);
nor U24223 (N_24223,N_23982,N_23171);
and U24224 (N_24224,N_23543,N_23967);
nor U24225 (N_24225,N_23666,N_23296);
nand U24226 (N_24226,N_22933,N_23168);
nand U24227 (N_24227,N_23987,N_23491);
or U24228 (N_24228,N_23424,N_22881);
and U24229 (N_24229,N_23134,N_23287);
and U24230 (N_24230,N_23428,N_23948);
nor U24231 (N_24231,N_23623,N_23093);
nor U24232 (N_24232,N_23579,N_23533);
nor U24233 (N_24233,N_23583,N_23049);
xnor U24234 (N_24234,N_22841,N_23392);
and U24235 (N_24235,N_23710,N_23076);
nand U24236 (N_24236,N_23769,N_22978);
xor U24237 (N_24237,N_23585,N_23151);
nand U24238 (N_24238,N_23981,N_23947);
xor U24239 (N_24239,N_23530,N_22899);
and U24240 (N_24240,N_22923,N_23872);
xnor U24241 (N_24241,N_23997,N_23840);
xnor U24242 (N_24242,N_23114,N_23858);
xnor U24243 (N_24243,N_23975,N_22897);
nor U24244 (N_24244,N_23911,N_23261);
xnor U24245 (N_24245,N_23016,N_23108);
nand U24246 (N_24246,N_23456,N_23496);
xor U24247 (N_24247,N_23345,N_23930);
and U24248 (N_24248,N_23673,N_23650);
xor U24249 (N_24249,N_23072,N_23055);
xor U24250 (N_24250,N_22961,N_23014);
nor U24251 (N_24251,N_23152,N_23520);
nand U24252 (N_24252,N_23869,N_23177);
xnor U24253 (N_24253,N_22800,N_23455);
or U24254 (N_24254,N_23293,N_23418);
xor U24255 (N_24255,N_23784,N_23409);
xor U24256 (N_24256,N_23504,N_23017);
nand U24257 (N_24257,N_23499,N_23719);
xnor U24258 (N_24258,N_23105,N_22813);
xnor U24259 (N_24259,N_23429,N_23367);
nor U24260 (N_24260,N_22994,N_23346);
and U24261 (N_24261,N_23745,N_23054);
and U24262 (N_24262,N_23433,N_23803);
or U24263 (N_24263,N_23935,N_23284);
nand U24264 (N_24264,N_23247,N_23223);
xor U24265 (N_24265,N_22939,N_23307);
or U24266 (N_24266,N_23926,N_23204);
and U24267 (N_24267,N_23235,N_23810);
nor U24268 (N_24268,N_23110,N_23646);
or U24269 (N_24269,N_23459,N_23206);
or U24270 (N_24270,N_23013,N_23633);
xor U24271 (N_24271,N_23555,N_22836);
nor U24272 (N_24272,N_23065,N_23047);
nor U24273 (N_24273,N_23780,N_23245);
nor U24274 (N_24274,N_23515,N_23026);
nand U24275 (N_24275,N_23406,N_23581);
or U24276 (N_24276,N_23654,N_23473);
nor U24277 (N_24277,N_23658,N_23069);
nor U24278 (N_24278,N_22928,N_23145);
xnor U24279 (N_24279,N_23467,N_23979);
xnor U24280 (N_24280,N_23132,N_23213);
or U24281 (N_24281,N_23308,N_23877);
nand U24282 (N_24282,N_23015,N_22824);
xor U24283 (N_24283,N_22826,N_23715);
and U24284 (N_24284,N_23552,N_22962);
xor U24285 (N_24285,N_23142,N_22837);
xnor U24286 (N_24286,N_23695,N_23083);
nor U24287 (N_24287,N_23426,N_23090);
nor U24288 (N_24288,N_23584,N_23370);
xor U24289 (N_24289,N_23749,N_23487);
nand U24290 (N_24290,N_23220,N_23466);
nor U24291 (N_24291,N_23529,N_23980);
xor U24292 (N_24292,N_22992,N_23618);
nand U24293 (N_24293,N_23609,N_23178);
nand U24294 (N_24294,N_23166,N_23464);
nand U24295 (N_24295,N_23449,N_23932);
and U24296 (N_24296,N_22867,N_23534);
and U24297 (N_24297,N_23880,N_23917);
or U24298 (N_24298,N_22807,N_23865);
nor U24299 (N_24299,N_23280,N_23077);
xnor U24300 (N_24300,N_22980,N_22976);
xor U24301 (N_24301,N_23486,N_23228);
and U24302 (N_24302,N_23009,N_23760);
xnor U24303 (N_24303,N_23901,N_23452);
or U24304 (N_24304,N_23988,N_23939);
nand U24305 (N_24305,N_23985,N_23866);
nand U24306 (N_24306,N_22925,N_23639);
and U24307 (N_24307,N_23567,N_22938);
nand U24308 (N_24308,N_22920,N_23670);
nand U24309 (N_24309,N_23750,N_23604);
and U24310 (N_24310,N_23681,N_23934);
or U24311 (N_24311,N_23271,N_23668);
or U24312 (N_24312,N_23944,N_23689);
xnor U24313 (N_24313,N_23115,N_23600);
xor U24314 (N_24314,N_23446,N_23400);
nor U24315 (N_24315,N_23826,N_23167);
and U24316 (N_24316,N_22940,N_23589);
and U24317 (N_24317,N_23545,N_22872);
and U24318 (N_24318,N_23775,N_22855);
xor U24319 (N_24319,N_23809,N_23506);
and U24320 (N_24320,N_23606,N_23970);
nand U24321 (N_24321,N_23720,N_23031);
and U24322 (N_24322,N_23348,N_22917);
xnor U24323 (N_24323,N_23873,N_22805);
nand U24324 (N_24324,N_22924,N_23557);
or U24325 (N_24325,N_22815,N_23471);
or U24326 (N_24326,N_23651,N_23329);
nor U24327 (N_24327,N_23251,N_23283);
and U24328 (N_24328,N_23088,N_23002);
and U24329 (N_24329,N_23388,N_22982);
and U24330 (N_24330,N_23126,N_22955);
nand U24331 (N_24331,N_23194,N_23057);
nor U24332 (N_24332,N_23730,N_23269);
or U24333 (N_24333,N_23290,N_23489);
and U24334 (N_24334,N_23806,N_23339);
xor U24335 (N_24335,N_23573,N_23211);
nand U24336 (N_24336,N_23106,N_23726);
and U24337 (N_24337,N_23198,N_23889);
nor U24338 (N_24338,N_23790,N_23154);
or U24339 (N_24339,N_23462,N_23170);
xor U24340 (N_24340,N_23686,N_23038);
or U24341 (N_24341,N_23075,N_22914);
nor U24342 (N_24342,N_23757,N_23441);
nand U24343 (N_24343,N_22905,N_23677);
and U24344 (N_24344,N_23931,N_23236);
nor U24345 (N_24345,N_23174,N_23133);
nand U24346 (N_24346,N_23572,N_22803);
and U24347 (N_24347,N_22818,N_22911);
and U24348 (N_24348,N_23892,N_23505);
and U24349 (N_24349,N_23306,N_23690);
xor U24350 (N_24350,N_22972,N_22844);
and U24351 (N_24351,N_22854,N_22842);
xor U24352 (N_24352,N_23834,N_23563);
nand U24353 (N_24353,N_23599,N_23811);
and U24354 (N_24354,N_23701,N_23787);
xor U24355 (N_24355,N_23850,N_23693);
and U24356 (N_24356,N_23558,N_23480);
or U24357 (N_24357,N_23356,N_23562);
or U24358 (N_24358,N_23986,N_23131);
xor U24359 (N_24359,N_23995,N_23640);
and U24360 (N_24360,N_23665,N_23159);
xor U24361 (N_24361,N_23888,N_23708);
or U24362 (N_24362,N_23954,N_23718);
and U24363 (N_24363,N_23253,N_23321);
nor U24364 (N_24364,N_22860,N_23461);
nand U24365 (N_24365,N_23871,N_23929);
nor U24366 (N_24366,N_23207,N_23886);
or U24367 (N_24367,N_23791,N_23625);
nor U24368 (N_24368,N_23798,N_23910);
and U24369 (N_24369,N_23045,N_22998);
and U24370 (N_24370,N_22981,N_23472);
nand U24371 (N_24371,N_22863,N_23959);
and U24372 (N_24372,N_22846,N_23612);
nand U24373 (N_24373,N_23265,N_23067);
and U24374 (N_24374,N_22821,N_23945);
nor U24375 (N_24375,N_22892,N_23991);
nor U24376 (N_24376,N_23816,N_23413);
nand U24377 (N_24377,N_22904,N_23839);
or U24378 (N_24378,N_23936,N_23390);
or U24379 (N_24379,N_23953,N_22809);
nor U24380 (N_24380,N_23022,N_23830);
nor U24381 (N_24381,N_23928,N_23593);
xor U24382 (N_24382,N_23727,N_23262);
nand U24383 (N_24383,N_23341,N_23135);
and U24384 (N_24384,N_23381,N_23254);
or U24385 (N_24385,N_23214,N_23000);
or U24386 (N_24386,N_23332,N_23343);
xor U24387 (N_24387,N_23199,N_23244);
nand U24388 (N_24388,N_23656,N_23620);
and U24389 (N_24389,N_22995,N_23759);
and U24390 (N_24390,N_23916,N_23193);
nor U24391 (N_24391,N_22910,N_23018);
and U24392 (N_24392,N_23973,N_23815);
nand U24393 (N_24393,N_23305,N_22943);
or U24394 (N_24394,N_23765,N_23782);
nor U24395 (N_24395,N_22888,N_23173);
and U24396 (N_24396,N_23333,N_22838);
or U24397 (N_24397,N_22936,N_23371);
nand U24398 (N_24398,N_23821,N_22968);
xnor U24399 (N_24399,N_23660,N_23685);
and U24400 (N_24400,N_23896,N_23309);
nor U24401 (N_24401,N_23965,N_22820);
or U24402 (N_24402,N_23238,N_23635);
and U24403 (N_24403,N_23521,N_22845);
nor U24404 (N_24404,N_23574,N_23379);
xnor U24405 (N_24405,N_23143,N_23494);
nand U24406 (N_24406,N_23792,N_23027);
or U24407 (N_24407,N_23438,N_23698);
xnor U24408 (N_24408,N_23636,N_23374);
nand U24409 (N_24409,N_23739,N_23421);
xor U24410 (N_24410,N_23577,N_23969);
and U24411 (N_24411,N_22882,N_23323);
or U24412 (N_24412,N_23358,N_23116);
xnor U24413 (N_24413,N_22832,N_23594);
nand U24414 (N_24414,N_23005,N_23224);
and U24415 (N_24415,N_22868,N_23508);
and U24416 (N_24416,N_23844,N_23189);
or U24417 (N_24417,N_23266,N_23766);
and U24418 (N_24418,N_22927,N_23957);
or U24419 (N_24419,N_23590,N_23270);
nand U24420 (N_24420,N_23602,N_23322);
and U24421 (N_24421,N_23282,N_23814);
xor U24422 (N_24422,N_23503,N_23854);
nor U24423 (N_24423,N_23347,N_23468);
or U24424 (N_24424,N_23793,N_23001);
or U24425 (N_24425,N_23401,N_23411);
or U24426 (N_24426,N_23813,N_23186);
nand U24427 (N_24427,N_22871,N_23783);
xor U24428 (N_24428,N_23829,N_23763);
xor U24429 (N_24429,N_23337,N_23230);
and U24430 (N_24430,N_23361,N_23086);
nor U24431 (N_24431,N_23607,N_22934);
xor U24432 (N_24432,N_23252,N_22823);
or U24433 (N_24433,N_23751,N_23394);
nor U24434 (N_24434,N_23373,N_23994);
and U24435 (N_24435,N_23420,N_23630);
nor U24436 (N_24436,N_22849,N_23838);
and U24437 (N_24437,N_22864,N_23407);
xor U24438 (N_24438,N_23395,N_23603);
and U24439 (N_24439,N_23203,N_23887);
or U24440 (N_24440,N_23377,N_23024);
nand U24441 (N_24441,N_23089,N_22945);
and U24442 (N_24442,N_22941,N_23702);
nor U24443 (N_24443,N_23112,N_23653);
nand U24444 (N_24444,N_23378,N_23818);
nand U24445 (N_24445,N_22926,N_23079);
or U24446 (N_24446,N_23063,N_23103);
xor U24447 (N_24447,N_23655,N_23318);
xor U24448 (N_24448,N_23042,N_23744);
xor U24449 (N_24449,N_23197,N_23925);
nor U24450 (N_24450,N_23435,N_23095);
and U24451 (N_24451,N_22891,N_23101);
xnor U24452 (N_24452,N_22959,N_23357);
nor U24453 (N_24453,N_23128,N_23458);
nor U24454 (N_24454,N_23919,N_23761);
and U24455 (N_24455,N_23657,N_23444);
xor U24456 (N_24456,N_23221,N_23768);
and U24457 (N_24457,N_23359,N_23774);
nand U24458 (N_24458,N_23588,N_22876);
xor U24459 (N_24459,N_23187,N_23427);
nand U24460 (N_24460,N_23688,N_22944);
and U24461 (N_24461,N_23124,N_23596);
nand U24462 (N_24462,N_23796,N_23680);
or U24463 (N_24463,N_23587,N_22890);
xor U24464 (N_24464,N_22947,N_23457);
nand U24465 (N_24465,N_23432,N_23139);
xnor U24466 (N_24466,N_23795,N_23231);
or U24467 (N_24467,N_23414,N_23770);
xor U24468 (N_24468,N_23164,N_22996);
or U24469 (N_24469,N_23396,N_23833);
or U24470 (N_24470,N_23921,N_23914);
and U24471 (N_24471,N_23387,N_23807);
nand U24472 (N_24472,N_22817,N_23906);
and U24473 (N_24473,N_23516,N_23200);
and U24474 (N_24474,N_23179,N_23222);
xor U24475 (N_24475,N_22840,N_23762);
xnor U24476 (N_24476,N_23882,N_23225);
nor U24477 (N_24477,N_22974,N_23436);
nor U24478 (N_24478,N_22915,N_23637);
and U24479 (N_24479,N_23902,N_22850);
nand U24480 (N_24480,N_22986,N_23039);
or U24481 (N_24481,N_23511,N_23288);
or U24482 (N_24482,N_22946,N_23978);
or U24483 (N_24483,N_23241,N_23267);
and U24484 (N_24484,N_23289,N_22848);
or U24485 (N_24485,N_23711,N_23741);
nand U24486 (N_24486,N_23748,N_23422);
nor U24487 (N_24487,N_23475,N_23595);
xor U24488 (N_24488,N_23325,N_23509);
nand U24489 (N_24489,N_23113,N_23661);
nor U24490 (N_24490,N_23812,N_23846);
nor U24491 (N_24491,N_23125,N_23542);
or U24492 (N_24492,N_23327,N_23302);
or U24493 (N_24493,N_23268,N_22877);
and U24494 (N_24494,N_23217,N_23808);
xor U24495 (N_24495,N_23163,N_23156);
nand U24496 (N_24496,N_23964,N_23528);
nor U24497 (N_24497,N_23393,N_23669);
and U24498 (N_24498,N_23399,N_23237);
nand U24499 (N_24499,N_22819,N_23616);
and U24500 (N_24500,N_23369,N_23391);
xor U24501 (N_24501,N_22900,N_23160);
or U24502 (N_24502,N_23123,N_23671);
and U24503 (N_24503,N_23493,N_23758);
nor U24504 (N_24504,N_23278,N_23820);
xor U24505 (N_24505,N_22893,N_23999);
or U24506 (N_24506,N_22843,N_23845);
nor U24507 (N_24507,N_22952,N_23832);
and U24508 (N_24508,N_23058,N_22929);
xnor U24509 (N_24509,N_23879,N_23303);
nand U24510 (N_24510,N_23883,N_23071);
xor U24511 (N_24511,N_22916,N_23497);
nand U24512 (N_24512,N_23096,N_22993);
or U24513 (N_24513,N_22931,N_23232);
nand U24514 (N_24514,N_23153,N_23961);
nor U24515 (N_24515,N_23924,N_23482);
xor U24516 (N_24516,N_23340,N_23915);
xor U24517 (N_24517,N_23538,N_22865);
or U24518 (N_24518,N_23571,N_23524);
xor U24519 (N_24519,N_23789,N_23495);
xor U24520 (N_24520,N_23626,N_23208);
or U24521 (N_24521,N_23059,N_23663);
or U24522 (N_24522,N_23119,N_23501);
xor U24523 (N_24523,N_23893,N_23242);
and U24524 (N_24524,N_23696,N_22997);
and U24525 (N_24525,N_23044,N_23205);
nand U24526 (N_24526,N_23227,N_22810);
and U24527 (N_24527,N_22979,N_23299);
nand U24528 (N_24528,N_23181,N_22887);
nor U24529 (N_24529,N_23852,N_23645);
or U24530 (N_24530,N_22885,N_23998);
xor U24531 (N_24531,N_23662,N_23894);
xor U24532 (N_24532,N_23118,N_23485);
nand U24533 (N_24533,N_22829,N_23034);
nand U24534 (N_24534,N_23311,N_23192);
and U24535 (N_24535,N_23073,N_23800);
or U24536 (N_24536,N_23856,N_22901);
nand U24537 (N_24537,N_23743,N_22801);
or U24538 (N_24538,N_23943,N_23564);
nor U24539 (N_24539,N_23291,N_23272);
or U24540 (N_24540,N_23098,N_23619);
xor U24541 (N_24541,N_23576,N_22922);
xnor U24542 (N_24542,N_23448,N_23993);
nand U24543 (N_24543,N_23706,N_23440);
nand U24544 (N_24544,N_23897,N_23659);
and U24545 (N_24545,N_23535,N_23694);
nand U24546 (N_24546,N_23175,N_23275);
xnor U24547 (N_24547,N_23183,N_23158);
xnor U24548 (N_24548,N_22883,N_23120);
nor U24549 (N_24549,N_23081,N_23779);
or U24550 (N_24550,N_23674,N_23130);
xnor U24551 (N_24551,N_23249,N_23443);
and U24552 (N_24552,N_23404,N_22853);
xnor U24553 (N_24553,N_23851,N_23425);
nand U24554 (N_24554,N_22834,N_23628);
nand U24555 (N_24555,N_23570,N_23544);
or U24556 (N_24556,N_22969,N_23050);
or U24557 (N_24557,N_22988,N_23100);
xnor U24558 (N_24558,N_23864,N_22808);
nor U24559 (N_24559,N_23169,N_23912);
nor U24560 (N_24560,N_23895,N_22814);
or U24561 (N_24561,N_23149,N_23740);
or U24562 (N_24562,N_22906,N_23752);
nand U24563 (N_24563,N_23502,N_22870);
or U24564 (N_24564,N_23831,N_23162);
nor U24565 (N_24565,N_23621,N_23962);
and U24566 (N_24566,N_23802,N_23717);
xor U24567 (N_24567,N_23569,N_23510);
nor U24568 (N_24568,N_23147,N_23541);
or U24569 (N_24569,N_23617,N_22812);
or U24570 (N_24570,N_23439,N_23209);
xor U24571 (N_24571,N_23918,N_23397);
or U24572 (N_24572,N_23233,N_23652);
nor U24573 (N_24573,N_23862,N_23575);
nor U24574 (N_24574,N_23389,N_23368);
nor U24575 (N_24575,N_23006,N_22896);
nor U24576 (N_24576,N_23684,N_23721);
and U24577 (N_24577,N_23771,N_23326);
nand U24578 (N_24578,N_23298,N_23825);
xnor U24579 (N_24579,N_23667,N_23453);
or U24580 (N_24580,N_23847,N_22971);
or U24581 (N_24581,N_23150,N_23767);
and U24582 (N_24582,N_22857,N_23519);
xor U24583 (N_24583,N_23682,N_23068);
xor U24584 (N_24584,N_23890,N_23631);
nor U24585 (N_24585,N_23056,N_22975);
and U24586 (N_24586,N_23725,N_22989);
or U24587 (N_24587,N_23146,N_23968);
xnor U24588 (N_24588,N_22852,N_23355);
and U24589 (N_24589,N_23423,N_22954);
nand U24590 (N_24590,N_23553,N_23121);
nor U24591 (N_24591,N_23712,N_23239);
nor U24592 (N_24592,N_22828,N_23512);
xor U24593 (N_24593,N_22950,N_22921);
nor U24594 (N_24594,N_23601,N_22965);
nand U24595 (N_24595,N_23477,N_23898);
nand U24596 (N_24596,N_23940,N_23876);
nor U24597 (N_24597,N_23064,N_23176);
and U24598 (N_24598,N_23041,N_22912);
xnor U24599 (N_24599,N_22970,N_23634);
nor U24600 (N_24600,N_23984,N_23336);
nor U24601 (N_24601,N_23550,N_23101);
nor U24602 (N_24602,N_22904,N_23632);
or U24603 (N_24603,N_23852,N_23819);
and U24604 (N_24604,N_22836,N_23365);
and U24605 (N_24605,N_22837,N_23390);
and U24606 (N_24606,N_23637,N_23217);
nor U24607 (N_24607,N_23539,N_23716);
xnor U24608 (N_24608,N_23406,N_23931);
nor U24609 (N_24609,N_23407,N_22935);
nor U24610 (N_24610,N_23916,N_23949);
nand U24611 (N_24611,N_23945,N_23203);
nor U24612 (N_24612,N_23255,N_23942);
xnor U24613 (N_24613,N_23948,N_23366);
nor U24614 (N_24614,N_23711,N_23733);
nor U24615 (N_24615,N_23264,N_23714);
xor U24616 (N_24616,N_23347,N_22867);
nand U24617 (N_24617,N_23973,N_23861);
nor U24618 (N_24618,N_23128,N_23881);
nor U24619 (N_24619,N_23610,N_23855);
and U24620 (N_24620,N_23733,N_23822);
nor U24621 (N_24621,N_22937,N_23285);
and U24622 (N_24622,N_23347,N_23757);
nand U24623 (N_24623,N_23596,N_22932);
nand U24624 (N_24624,N_23837,N_23303);
nor U24625 (N_24625,N_23168,N_23585);
and U24626 (N_24626,N_23298,N_22971);
xor U24627 (N_24627,N_23046,N_23544);
nor U24628 (N_24628,N_23756,N_23313);
nand U24629 (N_24629,N_23064,N_23838);
nor U24630 (N_24630,N_23705,N_23939);
or U24631 (N_24631,N_23725,N_23593);
and U24632 (N_24632,N_23383,N_23007);
nor U24633 (N_24633,N_23824,N_23426);
nor U24634 (N_24634,N_23108,N_23804);
or U24635 (N_24635,N_23055,N_23672);
nor U24636 (N_24636,N_23709,N_23681);
or U24637 (N_24637,N_22809,N_23053);
or U24638 (N_24638,N_23697,N_23417);
or U24639 (N_24639,N_23456,N_23492);
nand U24640 (N_24640,N_23991,N_23498);
or U24641 (N_24641,N_23376,N_23741);
and U24642 (N_24642,N_23698,N_23517);
and U24643 (N_24643,N_23805,N_23693);
nor U24644 (N_24644,N_23031,N_22910);
and U24645 (N_24645,N_22925,N_23072);
nand U24646 (N_24646,N_22954,N_23805);
or U24647 (N_24647,N_23057,N_23937);
nor U24648 (N_24648,N_23446,N_23125);
nor U24649 (N_24649,N_23743,N_23946);
xor U24650 (N_24650,N_23723,N_23998);
nor U24651 (N_24651,N_23196,N_23417);
or U24652 (N_24652,N_23292,N_23639);
nor U24653 (N_24653,N_23603,N_23593);
nand U24654 (N_24654,N_23481,N_22993);
nor U24655 (N_24655,N_23332,N_23209);
and U24656 (N_24656,N_23172,N_23895);
xnor U24657 (N_24657,N_23759,N_23708);
nor U24658 (N_24658,N_23613,N_23789);
or U24659 (N_24659,N_22820,N_23235);
xor U24660 (N_24660,N_23240,N_23642);
or U24661 (N_24661,N_23237,N_23061);
nor U24662 (N_24662,N_22918,N_23843);
nor U24663 (N_24663,N_23855,N_23598);
nand U24664 (N_24664,N_23415,N_23439);
and U24665 (N_24665,N_23015,N_23779);
or U24666 (N_24666,N_22801,N_23018);
or U24667 (N_24667,N_23922,N_23099);
xor U24668 (N_24668,N_23910,N_23338);
xor U24669 (N_24669,N_23590,N_23559);
xor U24670 (N_24670,N_23553,N_23619);
nor U24671 (N_24671,N_23009,N_23648);
or U24672 (N_24672,N_23700,N_23635);
xor U24673 (N_24673,N_23848,N_23501);
nor U24674 (N_24674,N_23722,N_23113);
nand U24675 (N_24675,N_23915,N_23884);
xnor U24676 (N_24676,N_23175,N_23789);
xnor U24677 (N_24677,N_23802,N_23118);
and U24678 (N_24678,N_22984,N_23591);
or U24679 (N_24679,N_23480,N_23929);
and U24680 (N_24680,N_23306,N_23006);
xnor U24681 (N_24681,N_23051,N_23661);
nor U24682 (N_24682,N_22935,N_23614);
or U24683 (N_24683,N_23120,N_23651);
or U24684 (N_24684,N_22985,N_23235);
nand U24685 (N_24685,N_23936,N_22836);
xor U24686 (N_24686,N_22841,N_23293);
or U24687 (N_24687,N_23539,N_23002);
and U24688 (N_24688,N_23210,N_23506);
nand U24689 (N_24689,N_23610,N_23595);
or U24690 (N_24690,N_23149,N_23079);
nand U24691 (N_24691,N_23467,N_22896);
nand U24692 (N_24692,N_23205,N_23571);
nand U24693 (N_24693,N_23985,N_22831);
xor U24694 (N_24694,N_23518,N_23196);
or U24695 (N_24695,N_23540,N_23282);
and U24696 (N_24696,N_23120,N_22846);
nor U24697 (N_24697,N_23729,N_22934);
nor U24698 (N_24698,N_23223,N_23036);
xor U24699 (N_24699,N_23896,N_22985);
nor U24700 (N_24700,N_23775,N_22880);
xor U24701 (N_24701,N_23463,N_23489);
nand U24702 (N_24702,N_23502,N_23048);
nor U24703 (N_24703,N_23071,N_23236);
nor U24704 (N_24704,N_23530,N_23293);
xnor U24705 (N_24705,N_23551,N_22994);
or U24706 (N_24706,N_23018,N_23925);
and U24707 (N_24707,N_23894,N_23352);
xnor U24708 (N_24708,N_22861,N_23480);
or U24709 (N_24709,N_23323,N_22948);
xnor U24710 (N_24710,N_23211,N_22942);
and U24711 (N_24711,N_23392,N_23301);
and U24712 (N_24712,N_22985,N_22809);
xnor U24713 (N_24713,N_23534,N_22862);
nand U24714 (N_24714,N_23202,N_23976);
xor U24715 (N_24715,N_23941,N_22877);
xor U24716 (N_24716,N_23547,N_22818);
xnor U24717 (N_24717,N_23654,N_23147);
nor U24718 (N_24718,N_23414,N_22880);
and U24719 (N_24719,N_23608,N_23732);
or U24720 (N_24720,N_23616,N_22848);
nor U24721 (N_24721,N_23452,N_22835);
or U24722 (N_24722,N_23426,N_23920);
nand U24723 (N_24723,N_23039,N_23493);
or U24724 (N_24724,N_22882,N_23685);
xor U24725 (N_24725,N_23257,N_23069);
nor U24726 (N_24726,N_23700,N_23146);
nor U24727 (N_24727,N_23938,N_23325);
and U24728 (N_24728,N_23967,N_22922);
xor U24729 (N_24729,N_22964,N_23461);
or U24730 (N_24730,N_23592,N_23010);
nor U24731 (N_24731,N_23212,N_23881);
and U24732 (N_24732,N_23876,N_23292);
nand U24733 (N_24733,N_23143,N_23665);
xnor U24734 (N_24734,N_23836,N_23540);
nor U24735 (N_24735,N_22980,N_22887);
nor U24736 (N_24736,N_23771,N_23590);
nand U24737 (N_24737,N_23673,N_23432);
nor U24738 (N_24738,N_23237,N_23455);
xor U24739 (N_24739,N_23238,N_23926);
nand U24740 (N_24740,N_23914,N_23610);
nand U24741 (N_24741,N_23881,N_23542);
xnor U24742 (N_24742,N_22805,N_22904);
or U24743 (N_24743,N_23809,N_23280);
nor U24744 (N_24744,N_23878,N_22982);
xor U24745 (N_24745,N_23514,N_23641);
nor U24746 (N_24746,N_23009,N_23945);
nand U24747 (N_24747,N_23173,N_23072);
nand U24748 (N_24748,N_23057,N_22928);
nor U24749 (N_24749,N_23782,N_22880);
and U24750 (N_24750,N_23201,N_23158);
and U24751 (N_24751,N_23925,N_22967);
or U24752 (N_24752,N_23246,N_22820);
nor U24753 (N_24753,N_23804,N_23046);
and U24754 (N_24754,N_23356,N_23993);
and U24755 (N_24755,N_22930,N_23015);
nand U24756 (N_24756,N_23069,N_23256);
and U24757 (N_24757,N_23226,N_22852);
xnor U24758 (N_24758,N_23783,N_22984);
xnor U24759 (N_24759,N_23191,N_23336);
nor U24760 (N_24760,N_23851,N_23628);
and U24761 (N_24761,N_22846,N_23870);
xnor U24762 (N_24762,N_22919,N_23689);
xor U24763 (N_24763,N_23246,N_23452);
nor U24764 (N_24764,N_23099,N_23269);
and U24765 (N_24765,N_23701,N_23752);
nor U24766 (N_24766,N_22887,N_23465);
or U24767 (N_24767,N_23683,N_23613);
or U24768 (N_24768,N_23364,N_23786);
xnor U24769 (N_24769,N_23753,N_23034);
and U24770 (N_24770,N_23689,N_23041);
or U24771 (N_24771,N_22936,N_23105);
or U24772 (N_24772,N_23973,N_23995);
xor U24773 (N_24773,N_22899,N_23920);
nand U24774 (N_24774,N_23091,N_23255);
and U24775 (N_24775,N_23606,N_23307);
nand U24776 (N_24776,N_23820,N_23769);
and U24777 (N_24777,N_23473,N_23214);
nand U24778 (N_24778,N_23187,N_23938);
or U24779 (N_24779,N_23260,N_23611);
or U24780 (N_24780,N_23263,N_23019);
nor U24781 (N_24781,N_22852,N_23834);
nor U24782 (N_24782,N_23490,N_23534);
or U24783 (N_24783,N_23419,N_23291);
and U24784 (N_24784,N_23564,N_22895);
xor U24785 (N_24785,N_23973,N_23498);
nor U24786 (N_24786,N_23788,N_23103);
nand U24787 (N_24787,N_23633,N_23486);
nand U24788 (N_24788,N_23412,N_23265);
xnor U24789 (N_24789,N_23830,N_23630);
and U24790 (N_24790,N_23212,N_23607);
or U24791 (N_24791,N_23017,N_23544);
nand U24792 (N_24792,N_23512,N_23649);
xor U24793 (N_24793,N_22920,N_23484);
nor U24794 (N_24794,N_23509,N_23218);
or U24795 (N_24795,N_23253,N_22825);
and U24796 (N_24796,N_23630,N_23590);
nand U24797 (N_24797,N_22878,N_23698);
xnor U24798 (N_24798,N_23794,N_23507);
nand U24799 (N_24799,N_23461,N_23226);
or U24800 (N_24800,N_23516,N_23839);
or U24801 (N_24801,N_23781,N_23197);
nand U24802 (N_24802,N_23816,N_22873);
xor U24803 (N_24803,N_23956,N_23540);
and U24804 (N_24804,N_23600,N_23076);
and U24805 (N_24805,N_23753,N_23896);
nand U24806 (N_24806,N_23743,N_22847);
or U24807 (N_24807,N_23760,N_22849);
and U24808 (N_24808,N_23654,N_23393);
or U24809 (N_24809,N_23180,N_22857);
and U24810 (N_24810,N_23665,N_23773);
or U24811 (N_24811,N_23570,N_23670);
and U24812 (N_24812,N_23266,N_23361);
or U24813 (N_24813,N_22884,N_23227);
or U24814 (N_24814,N_23768,N_23160);
xor U24815 (N_24815,N_23815,N_23534);
and U24816 (N_24816,N_23046,N_23930);
xor U24817 (N_24817,N_23687,N_23727);
nor U24818 (N_24818,N_23481,N_23759);
xor U24819 (N_24819,N_23453,N_23259);
xnor U24820 (N_24820,N_23630,N_23734);
and U24821 (N_24821,N_23142,N_23938);
nand U24822 (N_24822,N_23172,N_22926);
or U24823 (N_24823,N_23433,N_23720);
or U24824 (N_24824,N_23069,N_22819);
nor U24825 (N_24825,N_23436,N_23257);
and U24826 (N_24826,N_23973,N_23082);
xor U24827 (N_24827,N_23377,N_23774);
nor U24828 (N_24828,N_22904,N_23745);
and U24829 (N_24829,N_23464,N_23365);
nor U24830 (N_24830,N_23810,N_23448);
nand U24831 (N_24831,N_23875,N_23217);
nand U24832 (N_24832,N_23904,N_23308);
and U24833 (N_24833,N_23913,N_23469);
nor U24834 (N_24834,N_23764,N_23757);
or U24835 (N_24835,N_23353,N_22812);
or U24836 (N_24836,N_23148,N_23776);
or U24837 (N_24837,N_23437,N_23218);
nand U24838 (N_24838,N_22923,N_23720);
nor U24839 (N_24839,N_23060,N_23916);
nor U24840 (N_24840,N_23168,N_23813);
or U24841 (N_24841,N_22842,N_23224);
or U24842 (N_24842,N_22805,N_23038);
or U24843 (N_24843,N_23912,N_23407);
or U24844 (N_24844,N_23729,N_22936);
xor U24845 (N_24845,N_23572,N_23263);
and U24846 (N_24846,N_23580,N_23503);
xor U24847 (N_24847,N_23419,N_23175);
nor U24848 (N_24848,N_22917,N_23144);
nand U24849 (N_24849,N_23307,N_23616);
nand U24850 (N_24850,N_23652,N_23595);
nand U24851 (N_24851,N_23660,N_23216);
nor U24852 (N_24852,N_23096,N_23437);
and U24853 (N_24853,N_22940,N_22985);
or U24854 (N_24854,N_23228,N_23799);
nor U24855 (N_24855,N_23720,N_22818);
nand U24856 (N_24856,N_22871,N_23400);
nand U24857 (N_24857,N_23806,N_23859);
xor U24858 (N_24858,N_22846,N_23027);
nor U24859 (N_24859,N_23565,N_23197);
and U24860 (N_24860,N_23149,N_23861);
and U24861 (N_24861,N_23555,N_23413);
and U24862 (N_24862,N_23943,N_23742);
nand U24863 (N_24863,N_23961,N_23122);
xnor U24864 (N_24864,N_22906,N_23002);
nand U24865 (N_24865,N_23036,N_23200);
nor U24866 (N_24866,N_23441,N_23112);
nor U24867 (N_24867,N_22924,N_23772);
xnor U24868 (N_24868,N_23392,N_23828);
nand U24869 (N_24869,N_23700,N_23955);
and U24870 (N_24870,N_23974,N_23222);
nand U24871 (N_24871,N_23424,N_23477);
nand U24872 (N_24872,N_23217,N_23494);
nor U24873 (N_24873,N_23029,N_23769);
or U24874 (N_24874,N_23407,N_23478);
xor U24875 (N_24875,N_23877,N_23260);
and U24876 (N_24876,N_23717,N_23891);
and U24877 (N_24877,N_23823,N_23214);
and U24878 (N_24878,N_23905,N_23927);
nor U24879 (N_24879,N_23391,N_23725);
or U24880 (N_24880,N_23736,N_22849);
or U24881 (N_24881,N_23284,N_23461);
or U24882 (N_24882,N_22810,N_23113);
nand U24883 (N_24883,N_23520,N_23499);
xnor U24884 (N_24884,N_22934,N_23703);
and U24885 (N_24885,N_22828,N_23464);
or U24886 (N_24886,N_22898,N_23181);
nand U24887 (N_24887,N_23716,N_23958);
nand U24888 (N_24888,N_23059,N_22875);
or U24889 (N_24889,N_23936,N_22888);
nand U24890 (N_24890,N_23542,N_23717);
nor U24891 (N_24891,N_22887,N_23926);
xnor U24892 (N_24892,N_23564,N_22926);
and U24893 (N_24893,N_23165,N_23340);
nor U24894 (N_24894,N_23764,N_23218);
nor U24895 (N_24895,N_23096,N_23872);
nand U24896 (N_24896,N_23469,N_23208);
xnor U24897 (N_24897,N_23167,N_22828);
xor U24898 (N_24898,N_23849,N_23577);
and U24899 (N_24899,N_23721,N_23632);
and U24900 (N_24900,N_23090,N_23018);
or U24901 (N_24901,N_22932,N_23227);
nand U24902 (N_24902,N_23242,N_23385);
nor U24903 (N_24903,N_23242,N_23152);
or U24904 (N_24904,N_23904,N_23681);
nor U24905 (N_24905,N_23956,N_22873);
xor U24906 (N_24906,N_23005,N_23556);
nor U24907 (N_24907,N_23358,N_22855);
nor U24908 (N_24908,N_23239,N_22983);
or U24909 (N_24909,N_23992,N_23720);
nand U24910 (N_24910,N_23920,N_22891);
or U24911 (N_24911,N_22947,N_23796);
nor U24912 (N_24912,N_23219,N_23122);
xnor U24913 (N_24913,N_22997,N_23663);
xnor U24914 (N_24914,N_22957,N_23693);
nand U24915 (N_24915,N_23129,N_23606);
nor U24916 (N_24916,N_23048,N_23631);
nand U24917 (N_24917,N_23946,N_23202);
nand U24918 (N_24918,N_23644,N_23876);
xor U24919 (N_24919,N_23312,N_22924);
and U24920 (N_24920,N_23494,N_23726);
nor U24921 (N_24921,N_22857,N_23596);
nand U24922 (N_24922,N_23428,N_23310);
and U24923 (N_24923,N_23583,N_23188);
or U24924 (N_24924,N_23378,N_23713);
nor U24925 (N_24925,N_22902,N_23410);
xor U24926 (N_24926,N_23965,N_23121);
and U24927 (N_24927,N_23721,N_23705);
nand U24928 (N_24928,N_23672,N_22879);
nor U24929 (N_24929,N_23866,N_23169);
xnor U24930 (N_24930,N_22929,N_23699);
nor U24931 (N_24931,N_23479,N_23978);
nor U24932 (N_24932,N_22939,N_23085);
nand U24933 (N_24933,N_23539,N_23502);
and U24934 (N_24934,N_23784,N_23360);
and U24935 (N_24935,N_23537,N_22802);
and U24936 (N_24936,N_22960,N_23238);
xor U24937 (N_24937,N_23914,N_23297);
or U24938 (N_24938,N_23607,N_23165);
or U24939 (N_24939,N_23771,N_23164);
xor U24940 (N_24940,N_23703,N_23914);
nand U24941 (N_24941,N_23259,N_23998);
or U24942 (N_24942,N_23863,N_23198);
and U24943 (N_24943,N_23625,N_22949);
xor U24944 (N_24944,N_23284,N_23791);
xnor U24945 (N_24945,N_23832,N_22873);
nand U24946 (N_24946,N_23015,N_23244);
or U24947 (N_24947,N_23031,N_22892);
or U24948 (N_24948,N_23267,N_22996);
and U24949 (N_24949,N_23413,N_22908);
or U24950 (N_24950,N_22874,N_23882);
or U24951 (N_24951,N_22840,N_23733);
and U24952 (N_24952,N_23122,N_22809);
and U24953 (N_24953,N_23936,N_23255);
and U24954 (N_24954,N_23942,N_23060);
and U24955 (N_24955,N_23127,N_23839);
nand U24956 (N_24956,N_23910,N_23189);
nor U24957 (N_24957,N_23263,N_23523);
or U24958 (N_24958,N_23528,N_22824);
and U24959 (N_24959,N_23558,N_23867);
nor U24960 (N_24960,N_23230,N_22996);
or U24961 (N_24961,N_23104,N_23053);
xnor U24962 (N_24962,N_22840,N_23032);
nor U24963 (N_24963,N_23427,N_23284);
and U24964 (N_24964,N_23064,N_23698);
nand U24965 (N_24965,N_23855,N_22948);
and U24966 (N_24966,N_23205,N_23801);
nor U24967 (N_24967,N_23529,N_23091);
nand U24968 (N_24968,N_23639,N_23678);
and U24969 (N_24969,N_23259,N_23604);
or U24970 (N_24970,N_23665,N_23519);
nand U24971 (N_24971,N_22942,N_23378);
nor U24972 (N_24972,N_23794,N_23550);
xnor U24973 (N_24973,N_23203,N_23848);
and U24974 (N_24974,N_23184,N_23329);
or U24975 (N_24975,N_22822,N_23547);
xor U24976 (N_24976,N_22890,N_23576);
or U24977 (N_24977,N_23718,N_23767);
nor U24978 (N_24978,N_23547,N_23996);
and U24979 (N_24979,N_23527,N_23192);
or U24980 (N_24980,N_23710,N_23849);
or U24981 (N_24981,N_23760,N_23845);
and U24982 (N_24982,N_23191,N_22923);
or U24983 (N_24983,N_23121,N_22980);
nand U24984 (N_24984,N_23165,N_23760);
or U24985 (N_24985,N_23560,N_22937);
nor U24986 (N_24986,N_23678,N_22897);
and U24987 (N_24987,N_22853,N_23556);
xor U24988 (N_24988,N_23188,N_23954);
nor U24989 (N_24989,N_23136,N_23984);
and U24990 (N_24990,N_23318,N_22949);
and U24991 (N_24991,N_23736,N_23963);
nand U24992 (N_24992,N_23468,N_23456);
xnor U24993 (N_24993,N_23157,N_23009);
nand U24994 (N_24994,N_23210,N_23400);
xnor U24995 (N_24995,N_23492,N_23684);
nor U24996 (N_24996,N_22817,N_23498);
xnor U24997 (N_24997,N_23093,N_23308);
xnor U24998 (N_24998,N_23964,N_23339);
nand U24999 (N_24999,N_23291,N_23472);
nor U25000 (N_25000,N_22999,N_23675);
or U25001 (N_25001,N_23198,N_23989);
nand U25002 (N_25002,N_23372,N_23366);
nand U25003 (N_25003,N_23155,N_23812);
nor U25004 (N_25004,N_23339,N_23588);
and U25005 (N_25005,N_22870,N_22859);
or U25006 (N_25006,N_23140,N_23082);
nor U25007 (N_25007,N_23679,N_23708);
or U25008 (N_25008,N_22818,N_23270);
nand U25009 (N_25009,N_23913,N_23962);
nor U25010 (N_25010,N_23999,N_23598);
nor U25011 (N_25011,N_23261,N_23691);
nor U25012 (N_25012,N_23774,N_23493);
and U25013 (N_25013,N_23581,N_23849);
nor U25014 (N_25014,N_23724,N_22965);
or U25015 (N_25015,N_23860,N_23471);
nand U25016 (N_25016,N_23290,N_23458);
nor U25017 (N_25017,N_22892,N_23640);
or U25018 (N_25018,N_22884,N_23240);
or U25019 (N_25019,N_23890,N_23406);
xor U25020 (N_25020,N_23408,N_23037);
xnor U25021 (N_25021,N_23438,N_23876);
and U25022 (N_25022,N_23198,N_23515);
or U25023 (N_25023,N_23095,N_23622);
nor U25024 (N_25024,N_23252,N_23158);
nand U25025 (N_25025,N_23192,N_23418);
and U25026 (N_25026,N_23819,N_22918);
and U25027 (N_25027,N_23403,N_23808);
nand U25028 (N_25028,N_23722,N_22839);
and U25029 (N_25029,N_22861,N_23618);
xor U25030 (N_25030,N_23353,N_23008);
xnor U25031 (N_25031,N_23501,N_23866);
nor U25032 (N_25032,N_23604,N_23025);
nand U25033 (N_25033,N_23144,N_23947);
and U25034 (N_25034,N_23455,N_23073);
nor U25035 (N_25035,N_22910,N_23302);
and U25036 (N_25036,N_23072,N_23715);
nor U25037 (N_25037,N_23503,N_23924);
or U25038 (N_25038,N_23347,N_23512);
or U25039 (N_25039,N_23126,N_23511);
or U25040 (N_25040,N_23720,N_23071);
or U25041 (N_25041,N_22809,N_23506);
and U25042 (N_25042,N_23761,N_23943);
nor U25043 (N_25043,N_23213,N_22987);
or U25044 (N_25044,N_23216,N_23657);
nor U25045 (N_25045,N_23096,N_23129);
xor U25046 (N_25046,N_23976,N_23367);
nand U25047 (N_25047,N_23982,N_22830);
or U25048 (N_25048,N_23890,N_23902);
nor U25049 (N_25049,N_23282,N_23146);
and U25050 (N_25050,N_23972,N_23834);
or U25051 (N_25051,N_23210,N_23654);
nand U25052 (N_25052,N_23990,N_23413);
nor U25053 (N_25053,N_23727,N_23240);
or U25054 (N_25054,N_22967,N_23509);
xnor U25055 (N_25055,N_23292,N_22802);
or U25056 (N_25056,N_22970,N_23268);
nand U25057 (N_25057,N_23399,N_23861);
nand U25058 (N_25058,N_23990,N_23019);
or U25059 (N_25059,N_23037,N_23959);
nand U25060 (N_25060,N_23538,N_22910);
nand U25061 (N_25061,N_22889,N_23302);
and U25062 (N_25062,N_23353,N_23568);
xnor U25063 (N_25063,N_23655,N_22883);
nand U25064 (N_25064,N_23399,N_23964);
and U25065 (N_25065,N_23377,N_23347);
nor U25066 (N_25066,N_23221,N_23737);
and U25067 (N_25067,N_23864,N_22903);
and U25068 (N_25068,N_23877,N_23896);
nor U25069 (N_25069,N_23288,N_23562);
xnor U25070 (N_25070,N_23447,N_23574);
nand U25071 (N_25071,N_23262,N_23349);
nand U25072 (N_25072,N_23904,N_23609);
nor U25073 (N_25073,N_23471,N_23535);
or U25074 (N_25074,N_23954,N_23370);
and U25075 (N_25075,N_23726,N_23721);
or U25076 (N_25076,N_23959,N_23026);
xor U25077 (N_25077,N_23624,N_22920);
nand U25078 (N_25078,N_23977,N_22952);
xor U25079 (N_25079,N_23336,N_22920);
or U25080 (N_25080,N_23002,N_22907);
nand U25081 (N_25081,N_23518,N_23266);
or U25082 (N_25082,N_23804,N_22941);
and U25083 (N_25083,N_23908,N_23614);
nand U25084 (N_25084,N_22990,N_22902);
nand U25085 (N_25085,N_23753,N_23989);
xnor U25086 (N_25086,N_22886,N_23799);
or U25087 (N_25087,N_23030,N_23369);
and U25088 (N_25088,N_23507,N_23468);
nand U25089 (N_25089,N_23812,N_23345);
nand U25090 (N_25090,N_23635,N_22972);
nor U25091 (N_25091,N_23387,N_23077);
and U25092 (N_25092,N_23145,N_23828);
and U25093 (N_25093,N_23499,N_23456);
xnor U25094 (N_25094,N_23776,N_23916);
and U25095 (N_25095,N_22901,N_23600);
or U25096 (N_25096,N_23981,N_23297);
nor U25097 (N_25097,N_23472,N_23546);
nor U25098 (N_25098,N_23854,N_23343);
or U25099 (N_25099,N_23722,N_22937);
or U25100 (N_25100,N_23835,N_23893);
nor U25101 (N_25101,N_22909,N_23961);
nand U25102 (N_25102,N_23711,N_23138);
or U25103 (N_25103,N_23289,N_23006);
nand U25104 (N_25104,N_23177,N_23103);
or U25105 (N_25105,N_23146,N_22899);
xor U25106 (N_25106,N_23432,N_23501);
nand U25107 (N_25107,N_23103,N_23454);
nand U25108 (N_25108,N_23620,N_23851);
nor U25109 (N_25109,N_23379,N_23108);
nor U25110 (N_25110,N_23316,N_23737);
nand U25111 (N_25111,N_23043,N_23807);
or U25112 (N_25112,N_23557,N_23685);
nor U25113 (N_25113,N_23718,N_23772);
nand U25114 (N_25114,N_23746,N_23509);
and U25115 (N_25115,N_23585,N_22988);
or U25116 (N_25116,N_23923,N_23607);
or U25117 (N_25117,N_23273,N_23753);
nor U25118 (N_25118,N_23714,N_23129);
and U25119 (N_25119,N_23270,N_23824);
or U25120 (N_25120,N_23239,N_22861);
nor U25121 (N_25121,N_22916,N_23308);
nor U25122 (N_25122,N_22938,N_23173);
and U25123 (N_25123,N_22844,N_22989);
xor U25124 (N_25124,N_23601,N_23950);
xnor U25125 (N_25125,N_23907,N_23352);
nand U25126 (N_25126,N_22938,N_23400);
nand U25127 (N_25127,N_22997,N_23665);
nand U25128 (N_25128,N_23252,N_22944);
nor U25129 (N_25129,N_23404,N_23571);
nor U25130 (N_25130,N_23709,N_22926);
nand U25131 (N_25131,N_23330,N_23831);
or U25132 (N_25132,N_23606,N_23244);
nor U25133 (N_25133,N_23894,N_23095);
and U25134 (N_25134,N_23338,N_23818);
xnor U25135 (N_25135,N_23141,N_23283);
or U25136 (N_25136,N_23876,N_23336);
and U25137 (N_25137,N_23167,N_23520);
or U25138 (N_25138,N_23511,N_23863);
xnor U25139 (N_25139,N_23903,N_23912);
xnor U25140 (N_25140,N_23827,N_23443);
nand U25141 (N_25141,N_23804,N_23090);
nor U25142 (N_25142,N_23264,N_23262);
nor U25143 (N_25143,N_23241,N_23610);
nor U25144 (N_25144,N_23566,N_23145);
nor U25145 (N_25145,N_23618,N_22938);
nor U25146 (N_25146,N_23849,N_23142);
nor U25147 (N_25147,N_23102,N_23877);
and U25148 (N_25148,N_23241,N_23183);
and U25149 (N_25149,N_23249,N_23786);
nand U25150 (N_25150,N_23279,N_23359);
and U25151 (N_25151,N_23103,N_23292);
nor U25152 (N_25152,N_23831,N_23366);
and U25153 (N_25153,N_23231,N_23661);
or U25154 (N_25154,N_22847,N_23532);
or U25155 (N_25155,N_23255,N_23004);
nor U25156 (N_25156,N_23880,N_23678);
xnor U25157 (N_25157,N_22978,N_23624);
nand U25158 (N_25158,N_23319,N_23270);
or U25159 (N_25159,N_23098,N_23033);
and U25160 (N_25160,N_23073,N_23905);
nand U25161 (N_25161,N_22940,N_23078);
nor U25162 (N_25162,N_23953,N_23382);
and U25163 (N_25163,N_23703,N_23766);
xnor U25164 (N_25164,N_23204,N_23948);
and U25165 (N_25165,N_23299,N_22807);
and U25166 (N_25166,N_23793,N_23777);
xor U25167 (N_25167,N_23828,N_23548);
or U25168 (N_25168,N_22930,N_23744);
nand U25169 (N_25169,N_23701,N_23011);
nor U25170 (N_25170,N_23642,N_23198);
or U25171 (N_25171,N_23288,N_23343);
or U25172 (N_25172,N_22890,N_23474);
xnor U25173 (N_25173,N_23754,N_23471);
nand U25174 (N_25174,N_23044,N_23292);
nand U25175 (N_25175,N_23484,N_23677);
nand U25176 (N_25176,N_23522,N_23661);
and U25177 (N_25177,N_23860,N_23764);
nand U25178 (N_25178,N_23708,N_23352);
xor U25179 (N_25179,N_23338,N_23986);
or U25180 (N_25180,N_23302,N_23497);
xnor U25181 (N_25181,N_23090,N_22871);
or U25182 (N_25182,N_22889,N_23822);
or U25183 (N_25183,N_23808,N_23957);
nor U25184 (N_25184,N_23329,N_23010);
and U25185 (N_25185,N_23461,N_23110);
and U25186 (N_25186,N_22942,N_23880);
nand U25187 (N_25187,N_23800,N_23036);
xor U25188 (N_25188,N_22896,N_23518);
xnor U25189 (N_25189,N_23468,N_22927);
or U25190 (N_25190,N_23133,N_23313);
and U25191 (N_25191,N_23140,N_23448);
nor U25192 (N_25192,N_23157,N_22833);
nor U25193 (N_25193,N_23655,N_23543);
and U25194 (N_25194,N_22978,N_23658);
xnor U25195 (N_25195,N_23720,N_23501);
or U25196 (N_25196,N_23320,N_22851);
xor U25197 (N_25197,N_23470,N_23288);
and U25198 (N_25198,N_23594,N_23381);
or U25199 (N_25199,N_23265,N_23060);
nand U25200 (N_25200,N_24420,N_24760);
or U25201 (N_25201,N_24495,N_24563);
and U25202 (N_25202,N_24077,N_24357);
nand U25203 (N_25203,N_25006,N_25024);
xnor U25204 (N_25204,N_24430,N_24791);
nor U25205 (N_25205,N_25073,N_25121);
or U25206 (N_25206,N_24334,N_25017);
nor U25207 (N_25207,N_24953,N_24094);
nand U25208 (N_25208,N_24893,N_25101);
nand U25209 (N_25209,N_24050,N_24807);
and U25210 (N_25210,N_24510,N_24919);
or U25211 (N_25211,N_25088,N_24913);
or U25212 (N_25212,N_24287,N_24278);
xnor U25213 (N_25213,N_24058,N_24256);
or U25214 (N_25214,N_24659,N_24689);
xor U25215 (N_25215,N_24053,N_24894);
or U25216 (N_25216,N_24683,N_24819);
and U25217 (N_25217,N_24467,N_24498);
and U25218 (N_25218,N_24187,N_24194);
or U25219 (N_25219,N_24654,N_24246);
nor U25220 (N_25220,N_24567,N_25096);
or U25221 (N_25221,N_24959,N_24181);
and U25222 (N_25222,N_24290,N_24776);
nand U25223 (N_25223,N_24419,N_24485);
or U25224 (N_25224,N_24342,N_24642);
nand U25225 (N_25225,N_25156,N_24440);
or U25226 (N_25226,N_24190,N_25183);
or U25227 (N_25227,N_24458,N_25018);
and U25228 (N_25228,N_24782,N_24012);
and U25229 (N_25229,N_24320,N_24144);
and U25230 (N_25230,N_24191,N_25061);
xnor U25231 (N_25231,N_25192,N_24249);
xor U25232 (N_25232,N_24015,N_24716);
nor U25233 (N_25233,N_24656,N_24348);
or U25234 (N_25234,N_24277,N_24956);
nor U25235 (N_25235,N_24666,N_24182);
xor U25236 (N_25236,N_24992,N_24323);
xnor U25237 (N_25237,N_24099,N_24773);
xnor U25238 (N_25238,N_25196,N_24243);
or U25239 (N_25239,N_24818,N_24852);
xnor U25240 (N_25240,N_24925,N_24915);
or U25241 (N_25241,N_24155,N_24410);
nand U25242 (N_25242,N_24763,N_24984);
nand U25243 (N_25243,N_24667,N_24062);
nand U25244 (N_25244,N_25031,N_25152);
nor U25245 (N_25245,N_24281,N_24314);
or U25246 (N_25246,N_24756,N_24944);
xor U25247 (N_25247,N_24068,N_25055);
nand U25248 (N_25248,N_24907,N_24870);
nor U25249 (N_25249,N_25012,N_24384);
xnor U25250 (N_25250,N_24820,N_24890);
xnor U25251 (N_25251,N_24883,N_25130);
or U25252 (N_25252,N_24343,N_24031);
or U25253 (N_25253,N_24257,N_24914);
or U25254 (N_25254,N_24116,N_24680);
nor U25255 (N_25255,N_24599,N_24413);
nand U25256 (N_25256,N_24995,N_24799);
nand U25257 (N_25257,N_24552,N_24911);
nor U25258 (N_25258,N_24114,N_24235);
nand U25259 (N_25259,N_24878,N_24470);
nand U25260 (N_25260,N_24753,N_24073);
or U25261 (N_25261,N_24222,N_24273);
xor U25262 (N_25262,N_25009,N_24316);
nor U25263 (N_25263,N_24494,N_25159);
and U25264 (N_25264,N_24163,N_24950);
nand U25265 (N_25265,N_24091,N_24876);
and U25266 (N_25266,N_24771,N_24034);
nor U25267 (N_25267,N_24141,N_24690);
or U25268 (N_25268,N_24113,N_24267);
and U25269 (N_25269,N_24826,N_24695);
xor U25270 (N_25270,N_24906,N_25056);
nand U25271 (N_25271,N_24171,N_24108);
xnor U25272 (N_25272,N_24941,N_24239);
xnor U25273 (N_25273,N_24213,N_24721);
nor U25274 (N_25274,N_24322,N_24432);
and U25275 (N_25275,N_25100,N_24174);
and U25276 (N_25276,N_24702,N_24148);
or U25277 (N_25277,N_24715,N_24977);
xnor U25278 (N_25278,N_24139,N_24511);
and U25279 (N_25279,N_25072,N_24317);
or U25280 (N_25280,N_24220,N_24052);
or U25281 (N_25281,N_24755,N_25126);
nand U25282 (N_25282,N_24212,N_24547);
and U25283 (N_25283,N_24435,N_24304);
or U25284 (N_25284,N_24308,N_24669);
or U25285 (N_25285,N_25137,N_24581);
or U25286 (N_25286,N_24041,N_25112);
and U25287 (N_25287,N_25172,N_24026);
nor U25288 (N_25288,N_24143,N_24422);
nand U25289 (N_25289,N_25175,N_25180);
or U25290 (N_25290,N_25097,N_24045);
nand U25291 (N_25291,N_24169,N_24577);
nor U25292 (N_25292,N_24223,N_25066);
nand U25293 (N_25293,N_24491,N_24869);
or U25294 (N_25294,N_25118,N_24007);
and U25295 (N_25295,N_24529,N_24947);
and U25296 (N_25296,N_25092,N_24622);
and U25297 (N_25297,N_24728,N_25157);
or U25298 (N_25298,N_24887,N_24969);
and U25299 (N_25299,N_24983,N_25185);
nand U25300 (N_25300,N_24668,N_24391);
nor U25301 (N_25301,N_24395,N_24234);
and U25302 (N_25302,N_24135,N_24789);
or U25303 (N_25303,N_24298,N_24920);
and U25304 (N_25304,N_25188,N_24929);
xnor U25305 (N_25305,N_25090,N_24998);
xor U25306 (N_25306,N_24363,N_24710);
nor U25307 (N_25307,N_24792,N_24801);
nand U25308 (N_25308,N_24228,N_24089);
nand U25309 (N_25309,N_24922,N_24369);
or U25310 (N_25310,N_24788,N_24371);
and U25311 (N_25311,N_24479,N_24347);
and U25312 (N_25312,N_24918,N_24055);
and U25313 (N_25313,N_24978,N_25078);
nor U25314 (N_25314,N_24313,N_25085);
xnor U25315 (N_25315,N_24985,N_24100);
or U25316 (N_25316,N_24092,N_24211);
nand U25317 (N_25317,N_24924,N_24707);
nand U25318 (N_25318,N_24056,N_25014);
or U25319 (N_25319,N_24164,N_25174);
or U25320 (N_25320,N_24508,N_24200);
nand U25321 (N_25321,N_24974,N_24142);
or U25322 (N_25322,N_24451,N_24090);
and U25323 (N_25323,N_24406,N_24898);
or U25324 (N_25324,N_24589,N_24205);
xor U25325 (N_25325,N_24851,N_25178);
or U25326 (N_25326,N_24147,N_24445);
nor U25327 (N_25327,N_24216,N_24838);
or U25328 (N_25328,N_24473,N_25171);
and U25329 (N_25329,N_25140,N_24646);
or U25330 (N_25330,N_24717,N_24949);
nand U25331 (N_25331,N_24963,N_25060);
and U25332 (N_25332,N_24686,N_24916);
nand U25333 (N_25333,N_24688,N_24427);
nand U25334 (N_25334,N_25067,N_24166);
and U25335 (N_25335,N_24566,N_24575);
and U25336 (N_25336,N_24376,N_24812);
or U25337 (N_25337,N_24857,N_24507);
xor U25338 (N_25338,N_25036,N_24904);
or U25339 (N_25339,N_24633,N_24103);
or U25340 (N_25340,N_24475,N_25142);
nand U25341 (N_25341,N_24722,N_24122);
xnor U25342 (N_25342,N_24008,N_24647);
xnor U25343 (N_25343,N_24670,N_24258);
or U25344 (N_25344,N_24204,N_24382);
and U25345 (N_25345,N_24288,N_24970);
and U25346 (N_25346,N_25133,N_25021);
xor U25347 (N_25347,N_24285,N_24576);
nor U25348 (N_25348,N_24241,N_24570);
and U25349 (N_25349,N_24777,N_24331);
xnor U25350 (N_25350,N_24629,N_24390);
and U25351 (N_25351,N_24584,N_25162);
nor U25352 (N_25352,N_24452,N_24787);
xnor U25353 (N_25353,N_24879,N_25143);
xnor U25354 (N_25354,N_24889,N_24850);
nor U25355 (N_25355,N_25032,N_24627);
xor U25356 (N_25356,N_24875,N_24461);
xnor U25357 (N_25357,N_25045,N_24783);
xor U25358 (N_25358,N_24639,N_24083);
and U25359 (N_25359,N_24425,N_24151);
and U25360 (N_25360,N_24496,N_24608);
or U25361 (N_25361,N_24446,N_24559);
xnor U25362 (N_25362,N_24582,N_24110);
and U25363 (N_25363,N_25110,N_24571);
or U25364 (N_25364,N_24469,N_24042);
xor U25365 (N_25365,N_25164,N_24943);
nor U25366 (N_25366,N_24138,N_24810);
nand U25367 (N_25367,N_24772,N_25020);
and U25368 (N_25368,N_24196,N_24193);
or U25369 (N_25369,N_24214,N_25109);
and U25370 (N_25370,N_24655,N_25132);
nand U25371 (N_25371,N_25052,N_24940);
or U25372 (N_25372,N_24242,N_25046);
nor U25373 (N_25373,N_24672,N_24587);
nand U25374 (N_25374,N_25084,N_24134);
nor U25375 (N_25375,N_24534,N_24111);
nand U25376 (N_25376,N_24224,N_24043);
xnor U25377 (N_25377,N_24027,N_24831);
or U25378 (N_25378,N_24794,N_24136);
and U25379 (N_25379,N_24059,N_24928);
nor U25380 (N_25380,N_25022,N_24367);
nor U25381 (N_25381,N_25150,N_24676);
and U25382 (N_25382,N_25113,N_24518);
or U25383 (N_25383,N_25027,N_24610);
xor U25384 (N_25384,N_24407,N_24708);
nand U25385 (N_25385,N_24462,N_25059);
nand U25386 (N_25386,N_25161,N_24024);
xnor U25387 (N_25387,N_25102,N_24945);
nor U25388 (N_25388,N_24021,N_24609);
nand U25389 (N_25389,N_24523,N_24125);
nor U25390 (N_25390,N_24621,N_25124);
or U25391 (N_25391,N_24455,N_24209);
nand U25392 (N_25392,N_24449,N_24431);
or U25393 (N_25393,N_24847,N_24167);
nand U25394 (N_25394,N_25190,N_24279);
nand U25395 (N_25395,N_24364,N_24162);
nor U25396 (N_25396,N_24713,N_24798);
xor U25397 (N_25397,N_24635,N_24482);
nor U25398 (N_25398,N_24165,N_24860);
and U25399 (N_25399,N_24072,N_24653);
xnor U25400 (N_25400,N_24719,N_24591);
and U25401 (N_25401,N_24762,N_25015);
xor U25402 (N_25402,N_24515,N_24671);
nand U25403 (N_25403,N_24044,N_25079);
or U25404 (N_25404,N_24514,N_24490);
nor U25405 (N_25405,N_24814,N_24768);
nand U25406 (N_25406,N_24752,N_25122);
or U25407 (N_25407,N_24102,N_24555);
and U25408 (N_25408,N_24856,N_24868);
or U25409 (N_25409,N_24657,N_24551);
or U25410 (N_25410,N_24471,N_24502);
nand U25411 (N_25411,N_24971,N_24793);
xor U25412 (N_25412,N_24442,N_24892);
xnor U25413 (N_25413,N_24311,N_24675);
and U25414 (N_25414,N_24808,N_25075);
nor U25415 (N_25415,N_24176,N_24408);
and U25416 (N_25416,N_24538,N_24554);
nor U25417 (N_25417,N_24612,N_25039);
xnor U25418 (N_25418,N_24393,N_24806);
and U25419 (N_25419,N_25080,N_24037);
or U25420 (N_25420,N_24981,N_24416);
nand U25421 (N_25421,N_24834,N_24293);
nand U25422 (N_25422,N_24961,N_25194);
and U25423 (N_25423,N_24085,N_24699);
nor U25424 (N_25424,N_25123,N_24417);
xnor U25425 (N_25425,N_24254,N_25111);
or U25426 (N_25426,N_24816,N_24319);
and U25427 (N_25427,N_24556,N_24387);
or U25428 (N_25428,N_25070,N_24292);
xor U25429 (N_25429,N_24275,N_25103);
nor U25430 (N_25430,N_24268,N_25026);
xor U25431 (N_25431,N_24312,N_24450);
xnor U25432 (N_25432,N_24271,N_24607);
and U25433 (N_25433,N_25034,N_24412);
nand U25434 (N_25434,N_24486,N_24931);
nand U25435 (N_25435,N_24874,N_24714);
and U25436 (N_25436,N_24594,N_24561);
nand U25437 (N_25437,N_24010,N_24638);
nand U25438 (N_25438,N_24877,N_24968);
nand U25439 (N_25439,N_24624,N_24861);
or U25440 (N_25440,N_24660,N_24872);
xor U25441 (N_25441,N_24542,N_25002);
and U25442 (N_25442,N_25179,N_24780);
xor U25443 (N_25443,N_24185,N_24201);
xor U25444 (N_25444,N_24679,N_24528);
or U25445 (N_25445,N_24824,N_24039);
nor U25446 (N_25446,N_24465,N_24444);
nand U25447 (N_25447,N_24378,N_24140);
xnor U25448 (N_25448,N_24512,N_24900);
nand U25449 (N_25449,N_24404,N_24543);
and U25450 (N_25450,N_25141,N_24909);
xor U25451 (N_25451,N_24997,N_24521);
and U25452 (N_25452,N_25038,N_25003);
nand U25453 (N_25453,N_24453,N_24746);
nor U25454 (N_25454,N_24020,N_24177);
nand U25455 (N_25455,N_24385,N_24310);
nor U25456 (N_25456,N_24480,N_24456);
or U25457 (N_25457,N_24749,N_24937);
nor U25458 (N_25458,N_24013,N_25160);
nand U25459 (N_25459,N_24828,N_24305);
and U25460 (N_25460,N_24544,N_24373);
xor U25461 (N_25461,N_24006,N_24520);
nor U25462 (N_25462,N_24979,N_24955);
xnor U25463 (N_25463,N_25091,N_24345);
nor U25464 (N_25464,N_24705,N_24137);
nand U25465 (N_25465,N_24299,N_25004);
nor U25466 (N_25466,N_24226,N_25041);
or U25467 (N_25467,N_24586,N_25098);
or U25468 (N_25468,N_24358,N_25145);
or U25469 (N_25469,N_24614,N_25107);
or U25470 (N_25470,N_24886,N_24743);
or U25471 (N_25471,N_24082,N_24218);
xor U25472 (N_25472,N_24296,N_24558);
and U25473 (N_25473,N_24697,N_24179);
xnor U25474 (N_25474,N_25199,N_25125);
and U25475 (N_25475,N_24036,N_24127);
nor U25476 (N_25476,N_24232,N_24238);
nand U25477 (N_25477,N_24687,N_24063);
nand U25478 (N_25478,N_24074,N_24199);
nand U25479 (N_25479,N_24161,N_24797);
nand U25480 (N_25480,N_24380,N_25082);
nand U25481 (N_25481,N_24623,N_25153);
xor U25482 (N_25482,N_25104,N_24863);
or U25483 (N_25483,N_24723,N_24615);
and U25484 (N_25484,N_24854,N_24303);
nor U25485 (N_25485,N_24152,N_24805);
nand U25486 (N_25486,N_25115,N_24202);
xnor U25487 (N_25487,N_24328,N_24734);
nor U25488 (N_25488,N_24236,N_24078);
and U25489 (N_25489,N_24500,N_24002);
and U25490 (N_25490,N_24188,N_24901);
nor U25491 (N_25491,N_24645,N_24375);
nand U25492 (N_25492,N_24497,N_24712);
nor U25493 (N_25493,N_24982,N_24770);
or U25494 (N_25494,N_24175,N_24437);
and U25495 (N_25495,N_24389,N_24168);
nor U25496 (N_25496,N_24960,N_24405);
or U25497 (N_25497,N_24748,N_24862);
or U25498 (N_25498,N_24460,N_24180);
xor U25499 (N_25499,N_24291,N_24821);
or U25500 (N_25500,N_24372,N_24329);
nand U25501 (N_25501,N_24882,N_24952);
xor U25502 (N_25502,N_24517,N_24219);
nor U25503 (N_25503,N_24744,N_25037);
xnor U25504 (N_25504,N_24815,N_24733);
nor U25505 (N_25505,N_24619,N_24774);
nor U25506 (N_25506,N_24145,N_24421);
or U25507 (N_25507,N_24014,N_24738);
and U25508 (N_25508,N_24433,N_24912);
or U25509 (N_25509,N_24933,N_24764);
nand U25510 (N_25510,N_24921,N_24210);
or U25511 (N_25511,N_24183,N_24441);
nand U25512 (N_25512,N_25043,N_24597);
and U25513 (N_25513,N_24093,N_24240);
or U25514 (N_25514,N_25010,N_24084);
and U25515 (N_25515,N_24335,N_24418);
nor U25516 (N_25516,N_24637,N_24352);
nand U25517 (N_25517,N_24562,N_25093);
nor U25518 (N_25518,N_24107,N_24739);
nand U25519 (N_25519,N_24540,N_24694);
xnor U25520 (N_25520,N_24360,N_24098);
xor U25521 (N_25521,N_24905,N_24550);
xor U25522 (N_25522,N_25065,N_24402);
or U25523 (N_25523,N_24840,N_24079);
xor U25524 (N_25524,N_25069,N_25105);
and U25525 (N_25525,N_24761,N_24097);
nand U25526 (N_25526,N_25170,N_24344);
nand U25527 (N_25527,N_25001,N_24459);
xnor U25528 (N_25528,N_24972,N_24379);
nand U25529 (N_25529,N_24809,N_24665);
nand U25530 (N_25530,N_24018,N_24381);
or U25531 (N_25531,N_25129,N_24632);
and U25532 (N_25532,N_24936,N_24903);
and U25533 (N_25533,N_24750,N_24374);
or U25534 (N_25534,N_24252,N_24880);
xnor U25535 (N_25535,N_24778,N_24549);
or U25536 (N_25536,N_24326,N_24602);
xor U25537 (N_25537,N_24075,N_24192);
nor U25538 (N_25538,N_24172,N_25086);
nor U25539 (N_25539,N_25063,N_24560);
or U25540 (N_25540,N_24836,N_24030);
and U25541 (N_25541,N_24765,N_24255);
or U25542 (N_25542,N_24221,N_24966);
xnor U25543 (N_25543,N_24813,N_24366);
and U25544 (N_25544,N_24902,N_24829);
and U25545 (N_25545,N_24265,N_24701);
or U25546 (N_25546,N_24718,N_24737);
nor U25547 (N_25547,N_24546,N_24132);
nor U25548 (N_25548,N_25187,N_24917);
nor U25549 (N_25549,N_24259,N_24476);
and U25550 (N_25550,N_24307,N_24025);
nand U25551 (N_25551,N_24698,N_24726);
and U25552 (N_25552,N_24842,N_24759);
nor U25553 (N_25553,N_25033,N_24585);
or U25554 (N_25554,N_25131,N_24678);
nand U25555 (N_25555,N_24302,N_24150);
or U25556 (N_25556,N_24897,N_25182);
nand U25557 (N_25557,N_24859,N_24351);
nor U25558 (N_25558,N_25177,N_24853);
nand U25559 (N_25559,N_24117,N_25163);
nand U25560 (N_25560,N_24361,N_24409);
nand U25561 (N_25561,N_24684,N_24841);
nand U25562 (N_25562,N_24785,N_24855);
nand U25563 (N_25563,N_24871,N_24208);
nand U25564 (N_25564,N_24600,N_24336);
and U25565 (N_25565,N_25127,N_24505);
xnor U25566 (N_25566,N_25116,N_25184);
xnor U25567 (N_25567,N_24873,N_24827);
or U25568 (N_25568,N_25158,N_24341);
and U25569 (N_25569,N_24578,N_24965);
or U25570 (N_25570,N_24895,N_24681);
xor U25571 (N_25571,N_24595,N_24867);
and U25572 (N_25572,N_24839,N_24054);
or U25573 (N_25573,N_24617,N_24244);
and U25574 (N_25574,N_24439,N_25146);
nor U25575 (N_25575,N_25042,N_24910);
nand U25576 (N_25576,N_25197,N_24049);
nand U25577 (N_25577,N_24203,N_24325);
and U25578 (N_25578,N_24253,N_24081);
nor U25579 (N_25579,N_24038,N_24128);
xor U25580 (N_25580,N_25016,N_24489);
xor U25581 (N_25581,N_24962,N_24849);
and U25582 (N_25582,N_24133,N_24356);
nand U25583 (N_25583,N_24817,N_24926);
xnor U25584 (N_25584,N_24991,N_24332);
or U25585 (N_25585,N_24086,N_24368);
or U25586 (N_25586,N_24060,N_25198);
xnor U25587 (N_25587,N_24796,N_24330);
nor U25588 (N_25588,N_24740,N_24896);
xor U25589 (N_25589,N_24016,N_24158);
nand U25590 (N_25590,N_24397,N_24823);
nand U25591 (N_25591,N_25166,N_24438);
or U25592 (N_25592,N_25094,N_24539);
or U25593 (N_25593,N_25189,N_24758);
and U25594 (N_25594,N_24644,N_24386);
xor U25595 (N_25595,N_24009,N_24333);
and U25596 (N_25596,N_24598,N_24229);
xor U25597 (N_25597,N_24848,N_24530);
or U25598 (N_25598,N_24124,N_25068);
nand U25599 (N_25599,N_24383,N_24269);
nand U25600 (N_25600,N_24263,N_24548);
xor U25601 (N_25601,N_24786,N_24927);
nor U25602 (N_25602,N_24301,N_25193);
xor U25603 (N_25603,N_24251,N_25077);
and U25604 (N_25604,N_24579,N_24935);
or U25605 (N_25605,N_24477,N_24464);
nand U25606 (N_25606,N_24662,N_24939);
xor U25607 (N_25607,N_24975,N_24264);
nor U25608 (N_25608,N_25007,N_24651);
nand U25609 (N_25609,N_24938,N_24742);
xnor U25610 (N_25610,N_24023,N_24033);
and U25611 (N_25611,N_25195,N_24350);
nor U25612 (N_25612,N_24130,N_24664);
nor U25613 (N_25613,N_24596,N_24483);
and U25614 (N_25614,N_24362,N_24466);
and U25615 (N_25615,N_24000,N_24403);
xor U25616 (N_25616,N_24019,N_24973);
xor U25617 (N_25617,N_24028,N_24885);
and U25618 (N_25618,N_25044,N_24625);
and U25619 (N_25619,N_25147,N_24833);
xor U25620 (N_25620,N_24105,N_24423);
or U25621 (N_25621,N_24958,N_25099);
or U25622 (N_25622,N_24118,N_24711);
nor U25623 (N_25623,N_25030,N_24845);
nor U25624 (N_25624,N_24004,N_24643);
xor U25625 (N_25625,N_24565,N_24640);
and U25626 (N_25626,N_24706,N_24076);
nor U25627 (N_25627,N_24864,N_24757);
and U25628 (N_25628,N_24170,N_24631);
xnor U25629 (N_25629,N_24215,N_24198);
and U25630 (N_25630,N_24230,N_24994);
or U25631 (N_25631,N_24153,N_24583);
or U25632 (N_25632,N_24067,N_24365);
and U25633 (N_25633,N_24295,N_24022);
xnor U25634 (N_25634,N_24121,N_24283);
nand U25635 (N_25635,N_24724,N_25047);
nor U25636 (N_25636,N_24414,N_24231);
xnor U25637 (N_25637,N_24472,N_24865);
or U25638 (N_25638,N_24564,N_24096);
and U25639 (N_25639,N_24065,N_24468);
nor U25640 (N_25640,N_24248,N_24499);
or U25641 (N_25641,N_24154,N_24428);
nor U25642 (N_25642,N_25095,N_24411);
nand U25643 (N_25643,N_24131,N_25083);
nand U25644 (N_25644,N_24891,N_24399);
nor U25645 (N_25645,N_25005,N_24324);
and U25646 (N_25646,N_24106,N_24001);
and U25647 (N_25647,N_24747,N_24394);
nor U25648 (N_25648,N_24488,N_25186);
nor U25649 (N_25649,N_24173,N_24487);
nand U25650 (N_25650,N_24844,N_24272);
or U25651 (N_25651,N_24297,N_24159);
or U25652 (N_25652,N_25062,N_24519);
nor U25653 (N_25653,N_24703,N_24648);
and U25654 (N_25654,N_24524,N_24769);
xor U25655 (N_25655,N_25135,N_24531);
nand U25656 (N_25656,N_24605,N_24337);
nand U25657 (N_25657,N_25013,N_25028);
or U25658 (N_25658,N_24825,N_24047);
xnor U25659 (N_25659,N_24282,N_25035);
nand U25660 (N_25660,N_24156,N_25050);
and U25661 (N_25661,N_25058,N_24976);
nor U25662 (N_25662,N_24704,N_24730);
nand U25663 (N_25663,N_24513,N_25165);
nor U25664 (N_25664,N_24673,N_24447);
xor U25665 (N_25665,N_25053,N_24967);
or U25666 (N_25666,N_24501,N_24104);
nand U25667 (N_25667,N_24247,N_24064);
nand U25668 (N_25668,N_24005,N_24736);
xor U25669 (N_25669,N_24184,N_24709);
and U25670 (N_25670,N_24088,N_24040);
or U25671 (N_25671,N_24634,N_24318);
nand U25672 (N_25672,N_24795,N_24980);
xor U25673 (N_25673,N_24988,N_24729);
xnor U25674 (N_25674,N_24276,N_24934);
and U25675 (N_25675,N_24930,N_24115);
nand U25676 (N_25676,N_24781,N_24286);
nand U25677 (N_25677,N_24129,N_24593);
nor U25678 (N_25678,N_24948,N_24509);
nor U25679 (N_25679,N_24415,N_24745);
xnor U25680 (N_25680,N_24603,N_24537);
nand U25681 (N_25681,N_24463,N_24061);
xnor U25682 (N_25682,N_24630,N_24533);
or U25683 (N_25683,N_24964,N_24685);
nand U25684 (N_25684,N_24066,N_24436);
nand U25685 (N_25685,N_24993,N_24954);
or U25686 (N_25686,N_24658,N_24613);
xor U25687 (N_25687,N_24606,N_24484);
nand U25688 (N_25688,N_24951,N_25049);
nor U25689 (N_25689,N_24346,N_24720);
or U25690 (N_25690,N_24398,N_24569);
xnor U25691 (N_25691,N_24327,N_24588);
nor U25692 (N_25692,N_24990,N_24503);
and U25693 (N_25693,N_24641,N_24315);
or U25694 (N_25694,N_25087,N_24700);
and U25695 (N_25695,N_24035,N_24999);
or U25696 (N_25696,N_24693,N_25169);
or U25697 (N_25697,N_25138,N_24946);
xor U25698 (N_25698,N_24123,N_24207);
and U25699 (N_25699,N_25025,N_24830);
xor U25700 (N_25700,N_24652,N_24899);
nand U25701 (N_25701,N_24957,N_24618);
xor U25702 (N_25702,N_24811,N_24696);
or U25703 (N_25703,N_25106,N_24822);
xor U25704 (N_25704,N_24048,N_24775);
and U25705 (N_25705,N_24359,N_24580);
xor U25706 (N_25706,N_24274,N_24766);
nand U25707 (N_25707,N_25076,N_24197);
nand U25708 (N_25708,N_25114,N_24800);
nor U25709 (N_25709,N_24426,N_25181);
nand U25710 (N_25710,N_24545,N_24835);
or U25711 (N_25711,N_24029,N_24881);
xor U25712 (N_25712,N_24604,N_24535);
xnor U25713 (N_25713,N_24186,N_25176);
nand U25714 (N_25714,N_24392,N_24069);
nor U25715 (N_25715,N_24626,N_24837);
nor U25716 (N_25716,N_24126,N_24011);
nor U25717 (N_25717,N_24516,N_24932);
or U25718 (N_25718,N_25119,N_24087);
and U25719 (N_25719,N_24732,N_24017);
or U25720 (N_25720,N_24250,N_24057);
and U25721 (N_25721,N_24846,N_24590);
xnor U25722 (N_25722,N_24741,N_24987);
or U25723 (N_25723,N_24616,N_24306);
and U25724 (N_25724,N_24506,N_24112);
or U25725 (N_25725,N_24400,N_24650);
nor U25726 (N_25726,N_24843,N_24429);
xor U25727 (N_25727,N_24051,N_24522);
or U25728 (N_25728,N_25108,N_24481);
and U25729 (N_25729,N_25019,N_24611);
xnor U25730 (N_25730,N_24095,N_24266);
nand U25731 (N_25731,N_24474,N_24443);
or U25732 (N_25732,N_25057,N_24178);
xnor U25733 (N_25733,N_24986,N_24492);
and U25734 (N_25734,N_24080,N_25117);
nor U25735 (N_25735,N_24284,N_25136);
nand U25736 (N_25736,N_24541,N_25081);
nand U25737 (N_25737,N_24189,N_24270);
or U25738 (N_25738,N_24572,N_25023);
or U25739 (N_25739,N_24434,N_24804);
or U25740 (N_25740,N_24620,N_25168);
and U25741 (N_25741,N_25148,N_24691);
and U25742 (N_25742,N_25051,N_24070);
xnor U25743 (N_25743,N_24923,N_24233);
nor U25744 (N_25744,N_24339,N_24553);
nor U25745 (N_25745,N_25154,N_25167);
nor U25746 (N_25746,N_24206,N_24454);
or U25747 (N_25747,N_24349,N_24803);
or U25748 (N_25748,N_24260,N_24888);
and U25749 (N_25749,N_24526,N_24309);
and U25750 (N_25750,N_24751,N_24388);
nand U25751 (N_25751,N_24790,N_25029);
or U25752 (N_25752,N_25000,N_24767);
nand U25753 (N_25753,N_25064,N_24802);
xor U25754 (N_25754,N_24727,N_24109);
nand U25755 (N_25755,N_24663,N_24525);
xor U25756 (N_25756,N_24225,N_25151);
nand U25757 (N_25757,N_24294,N_24448);
xor U25758 (N_25758,N_24592,N_24504);
nor U25759 (N_25759,N_24353,N_24731);
nor U25760 (N_25760,N_24338,N_24568);
and U25761 (N_25761,N_24377,N_24649);
nor U25762 (N_25762,N_24457,N_24478);
and U25763 (N_25763,N_24157,N_24527);
and U25764 (N_25764,N_24262,N_24661);
nor U25765 (N_25765,N_24401,N_24942);
and U25766 (N_25766,N_25008,N_25120);
nand U25767 (N_25767,N_24784,N_24280);
nand U25768 (N_25768,N_24340,N_24227);
and U25769 (N_25769,N_25074,N_24101);
or U25770 (N_25770,N_25071,N_24160);
nor U25771 (N_25771,N_24354,N_24725);
or U25772 (N_25772,N_24321,N_24119);
and U25773 (N_25773,N_25191,N_24908);
nor U25774 (N_25774,N_24601,N_24536);
or U25775 (N_25775,N_25149,N_24866);
and U25776 (N_25776,N_24682,N_25173);
nand U25777 (N_25777,N_24636,N_24355);
xor U25778 (N_25778,N_24832,N_24989);
nand U25779 (N_25779,N_25128,N_24628);
xor U25780 (N_25780,N_24120,N_24032);
or U25781 (N_25781,N_25048,N_24370);
or U25782 (N_25782,N_24573,N_24754);
and U25783 (N_25783,N_24237,N_24674);
nand U25784 (N_25784,N_24149,N_25054);
nand U25785 (N_25785,N_25139,N_25040);
nand U25786 (N_25786,N_24261,N_24071);
and U25787 (N_25787,N_24300,N_25089);
or U25788 (N_25788,N_24396,N_24735);
or U25789 (N_25789,N_24557,N_25011);
nand U25790 (N_25790,N_25134,N_24146);
nand U25791 (N_25791,N_24289,N_24677);
nand U25792 (N_25792,N_24493,N_24424);
and U25793 (N_25793,N_24046,N_24195);
xnor U25794 (N_25794,N_24779,N_24884);
xnor U25795 (N_25795,N_24003,N_24217);
nand U25796 (N_25796,N_24245,N_24858);
xor U25797 (N_25797,N_24996,N_25155);
and U25798 (N_25798,N_25144,N_24532);
nand U25799 (N_25799,N_24692,N_24574);
nor U25800 (N_25800,N_24990,N_24188);
xor U25801 (N_25801,N_25148,N_24640);
nor U25802 (N_25802,N_24265,N_24781);
and U25803 (N_25803,N_24715,N_24544);
nor U25804 (N_25804,N_24681,N_24164);
nand U25805 (N_25805,N_24342,N_24273);
or U25806 (N_25806,N_24319,N_24507);
nand U25807 (N_25807,N_24102,N_25095);
nand U25808 (N_25808,N_24669,N_24250);
nand U25809 (N_25809,N_24622,N_24695);
nor U25810 (N_25810,N_24772,N_24625);
nand U25811 (N_25811,N_24138,N_24682);
nand U25812 (N_25812,N_24222,N_24359);
nor U25813 (N_25813,N_24852,N_25021);
nand U25814 (N_25814,N_24877,N_24162);
xor U25815 (N_25815,N_24099,N_24655);
nor U25816 (N_25816,N_24183,N_24452);
nand U25817 (N_25817,N_24528,N_24253);
and U25818 (N_25818,N_24810,N_24497);
nor U25819 (N_25819,N_24822,N_24027);
nand U25820 (N_25820,N_24637,N_24482);
or U25821 (N_25821,N_25130,N_25137);
and U25822 (N_25822,N_24724,N_24743);
xor U25823 (N_25823,N_24874,N_24322);
or U25824 (N_25824,N_24795,N_24508);
nand U25825 (N_25825,N_24710,N_25162);
and U25826 (N_25826,N_24715,N_24948);
nor U25827 (N_25827,N_24398,N_24816);
nand U25828 (N_25828,N_24465,N_25155);
nor U25829 (N_25829,N_24345,N_24654);
or U25830 (N_25830,N_24359,N_24915);
and U25831 (N_25831,N_24494,N_24472);
or U25832 (N_25832,N_24542,N_24396);
and U25833 (N_25833,N_24626,N_24394);
nand U25834 (N_25834,N_24213,N_24266);
and U25835 (N_25835,N_24478,N_24178);
or U25836 (N_25836,N_24144,N_25190);
xnor U25837 (N_25837,N_24258,N_25010);
and U25838 (N_25838,N_24709,N_24571);
or U25839 (N_25839,N_24565,N_24376);
nor U25840 (N_25840,N_24166,N_24966);
or U25841 (N_25841,N_24922,N_24523);
xnor U25842 (N_25842,N_24916,N_24615);
or U25843 (N_25843,N_24249,N_24192);
nor U25844 (N_25844,N_25187,N_25066);
xnor U25845 (N_25845,N_24297,N_24288);
or U25846 (N_25846,N_24813,N_25121);
nor U25847 (N_25847,N_24486,N_24045);
nand U25848 (N_25848,N_24966,N_24099);
or U25849 (N_25849,N_24431,N_24823);
xnor U25850 (N_25850,N_24137,N_24871);
nand U25851 (N_25851,N_24863,N_25186);
nand U25852 (N_25852,N_24245,N_24208);
xor U25853 (N_25853,N_24661,N_24343);
or U25854 (N_25854,N_25143,N_25074);
nand U25855 (N_25855,N_24730,N_24594);
xnor U25856 (N_25856,N_24575,N_24516);
nor U25857 (N_25857,N_24582,N_24214);
and U25858 (N_25858,N_24402,N_24496);
nor U25859 (N_25859,N_24403,N_24840);
nand U25860 (N_25860,N_25093,N_24919);
or U25861 (N_25861,N_24187,N_24430);
nor U25862 (N_25862,N_24671,N_24733);
nand U25863 (N_25863,N_25060,N_24322);
xnor U25864 (N_25864,N_24552,N_25082);
xor U25865 (N_25865,N_24014,N_25134);
and U25866 (N_25866,N_24204,N_24827);
and U25867 (N_25867,N_24323,N_24590);
xnor U25868 (N_25868,N_24903,N_24311);
or U25869 (N_25869,N_24829,N_24144);
nor U25870 (N_25870,N_24503,N_24936);
nor U25871 (N_25871,N_24820,N_24277);
nand U25872 (N_25872,N_24149,N_24813);
or U25873 (N_25873,N_25083,N_24766);
and U25874 (N_25874,N_24980,N_24136);
and U25875 (N_25875,N_24142,N_24105);
nor U25876 (N_25876,N_24523,N_24433);
and U25877 (N_25877,N_25044,N_24735);
xnor U25878 (N_25878,N_25188,N_24232);
nand U25879 (N_25879,N_24570,N_24114);
nand U25880 (N_25880,N_24636,N_24575);
and U25881 (N_25881,N_24935,N_24971);
nor U25882 (N_25882,N_24824,N_24274);
or U25883 (N_25883,N_24343,N_24241);
nor U25884 (N_25884,N_24572,N_24355);
nand U25885 (N_25885,N_24451,N_24365);
and U25886 (N_25886,N_24654,N_24392);
or U25887 (N_25887,N_24008,N_25048);
or U25888 (N_25888,N_25164,N_24370);
nand U25889 (N_25889,N_24508,N_24048);
nor U25890 (N_25890,N_24800,N_24022);
or U25891 (N_25891,N_24874,N_25159);
and U25892 (N_25892,N_24708,N_24744);
nor U25893 (N_25893,N_24182,N_24729);
nand U25894 (N_25894,N_24256,N_24039);
and U25895 (N_25895,N_24117,N_25151);
or U25896 (N_25896,N_24366,N_25063);
xnor U25897 (N_25897,N_25184,N_24161);
and U25898 (N_25898,N_25084,N_24579);
nor U25899 (N_25899,N_24543,N_24599);
or U25900 (N_25900,N_24315,N_24221);
and U25901 (N_25901,N_24629,N_24048);
nor U25902 (N_25902,N_25168,N_25019);
or U25903 (N_25903,N_24695,N_24216);
or U25904 (N_25904,N_25103,N_24785);
nand U25905 (N_25905,N_24109,N_24675);
and U25906 (N_25906,N_24424,N_24257);
or U25907 (N_25907,N_24919,N_24072);
and U25908 (N_25908,N_24987,N_24091);
xor U25909 (N_25909,N_24551,N_24573);
nand U25910 (N_25910,N_24016,N_24660);
or U25911 (N_25911,N_24418,N_24659);
nand U25912 (N_25912,N_24851,N_24589);
or U25913 (N_25913,N_25180,N_24877);
nor U25914 (N_25914,N_24209,N_24680);
or U25915 (N_25915,N_24358,N_25158);
and U25916 (N_25916,N_24675,N_24404);
nor U25917 (N_25917,N_24446,N_24692);
xnor U25918 (N_25918,N_24366,N_24659);
xnor U25919 (N_25919,N_24580,N_24726);
xnor U25920 (N_25920,N_24700,N_25019);
xnor U25921 (N_25921,N_24296,N_24356);
nand U25922 (N_25922,N_24738,N_24292);
or U25923 (N_25923,N_24864,N_24248);
or U25924 (N_25924,N_24311,N_24593);
or U25925 (N_25925,N_24456,N_24908);
and U25926 (N_25926,N_24291,N_24737);
and U25927 (N_25927,N_24452,N_24467);
and U25928 (N_25928,N_24604,N_24716);
xnor U25929 (N_25929,N_24543,N_24679);
or U25930 (N_25930,N_24446,N_25165);
nand U25931 (N_25931,N_24306,N_25166);
and U25932 (N_25932,N_24747,N_24279);
and U25933 (N_25933,N_24202,N_24121);
or U25934 (N_25934,N_24416,N_24385);
xor U25935 (N_25935,N_24500,N_24516);
xnor U25936 (N_25936,N_24711,N_24057);
nand U25937 (N_25937,N_24507,N_24268);
and U25938 (N_25938,N_24360,N_24462);
xnor U25939 (N_25939,N_24471,N_24038);
and U25940 (N_25940,N_24155,N_24788);
nand U25941 (N_25941,N_24709,N_24820);
nand U25942 (N_25942,N_24625,N_24278);
nand U25943 (N_25943,N_24432,N_24115);
nor U25944 (N_25944,N_24492,N_24955);
and U25945 (N_25945,N_24236,N_24083);
nand U25946 (N_25946,N_24400,N_24852);
nand U25947 (N_25947,N_24695,N_24599);
nor U25948 (N_25948,N_24998,N_24638);
nor U25949 (N_25949,N_24016,N_25175);
or U25950 (N_25950,N_24124,N_24318);
nor U25951 (N_25951,N_24160,N_24164);
and U25952 (N_25952,N_24288,N_24749);
nand U25953 (N_25953,N_24551,N_24962);
or U25954 (N_25954,N_25140,N_24161);
or U25955 (N_25955,N_24852,N_24361);
and U25956 (N_25956,N_24992,N_24300);
xor U25957 (N_25957,N_24152,N_24739);
or U25958 (N_25958,N_24627,N_24127);
and U25959 (N_25959,N_25114,N_25066);
and U25960 (N_25960,N_25031,N_24226);
and U25961 (N_25961,N_24647,N_24811);
and U25962 (N_25962,N_24548,N_24995);
and U25963 (N_25963,N_24857,N_24318);
and U25964 (N_25964,N_24183,N_24971);
nand U25965 (N_25965,N_24092,N_24193);
or U25966 (N_25966,N_25153,N_24180);
and U25967 (N_25967,N_24393,N_24568);
xor U25968 (N_25968,N_24144,N_24032);
nand U25969 (N_25969,N_24798,N_24454);
xor U25970 (N_25970,N_24576,N_24700);
or U25971 (N_25971,N_25089,N_24893);
or U25972 (N_25972,N_25005,N_24100);
and U25973 (N_25973,N_24810,N_24144);
and U25974 (N_25974,N_25116,N_24080);
xor U25975 (N_25975,N_24781,N_25096);
or U25976 (N_25976,N_25198,N_24176);
nand U25977 (N_25977,N_24511,N_24600);
nand U25978 (N_25978,N_24269,N_24644);
and U25979 (N_25979,N_24399,N_24759);
xnor U25980 (N_25980,N_24814,N_24987);
or U25981 (N_25981,N_24038,N_24812);
or U25982 (N_25982,N_24561,N_24582);
and U25983 (N_25983,N_24424,N_24811);
xnor U25984 (N_25984,N_24730,N_24616);
and U25985 (N_25985,N_24877,N_24712);
or U25986 (N_25986,N_24806,N_24528);
nand U25987 (N_25987,N_24302,N_24598);
xor U25988 (N_25988,N_24282,N_24677);
nand U25989 (N_25989,N_24175,N_24507);
xnor U25990 (N_25990,N_24295,N_24217);
and U25991 (N_25991,N_24592,N_24024);
xnor U25992 (N_25992,N_24459,N_24494);
xnor U25993 (N_25993,N_24583,N_24521);
nand U25994 (N_25994,N_24517,N_25171);
and U25995 (N_25995,N_25147,N_24029);
xnor U25996 (N_25996,N_24760,N_24417);
xnor U25997 (N_25997,N_24260,N_24369);
and U25998 (N_25998,N_25068,N_24044);
nor U25999 (N_25999,N_25145,N_24325);
nor U26000 (N_26000,N_24655,N_25180);
and U26001 (N_26001,N_25132,N_25195);
nor U26002 (N_26002,N_24332,N_24134);
xnor U26003 (N_26003,N_24646,N_24804);
xor U26004 (N_26004,N_24210,N_24194);
xor U26005 (N_26005,N_24883,N_24987);
xnor U26006 (N_26006,N_24484,N_24614);
or U26007 (N_26007,N_24285,N_24019);
nand U26008 (N_26008,N_25112,N_24392);
nand U26009 (N_26009,N_24055,N_24403);
and U26010 (N_26010,N_24888,N_24671);
nand U26011 (N_26011,N_25163,N_24466);
or U26012 (N_26012,N_24843,N_24745);
or U26013 (N_26013,N_24152,N_24728);
nor U26014 (N_26014,N_25075,N_24190);
and U26015 (N_26015,N_24754,N_24685);
nor U26016 (N_26016,N_25065,N_24040);
nor U26017 (N_26017,N_24954,N_24639);
nor U26018 (N_26018,N_24214,N_24003);
xor U26019 (N_26019,N_24845,N_25098);
and U26020 (N_26020,N_24777,N_24537);
nor U26021 (N_26021,N_24556,N_25086);
or U26022 (N_26022,N_24958,N_24499);
nand U26023 (N_26023,N_24975,N_24079);
and U26024 (N_26024,N_24334,N_24481);
and U26025 (N_26025,N_24718,N_24241);
and U26026 (N_26026,N_24866,N_24717);
or U26027 (N_26027,N_25102,N_24875);
nor U26028 (N_26028,N_24985,N_24199);
and U26029 (N_26029,N_25003,N_24335);
or U26030 (N_26030,N_25019,N_25146);
nor U26031 (N_26031,N_24519,N_24725);
nor U26032 (N_26032,N_24064,N_24849);
or U26033 (N_26033,N_24106,N_24320);
and U26034 (N_26034,N_24472,N_25146);
or U26035 (N_26035,N_24844,N_24908);
xor U26036 (N_26036,N_24327,N_24081);
nor U26037 (N_26037,N_24349,N_24258);
and U26038 (N_26038,N_25125,N_24739);
and U26039 (N_26039,N_25084,N_24655);
xnor U26040 (N_26040,N_24408,N_24561);
or U26041 (N_26041,N_25049,N_25179);
nand U26042 (N_26042,N_24321,N_24572);
and U26043 (N_26043,N_24768,N_24017);
nand U26044 (N_26044,N_24320,N_24171);
nor U26045 (N_26045,N_24793,N_24791);
xnor U26046 (N_26046,N_24377,N_25069);
xnor U26047 (N_26047,N_25155,N_24173);
and U26048 (N_26048,N_24894,N_24607);
xnor U26049 (N_26049,N_24954,N_24362);
and U26050 (N_26050,N_24844,N_25182);
or U26051 (N_26051,N_24725,N_24381);
or U26052 (N_26052,N_24025,N_25017);
and U26053 (N_26053,N_24746,N_24190);
xnor U26054 (N_26054,N_25103,N_24042);
nand U26055 (N_26055,N_24559,N_24595);
nor U26056 (N_26056,N_25031,N_24311);
nor U26057 (N_26057,N_24353,N_24120);
or U26058 (N_26058,N_24760,N_24647);
nor U26059 (N_26059,N_24093,N_24197);
xnor U26060 (N_26060,N_24291,N_24475);
or U26061 (N_26061,N_24865,N_24927);
xnor U26062 (N_26062,N_24862,N_24294);
xor U26063 (N_26063,N_25096,N_25134);
or U26064 (N_26064,N_25155,N_24012);
or U26065 (N_26065,N_24289,N_24535);
xor U26066 (N_26066,N_24365,N_24804);
xnor U26067 (N_26067,N_24088,N_24189);
nand U26068 (N_26068,N_24295,N_24761);
nand U26069 (N_26069,N_24645,N_24000);
nand U26070 (N_26070,N_25089,N_24237);
nand U26071 (N_26071,N_24949,N_24652);
nor U26072 (N_26072,N_24987,N_25108);
nand U26073 (N_26073,N_24621,N_25166);
nor U26074 (N_26074,N_24333,N_24751);
xor U26075 (N_26075,N_24738,N_24016);
or U26076 (N_26076,N_24876,N_24070);
nand U26077 (N_26077,N_24689,N_24989);
or U26078 (N_26078,N_25154,N_24045);
nand U26079 (N_26079,N_25094,N_24639);
nor U26080 (N_26080,N_25163,N_24619);
and U26081 (N_26081,N_24729,N_24940);
and U26082 (N_26082,N_24096,N_24749);
nor U26083 (N_26083,N_24024,N_24856);
and U26084 (N_26084,N_24722,N_24021);
xnor U26085 (N_26085,N_24890,N_24299);
or U26086 (N_26086,N_24630,N_24262);
nor U26087 (N_26087,N_24506,N_24774);
xor U26088 (N_26088,N_24805,N_24234);
nand U26089 (N_26089,N_24894,N_24540);
or U26090 (N_26090,N_24970,N_24210);
nand U26091 (N_26091,N_24660,N_24014);
nor U26092 (N_26092,N_24204,N_24114);
or U26093 (N_26093,N_24593,N_24683);
or U26094 (N_26094,N_24439,N_24978);
or U26095 (N_26095,N_24604,N_24741);
nand U26096 (N_26096,N_25194,N_24839);
and U26097 (N_26097,N_24492,N_24242);
xor U26098 (N_26098,N_25137,N_24363);
and U26099 (N_26099,N_24844,N_24551);
xnor U26100 (N_26100,N_24199,N_25055);
or U26101 (N_26101,N_24013,N_24298);
nor U26102 (N_26102,N_24044,N_24632);
nand U26103 (N_26103,N_24746,N_24637);
and U26104 (N_26104,N_24834,N_24582);
and U26105 (N_26105,N_24589,N_24462);
or U26106 (N_26106,N_25095,N_24881);
or U26107 (N_26107,N_24554,N_24697);
nand U26108 (N_26108,N_24641,N_25019);
nor U26109 (N_26109,N_24590,N_24648);
nor U26110 (N_26110,N_25042,N_24155);
and U26111 (N_26111,N_24535,N_24742);
xor U26112 (N_26112,N_25027,N_24951);
nand U26113 (N_26113,N_24007,N_25010);
xor U26114 (N_26114,N_24454,N_25171);
and U26115 (N_26115,N_24016,N_25169);
xnor U26116 (N_26116,N_24838,N_24350);
and U26117 (N_26117,N_25063,N_24648);
or U26118 (N_26118,N_24868,N_24158);
and U26119 (N_26119,N_24746,N_24248);
nand U26120 (N_26120,N_24718,N_24054);
and U26121 (N_26121,N_24595,N_24954);
nor U26122 (N_26122,N_25168,N_24398);
and U26123 (N_26123,N_24765,N_24700);
and U26124 (N_26124,N_24416,N_24972);
and U26125 (N_26125,N_24597,N_24566);
xnor U26126 (N_26126,N_24397,N_25126);
xor U26127 (N_26127,N_24559,N_24790);
or U26128 (N_26128,N_24926,N_24147);
nand U26129 (N_26129,N_24515,N_24155);
xor U26130 (N_26130,N_24084,N_24270);
and U26131 (N_26131,N_25167,N_24511);
nor U26132 (N_26132,N_24346,N_24349);
and U26133 (N_26133,N_24831,N_24164);
nor U26134 (N_26134,N_24274,N_25089);
or U26135 (N_26135,N_24402,N_24983);
xor U26136 (N_26136,N_24613,N_25027);
nand U26137 (N_26137,N_25136,N_24829);
xor U26138 (N_26138,N_24024,N_24902);
and U26139 (N_26139,N_24880,N_25059);
nand U26140 (N_26140,N_24836,N_24658);
and U26141 (N_26141,N_24516,N_24298);
nand U26142 (N_26142,N_24283,N_25175);
xnor U26143 (N_26143,N_24495,N_24791);
xor U26144 (N_26144,N_24711,N_24992);
xnor U26145 (N_26145,N_24405,N_24917);
nand U26146 (N_26146,N_24135,N_24982);
nor U26147 (N_26147,N_24040,N_24552);
nor U26148 (N_26148,N_24526,N_24823);
and U26149 (N_26149,N_24975,N_24771);
nor U26150 (N_26150,N_25166,N_24223);
xor U26151 (N_26151,N_24872,N_24600);
nand U26152 (N_26152,N_25198,N_24200);
nand U26153 (N_26153,N_24888,N_24616);
and U26154 (N_26154,N_25133,N_25008);
xor U26155 (N_26155,N_24692,N_24135);
xor U26156 (N_26156,N_24877,N_24331);
nand U26157 (N_26157,N_24485,N_24502);
xor U26158 (N_26158,N_25160,N_24677);
and U26159 (N_26159,N_24725,N_24355);
nand U26160 (N_26160,N_24506,N_24507);
xor U26161 (N_26161,N_24120,N_24339);
xnor U26162 (N_26162,N_25018,N_24316);
or U26163 (N_26163,N_24668,N_24968);
nor U26164 (N_26164,N_24887,N_24133);
or U26165 (N_26165,N_24610,N_24813);
and U26166 (N_26166,N_24659,N_24431);
or U26167 (N_26167,N_24282,N_24502);
nand U26168 (N_26168,N_24235,N_24152);
or U26169 (N_26169,N_24131,N_24622);
xor U26170 (N_26170,N_24804,N_24172);
and U26171 (N_26171,N_24500,N_25186);
and U26172 (N_26172,N_24402,N_24117);
and U26173 (N_26173,N_25020,N_25191);
xor U26174 (N_26174,N_24249,N_25154);
nor U26175 (N_26175,N_24088,N_24120);
or U26176 (N_26176,N_24277,N_24202);
nor U26177 (N_26177,N_25178,N_24347);
and U26178 (N_26178,N_25154,N_24265);
xnor U26179 (N_26179,N_24982,N_24338);
or U26180 (N_26180,N_24043,N_24847);
and U26181 (N_26181,N_24329,N_24599);
nand U26182 (N_26182,N_24920,N_24036);
nand U26183 (N_26183,N_24764,N_24425);
or U26184 (N_26184,N_24740,N_24723);
xnor U26185 (N_26185,N_24003,N_24313);
and U26186 (N_26186,N_24133,N_24166);
or U26187 (N_26187,N_24724,N_24094);
nor U26188 (N_26188,N_24299,N_24971);
or U26189 (N_26189,N_24386,N_24572);
and U26190 (N_26190,N_24052,N_24818);
and U26191 (N_26191,N_24497,N_25108);
or U26192 (N_26192,N_24279,N_24788);
nor U26193 (N_26193,N_24689,N_24183);
and U26194 (N_26194,N_24497,N_24112);
nand U26195 (N_26195,N_24945,N_24222);
nand U26196 (N_26196,N_24613,N_24867);
and U26197 (N_26197,N_25187,N_24969);
nand U26198 (N_26198,N_24759,N_24943);
nor U26199 (N_26199,N_24313,N_24396);
or U26200 (N_26200,N_24170,N_24195);
nor U26201 (N_26201,N_24318,N_25168);
nor U26202 (N_26202,N_24363,N_24730);
xnor U26203 (N_26203,N_25056,N_24854);
nor U26204 (N_26204,N_24882,N_24736);
xnor U26205 (N_26205,N_24987,N_24786);
and U26206 (N_26206,N_25155,N_25022);
or U26207 (N_26207,N_24754,N_24662);
nor U26208 (N_26208,N_24866,N_24801);
nand U26209 (N_26209,N_24857,N_24520);
and U26210 (N_26210,N_24656,N_24277);
or U26211 (N_26211,N_24629,N_24253);
nor U26212 (N_26212,N_24044,N_25009);
nand U26213 (N_26213,N_24253,N_24082);
nand U26214 (N_26214,N_24138,N_24417);
xnor U26215 (N_26215,N_24964,N_25103);
and U26216 (N_26216,N_24486,N_24606);
xor U26217 (N_26217,N_24202,N_25182);
or U26218 (N_26218,N_24560,N_24163);
and U26219 (N_26219,N_25174,N_24731);
nand U26220 (N_26220,N_25189,N_24796);
nand U26221 (N_26221,N_24550,N_24011);
nor U26222 (N_26222,N_24422,N_24751);
and U26223 (N_26223,N_24068,N_24806);
xnor U26224 (N_26224,N_25182,N_25049);
and U26225 (N_26225,N_24268,N_24109);
xnor U26226 (N_26226,N_24822,N_24841);
nor U26227 (N_26227,N_24983,N_24353);
xnor U26228 (N_26228,N_24012,N_25116);
nor U26229 (N_26229,N_24255,N_25102);
nand U26230 (N_26230,N_24635,N_24127);
nor U26231 (N_26231,N_25023,N_24583);
nand U26232 (N_26232,N_25060,N_24388);
xnor U26233 (N_26233,N_24769,N_24757);
and U26234 (N_26234,N_24329,N_24505);
or U26235 (N_26235,N_25070,N_25192);
nand U26236 (N_26236,N_24695,N_24843);
or U26237 (N_26237,N_24532,N_24564);
xor U26238 (N_26238,N_24648,N_24135);
nand U26239 (N_26239,N_25022,N_24700);
and U26240 (N_26240,N_25079,N_24339);
or U26241 (N_26241,N_24632,N_24997);
xor U26242 (N_26242,N_24507,N_24970);
nor U26243 (N_26243,N_24016,N_24840);
nand U26244 (N_26244,N_24016,N_24353);
nand U26245 (N_26245,N_24920,N_24310);
xnor U26246 (N_26246,N_24608,N_24987);
nand U26247 (N_26247,N_24138,N_24365);
xnor U26248 (N_26248,N_24024,N_24930);
or U26249 (N_26249,N_24358,N_25089);
and U26250 (N_26250,N_24437,N_24812);
nor U26251 (N_26251,N_24696,N_24767);
and U26252 (N_26252,N_24252,N_24036);
nand U26253 (N_26253,N_24470,N_24041);
xnor U26254 (N_26254,N_24989,N_24602);
xnor U26255 (N_26255,N_24753,N_24301);
xor U26256 (N_26256,N_25053,N_24121);
xnor U26257 (N_26257,N_24116,N_24785);
or U26258 (N_26258,N_24387,N_24248);
nand U26259 (N_26259,N_24295,N_24657);
xor U26260 (N_26260,N_24076,N_24573);
or U26261 (N_26261,N_24839,N_24986);
nand U26262 (N_26262,N_24755,N_24012);
and U26263 (N_26263,N_24330,N_24999);
xnor U26264 (N_26264,N_24184,N_24416);
nor U26265 (N_26265,N_24971,N_24446);
nor U26266 (N_26266,N_24742,N_24769);
nor U26267 (N_26267,N_24967,N_24081);
or U26268 (N_26268,N_24716,N_24102);
nand U26269 (N_26269,N_25132,N_24077);
xor U26270 (N_26270,N_24113,N_24983);
nor U26271 (N_26271,N_24744,N_24662);
xor U26272 (N_26272,N_24876,N_24256);
or U26273 (N_26273,N_25027,N_24373);
and U26274 (N_26274,N_24184,N_24649);
and U26275 (N_26275,N_24816,N_24082);
and U26276 (N_26276,N_24594,N_24702);
or U26277 (N_26277,N_24281,N_24074);
xor U26278 (N_26278,N_24016,N_24549);
xor U26279 (N_26279,N_24964,N_24233);
and U26280 (N_26280,N_24661,N_24461);
nand U26281 (N_26281,N_24247,N_24119);
nor U26282 (N_26282,N_25133,N_25184);
or U26283 (N_26283,N_24233,N_24899);
xor U26284 (N_26284,N_24348,N_24893);
or U26285 (N_26285,N_24597,N_25045);
and U26286 (N_26286,N_24568,N_24252);
nand U26287 (N_26287,N_24114,N_24382);
nand U26288 (N_26288,N_24195,N_24596);
nor U26289 (N_26289,N_24901,N_24423);
xnor U26290 (N_26290,N_25103,N_24434);
nor U26291 (N_26291,N_25166,N_24314);
nand U26292 (N_26292,N_24985,N_24587);
nor U26293 (N_26293,N_24176,N_24719);
xnor U26294 (N_26294,N_24578,N_24423);
and U26295 (N_26295,N_25090,N_24331);
nand U26296 (N_26296,N_24808,N_24928);
xor U26297 (N_26297,N_24384,N_24804);
nand U26298 (N_26298,N_24150,N_24542);
or U26299 (N_26299,N_24498,N_24158);
nor U26300 (N_26300,N_24014,N_24425);
and U26301 (N_26301,N_24794,N_24343);
and U26302 (N_26302,N_24634,N_24260);
and U26303 (N_26303,N_25196,N_24601);
and U26304 (N_26304,N_24896,N_24182);
and U26305 (N_26305,N_24356,N_25024);
nor U26306 (N_26306,N_25085,N_24179);
nor U26307 (N_26307,N_24013,N_24431);
nor U26308 (N_26308,N_24447,N_24376);
or U26309 (N_26309,N_24813,N_24984);
xor U26310 (N_26310,N_25063,N_24303);
nor U26311 (N_26311,N_24829,N_24692);
xor U26312 (N_26312,N_24659,N_24164);
nor U26313 (N_26313,N_24314,N_24498);
nand U26314 (N_26314,N_24815,N_25152);
nor U26315 (N_26315,N_24353,N_24257);
nand U26316 (N_26316,N_24904,N_24378);
and U26317 (N_26317,N_24762,N_24894);
nor U26318 (N_26318,N_24207,N_24237);
or U26319 (N_26319,N_25134,N_24925);
nor U26320 (N_26320,N_25188,N_24654);
and U26321 (N_26321,N_24785,N_24685);
or U26322 (N_26322,N_24957,N_24309);
or U26323 (N_26323,N_24374,N_25157);
nor U26324 (N_26324,N_25027,N_24379);
nand U26325 (N_26325,N_24799,N_24596);
or U26326 (N_26326,N_24394,N_24729);
or U26327 (N_26327,N_24930,N_24834);
or U26328 (N_26328,N_24968,N_25136);
xnor U26329 (N_26329,N_24200,N_24868);
xor U26330 (N_26330,N_24369,N_24832);
or U26331 (N_26331,N_25010,N_24482);
nand U26332 (N_26332,N_24687,N_24548);
xor U26333 (N_26333,N_24551,N_24126);
xnor U26334 (N_26334,N_24048,N_24326);
or U26335 (N_26335,N_24865,N_24138);
or U26336 (N_26336,N_24811,N_24224);
and U26337 (N_26337,N_24462,N_24581);
nand U26338 (N_26338,N_24213,N_25123);
or U26339 (N_26339,N_24948,N_24154);
or U26340 (N_26340,N_24937,N_24959);
nand U26341 (N_26341,N_24483,N_24205);
or U26342 (N_26342,N_24979,N_24103);
xor U26343 (N_26343,N_25082,N_24251);
xor U26344 (N_26344,N_24666,N_24617);
and U26345 (N_26345,N_24895,N_24387);
and U26346 (N_26346,N_24830,N_24500);
xor U26347 (N_26347,N_24790,N_24035);
xor U26348 (N_26348,N_24734,N_24028);
xnor U26349 (N_26349,N_24010,N_25031);
or U26350 (N_26350,N_24494,N_24980);
nand U26351 (N_26351,N_25097,N_24468);
nand U26352 (N_26352,N_24129,N_25031);
nor U26353 (N_26353,N_24068,N_24287);
and U26354 (N_26354,N_24337,N_24660);
or U26355 (N_26355,N_24932,N_24433);
xnor U26356 (N_26356,N_25159,N_24670);
nor U26357 (N_26357,N_24885,N_24136);
xor U26358 (N_26358,N_24395,N_24542);
xor U26359 (N_26359,N_24668,N_24573);
xnor U26360 (N_26360,N_25075,N_25176);
and U26361 (N_26361,N_24022,N_24286);
nor U26362 (N_26362,N_24650,N_24507);
nand U26363 (N_26363,N_24531,N_24137);
or U26364 (N_26364,N_24631,N_24240);
or U26365 (N_26365,N_24402,N_24981);
xnor U26366 (N_26366,N_24472,N_24754);
or U26367 (N_26367,N_24262,N_24575);
xor U26368 (N_26368,N_24336,N_24820);
nand U26369 (N_26369,N_24045,N_24580);
and U26370 (N_26370,N_24690,N_25184);
or U26371 (N_26371,N_24744,N_24867);
xor U26372 (N_26372,N_24224,N_25164);
or U26373 (N_26373,N_24515,N_24778);
or U26374 (N_26374,N_24055,N_24722);
xor U26375 (N_26375,N_24519,N_24016);
and U26376 (N_26376,N_24560,N_24645);
nor U26377 (N_26377,N_24841,N_24557);
and U26378 (N_26378,N_24147,N_24788);
nand U26379 (N_26379,N_24288,N_24187);
and U26380 (N_26380,N_24836,N_24410);
xnor U26381 (N_26381,N_24084,N_24790);
or U26382 (N_26382,N_24882,N_24903);
or U26383 (N_26383,N_25038,N_25049);
xor U26384 (N_26384,N_24827,N_24553);
or U26385 (N_26385,N_24064,N_24381);
or U26386 (N_26386,N_24948,N_24613);
xor U26387 (N_26387,N_24812,N_24321);
nand U26388 (N_26388,N_25140,N_24657);
nand U26389 (N_26389,N_25194,N_24028);
and U26390 (N_26390,N_25096,N_24145);
nor U26391 (N_26391,N_25083,N_24860);
xnor U26392 (N_26392,N_24297,N_24327);
xor U26393 (N_26393,N_24385,N_24482);
xnor U26394 (N_26394,N_24792,N_25198);
nand U26395 (N_26395,N_24708,N_24837);
xor U26396 (N_26396,N_24017,N_24063);
or U26397 (N_26397,N_24528,N_24422);
xnor U26398 (N_26398,N_24992,N_24152);
and U26399 (N_26399,N_24136,N_25111);
nand U26400 (N_26400,N_25376,N_25602);
nor U26401 (N_26401,N_25554,N_25393);
nor U26402 (N_26402,N_25616,N_25477);
nor U26403 (N_26403,N_25652,N_26368);
xnor U26404 (N_26404,N_25954,N_25441);
nor U26405 (N_26405,N_25632,N_25360);
xor U26406 (N_26406,N_25714,N_25359);
or U26407 (N_26407,N_26021,N_25298);
nand U26408 (N_26408,N_26351,N_25678);
or U26409 (N_26409,N_25504,N_25494);
xnor U26410 (N_26410,N_26081,N_25532);
nor U26411 (N_26411,N_26288,N_25621);
nor U26412 (N_26412,N_25261,N_25580);
nand U26413 (N_26413,N_25709,N_25603);
or U26414 (N_26414,N_25465,N_25863);
nor U26415 (N_26415,N_26172,N_25710);
nand U26416 (N_26416,N_26255,N_25481);
nand U26417 (N_26417,N_25623,N_26382);
and U26418 (N_26418,N_25620,N_25776);
or U26419 (N_26419,N_25218,N_25242);
or U26420 (N_26420,N_25949,N_25646);
nand U26421 (N_26421,N_25633,N_25878);
and U26422 (N_26422,N_25936,N_25392);
nor U26423 (N_26423,N_25841,N_25537);
nor U26424 (N_26424,N_25593,N_25794);
and U26425 (N_26425,N_25337,N_25831);
nor U26426 (N_26426,N_25557,N_25752);
xor U26427 (N_26427,N_25284,N_25358);
and U26428 (N_26428,N_25422,N_25350);
nand U26429 (N_26429,N_25318,N_25340);
and U26430 (N_26430,N_25275,N_25899);
xnor U26431 (N_26431,N_25904,N_26377);
and U26432 (N_26432,N_25201,N_25812);
nand U26433 (N_26433,N_25470,N_26293);
nor U26434 (N_26434,N_26367,N_25976);
xor U26435 (N_26435,N_26389,N_25849);
nor U26436 (N_26436,N_26101,N_25496);
or U26437 (N_26437,N_26272,N_26245);
nor U26438 (N_26438,N_25706,N_26342);
xnor U26439 (N_26439,N_25757,N_25250);
and U26440 (N_26440,N_25444,N_25323);
nor U26441 (N_26441,N_26123,N_25892);
nand U26442 (N_26442,N_25845,N_25839);
nor U26443 (N_26443,N_25826,N_25973);
nor U26444 (N_26444,N_25853,N_25395);
xnor U26445 (N_26445,N_25263,N_25805);
and U26446 (N_26446,N_25735,N_26158);
xnor U26447 (N_26447,N_26063,N_25338);
and U26448 (N_26448,N_25804,N_26004);
xnor U26449 (N_26449,N_25549,N_25431);
nor U26450 (N_26450,N_25448,N_26070);
xnor U26451 (N_26451,N_25208,N_26269);
xor U26452 (N_26452,N_26187,N_25858);
xor U26453 (N_26453,N_25488,N_26059);
nor U26454 (N_26454,N_25993,N_26332);
or U26455 (N_26455,N_26373,N_25851);
and U26456 (N_26456,N_25894,N_25437);
xnor U26457 (N_26457,N_25344,N_25627);
or U26458 (N_26458,N_25665,N_26064);
xor U26459 (N_26459,N_25267,N_25762);
and U26460 (N_26460,N_25558,N_25378);
nand U26461 (N_26461,N_26054,N_25864);
nor U26462 (N_26462,N_26282,N_25923);
and U26463 (N_26463,N_26216,N_25372);
nand U26464 (N_26464,N_26111,N_25988);
nor U26465 (N_26465,N_25875,N_25562);
or U26466 (N_26466,N_25870,N_25888);
or U26467 (N_26467,N_25950,N_25205);
nand U26468 (N_26468,N_25925,N_25679);
and U26469 (N_26469,N_25837,N_26166);
xor U26470 (N_26470,N_26058,N_25290);
or U26471 (N_26471,N_25262,N_26193);
and U26472 (N_26472,N_25381,N_25962);
xnor U26473 (N_26473,N_26364,N_25765);
xnor U26474 (N_26474,N_25650,N_26203);
and U26475 (N_26475,N_25671,N_26195);
and U26476 (N_26476,N_25749,N_25584);
or U26477 (N_26477,N_26122,N_26258);
or U26478 (N_26478,N_25386,N_25803);
nand U26479 (N_26479,N_25717,N_26378);
or U26480 (N_26480,N_26285,N_25916);
nand U26481 (N_26481,N_26083,N_26208);
and U26482 (N_26482,N_26205,N_26197);
nand U26483 (N_26483,N_26394,N_25824);
nor U26484 (N_26484,N_25642,N_25215);
xnor U26485 (N_26485,N_25969,N_26279);
and U26486 (N_26486,N_26042,N_25777);
nor U26487 (N_26487,N_25618,N_25221);
nand U26488 (N_26488,N_25978,N_26225);
and U26489 (N_26489,N_25756,N_26136);
or U26490 (N_26490,N_25860,N_25301);
or U26491 (N_26491,N_26170,N_26214);
nor U26492 (N_26492,N_25921,N_25458);
or U26493 (N_26493,N_25544,N_26086);
or U26494 (N_26494,N_25834,N_26008);
nand U26495 (N_26495,N_25963,N_25946);
nand U26496 (N_26496,N_26137,N_26322);
nand U26497 (N_26497,N_25428,N_25825);
nand U26498 (N_26498,N_25495,N_26217);
nor U26499 (N_26499,N_25595,N_25576);
xor U26500 (N_26500,N_25232,N_25235);
and U26501 (N_26501,N_26385,N_25429);
and U26502 (N_26502,N_25877,N_25833);
nand U26503 (N_26503,N_25760,N_26333);
xor U26504 (N_26504,N_25772,N_26221);
and U26505 (N_26505,N_25604,N_26125);
and U26506 (N_26506,N_25855,N_25506);
nor U26507 (N_26507,N_26301,N_25952);
and U26508 (N_26508,N_25503,N_25572);
or U26509 (N_26509,N_25659,N_26192);
nor U26510 (N_26510,N_26189,N_26151);
or U26511 (N_26511,N_25673,N_25666);
nor U26512 (N_26512,N_26200,N_26387);
and U26513 (N_26513,N_25471,N_25599);
nand U26514 (N_26514,N_25516,N_25510);
nand U26515 (N_26515,N_26253,N_25586);
nand U26516 (N_26516,N_25613,N_25405);
nor U26517 (N_26517,N_25223,N_25548);
nand U26518 (N_26518,N_26390,N_25754);
or U26519 (N_26519,N_26283,N_25647);
nand U26520 (N_26520,N_25414,N_26060);
xor U26521 (N_26521,N_25887,N_25725);
xnor U26522 (N_26522,N_25367,N_26291);
and U26523 (N_26523,N_26061,N_26011);
and U26524 (N_26524,N_25260,N_26198);
or U26525 (N_26525,N_25243,N_25382);
or U26526 (N_26526,N_25575,N_25332);
or U26527 (N_26527,N_25225,N_26260);
or U26528 (N_26528,N_25748,N_26132);
xor U26529 (N_26529,N_25288,N_26399);
nor U26530 (N_26530,N_25913,N_25662);
nor U26531 (N_26531,N_25715,N_25891);
and U26532 (N_26532,N_25509,N_25230);
xor U26533 (N_26533,N_25823,N_26355);
nor U26534 (N_26534,N_26268,N_25838);
xnor U26535 (N_26535,N_26133,N_25202);
and U26536 (N_26536,N_25655,N_25700);
nand U26537 (N_26537,N_25570,N_25564);
or U26538 (N_26538,N_25307,N_25396);
nand U26539 (N_26539,N_25964,N_25265);
xnor U26540 (N_26540,N_25846,N_25308);
and U26541 (N_26541,N_25545,N_26048);
nor U26542 (N_26542,N_25327,N_26139);
nand U26543 (N_26543,N_25240,N_26173);
or U26544 (N_26544,N_25412,N_26196);
nand U26545 (N_26545,N_25746,N_26178);
nor U26546 (N_26546,N_25417,N_25380);
nand U26547 (N_26547,N_26243,N_26085);
and U26548 (N_26548,N_25722,N_26311);
xnor U26549 (N_26549,N_26160,N_25445);
nor U26550 (N_26550,N_26091,N_25986);
or U26551 (N_26551,N_25727,N_25568);
and U26552 (N_26552,N_25355,N_25733);
nand U26553 (N_26553,N_26068,N_26033);
nor U26554 (N_26554,N_25786,N_25842);
and U26555 (N_26555,N_25353,N_26384);
xnor U26556 (N_26556,N_25938,N_26300);
nand U26557 (N_26557,N_26116,N_26357);
nor U26558 (N_26558,N_25672,N_26179);
and U26559 (N_26559,N_26380,N_25500);
and U26560 (N_26560,N_25867,N_25948);
or U26561 (N_26561,N_26396,N_25712);
or U26562 (N_26562,N_25419,N_25487);
or U26563 (N_26563,N_26098,N_25291);
or U26564 (N_26564,N_26002,N_25497);
or U26565 (N_26565,N_26248,N_26128);
and U26566 (N_26566,N_26340,N_25645);
xor U26567 (N_26567,N_25657,N_25912);
nand U26568 (N_26568,N_25987,N_25363);
or U26569 (N_26569,N_25521,N_25279);
nand U26570 (N_26570,N_25896,N_26249);
or U26571 (N_26571,N_25493,N_25984);
xor U26572 (N_26572,N_25769,N_25957);
nor U26573 (N_26573,N_25526,N_25609);
and U26574 (N_26574,N_26035,N_25744);
and U26575 (N_26575,N_26257,N_26287);
or U26576 (N_26576,N_25394,N_25383);
and U26577 (N_26577,N_25224,N_25587);
nand U26578 (N_26578,N_25583,N_25880);
or U26579 (N_26579,N_25995,N_26330);
nand U26580 (N_26580,N_26171,N_25955);
xnor U26581 (N_26581,N_26107,N_26202);
nor U26582 (N_26582,N_26090,N_25681);
or U26583 (N_26583,N_25610,N_25607);
nand U26584 (N_26584,N_25767,N_26310);
and U26585 (N_26585,N_25897,N_25443);
nor U26586 (N_26586,N_25654,N_26262);
or U26587 (N_26587,N_25430,N_26201);
nor U26588 (N_26588,N_26052,N_25553);
and U26589 (N_26589,N_25226,N_25336);
nand U26590 (N_26590,N_25764,N_26356);
nand U26591 (N_26591,N_25810,N_26360);
nand U26592 (N_26592,N_26317,N_25835);
xor U26593 (N_26593,N_25909,N_25552);
and U26594 (N_26594,N_26102,N_26155);
xnor U26595 (N_26595,N_26199,N_25670);
xor U26596 (N_26596,N_26038,N_25425);
nand U26597 (N_26597,N_25569,N_25528);
nor U26598 (N_26598,N_25361,N_26273);
or U26599 (N_26599,N_26206,N_25438);
nor U26600 (N_26600,N_25668,N_26324);
xor U26601 (N_26601,N_25677,N_25342);
nand U26602 (N_26602,N_26302,N_26131);
and U26603 (N_26603,N_25859,N_26219);
nand U26604 (N_26604,N_25499,N_25740);
nor U26605 (N_26605,N_25844,N_25763);
and U26606 (N_26606,N_25815,N_25424);
nor U26607 (N_26607,N_26082,N_26162);
or U26608 (N_26608,N_26354,N_25876);
and U26609 (N_26609,N_25309,N_25693);
or U26610 (N_26610,N_26120,N_26210);
nor U26611 (N_26611,N_25641,N_25403);
xnor U26612 (N_26612,N_25703,N_25771);
nand U26613 (N_26613,N_26065,N_26218);
or U26614 (N_26614,N_25782,N_25498);
xnor U26615 (N_26615,N_26144,N_25959);
and U26616 (N_26616,N_25734,N_25565);
xor U26617 (N_26617,N_25994,N_25287);
nand U26618 (N_26618,N_25902,N_26175);
and U26619 (N_26619,N_25966,N_26298);
nor U26620 (N_26620,N_26365,N_26150);
or U26621 (N_26621,N_25289,N_25321);
and U26622 (N_26622,N_25302,N_25517);
xnor U26623 (N_26623,N_26176,N_26154);
xor U26624 (N_26624,N_26013,N_26229);
or U26625 (N_26625,N_25639,N_26174);
or U26626 (N_26626,N_25371,N_25648);
and U26627 (N_26627,N_25408,N_25625);
xnor U26628 (N_26628,N_26049,N_25300);
nor U26629 (N_26629,N_25379,N_26278);
nand U26630 (N_26630,N_25295,N_25550);
nand U26631 (N_26631,N_25566,N_26321);
nand U26632 (N_26632,N_25972,N_25981);
nor U26633 (N_26633,N_26118,N_26295);
nand U26634 (N_26634,N_25320,N_25316);
or U26635 (N_26635,N_25945,N_26006);
nand U26636 (N_26636,N_25432,N_25911);
nor U26637 (N_26637,N_26207,N_25898);
xnor U26638 (N_26638,N_26010,N_25614);
and U26639 (N_26639,N_25254,N_25691);
and U26640 (N_26640,N_25389,N_25463);
xor U26641 (N_26641,N_25871,N_25390);
or U26642 (N_26642,N_25426,N_25501);
and U26643 (N_26643,N_26169,N_26397);
nor U26644 (N_26644,N_26126,N_26240);
nor U26645 (N_26645,N_25890,N_26350);
and U26646 (N_26646,N_26050,N_26388);
nand U26647 (N_26647,N_26029,N_25720);
nand U26648 (N_26648,N_25385,N_25731);
or U26649 (N_26649,N_26246,N_26129);
nor U26650 (N_26650,N_25418,N_25440);
and U26651 (N_26651,N_26164,N_25792);
nand U26652 (N_26652,N_26096,N_25663);
xor U26653 (N_26653,N_25507,N_25882);
nand U26654 (N_26654,N_25236,N_25556);
nor U26655 (N_26655,N_25827,N_26093);
nand U26656 (N_26656,N_26275,N_25785);
xor U26657 (N_26657,N_25559,N_25585);
and U26658 (N_26658,N_25352,N_25365);
and U26659 (N_26659,N_25539,N_25920);
nand U26660 (N_26660,N_25612,N_25253);
nor U26661 (N_26661,N_26184,N_25271);
nor U26662 (N_26662,N_25811,N_26352);
or U26663 (N_26663,N_25282,N_25377);
nor U26664 (N_26664,N_26109,N_25272);
and U26665 (N_26665,N_25578,N_25798);
and U26666 (N_26666,N_26336,N_26308);
nor U26667 (N_26667,N_26159,N_26034);
and U26668 (N_26668,N_25206,N_25857);
or U26669 (N_26669,N_25992,N_26392);
or U26670 (N_26670,N_25968,N_25335);
nor U26671 (N_26671,N_25312,N_25530);
nand U26672 (N_26672,N_26239,N_26023);
xnor U26673 (N_26673,N_25281,N_26067);
xor U26674 (N_26674,N_25695,N_26265);
or U26675 (N_26675,N_25442,N_25346);
xor U26676 (N_26676,N_25998,N_25914);
nor U26677 (N_26677,N_25436,N_25928);
and U26678 (N_26678,N_25906,N_26250);
nor U26679 (N_26679,N_25415,N_25401);
or U26680 (N_26680,N_25357,N_26233);
nor U26681 (N_26681,N_25364,N_25941);
or U26682 (N_26682,N_25822,N_25758);
xnor U26683 (N_26683,N_26104,N_26080);
nand U26684 (N_26684,N_25630,N_25277);
nor U26685 (N_26685,N_26000,N_25929);
nor U26686 (N_26686,N_25214,N_25582);
xnor U26687 (N_26687,N_25664,N_25333);
or U26688 (N_26688,N_26106,N_25283);
nor U26689 (N_26689,N_25362,N_26167);
xor U26690 (N_26690,N_26103,N_25908);
and U26691 (N_26691,N_25667,N_26231);
nand U26692 (N_26692,N_25563,N_25791);
xnor U26693 (N_26693,N_26237,N_25699);
nand U26694 (N_26694,N_25370,N_26088);
nor U26695 (N_26695,N_25435,N_26186);
xnor U26696 (N_26696,N_26028,N_25369);
and U26697 (N_26697,N_25345,N_25656);
xnor U26698 (N_26698,N_25761,N_25339);
xor U26699 (N_26699,N_25200,N_25674);
or U26700 (N_26700,N_25644,N_25601);
or U26701 (N_26701,N_25325,N_26274);
xnor U26702 (N_26702,N_26306,N_26121);
nand U26703 (N_26703,N_26062,N_25464);
nor U26704 (N_26704,N_26353,N_25522);
or U26705 (N_26705,N_25391,N_25527);
xnor U26706 (N_26706,N_25806,N_25286);
or U26707 (N_26707,N_26043,N_26320);
and U26708 (N_26708,N_25915,N_26134);
xnor U26709 (N_26709,N_25533,N_25523);
nand U26710 (N_26710,N_25518,N_25457);
nand U26711 (N_26711,N_26358,N_25455);
or U26712 (N_26712,N_25466,N_25683);
or U26713 (N_26713,N_26053,N_25297);
xor U26714 (N_26714,N_26057,N_25347);
or U26715 (N_26715,N_25799,N_25918);
or U26716 (N_26716,N_25797,N_26039);
and U26717 (N_26717,N_25937,N_25713);
nand U26718 (N_26718,N_25807,N_26071);
nor U26719 (N_26719,N_25989,N_25483);
nand U26720 (N_26720,N_26228,N_25315);
and U26721 (N_26721,N_26267,N_25474);
nand U26722 (N_26722,N_25975,N_25547);
nor U26723 (N_26723,N_26323,N_25728);
xor U26724 (N_26724,N_25747,N_26119);
and U26725 (N_26725,N_26095,N_25447);
nor U26726 (N_26726,N_26326,N_25433);
nor U26727 (N_26727,N_26190,N_25883);
and U26728 (N_26728,N_25942,N_25680);
or U26729 (N_26729,N_26152,N_25306);
nand U26730 (N_26730,N_25723,N_25828);
nor U26731 (N_26731,N_25524,N_25567);
and U26732 (N_26732,N_26303,N_25268);
or U26733 (N_26733,N_26227,N_26180);
nand U26734 (N_26734,N_25446,N_25985);
xnor U26735 (N_26735,N_26281,N_25856);
nor U26736 (N_26736,N_25231,N_25965);
and U26737 (N_26737,N_26215,N_25884);
nand U26738 (N_26738,N_25751,N_26232);
and U26739 (N_26739,N_26305,N_25800);
nor U26740 (N_26740,N_26224,N_25531);
xnor U26741 (N_26741,N_25203,N_26191);
and U26742 (N_26742,N_25220,N_26117);
and U26743 (N_26743,N_25227,N_26020);
and U26744 (N_26744,N_25900,N_25449);
nand U26745 (N_26745,N_25490,N_26108);
nand U26746 (N_26746,N_25745,N_26369);
and U26747 (N_26747,N_25637,N_26127);
or U26748 (N_26748,N_26211,N_26325);
or U26749 (N_26749,N_25788,N_25692);
and U26750 (N_26750,N_26209,N_25233);
and U26751 (N_26751,N_25388,N_26114);
nor U26752 (N_26752,N_26014,N_25893);
xnor U26753 (N_26753,N_25492,N_26296);
xnor U26754 (N_26754,N_25249,N_26348);
nor U26755 (N_26755,N_25421,N_26316);
nor U26756 (N_26756,N_25830,N_25829);
and U26757 (N_26757,N_25718,N_25775);
nand U26758 (N_26758,N_26007,N_25551);
or U26759 (N_26759,N_26012,N_25927);
and U26760 (N_26760,N_25351,N_26236);
xnor U26761 (N_26761,N_25980,N_25624);
nor U26762 (N_26762,N_26056,N_26076);
xnor U26763 (N_26763,N_25635,N_25311);
and U26764 (N_26764,N_25768,N_25467);
and U26765 (N_26765,N_25273,N_25328);
xor U26766 (N_26766,N_25590,N_25759);
and U26767 (N_26767,N_25374,N_25259);
xor U26768 (N_26768,N_26100,N_26110);
xnor U26769 (N_26769,N_25809,N_26318);
xor U26770 (N_26770,N_26094,N_25237);
nor U26771 (N_26771,N_25475,N_26188);
or U26772 (N_26772,N_25598,N_25636);
nor U26773 (N_26773,N_26266,N_25879);
or U26774 (N_26774,N_25750,N_26040);
nor U26775 (N_26775,N_25519,N_26078);
and U26776 (N_26776,N_25373,N_25462);
xor U26777 (N_26777,N_25411,N_25708);
and U26778 (N_26778,N_26194,N_26147);
or U26779 (N_26779,N_25472,N_26280);
xor U26780 (N_26780,N_25238,N_26124);
nor U26781 (N_26781,N_25903,N_25579);
xnor U26782 (N_26782,N_25862,N_25732);
and U26783 (N_26783,N_25515,N_25869);
nor U26784 (N_26784,N_25698,N_25951);
and U26785 (N_26785,N_26112,N_25400);
or U26786 (N_26786,N_25406,N_26286);
nand U26787 (N_26787,N_26181,N_26341);
xnor U26788 (N_26788,N_26045,N_25269);
nand U26789 (N_26789,N_25592,N_25622);
or U26790 (N_26790,N_26157,N_26372);
nor U26791 (N_26791,N_25217,N_26223);
and U26792 (N_26792,N_25881,N_26335);
and U26793 (N_26793,N_26289,N_25931);
nor U26794 (N_26794,N_25591,N_26140);
and U26795 (N_26795,N_25409,N_25330);
and U26796 (N_26796,N_26230,N_25478);
nor U26797 (N_26797,N_26030,N_25485);
nand U26798 (N_26798,N_26182,N_26032);
nand U26799 (N_26799,N_25276,N_26115);
and U26800 (N_26800,N_25280,N_25264);
or U26801 (N_26801,N_25460,N_25454);
nand U26802 (N_26802,N_25778,N_26163);
nand U26803 (N_26803,N_25971,N_26242);
xor U26804 (N_26804,N_25600,N_26251);
nor U26805 (N_26805,N_25917,N_25534);
xor U26806 (N_26806,N_26073,N_25305);
nand U26807 (N_26807,N_25482,N_25402);
and U26808 (N_26808,N_25239,N_25529);
xnor U26809 (N_26809,N_25737,N_25983);
nand U26810 (N_26810,N_25682,N_25687);
nand U26811 (N_26811,N_25322,N_25716);
nand U26812 (N_26812,N_25427,N_25560);
and U26813 (N_26813,N_25638,N_25817);
nand U26814 (N_26814,N_26222,N_26046);
nor U26815 (N_26815,N_25514,N_26292);
nand U26816 (N_26816,N_26277,N_25541);
nor U26817 (N_26817,N_26376,N_26024);
and U26818 (N_26818,N_25719,N_25991);
or U26819 (N_26819,N_25940,N_26141);
nand U26820 (N_26820,N_25407,N_25901);
or U26821 (N_26821,N_25802,N_25658);
and U26822 (N_26822,N_25990,N_26226);
nand U26823 (N_26823,N_26135,N_25707);
nand U26824 (N_26824,N_25615,N_26247);
nand U26825 (N_26825,N_25821,N_25468);
and U26826 (N_26826,N_25690,N_25736);
nor U26827 (N_26827,N_25953,N_25354);
nand U26828 (N_26828,N_26363,N_25423);
and U26829 (N_26829,N_25606,N_26148);
and U26830 (N_26830,N_25619,N_25329);
nand U26831 (N_26831,N_26386,N_25491);
or U26832 (N_26832,N_25781,N_25384);
and U26833 (N_26833,N_26204,N_25452);
nand U26834 (N_26834,N_26374,N_25854);
nor U26835 (N_26835,N_26009,N_25605);
nor U26836 (N_26836,N_25872,N_25451);
or U26837 (N_26837,N_26312,N_25935);
xnor U26838 (N_26838,N_26313,N_25244);
nand U26839 (N_26839,N_25790,N_25933);
nand U26840 (N_26840,N_26074,N_25304);
nor U26841 (N_26841,N_25484,N_25661);
or U26842 (N_26842,N_25944,N_25251);
and U26843 (N_26843,N_25922,N_25278);
nor U26844 (N_26844,N_25868,N_25813);
xnor U26845 (N_26845,N_26344,N_26375);
xnor U26846 (N_26846,N_25476,N_25697);
and U26847 (N_26847,N_26361,N_25439);
xnor U26848 (N_26848,N_25513,N_26270);
nand U26849 (N_26849,N_25368,N_26213);
or U26850 (N_26850,N_25577,N_26016);
and U26851 (N_26851,N_26212,N_25511);
nor U26852 (N_26852,N_25207,N_25865);
or U26853 (N_26853,N_25729,N_25816);
or U26854 (N_26854,N_25686,N_25974);
nor U26855 (N_26855,N_26347,N_25970);
xnor U26856 (N_26856,N_26327,N_26328);
and U26857 (N_26857,N_25960,N_26234);
nand U26858 (N_26858,N_25486,N_25588);
nand U26859 (N_26859,N_25404,N_26331);
nor U26860 (N_26860,N_26001,N_26339);
or U26861 (N_26861,N_26349,N_25314);
nand U26862 (N_26862,N_25934,N_25705);
and U26863 (N_26863,N_25398,N_25787);
and U26864 (N_26864,N_25505,N_25555);
or U26865 (N_26865,N_26290,N_25753);
nand U26866 (N_26866,N_25310,N_25581);
and U26867 (N_26867,N_25543,N_26003);
or U26868 (N_26868,N_26299,N_26105);
nor U26869 (N_26869,N_26022,N_25343);
or U26870 (N_26870,N_26142,N_25689);
nand U26871 (N_26871,N_25926,N_25649);
nand U26872 (N_26872,N_25416,N_25459);
nor U26873 (N_26873,N_26359,N_25397);
and U26874 (N_26874,N_25296,N_25818);
or U26875 (N_26875,N_25956,N_25245);
nor U26876 (N_26876,N_25589,N_26362);
nand U26877 (N_26877,N_26264,N_26084);
and U26878 (N_26878,N_25349,N_26113);
xnor U26879 (N_26879,N_26026,N_25608);
or U26880 (N_26880,N_25410,N_26047);
and U26881 (N_26881,N_25808,N_25596);
xor U26882 (N_26882,N_25675,N_25341);
or U26883 (N_26883,N_25246,N_25561);
nor U26884 (N_26884,N_25780,N_26315);
or U26885 (N_26885,N_25525,N_25209);
or U26886 (N_26886,N_26244,N_25299);
or U26887 (N_26887,N_25469,N_26075);
nor U26888 (N_26888,N_26055,N_25536);
nor U26889 (N_26889,N_26370,N_25979);
nand U26890 (N_26890,N_26037,N_25651);
and U26891 (N_26891,N_25266,N_25861);
nand U26892 (N_26892,N_25617,N_25324);
and U26893 (N_26893,N_25784,N_25255);
nor U26894 (N_26894,N_25241,N_25795);
xnor U26895 (N_26895,N_26145,N_25852);
nor U26896 (N_26896,N_25258,N_25634);
nor U26897 (N_26897,N_26165,N_25947);
and U26898 (N_26898,N_25694,N_26252);
nor U26899 (N_26899,N_26031,N_26383);
and U26900 (N_26900,N_25766,N_25755);
xor U26901 (N_26901,N_25943,N_25628);
nand U26902 (N_26902,N_26338,N_25274);
and U26903 (N_26903,N_26069,N_25520);
nor U26904 (N_26904,N_25542,N_26276);
xor U26905 (N_26905,N_26337,N_25704);
or U26906 (N_26906,N_25819,N_26256);
nor U26907 (N_26907,N_25247,N_26261);
xor U26908 (N_26908,N_26271,N_26177);
nand U26909 (N_26909,N_26381,N_26238);
xnor U26910 (N_26910,N_25997,N_25229);
or U26911 (N_26911,N_25783,N_26398);
xor U26912 (N_26912,N_25688,N_25905);
or U26913 (N_26913,N_25387,N_25676);
nor U26914 (N_26914,N_26314,N_25640);
or U26915 (N_26915,N_25631,N_25453);
nor U26916 (N_26916,N_25270,N_25885);
xor U26917 (N_26917,N_25910,N_26254);
or U26918 (N_26918,N_25294,N_26235);
xnor U26919 (N_26919,N_26343,N_25216);
nand U26920 (N_26920,N_25770,N_26072);
nor U26921 (N_26921,N_25702,N_25907);
and U26922 (N_26922,N_26099,N_25234);
nand U26923 (N_26923,N_25774,N_25886);
or U26924 (N_26924,N_25546,N_26346);
xnor U26925 (N_26925,N_26345,N_25456);
or U26926 (N_26926,N_26183,N_25643);
nand U26927 (N_26927,N_25248,N_25789);
nand U26928 (N_26928,N_25331,N_25573);
and U26929 (N_26929,N_25512,N_25696);
and U26930 (N_26930,N_25538,N_25874);
nand U26931 (N_26931,N_25961,N_25366);
or U26932 (N_26932,N_26393,N_26077);
or U26933 (N_26933,N_25848,N_25873);
nor U26934 (N_26934,N_25375,N_25866);
nand U26935 (N_26935,N_25502,N_26051);
and U26936 (N_26936,N_25814,N_25684);
and U26937 (N_26937,N_25574,N_25730);
nand U26938 (N_26938,N_25319,N_25724);
nor U26939 (N_26939,N_25212,N_25629);
nand U26940 (N_26940,N_25996,N_25626);
xor U26941 (N_26941,N_25741,N_25738);
nand U26942 (N_26942,N_25348,N_26307);
nor U26943 (N_26943,N_25450,N_25334);
and U26944 (N_26944,N_26297,N_25939);
nand U26945 (N_26945,N_25889,N_25210);
xor U26946 (N_26946,N_26395,N_26185);
nand U26947 (N_26947,N_25480,N_25843);
or U26948 (N_26948,N_25508,N_25820);
nand U26949 (N_26949,N_26259,N_26391);
xnor U26950 (N_26950,N_26146,N_25540);
and U26951 (N_26951,N_25660,N_26156);
xor U26952 (N_26952,N_25413,N_25977);
nor U26953 (N_26953,N_26153,N_25292);
nor U26954 (N_26954,N_25356,N_25721);
and U26955 (N_26955,N_25213,N_25597);
nor U26956 (N_26956,N_25999,N_26379);
nand U26957 (N_26957,N_26371,N_25832);
and U26958 (N_26958,N_25982,N_26329);
and U26959 (N_26959,N_26017,N_25256);
xnor U26960 (N_26960,N_26366,N_25420);
nand U26961 (N_26961,N_25461,N_25796);
and U26962 (N_26962,N_26041,N_25252);
or U26963 (N_26963,N_26263,N_25326);
xnor U26964 (N_26964,N_25489,N_25793);
and U26965 (N_26965,N_25701,N_25535);
nand U26966 (N_26966,N_25836,N_25399);
nor U26967 (N_26967,N_25571,N_26334);
and U26968 (N_26968,N_25924,N_26168);
and U26969 (N_26969,N_26097,N_26309);
or U26970 (N_26970,N_25434,N_25228);
nand U26971 (N_26971,N_25653,N_26143);
and U26972 (N_26972,N_25211,N_26294);
and U26973 (N_26973,N_25473,N_26284);
or U26974 (N_26974,N_25932,N_25611);
nand U26975 (N_26975,N_26130,N_25313);
xor U26976 (N_26976,N_25669,N_26036);
nand U26977 (N_26977,N_26304,N_26079);
and U26978 (N_26978,N_25779,N_26220);
nand U26979 (N_26979,N_25711,N_25594);
xor U26980 (N_26980,N_25742,N_25685);
nor U26981 (N_26981,N_26092,N_25739);
nor U26982 (N_26982,N_25847,N_25479);
xor U26983 (N_26983,N_26005,N_25743);
nor U26984 (N_26984,N_25840,N_26149);
and U26985 (N_26985,N_26138,N_26025);
or U26986 (N_26986,N_25958,N_25317);
and U26987 (N_26987,N_25222,N_25850);
and U26988 (N_26988,N_25204,N_25895);
nor U26989 (N_26989,N_25293,N_26066);
nor U26990 (N_26990,N_25219,N_26319);
and U26991 (N_26991,N_25726,N_26161);
xnor U26992 (N_26992,N_25303,N_26087);
nor U26993 (N_26993,N_25919,N_26027);
and U26994 (N_26994,N_25773,N_26018);
or U26995 (N_26995,N_26019,N_25967);
or U26996 (N_26996,N_26241,N_25930);
or U26997 (N_26997,N_26015,N_26044);
xor U26998 (N_26998,N_25801,N_25257);
and U26999 (N_26999,N_26089,N_25285);
and U27000 (N_27000,N_26019,N_25258);
xor U27001 (N_27001,N_26068,N_26106);
nand U27002 (N_27002,N_25965,N_25404);
or U27003 (N_27003,N_26014,N_26132);
or U27004 (N_27004,N_25467,N_25696);
nand U27005 (N_27005,N_25732,N_25314);
nor U27006 (N_27006,N_25218,N_25399);
and U27007 (N_27007,N_25782,N_25286);
nor U27008 (N_27008,N_26111,N_26002);
xor U27009 (N_27009,N_26323,N_25493);
nor U27010 (N_27010,N_25463,N_26228);
or U27011 (N_27011,N_26298,N_26264);
nor U27012 (N_27012,N_26342,N_25255);
or U27013 (N_27013,N_25380,N_25415);
nor U27014 (N_27014,N_26121,N_26230);
nor U27015 (N_27015,N_26196,N_25583);
or U27016 (N_27016,N_25856,N_25266);
nand U27017 (N_27017,N_25802,N_25751);
nor U27018 (N_27018,N_26240,N_26171);
nor U27019 (N_27019,N_26028,N_26068);
nor U27020 (N_27020,N_26357,N_26038);
or U27021 (N_27021,N_25950,N_25747);
or U27022 (N_27022,N_25453,N_25398);
or U27023 (N_27023,N_25310,N_25926);
xor U27024 (N_27024,N_25253,N_26074);
or U27025 (N_27025,N_25491,N_25303);
or U27026 (N_27026,N_26018,N_25793);
nor U27027 (N_27027,N_25370,N_26135);
xor U27028 (N_27028,N_26191,N_26277);
and U27029 (N_27029,N_25559,N_26204);
nor U27030 (N_27030,N_26075,N_26216);
nand U27031 (N_27031,N_26213,N_26136);
nand U27032 (N_27032,N_26340,N_26182);
xor U27033 (N_27033,N_25677,N_26315);
nand U27034 (N_27034,N_26036,N_26114);
or U27035 (N_27035,N_26221,N_25440);
or U27036 (N_27036,N_26030,N_26080);
nand U27037 (N_27037,N_25746,N_25501);
nor U27038 (N_27038,N_26320,N_25732);
xnor U27039 (N_27039,N_26297,N_25866);
nor U27040 (N_27040,N_26248,N_25656);
nand U27041 (N_27041,N_25264,N_25230);
and U27042 (N_27042,N_25661,N_25268);
or U27043 (N_27043,N_25426,N_25871);
and U27044 (N_27044,N_25270,N_26197);
nand U27045 (N_27045,N_25840,N_25793);
nand U27046 (N_27046,N_25490,N_25947);
xor U27047 (N_27047,N_25976,N_26087);
nor U27048 (N_27048,N_26356,N_25944);
nor U27049 (N_27049,N_26079,N_25580);
nor U27050 (N_27050,N_26124,N_25451);
xor U27051 (N_27051,N_25613,N_26108);
nand U27052 (N_27052,N_25577,N_25300);
nor U27053 (N_27053,N_25631,N_26399);
or U27054 (N_27054,N_25891,N_25773);
xor U27055 (N_27055,N_25565,N_26192);
xnor U27056 (N_27056,N_25401,N_25569);
xor U27057 (N_27057,N_25506,N_26035);
nor U27058 (N_27058,N_25671,N_25711);
and U27059 (N_27059,N_26298,N_25670);
or U27060 (N_27060,N_25778,N_25278);
xnor U27061 (N_27061,N_25604,N_26170);
and U27062 (N_27062,N_25456,N_25524);
nor U27063 (N_27063,N_26027,N_26083);
and U27064 (N_27064,N_25812,N_26042);
nor U27065 (N_27065,N_25295,N_26368);
or U27066 (N_27066,N_25500,N_26225);
or U27067 (N_27067,N_25688,N_26047);
or U27068 (N_27068,N_26062,N_25735);
nor U27069 (N_27069,N_26297,N_25792);
nand U27070 (N_27070,N_25396,N_25904);
or U27071 (N_27071,N_25644,N_25649);
or U27072 (N_27072,N_25811,N_26190);
nand U27073 (N_27073,N_25234,N_25729);
nor U27074 (N_27074,N_25467,N_25692);
or U27075 (N_27075,N_25721,N_25845);
and U27076 (N_27076,N_25991,N_25662);
nor U27077 (N_27077,N_26375,N_25227);
xnor U27078 (N_27078,N_26254,N_25403);
and U27079 (N_27079,N_25427,N_26005);
nor U27080 (N_27080,N_26367,N_25504);
or U27081 (N_27081,N_25370,N_25623);
nor U27082 (N_27082,N_26008,N_25309);
nand U27083 (N_27083,N_26143,N_25856);
nand U27084 (N_27084,N_26331,N_25645);
xnor U27085 (N_27085,N_26066,N_25433);
nor U27086 (N_27086,N_25409,N_25200);
or U27087 (N_27087,N_25713,N_25323);
nand U27088 (N_27088,N_26244,N_25401);
nor U27089 (N_27089,N_25958,N_26283);
xnor U27090 (N_27090,N_25533,N_25420);
xnor U27091 (N_27091,N_25908,N_25898);
and U27092 (N_27092,N_25749,N_26274);
nor U27093 (N_27093,N_25436,N_26189);
xnor U27094 (N_27094,N_26388,N_25820);
nand U27095 (N_27095,N_25868,N_26228);
nor U27096 (N_27096,N_25858,N_26327);
nor U27097 (N_27097,N_26026,N_25960);
nand U27098 (N_27098,N_26293,N_25507);
or U27099 (N_27099,N_26205,N_26043);
nor U27100 (N_27100,N_26344,N_26354);
nor U27101 (N_27101,N_25209,N_26330);
nand U27102 (N_27102,N_25889,N_26280);
xor U27103 (N_27103,N_25639,N_26037);
or U27104 (N_27104,N_25864,N_25219);
xnor U27105 (N_27105,N_25701,N_25495);
nand U27106 (N_27106,N_26166,N_26164);
nor U27107 (N_27107,N_25824,N_25287);
nand U27108 (N_27108,N_25708,N_25927);
nor U27109 (N_27109,N_26288,N_25340);
xnor U27110 (N_27110,N_25910,N_26305);
or U27111 (N_27111,N_25591,N_26009);
nand U27112 (N_27112,N_26270,N_25537);
xor U27113 (N_27113,N_25920,N_26249);
and U27114 (N_27114,N_26235,N_26130);
and U27115 (N_27115,N_25755,N_25308);
nand U27116 (N_27116,N_26149,N_26187);
xnor U27117 (N_27117,N_25670,N_26159);
and U27118 (N_27118,N_25399,N_26221);
nor U27119 (N_27119,N_26108,N_25356);
xor U27120 (N_27120,N_26292,N_25609);
or U27121 (N_27121,N_25585,N_26316);
xnor U27122 (N_27122,N_25966,N_25266);
or U27123 (N_27123,N_25367,N_25665);
xor U27124 (N_27124,N_26298,N_25774);
and U27125 (N_27125,N_26160,N_25706);
nand U27126 (N_27126,N_26290,N_25503);
nor U27127 (N_27127,N_25590,N_25784);
nand U27128 (N_27128,N_26306,N_25638);
xor U27129 (N_27129,N_26061,N_25639);
or U27130 (N_27130,N_26045,N_26088);
and U27131 (N_27131,N_25705,N_25977);
nand U27132 (N_27132,N_26052,N_26279);
and U27133 (N_27133,N_25807,N_25728);
nand U27134 (N_27134,N_26111,N_26238);
nor U27135 (N_27135,N_25961,N_25667);
nand U27136 (N_27136,N_25593,N_25404);
or U27137 (N_27137,N_26253,N_25818);
or U27138 (N_27138,N_25478,N_26051);
and U27139 (N_27139,N_25603,N_26064);
or U27140 (N_27140,N_25507,N_25969);
nand U27141 (N_27141,N_25209,N_26320);
and U27142 (N_27142,N_25936,N_26216);
xor U27143 (N_27143,N_25536,N_25621);
xnor U27144 (N_27144,N_25534,N_26282);
nor U27145 (N_27145,N_26203,N_25294);
xor U27146 (N_27146,N_25778,N_25932);
or U27147 (N_27147,N_25640,N_25375);
nand U27148 (N_27148,N_26025,N_26379);
xnor U27149 (N_27149,N_25813,N_26137);
or U27150 (N_27150,N_26242,N_26387);
nor U27151 (N_27151,N_25484,N_25696);
nor U27152 (N_27152,N_25552,N_25342);
nand U27153 (N_27153,N_25712,N_26200);
and U27154 (N_27154,N_26144,N_26109);
or U27155 (N_27155,N_25927,N_26057);
nor U27156 (N_27156,N_25657,N_25238);
xor U27157 (N_27157,N_26117,N_25316);
or U27158 (N_27158,N_25473,N_25958);
or U27159 (N_27159,N_25341,N_25475);
or U27160 (N_27160,N_26224,N_25583);
and U27161 (N_27161,N_25864,N_25443);
or U27162 (N_27162,N_25626,N_25943);
nor U27163 (N_27163,N_25851,N_25360);
nand U27164 (N_27164,N_25753,N_25346);
and U27165 (N_27165,N_25850,N_25990);
xnor U27166 (N_27166,N_25593,N_26254);
nor U27167 (N_27167,N_25318,N_25512);
nor U27168 (N_27168,N_25596,N_25490);
nor U27169 (N_27169,N_26291,N_25913);
and U27170 (N_27170,N_26298,N_25918);
and U27171 (N_27171,N_25891,N_25339);
or U27172 (N_27172,N_25621,N_25295);
nand U27173 (N_27173,N_25492,N_25623);
and U27174 (N_27174,N_25928,N_25485);
xnor U27175 (N_27175,N_26020,N_25416);
nor U27176 (N_27176,N_25416,N_25721);
or U27177 (N_27177,N_25526,N_26232);
nand U27178 (N_27178,N_25508,N_25445);
nand U27179 (N_27179,N_26331,N_25457);
and U27180 (N_27180,N_25343,N_25446);
nor U27181 (N_27181,N_25419,N_25434);
nand U27182 (N_27182,N_25386,N_25659);
and U27183 (N_27183,N_25899,N_26200);
nand U27184 (N_27184,N_25561,N_26353);
xor U27185 (N_27185,N_26144,N_25463);
nor U27186 (N_27186,N_25736,N_26120);
or U27187 (N_27187,N_26387,N_26193);
xnor U27188 (N_27188,N_25517,N_25551);
or U27189 (N_27189,N_25559,N_25421);
nand U27190 (N_27190,N_25556,N_26067);
nor U27191 (N_27191,N_25763,N_25668);
xnor U27192 (N_27192,N_25533,N_25408);
and U27193 (N_27193,N_25817,N_25291);
xor U27194 (N_27194,N_25735,N_25578);
xnor U27195 (N_27195,N_25595,N_26068);
xnor U27196 (N_27196,N_25727,N_25258);
and U27197 (N_27197,N_25539,N_26241);
xor U27198 (N_27198,N_25766,N_25230);
or U27199 (N_27199,N_25690,N_26229);
or U27200 (N_27200,N_26366,N_25963);
nand U27201 (N_27201,N_25495,N_25727);
nor U27202 (N_27202,N_26302,N_25628);
xor U27203 (N_27203,N_25537,N_25671);
or U27204 (N_27204,N_25634,N_25526);
or U27205 (N_27205,N_25455,N_25816);
nor U27206 (N_27206,N_25292,N_25998);
nand U27207 (N_27207,N_25622,N_26139);
or U27208 (N_27208,N_25796,N_25663);
or U27209 (N_27209,N_26315,N_25958);
xor U27210 (N_27210,N_25949,N_25601);
nand U27211 (N_27211,N_26353,N_25477);
nor U27212 (N_27212,N_25824,N_25926);
nand U27213 (N_27213,N_25446,N_26110);
and U27214 (N_27214,N_25591,N_25659);
or U27215 (N_27215,N_25501,N_26328);
nor U27216 (N_27216,N_25501,N_25644);
nor U27217 (N_27217,N_26131,N_26197);
and U27218 (N_27218,N_25323,N_25967);
and U27219 (N_27219,N_25294,N_25218);
nand U27220 (N_27220,N_25677,N_25592);
nor U27221 (N_27221,N_25373,N_26237);
nor U27222 (N_27222,N_25729,N_25978);
nand U27223 (N_27223,N_25759,N_25420);
xnor U27224 (N_27224,N_25663,N_25790);
nor U27225 (N_27225,N_25640,N_25702);
and U27226 (N_27226,N_25533,N_25467);
nand U27227 (N_27227,N_25561,N_26219);
nand U27228 (N_27228,N_25877,N_25752);
nor U27229 (N_27229,N_25255,N_25522);
nand U27230 (N_27230,N_25614,N_25920);
xor U27231 (N_27231,N_25645,N_25360);
and U27232 (N_27232,N_26143,N_25724);
and U27233 (N_27233,N_25945,N_25675);
or U27234 (N_27234,N_25852,N_25912);
nand U27235 (N_27235,N_25747,N_25347);
and U27236 (N_27236,N_25990,N_25409);
nor U27237 (N_27237,N_25381,N_26035);
xor U27238 (N_27238,N_25834,N_25696);
or U27239 (N_27239,N_25867,N_26293);
and U27240 (N_27240,N_25756,N_26159);
nor U27241 (N_27241,N_26376,N_25299);
xor U27242 (N_27242,N_25878,N_25742);
xor U27243 (N_27243,N_26272,N_25511);
xnor U27244 (N_27244,N_25902,N_25315);
or U27245 (N_27245,N_26319,N_25216);
and U27246 (N_27246,N_25780,N_26042);
and U27247 (N_27247,N_26298,N_26386);
xnor U27248 (N_27248,N_25299,N_25483);
or U27249 (N_27249,N_26374,N_25659);
and U27250 (N_27250,N_26361,N_25397);
and U27251 (N_27251,N_26150,N_25511);
xor U27252 (N_27252,N_26366,N_25771);
nand U27253 (N_27253,N_26160,N_25451);
xnor U27254 (N_27254,N_26348,N_26147);
and U27255 (N_27255,N_25720,N_26398);
xnor U27256 (N_27256,N_26261,N_25858);
nand U27257 (N_27257,N_25664,N_26374);
nor U27258 (N_27258,N_26329,N_26336);
nand U27259 (N_27259,N_25957,N_26234);
and U27260 (N_27260,N_25641,N_26100);
or U27261 (N_27261,N_26010,N_26002);
nand U27262 (N_27262,N_26325,N_26040);
or U27263 (N_27263,N_26285,N_25220);
nand U27264 (N_27264,N_25822,N_26343);
nand U27265 (N_27265,N_25467,N_26366);
nand U27266 (N_27266,N_25681,N_25492);
or U27267 (N_27267,N_26253,N_26079);
nand U27268 (N_27268,N_25926,N_26269);
and U27269 (N_27269,N_25288,N_25425);
or U27270 (N_27270,N_25676,N_25961);
nor U27271 (N_27271,N_26122,N_26091);
nor U27272 (N_27272,N_25709,N_25357);
nand U27273 (N_27273,N_26000,N_26315);
or U27274 (N_27274,N_26101,N_25405);
or U27275 (N_27275,N_26221,N_26153);
and U27276 (N_27276,N_26188,N_25427);
or U27277 (N_27277,N_26020,N_25756);
xor U27278 (N_27278,N_25472,N_26253);
and U27279 (N_27279,N_25595,N_25280);
and U27280 (N_27280,N_25691,N_25942);
or U27281 (N_27281,N_25698,N_25858);
nand U27282 (N_27282,N_25401,N_26368);
or U27283 (N_27283,N_25639,N_25871);
and U27284 (N_27284,N_25715,N_26311);
xnor U27285 (N_27285,N_26273,N_25543);
xor U27286 (N_27286,N_26361,N_25304);
nand U27287 (N_27287,N_25715,N_25298);
and U27288 (N_27288,N_25765,N_25744);
nor U27289 (N_27289,N_26295,N_25582);
xor U27290 (N_27290,N_25450,N_25208);
nor U27291 (N_27291,N_25524,N_25727);
xnor U27292 (N_27292,N_25916,N_25339);
or U27293 (N_27293,N_25576,N_26151);
nand U27294 (N_27294,N_25343,N_25317);
nand U27295 (N_27295,N_25461,N_26339);
or U27296 (N_27296,N_25649,N_25463);
or U27297 (N_27297,N_25817,N_26240);
nand U27298 (N_27298,N_25441,N_25572);
or U27299 (N_27299,N_25937,N_26121);
and U27300 (N_27300,N_25550,N_26348);
xnor U27301 (N_27301,N_25888,N_25993);
and U27302 (N_27302,N_25535,N_26042);
and U27303 (N_27303,N_26315,N_26234);
nand U27304 (N_27304,N_25358,N_26347);
nand U27305 (N_27305,N_25773,N_25832);
nand U27306 (N_27306,N_26124,N_26250);
nand U27307 (N_27307,N_25275,N_25830);
and U27308 (N_27308,N_26215,N_25407);
nand U27309 (N_27309,N_25282,N_26066);
nand U27310 (N_27310,N_26385,N_25874);
or U27311 (N_27311,N_25310,N_26163);
nor U27312 (N_27312,N_26010,N_25984);
nand U27313 (N_27313,N_25642,N_25852);
or U27314 (N_27314,N_25381,N_26385);
xor U27315 (N_27315,N_26092,N_26241);
xor U27316 (N_27316,N_25724,N_26203);
xnor U27317 (N_27317,N_26240,N_26297);
nand U27318 (N_27318,N_25663,N_26011);
and U27319 (N_27319,N_25919,N_25621);
nand U27320 (N_27320,N_26005,N_25883);
xnor U27321 (N_27321,N_26038,N_25499);
nor U27322 (N_27322,N_25499,N_25335);
or U27323 (N_27323,N_25246,N_25352);
and U27324 (N_27324,N_25385,N_25226);
xor U27325 (N_27325,N_25882,N_25301);
and U27326 (N_27326,N_25608,N_25319);
and U27327 (N_27327,N_25366,N_25259);
and U27328 (N_27328,N_25590,N_25683);
nor U27329 (N_27329,N_26048,N_25554);
nand U27330 (N_27330,N_26398,N_26399);
and U27331 (N_27331,N_26001,N_26015);
nand U27332 (N_27332,N_25222,N_26358);
nand U27333 (N_27333,N_25249,N_25527);
or U27334 (N_27334,N_26204,N_25961);
or U27335 (N_27335,N_26259,N_26175);
and U27336 (N_27336,N_25455,N_25248);
xor U27337 (N_27337,N_25735,N_26385);
and U27338 (N_27338,N_25570,N_25551);
nor U27339 (N_27339,N_26186,N_25233);
nor U27340 (N_27340,N_26089,N_26354);
nand U27341 (N_27341,N_26004,N_26007);
xnor U27342 (N_27342,N_26138,N_26258);
nand U27343 (N_27343,N_25553,N_26173);
nor U27344 (N_27344,N_26217,N_25515);
and U27345 (N_27345,N_26029,N_26315);
nand U27346 (N_27346,N_25225,N_25316);
and U27347 (N_27347,N_25671,N_26180);
or U27348 (N_27348,N_25576,N_26168);
nand U27349 (N_27349,N_25482,N_25745);
nand U27350 (N_27350,N_25950,N_25716);
or U27351 (N_27351,N_26171,N_26310);
or U27352 (N_27352,N_26198,N_25894);
and U27353 (N_27353,N_26072,N_25758);
xor U27354 (N_27354,N_25930,N_25648);
or U27355 (N_27355,N_25417,N_25288);
nand U27356 (N_27356,N_25773,N_25215);
nor U27357 (N_27357,N_25218,N_26316);
nand U27358 (N_27358,N_25581,N_25317);
nand U27359 (N_27359,N_26221,N_25669);
nand U27360 (N_27360,N_26047,N_25243);
nand U27361 (N_27361,N_25605,N_25216);
or U27362 (N_27362,N_26164,N_25205);
and U27363 (N_27363,N_26384,N_26107);
or U27364 (N_27364,N_25934,N_25996);
nand U27365 (N_27365,N_26064,N_25674);
nand U27366 (N_27366,N_25214,N_25451);
nand U27367 (N_27367,N_25766,N_25301);
nor U27368 (N_27368,N_25979,N_26140);
and U27369 (N_27369,N_26057,N_25813);
and U27370 (N_27370,N_25635,N_26210);
nor U27371 (N_27371,N_25954,N_25765);
nor U27372 (N_27372,N_26192,N_25399);
nand U27373 (N_27373,N_25225,N_26347);
or U27374 (N_27374,N_26172,N_26354);
nor U27375 (N_27375,N_25598,N_26185);
xor U27376 (N_27376,N_26222,N_25253);
xor U27377 (N_27377,N_26321,N_25240);
nand U27378 (N_27378,N_25657,N_25348);
and U27379 (N_27379,N_26246,N_26123);
and U27380 (N_27380,N_26324,N_25487);
or U27381 (N_27381,N_25497,N_25316);
xnor U27382 (N_27382,N_25320,N_25322);
xnor U27383 (N_27383,N_26217,N_25605);
nand U27384 (N_27384,N_25733,N_26254);
xnor U27385 (N_27385,N_25705,N_25751);
nand U27386 (N_27386,N_25933,N_26080);
nor U27387 (N_27387,N_25358,N_26242);
or U27388 (N_27388,N_25403,N_25377);
nor U27389 (N_27389,N_26261,N_25339);
and U27390 (N_27390,N_25446,N_26104);
or U27391 (N_27391,N_25702,N_26238);
or U27392 (N_27392,N_25953,N_25217);
nor U27393 (N_27393,N_25352,N_25772);
xor U27394 (N_27394,N_25864,N_25231);
nand U27395 (N_27395,N_25955,N_25345);
nand U27396 (N_27396,N_25858,N_25884);
or U27397 (N_27397,N_25933,N_25271);
nor U27398 (N_27398,N_25200,N_26196);
nand U27399 (N_27399,N_25240,N_25417);
xnor U27400 (N_27400,N_25924,N_25968);
xnor U27401 (N_27401,N_25898,N_25568);
and U27402 (N_27402,N_25834,N_25551);
nand U27403 (N_27403,N_25316,N_25706);
or U27404 (N_27404,N_25367,N_25288);
nand U27405 (N_27405,N_26342,N_25772);
or U27406 (N_27406,N_25206,N_26090);
nand U27407 (N_27407,N_25531,N_25843);
or U27408 (N_27408,N_25253,N_26327);
nand U27409 (N_27409,N_25233,N_25310);
xnor U27410 (N_27410,N_25585,N_25697);
nand U27411 (N_27411,N_25644,N_26048);
and U27412 (N_27412,N_26078,N_25676);
xnor U27413 (N_27413,N_25777,N_25291);
xor U27414 (N_27414,N_26209,N_26295);
and U27415 (N_27415,N_26333,N_25931);
or U27416 (N_27416,N_25201,N_25699);
nand U27417 (N_27417,N_25478,N_26118);
and U27418 (N_27418,N_26360,N_25834);
nor U27419 (N_27419,N_25852,N_25951);
nor U27420 (N_27420,N_25791,N_25362);
xnor U27421 (N_27421,N_26070,N_26230);
xor U27422 (N_27422,N_25789,N_25826);
nand U27423 (N_27423,N_25983,N_26071);
and U27424 (N_27424,N_25211,N_25881);
and U27425 (N_27425,N_25857,N_25513);
xnor U27426 (N_27426,N_26282,N_25889);
nand U27427 (N_27427,N_26113,N_25498);
nor U27428 (N_27428,N_25845,N_25706);
and U27429 (N_27429,N_25263,N_25865);
xor U27430 (N_27430,N_26270,N_26083);
nand U27431 (N_27431,N_26341,N_25848);
nor U27432 (N_27432,N_26233,N_25786);
nor U27433 (N_27433,N_26340,N_25727);
nand U27434 (N_27434,N_25240,N_26361);
and U27435 (N_27435,N_25343,N_25260);
nor U27436 (N_27436,N_25267,N_25748);
xor U27437 (N_27437,N_25424,N_25278);
and U27438 (N_27438,N_25724,N_25460);
nand U27439 (N_27439,N_26064,N_26007);
xnor U27440 (N_27440,N_26018,N_25762);
or U27441 (N_27441,N_26387,N_26118);
xnor U27442 (N_27442,N_26010,N_25692);
nand U27443 (N_27443,N_26323,N_26010);
nor U27444 (N_27444,N_25522,N_26300);
xnor U27445 (N_27445,N_25726,N_25206);
and U27446 (N_27446,N_26358,N_25264);
xnor U27447 (N_27447,N_25972,N_25417);
xnor U27448 (N_27448,N_25877,N_26076);
nor U27449 (N_27449,N_25760,N_25998);
and U27450 (N_27450,N_25776,N_26230);
xnor U27451 (N_27451,N_25433,N_25779);
or U27452 (N_27452,N_25908,N_26284);
nor U27453 (N_27453,N_26323,N_25400);
or U27454 (N_27454,N_26138,N_25462);
or U27455 (N_27455,N_25972,N_26026);
or U27456 (N_27456,N_26263,N_25963);
nand U27457 (N_27457,N_26111,N_26204);
and U27458 (N_27458,N_25257,N_25477);
or U27459 (N_27459,N_25908,N_26374);
xnor U27460 (N_27460,N_25807,N_25375);
and U27461 (N_27461,N_26184,N_26341);
nor U27462 (N_27462,N_25326,N_26128);
nand U27463 (N_27463,N_25220,N_25954);
nand U27464 (N_27464,N_25928,N_25387);
xnor U27465 (N_27465,N_25602,N_25972);
nor U27466 (N_27466,N_25254,N_25295);
or U27467 (N_27467,N_25986,N_25238);
or U27468 (N_27468,N_25473,N_25947);
and U27469 (N_27469,N_25903,N_26051);
and U27470 (N_27470,N_25203,N_25216);
nor U27471 (N_27471,N_25818,N_26101);
xor U27472 (N_27472,N_26057,N_26245);
or U27473 (N_27473,N_25551,N_25734);
nand U27474 (N_27474,N_25755,N_25875);
or U27475 (N_27475,N_25533,N_25282);
or U27476 (N_27476,N_25390,N_25904);
nand U27477 (N_27477,N_25553,N_25399);
xor U27478 (N_27478,N_26381,N_26009);
xnor U27479 (N_27479,N_26126,N_25285);
nor U27480 (N_27480,N_25868,N_25615);
and U27481 (N_27481,N_25751,N_25400);
and U27482 (N_27482,N_25334,N_25335);
and U27483 (N_27483,N_26183,N_26022);
and U27484 (N_27484,N_26181,N_25654);
or U27485 (N_27485,N_25582,N_25222);
nor U27486 (N_27486,N_26060,N_25745);
nand U27487 (N_27487,N_25225,N_25496);
or U27488 (N_27488,N_25999,N_26293);
or U27489 (N_27489,N_26246,N_26103);
or U27490 (N_27490,N_26218,N_25892);
nor U27491 (N_27491,N_25685,N_25870);
nor U27492 (N_27492,N_25623,N_25653);
nor U27493 (N_27493,N_26268,N_26040);
nand U27494 (N_27494,N_25576,N_25451);
nor U27495 (N_27495,N_26092,N_25911);
xnor U27496 (N_27496,N_25547,N_26386);
xnor U27497 (N_27497,N_25560,N_26031);
nor U27498 (N_27498,N_26385,N_25479);
and U27499 (N_27499,N_26361,N_26321);
nor U27500 (N_27500,N_26300,N_25902);
xor U27501 (N_27501,N_26315,N_25735);
nor U27502 (N_27502,N_25904,N_25986);
nand U27503 (N_27503,N_25250,N_25701);
xnor U27504 (N_27504,N_26294,N_25968);
nor U27505 (N_27505,N_26266,N_25978);
nor U27506 (N_27506,N_25574,N_26122);
and U27507 (N_27507,N_26003,N_25954);
xor U27508 (N_27508,N_25289,N_25505);
nor U27509 (N_27509,N_26344,N_25806);
or U27510 (N_27510,N_26269,N_26003);
nor U27511 (N_27511,N_25730,N_25776);
xor U27512 (N_27512,N_26330,N_26343);
or U27513 (N_27513,N_25620,N_25560);
xnor U27514 (N_27514,N_26017,N_25785);
nand U27515 (N_27515,N_25221,N_25939);
and U27516 (N_27516,N_26155,N_26005);
and U27517 (N_27517,N_25343,N_26362);
or U27518 (N_27518,N_26119,N_25472);
and U27519 (N_27519,N_25923,N_26319);
nand U27520 (N_27520,N_25820,N_26023);
xnor U27521 (N_27521,N_26246,N_25848);
nor U27522 (N_27522,N_25534,N_25702);
or U27523 (N_27523,N_25759,N_26094);
and U27524 (N_27524,N_26274,N_25279);
nand U27525 (N_27525,N_26015,N_25460);
or U27526 (N_27526,N_25483,N_25618);
nor U27527 (N_27527,N_25344,N_25531);
or U27528 (N_27528,N_26241,N_25397);
xnor U27529 (N_27529,N_25660,N_25567);
and U27530 (N_27530,N_25368,N_25360);
xnor U27531 (N_27531,N_25805,N_26209);
xor U27532 (N_27532,N_25987,N_25515);
nand U27533 (N_27533,N_26180,N_26077);
nand U27534 (N_27534,N_25387,N_25925);
xnor U27535 (N_27535,N_25227,N_26233);
and U27536 (N_27536,N_25251,N_25902);
nor U27537 (N_27537,N_25279,N_25764);
and U27538 (N_27538,N_25922,N_25353);
nand U27539 (N_27539,N_25293,N_26104);
xnor U27540 (N_27540,N_26293,N_25579);
xnor U27541 (N_27541,N_26337,N_25801);
nand U27542 (N_27542,N_25316,N_25504);
or U27543 (N_27543,N_25709,N_25733);
xor U27544 (N_27544,N_26226,N_25358);
nor U27545 (N_27545,N_26183,N_26250);
and U27546 (N_27546,N_26060,N_25525);
xor U27547 (N_27547,N_25639,N_26014);
nor U27548 (N_27548,N_25210,N_26231);
nand U27549 (N_27549,N_25280,N_25687);
xnor U27550 (N_27550,N_26188,N_26273);
nor U27551 (N_27551,N_25471,N_26158);
nor U27552 (N_27552,N_25869,N_25864);
nand U27553 (N_27553,N_25590,N_25882);
and U27554 (N_27554,N_25553,N_25622);
and U27555 (N_27555,N_25483,N_25869);
nand U27556 (N_27556,N_25544,N_26081);
nand U27557 (N_27557,N_25684,N_25375);
nand U27558 (N_27558,N_25381,N_25336);
or U27559 (N_27559,N_25874,N_25352);
or U27560 (N_27560,N_25826,N_26393);
or U27561 (N_27561,N_26179,N_25894);
nor U27562 (N_27562,N_25966,N_26248);
nor U27563 (N_27563,N_26053,N_25540);
nand U27564 (N_27564,N_26107,N_26259);
nor U27565 (N_27565,N_25985,N_26224);
nor U27566 (N_27566,N_25934,N_26201);
or U27567 (N_27567,N_25544,N_25804);
or U27568 (N_27568,N_25763,N_25749);
and U27569 (N_27569,N_25614,N_26255);
or U27570 (N_27570,N_25220,N_25857);
or U27571 (N_27571,N_25278,N_26157);
nand U27572 (N_27572,N_26114,N_25883);
or U27573 (N_27573,N_26292,N_25887);
and U27574 (N_27574,N_26380,N_26225);
xnor U27575 (N_27575,N_26242,N_25966);
nor U27576 (N_27576,N_25801,N_25936);
xor U27577 (N_27577,N_26090,N_25232);
or U27578 (N_27578,N_25814,N_25234);
nor U27579 (N_27579,N_25947,N_25474);
nand U27580 (N_27580,N_25314,N_25670);
nor U27581 (N_27581,N_26240,N_25546);
or U27582 (N_27582,N_25965,N_25452);
nand U27583 (N_27583,N_25761,N_25984);
and U27584 (N_27584,N_26015,N_26355);
xor U27585 (N_27585,N_25915,N_25582);
nand U27586 (N_27586,N_26041,N_26306);
or U27587 (N_27587,N_25359,N_26086);
xor U27588 (N_27588,N_25405,N_25475);
nand U27589 (N_27589,N_25419,N_25916);
nor U27590 (N_27590,N_26225,N_25466);
xor U27591 (N_27591,N_26207,N_26081);
or U27592 (N_27592,N_25708,N_26339);
nand U27593 (N_27593,N_25417,N_26069);
nor U27594 (N_27594,N_25289,N_26252);
xor U27595 (N_27595,N_26220,N_26008);
and U27596 (N_27596,N_26337,N_26105);
xnor U27597 (N_27597,N_25832,N_25423);
nor U27598 (N_27598,N_25730,N_26364);
xnor U27599 (N_27599,N_25459,N_25889);
xor U27600 (N_27600,N_27383,N_26556);
nor U27601 (N_27601,N_27376,N_26948);
xor U27602 (N_27602,N_27360,N_26659);
nand U27603 (N_27603,N_26786,N_27177);
xnor U27604 (N_27604,N_26779,N_26692);
nand U27605 (N_27605,N_26686,N_27489);
and U27606 (N_27606,N_26977,N_26730);
nor U27607 (N_27607,N_26433,N_26896);
xnor U27608 (N_27608,N_26778,N_27029);
and U27609 (N_27609,N_27362,N_27225);
xnor U27610 (N_27610,N_27413,N_27438);
and U27611 (N_27611,N_26849,N_26437);
nand U27612 (N_27612,N_27369,N_26402);
or U27613 (N_27613,N_27488,N_26997);
nand U27614 (N_27614,N_26870,N_26553);
xnor U27615 (N_27615,N_26625,N_26712);
and U27616 (N_27616,N_26578,N_27178);
xnor U27617 (N_27617,N_27444,N_26764);
nor U27618 (N_27618,N_26755,N_26975);
nand U27619 (N_27619,N_27430,N_27135);
nor U27620 (N_27620,N_26689,N_26912);
nor U27621 (N_27621,N_26528,N_27211);
nand U27622 (N_27622,N_26966,N_26717);
nand U27623 (N_27623,N_26781,N_27311);
nand U27624 (N_27624,N_26508,N_26559);
nor U27625 (N_27625,N_27401,N_26996);
nor U27626 (N_27626,N_26859,N_26926);
and U27627 (N_27627,N_26703,N_27270);
and U27628 (N_27628,N_27012,N_26493);
and U27629 (N_27629,N_26964,N_26872);
xor U27630 (N_27630,N_26843,N_27333);
nor U27631 (N_27631,N_26456,N_26737);
or U27632 (N_27632,N_27374,N_26706);
and U27633 (N_27633,N_26688,N_26491);
xnor U27634 (N_27634,N_26435,N_27336);
and U27635 (N_27635,N_26772,N_27290);
xor U27636 (N_27636,N_27396,N_26609);
nand U27637 (N_27637,N_26457,N_27384);
xor U27638 (N_27638,N_27160,N_27163);
and U27639 (N_27639,N_26807,N_26665);
nand U27640 (N_27640,N_27260,N_26969);
xor U27641 (N_27641,N_27455,N_27089);
xnor U27642 (N_27642,N_26763,N_27036);
and U27643 (N_27643,N_26761,N_26630);
nor U27644 (N_27644,N_27134,N_26418);
nand U27645 (N_27645,N_27068,N_27133);
nor U27646 (N_27646,N_27596,N_27501);
xnor U27647 (N_27647,N_27569,N_27080);
xor U27648 (N_27648,N_26681,N_27512);
nor U27649 (N_27649,N_27052,N_27033);
xnor U27650 (N_27650,N_26573,N_27576);
and U27651 (N_27651,N_26612,N_26666);
nor U27652 (N_27652,N_27355,N_26751);
xnor U27653 (N_27653,N_26978,N_26592);
and U27654 (N_27654,N_26757,N_26961);
and U27655 (N_27655,N_26511,N_26902);
and U27656 (N_27656,N_26434,N_26588);
nand U27657 (N_27657,N_27233,N_27166);
nor U27658 (N_27658,N_26711,N_27300);
nand U27659 (N_27659,N_26445,N_27461);
xnor U27660 (N_27660,N_26488,N_26444);
nand U27661 (N_27661,N_26981,N_27475);
and U27662 (N_27662,N_26601,N_26947);
nand U27663 (N_27663,N_26586,N_27456);
xnor U27664 (N_27664,N_26576,N_26503);
or U27665 (N_27665,N_27168,N_26669);
and U27666 (N_27666,N_27185,N_26982);
nor U27667 (N_27667,N_27464,N_26621);
nand U27668 (N_27668,N_27148,N_27516);
and U27669 (N_27669,N_26985,N_27105);
xnor U27670 (N_27670,N_26745,N_27193);
or U27671 (N_27671,N_26863,N_26959);
nand U27672 (N_27672,N_27146,N_27329);
xor U27673 (N_27673,N_27494,N_27522);
or U27674 (N_27674,N_27305,N_26547);
nor U27675 (N_27675,N_27157,N_27531);
and U27676 (N_27676,N_27171,N_27428);
and U27677 (N_27677,N_26722,N_26837);
or U27678 (N_27678,N_27212,N_27010);
and U27679 (N_27679,N_27139,N_27370);
nand U27680 (N_27680,N_27429,N_27125);
and U27681 (N_27681,N_26844,N_26585);
nor U27682 (N_27682,N_27126,N_27006);
nor U27683 (N_27683,N_27122,N_26847);
and U27684 (N_27684,N_27152,N_27007);
nor U27685 (N_27685,N_27434,N_27041);
or U27686 (N_27686,N_27504,N_26638);
nand U27687 (N_27687,N_26683,N_26853);
or U27688 (N_27688,N_26841,N_26965);
and U27689 (N_27689,N_26930,N_27457);
nand U27690 (N_27690,N_27321,N_27109);
and U27691 (N_27691,N_26526,N_26879);
and U27692 (N_27692,N_27322,N_27317);
nand U27693 (N_27693,N_27519,N_26685);
nand U27694 (N_27694,N_26980,N_26955);
nand U27695 (N_27695,N_27348,N_26939);
nand U27696 (N_27696,N_26998,N_26992);
xor U27697 (N_27697,N_26700,N_27053);
nand U27698 (N_27698,N_26538,N_26798);
nand U27699 (N_27699,N_26424,N_26584);
xnor U27700 (N_27700,N_27441,N_27031);
nor U27701 (N_27701,N_27580,N_27116);
and U27702 (N_27702,N_27480,N_27502);
or U27703 (N_27703,N_27045,N_26794);
nor U27704 (N_27704,N_27448,N_26835);
xor U27705 (N_27705,N_27373,N_26554);
nor U27706 (N_27706,N_27078,N_27275);
nor U27707 (N_27707,N_27055,N_26639);
and U27708 (N_27708,N_26884,N_26525);
and U27709 (N_27709,N_27297,N_26651);
and U27710 (N_27710,N_26723,N_27472);
nor U27711 (N_27711,N_27402,N_27347);
xor U27712 (N_27712,N_27106,N_26495);
nor U27713 (N_27713,N_27537,N_27183);
xor U27714 (N_27714,N_27386,N_26768);
nor U27715 (N_27715,N_26986,N_26851);
and U27716 (N_27716,N_26820,N_26658);
nor U27717 (N_27717,N_26512,N_27087);
nand U27718 (N_27718,N_27389,N_26784);
nand U27719 (N_27719,N_27553,N_27539);
or U27720 (N_27720,N_27289,N_26549);
and U27721 (N_27721,N_27548,N_27412);
and U27722 (N_27722,N_27063,N_26782);
or U27723 (N_27723,N_26958,N_27190);
or U27724 (N_27724,N_27547,N_27247);
nand U27725 (N_27725,N_26480,N_27584);
nand U27726 (N_27726,N_26829,N_27001);
and U27727 (N_27727,N_27021,N_27182);
and U27728 (N_27728,N_26832,N_27567);
nand U27729 (N_27729,N_27077,N_26860);
nand U27730 (N_27730,N_27435,N_26811);
and U27731 (N_27731,N_26888,N_26803);
or U27732 (N_27732,N_27020,N_26759);
nor U27733 (N_27733,N_26485,N_27064);
and U27734 (N_27734,N_26756,N_27170);
or U27735 (N_27735,N_26569,N_26725);
nand U27736 (N_27736,N_27418,N_26881);
or U27737 (N_27737,N_27127,N_27030);
or U27738 (N_27738,N_26889,N_26758);
nand U27739 (N_27739,N_27459,N_27156);
or U27740 (N_27740,N_27218,N_26441);
and U27741 (N_27741,N_27203,N_26627);
nor U27742 (N_27742,N_26901,N_26907);
xnor U27743 (N_27743,N_26857,N_27091);
or U27744 (N_27744,N_26645,N_26661);
nor U27745 (N_27745,N_27253,N_26461);
xor U27746 (N_27746,N_27585,N_27381);
nand U27747 (N_27747,N_26475,N_26925);
nand U27748 (N_27748,N_27235,N_27194);
nor U27749 (N_27749,N_27568,N_26810);
and U27750 (N_27750,N_26915,N_27479);
and U27751 (N_27751,N_26482,N_27111);
and U27752 (N_27752,N_26505,N_26951);
nor U27753 (N_27753,N_27346,N_26905);
nor U27754 (N_27754,N_26701,N_26417);
or U27755 (N_27755,N_27299,N_27529);
or U27756 (N_27756,N_27560,N_27312);
and U27757 (N_27757,N_26571,N_27083);
or U27758 (N_27758,N_27236,N_26924);
nor U27759 (N_27759,N_26776,N_26492);
nand U27760 (N_27760,N_27257,N_26671);
and U27761 (N_27761,N_27433,N_26945);
nor U27762 (N_27762,N_27535,N_27285);
xnor U27763 (N_27763,N_26497,N_27060);
or U27764 (N_27764,N_27103,N_26770);
nand U27765 (N_27765,N_26806,N_27250);
nand U27766 (N_27766,N_26773,N_26421);
xnor U27767 (N_27767,N_27432,N_27579);
nor U27768 (N_27768,N_26419,N_27491);
nor U27769 (N_27769,N_27069,N_26777);
nor U27770 (N_27770,N_26960,N_27410);
nand U27771 (N_27771,N_27061,N_27387);
and U27772 (N_27772,N_27405,N_27566);
or U27773 (N_27773,N_26679,N_26801);
and U27774 (N_27774,N_27352,N_26771);
or U27775 (N_27775,N_27406,N_27093);
or U27776 (N_27776,N_27572,N_26707);
and U27777 (N_27777,N_27356,N_27308);
nand U27778 (N_27778,N_26504,N_27378);
or U27779 (N_27779,N_26510,N_26993);
nor U27780 (N_27780,N_26611,N_27481);
xnor U27781 (N_27781,N_27325,N_27104);
or U27782 (N_27782,N_26566,N_26478);
or U27783 (N_27783,N_26551,N_27174);
nor U27784 (N_27784,N_26854,N_26675);
nand U27785 (N_27785,N_27540,N_27145);
and U27786 (N_27786,N_27578,N_26414);
or U27787 (N_27787,N_26463,N_26867);
xor U27788 (N_27788,N_27533,N_27188);
and U27789 (N_27789,N_26727,N_27016);
nor U27790 (N_27790,N_26775,N_27581);
or U27791 (N_27791,N_27117,N_26868);
xnor U27792 (N_27792,N_26968,N_27261);
nor U27793 (N_27793,N_26670,N_26911);
and U27794 (N_27794,N_27124,N_26608);
xor U27795 (N_27795,N_26941,N_27474);
nor U27796 (N_27796,N_27119,N_27266);
and U27797 (N_27797,N_27202,N_27380);
and U27798 (N_27798,N_27196,N_26502);
nor U27799 (N_27799,N_27513,N_27478);
and U27800 (N_27800,N_26999,N_27268);
xor U27801 (N_27801,N_26967,N_27408);
and U27802 (N_27802,N_27315,N_26691);
nor U27803 (N_27803,N_27096,N_26438);
or U27804 (N_27804,N_26827,N_27573);
and U27805 (N_27805,N_26793,N_27227);
and U27806 (N_27806,N_27546,N_27199);
nand U27807 (N_27807,N_26788,N_27192);
and U27808 (N_27808,N_27217,N_27331);
xor U27809 (N_27809,N_27110,N_27128);
nand U27810 (N_27810,N_27267,N_27138);
and U27811 (N_27811,N_27240,N_26732);
nand U27812 (N_27812,N_26876,N_27019);
or U27813 (N_27813,N_27027,N_27467);
or U27814 (N_27814,N_27463,N_27309);
xnor U27815 (N_27815,N_27047,N_26410);
nand U27816 (N_27816,N_27208,N_27051);
nand U27817 (N_27817,N_26921,N_26971);
xnor U27818 (N_27818,N_26555,N_27294);
and U27819 (N_27819,N_26979,N_26957);
or U27820 (N_27820,N_26697,N_27214);
and U27821 (N_27821,N_26815,N_26831);
or U27822 (N_27822,N_27070,N_27044);
and U27823 (N_27823,N_26606,N_26818);
nor U27824 (N_27824,N_26878,N_27179);
and U27825 (N_27825,N_27351,N_27427);
nand U27826 (N_27826,N_26680,N_26792);
and U27827 (N_27827,N_26411,N_26486);
and U27828 (N_27828,N_27219,N_27498);
or U27829 (N_27829,N_27372,N_27079);
xnor U27830 (N_27830,N_26933,N_26822);
nor U27831 (N_27831,N_27514,N_27525);
xor U27832 (N_27832,N_26436,N_27132);
and U27833 (N_27833,N_27407,N_27364);
nand U27834 (N_27834,N_26604,N_27411);
or U27835 (N_27835,N_26626,N_26649);
or U27836 (N_27836,N_27436,N_27147);
or U27837 (N_27837,N_26581,N_26442);
nor U27838 (N_27838,N_27082,N_27292);
nor U27839 (N_27839,N_27162,N_26534);
xor U27840 (N_27840,N_27011,N_26970);
or U27841 (N_27841,N_27536,N_27353);
nor U27842 (N_27842,N_26826,N_27226);
or U27843 (N_27843,N_27420,N_27142);
and U27844 (N_27844,N_27040,N_27088);
xnor U27845 (N_27845,N_27090,N_27186);
nor U27846 (N_27846,N_27151,N_26423);
nor U27847 (N_27847,N_27258,N_27107);
nand U27848 (N_27848,N_27035,N_27549);
xor U27849 (N_27849,N_26940,N_26962);
or U27850 (N_27850,N_27446,N_26883);
xor U27851 (N_27851,N_26575,N_27158);
nand U27852 (N_27852,N_26949,N_27555);
nand U27853 (N_27853,N_26875,N_27517);
xor U27854 (N_27854,N_26650,N_27154);
nor U27855 (N_27855,N_26568,N_27014);
xor U27856 (N_27856,N_27367,N_26674);
nor U27857 (N_27857,N_27101,N_26895);
xor U27858 (N_27858,N_26774,N_26744);
nand U27859 (N_27859,N_26963,N_26714);
and U27860 (N_27860,N_27447,N_27454);
xnor U27861 (N_27861,N_27506,N_26540);
or U27862 (N_27862,N_27224,N_27097);
or U27863 (N_27863,N_26459,N_26563);
nand U27864 (N_27864,N_27487,N_26432);
nand U27865 (N_27865,N_27590,N_27009);
xnor U27866 (N_27866,N_27440,N_26546);
xnor U27867 (N_27867,N_27123,N_26631);
nand U27868 (N_27868,N_27120,N_27332);
and U27869 (N_27869,N_27222,N_27262);
or U27870 (N_27870,N_27198,N_27485);
xnor U27871 (N_27871,N_26791,N_26995);
xor U27872 (N_27872,N_26765,N_26451);
nor U27873 (N_27873,N_26467,N_27050);
and U27874 (N_27874,N_27167,N_27425);
or U27875 (N_27875,N_27594,N_27283);
nor U27876 (N_27876,N_26616,N_27215);
nand U27877 (N_27877,N_27076,N_27164);
nor U27878 (N_27878,N_26603,N_27562);
or U27879 (N_27879,N_26989,N_26787);
xor U27880 (N_27880,N_26729,N_27234);
nor U27881 (N_27881,N_27191,N_26544);
and U27882 (N_27882,N_26426,N_26531);
and U27883 (N_27883,N_26809,N_27541);
nand U27884 (N_27884,N_26413,N_27205);
nand U27885 (N_27885,N_26590,N_27523);
nor U27886 (N_27886,N_27518,N_26936);
nand U27887 (N_27887,N_27098,N_27200);
or U27888 (N_27888,N_27210,N_26660);
and U27889 (N_27889,N_27169,N_27319);
and U27890 (N_27890,N_27054,N_26690);
and U27891 (N_27891,N_27484,N_26425);
nand U27892 (N_27892,N_27180,N_26931);
and U27893 (N_27893,N_27231,N_27005);
nor U27894 (N_27894,N_27558,N_27273);
or U27895 (N_27895,N_26668,N_27397);
nand U27896 (N_27896,N_27589,N_26570);
or U27897 (N_27897,N_26944,N_26613);
xor U27898 (N_27898,N_26494,N_26535);
nor U27899 (N_27899,N_26583,N_27471);
nor U27900 (N_27900,N_27335,N_26481);
nand U27901 (N_27901,N_26916,N_27328);
xnor U27902 (N_27902,N_26738,N_27286);
nand U27903 (N_27903,N_27511,N_26522);
nor U27904 (N_27904,N_27577,N_26762);
xnor U27905 (N_27905,N_27449,N_26715);
nand U27906 (N_27906,N_26500,N_26487);
nor U27907 (N_27907,N_26599,N_26848);
or U27908 (N_27908,N_27062,N_27206);
and U27909 (N_27909,N_26596,N_26724);
nor U27910 (N_27910,N_26695,N_27342);
nor U27911 (N_27911,N_27431,N_26702);
or U27912 (N_27912,N_26842,N_26892);
and U27913 (N_27913,N_27495,N_27269);
nand U27914 (N_27914,N_26932,N_26850);
or U27915 (N_27915,N_27306,N_27582);
or U27916 (N_27916,N_27189,N_26430);
or U27917 (N_27917,N_27417,N_27338);
xor U27918 (N_27918,N_26489,N_27149);
xor U27919 (N_27919,N_27004,N_27223);
and U27920 (N_27920,N_26943,N_26731);
nor U27921 (N_27921,N_27293,N_26469);
and U27922 (N_27922,N_27008,N_26973);
or U27923 (N_27923,N_26465,N_27039);
or U27924 (N_27924,N_26552,N_26785);
xor U27925 (N_27925,N_27271,N_26622);
xnor U27926 (N_27926,N_27074,N_26484);
or U27927 (N_27927,N_26509,N_27144);
nor U27928 (N_27928,N_26862,N_27112);
or U27929 (N_27929,N_26629,N_27359);
or U27930 (N_27930,N_27287,N_27221);
xor U27931 (N_27931,N_26748,N_26874);
nand U27932 (N_27932,N_26769,N_26856);
and U27933 (N_27933,N_27175,N_26640);
nor U27934 (N_27934,N_27303,N_26923);
nand U27935 (N_27935,N_26427,N_26672);
xnor U27936 (N_27936,N_26713,N_26917);
and U27937 (N_27937,N_26514,N_26635);
or U27938 (N_27938,N_26682,N_26663);
and U27939 (N_27939,N_26646,N_27515);
nor U27940 (N_27940,N_27363,N_27242);
or U27941 (N_27941,N_26684,N_27365);
and U27942 (N_27942,N_26913,N_27023);
and U27943 (N_27943,N_27252,N_26972);
or U27944 (N_27944,N_27341,N_27318);
or U27945 (N_27945,N_26813,N_26483);
xor U27946 (N_27946,N_26550,N_26466);
nand U27947 (N_27947,N_26752,N_27057);
xor U27948 (N_27948,N_27483,N_26886);
or U27949 (N_27949,N_27571,N_27377);
or U27950 (N_27950,N_27368,N_26634);
xor U27951 (N_27951,N_27395,N_27113);
nand U27952 (N_27952,N_27534,N_26935);
nand U27953 (N_27953,N_27295,N_27390);
and U27954 (N_27954,N_26796,N_26942);
or U27955 (N_27955,N_26865,N_27557);
nand U27956 (N_27956,N_26641,N_26447);
nand U27957 (N_27957,N_26677,N_26934);
nand U27958 (N_27958,N_27419,N_27583);
or U27959 (N_27959,N_26946,N_26416);
nor U27960 (N_27960,N_26882,N_26643);
or U27961 (N_27961,N_27423,N_27251);
or U27962 (N_27962,N_26767,N_26443);
or U27963 (N_27963,N_27476,N_27505);
or U27964 (N_27964,N_27081,N_26548);
nand U27965 (N_27965,N_26821,N_26938);
nand U27966 (N_27966,N_26477,N_26516);
and U27967 (N_27967,N_27422,N_27002);
nand U27968 (N_27968,N_27593,N_27099);
or U27969 (N_27969,N_27161,N_26657);
nor U27970 (N_27970,N_26908,N_27284);
nor U27971 (N_27971,N_26633,N_26446);
or U27972 (N_27972,N_27141,N_27334);
nand U27973 (N_27973,N_27028,N_27032);
nor U27974 (N_27974,N_26464,N_27598);
and U27975 (N_27975,N_27100,N_27366);
nand U27976 (N_27976,N_27400,N_26840);
and U27977 (N_27977,N_26579,N_26401);
nand U27978 (N_27978,N_26754,N_26450);
nor U27979 (N_27979,N_26833,N_26667);
nand U27980 (N_27980,N_26812,N_27458);
nand U27981 (N_27981,N_26716,N_27220);
xnor U27982 (N_27982,N_27043,N_26705);
and U27983 (N_27983,N_26743,N_27072);
or U27984 (N_27984,N_26561,N_27049);
nand U27985 (N_27985,N_27597,N_26536);
nor U27986 (N_27986,N_27246,N_26687);
nor U27987 (N_27987,N_26617,N_27108);
or U27988 (N_27988,N_26834,N_27394);
xnor U27989 (N_27989,N_26676,N_26709);
xnor U27990 (N_27990,N_27451,N_26449);
nor U27991 (N_27991,N_26736,N_26653);
nand U27992 (N_27992,N_27195,N_27361);
nand U27993 (N_27993,N_26518,N_27263);
nand U27994 (N_27994,N_27453,N_27131);
or U27995 (N_27995,N_26598,N_27288);
nand U27996 (N_27996,N_26718,N_26839);
and U27997 (N_27997,N_27313,N_26864);
and U27998 (N_27998,N_27013,N_27496);
nand U27999 (N_27999,N_27048,N_27017);
nand U28000 (N_28000,N_26532,N_27278);
or U28001 (N_28001,N_26918,N_27000);
or U28002 (N_28002,N_26866,N_27526);
xnor U28003 (N_28003,N_26797,N_27038);
xnor U28004 (N_28004,N_27296,N_26869);
and U28005 (N_28005,N_27528,N_27298);
xnor U28006 (N_28006,N_26900,N_26830);
xnor U28007 (N_28007,N_26708,N_27274);
xor U28008 (N_28008,N_27532,N_26490);
nor U28009 (N_28009,N_27507,N_26473);
nor U28010 (N_28010,N_26790,N_26479);
and U28011 (N_28011,N_27550,N_26476);
and U28012 (N_28012,N_26861,N_26929);
nor U28013 (N_28013,N_26597,N_26824);
nand U28014 (N_28014,N_27241,N_27150);
xor U28015 (N_28015,N_27340,N_26648);
and U28016 (N_28016,N_26422,N_26880);
or U28017 (N_28017,N_26565,N_26922);
xnor U28018 (N_28018,N_27486,N_26783);
or U28019 (N_28019,N_26799,N_27323);
nor U28020 (N_28020,N_27304,N_26795);
or U28021 (N_28021,N_27026,N_26956);
and U28022 (N_28022,N_27204,N_26620);
nor U28023 (N_28023,N_27239,N_26564);
nor U28024 (N_28024,N_26823,N_26440);
nand U28025 (N_28025,N_26742,N_27248);
xnor U28026 (N_28026,N_27058,N_27337);
and U28027 (N_28027,N_26976,N_27563);
and U28028 (N_28028,N_26400,N_26927);
nor U28029 (N_28029,N_27244,N_27375);
or U28030 (N_28030,N_26726,N_27159);
nand U28031 (N_28031,N_27482,N_27470);
nand U28032 (N_28032,N_27326,N_26808);
or U28033 (N_28033,N_26524,N_26453);
or U28034 (N_28034,N_27084,N_27114);
xor U28035 (N_28035,N_27176,N_26740);
nor U28036 (N_28036,N_27165,N_26455);
and U28037 (N_28037,N_26513,N_26560);
or U28038 (N_28038,N_26699,N_26928);
nand U28039 (N_28039,N_27442,N_26873);
nand U28040 (N_28040,N_26950,N_26952);
nand U28041 (N_28041,N_27073,N_27468);
nand U28042 (N_28042,N_26470,N_27493);
xor U28043 (N_28043,N_26733,N_26619);
nand U28044 (N_28044,N_26409,N_26694);
xor U28045 (N_28045,N_27385,N_26587);
nor U28046 (N_28046,N_26909,N_27379);
nand U28047 (N_28047,N_27524,N_27085);
nand U28048 (N_28048,N_27279,N_26836);
or U28049 (N_28049,N_27249,N_27586);
xor U28050 (N_28050,N_26728,N_26910);
xnor U28051 (N_28051,N_27424,N_26580);
nand U28052 (N_28052,N_27439,N_27022);
xor U28053 (N_28053,N_26623,N_26507);
or U28054 (N_28054,N_26766,N_27129);
nor U28055 (N_28055,N_27243,N_26593);
xnor U28056 (N_28056,N_26953,N_26838);
nor U28057 (N_28057,N_26595,N_26533);
or U28058 (N_28058,N_26523,N_27265);
and U28059 (N_28059,N_27067,N_27460);
nand U28060 (N_28060,N_27403,N_27499);
nand U28061 (N_28061,N_26814,N_27350);
nand U28062 (N_28062,N_26458,N_26893);
nor U28063 (N_28063,N_26412,N_27018);
nand U28064 (N_28064,N_26819,N_27393);
nand U28065 (N_28065,N_26735,N_26618);
nand U28066 (N_28066,N_27530,N_27237);
and U28067 (N_28067,N_27230,N_27254);
and U28068 (N_28068,N_27509,N_26656);
nor U28069 (N_28069,N_27184,N_27354);
or U28070 (N_28070,N_27565,N_26460);
nand U28071 (N_28071,N_26904,N_26739);
nand U28072 (N_28072,N_26589,N_27349);
and U28073 (N_28073,N_27056,N_27197);
xnor U28074 (N_28074,N_26415,N_26655);
nand U28075 (N_28075,N_27255,N_26698);
nor U28076 (N_28076,N_26845,N_27592);
and U28077 (N_28077,N_26802,N_27465);
nand U28078 (N_28078,N_26600,N_27551);
and U28079 (N_28079,N_26429,N_26899);
and U28080 (N_28080,N_26920,N_26846);
xor U28081 (N_28081,N_27201,N_26898);
xnor U28082 (N_28082,N_27209,N_26987);
or U28083 (N_28083,N_27143,N_26983);
xor U28084 (N_28084,N_27320,N_26501);
and U28085 (N_28085,N_26517,N_26541);
and U28086 (N_28086,N_27382,N_26984);
nor U28087 (N_28087,N_26780,N_27115);
xnor U28088 (N_28088,N_26805,N_27015);
and U28089 (N_28089,N_27556,N_26804);
or U28090 (N_28090,N_27398,N_27259);
or U28091 (N_28091,N_27095,N_27291);
xor U28092 (N_28092,N_26448,N_27399);
and U28093 (N_28093,N_27301,N_27450);
nor U28094 (N_28094,N_26591,N_27130);
or U28095 (N_28095,N_27042,N_26527);
nand U28096 (N_28096,N_26919,N_26471);
and U28097 (N_28097,N_27121,N_27272);
nor U28098 (N_28098,N_26615,N_27545);
nand U28099 (N_28099,N_27345,N_26871);
xnor U28100 (N_28100,N_26624,N_26858);
nor U28101 (N_28101,N_27207,N_27034);
xnor U28102 (N_28102,N_27046,N_27086);
nor U28103 (N_28103,N_26407,N_27527);
nand U28104 (N_28104,N_27538,N_27140);
xnor U28105 (N_28105,N_27559,N_27564);
nor U28106 (N_28106,N_26704,N_27216);
xnor U28107 (N_28107,N_26428,N_27229);
or U28108 (N_28108,N_26521,N_27500);
or U28109 (N_28109,N_26605,N_26496);
nor U28110 (N_28110,N_26750,N_26800);
and U28111 (N_28111,N_26582,N_26825);
and U28112 (N_28112,N_26673,N_26577);
or U28113 (N_28113,N_27264,N_26741);
nor U28114 (N_28114,N_26789,N_26567);
xnor U28115 (N_28115,N_27302,N_27187);
xor U28116 (N_28116,N_26678,N_26602);
xor U28117 (N_28117,N_27595,N_27443);
and U28118 (N_28118,N_27344,N_27094);
xnor U28119 (N_28119,N_26644,N_26468);
and U28120 (N_28120,N_26937,N_26607);
nand U28121 (N_28121,N_26452,N_26894);
nand U28122 (N_28122,N_27153,N_26914);
xor U28123 (N_28123,N_26990,N_27037);
nor U28124 (N_28124,N_26817,N_26439);
nand U28125 (N_28125,N_26647,N_27426);
xnor U28126 (N_28126,N_27213,N_27599);
nor U28127 (N_28127,N_27059,N_27339);
nor U28128 (N_28128,N_27575,N_26562);
nor U28129 (N_28129,N_27415,N_27324);
xor U28130 (N_28130,N_27277,N_26462);
or U28131 (N_28131,N_27574,N_27437);
or U28132 (N_28132,N_27358,N_26721);
xor U28133 (N_28133,N_26887,N_26557);
nor U28134 (N_28134,N_27552,N_26537);
nor U28135 (N_28135,N_26852,N_26542);
nor U28136 (N_28136,N_27404,N_27543);
and U28137 (N_28137,N_27075,N_26406);
nand U28138 (N_28138,N_27024,N_26720);
xnor U28139 (N_28139,N_27416,N_26499);
or U28140 (N_28140,N_27357,N_26614);
xor U28141 (N_28141,N_27371,N_27473);
or U28142 (N_28142,N_27118,N_27409);
or U28143 (N_28143,N_27490,N_26408);
nor U28144 (N_28144,N_27256,N_27092);
and U28145 (N_28145,N_27492,N_26662);
xor U28146 (N_28146,N_27025,N_26747);
nor U28147 (N_28147,N_26654,N_27542);
xor U28148 (N_28148,N_26520,N_26405);
nor U28149 (N_28149,N_26719,N_26420);
nor U28150 (N_28150,N_27276,N_27071);
xnor U28151 (N_28151,N_26816,N_27307);
nor U28152 (N_28152,N_27065,N_26572);
and U28153 (N_28153,N_26890,N_27003);
nand U28154 (N_28154,N_26530,N_26746);
or U28155 (N_28155,N_27066,N_27310);
and U28156 (N_28156,N_27544,N_27497);
and U28157 (N_28157,N_26403,N_26506);
or U28158 (N_28158,N_27445,N_27228);
xor U28159 (N_28159,N_26431,N_27281);
and U28160 (N_28160,N_27508,N_26991);
xor U28161 (N_28161,N_27587,N_27561);
nand U28162 (N_28162,N_26664,N_27282);
nand U28163 (N_28163,N_27452,N_26539);
and U28164 (N_28164,N_27172,N_27181);
nor U28165 (N_28165,N_26472,N_27510);
nor U28166 (N_28166,N_26897,N_27388);
or U28167 (N_28167,N_27462,N_26574);
xnor U28168 (N_28168,N_26642,N_27591);
nor U28169 (N_28169,N_27391,N_26749);
and U28170 (N_28170,N_26519,N_27503);
and U28171 (N_28171,N_26903,N_27330);
and U28172 (N_28172,N_27173,N_26636);
and U28173 (N_28173,N_27588,N_27469);
nor U28174 (N_28174,N_26474,N_26696);
and U28175 (N_28175,N_27155,N_27521);
and U28176 (N_28176,N_26610,N_27477);
xor U28177 (N_28177,N_26404,N_26760);
xor U28178 (N_28178,N_26543,N_26545);
nand U28179 (N_28179,N_26954,N_27232);
nor U28180 (N_28180,N_27238,N_26454);
and U28181 (N_28181,N_27327,N_27570);
xor U28182 (N_28182,N_26558,N_27316);
and U28183 (N_28183,N_26637,N_26710);
nand U28184 (N_28184,N_26828,N_26734);
and U28185 (N_28185,N_26632,N_27343);
nand U28186 (N_28186,N_26891,N_27102);
nand U28187 (N_28187,N_26693,N_26628);
nor U28188 (N_28188,N_26515,N_26906);
nor U28189 (N_28189,N_27280,N_26594);
or U28190 (N_28190,N_26855,N_27466);
xor U28191 (N_28191,N_27137,N_27421);
or U28192 (N_28192,N_26885,N_27554);
xnor U28193 (N_28193,N_27520,N_27245);
and U28194 (N_28194,N_26529,N_26652);
xor U28195 (N_28195,N_27392,N_26988);
nor U28196 (N_28196,N_27314,N_26498);
and U28197 (N_28197,N_27414,N_26974);
nand U28198 (N_28198,N_26877,N_26753);
nor U28199 (N_28199,N_26994,N_27136);
nand U28200 (N_28200,N_27112,N_26735);
and U28201 (N_28201,N_26966,N_26506);
or U28202 (N_28202,N_26795,N_26880);
and U28203 (N_28203,N_26790,N_26803);
nand U28204 (N_28204,N_26957,N_26581);
nand U28205 (N_28205,N_26800,N_26577);
xnor U28206 (N_28206,N_26577,N_27058);
nor U28207 (N_28207,N_26640,N_26686);
nand U28208 (N_28208,N_26468,N_27581);
and U28209 (N_28209,N_27551,N_27060);
nor U28210 (N_28210,N_27123,N_27289);
or U28211 (N_28211,N_27359,N_27423);
nand U28212 (N_28212,N_26584,N_27225);
or U28213 (N_28213,N_27246,N_26439);
xor U28214 (N_28214,N_26997,N_27104);
xnor U28215 (N_28215,N_26935,N_26670);
nand U28216 (N_28216,N_27347,N_26999);
or U28217 (N_28217,N_27436,N_26451);
xnor U28218 (N_28218,N_26553,N_26473);
nand U28219 (N_28219,N_26649,N_27345);
and U28220 (N_28220,N_27434,N_27133);
and U28221 (N_28221,N_26572,N_26582);
or U28222 (N_28222,N_27258,N_26658);
nand U28223 (N_28223,N_26957,N_26671);
and U28224 (N_28224,N_26712,N_26417);
xor U28225 (N_28225,N_27000,N_27535);
xnor U28226 (N_28226,N_27296,N_27149);
xor U28227 (N_28227,N_27221,N_26640);
nor U28228 (N_28228,N_27232,N_26450);
and U28229 (N_28229,N_27475,N_26912);
or U28230 (N_28230,N_26493,N_26405);
nor U28231 (N_28231,N_26623,N_27389);
and U28232 (N_28232,N_27138,N_27430);
nand U28233 (N_28233,N_26638,N_26651);
xor U28234 (N_28234,N_27431,N_26785);
and U28235 (N_28235,N_26830,N_26922);
nand U28236 (N_28236,N_27163,N_27504);
nand U28237 (N_28237,N_26703,N_27103);
nor U28238 (N_28238,N_27026,N_27093);
xnor U28239 (N_28239,N_27245,N_27423);
nand U28240 (N_28240,N_26525,N_27150);
xor U28241 (N_28241,N_26744,N_26478);
xor U28242 (N_28242,N_26994,N_26440);
xnor U28243 (N_28243,N_26508,N_27437);
nand U28244 (N_28244,N_27308,N_27019);
xor U28245 (N_28245,N_26723,N_26725);
nor U28246 (N_28246,N_27279,N_26570);
nand U28247 (N_28247,N_26800,N_27281);
nor U28248 (N_28248,N_27452,N_26448);
xor U28249 (N_28249,N_27048,N_26802);
xor U28250 (N_28250,N_26995,N_26991);
nand U28251 (N_28251,N_27393,N_27598);
nor U28252 (N_28252,N_26442,N_27370);
nor U28253 (N_28253,N_26851,N_27582);
nand U28254 (N_28254,N_26561,N_27204);
and U28255 (N_28255,N_26898,N_26430);
nor U28256 (N_28256,N_26509,N_26727);
xor U28257 (N_28257,N_27098,N_27021);
nor U28258 (N_28258,N_27579,N_26438);
nor U28259 (N_28259,N_26827,N_26571);
nand U28260 (N_28260,N_27372,N_26707);
xnor U28261 (N_28261,N_27042,N_26543);
and U28262 (N_28262,N_27134,N_27251);
or U28263 (N_28263,N_26873,N_27047);
nand U28264 (N_28264,N_27475,N_27024);
and U28265 (N_28265,N_27577,N_27525);
and U28266 (N_28266,N_26741,N_27410);
xnor U28267 (N_28267,N_27361,N_27036);
and U28268 (N_28268,N_27344,N_26425);
and U28269 (N_28269,N_27009,N_26632);
xor U28270 (N_28270,N_27356,N_26471);
nor U28271 (N_28271,N_26471,N_27048);
nand U28272 (N_28272,N_27522,N_26964);
nand U28273 (N_28273,N_26528,N_26619);
or U28274 (N_28274,N_26423,N_26910);
or U28275 (N_28275,N_26718,N_26840);
nor U28276 (N_28276,N_26421,N_26951);
and U28277 (N_28277,N_27339,N_27244);
xor U28278 (N_28278,N_27550,N_27250);
xnor U28279 (N_28279,N_27587,N_27566);
nor U28280 (N_28280,N_27589,N_27056);
or U28281 (N_28281,N_26745,N_26880);
nand U28282 (N_28282,N_26701,N_27031);
and U28283 (N_28283,N_26649,N_27175);
nor U28284 (N_28284,N_27363,N_26705);
xnor U28285 (N_28285,N_27426,N_27559);
and U28286 (N_28286,N_27113,N_26534);
xor U28287 (N_28287,N_27531,N_27537);
xor U28288 (N_28288,N_26859,N_27205);
and U28289 (N_28289,N_27329,N_26483);
nor U28290 (N_28290,N_26564,N_27446);
xnor U28291 (N_28291,N_27085,N_27167);
nand U28292 (N_28292,N_26685,N_26893);
nand U28293 (N_28293,N_27228,N_27174);
nor U28294 (N_28294,N_27221,N_27336);
nor U28295 (N_28295,N_26470,N_27278);
nor U28296 (N_28296,N_27012,N_27534);
nand U28297 (N_28297,N_27363,N_26953);
nor U28298 (N_28298,N_27258,N_27112);
and U28299 (N_28299,N_27314,N_27093);
or U28300 (N_28300,N_26887,N_26870);
or U28301 (N_28301,N_27338,N_27202);
or U28302 (N_28302,N_26674,N_26419);
and U28303 (N_28303,N_27280,N_27497);
nor U28304 (N_28304,N_26680,N_26563);
and U28305 (N_28305,N_27356,N_26701);
and U28306 (N_28306,N_26590,N_26513);
xnor U28307 (N_28307,N_27152,N_26403);
or U28308 (N_28308,N_27337,N_27260);
and U28309 (N_28309,N_27497,N_27233);
or U28310 (N_28310,N_26725,N_27025);
nor U28311 (N_28311,N_27538,N_26850);
nor U28312 (N_28312,N_26867,N_26637);
or U28313 (N_28313,N_27435,N_27547);
and U28314 (N_28314,N_26446,N_26852);
xnor U28315 (N_28315,N_27592,N_27225);
or U28316 (N_28316,N_26737,N_26670);
xor U28317 (N_28317,N_27300,N_27598);
nand U28318 (N_28318,N_27163,N_26424);
or U28319 (N_28319,N_27527,N_26762);
nor U28320 (N_28320,N_27179,N_27103);
and U28321 (N_28321,N_26967,N_26913);
and U28322 (N_28322,N_26645,N_26793);
xnor U28323 (N_28323,N_26708,N_27116);
or U28324 (N_28324,N_26468,N_26736);
nor U28325 (N_28325,N_26895,N_26570);
and U28326 (N_28326,N_26992,N_27293);
or U28327 (N_28327,N_27187,N_27400);
and U28328 (N_28328,N_26425,N_26733);
nor U28329 (N_28329,N_26779,N_26491);
nand U28330 (N_28330,N_27200,N_27289);
nor U28331 (N_28331,N_26611,N_26480);
xor U28332 (N_28332,N_27203,N_27182);
xor U28333 (N_28333,N_27504,N_27113);
nor U28334 (N_28334,N_26749,N_26899);
nand U28335 (N_28335,N_26983,N_26802);
xnor U28336 (N_28336,N_26997,N_26409);
and U28337 (N_28337,N_26764,N_27210);
and U28338 (N_28338,N_27287,N_26683);
nand U28339 (N_28339,N_27535,N_27341);
xor U28340 (N_28340,N_27028,N_27316);
xor U28341 (N_28341,N_26695,N_26527);
and U28342 (N_28342,N_26589,N_27408);
and U28343 (N_28343,N_26475,N_26839);
and U28344 (N_28344,N_26409,N_26843);
xnor U28345 (N_28345,N_27214,N_26862);
and U28346 (N_28346,N_27382,N_26688);
or U28347 (N_28347,N_27586,N_27392);
xor U28348 (N_28348,N_27228,N_27258);
and U28349 (N_28349,N_26732,N_26824);
xnor U28350 (N_28350,N_27411,N_26623);
xor U28351 (N_28351,N_26956,N_26483);
nand U28352 (N_28352,N_26873,N_26616);
and U28353 (N_28353,N_27284,N_27351);
and U28354 (N_28354,N_27147,N_27445);
xor U28355 (N_28355,N_27262,N_27250);
nand U28356 (N_28356,N_27052,N_27105);
nand U28357 (N_28357,N_27561,N_27474);
or U28358 (N_28358,N_27258,N_26899);
nand U28359 (N_28359,N_26471,N_26976);
nand U28360 (N_28360,N_26772,N_27042);
xor U28361 (N_28361,N_27128,N_26659);
nand U28362 (N_28362,N_27591,N_27194);
or U28363 (N_28363,N_26662,N_26808);
and U28364 (N_28364,N_27592,N_26708);
nand U28365 (N_28365,N_27277,N_26915);
or U28366 (N_28366,N_27226,N_26815);
nor U28367 (N_28367,N_27451,N_26791);
nand U28368 (N_28368,N_26787,N_27139);
nand U28369 (N_28369,N_27309,N_27384);
and U28370 (N_28370,N_27215,N_27037);
nand U28371 (N_28371,N_27594,N_27312);
nor U28372 (N_28372,N_26816,N_27430);
nor U28373 (N_28373,N_26417,N_26501);
nand U28374 (N_28374,N_27292,N_26529);
and U28375 (N_28375,N_27347,N_27467);
or U28376 (N_28376,N_27305,N_26900);
nand U28377 (N_28377,N_26593,N_26492);
nor U28378 (N_28378,N_26678,N_26621);
xor U28379 (N_28379,N_27528,N_26660);
nand U28380 (N_28380,N_27225,N_27182);
xor U28381 (N_28381,N_27166,N_27043);
xor U28382 (N_28382,N_26547,N_27501);
nor U28383 (N_28383,N_26713,N_27232);
nor U28384 (N_28384,N_27113,N_27168);
nand U28385 (N_28385,N_26988,N_27240);
or U28386 (N_28386,N_26714,N_26678);
or U28387 (N_28387,N_26417,N_26421);
xor U28388 (N_28388,N_26715,N_26925);
nand U28389 (N_28389,N_26406,N_27067);
and U28390 (N_28390,N_27405,N_27565);
xnor U28391 (N_28391,N_27120,N_26567);
nand U28392 (N_28392,N_26948,N_26852);
and U28393 (N_28393,N_27355,N_27300);
xor U28394 (N_28394,N_27028,N_26938);
nand U28395 (N_28395,N_26689,N_26633);
and U28396 (N_28396,N_26773,N_27021);
xnor U28397 (N_28397,N_27220,N_26759);
and U28398 (N_28398,N_26600,N_27359);
nor U28399 (N_28399,N_26953,N_26621);
xor U28400 (N_28400,N_26848,N_26762);
xnor U28401 (N_28401,N_26452,N_26889);
or U28402 (N_28402,N_27165,N_26754);
xnor U28403 (N_28403,N_27449,N_26800);
nor U28404 (N_28404,N_27160,N_27258);
nor U28405 (N_28405,N_27303,N_26978);
nor U28406 (N_28406,N_27085,N_27455);
nand U28407 (N_28407,N_26621,N_27244);
nor U28408 (N_28408,N_27273,N_26873);
nor U28409 (N_28409,N_26587,N_26405);
xnor U28410 (N_28410,N_26881,N_26601);
nor U28411 (N_28411,N_26927,N_27571);
nor U28412 (N_28412,N_26585,N_26965);
nor U28413 (N_28413,N_26989,N_26448);
and U28414 (N_28414,N_26520,N_26751);
or U28415 (N_28415,N_27234,N_27418);
nor U28416 (N_28416,N_27546,N_26479);
nor U28417 (N_28417,N_26575,N_27371);
or U28418 (N_28418,N_26476,N_27542);
and U28419 (N_28419,N_26786,N_27240);
xor U28420 (N_28420,N_26909,N_26448);
or U28421 (N_28421,N_27502,N_27075);
and U28422 (N_28422,N_26840,N_27590);
and U28423 (N_28423,N_26930,N_27304);
and U28424 (N_28424,N_26998,N_27164);
nor U28425 (N_28425,N_26642,N_27552);
nand U28426 (N_28426,N_26956,N_26410);
and U28427 (N_28427,N_26779,N_26724);
nand U28428 (N_28428,N_27592,N_26673);
and U28429 (N_28429,N_27569,N_26709);
nor U28430 (N_28430,N_26570,N_26524);
and U28431 (N_28431,N_26419,N_27482);
nor U28432 (N_28432,N_27584,N_27023);
xor U28433 (N_28433,N_27514,N_26856);
nor U28434 (N_28434,N_27306,N_26632);
and U28435 (N_28435,N_26753,N_27420);
and U28436 (N_28436,N_26672,N_26977);
nand U28437 (N_28437,N_27454,N_26489);
xor U28438 (N_28438,N_27353,N_26468);
nor U28439 (N_28439,N_27144,N_27347);
or U28440 (N_28440,N_27599,N_27252);
or U28441 (N_28441,N_26857,N_27252);
and U28442 (N_28442,N_27553,N_26886);
nor U28443 (N_28443,N_26520,N_26740);
or U28444 (N_28444,N_26993,N_27172);
xor U28445 (N_28445,N_26440,N_26627);
or U28446 (N_28446,N_26653,N_27368);
and U28447 (N_28447,N_26457,N_26745);
or U28448 (N_28448,N_26754,N_26591);
nand U28449 (N_28449,N_27205,N_26953);
nor U28450 (N_28450,N_26847,N_26585);
xnor U28451 (N_28451,N_26427,N_27219);
nand U28452 (N_28452,N_26940,N_26747);
nand U28453 (N_28453,N_27443,N_27369);
and U28454 (N_28454,N_26977,N_27118);
or U28455 (N_28455,N_26607,N_26691);
or U28456 (N_28456,N_27539,N_26674);
nor U28457 (N_28457,N_27252,N_26885);
nor U28458 (N_28458,N_26937,N_27399);
and U28459 (N_28459,N_26489,N_27208);
xnor U28460 (N_28460,N_26566,N_26997);
and U28461 (N_28461,N_26894,N_26747);
nor U28462 (N_28462,N_27586,N_27283);
xnor U28463 (N_28463,N_27437,N_26840);
nor U28464 (N_28464,N_27364,N_26519);
or U28465 (N_28465,N_26488,N_27130);
nor U28466 (N_28466,N_27377,N_27553);
nand U28467 (N_28467,N_26686,N_26671);
and U28468 (N_28468,N_27378,N_27282);
nor U28469 (N_28469,N_27294,N_26904);
xnor U28470 (N_28470,N_26687,N_27332);
xnor U28471 (N_28471,N_26756,N_27113);
or U28472 (N_28472,N_26926,N_26426);
xnor U28473 (N_28473,N_26727,N_26685);
xnor U28474 (N_28474,N_26934,N_27557);
or U28475 (N_28475,N_26855,N_27248);
or U28476 (N_28476,N_27499,N_27006);
xnor U28477 (N_28477,N_27364,N_26441);
nor U28478 (N_28478,N_27412,N_26533);
nor U28479 (N_28479,N_26684,N_26913);
and U28480 (N_28480,N_27416,N_27214);
xnor U28481 (N_28481,N_27228,N_27240);
or U28482 (N_28482,N_27565,N_26966);
nand U28483 (N_28483,N_27593,N_26757);
nand U28484 (N_28484,N_27393,N_26839);
and U28485 (N_28485,N_27173,N_26724);
or U28486 (N_28486,N_26889,N_27137);
nor U28487 (N_28487,N_26417,N_26424);
nand U28488 (N_28488,N_26914,N_26436);
xor U28489 (N_28489,N_26984,N_27570);
and U28490 (N_28490,N_27032,N_26541);
nand U28491 (N_28491,N_27542,N_27193);
and U28492 (N_28492,N_27512,N_27336);
nand U28493 (N_28493,N_26621,N_27086);
xnor U28494 (N_28494,N_26898,N_26887);
nand U28495 (N_28495,N_26825,N_27550);
xor U28496 (N_28496,N_27564,N_27056);
xnor U28497 (N_28497,N_27296,N_27259);
nand U28498 (N_28498,N_27384,N_26476);
xnor U28499 (N_28499,N_26458,N_26798);
nand U28500 (N_28500,N_26580,N_27563);
nor U28501 (N_28501,N_26850,N_26920);
nand U28502 (N_28502,N_27572,N_26982);
nand U28503 (N_28503,N_27525,N_27053);
or U28504 (N_28504,N_27322,N_26668);
xnor U28505 (N_28505,N_27456,N_27479);
or U28506 (N_28506,N_26690,N_26764);
nand U28507 (N_28507,N_27452,N_26813);
or U28508 (N_28508,N_26805,N_26673);
or U28509 (N_28509,N_27081,N_27555);
xnor U28510 (N_28510,N_26838,N_27589);
xor U28511 (N_28511,N_26700,N_27421);
nand U28512 (N_28512,N_26519,N_27241);
and U28513 (N_28513,N_27399,N_27520);
or U28514 (N_28514,N_27025,N_27173);
nor U28515 (N_28515,N_26546,N_26455);
nand U28516 (N_28516,N_26964,N_26863);
or U28517 (N_28517,N_26502,N_26824);
and U28518 (N_28518,N_26422,N_26413);
xnor U28519 (N_28519,N_26535,N_26879);
nor U28520 (N_28520,N_27286,N_27585);
nor U28521 (N_28521,N_26616,N_27586);
or U28522 (N_28522,N_27383,N_26429);
and U28523 (N_28523,N_26890,N_26889);
and U28524 (N_28524,N_26463,N_27462);
nor U28525 (N_28525,N_26850,N_27158);
and U28526 (N_28526,N_26890,N_27475);
or U28527 (N_28527,N_27116,N_26532);
or U28528 (N_28528,N_26675,N_26893);
nand U28529 (N_28529,N_26638,N_26529);
and U28530 (N_28530,N_26585,N_26724);
nor U28531 (N_28531,N_27414,N_26893);
nor U28532 (N_28532,N_26893,N_27256);
xnor U28533 (N_28533,N_26443,N_27591);
nand U28534 (N_28534,N_27426,N_26697);
or U28535 (N_28535,N_26731,N_27110);
nor U28536 (N_28536,N_26591,N_26812);
nand U28537 (N_28537,N_27134,N_26674);
xnor U28538 (N_28538,N_27045,N_26905);
or U28539 (N_28539,N_27409,N_27213);
or U28540 (N_28540,N_26697,N_26821);
and U28541 (N_28541,N_27014,N_26798);
and U28542 (N_28542,N_27344,N_27049);
nand U28543 (N_28543,N_27471,N_26783);
nor U28544 (N_28544,N_27025,N_26912);
nor U28545 (N_28545,N_27127,N_26711);
xnor U28546 (N_28546,N_27161,N_26690);
and U28547 (N_28547,N_27381,N_27564);
and U28548 (N_28548,N_27284,N_26980);
or U28549 (N_28549,N_26913,N_26679);
xnor U28550 (N_28550,N_27555,N_26924);
nand U28551 (N_28551,N_26574,N_26695);
and U28552 (N_28552,N_26487,N_26418);
or U28553 (N_28553,N_26950,N_26527);
xnor U28554 (N_28554,N_26892,N_26492);
or U28555 (N_28555,N_26657,N_27429);
xnor U28556 (N_28556,N_26978,N_27372);
and U28557 (N_28557,N_27118,N_26842);
xnor U28558 (N_28558,N_27249,N_26866);
or U28559 (N_28559,N_27584,N_26878);
or U28560 (N_28560,N_26742,N_27263);
and U28561 (N_28561,N_27048,N_27227);
or U28562 (N_28562,N_26642,N_27121);
or U28563 (N_28563,N_26808,N_27339);
nand U28564 (N_28564,N_27260,N_27329);
xnor U28565 (N_28565,N_27596,N_27586);
nor U28566 (N_28566,N_27419,N_26847);
and U28567 (N_28567,N_26916,N_26774);
or U28568 (N_28568,N_27468,N_26823);
and U28569 (N_28569,N_26521,N_26955);
xor U28570 (N_28570,N_26852,N_27074);
nor U28571 (N_28571,N_26917,N_27027);
and U28572 (N_28572,N_27238,N_27533);
and U28573 (N_28573,N_26760,N_26898);
xnor U28574 (N_28574,N_27349,N_27510);
nand U28575 (N_28575,N_27416,N_26767);
or U28576 (N_28576,N_27152,N_26936);
or U28577 (N_28577,N_27282,N_27324);
xor U28578 (N_28578,N_27410,N_26433);
nand U28579 (N_28579,N_27445,N_27459);
nor U28580 (N_28580,N_27255,N_27086);
xor U28581 (N_28581,N_27145,N_26943);
nand U28582 (N_28582,N_27078,N_27489);
nand U28583 (N_28583,N_26976,N_26743);
or U28584 (N_28584,N_27567,N_27282);
or U28585 (N_28585,N_26828,N_26822);
nand U28586 (N_28586,N_27230,N_26403);
nand U28587 (N_28587,N_27553,N_27069);
nand U28588 (N_28588,N_26625,N_27412);
or U28589 (N_28589,N_26585,N_27345);
xnor U28590 (N_28590,N_27062,N_27566);
xor U28591 (N_28591,N_27106,N_27311);
or U28592 (N_28592,N_26475,N_27288);
nor U28593 (N_28593,N_27442,N_26578);
nor U28594 (N_28594,N_26560,N_26448);
and U28595 (N_28595,N_27109,N_27000);
xor U28596 (N_28596,N_26957,N_26970);
or U28597 (N_28597,N_26436,N_26754);
nand U28598 (N_28598,N_27049,N_27471);
nand U28599 (N_28599,N_26412,N_27168);
nand U28600 (N_28600,N_26463,N_26753);
nand U28601 (N_28601,N_26559,N_26934);
nor U28602 (N_28602,N_26776,N_27417);
or U28603 (N_28603,N_27069,N_27313);
nor U28604 (N_28604,N_26955,N_26573);
nor U28605 (N_28605,N_26715,N_27034);
xor U28606 (N_28606,N_26450,N_26987);
nor U28607 (N_28607,N_26538,N_27475);
xor U28608 (N_28608,N_27370,N_27377);
and U28609 (N_28609,N_26831,N_26996);
and U28610 (N_28610,N_26736,N_26561);
or U28611 (N_28611,N_27546,N_27001);
and U28612 (N_28612,N_27585,N_27141);
xnor U28613 (N_28613,N_27376,N_27000);
nor U28614 (N_28614,N_26951,N_26435);
nor U28615 (N_28615,N_27589,N_27110);
nor U28616 (N_28616,N_27182,N_27242);
or U28617 (N_28617,N_26870,N_26627);
and U28618 (N_28618,N_27507,N_26530);
and U28619 (N_28619,N_27297,N_27147);
and U28620 (N_28620,N_26422,N_27535);
nor U28621 (N_28621,N_27400,N_26750);
or U28622 (N_28622,N_26947,N_27498);
nor U28623 (N_28623,N_27571,N_26892);
nor U28624 (N_28624,N_27209,N_26717);
xnor U28625 (N_28625,N_27148,N_26495);
and U28626 (N_28626,N_26821,N_27166);
nand U28627 (N_28627,N_26730,N_26578);
nor U28628 (N_28628,N_27230,N_27407);
and U28629 (N_28629,N_27085,N_27101);
xor U28630 (N_28630,N_27492,N_27315);
or U28631 (N_28631,N_26654,N_27380);
xor U28632 (N_28632,N_27070,N_26810);
xnor U28633 (N_28633,N_27418,N_26898);
and U28634 (N_28634,N_26911,N_27098);
or U28635 (N_28635,N_27407,N_27494);
nor U28636 (N_28636,N_27180,N_27459);
nor U28637 (N_28637,N_27273,N_26791);
nand U28638 (N_28638,N_26712,N_26687);
xor U28639 (N_28639,N_26510,N_27161);
nor U28640 (N_28640,N_27289,N_27295);
or U28641 (N_28641,N_27460,N_27099);
nor U28642 (N_28642,N_27130,N_27503);
xor U28643 (N_28643,N_26711,N_26850);
and U28644 (N_28644,N_27324,N_26623);
nand U28645 (N_28645,N_26897,N_26952);
or U28646 (N_28646,N_27100,N_26931);
and U28647 (N_28647,N_26512,N_26980);
and U28648 (N_28648,N_26930,N_27280);
nand U28649 (N_28649,N_26416,N_27195);
xnor U28650 (N_28650,N_26572,N_27523);
nor U28651 (N_28651,N_26556,N_26968);
xor U28652 (N_28652,N_27106,N_27459);
or U28653 (N_28653,N_27046,N_27174);
and U28654 (N_28654,N_27281,N_27004);
and U28655 (N_28655,N_26840,N_26516);
nor U28656 (N_28656,N_27069,N_27289);
nand U28657 (N_28657,N_27510,N_26758);
or U28658 (N_28658,N_26929,N_26426);
or U28659 (N_28659,N_27301,N_27261);
or U28660 (N_28660,N_26799,N_26844);
nor U28661 (N_28661,N_26804,N_27454);
and U28662 (N_28662,N_26479,N_27509);
and U28663 (N_28663,N_26967,N_26836);
nand U28664 (N_28664,N_27400,N_27551);
and U28665 (N_28665,N_26695,N_26819);
nor U28666 (N_28666,N_26791,N_27285);
and U28667 (N_28667,N_26594,N_26778);
nand U28668 (N_28668,N_27135,N_26989);
and U28669 (N_28669,N_27474,N_26890);
nor U28670 (N_28670,N_26667,N_26791);
xor U28671 (N_28671,N_27418,N_27498);
nor U28672 (N_28672,N_26688,N_26669);
nor U28673 (N_28673,N_26953,N_27283);
or U28674 (N_28674,N_26456,N_27446);
xor U28675 (N_28675,N_26938,N_26735);
xor U28676 (N_28676,N_27417,N_26603);
or U28677 (N_28677,N_26747,N_26848);
nor U28678 (N_28678,N_27499,N_26751);
nand U28679 (N_28679,N_26516,N_27060);
and U28680 (N_28680,N_26718,N_27035);
nor U28681 (N_28681,N_26655,N_26982);
nor U28682 (N_28682,N_27229,N_26707);
or U28683 (N_28683,N_26751,N_26578);
nor U28684 (N_28684,N_27083,N_26402);
xor U28685 (N_28685,N_26927,N_27417);
or U28686 (N_28686,N_27286,N_26978);
nor U28687 (N_28687,N_26605,N_27328);
xnor U28688 (N_28688,N_26762,N_27503);
and U28689 (N_28689,N_26401,N_27563);
and U28690 (N_28690,N_27066,N_27326);
and U28691 (N_28691,N_27044,N_26970);
nand U28692 (N_28692,N_26594,N_27164);
and U28693 (N_28693,N_26556,N_27452);
and U28694 (N_28694,N_26834,N_27214);
or U28695 (N_28695,N_27147,N_27158);
nand U28696 (N_28696,N_26885,N_27597);
or U28697 (N_28697,N_27450,N_26403);
and U28698 (N_28698,N_27195,N_26588);
xnor U28699 (N_28699,N_26843,N_27244);
xnor U28700 (N_28700,N_27376,N_26963);
and U28701 (N_28701,N_27327,N_26494);
nand U28702 (N_28702,N_26401,N_26915);
and U28703 (N_28703,N_27105,N_26593);
nor U28704 (N_28704,N_27469,N_26906);
nand U28705 (N_28705,N_27387,N_26445);
and U28706 (N_28706,N_26846,N_27157);
or U28707 (N_28707,N_26694,N_27243);
nand U28708 (N_28708,N_26778,N_27554);
and U28709 (N_28709,N_26463,N_26811);
nor U28710 (N_28710,N_26545,N_27351);
or U28711 (N_28711,N_27307,N_26616);
and U28712 (N_28712,N_27423,N_27597);
nand U28713 (N_28713,N_26848,N_27219);
nand U28714 (N_28714,N_26403,N_26766);
xnor U28715 (N_28715,N_26725,N_26748);
nor U28716 (N_28716,N_27543,N_27107);
or U28717 (N_28717,N_26654,N_26768);
and U28718 (N_28718,N_26855,N_27370);
and U28719 (N_28719,N_26904,N_26576);
nor U28720 (N_28720,N_27590,N_26628);
xnor U28721 (N_28721,N_26603,N_26960);
and U28722 (N_28722,N_26821,N_27077);
nor U28723 (N_28723,N_26741,N_26816);
nand U28724 (N_28724,N_27195,N_26744);
nor U28725 (N_28725,N_26592,N_27242);
nor U28726 (N_28726,N_26432,N_27527);
nor U28727 (N_28727,N_27243,N_26642);
nor U28728 (N_28728,N_26607,N_27353);
and U28729 (N_28729,N_27562,N_27388);
and U28730 (N_28730,N_26834,N_26865);
and U28731 (N_28731,N_27197,N_27502);
nor U28732 (N_28732,N_26979,N_26873);
or U28733 (N_28733,N_27527,N_26586);
nand U28734 (N_28734,N_27086,N_27402);
nand U28735 (N_28735,N_27194,N_27532);
or U28736 (N_28736,N_26873,N_27320);
and U28737 (N_28737,N_27034,N_26957);
nor U28738 (N_28738,N_27315,N_26478);
or U28739 (N_28739,N_26646,N_27040);
xor U28740 (N_28740,N_26862,N_27154);
and U28741 (N_28741,N_27205,N_26717);
nor U28742 (N_28742,N_26602,N_27059);
and U28743 (N_28743,N_27233,N_26521);
xnor U28744 (N_28744,N_26659,N_26486);
or U28745 (N_28745,N_27060,N_26698);
or U28746 (N_28746,N_27374,N_26880);
nor U28747 (N_28747,N_27097,N_26429);
nor U28748 (N_28748,N_27217,N_26512);
and U28749 (N_28749,N_26979,N_27443);
nor U28750 (N_28750,N_27264,N_27167);
nand U28751 (N_28751,N_27395,N_27433);
nand U28752 (N_28752,N_27594,N_26615);
and U28753 (N_28753,N_26796,N_27359);
nand U28754 (N_28754,N_26718,N_27242);
nor U28755 (N_28755,N_26645,N_27447);
nand U28756 (N_28756,N_27185,N_27422);
or U28757 (N_28757,N_27104,N_27484);
xnor U28758 (N_28758,N_26911,N_26729);
xor U28759 (N_28759,N_27183,N_27109);
nand U28760 (N_28760,N_26557,N_26830);
and U28761 (N_28761,N_27036,N_26859);
xor U28762 (N_28762,N_26573,N_27340);
nand U28763 (N_28763,N_27501,N_27096);
and U28764 (N_28764,N_26556,N_26880);
nand U28765 (N_28765,N_27469,N_27113);
nor U28766 (N_28766,N_26558,N_26735);
nor U28767 (N_28767,N_26788,N_26849);
nor U28768 (N_28768,N_26628,N_27532);
nor U28769 (N_28769,N_26763,N_26471);
nand U28770 (N_28770,N_26848,N_27563);
or U28771 (N_28771,N_26519,N_27177);
nand U28772 (N_28772,N_26511,N_27376);
and U28773 (N_28773,N_26534,N_26897);
nand U28774 (N_28774,N_27193,N_26479);
xnor U28775 (N_28775,N_26561,N_26753);
nor U28776 (N_28776,N_26847,N_27581);
nor U28777 (N_28777,N_27127,N_27431);
xnor U28778 (N_28778,N_26483,N_26746);
xor U28779 (N_28779,N_26975,N_27476);
or U28780 (N_28780,N_26765,N_27357);
xor U28781 (N_28781,N_26841,N_26809);
or U28782 (N_28782,N_27423,N_27350);
nand U28783 (N_28783,N_27365,N_27182);
xor U28784 (N_28784,N_26915,N_26671);
nor U28785 (N_28785,N_26902,N_27361);
nand U28786 (N_28786,N_27145,N_26668);
and U28787 (N_28787,N_27485,N_27173);
and U28788 (N_28788,N_26891,N_26750);
nor U28789 (N_28789,N_27394,N_27197);
and U28790 (N_28790,N_26750,N_27394);
and U28791 (N_28791,N_27513,N_26413);
nor U28792 (N_28792,N_26557,N_26921);
and U28793 (N_28793,N_26780,N_27169);
nor U28794 (N_28794,N_26802,N_26544);
and U28795 (N_28795,N_26545,N_26536);
nor U28796 (N_28796,N_26863,N_27159);
nor U28797 (N_28797,N_27583,N_26519);
and U28798 (N_28798,N_26889,N_27011);
nor U28799 (N_28799,N_26870,N_26444);
and U28800 (N_28800,N_27870,N_28504);
nor U28801 (N_28801,N_28724,N_28509);
nor U28802 (N_28802,N_27905,N_27614);
xor U28803 (N_28803,N_28613,N_28384);
nor U28804 (N_28804,N_27824,N_27907);
and U28805 (N_28805,N_28661,N_27897);
nand U28806 (N_28806,N_27840,N_28664);
and U28807 (N_28807,N_28420,N_28428);
or U28808 (N_28808,N_28640,N_28796);
or U28809 (N_28809,N_27657,N_28487);
nor U28810 (N_28810,N_28149,N_28503);
and U28811 (N_28811,N_27927,N_27943);
or U28812 (N_28812,N_27650,N_28175);
nand U28813 (N_28813,N_27857,N_28647);
and U28814 (N_28814,N_28635,N_27851);
and U28815 (N_28815,N_28329,N_27749);
or U28816 (N_28816,N_27909,N_28601);
or U28817 (N_28817,N_28666,N_28489);
and U28818 (N_28818,N_28760,N_28683);
and U28819 (N_28819,N_28399,N_27834);
nand U28820 (N_28820,N_28014,N_28729);
xor U28821 (N_28821,N_27859,N_28153);
nand U28822 (N_28822,N_28270,N_28646);
xor U28823 (N_28823,N_28061,N_27699);
xnor U28824 (N_28824,N_28056,N_28543);
nor U28825 (N_28825,N_28511,N_28449);
nand U28826 (N_28826,N_28387,N_28629);
xor U28827 (N_28827,N_28377,N_28138);
nand U28828 (N_28828,N_28459,N_27773);
and U28829 (N_28829,N_28063,N_28677);
and U28830 (N_28830,N_28461,N_28542);
xnor U28831 (N_28831,N_28260,N_28164);
xnor U28832 (N_28832,N_27663,N_27873);
and U28833 (N_28833,N_28478,N_27777);
nor U28834 (N_28834,N_28572,N_27829);
nand U28835 (N_28835,N_27816,N_27629);
nand U28836 (N_28836,N_28367,N_28722);
nand U28837 (N_28837,N_27640,N_28773);
xor U28838 (N_28838,N_27849,N_28473);
or U28839 (N_28839,N_28077,N_28475);
xor U28840 (N_28840,N_28448,N_28727);
and U28841 (N_28841,N_28158,N_28110);
or U28842 (N_28842,N_28404,N_27940);
and U28843 (N_28843,N_27702,N_28551);
and U28844 (N_28844,N_27884,N_28105);
and U28845 (N_28845,N_27769,N_28049);
nor U28846 (N_28846,N_27692,N_28782);
xnor U28847 (N_28847,N_27715,N_28029);
nor U28848 (N_28848,N_28172,N_27904);
and U28849 (N_28849,N_27659,N_27833);
xnor U28850 (N_28850,N_28240,N_27809);
and U28851 (N_28851,N_27936,N_27838);
or U28852 (N_28852,N_27805,N_28765);
and U28853 (N_28853,N_27881,N_28741);
xnor U28854 (N_28854,N_28257,N_28691);
and U28855 (N_28855,N_28232,N_28290);
nor U28856 (N_28856,N_28292,N_28781);
or U28857 (N_28857,N_27989,N_28332);
and U28858 (N_28858,N_27780,N_28090);
nand U28859 (N_28859,N_27845,N_27995);
nand U28860 (N_28860,N_28253,N_28454);
xor U28861 (N_28861,N_28313,N_28753);
nand U28862 (N_28862,N_28395,N_28467);
nand U28863 (N_28863,N_27795,N_28327);
or U28864 (N_28864,N_27818,N_27768);
nor U28865 (N_28865,N_28492,N_28508);
nand U28866 (N_28866,N_27766,N_28651);
or U28867 (N_28867,N_28092,N_27804);
nor U28868 (N_28868,N_28097,N_28343);
xnor U28869 (N_28869,N_28099,N_28345);
nand U28870 (N_28870,N_27622,N_27690);
nor U28871 (N_28871,N_28565,N_27667);
xor U28872 (N_28872,N_27977,N_28293);
nor U28873 (N_28873,N_28669,N_28177);
and U28874 (N_28874,N_28463,N_28549);
xnor U28875 (N_28875,N_28003,N_28122);
or U28876 (N_28876,N_28389,N_28414);
nand U28877 (N_28877,N_28268,N_27979);
nand U28878 (N_28878,N_28010,N_28366);
and U28879 (N_28879,N_28225,N_28456);
nand U28880 (N_28880,N_27695,N_28062);
nand U28881 (N_28881,N_28198,N_28152);
or U28882 (N_28882,N_28300,N_27661);
nor U28883 (N_28883,N_28445,N_27643);
nor U28884 (N_28884,N_27608,N_28533);
nand U28885 (N_28885,N_28314,N_27826);
or U28886 (N_28886,N_28479,N_27700);
or U28887 (N_28887,N_28307,N_27903);
and U28888 (N_28888,N_28150,N_28402);
nand U28889 (N_28889,N_28556,N_28440);
xor U28890 (N_28890,N_28562,N_27978);
and U28891 (N_28891,N_28596,N_28560);
nand U28892 (N_28892,N_28318,N_28320);
or U28893 (N_28893,N_28604,N_28712);
nor U28894 (N_28894,N_27815,N_28338);
nand U28895 (N_28895,N_28372,N_28554);
xor U28896 (N_28896,N_27937,N_28221);
nand U28897 (N_28897,N_27616,N_27958);
nor U28898 (N_28898,N_27919,N_28256);
nor U28899 (N_28899,N_28794,N_28631);
nand U28900 (N_28900,N_28047,N_28627);
nor U28901 (N_28901,N_27736,N_27878);
xor U28902 (N_28902,N_28176,N_28133);
nand U28903 (N_28903,N_27609,N_28595);
and U28904 (N_28904,N_28706,N_28248);
nand U28905 (N_28905,N_28227,N_28762);
and U28906 (N_28906,N_28477,N_28183);
or U28907 (N_28907,N_28582,N_28263);
xnor U28908 (N_28908,N_28375,N_28025);
and U28909 (N_28909,N_28184,N_28084);
nor U28910 (N_28910,N_28458,N_27679);
xor U28911 (N_28911,N_28048,N_28797);
xnor U28912 (N_28912,N_27678,N_28380);
nor U28913 (N_28913,N_28472,N_28589);
nand U28914 (N_28914,N_28371,N_28685);
or U28915 (N_28915,N_27868,N_28165);
nor U28916 (N_28916,N_28082,N_28648);
and U28917 (N_28917,N_27645,N_27844);
nand U28918 (N_28918,N_28173,N_27847);
or U28919 (N_28919,N_27987,N_27775);
nor U28920 (N_28920,N_28587,N_27921);
nand U28921 (N_28921,N_28137,N_28787);
nand U28922 (N_28922,N_27632,N_28022);
nand U28923 (N_28923,N_27902,N_28139);
and U28924 (N_28924,N_28548,N_27644);
nand U28925 (N_28925,N_27882,N_27788);
nand U28926 (N_28926,N_27942,N_28308);
and U28927 (N_28927,N_28089,N_28547);
or U28928 (N_28928,N_28255,N_28754);
xor U28929 (N_28929,N_27637,N_28728);
nand U28930 (N_28930,N_28605,N_27660);
nor U28931 (N_28931,N_27993,N_28622);
nand U28932 (N_28932,N_27781,N_28649);
or U28933 (N_28933,N_27717,N_28570);
nor U28934 (N_28934,N_28681,N_28252);
nand U28935 (N_28935,N_27689,N_27801);
or U28936 (N_28936,N_27891,N_27999);
xnor U28937 (N_28937,N_27928,N_27716);
nor U28938 (N_28938,N_28671,N_28378);
nand U28939 (N_28939,N_28316,N_28439);
nand U28940 (N_28940,N_28045,N_28597);
or U28941 (N_28941,N_28333,N_27742);
nand U28942 (N_28942,N_28668,N_28228);
nand U28943 (N_28943,N_28085,N_27725);
nor U28944 (N_28944,N_28740,N_27668);
nor U28945 (N_28945,N_28073,N_27662);
or U28946 (N_28946,N_28659,N_28219);
or U28947 (N_28947,N_28331,N_28296);
nor U28948 (N_28948,N_28058,N_28055);
or U28949 (N_28949,N_28295,N_28438);
and U28950 (N_28950,N_28321,N_27831);
nor U28951 (N_28951,N_28123,N_28732);
and U28952 (N_28952,N_27635,N_28069);
nor U28953 (N_28953,N_28695,N_28767);
nor U28954 (N_28954,N_28455,N_28434);
or U28955 (N_28955,N_28127,N_28534);
nor U28956 (N_28956,N_28027,N_28159);
or U28957 (N_28957,N_28625,N_27710);
nand U28958 (N_28958,N_28720,N_27997);
or U28959 (N_28959,N_28580,N_27743);
nor U28960 (N_28960,N_28746,N_27895);
xor U28961 (N_28961,N_27729,N_28054);
xnor U28962 (N_28962,N_28311,N_28118);
and U28963 (N_28963,N_28262,N_28405);
xnor U28964 (N_28964,N_28744,N_28761);
nor U28965 (N_28965,N_28067,N_28120);
nand U28966 (N_28966,N_28617,N_28381);
xor U28967 (N_28967,N_28349,N_28267);
nand U28968 (N_28968,N_28093,N_28654);
nand U28969 (N_28969,N_28522,N_28491);
nor U28970 (N_28970,N_27855,N_28644);
and U28971 (N_28971,N_27984,N_27797);
xnor U28972 (N_28972,N_27906,N_28297);
and U28973 (N_28973,N_28106,N_28476);
nand U28974 (N_28974,N_28355,N_27794);
and U28975 (N_28975,N_27688,N_27861);
or U28976 (N_28976,N_27938,N_28751);
or U28977 (N_28977,N_28312,N_28168);
nor U28978 (N_28978,N_28694,N_27951);
xor U28979 (N_28979,N_28687,N_28271);
xor U28980 (N_28980,N_27812,N_28189);
and U28981 (N_28981,N_28236,N_27759);
or U28982 (N_28982,N_28600,N_28140);
nand U28983 (N_28983,N_28680,N_28098);
nor U28984 (N_28984,N_28146,N_28030);
nand U28985 (N_28985,N_28305,N_27693);
nand U28986 (N_28986,N_28024,N_27980);
xor U28987 (N_28987,N_28771,N_27606);
nand U28988 (N_28988,N_27955,N_27627);
or U28989 (N_28989,N_28336,N_28566);
xnor U28990 (N_28990,N_27724,N_28230);
and U28991 (N_28991,N_28264,N_27848);
nor U28992 (N_28992,N_28624,N_28663);
nor U28993 (N_28993,N_28702,N_28734);
or U28994 (N_28994,N_28167,N_27704);
nor U28995 (N_28995,N_27968,N_27867);
or U28996 (N_28996,N_28550,N_27875);
xnor U28997 (N_28997,N_27837,N_28507);
and U28998 (N_28998,N_28546,N_28482);
nor U28999 (N_28999,N_28537,N_28209);
or U29000 (N_29000,N_28633,N_28246);
nor U29001 (N_29001,N_28682,N_28493);
nor U29002 (N_29002,N_28460,N_28079);
xor U29003 (N_29003,N_28719,N_28770);
xor U29004 (N_29004,N_28362,N_27723);
nand U29005 (N_29005,N_28224,N_28116);
nand U29006 (N_29006,N_27711,N_28360);
xnor U29007 (N_29007,N_28501,N_27750);
xnor U29008 (N_29008,N_27648,N_27880);
nand U29009 (N_29009,N_27866,N_28788);
and U29010 (N_29010,N_28718,N_27941);
xor U29011 (N_29011,N_28019,N_28406);
xnor U29012 (N_29012,N_28050,N_27888);
nand U29013 (N_29013,N_28148,N_28057);
nand U29014 (N_29014,N_28287,N_27713);
nor U29015 (N_29015,N_28160,N_28278);
or U29016 (N_29016,N_28711,N_27877);
or U29017 (N_29017,N_28128,N_28361);
xor U29018 (N_29018,N_28608,N_27754);
nand U29019 (N_29019,N_28621,N_28188);
xor U29020 (N_29020,N_28407,N_28131);
nand U29021 (N_29021,N_28016,N_27944);
nand U29022 (N_29022,N_27952,N_28298);
or U29023 (N_29023,N_28238,N_28656);
nor U29024 (N_29024,N_28390,N_27820);
or U29025 (N_29025,N_27746,N_28576);
or U29026 (N_29026,N_28759,N_28632);
xnor U29027 (N_29027,N_27915,N_28408);
or U29028 (N_29028,N_27654,N_28514);
and U29029 (N_29029,N_28202,N_27854);
and U29030 (N_29030,N_27747,N_28041);
nor U29031 (N_29031,N_27929,N_28036);
nor U29032 (N_29032,N_28039,N_27740);
and U29033 (N_29033,N_28452,N_27974);
nand U29034 (N_29034,N_28005,N_28721);
nand U29035 (N_29035,N_27651,N_27959);
xor U29036 (N_29036,N_28330,N_27810);
nand U29037 (N_29037,N_28700,N_28777);
nor U29038 (N_29038,N_28675,N_27842);
and U29039 (N_29039,N_28279,N_27862);
and U29040 (N_29040,N_28657,N_28713);
and U29041 (N_29041,N_28552,N_28265);
nor U29042 (N_29042,N_27619,N_28690);
nand U29043 (N_29043,N_28409,N_28142);
and U29044 (N_29044,N_28614,N_28525);
or U29045 (N_29045,N_28334,N_27760);
xor U29046 (N_29046,N_28778,N_28358);
and U29047 (N_29047,N_27735,N_27680);
or U29048 (N_29048,N_28353,N_27696);
nor U29049 (N_29049,N_28784,N_27835);
or U29050 (N_29050,N_27966,N_27767);
nor U29051 (N_29051,N_28021,N_27954);
and U29052 (N_29052,N_28171,N_28400);
nor U29053 (N_29053,N_27634,N_28394);
or U29054 (N_29054,N_28516,N_28786);
and U29055 (N_29055,N_27791,N_27939);
and U29056 (N_29056,N_27892,N_28103);
and U29057 (N_29057,N_27603,N_28203);
and U29058 (N_29058,N_28433,N_28348);
or U29059 (N_29059,N_28688,N_28347);
nor U29060 (N_29060,N_28444,N_28446);
nor U29061 (N_29061,N_27967,N_28524);
or U29062 (N_29062,N_28009,N_28650);
and U29063 (N_29063,N_28506,N_28040);
and U29064 (N_29064,N_28337,N_28785);
xnor U29065 (N_29065,N_27806,N_27910);
xnor U29066 (N_29066,N_27817,N_27613);
xnor U29067 (N_29067,N_28234,N_28363);
xor U29068 (N_29068,N_28065,N_27828);
nand U29069 (N_29069,N_28519,N_28497);
or U29070 (N_29070,N_27789,N_28679);
and U29071 (N_29071,N_28261,N_28204);
or U29072 (N_29072,N_27807,N_27879);
nand U29073 (N_29073,N_28350,N_28151);
or U29074 (N_29074,N_28113,N_27626);
nor U29075 (N_29075,N_28156,N_27719);
or U29076 (N_29076,N_28276,N_27790);
nand U29077 (N_29077,N_28386,N_27886);
nand U29078 (N_29078,N_28415,N_27658);
and U29079 (N_29079,N_28447,N_27948);
or U29080 (N_29080,N_28779,N_28764);
xnor U29081 (N_29081,N_28726,N_28294);
nand U29082 (N_29082,N_27822,N_28170);
and U29083 (N_29083,N_28699,N_27639);
xnor U29084 (N_29084,N_28563,N_28523);
or U29085 (N_29085,N_28707,N_28214);
and U29086 (N_29086,N_27962,N_27776);
nand U29087 (N_29087,N_28042,N_28291);
nor U29088 (N_29088,N_27786,N_27893);
and U29089 (N_29089,N_27774,N_28239);
and U29090 (N_29090,N_27761,N_28020);
nand U29091 (N_29091,N_27687,N_28017);
or U29092 (N_29092,N_28450,N_28038);
nor U29093 (N_29093,N_27874,N_28145);
nor U29094 (N_29094,N_28569,N_28008);
or U29095 (N_29095,N_28306,N_28403);
or U29096 (N_29096,N_27894,N_28325);
nand U29097 (N_29097,N_28028,N_28574);
nand U29098 (N_29098,N_28639,N_27755);
xor U29099 (N_29099,N_27675,N_28432);
or U29100 (N_29100,N_28465,N_28701);
nand U29101 (N_29101,N_27947,N_28485);
or U29102 (N_29102,N_27839,N_28737);
xor U29103 (N_29103,N_28319,N_28692);
xnor U29104 (N_29104,N_28775,N_27926);
nand U29105 (N_29105,N_28244,N_27996);
nand U29106 (N_29106,N_28317,N_28359);
or U29107 (N_29107,N_27670,N_28101);
nand U29108 (N_29108,N_27686,N_28541);
xor U29109 (N_29109,N_28466,N_27757);
nand U29110 (N_29110,N_27738,N_28015);
xnor U29111 (N_29111,N_28364,N_28286);
and U29112 (N_29112,N_27808,N_28354);
nor U29113 (N_29113,N_28231,N_27932);
nand U29114 (N_29114,N_28792,N_28626);
nor U29115 (N_29115,N_28108,N_28174);
and U29116 (N_29116,N_27985,N_28095);
nand U29117 (N_29117,N_28419,N_28559);
xnor U29118 (N_29118,N_28072,N_28588);
nand U29119 (N_29119,N_27751,N_27796);
xnor U29120 (N_29120,N_28495,N_27771);
nand U29121 (N_29121,N_28324,N_28119);
nor U29122 (N_29122,N_28068,N_28735);
nand U29123 (N_29123,N_28610,N_28284);
or U29124 (N_29124,N_27744,N_28370);
and U29125 (N_29125,N_28299,N_27602);
nand U29126 (N_29126,N_28579,N_28612);
or U29127 (N_29127,N_27956,N_27722);
and U29128 (N_29128,N_27672,N_28141);
nor U29129 (N_29129,N_28289,N_28592);
nor U29130 (N_29130,N_27961,N_28422);
or U29131 (N_29131,N_27832,N_28081);
nor U29132 (N_29132,N_28532,N_28273);
xnor U29133 (N_29133,N_28277,N_28206);
nor U29134 (N_29134,N_28684,N_27728);
nand U29135 (N_29135,N_28584,N_28107);
and U29136 (N_29136,N_27707,N_28705);
nor U29137 (N_29137,N_27908,N_28529);
nand U29138 (N_29138,N_28346,N_27841);
nand U29139 (N_29139,N_28443,N_28453);
xor U29140 (N_29140,N_28637,N_28396);
nor U29141 (N_29141,N_28667,N_28531);
nand U29142 (N_29142,N_27714,N_28615);
and U29143 (N_29143,N_28033,N_27930);
nand U29144 (N_29144,N_27988,N_28540);
or U29145 (N_29145,N_27630,N_27933);
nand U29146 (N_29146,N_27949,N_28638);
or U29147 (N_29147,N_28673,N_28620);
nor U29148 (N_29148,N_27901,N_27918);
or U29149 (N_29149,N_28623,N_28544);
nor U29150 (N_29150,N_27986,N_28076);
and U29151 (N_29151,N_27981,N_28192);
nand U29152 (N_29152,N_28205,N_27653);
nand U29153 (N_29153,N_28288,N_28066);
and U29154 (N_29154,N_28530,N_27813);
nor U29155 (N_29155,N_28104,N_27727);
nor U29156 (N_29156,N_28498,N_28074);
nor U29157 (N_29157,N_28335,N_27684);
and U29158 (N_29158,N_27682,N_28512);
xor U29159 (N_29159,N_28616,N_28742);
xor U29160 (N_29160,N_28147,N_28745);
xnor U29161 (N_29161,N_27946,N_27957);
nor U29162 (N_29162,N_28609,N_27628);
or U29163 (N_29163,N_28000,N_27655);
xor U29164 (N_29164,N_28383,N_28653);
or U29165 (N_29165,N_28490,N_28630);
xnor U29166 (N_29166,N_28769,N_28750);
nand U29167 (N_29167,N_28179,N_28266);
or U29168 (N_29168,N_28739,N_28725);
nor U29169 (N_29169,N_28578,N_27764);
and U29170 (N_29170,N_28303,N_28006);
nor U29171 (N_29171,N_28094,N_27890);
and U29172 (N_29172,N_28032,N_27992);
or U29173 (N_29173,N_27708,N_27853);
xor U29174 (N_29174,N_27726,N_27638);
nand U29175 (N_29175,N_27681,N_28323);
and U29176 (N_29176,N_28583,N_28553);
xnor U29177 (N_29177,N_28708,N_27610);
nand U29178 (N_29178,N_28195,N_27647);
nor U29179 (N_29179,N_28714,N_27782);
nand U29180 (N_29180,N_27922,N_28393);
or U29181 (N_29181,N_28568,N_27636);
nand U29182 (N_29182,N_28237,N_28674);
or U29183 (N_29183,N_27964,N_28114);
nor U29184 (N_29184,N_28696,N_27931);
or U29185 (N_29185,N_28451,N_27912);
or U29186 (N_29186,N_28571,N_27970);
and U29187 (N_29187,N_28199,N_27983);
or U29188 (N_29188,N_28431,N_27718);
xor U29189 (N_29189,N_28643,N_28281);
nor U29190 (N_29190,N_27617,N_27664);
nor U29191 (N_29191,N_28749,N_27683);
xnor U29192 (N_29192,N_28710,N_28539);
nand U29193 (N_29193,N_28689,N_28783);
nand U29194 (N_29194,N_28756,N_27802);
or U29195 (N_29195,N_27863,N_28196);
nor U29196 (N_29196,N_28339,N_27846);
nand U29197 (N_29197,N_28129,N_27913);
or U29198 (N_29198,N_28418,N_28518);
nor U29199 (N_29199,N_28310,N_27739);
nand U29200 (N_29200,N_28703,N_28013);
or U29201 (N_29201,N_28018,N_27914);
and U29202 (N_29202,N_28426,N_28373);
or U29203 (N_29203,N_28411,N_27830);
and U29204 (N_29204,N_28427,N_27803);
xor U29205 (N_29205,N_27994,N_28130);
or U29206 (N_29206,N_28088,N_28037);
xor U29207 (N_29207,N_27973,N_28144);
nor U29208 (N_29208,N_28730,N_28215);
or U29209 (N_29209,N_28193,N_28315);
or U29210 (N_29210,N_27712,N_28111);
nor U29211 (N_29211,N_28070,N_28619);
and U29212 (N_29212,N_27772,N_28468);
xnor U29213 (N_29213,N_28046,N_28747);
xnor U29214 (N_29214,N_27612,N_27623);
or U29215 (N_29215,N_27872,N_28031);
and U29216 (N_29216,N_28247,N_28527);
nand U29217 (N_29217,N_28210,N_28216);
nor U29218 (N_29218,N_28200,N_27770);
xor U29219 (N_29219,N_28220,N_28698);
xnor U29220 (N_29220,N_28471,N_28510);
and U29221 (N_29221,N_28437,N_28011);
xnor U29222 (N_29222,N_28716,N_27756);
and U29223 (N_29223,N_28494,N_27825);
nand U29224 (N_29224,N_27945,N_28382);
nor U29225 (N_29225,N_28258,N_28328);
xnor U29226 (N_29226,N_28241,N_27709);
and U29227 (N_29227,N_28480,N_27969);
nand U29228 (N_29228,N_28717,N_28197);
nand U29229 (N_29229,N_28789,N_28526);
or U29230 (N_29230,N_28567,N_27779);
nor U29231 (N_29231,N_28269,N_28483);
nor U29232 (N_29232,N_27674,N_27911);
xnor U29233 (N_29233,N_27652,N_27827);
nor U29234 (N_29234,N_28564,N_28059);
nand U29235 (N_29235,N_28686,N_28520);
nor U29236 (N_29236,N_27864,N_28233);
xnor U29237 (N_29237,N_28435,N_28182);
xor U29238 (N_29238,N_28505,N_28259);
and U29239 (N_29239,N_28774,N_27889);
nand U29240 (N_29240,N_28416,N_28154);
nand U29241 (N_29241,N_27963,N_28190);
nor U29242 (N_29242,N_28581,N_28161);
nand U29243 (N_29243,N_28577,N_28723);
and U29244 (N_29244,N_28376,N_27856);
nand U29245 (N_29245,N_28136,N_28528);
xnor U29246 (N_29246,N_28342,N_28251);
nand U29247 (N_29247,N_28155,N_27656);
nand U29248 (N_29248,N_27646,N_27852);
xnor U29249 (N_29249,N_28002,N_27685);
nor U29250 (N_29250,N_28704,N_28590);
xor U29251 (N_29251,N_28007,N_27720);
and U29252 (N_29252,N_28469,N_27666);
xnor U29253 (N_29253,N_28423,N_28515);
or U29254 (N_29254,N_28709,N_27998);
nand U29255 (N_29255,N_28162,N_28121);
nand U29256 (N_29256,N_28201,N_28517);
nand U29257 (N_29257,N_28207,N_27896);
xor U29258 (N_29258,N_27982,N_28186);
xnor U29259 (N_29259,N_28178,N_27748);
nand U29260 (N_29260,N_28598,N_28486);
nand U29261 (N_29261,N_28226,N_28628);
xor U29262 (N_29262,N_27850,N_28500);
or U29263 (N_29263,N_27649,N_28272);
nand U29264 (N_29264,N_27621,N_27836);
xor U29265 (N_29265,N_28593,N_27676);
nor U29266 (N_29266,N_28034,N_27631);
nand U29267 (N_29267,N_28341,N_27758);
xor U29268 (N_29268,N_28391,N_28398);
nor U29269 (N_29269,N_28457,N_27843);
and U29270 (N_29270,N_27620,N_28424);
and U29271 (N_29271,N_28245,N_27604);
and U29272 (N_29272,N_28502,N_28185);
and U29273 (N_29273,N_28309,N_28365);
nor U29274 (N_29274,N_28181,N_27721);
nor U29275 (N_29275,N_28743,N_28132);
or U29276 (N_29276,N_27615,N_28344);
and U29277 (N_29277,N_28080,N_27865);
xnor U29278 (N_29278,N_27923,N_28545);
and U29279 (N_29279,N_28274,N_27618);
nor U29280 (N_29280,N_28078,N_28462);
or U29281 (N_29281,N_27697,N_27800);
or U29282 (N_29282,N_27976,N_28096);
xor U29283 (N_29283,N_27899,N_27732);
nand U29284 (N_29284,N_28026,N_27799);
nor U29285 (N_29285,N_28397,N_27787);
or U29286 (N_29286,N_27734,N_28223);
xnor U29287 (N_29287,N_28212,N_28004);
or U29288 (N_29288,N_28060,N_28768);
nand U29289 (N_29289,N_27972,N_28693);
nor U29290 (N_29290,N_28369,N_28755);
and U29291 (N_29291,N_27925,N_28499);
xor U29292 (N_29292,N_28586,N_28793);
and U29293 (N_29293,N_27821,N_28087);
nand U29294 (N_29294,N_28736,N_28618);
and U29295 (N_29295,N_28044,N_27819);
nand U29296 (N_29296,N_27953,N_28351);
nor U29297 (N_29297,N_27763,N_28208);
nand U29298 (N_29298,N_28109,N_27887);
xnor U29299 (N_29299,N_28748,N_28218);
and U29300 (N_29300,N_28421,N_27823);
or U29301 (N_29301,N_28180,N_27858);
xor U29302 (N_29302,N_28429,N_28143);
and U29303 (N_29303,N_28135,N_28023);
or U29304 (N_29304,N_27778,N_28001);
or U29305 (N_29305,N_28388,N_28213);
nand U29306 (N_29306,N_28470,N_28738);
and U29307 (N_29307,N_28634,N_27745);
xnor U29308 (N_29308,N_28573,N_27991);
nand U29309 (N_29309,N_28282,N_28157);
and U29310 (N_29310,N_28464,N_28166);
xor U29311 (N_29311,N_27605,N_27737);
xnor U29312 (N_29312,N_28536,N_28670);
xor U29313 (N_29313,N_28752,N_28322);
xnor U29314 (N_29314,N_28798,N_27611);
or U29315 (N_29315,N_28283,N_27916);
nand U29316 (N_29316,N_27600,N_27965);
nor U29317 (N_29317,N_28697,N_27673);
nand U29318 (N_29318,N_28474,N_27935);
or U29319 (N_29319,N_28254,N_28126);
or U29320 (N_29320,N_27607,N_28557);
nor U29321 (N_29321,N_28585,N_28763);
xor U29322 (N_29322,N_28187,N_28115);
or U29323 (N_29323,N_27814,N_28636);
nor U29324 (N_29324,N_27731,N_27741);
nand U29325 (N_29325,N_28642,N_28012);
xnor U29326 (N_29326,N_27975,N_28425);
and U29327 (N_29327,N_28217,N_28413);
nor U29328 (N_29328,N_28733,N_28496);
nor U29329 (N_29329,N_28356,N_27798);
and U29330 (N_29330,N_28280,N_27885);
and U29331 (N_29331,N_28385,N_27793);
nand U29332 (N_29332,N_28538,N_27785);
xor U29333 (N_29333,N_28758,N_28043);
or U29334 (N_29334,N_27860,N_28780);
and U29335 (N_29335,N_28053,N_27876);
or U29336 (N_29336,N_28194,N_28558);
or U29337 (N_29337,N_27698,N_27898);
nor U29338 (N_29338,N_28655,N_27883);
nand U29339 (N_29339,N_28555,N_27633);
and U29340 (N_29340,N_28591,N_28575);
and U29341 (N_29341,N_27691,N_27730);
nor U29342 (N_29342,N_28513,N_28235);
nor U29343 (N_29343,N_27703,N_28285);
nor U29344 (N_29344,N_28606,N_28117);
or U29345 (N_29345,N_28481,N_27869);
xor U29346 (N_29346,N_28249,N_28672);
or U29347 (N_29347,N_28790,N_27990);
and U29348 (N_29348,N_28124,N_27625);
and U29349 (N_29349,N_28275,N_28250);
or U29350 (N_29350,N_28795,N_28125);
and U29351 (N_29351,N_28222,N_28561);
nand U29352 (N_29352,N_27783,N_27811);
and U29353 (N_29353,N_28658,N_28035);
and U29354 (N_29354,N_28430,N_27669);
nor U29355 (N_29355,N_28086,N_28064);
or U29356 (N_29356,N_27752,N_28607);
and U29357 (N_29357,N_27701,N_27917);
nor U29358 (N_29358,N_28301,N_28191);
and U29359 (N_29359,N_28243,N_27705);
or U29360 (N_29360,N_28083,N_28242);
nand U29361 (N_29361,N_28594,N_28611);
nor U29362 (N_29362,N_28304,N_27871);
and U29363 (N_29363,N_28410,N_28488);
xor U29364 (N_29364,N_28352,N_28102);
and U29365 (N_29365,N_28392,N_27971);
nor U29366 (N_29366,N_27601,N_28100);
or U29367 (N_29367,N_28051,N_27733);
and U29368 (N_29368,N_28521,N_28052);
nor U29369 (N_29369,N_28229,N_27671);
and U29370 (N_29370,N_28112,N_28401);
nor U29371 (N_29371,N_27694,N_28368);
or U29372 (N_29372,N_27960,N_28302);
xor U29373 (N_29373,N_28791,N_28379);
nand U29374 (N_29374,N_27950,N_27624);
nand U29375 (N_29375,N_28436,N_27920);
or U29376 (N_29376,N_27677,N_27924);
nor U29377 (N_29377,N_28641,N_28417);
and U29378 (N_29378,N_28776,N_28134);
nor U29379 (N_29379,N_28075,N_28662);
and U29380 (N_29380,N_28340,N_28678);
nor U29381 (N_29381,N_27753,N_28715);
xnor U29382 (N_29382,N_28169,N_28357);
nor U29383 (N_29383,N_27934,N_28163);
xor U29384 (N_29384,N_27641,N_27792);
nand U29385 (N_29385,N_28599,N_27762);
nor U29386 (N_29386,N_28602,N_27642);
or U29387 (N_29387,N_28071,N_27765);
nor U29388 (N_29388,N_28731,N_27900);
and U29389 (N_29389,N_28645,N_28484);
and U29390 (N_29390,N_28211,N_27665);
nand U29391 (N_29391,N_28676,N_27706);
or U29392 (N_29392,N_28665,N_28442);
and U29393 (N_29393,N_28603,N_27784);
xnor U29394 (N_29394,N_28757,N_28652);
xor U29395 (N_29395,N_28660,N_28091);
xor U29396 (N_29396,N_28412,N_28441);
and U29397 (N_29397,N_28772,N_28766);
nand U29398 (N_29398,N_28326,N_28799);
nand U29399 (N_29399,N_28535,N_28374);
and U29400 (N_29400,N_27781,N_28643);
nor U29401 (N_29401,N_28618,N_28598);
or U29402 (N_29402,N_27957,N_28533);
xnor U29403 (N_29403,N_27905,N_28435);
and U29404 (N_29404,N_27684,N_27657);
xnor U29405 (N_29405,N_28716,N_28574);
and U29406 (N_29406,N_27821,N_28627);
xor U29407 (N_29407,N_28396,N_28061);
nor U29408 (N_29408,N_28072,N_28795);
and U29409 (N_29409,N_28592,N_28053);
nand U29410 (N_29410,N_28345,N_28711);
or U29411 (N_29411,N_28070,N_27663);
nand U29412 (N_29412,N_28613,N_28238);
nand U29413 (N_29413,N_28090,N_27789);
or U29414 (N_29414,N_27786,N_28079);
nand U29415 (N_29415,N_28251,N_28137);
and U29416 (N_29416,N_28689,N_27696);
nand U29417 (N_29417,N_28682,N_27853);
or U29418 (N_29418,N_27950,N_27911);
nand U29419 (N_29419,N_28453,N_28286);
xor U29420 (N_29420,N_28543,N_27700);
and U29421 (N_29421,N_28184,N_27933);
xnor U29422 (N_29422,N_27736,N_27613);
and U29423 (N_29423,N_28220,N_27604);
nor U29424 (N_29424,N_28745,N_28576);
or U29425 (N_29425,N_27814,N_27797);
nor U29426 (N_29426,N_28127,N_28032);
or U29427 (N_29427,N_27792,N_28331);
nand U29428 (N_29428,N_28352,N_27743);
nand U29429 (N_29429,N_28301,N_28651);
nor U29430 (N_29430,N_28316,N_28181);
nand U29431 (N_29431,N_28271,N_28332);
or U29432 (N_29432,N_28278,N_28589);
or U29433 (N_29433,N_28572,N_28063);
and U29434 (N_29434,N_27633,N_27942);
or U29435 (N_29435,N_27855,N_28329);
or U29436 (N_29436,N_28630,N_27697);
nor U29437 (N_29437,N_28259,N_27611);
xnor U29438 (N_29438,N_28372,N_28528);
nor U29439 (N_29439,N_28298,N_28557);
nor U29440 (N_29440,N_28375,N_28109);
and U29441 (N_29441,N_28725,N_28194);
xnor U29442 (N_29442,N_27656,N_28114);
or U29443 (N_29443,N_27953,N_28450);
or U29444 (N_29444,N_28620,N_28699);
and U29445 (N_29445,N_28188,N_27672);
xor U29446 (N_29446,N_27962,N_28154);
or U29447 (N_29447,N_28229,N_27978);
nor U29448 (N_29448,N_27995,N_27773);
or U29449 (N_29449,N_27809,N_28632);
or U29450 (N_29450,N_28627,N_28100);
and U29451 (N_29451,N_28579,N_28716);
and U29452 (N_29452,N_27712,N_28032);
xor U29453 (N_29453,N_27773,N_28151);
nor U29454 (N_29454,N_27969,N_28097);
nand U29455 (N_29455,N_28303,N_28718);
nor U29456 (N_29456,N_27794,N_28476);
and U29457 (N_29457,N_27770,N_28260);
nor U29458 (N_29458,N_27658,N_28343);
nor U29459 (N_29459,N_28607,N_28346);
xnor U29460 (N_29460,N_27750,N_28166);
nor U29461 (N_29461,N_27958,N_28299);
nor U29462 (N_29462,N_28409,N_28695);
nand U29463 (N_29463,N_27896,N_28242);
or U29464 (N_29464,N_27670,N_28381);
and U29465 (N_29465,N_28167,N_27623);
and U29466 (N_29466,N_27940,N_27824);
nor U29467 (N_29467,N_28047,N_28547);
and U29468 (N_29468,N_27988,N_28764);
nor U29469 (N_29469,N_27617,N_28485);
xnor U29470 (N_29470,N_28432,N_27609);
xor U29471 (N_29471,N_28133,N_27895);
nand U29472 (N_29472,N_28310,N_27843);
or U29473 (N_29473,N_27913,N_28673);
nor U29474 (N_29474,N_27888,N_27754);
xor U29475 (N_29475,N_27764,N_27750);
xnor U29476 (N_29476,N_28266,N_27977);
and U29477 (N_29477,N_28623,N_27757);
or U29478 (N_29478,N_28319,N_28717);
nor U29479 (N_29479,N_28653,N_27924);
xor U29480 (N_29480,N_27656,N_28324);
nand U29481 (N_29481,N_28373,N_28544);
nand U29482 (N_29482,N_28369,N_27949);
and U29483 (N_29483,N_27685,N_27840);
nor U29484 (N_29484,N_28218,N_28124);
or U29485 (N_29485,N_27952,N_28746);
or U29486 (N_29486,N_28697,N_28507);
xnor U29487 (N_29487,N_28345,N_28485);
and U29488 (N_29488,N_28501,N_28699);
xor U29489 (N_29489,N_28699,N_28444);
or U29490 (N_29490,N_27952,N_28558);
nand U29491 (N_29491,N_27637,N_27726);
nor U29492 (N_29492,N_28772,N_28604);
or U29493 (N_29493,N_27996,N_28014);
or U29494 (N_29494,N_28132,N_28799);
nand U29495 (N_29495,N_28048,N_28441);
nand U29496 (N_29496,N_28653,N_28376);
and U29497 (N_29497,N_27639,N_28626);
nor U29498 (N_29498,N_28533,N_28105);
xor U29499 (N_29499,N_27716,N_28127);
nand U29500 (N_29500,N_27696,N_28406);
nor U29501 (N_29501,N_28207,N_28404);
nor U29502 (N_29502,N_28706,N_28621);
and U29503 (N_29503,N_28676,N_28169);
or U29504 (N_29504,N_28594,N_28329);
nand U29505 (N_29505,N_28131,N_27643);
nor U29506 (N_29506,N_28098,N_28522);
nand U29507 (N_29507,N_28327,N_28082);
or U29508 (N_29508,N_27691,N_27692);
nor U29509 (N_29509,N_27990,N_28500);
nand U29510 (N_29510,N_28008,N_27612);
nor U29511 (N_29511,N_28602,N_28647);
or U29512 (N_29512,N_27879,N_28752);
nor U29513 (N_29513,N_28428,N_27878);
or U29514 (N_29514,N_28790,N_28333);
or U29515 (N_29515,N_28685,N_27908);
xor U29516 (N_29516,N_27756,N_28472);
or U29517 (N_29517,N_27740,N_28180);
xnor U29518 (N_29518,N_28026,N_28317);
nand U29519 (N_29519,N_27757,N_28383);
or U29520 (N_29520,N_28725,N_28006);
or U29521 (N_29521,N_28436,N_28002);
nand U29522 (N_29522,N_28273,N_28297);
or U29523 (N_29523,N_28085,N_28320);
and U29524 (N_29524,N_27743,N_27600);
nand U29525 (N_29525,N_28271,N_28688);
xnor U29526 (N_29526,N_28398,N_27736);
xor U29527 (N_29527,N_28524,N_27915);
or U29528 (N_29528,N_27691,N_27816);
or U29529 (N_29529,N_28060,N_28305);
nor U29530 (N_29530,N_28274,N_28282);
nor U29531 (N_29531,N_28584,N_27712);
xnor U29532 (N_29532,N_28245,N_28620);
and U29533 (N_29533,N_28665,N_28069);
or U29534 (N_29534,N_28730,N_28768);
and U29535 (N_29535,N_27868,N_27651);
or U29536 (N_29536,N_28066,N_27708);
nand U29537 (N_29537,N_28111,N_27606);
nor U29538 (N_29538,N_28760,N_27944);
nand U29539 (N_29539,N_28453,N_27975);
nand U29540 (N_29540,N_28550,N_28555);
nand U29541 (N_29541,N_28383,N_27775);
nand U29542 (N_29542,N_28638,N_28641);
xor U29543 (N_29543,N_28038,N_27898);
and U29544 (N_29544,N_28597,N_28135);
xnor U29545 (N_29545,N_28230,N_28332);
and U29546 (N_29546,N_28369,N_28031);
xnor U29547 (N_29547,N_28367,N_28470);
or U29548 (N_29548,N_28144,N_28384);
or U29549 (N_29549,N_28306,N_27956);
xor U29550 (N_29550,N_28681,N_28306);
and U29551 (N_29551,N_27789,N_27688);
nor U29552 (N_29552,N_28235,N_27780);
nor U29553 (N_29553,N_28749,N_28338);
or U29554 (N_29554,N_28043,N_28465);
and U29555 (N_29555,N_28491,N_28164);
or U29556 (N_29556,N_28233,N_28542);
nor U29557 (N_29557,N_28162,N_28056);
or U29558 (N_29558,N_27679,N_27977);
xor U29559 (N_29559,N_28471,N_28746);
and U29560 (N_29560,N_27676,N_28785);
or U29561 (N_29561,N_27878,N_28333);
xnor U29562 (N_29562,N_28685,N_28714);
or U29563 (N_29563,N_28044,N_28773);
nand U29564 (N_29564,N_28792,N_28673);
xor U29565 (N_29565,N_28163,N_27961);
nand U29566 (N_29566,N_28084,N_28545);
nor U29567 (N_29567,N_28653,N_27841);
nor U29568 (N_29568,N_27787,N_28200);
nand U29569 (N_29569,N_28005,N_27645);
xor U29570 (N_29570,N_28328,N_28769);
nor U29571 (N_29571,N_28382,N_27980);
nand U29572 (N_29572,N_28147,N_28244);
nand U29573 (N_29573,N_28189,N_28246);
xor U29574 (N_29574,N_27717,N_27740);
nand U29575 (N_29575,N_28423,N_28089);
xnor U29576 (N_29576,N_28427,N_28244);
and U29577 (N_29577,N_28706,N_28776);
and U29578 (N_29578,N_28482,N_28545);
or U29579 (N_29579,N_28323,N_28269);
and U29580 (N_29580,N_28083,N_28363);
nand U29581 (N_29581,N_27789,N_28147);
nor U29582 (N_29582,N_27845,N_27726);
and U29583 (N_29583,N_27913,N_28220);
nor U29584 (N_29584,N_28280,N_28204);
and U29585 (N_29585,N_27638,N_28173);
xor U29586 (N_29586,N_28389,N_28025);
nand U29587 (N_29587,N_28374,N_28493);
or U29588 (N_29588,N_28799,N_28551);
and U29589 (N_29589,N_28481,N_28453);
or U29590 (N_29590,N_27708,N_28634);
and U29591 (N_29591,N_27818,N_27608);
and U29592 (N_29592,N_28600,N_28024);
nor U29593 (N_29593,N_27636,N_28496);
xnor U29594 (N_29594,N_28729,N_28535);
or U29595 (N_29595,N_28498,N_27707);
or U29596 (N_29596,N_27710,N_27683);
or U29597 (N_29597,N_27727,N_28217);
nand U29598 (N_29598,N_27953,N_28688);
or U29599 (N_29599,N_27995,N_27627);
and U29600 (N_29600,N_27664,N_28147);
or U29601 (N_29601,N_27703,N_27809);
and U29602 (N_29602,N_28439,N_27892);
and U29603 (N_29603,N_28191,N_28134);
and U29604 (N_29604,N_27886,N_28277);
and U29605 (N_29605,N_27815,N_27686);
nand U29606 (N_29606,N_27615,N_28470);
nor U29607 (N_29607,N_28601,N_28144);
nand U29608 (N_29608,N_28452,N_27691);
or U29609 (N_29609,N_27970,N_27767);
xor U29610 (N_29610,N_28242,N_27682);
xor U29611 (N_29611,N_28634,N_28136);
nand U29612 (N_29612,N_28686,N_28397);
xor U29613 (N_29613,N_28512,N_28796);
nand U29614 (N_29614,N_28236,N_27911);
xnor U29615 (N_29615,N_28671,N_27799);
or U29616 (N_29616,N_28739,N_28081);
xnor U29617 (N_29617,N_28438,N_27640);
nor U29618 (N_29618,N_28360,N_28647);
or U29619 (N_29619,N_28770,N_28379);
nor U29620 (N_29620,N_28305,N_28725);
or U29621 (N_29621,N_27698,N_28784);
xnor U29622 (N_29622,N_28601,N_28561);
nand U29623 (N_29623,N_28619,N_28393);
xor U29624 (N_29624,N_28326,N_28444);
nand U29625 (N_29625,N_28333,N_28263);
and U29626 (N_29626,N_27817,N_28051);
or U29627 (N_29627,N_27808,N_28096);
nor U29628 (N_29628,N_28639,N_28296);
nor U29629 (N_29629,N_27709,N_28106);
nor U29630 (N_29630,N_27728,N_28326);
nand U29631 (N_29631,N_28024,N_27635);
and U29632 (N_29632,N_28576,N_27805);
nor U29633 (N_29633,N_28780,N_27650);
or U29634 (N_29634,N_28050,N_28437);
xor U29635 (N_29635,N_28779,N_28602);
or U29636 (N_29636,N_28335,N_27907);
nand U29637 (N_29637,N_27753,N_27890);
or U29638 (N_29638,N_28031,N_27979);
nor U29639 (N_29639,N_28647,N_28379);
and U29640 (N_29640,N_27678,N_28415);
nor U29641 (N_29641,N_28625,N_28579);
nor U29642 (N_29642,N_28240,N_28455);
nor U29643 (N_29643,N_28435,N_28737);
nand U29644 (N_29644,N_28222,N_28628);
or U29645 (N_29645,N_28045,N_28486);
xnor U29646 (N_29646,N_28495,N_28015);
xor U29647 (N_29647,N_28721,N_27966);
and U29648 (N_29648,N_27669,N_27839);
nor U29649 (N_29649,N_28762,N_28540);
nand U29650 (N_29650,N_28409,N_27924);
xor U29651 (N_29651,N_27831,N_28734);
and U29652 (N_29652,N_27626,N_28640);
nand U29653 (N_29653,N_28068,N_28312);
or U29654 (N_29654,N_28577,N_27837);
nor U29655 (N_29655,N_27738,N_28698);
nand U29656 (N_29656,N_27895,N_28566);
nor U29657 (N_29657,N_27791,N_27946);
or U29658 (N_29658,N_28142,N_27788);
xnor U29659 (N_29659,N_27608,N_27700);
or U29660 (N_29660,N_28700,N_28417);
nand U29661 (N_29661,N_28131,N_28318);
nand U29662 (N_29662,N_28636,N_28525);
and U29663 (N_29663,N_28182,N_28710);
or U29664 (N_29664,N_28268,N_28571);
nand U29665 (N_29665,N_28084,N_27843);
nor U29666 (N_29666,N_28605,N_28546);
nor U29667 (N_29667,N_28781,N_28101);
nand U29668 (N_29668,N_27838,N_28721);
nor U29669 (N_29669,N_28064,N_28243);
or U29670 (N_29670,N_28043,N_27868);
or U29671 (N_29671,N_28568,N_28204);
nor U29672 (N_29672,N_28763,N_28147);
xnor U29673 (N_29673,N_28382,N_28793);
or U29674 (N_29674,N_28746,N_28000);
nor U29675 (N_29675,N_28339,N_27827);
nand U29676 (N_29676,N_28272,N_27962);
or U29677 (N_29677,N_28419,N_28053);
or U29678 (N_29678,N_28132,N_28133);
nor U29679 (N_29679,N_28161,N_27653);
and U29680 (N_29680,N_28292,N_28183);
xnor U29681 (N_29681,N_27741,N_28187);
nor U29682 (N_29682,N_28574,N_27758);
and U29683 (N_29683,N_28168,N_28758);
and U29684 (N_29684,N_28322,N_27706);
xor U29685 (N_29685,N_28616,N_27852);
nor U29686 (N_29686,N_28343,N_27998);
nand U29687 (N_29687,N_28321,N_27847);
or U29688 (N_29688,N_28137,N_28676);
nand U29689 (N_29689,N_28344,N_27669);
and U29690 (N_29690,N_27657,N_28382);
nand U29691 (N_29691,N_27697,N_27912);
nand U29692 (N_29692,N_28069,N_27627);
nor U29693 (N_29693,N_27665,N_27938);
or U29694 (N_29694,N_28106,N_28519);
nor U29695 (N_29695,N_28505,N_28052);
xnor U29696 (N_29696,N_27801,N_27722);
nand U29697 (N_29697,N_28327,N_28708);
or U29698 (N_29698,N_28726,N_27705);
and U29699 (N_29699,N_27893,N_28048);
or U29700 (N_29700,N_28772,N_28510);
nor U29701 (N_29701,N_28209,N_28325);
or U29702 (N_29702,N_27771,N_28765);
nand U29703 (N_29703,N_27965,N_28141);
xnor U29704 (N_29704,N_28609,N_27818);
nand U29705 (N_29705,N_28035,N_27962);
nor U29706 (N_29706,N_28053,N_27703);
and U29707 (N_29707,N_28071,N_28672);
nor U29708 (N_29708,N_27926,N_28210);
or U29709 (N_29709,N_27895,N_28705);
and U29710 (N_29710,N_28421,N_27836);
and U29711 (N_29711,N_28297,N_28311);
or U29712 (N_29712,N_28620,N_28309);
or U29713 (N_29713,N_27765,N_28415);
or U29714 (N_29714,N_28422,N_27902);
or U29715 (N_29715,N_27617,N_27686);
and U29716 (N_29716,N_27900,N_27895);
xnor U29717 (N_29717,N_27977,N_28493);
or U29718 (N_29718,N_28173,N_28000);
nand U29719 (N_29719,N_27607,N_27647);
or U29720 (N_29720,N_28684,N_28161);
nor U29721 (N_29721,N_28189,N_27621);
or U29722 (N_29722,N_28191,N_28282);
nor U29723 (N_29723,N_27915,N_28579);
nand U29724 (N_29724,N_28798,N_28294);
xnor U29725 (N_29725,N_28361,N_27847);
and U29726 (N_29726,N_28739,N_28385);
nor U29727 (N_29727,N_28207,N_28026);
xor U29728 (N_29728,N_28031,N_27792);
xor U29729 (N_29729,N_28652,N_28787);
nor U29730 (N_29730,N_28667,N_27841);
and U29731 (N_29731,N_28097,N_28458);
xor U29732 (N_29732,N_28632,N_28085);
and U29733 (N_29733,N_28707,N_27951);
nor U29734 (N_29734,N_28439,N_28321);
nor U29735 (N_29735,N_27968,N_28591);
or U29736 (N_29736,N_28142,N_28752);
nand U29737 (N_29737,N_28172,N_28752);
or U29738 (N_29738,N_28541,N_28793);
and U29739 (N_29739,N_27976,N_28064);
nor U29740 (N_29740,N_28473,N_28673);
or U29741 (N_29741,N_27832,N_28375);
nand U29742 (N_29742,N_28564,N_28457);
nand U29743 (N_29743,N_28238,N_28696);
nand U29744 (N_29744,N_28656,N_27715);
nand U29745 (N_29745,N_28186,N_28061);
and U29746 (N_29746,N_27639,N_27975);
and U29747 (N_29747,N_27728,N_27730);
and U29748 (N_29748,N_28000,N_28224);
and U29749 (N_29749,N_27601,N_27972);
nor U29750 (N_29750,N_28071,N_27768);
and U29751 (N_29751,N_27987,N_27934);
xnor U29752 (N_29752,N_27850,N_27834);
and U29753 (N_29753,N_27935,N_27946);
nor U29754 (N_29754,N_28617,N_27657);
or U29755 (N_29755,N_28754,N_28238);
and U29756 (N_29756,N_28174,N_28571);
and U29757 (N_29757,N_28450,N_28630);
and U29758 (N_29758,N_28021,N_27982);
and U29759 (N_29759,N_28070,N_27742);
xor U29760 (N_29760,N_28433,N_27959);
and U29761 (N_29761,N_27626,N_27677);
nand U29762 (N_29762,N_28362,N_27906);
or U29763 (N_29763,N_27625,N_28688);
nand U29764 (N_29764,N_28588,N_28472);
nand U29765 (N_29765,N_28292,N_28342);
nor U29766 (N_29766,N_28402,N_28618);
nor U29767 (N_29767,N_28442,N_27809);
or U29768 (N_29768,N_28038,N_28226);
nand U29769 (N_29769,N_28221,N_28268);
xnor U29770 (N_29770,N_28160,N_28267);
nor U29771 (N_29771,N_28479,N_27744);
nor U29772 (N_29772,N_27985,N_28286);
or U29773 (N_29773,N_28496,N_28057);
nand U29774 (N_29774,N_27723,N_28345);
or U29775 (N_29775,N_28001,N_28204);
and U29776 (N_29776,N_28371,N_28660);
xnor U29777 (N_29777,N_27888,N_27865);
xnor U29778 (N_29778,N_28466,N_27646);
and U29779 (N_29779,N_28736,N_27904);
nand U29780 (N_29780,N_28786,N_27756);
or U29781 (N_29781,N_27690,N_27790);
or U29782 (N_29782,N_28002,N_28777);
xnor U29783 (N_29783,N_27959,N_27696);
nor U29784 (N_29784,N_27730,N_28059);
nand U29785 (N_29785,N_28709,N_27934);
nor U29786 (N_29786,N_27711,N_27673);
nor U29787 (N_29787,N_28679,N_27700);
nor U29788 (N_29788,N_28128,N_28764);
or U29789 (N_29789,N_27959,N_28334);
xor U29790 (N_29790,N_27916,N_27605);
xnor U29791 (N_29791,N_27706,N_28524);
and U29792 (N_29792,N_27961,N_28571);
nand U29793 (N_29793,N_28517,N_28196);
nand U29794 (N_29794,N_28423,N_28273);
xor U29795 (N_29795,N_28194,N_28544);
or U29796 (N_29796,N_27879,N_28442);
nor U29797 (N_29797,N_28178,N_28490);
or U29798 (N_29798,N_27753,N_28527);
xnor U29799 (N_29799,N_28291,N_28543);
nor U29800 (N_29800,N_27883,N_28125);
or U29801 (N_29801,N_27855,N_27748);
or U29802 (N_29802,N_27639,N_28644);
nor U29803 (N_29803,N_28695,N_28299);
nand U29804 (N_29804,N_28223,N_27999);
nand U29805 (N_29805,N_27841,N_28519);
xor U29806 (N_29806,N_28221,N_28702);
nor U29807 (N_29807,N_27628,N_27686);
nand U29808 (N_29808,N_27658,N_27755);
nor U29809 (N_29809,N_28153,N_27861);
nand U29810 (N_29810,N_28726,N_28619);
xor U29811 (N_29811,N_28766,N_27864);
and U29812 (N_29812,N_28107,N_28266);
and U29813 (N_29813,N_28346,N_27668);
xor U29814 (N_29814,N_28550,N_28399);
xor U29815 (N_29815,N_27914,N_28752);
and U29816 (N_29816,N_27729,N_27640);
nand U29817 (N_29817,N_28609,N_28238);
nor U29818 (N_29818,N_27638,N_27945);
or U29819 (N_29819,N_27802,N_27719);
and U29820 (N_29820,N_27859,N_28486);
xor U29821 (N_29821,N_28564,N_27856);
and U29822 (N_29822,N_28760,N_27748);
xnor U29823 (N_29823,N_28769,N_28716);
xor U29824 (N_29824,N_28525,N_27991);
xnor U29825 (N_29825,N_28234,N_27786);
xnor U29826 (N_29826,N_28366,N_27804);
nor U29827 (N_29827,N_28637,N_28656);
xor U29828 (N_29828,N_28019,N_28287);
nor U29829 (N_29829,N_28403,N_28687);
nor U29830 (N_29830,N_28697,N_28405);
nand U29831 (N_29831,N_28625,N_28740);
xor U29832 (N_29832,N_28700,N_28105);
xor U29833 (N_29833,N_28314,N_27968);
and U29834 (N_29834,N_28169,N_28519);
nand U29835 (N_29835,N_28354,N_27846);
nor U29836 (N_29836,N_27985,N_28284);
xor U29837 (N_29837,N_28140,N_28636);
nand U29838 (N_29838,N_28394,N_27962);
or U29839 (N_29839,N_27812,N_28783);
nand U29840 (N_29840,N_27864,N_27809);
xor U29841 (N_29841,N_28191,N_28166);
nand U29842 (N_29842,N_28455,N_28641);
xnor U29843 (N_29843,N_28253,N_27754);
nor U29844 (N_29844,N_28264,N_27886);
nand U29845 (N_29845,N_28753,N_27720);
xnor U29846 (N_29846,N_27990,N_28359);
nor U29847 (N_29847,N_28570,N_28632);
xor U29848 (N_29848,N_27721,N_27955);
or U29849 (N_29849,N_27800,N_27658);
nand U29850 (N_29850,N_28227,N_28160);
nor U29851 (N_29851,N_28569,N_27661);
xnor U29852 (N_29852,N_28126,N_27673);
xor U29853 (N_29853,N_28424,N_28225);
nor U29854 (N_29854,N_28487,N_28226);
nor U29855 (N_29855,N_28152,N_28419);
nand U29856 (N_29856,N_28693,N_28146);
nand U29857 (N_29857,N_27983,N_28161);
or U29858 (N_29858,N_28693,N_27799);
nand U29859 (N_29859,N_28410,N_27982);
nor U29860 (N_29860,N_28549,N_27734);
nand U29861 (N_29861,N_27806,N_28617);
nor U29862 (N_29862,N_28705,N_28715);
xor U29863 (N_29863,N_28417,N_28193);
nor U29864 (N_29864,N_28303,N_28371);
and U29865 (N_29865,N_28580,N_27880);
or U29866 (N_29866,N_28096,N_28226);
or U29867 (N_29867,N_28758,N_27822);
nor U29868 (N_29868,N_27909,N_28380);
xnor U29869 (N_29869,N_28219,N_28443);
nor U29870 (N_29870,N_28140,N_28791);
nor U29871 (N_29871,N_28553,N_27654);
and U29872 (N_29872,N_28636,N_28730);
or U29873 (N_29873,N_27707,N_28570);
nand U29874 (N_29874,N_28567,N_27825);
and U29875 (N_29875,N_28483,N_28592);
or U29876 (N_29876,N_27860,N_28653);
nand U29877 (N_29877,N_27665,N_28266);
nand U29878 (N_29878,N_28339,N_27947);
xor U29879 (N_29879,N_27770,N_27971);
xnor U29880 (N_29880,N_28490,N_28518);
nor U29881 (N_29881,N_28710,N_28724);
and U29882 (N_29882,N_27699,N_28309);
nor U29883 (N_29883,N_27872,N_28047);
and U29884 (N_29884,N_28508,N_27628);
xor U29885 (N_29885,N_28104,N_27607);
nor U29886 (N_29886,N_28275,N_27818);
and U29887 (N_29887,N_28005,N_28218);
nand U29888 (N_29888,N_28084,N_28027);
nor U29889 (N_29889,N_28527,N_28014);
xnor U29890 (N_29890,N_28788,N_28240);
and U29891 (N_29891,N_28033,N_28456);
and U29892 (N_29892,N_27895,N_27827);
xor U29893 (N_29893,N_28071,N_28394);
or U29894 (N_29894,N_28048,N_28045);
nand U29895 (N_29895,N_27831,N_27626);
nand U29896 (N_29896,N_28327,N_28140);
or U29897 (N_29897,N_27747,N_28243);
nor U29898 (N_29898,N_28485,N_27785);
nor U29899 (N_29899,N_28615,N_28224);
or U29900 (N_29900,N_27971,N_28792);
nor U29901 (N_29901,N_27847,N_27859);
nand U29902 (N_29902,N_28637,N_27819);
nor U29903 (N_29903,N_28633,N_27635);
and U29904 (N_29904,N_28443,N_28785);
or U29905 (N_29905,N_28728,N_27605);
and U29906 (N_29906,N_27699,N_28183);
nand U29907 (N_29907,N_27954,N_27912);
or U29908 (N_29908,N_28587,N_27907);
nor U29909 (N_29909,N_28221,N_27793);
nor U29910 (N_29910,N_28230,N_27796);
and U29911 (N_29911,N_28005,N_28647);
nor U29912 (N_29912,N_28019,N_28096);
xor U29913 (N_29913,N_28166,N_28102);
nor U29914 (N_29914,N_27659,N_27800);
nor U29915 (N_29915,N_27780,N_28424);
or U29916 (N_29916,N_28033,N_27736);
xor U29917 (N_29917,N_28698,N_28231);
and U29918 (N_29918,N_28385,N_28026);
and U29919 (N_29919,N_28384,N_27841);
xnor U29920 (N_29920,N_27636,N_28265);
xor U29921 (N_29921,N_27996,N_28554);
xnor U29922 (N_29922,N_28037,N_28307);
nand U29923 (N_29923,N_27832,N_28620);
and U29924 (N_29924,N_28133,N_28614);
or U29925 (N_29925,N_27783,N_27666);
and U29926 (N_29926,N_28156,N_28545);
xnor U29927 (N_29927,N_28290,N_28266);
or U29928 (N_29928,N_27966,N_28536);
nand U29929 (N_29929,N_27898,N_27982);
or U29930 (N_29930,N_28601,N_27647);
nor U29931 (N_29931,N_28254,N_28700);
or U29932 (N_29932,N_28195,N_28717);
or U29933 (N_29933,N_28420,N_27759);
nor U29934 (N_29934,N_27656,N_27960);
or U29935 (N_29935,N_28352,N_28054);
nand U29936 (N_29936,N_28162,N_28603);
nor U29937 (N_29937,N_28450,N_28524);
nor U29938 (N_29938,N_28257,N_28625);
xnor U29939 (N_29939,N_28642,N_28208);
nor U29940 (N_29940,N_28567,N_27796);
xor U29941 (N_29941,N_28087,N_28486);
xor U29942 (N_29942,N_28247,N_28251);
or U29943 (N_29943,N_28017,N_28677);
xor U29944 (N_29944,N_27644,N_28601);
and U29945 (N_29945,N_28432,N_28386);
nor U29946 (N_29946,N_28458,N_27974);
or U29947 (N_29947,N_27605,N_28189);
or U29948 (N_29948,N_28686,N_27655);
or U29949 (N_29949,N_28147,N_28121);
and U29950 (N_29950,N_28663,N_27638);
and U29951 (N_29951,N_28592,N_28513);
or U29952 (N_29952,N_28658,N_28583);
or U29953 (N_29953,N_28576,N_28322);
nor U29954 (N_29954,N_27690,N_27757);
nand U29955 (N_29955,N_28470,N_27798);
nand U29956 (N_29956,N_27800,N_28207);
nor U29957 (N_29957,N_27634,N_28154);
or U29958 (N_29958,N_28466,N_27917);
or U29959 (N_29959,N_28419,N_28122);
and U29960 (N_29960,N_27612,N_28501);
nand U29961 (N_29961,N_27946,N_27781);
or U29962 (N_29962,N_28247,N_28607);
nand U29963 (N_29963,N_27709,N_28783);
nor U29964 (N_29964,N_27823,N_28386);
xnor U29965 (N_29965,N_27648,N_28364);
xor U29966 (N_29966,N_28680,N_27824);
nor U29967 (N_29967,N_27986,N_28470);
nand U29968 (N_29968,N_28777,N_27695);
or U29969 (N_29969,N_28134,N_28643);
and U29970 (N_29970,N_28023,N_27642);
nand U29971 (N_29971,N_28736,N_28141);
or U29972 (N_29972,N_28380,N_28559);
nand U29973 (N_29973,N_27919,N_27939);
and U29974 (N_29974,N_27819,N_28037);
nor U29975 (N_29975,N_28212,N_27663);
nor U29976 (N_29976,N_28787,N_28219);
and U29977 (N_29977,N_28162,N_27613);
and U29978 (N_29978,N_28610,N_28615);
nor U29979 (N_29979,N_28257,N_28694);
and U29980 (N_29980,N_27683,N_27653);
and U29981 (N_29981,N_27959,N_27716);
nand U29982 (N_29982,N_28589,N_27693);
or U29983 (N_29983,N_27831,N_28319);
nand U29984 (N_29984,N_28376,N_27968);
and U29985 (N_29985,N_28320,N_27996);
and U29986 (N_29986,N_28545,N_28497);
xor U29987 (N_29987,N_27826,N_28401);
or U29988 (N_29988,N_28695,N_28437);
xnor U29989 (N_29989,N_28561,N_28650);
xnor U29990 (N_29990,N_27721,N_28422);
xnor U29991 (N_29991,N_28288,N_28474);
and U29992 (N_29992,N_28585,N_28128);
or U29993 (N_29993,N_27737,N_28755);
nand U29994 (N_29994,N_27710,N_28385);
nor U29995 (N_29995,N_28088,N_28562);
nor U29996 (N_29996,N_28246,N_27922);
or U29997 (N_29997,N_28096,N_28693);
xnor U29998 (N_29998,N_28573,N_28444);
xnor U29999 (N_29999,N_28177,N_27910);
nor UO_0 (O_0,N_29879,N_29571);
nand UO_1 (O_1,N_29679,N_29485);
xnor UO_2 (O_2,N_28814,N_29740);
and UO_3 (O_3,N_29769,N_29018);
xor UO_4 (O_4,N_28866,N_29764);
or UO_5 (O_5,N_29731,N_29326);
and UO_6 (O_6,N_29661,N_28869);
nand UO_7 (O_7,N_29974,N_29623);
xnor UO_8 (O_8,N_29413,N_29736);
nand UO_9 (O_9,N_29927,N_29705);
and UO_10 (O_10,N_29333,N_29167);
nor UO_11 (O_11,N_29634,N_29351);
nand UO_12 (O_12,N_29364,N_28872);
nor UO_13 (O_13,N_29394,N_29063);
xnor UO_14 (O_14,N_29117,N_29432);
and UO_15 (O_15,N_29531,N_29497);
or UO_16 (O_16,N_29620,N_29763);
and UO_17 (O_17,N_29194,N_29986);
nand UO_18 (O_18,N_29648,N_29630);
and UO_19 (O_19,N_29170,N_29469);
nor UO_20 (O_20,N_29988,N_29857);
nor UO_21 (O_21,N_29292,N_29866);
nand UO_22 (O_22,N_29185,N_29157);
and UO_23 (O_23,N_28870,N_29835);
nor UO_24 (O_24,N_29340,N_28988);
xnor UO_25 (O_25,N_29047,N_29955);
and UO_26 (O_26,N_29462,N_29999);
xnor UO_27 (O_27,N_29206,N_29884);
nand UO_28 (O_28,N_29732,N_29041);
nor UO_29 (O_29,N_28820,N_29408);
nor UO_30 (O_30,N_29628,N_29823);
nor UO_31 (O_31,N_29320,N_29304);
and UO_32 (O_32,N_29098,N_29481);
nor UO_33 (O_33,N_29779,N_29298);
nor UO_34 (O_34,N_29305,N_29338);
xor UO_35 (O_35,N_29443,N_29285);
or UO_36 (O_36,N_29989,N_29971);
and UO_37 (O_37,N_29112,N_29796);
nand UO_38 (O_38,N_29187,N_29471);
and UO_39 (O_39,N_28995,N_28977);
or UO_40 (O_40,N_29213,N_28975);
xnor UO_41 (O_41,N_28837,N_29398);
nand UO_42 (O_42,N_29843,N_29150);
and UO_43 (O_43,N_29091,N_29093);
xor UO_44 (O_44,N_29082,N_29390);
nor UO_45 (O_45,N_29864,N_29061);
nand UO_46 (O_46,N_29528,N_29113);
and UO_47 (O_47,N_28928,N_29703);
and UO_48 (O_48,N_29611,N_28822);
and UO_49 (O_49,N_29165,N_29572);
or UO_50 (O_50,N_29179,N_29361);
or UO_51 (O_51,N_29455,N_29071);
and UO_52 (O_52,N_29598,N_28941);
xor UO_53 (O_53,N_29174,N_29141);
xnor UO_54 (O_54,N_29938,N_29537);
and UO_55 (O_55,N_29555,N_29618);
xnor UO_56 (O_56,N_29677,N_29559);
nor UO_57 (O_57,N_29714,N_29895);
nor UO_58 (O_58,N_29011,N_28816);
xnor UO_59 (O_59,N_29553,N_29060);
xor UO_60 (O_60,N_29662,N_29614);
and UO_61 (O_61,N_29266,N_29586);
xor UO_62 (O_62,N_29981,N_29059);
or UO_63 (O_63,N_28905,N_29655);
xnor UO_64 (O_64,N_29871,N_28852);
nor UO_65 (O_65,N_29388,N_28960);
or UO_66 (O_66,N_29079,N_29022);
nor UO_67 (O_67,N_29268,N_28901);
xnor UO_68 (O_68,N_29429,N_28921);
nor UO_69 (O_69,N_29793,N_29335);
nor UO_70 (O_70,N_29270,N_28855);
nand UO_71 (O_71,N_29133,N_29104);
nand UO_72 (O_72,N_29277,N_29842);
or UO_73 (O_73,N_29501,N_29651);
nand UO_74 (O_74,N_29342,N_29504);
xor UO_75 (O_75,N_29735,N_29996);
xor UO_76 (O_76,N_29128,N_29175);
or UO_77 (O_77,N_28970,N_28850);
and UO_78 (O_78,N_29404,N_29665);
xnor UO_79 (O_79,N_29992,N_29296);
and UO_80 (O_80,N_29554,N_29575);
and UO_81 (O_81,N_29035,N_29543);
or UO_82 (O_82,N_29858,N_29368);
or UO_83 (O_83,N_29287,N_28823);
and UO_84 (O_84,N_29813,N_29393);
nand UO_85 (O_85,N_29660,N_29513);
nor UO_86 (O_86,N_28839,N_29419);
or UO_87 (O_87,N_28965,N_28818);
or UO_88 (O_88,N_29007,N_29932);
and UO_89 (O_89,N_29182,N_29682);
or UO_90 (O_90,N_29297,N_28896);
xor UO_91 (O_91,N_29158,N_29922);
or UO_92 (O_92,N_29567,N_29028);
xor UO_93 (O_93,N_28914,N_29283);
xnor UO_94 (O_94,N_29905,N_29057);
nor UO_95 (O_95,N_29363,N_29610);
xnor UO_96 (O_96,N_29307,N_29316);
or UO_97 (O_97,N_29897,N_29839);
and UO_98 (O_98,N_29903,N_28813);
nor UO_99 (O_99,N_29696,N_28880);
or UO_100 (O_100,N_29697,N_28978);
xor UO_101 (O_101,N_29138,N_29994);
and UO_102 (O_102,N_29916,N_29299);
or UO_103 (O_103,N_28930,N_29937);
xnor UO_104 (O_104,N_29445,N_28885);
or UO_105 (O_105,N_28824,N_29780);
nand UO_106 (O_106,N_29952,N_29750);
nor UO_107 (O_107,N_29433,N_29540);
or UO_108 (O_108,N_29005,N_29849);
xor UO_109 (O_109,N_28926,N_28927);
nand UO_110 (O_110,N_29476,N_29101);
nor UO_111 (O_111,N_29600,N_29426);
nor UO_112 (O_112,N_29192,N_28856);
nand UO_113 (O_113,N_29350,N_29810);
or UO_114 (O_114,N_29089,N_28805);
and UO_115 (O_115,N_29243,N_29886);
xnor UO_116 (O_116,N_29414,N_29558);
and UO_117 (O_117,N_29752,N_28831);
or UO_118 (O_118,N_29303,N_29578);
and UO_119 (O_119,N_29218,N_29377);
nand UO_120 (O_120,N_29759,N_29959);
and UO_121 (O_121,N_29009,N_29654);
xnor UO_122 (O_122,N_29819,N_28952);
nand UO_123 (O_123,N_28834,N_29765);
and UO_124 (O_124,N_29706,N_29470);
nor UO_125 (O_125,N_29692,N_28929);
nand UO_126 (O_126,N_28990,N_29379);
and UO_127 (O_127,N_29427,N_29638);
nor UO_128 (O_128,N_28807,N_29902);
xnor UO_129 (O_129,N_28985,N_28851);
and UO_130 (O_130,N_28806,N_28833);
xnor UO_131 (O_131,N_29392,N_29383);
or UO_132 (O_132,N_29925,N_29210);
xnor UO_133 (O_133,N_29695,N_29286);
nand UO_134 (O_134,N_28871,N_28948);
nand UO_135 (O_135,N_29171,N_28974);
nand UO_136 (O_136,N_29755,N_29500);
nand UO_137 (O_137,N_29778,N_29967);
nor UO_138 (O_138,N_29139,N_29593);
nor UO_139 (O_139,N_29930,N_28966);
xor UO_140 (O_140,N_29597,N_29710);
or UO_141 (O_141,N_29026,N_29920);
and UO_142 (O_142,N_28991,N_28810);
xor UO_143 (O_143,N_29107,N_29966);
nand UO_144 (O_144,N_28876,N_29233);
xor UO_145 (O_145,N_29362,N_29459);
xor UO_146 (O_146,N_28875,N_29596);
xnor UO_147 (O_147,N_28981,N_28846);
xor UO_148 (O_148,N_29817,N_29032);
nand UO_149 (O_149,N_29818,N_29207);
or UO_150 (O_150,N_29657,N_29936);
nor UO_151 (O_151,N_29948,N_28865);
nor UO_152 (O_152,N_29223,N_29904);
and UO_153 (O_153,N_29401,N_28946);
or UO_154 (O_154,N_29950,N_29105);
nor UO_155 (O_155,N_29330,N_29797);
nand UO_156 (O_156,N_29530,N_29457);
nand UO_157 (O_157,N_29081,N_29766);
xor UO_158 (O_158,N_29040,N_29183);
or UO_159 (O_159,N_29100,N_29672);
xor UO_160 (O_160,N_29295,N_29613);
nand UO_161 (O_161,N_29365,N_29702);
and UO_162 (O_162,N_29760,N_29532);
and UO_163 (O_163,N_29560,N_29716);
xnor UO_164 (O_164,N_29012,N_29514);
nor UO_165 (O_165,N_29585,N_28924);
or UO_166 (O_166,N_29900,N_29131);
and UO_167 (O_167,N_29804,N_29375);
and UO_168 (O_168,N_29162,N_29521);
nand UO_169 (O_169,N_29889,N_29870);
nand UO_170 (O_170,N_29946,N_29331);
and UO_171 (O_171,N_28940,N_29641);
nand UO_172 (O_172,N_29496,N_29355);
xor UO_173 (O_173,N_29491,N_29958);
nand UO_174 (O_174,N_29747,N_29727);
nor UO_175 (O_175,N_29255,N_29836);
nor UO_176 (O_176,N_29119,N_29888);
nor UO_177 (O_177,N_29229,N_29873);
nand UO_178 (O_178,N_28878,N_29973);
nand UO_179 (O_179,N_29405,N_29947);
nand UO_180 (O_180,N_29103,N_29826);
nand UO_181 (O_181,N_29647,N_28910);
or UO_182 (O_182,N_28933,N_29738);
xor UO_183 (O_183,N_29939,N_29056);
nand UO_184 (O_184,N_28853,N_29008);
and UO_185 (O_185,N_29809,N_29454);
xnor UO_186 (O_186,N_29734,N_29058);
nand UO_187 (O_187,N_29371,N_29686);
nor UO_188 (O_188,N_29325,N_29701);
or UO_189 (O_189,N_29482,N_29953);
and UO_190 (O_190,N_29196,N_29694);
or UO_191 (O_191,N_29359,N_29965);
xnor UO_192 (O_192,N_29717,N_29786);
xnor UO_193 (O_193,N_29762,N_29632);
nand UO_194 (O_194,N_29653,N_29267);
nand UO_195 (O_195,N_28889,N_29945);
nor UO_196 (O_196,N_29507,N_29699);
xnor UO_197 (O_197,N_29017,N_29667);
nor UO_198 (O_198,N_29991,N_29739);
nor UO_199 (O_199,N_28947,N_29577);
nor UO_200 (O_200,N_29110,N_29216);
nand UO_201 (O_201,N_29396,N_29792);
nor UO_202 (O_202,N_28968,N_28882);
xor UO_203 (O_203,N_28913,N_29681);
nand UO_204 (O_204,N_28916,N_29534);
and UO_205 (O_205,N_29372,N_29837);
nor UO_206 (O_206,N_29652,N_29424);
nand UO_207 (O_207,N_29391,N_29376);
xor UO_208 (O_208,N_28979,N_29006);
nor UO_209 (O_209,N_29848,N_29129);
nor UO_210 (O_210,N_29893,N_29834);
xnor UO_211 (O_211,N_28939,N_29417);
nor UO_212 (O_212,N_29146,N_29689);
or UO_213 (O_213,N_29294,N_29815);
xor UO_214 (O_214,N_29195,N_29415);
nand UO_215 (O_215,N_29197,N_29982);
nand UO_216 (O_216,N_29944,N_29990);
or UO_217 (O_217,N_29328,N_29399);
nor UO_218 (O_218,N_28893,N_28817);
or UO_219 (O_219,N_29010,N_29998);
nor UO_220 (O_220,N_29219,N_28992);
or UO_221 (O_221,N_29776,N_29193);
nand UO_222 (O_222,N_29224,N_29409);
nor UO_223 (O_223,N_29386,N_28879);
and UO_224 (O_224,N_29172,N_29087);
or UO_225 (O_225,N_29931,N_29186);
nand UO_226 (O_226,N_28842,N_29924);
nor UO_227 (O_227,N_29599,N_29088);
nor UO_228 (O_228,N_29257,N_29321);
nor UO_229 (O_229,N_29512,N_29220);
and UO_230 (O_230,N_28890,N_29544);
and UO_231 (O_231,N_29824,N_29538);
nand UO_232 (O_232,N_29024,N_29607);
nor UO_233 (O_233,N_28958,N_29700);
or UO_234 (O_234,N_28997,N_28804);
nand UO_235 (O_235,N_29083,N_29830);
nand UO_236 (O_236,N_28937,N_29214);
and UO_237 (O_237,N_29642,N_29301);
nand UO_238 (O_238,N_29909,N_28987);
nor UO_239 (O_239,N_29217,N_29878);
xor UO_240 (O_240,N_29027,N_29136);
nand UO_241 (O_241,N_29524,N_29366);
nor UO_242 (O_242,N_29844,N_29256);
xnor UO_243 (O_243,N_29676,N_29042);
nand UO_244 (O_244,N_29502,N_29520);
nand UO_245 (O_245,N_29908,N_29322);
nand UO_246 (O_246,N_29664,N_29108);
nor UO_247 (O_247,N_29438,N_28830);
nand UO_248 (O_248,N_29671,N_29777);
nand UO_249 (O_249,N_29451,N_29806);
and UO_250 (O_250,N_28858,N_29095);
or UO_251 (O_251,N_29789,N_29508);
nor UO_252 (O_252,N_29487,N_29984);
xor UO_253 (O_253,N_29016,N_29280);
and UO_254 (O_254,N_29788,N_29822);
or UO_255 (O_255,N_29977,N_29282);
nand UO_256 (O_256,N_29166,N_29891);
and UO_257 (O_257,N_29724,N_29592);
xnor UO_258 (O_258,N_29475,N_28920);
xor UO_259 (O_259,N_29120,N_28838);
and UO_260 (O_260,N_29983,N_28993);
nor UO_261 (O_261,N_28969,N_29687);
and UO_262 (O_262,N_29072,N_29646);
nor UO_263 (O_263,N_29494,N_29854);
or UO_264 (O_264,N_29400,N_29782);
nand UO_265 (O_265,N_28801,N_29872);
nand UO_266 (O_266,N_28938,N_28959);
nor UO_267 (O_267,N_29463,N_29021);
xnor UO_268 (O_268,N_29637,N_29617);
nor UO_269 (O_269,N_28945,N_29013);
nand UO_270 (O_270,N_29441,N_29847);
nor UO_271 (O_271,N_29595,N_29626);
xor UO_272 (O_272,N_29343,N_29771);
nand UO_273 (O_273,N_29728,N_29160);
nor UO_274 (O_274,N_29410,N_29352);
xnor UO_275 (O_275,N_29756,N_28955);
nor UO_276 (O_276,N_28912,N_29180);
nand UO_277 (O_277,N_29754,N_29411);
xor UO_278 (O_278,N_29923,N_29204);
or UO_279 (O_279,N_29465,N_29020);
xnor UO_280 (O_280,N_29985,N_28891);
nor UO_281 (O_281,N_29801,N_29142);
xor UO_282 (O_282,N_29940,N_29550);
and UO_283 (O_283,N_29275,N_29498);
and UO_284 (O_284,N_29918,N_29484);
nor UO_285 (O_285,N_29054,N_29300);
nor UO_286 (O_286,N_29407,N_29045);
nand UO_287 (O_287,N_28903,N_29643);
xor UO_288 (O_288,N_29838,N_29161);
nand UO_289 (O_289,N_29862,N_29566);
and UO_290 (O_290,N_28815,N_29656);
and UO_291 (O_291,N_29264,N_29529);
and UO_292 (O_292,N_29506,N_29458);
xor UO_293 (O_293,N_29489,N_29143);
nor UO_294 (O_294,N_29680,N_29068);
or UO_295 (O_295,N_29044,N_29808);
nor UO_296 (O_296,N_29278,N_29499);
or UO_297 (O_297,N_29076,N_29025);
or UO_298 (O_298,N_29684,N_29370);
nor UO_299 (O_299,N_29608,N_29406);
nand UO_300 (O_300,N_29894,N_29997);
xor UO_301 (O_301,N_29743,N_28971);
and UO_302 (O_302,N_29188,N_29437);
xor UO_303 (O_303,N_28906,N_29271);
or UO_304 (O_304,N_29159,N_29052);
xor UO_305 (O_305,N_29466,N_28847);
and UO_306 (O_306,N_29825,N_29601);
nor UO_307 (O_307,N_28973,N_29516);
nor UO_308 (O_308,N_29725,N_29645);
xnor UO_309 (O_309,N_29688,N_28923);
or UO_310 (O_310,N_29704,N_29230);
nand UO_311 (O_311,N_29957,N_29348);
nor UO_312 (O_312,N_28976,N_29757);
nor UO_313 (O_313,N_28898,N_28907);
nand UO_314 (O_314,N_29783,N_29452);
nor UO_315 (O_315,N_28809,N_29073);
xnor UO_316 (O_316,N_29718,N_29004);
nor UO_317 (O_317,N_29561,N_29075);
nand UO_318 (O_318,N_29053,N_29852);
or UO_319 (O_319,N_29951,N_29883);
nor UO_320 (O_320,N_29263,N_29448);
or UO_321 (O_321,N_29774,N_29163);
or UO_322 (O_322,N_29876,N_29055);
nand UO_323 (O_323,N_29323,N_29354);
nor UO_324 (O_324,N_29851,N_28884);
nand UO_325 (O_325,N_28825,N_29861);
nor UO_326 (O_326,N_28840,N_29031);
or UO_327 (O_327,N_29910,N_28962);
nand UO_328 (O_328,N_28835,N_29802);
or UO_329 (O_329,N_28881,N_29557);
nor UO_330 (O_330,N_29935,N_28859);
or UO_331 (O_331,N_29753,N_29449);
and UO_332 (O_332,N_29892,N_29033);
nor UO_333 (O_333,N_29358,N_29503);
nand UO_334 (O_334,N_29832,N_29023);
nand UO_335 (O_335,N_29134,N_29302);
xnor UO_336 (O_336,N_29001,N_28808);
nand UO_337 (O_337,N_28849,N_29890);
nand UO_338 (O_338,N_29336,N_29418);
xor UO_339 (O_339,N_29464,N_28802);
nor UO_340 (O_340,N_29546,N_29240);
nor UO_341 (O_341,N_29238,N_28800);
or UO_342 (O_342,N_29430,N_29209);
or UO_343 (O_343,N_28867,N_29145);
nand UO_344 (O_344,N_29781,N_29722);
and UO_345 (O_345,N_29833,N_29914);
or UO_346 (O_346,N_28980,N_29106);
or UO_347 (O_347,N_29666,N_29226);
or UO_348 (O_348,N_29311,N_28989);
nand UO_349 (O_349,N_29199,N_29976);
nand UO_350 (O_350,N_29200,N_29373);
and UO_351 (O_351,N_29744,N_29719);
and UO_352 (O_352,N_29591,N_29190);
nor UO_353 (O_353,N_29840,N_29477);
xor UO_354 (O_354,N_29074,N_29709);
or UO_355 (O_355,N_29215,N_29245);
and UO_356 (O_356,N_28843,N_29621);
xor UO_357 (O_357,N_29259,N_29422);
or UO_358 (O_358,N_28899,N_29556);
xnor UO_359 (O_359,N_29313,N_29616);
nand UO_360 (O_360,N_29602,N_29212);
nand UO_361 (O_361,N_28922,N_29960);
nand UO_362 (O_362,N_29549,N_29085);
nor UO_363 (O_363,N_29000,N_28996);
nand UO_364 (O_364,N_29490,N_29587);
nor UO_365 (O_365,N_29551,N_29683);
xnor UO_366 (O_366,N_29019,N_29887);
and UO_367 (O_367,N_29912,N_29594);
nor UO_368 (O_368,N_29547,N_29720);
or UO_369 (O_369,N_29048,N_29880);
nand UO_370 (O_370,N_29674,N_29254);
nor UO_371 (O_371,N_29062,N_29712);
xnor UO_372 (O_372,N_29367,N_29673);
xnor UO_373 (O_373,N_29246,N_28982);
nor UO_374 (O_374,N_29345,N_29533);
nor UO_375 (O_375,N_28999,N_28918);
and UO_376 (O_376,N_29580,N_29576);
nand UO_377 (O_377,N_28964,N_29369);
and UO_378 (O_378,N_29114,N_29177);
xnor UO_379 (O_379,N_29541,N_29269);
nand UO_380 (O_380,N_29065,N_29588);
and UO_381 (O_381,N_29517,N_29154);
xor UO_382 (O_382,N_29926,N_29315);
nand UO_383 (O_383,N_29942,N_29856);
or UO_384 (O_384,N_29590,N_28886);
and UO_385 (O_385,N_28949,N_29241);
or UO_386 (O_386,N_29751,N_29868);
and UO_387 (O_387,N_29488,N_29374);
nand UO_388 (O_388,N_29511,N_28909);
or UO_389 (O_389,N_29510,N_29746);
and UO_390 (O_390,N_28915,N_29066);
and UO_391 (O_391,N_29569,N_28956);
or UO_392 (O_392,N_29135,N_29542);
and UO_393 (O_393,N_28863,N_29144);
and UO_394 (O_394,N_29795,N_29583);
or UO_395 (O_395,N_28892,N_29030);
or UO_396 (O_396,N_29568,N_29231);
nor UO_397 (O_397,N_29874,N_28986);
nor UO_398 (O_398,N_29347,N_29669);
nor UO_399 (O_399,N_29262,N_28967);
nor UO_400 (O_400,N_29225,N_29049);
or UO_401 (O_401,N_29385,N_29650);
and UO_402 (O_402,N_29064,N_29198);
and UO_403 (O_403,N_28994,N_29726);
nor UO_404 (O_404,N_28895,N_29798);
and UO_405 (O_405,N_29395,N_29312);
xor UO_406 (O_406,N_29324,N_28911);
and UO_407 (O_407,N_29954,N_29658);
or UO_408 (O_408,N_28868,N_29865);
nand UO_409 (O_409,N_29084,N_29222);
xnor UO_410 (O_410,N_29799,N_29609);
and UO_411 (O_411,N_29360,N_29397);
nor UO_412 (O_412,N_29439,N_29527);
nand UO_413 (O_413,N_29811,N_29251);
or UO_414 (O_414,N_29132,N_29639);
xor UO_415 (O_415,N_29289,N_29729);
and UO_416 (O_416,N_29234,N_29619);
nor UO_417 (O_417,N_29612,N_29434);
nor UO_418 (O_418,N_29941,N_29147);
nor UO_419 (O_419,N_29067,N_28844);
or UO_420 (O_420,N_29094,N_29814);
or UO_421 (O_421,N_29221,N_29339);
nor UO_422 (O_422,N_29090,N_29123);
nand UO_423 (O_423,N_29308,N_29603);
and UO_424 (O_424,N_29425,N_28861);
or UO_425 (O_425,N_29963,N_29353);
nor UO_426 (O_426,N_29253,N_28932);
and UO_427 (O_427,N_28957,N_29293);
xor UO_428 (O_428,N_29428,N_29495);
nor UO_429 (O_429,N_29440,N_29730);
nand UO_430 (O_430,N_29472,N_29522);
xor UO_431 (O_431,N_29745,N_29127);
nor UO_432 (O_432,N_29970,N_29151);
nor UO_433 (O_433,N_29378,N_29461);
nand UO_434 (O_434,N_29535,N_29911);
or UO_435 (O_435,N_29096,N_29118);
xor UO_436 (O_436,N_29334,N_29260);
or UO_437 (O_437,N_29790,N_29102);
or UO_438 (O_438,N_29480,N_28803);
nand UO_439 (O_439,N_29203,N_29423);
nand UO_440 (O_440,N_29562,N_29281);
nor UO_441 (O_441,N_29121,N_29309);
and UO_442 (O_442,N_29479,N_29919);
xnor UO_443 (O_443,N_28877,N_29152);
or UO_444 (O_444,N_29794,N_29855);
nor UO_445 (O_445,N_29625,N_29721);
or UO_446 (O_446,N_29468,N_29934);
xor UO_447 (O_447,N_28961,N_29034);
xor UO_448 (O_448,N_29306,N_29772);
and UO_449 (O_449,N_29412,N_29173);
xnor UO_450 (O_450,N_29708,N_28984);
and UO_451 (O_451,N_29713,N_29509);
nor UO_452 (O_452,N_29124,N_29467);
xnor UO_453 (O_453,N_29615,N_28897);
nand UO_454 (O_454,N_29381,N_29014);
nor UO_455 (O_455,N_29332,N_29898);
xor UO_456 (O_456,N_29629,N_29928);
and UO_457 (O_457,N_28998,N_29130);
nand UO_458 (O_458,N_28919,N_29933);
nand UO_459 (O_459,N_28972,N_29092);
or UO_460 (O_460,N_29707,N_29015);
and UO_461 (O_461,N_28841,N_29232);
or UO_462 (O_462,N_29962,N_29337);
and UO_463 (O_463,N_28904,N_29149);
xnor UO_464 (O_464,N_29787,N_29274);
xnor UO_465 (O_465,N_29450,N_29693);
nor UO_466 (O_466,N_29137,N_29279);
nand UO_467 (O_467,N_29805,N_29917);
xnor UO_468 (O_468,N_28821,N_29205);
or UO_469 (O_469,N_29273,N_29248);
or UO_470 (O_470,N_28864,N_29344);
nor UO_471 (O_471,N_29447,N_29515);
nand UO_472 (O_472,N_29519,N_28925);
xnor UO_473 (O_473,N_29649,N_29564);
nor UO_474 (O_474,N_29228,N_29478);
nand UO_475 (O_475,N_29431,N_29247);
nor UO_476 (O_476,N_29505,N_29968);
nand UO_477 (O_477,N_29901,N_29288);
nor UO_478 (O_478,N_29906,N_28812);
nor UO_479 (O_479,N_29723,N_29444);
nor UO_480 (O_480,N_29111,N_28954);
nor UO_481 (O_481,N_29659,N_29181);
and UO_482 (O_482,N_29622,N_29156);
xor UO_483 (O_483,N_28900,N_29812);
or UO_484 (O_484,N_29080,N_29474);
nand UO_485 (O_485,N_29964,N_29853);
and UO_486 (O_486,N_29969,N_28832);
or UO_487 (O_487,N_29319,N_29733);
nor UO_488 (O_488,N_29624,N_29863);
or UO_489 (O_489,N_29829,N_29357);
xnor UO_490 (O_490,N_29473,N_28854);
nor UO_491 (O_491,N_29038,N_29627);
nor UO_492 (O_492,N_29276,N_28873);
xnor UO_493 (O_493,N_29109,N_28917);
xnor UO_494 (O_494,N_29800,N_29526);
and UO_495 (O_495,N_29237,N_29046);
and UO_496 (O_496,N_29168,N_29767);
and UO_497 (O_497,N_29148,N_29961);
and UO_498 (O_498,N_29184,N_29972);
or UO_499 (O_499,N_29929,N_28983);
nor UO_500 (O_500,N_29993,N_29387);
nor UO_501 (O_501,N_29606,N_29483);
xnor UO_502 (O_502,N_29860,N_29420);
and UO_503 (O_503,N_29978,N_29690);
nor UO_504 (O_504,N_29202,N_29885);
nand UO_505 (O_505,N_29003,N_29631);
xnor UO_506 (O_506,N_29211,N_29956);
xnor UO_507 (O_507,N_29029,N_29164);
and UO_508 (O_508,N_28894,N_29069);
xor UO_509 (O_509,N_29346,N_29758);
and UO_510 (O_510,N_29741,N_29327);
or UO_511 (O_511,N_28883,N_29349);
and UO_512 (O_512,N_29584,N_29867);
or UO_513 (O_513,N_29460,N_29317);
xor UO_514 (O_514,N_29896,N_29775);
nand UO_515 (O_515,N_29518,N_29841);
and UO_516 (O_516,N_29421,N_29272);
or UO_517 (O_517,N_29265,N_29882);
xnor UO_518 (O_518,N_29122,N_28811);
xor UO_519 (O_519,N_29077,N_29949);
or UO_520 (O_520,N_29770,N_29402);
xnor UO_521 (O_521,N_29821,N_29536);
or UO_522 (O_522,N_29249,N_28951);
nand UO_523 (O_523,N_29899,N_28902);
and UO_524 (O_524,N_29002,N_29605);
or UO_525 (O_525,N_28908,N_29178);
xnor UO_526 (O_526,N_29341,N_29051);
xnor UO_527 (O_527,N_29563,N_28862);
nor UO_528 (O_528,N_29436,N_29176);
and UO_529 (O_529,N_29749,N_29250);
xor UO_530 (O_530,N_29140,N_29493);
nand UO_531 (O_531,N_29525,N_29565);
xnor UO_532 (O_532,N_29227,N_28887);
nand UO_533 (O_533,N_28819,N_29201);
and UO_534 (O_534,N_29456,N_29258);
and UO_535 (O_535,N_29907,N_29845);
and UO_536 (O_536,N_28935,N_29827);
xor UO_537 (O_537,N_29574,N_29711);
or UO_538 (O_538,N_29633,N_29670);
and UO_539 (O_539,N_29453,N_29913);
or UO_540 (O_540,N_29877,N_29078);
nand UO_541 (O_541,N_29492,N_29640);
xor UO_542 (O_542,N_29773,N_29403);
or UO_543 (O_543,N_28953,N_29604);
or UO_544 (O_544,N_29329,N_29486);
xnor UO_545 (O_545,N_28936,N_29115);
nand UO_546 (O_546,N_29442,N_28943);
xnor UO_547 (O_547,N_29668,N_29552);
and UO_548 (O_548,N_28931,N_29291);
or UO_549 (O_549,N_29539,N_29043);
xnor UO_550 (O_550,N_29189,N_28845);
nand UO_551 (O_551,N_28860,N_29678);
or UO_552 (O_552,N_29987,N_29995);
nand UO_553 (O_553,N_29389,N_29037);
and UO_554 (O_554,N_28826,N_29582);
or UO_555 (O_555,N_29242,N_29715);
and UO_556 (O_556,N_29070,N_29831);
and UO_557 (O_557,N_29698,N_29975);
and UO_558 (O_558,N_29675,N_29155);
and UO_559 (O_559,N_29816,N_29039);
and UO_560 (O_560,N_29153,N_29290);
nand UO_561 (O_561,N_29881,N_28888);
nor UO_562 (O_562,N_29523,N_28857);
nor UO_563 (O_563,N_29097,N_29356);
xor UO_564 (O_564,N_29570,N_29036);
xnor UO_565 (O_565,N_29435,N_28829);
or UO_566 (O_566,N_29284,N_29589);
nor UO_567 (O_567,N_29050,N_29244);
nor UO_568 (O_568,N_29875,N_29573);
xor UO_569 (O_569,N_28848,N_29980);
or UO_570 (O_570,N_28828,N_29803);
nand UO_571 (O_571,N_29416,N_29828);
nor UO_572 (O_572,N_29239,N_29807);
or UO_573 (O_573,N_29784,N_28836);
nor UO_574 (O_574,N_29235,N_29915);
nor UO_575 (O_575,N_29791,N_29820);
xnor UO_576 (O_576,N_29380,N_28874);
nand UO_577 (O_577,N_29252,N_29742);
or UO_578 (O_578,N_29636,N_29384);
and UO_579 (O_579,N_29579,N_29099);
xnor UO_580 (O_580,N_29169,N_29310);
or UO_581 (O_581,N_28827,N_29191);
nand UO_582 (O_582,N_29785,N_29644);
nor UO_583 (O_583,N_29116,N_29314);
xor UO_584 (O_584,N_29859,N_28934);
xor UO_585 (O_585,N_29663,N_28950);
nand UO_586 (O_586,N_29979,N_29691);
xnor UO_587 (O_587,N_29737,N_29869);
nand UO_588 (O_588,N_28944,N_29921);
nor UO_589 (O_589,N_29768,N_29545);
or UO_590 (O_590,N_29685,N_29850);
and UO_591 (O_591,N_29446,N_29236);
and UO_592 (O_592,N_29086,N_29548);
xor UO_593 (O_593,N_29846,N_29635);
xnor UO_594 (O_594,N_29581,N_29761);
xnor UO_595 (O_595,N_29261,N_28963);
or UO_596 (O_596,N_29126,N_29208);
nor UO_597 (O_597,N_28942,N_29318);
xor UO_598 (O_598,N_29382,N_29748);
and UO_599 (O_599,N_29125,N_29943);
or UO_600 (O_600,N_29900,N_29175);
xor UO_601 (O_601,N_29862,N_28963);
nand UO_602 (O_602,N_29669,N_29439);
nor UO_603 (O_603,N_28876,N_29275);
and UO_604 (O_604,N_29761,N_28878);
nor UO_605 (O_605,N_28804,N_29894);
or UO_606 (O_606,N_29067,N_29556);
nor UO_607 (O_607,N_29072,N_29304);
and UO_608 (O_608,N_29048,N_28919);
nand UO_609 (O_609,N_29724,N_29938);
or UO_610 (O_610,N_29322,N_28834);
nor UO_611 (O_611,N_29127,N_29638);
and UO_612 (O_612,N_29208,N_29015);
or UO_613 (O_613,N_29010,N_29913);
xor UO_614 (O_614,N_29148,N_29668);
and UO_615 (O_615,N_29158,N_29008);
nand UO_616 (O_616,N_28977,N_29074);
nand UO_617 (O_617,N_28848,N_29605);
nor UO_618 (O_618,N_29520,N_29973);
nor UO_619 (O_619,N_29950,N_29681);
or UO_620 (O_620,N_28928,N_29272);
xnor UO_621 (O_621,N_29957,N_29482);
nor UO_622 (O_622,N_29051,N_28991);
nand UO_623 (O_623,N_28822,N_29617);
and UO_624 (O_624,N_29565,N_29638);
xor UO_625 (O_625,N_28949,N_29623);
or UO_626 (O_626,N_29482,N_28851);
nor UO_627 (O_627,N_28921,N_29477);
and UO_628 (O_628,N_29673,N_28935);
xor UO_629 (O_629,N_29884,N_29689);
xnor UO_630 (O_630,N_28846,N_28808);
nand UO_631 (O_631,N_28938,N_29083);
nor UO_632 (O_632,N_29971,N_28961);
or UO_633 (O_633,N_28848,N_29551);
nor UO_634 (O_634,N_29824,N_29272);
nor UO_635 (O_635,N_29251,N_29632);
or UO_636 (O_636,N_29778,N_29626);
xor UO_637 (O_637,N_29409,N_29516);
nand UO_638 (O_638,N_29341,N_29404);
xor UO_639 (O_639,N_29919,N_29166);
xnor UO_640 (O_640,N_29185,N_29750);
nor UO_641 (O_641,N_29253,N_29861);
xor UO_642 (O_642,N_29824,N_28947);
and UO_643 (O_643,N_29772,N_29916);
or UO_644 (O_644,N_29943,N_29791);
nor UO_645 (O_645,N_29952,N_29529);
nor UO_646 (O_646,N_29163,N_29804);
xnor UO_647 (O_647,N_29475,N_29859);
nand UO_648 (O_648,N_29404,N_29095);
xnor UO_649 (O_649,N_29821,N_29384);
or UO_650 (O_650,N_28928,N_29267);
nor UO_651 (O_651,N_29217,N_28856);
nor UO_652 (O_652,N_29931,N_29523);
or UO_653 (O_653,N_29814,N_29555);
and UO_654 (O_654,N_29252,N_29465);
nor UO_655 (O_655,N_29837,N_29317);
or UO_656 (O_656,N_29768,N_29943);
nor UO_657 (O_657,N_29863,N_29797);
and UO_658 (O_658,N_29171,N_29088);
nor UO_659 (O_659,N_28865,N_29039);
or UO_660 (O_660,N_29661,N_29534);
and UO_661 (O_661,N_29009,N_28842);
nand UO_662 (O_662,N_29187,N_28983);
or UO_663 (O_663,N_29484,N_29199);
nor UO_664 (O_664,N_29876,N_29634);
nand UO_665 (O_665,N_29475,N_29941);
xnor UO_666 (O_666,N_29062,N_29103);
xor UO_667 (O_667,N_29549,N_29268);
nor UO_668 (O_668,N_28812,N_29126);
nor UO_669 (O_669,N_29113,N_29613);
or UO_670 (O_670,N_29546,N_29683);
nor UO_671 (O_671,N_29500,N_29740);
and UO_672 (O_672,N_29076,N_29672);
xnor UO_673 (O_673,N_29019,N_29471);
or UO_674 (O_674,N_29832,N_29553);
nand UO_675 (O_675,N_29597,N_29937);
nor UO_676 (O_676,N_29333,N_29701);
nor UO_677 (O_677,N_29259,N_29915);
xnor UO_678 (O_678,N_29615,N_29657);
and UO_679 (O_679,N_29351,N_29791);
or UO_680 (O_680,N_28837,N_29336);
nor UO_681 (O_681,N_29172,N_29361);
or UO_682 (O_682,N_29056,N_29934);
nor UO_683 (O_683,N_29276,N_29228);
xnor UO_684 (O_684,N_29329,N_29339);
xor UO_685 (O_685,N_29683,N_29565);
nor UO_686 (O_686,N_29103,N_29104);
nand UO_687 (O_687,N_29707,N_28918);
and UO_688 (O_688,N_29446,N_28817);
or UO_689 (O_689,N_29366,N_29912);
nor UO_690 (O_690,N_29536,N_29289);
xor UO_691 (O_691,N_29190,N_29269);
and UO_692 (O_692,N_29612,N_29752);
or UO_693 (O_693,N_29868,N_29340);
or UO_694 (O_694,N_29412,N_28803);
and UO_695 (O_695,N_29485,N_29601);
nand UO_696 (O_696,N_29636,N_29631);
nand UO_697 (O_697,N_29265,N_29419);
and UO_698 (O_698,N_28902,N_29067);
or UO_699 (O_699,N_29665,N_29597);
nand UO_700 (O_700,N_29626,N_29189);
and UO_701 (O_701,N_28862,N_29434);
xnor UO_702 (O_702,N_29752,N_29316);
nand UO_703 (O_703,N_29404,N_28814);
nor UO_704 (O_704,N_29942,N_29044);
xor UO_705 (O_705,N_29305,N_29942);
or UO_706 (O_706,N_29243,N_29460);
nand UO_707 (O_707,N_29450,N_29958);
nor UO_708 (O_708,N_29780,N_29489);
nor UO_709 (O_709,N_29839,N_29777);
nand UO_710 (O_710,N_29275,N_28829);
xor UO_711 (O_711,N_28991,N_29104);
nor UO_712 (O_712,N_29783,N_29921);
xor UO_713 (O_713,N_29827,N_29703);
or UO_714 (O_714,N_29682,N_29642);
and UO_715 (O_715,N_29927,N_29744);
xnor UO_716 (O_716,N_29815,N_29249);
and UO_717 (O_717,N_29899,N_29739);
nor UO_718 (O_718,N_29517,N_29047);
nor UO_719 (O_719,N_29491,N_29180);
xor UO_720 (O_720,N_29569,N_29586);
nand UO_721 (O_721,N_29374,N_29432);
or UO_722 (O_722,N_28865,N_29359);
xnor UO_723 (O_723,N_29542,N_28975);
nor UO_724 (O_724,N_29034,N_29661);
and UO_725 (O_725,N_29999,N_29714);
and UO_726 (O_726,N_28839,N_29812);
xnor UO_727 (O_727,N_29138,N_29635);
nor UO_728 (O_728,N_29380,N_29993);
or UO_729 (O_729,N_29837,N_29514);
xor UO_730 (O_730,N_28804,N_29350);
and UO_731 (O_731,N_29196,N_29551);
and UO_732 (O_732,N_29514,N_29678);
or UO_733 (O_733,N_29002,N_29607);
nor UO_734 (O_734,N_29979,N_29920);
xnor UO_735 (O_735,N_29596,N_29449);
nor UO_736 (O_736,N_28890,N_29267);
and UO_737 (O_737,N_29371,N_29889);
and UO_738 (O_738,N_29152,N_29173);
or UO_739 (O_739,N_29765,N_29202);
xnor UO_740 (O_740,N_29187,N_29585);
nand UO_741 (O_741,N_29527,N_29832);
and UO_742 (O_742,N_29673,N_29275);
or UO_743 (O_743,N_29376,N_29011);
nor UO_744 (O_744,N_29887,N_29076);
and UO_745 (O_745,N_29361,N_29416);
nand UO_746 (O_746,N_29001,N_29984);
nand UO_747 (O_747,N_29822,N_29217);
nor UO_748 (O_748,N_29262,N_29606);
nor UO_749 (O_749,N_29396,N_29373);
nand UO_750 (O_750,N_29048,N_28826);
nor UO_751 (O_751,N_29169,N_29649);
and UO_752 (O_752,N_29656,N_29887);
and UO_753 (O_753,N_29593,N_29972);
or UO_754 (O_754,N_29279,N_29338);
or UO_755 (O_755,N_29193,N_29859);
or UO_756 (O_756,N_28969,N_29190);
xor UO_757 (O_757,N_29583,N_29207);
nand UO_758 (O_758,N_28925,N_28893);
and UO_759 (O_759,N_29294,N_29536);
nand UO_760 (O_760,N_29590,N_29915);
nor UO_761 (O_761,N_29787,N_29564);
or UO_762 (O_762,N_29215,N_29896);
and UO_763 (O_763,N_29946,N_29865);
and UO_764 (O_764,N_29165,N_29901);
and UO_765 (O_765,N_28951,N_28868);
nand UO_766 (O_766,N_29861,N_28877);
nand UO_767 (O_767,N_29663,N_29999);
xnor UO_768 (O_768,N_29266,N_29400);
and UO_769 (O_769,N_29241,N_28807);
or UO_770 (O_770,N_29191,N_28993);
xor UO_771 (O_771,N_28812,N_29797);
nor UO_772 (O_772,N_28903,N_29926);
and UO_773 (O_773,N_29001,N_29967);
and UO_774 (O_774,N_29129,N_29716);
and UO_775 (O_775,N_29756,N_29921);
nor UO_776 (O_776,N_29823,N_29254);
and UO_777 (O_777,N_28818,N_29548);
nor UO_778 (O_778,N_29110,N_29528);
xor UO_779 (O_779,N_29223,N_29423);
xnor UO_780 (O_780,N_29327,N_28846);
and UO_781 (O_781,N_29368,N_29285);
nand UO_782 (O_782,N_29463,N_29708);
xor UO_783 (O_783,N_29628,N_29107);
xor UO_784 (O_784,N_28853,N_29694);
nand UO_785 (O_785,N_29749,N_28939);
or UO_786 (O_786,N_29816,N_29498);
xor UO_787 (O_787,N_29705,N_28847);
nor UO_788 (O_788,N_29637,N_29466);
nand UO_789 (O_789,N_29543,N_29755);
nor UO_790 (O_790,N_29539,N_29429);
or UO_791 (O_791,N_29092,N_29410);
nand UO_792 (O_792,N_29470,N_29038);
nand UO_793 (O_793,N_29197,N_29757);
xnor UO_794 (O_794,N_29682,N_29928);
xnor UO_795 (O_795,N_29484,N_29583);
nand UO_796 (O_796,N_29673,N_29041);
and UO_797 (O_797,N_29810,N_28870);
nand UO_798 (O_798,N_29151,N_29203);
xor UO_799 (O_799,N_29258,N_29289);
nand UO_800 (O_800,N_29601,N_29787);
and UO_801 (O_801,N_29305,N_28939);
or UO_802 (O_802,N_29038,N_28826);
nand UO_803 (O_803,N_29856,N_29071);
xor UO_804 (O_804,N_29024,N_29255);
and UO_805 (O_805,N_29750,N_29799);
xnor UO_806 (O_806,N_29789,N_29329);
and UO_807 (O_807,N_28913,N_29719);
nand UO_808 (O_808,N_29218,N_29454);
nand UO_809 (O_809,N_29961,N_28959);
nand UO_810 (O_810,N_29539,N_28992);
nor UO_811 (O_811,N_29796,N_29905);
or UO_812 (O_812,N_29511,N_29672);
xor UO_813 (O_813,N_29024,N_29659);
nand UO_814 (O_814,N_29190,N_29371);
xnor UO_815 (O_815,N_28807,N_28860);
or UO_816 (O_816,N_29119,N_29331);
nand UO_817 (O_817,N_29741,N_29537);
nand UO_818 (O_818,N_29657,N_29014);
nor UO_819 (O_819,N_29606,N_29301);
xor UO_820 (O_820,N_29370,N_29765);
nand UO_821 (O_821,N_29413,N_29893);
nor UO_822 (O_822,N_29854,N_29852);
or UO_823 (O_823,N_28820,N_29802);
xor UO_824 (O_824,N_29261,N_29440);
and UO_825 (O_825,N_29723,N_29728);
nand UO_826 (O_826,N_29017,N_29140);
nand UO_827 (O_827,N_29386,N_29376);
xor UO_828 (O_828,N_28899,N_29762);
nand UO_829 (O_829,N_29349,N_29227);
xor UO_830 (O_830,N_28814,N_29294);
nor UO_831 (O_831,N_29514,N_29696);
xor UO_832 (O_832,N_29657,N_28847);
or UO_833 (O_833,N_29260,N_28935);
xor UO_834 (O_834,N_29396,N_29241);
xnor UO_835 (O_835,N_29205,N_29541);
nor UO_836 (O_836,N_29351,N_29188);
nand UO_837 (O_837,N_29794,N_28998);
nand UO_838 (O_838,N_28906,N_29925);
xnor UO_839 (O_839,N_29575,N_29817);
and UO_840 (O_840,N_29483,N_29304);
and UO_841 (O_841,N_29935,N_29535);
xnor UO_842 (O_842,N_29156,N_29492);
xor UO_843 (O_843,N_29473,N_29916);
and UO_844 (O_844,N_29985,N_29972);
xnor UO_845 (O_845,N_29027,N_29773);
nand UO_846 (O_846,N_29482,N_29854);
or UO_847 (O_847,N_29337,N_28869);
nor UO_848 (O_848,N_29087,N_29259);
nor UO_849 (O_849,N_29350,N_28864);
or UO_850 (O_850,N_29705,N_29980);
and UO_851 (O_851,N_29428,N_29250);
or UO_852 (O_852,N_29370,N_29336);
and UO_853 (O_853,N_29110,N_29733);
xor UO_854 (O_854,N_28901,N_29830);
nor UO_855 (O_855,N_29123,N_29331);
and UO_856 (O_856,N_29422,N_29749);
nand UO_857 (O_857,N_29470,N_29337);
xor UO_858 (O_858,N_29739,N_29309);
nand UO_859 (O_859,N_29034,N_29041);
nand UO_860 (O_860,N_29944,N_29060);
or UO_861 (O_861,N_29182,N_29977);
nand UO_862 (O_862,N_29406,N_29766);
xor UO_863 (O_863,N_29407,N_29589);
or UO_864 (O_864,N_29333,N_28873);
nand UO_865 (O_865,N_29365,N_29775);
xor UO_866 (O_866,N_29545,N_28846);
or UO_867 (O_867,N_29955,N_29882);
nor UO_868 (O_868,N_29074,N_28844);
nand UO_869 (O_869,N_29036,N_29891);
or UO_870 (O_870,N_28841,N_29550);
nor UO_871 (O_871,N_29828,N_29490);
and UO_872 (O_872,N_29976,N_29395);
nand UO_873 (O_873,N_29315,N_28923);
nand UO_874 (O_874,N_29881,N_29644);
xnor UO_875 (O_875,N_29992,N_29993);
and UO_876 (O_876,N_29391,N_29748);
and UO_877 (O_877,N_29612,N_28942);
or UO_878 (O_878,N_28827,N_29021);
xor UO_879 (O_879,N_29472,N_29726);
xnor UO_880 (O_880,N_29469,N_29679);
xor UO_881 (O_881,N_28931,N_29214);
nand UO_882 (O_882,N_29565,N_29332);
nand UO_883 (O_883,N_29083,N_29723);
and UO_884 (O_884,N_28990,N_29056);
or UO_885 (O_885,N_29782,N_28849);
nand UO_886 (O_886,N_28890,N_29538);
nor UO_887 (O_887,N_29978,N_28823);
nand UO_888 (O_888,N_29021,N_28915);
or UO_889 (O_889,N_29043,N_29831);
nor UO_890 (O_890,N_29708,N_29282);
and UO_891 (O_891,N_28925,N_29604);
or UO_892 (O_892,N_29390,N_28952);
and UO_893 (O_893,N_29960,N_29578);
and UO_894 (O_894,N_29847,N_29442);
xor UO_895 (O_895,N_29101,N_29399);
xnor UO_896 (O_896,N_29087,N_29341);
nor UO_897 (O_897,N_29413,N_29601);
and UO_898 (O_898,N_29394,N_29713);
nor UO_899 (O_899,N_29456,N_29858);
nand UO_900 (O_900,N_29859,N_29452);
and UO_901 (O_901,N_29354,N_29285);
nor UO_902 (O_902,N_29434,N_29350);
nor UO_903 (O_903,N_29981,N_29638);
nor UO_904 (O_904,N_29564,N_29665);
nor UO_905 (O_905,N_29424,N_29140);
or UO_906 (O_906,N_29082,N_29509);
nand UO_907 (O_907,N_29461,N_28928);
xor UO_908 (O_908,N_29014,N_29476);
and UO_909 (O_909,N_28967,N_29350);
nor UO_910 (O_910,N_29053,N_28896);
nor UO_911 (O_911,N_29399,N_29512);
or UO_912 (O_912,N_28991,N_29836);
or UO_913 (O_913,N_29665,N_29979);
xor UO_914 (O_914,N_29029,N_29045);
nand UO_915 (O_915,N_29933,N_28962);
nand UO_916 (O_916,N_29413,N_29762);
xnor UO_917 (O_917,N_29046,N_29345);
nor UO_918 (O_918,N_29013,N_29709);
nand UO_919 (O_919,N_29935,N_29417);
xor UO_920 (O_920,N_29846,N_29565);
or UO_921 (O_921,N_28893,N_29708);
nand UO_922 (O_922,N_29599,N_28887);
xor UO_923 (O_923,N_29005,N_29301);
or UO_924 (O_924,N_28962,N_29724);
nand UO_925 (O_925,N_29780,N_29158);
nand UO_926 (O_926,N_29559,N_29933);
nand UO_927 (O_927,N_29790,N_29161);
nor UO_928 (O_928,N_29541,N_29418);
xnor UO_929 (O_929,N_29907,N_29975);
nor UO_930 (O_930,N_28991,N_29785);
and UO_931 (O_931,N_29509,N_29896);
nand UO_932 (O_932,N_29471,N_28969);
nor UO_933 (O_933,N_29626,N_29510);
nand UO_934 (O_934,N_29481,N_29558);
xnor UO_935 (O_935,N_29074,N_29368);
or UO_936 (O_936,N_29561,N_28833);
nor UO_937 (O_937,N_29136,N_28848);
nor UO_938 (O_938,N_29117,N_29946);
nand UO_939 (O_939,N_29084,N_29383);
nand UO_940 (O_940,N_29943,N_29119);
and UO_941 (O_941,N_29270,N_29233);
nor UO_942 (O_942,N_29935,N_29161);
and UO_943 (O_943,N_29932,N_29058);
nor UO_944 (O_944,N_29816,N_29219);
nand UO_945 (O_945,N_29894,N_29000);
or UO_946 (O_946,N_29780,N_29939);
nand UO_947 (O_947,N_28824,N_29452);
nand UO_948 (O_948,N_29072,N_29891);
nand UO_949 (O_949,N_29154,N_29017);
or UO_950 (O_950,N_29390,N_29426);
xnor UO_951 (O_951,N_29572,N_29845);
nor UO_952 (O_952,N_29941,N_29429);
xor UO_953 (O_953,N_29519,N_29418);
or UO_954 (O_954,N_29124,N_29085);
nand UO_955 (O_955,N_29984,N_29425);
and UO_956 (O_956,N_29096,N_29941);
xor UO_957 (O_957,N_29204,N_29637);
or UO_958 (O_958,N_29895,N_29808);
and UO_959 (O_959,N_29636,N_29640);
xor UO_960 (O_960,N_29992,N_29694);
or UO_961 (O_961,N_29271,N_28884);
nor UO_962 (O_962,N_29417,N_28983);
and UO_963 (O_963,N_29495,N_29963);
and UO_964 (O_964,N_28968,N_29253);
nand UO_965 (O_965,N_28853,N_29067);
nor UO_966 (O_966,N_29213,N_28918);
or UO_967 (O_967,N_29181,N_28934);
and UO_968 (O_968,N_29391,N_29290);
xnor UO_969 (O_969,N_29725,N_28854);
or UO_970 (O_970,N_29120,N_29681);
or UO_971 (O_971,N_29732,N_29413);
xor UO_972 (O_972,N_28903,N_29797);
and UO_973 (O_973,N_29375,N_29627);
or UO_974 (O_974,N_28866,N_28875);
or UO_975 (O_975,N_28942,N_29550);
nand UO_976 (O_976,N_29047,N_29457);
and UO_977 (O_977,N_29862,N_29467);
nand UO_978 (O_978,N_29356,N_29812);
nand UO_979 (O_979,N_29088,N_29395);
and UO_980 (O_980,N_28918,N_29484);
and UO_981 (O_981,N_29503,N_28875);
and UO_982 (O_982,N_29726,N_28979);
or UO_983 (O_983,N_29479,N_29117);
and UO_984 (O_984,N_29798,N_29821);
nor UO_985 (O_985,N_28951,N_29615);
nor UO_986 (O_986,N_29911,N_28984);
or UO_987 (O_987,N_29932,N_28810);
nor UO_988 (O_988,N_29467,N_29755);
xor UO_989 (O_989,N_29995,N_29916);
nand UO_990 (O_990,N_29057,N_29190);
and UO_991 (O_991,N_29646,N_29453);
or UO_992 (O_992,N_29057,N_28883);
or UO_993 (O_993,N_28976,N_29410);
nand UO_994 (O_994,N_29931,N_29481);
and UO_995 (O_995,N_28890,N_29341);
or UO_996 (O_996,N_29869,N_29003);
nand UO_997 (O_997,N_29640,N_28933);
nor UO_998 (O_998,N_28937,N_29791);
xnor UO_999 (O_999,N_29425,N_29752);
or UO_1000 (O_1000,N_29118,N_29967);
and UO_1001 (O_1001,N_29732,N_28937);
xnor UO_1002 (O_1002,N_29497,N_28899);
or UO_1003 (O_1003,N_28850,N_29857);
nor UO_1004 (O_1004,N_28981,N_29627);
or UO_1005 (O_1005,N_29867,N_28998);
nor UO_1006 (O_1006,N_29844,N_29862);
and UO_1007 (O_1007,N_29929,N_29778);
nor UO_1008 (O_1008,N_29689,N_29443);
nand UO_1009 (O_1009,N_29712,N_29714);
nor UO_1010 (O_1010,N_29016,N_29508);
nand UO_1011 (O_1011,N_28883,N_29519);
and UO_1012 (O_1012,N_29082,N_29701);
nor UO_1013 (O_1013,N_29644,N_29066);
xnor UO_1014 (O_1014,N_29428,N_28928);
nor UO_1015 (O_1015,N_29200,N_29672);
or UO_1016 (O_1016,N_29446,N_29487);
nor UO_1017 (O_1017,N_29200,N_29078);
xnor UO_1018 (O_1018,N_29737,N_29271);
and UO_1019 (O_1019,N_29086,N_29045);
or UO_1020 (O_1020,N_29148,N_29129);
and UO_1021 (O_1021,N_29969,N_28865);
and UO_1022 (O_1022,N_29755,N_28991);
xnor UO_1023 (O_1023,N_29636,N_28869);
nand UO_1024 (O_1024,N_29668,N_28922);
nor UO_1025 (O_1025,N_29192,N_29167);
nor UO_1026 (O_1026,N_29226,N_29237);
and UO_1027 (O_1027,N_29814,N_29049);
and UO_1028 (O_1028,N_29424,N_28978);
nor UO_1029 (O_1029,N_29332,N_29971);
and UO_1030 (O_1030,N_29623,N_29235);
xor UO_1031 (O_1031,N_29532,N_29528);
or UO_1032 (O_1032,N_29892,N_29765);
nand UO_1033 (O_1033,N_29651,N_29230);
nor UO_1034 (O_1034,N_29133,N_29671);
or UO_1035 (O_1035,N_29761,N_29619);
nand UO_1036 (O_1036,N_29409,N_28917);
nand UO_1037 (O_1037,N_28816,N_29243);
nor UO_1038 (O_1038,N_28811,N_29091);
nor UO_1039 (O_1039,N_29606,N_29579);
and UO_1040 (O_1040,N_29162,N_29798);
and UO_1041 (O_1041,N_29236,N_29026);
xor UO_1042 (O_1042,N_29269,N_29089);
nor UO_1043 (O_1043,N_28882,N_29043);
nor UO_1044 (O_1044,N_29310,N_29254);
and UO_1045 (O_1045,N_29242,N_28809);
xnor UO_1046 (O_1046,N_29806,N_29377);
and UO_1047 (O_1047,N_28957,N_29569);
nor UO_1048 (O_1048,N_29794,N_29254);
nor UO_1049 (O_1049,N_29620,N_29382);
and UO_1050 (O_1050,N_29853,N_29844);
nand UO_1051 (O_1051,N_29327,N_28876);
or UO_1052 (O_1052,N_29831,N_29400);
or UO_1053 (O_1053,N_28898,N_29763);
and UO_1054 (O_1054,N_29546,N_29032);
or UO_1055 (O_1055,N_29344,N_28862);
nor UO_1056 (O_1056,N_28884,N_29017);
and UO_1057 (O_1057,N_28979,N_29946);
or UO_1058 (O_1058,N_29182,N_28926);
or UO_1059 (O_1059,N_29531,N_29060);
nor UO_1060 (O_1060,N_28849,N_29818);
or UO_1061 (O_1061,N_29118,N_29675);
nand UO_1062 (O_1062,N_29088,N_29882);
or UO_1063 (O_1063,N_29834,N_29091);
nand UO_1064 (O_1064,N_29545,N_29179);
or UO_1065 (O_1065,N_29682,N_29894);
nor UO_1066 (O_1066,N_29370,N_29766);
and UO_1067 (O_1067,N_29995,N_29510);
xor UO_1068 (O_1068,N_29123,N_29307);
nand UO_1069 (O_1069,N_29442,N_29852);
xnor UO_1070 (O_1070,N_29264,N_28971);
xor UO_1071 (O_1071,N_29044,N_29881);
or UO_1072 (O_1072,N_29271,N_29375);
and UO_1073 (O_1073,N_29551,N_29326);
and UO_1074 (O_1074,N_29107,N_29048);
xor UO_1075 (O_1075,N_29045,N_29455);
and UO_1076 (O_1076,N_29343,N_29607);
nand UO_1077 (O_1077,N_29254,N_29051);
nand UO_1078 (O_1078,N_29363,N_29292);
xor UO_1079 (O_1079,N_29794,N_28859);
xnor UO_1080 (O_1080,N_29828,N_29284);
nor UO_1081 (O_1081,N_29272,N_28910);
nand UO_1082 (O_1082,N_29622,N_29458);
or UO_1083 (O_1083,N_29226,N_29150);
nor UO_1084 (O_1084,N_28825,N_29394);
and UO_1085 (O_1085,N_29346,N_29381);
or UO_1086 (O_1086,N_29666,N_29124);
nor UO_1087 (O_1087,N_29953,N_29251);
or UO_1088 (O_1088,N_29086,N_29078);
or UO_1089 (O_1089,N_28886,N_29994);
and UO_1090 (O_1090,N_29216,N_29616);
nor UO_1091 (O_1091,N_28936,N_29522);
xnor UO_1092 (O_1092,N_29272,N_29610);
and UO_1093 (O_1093,N_29700,N_29740);
nand UO_1094 (O_1094,N_29729,N_29989);
and UO_1095 (O_1095,N_29700,N_29624);
or UO_1096 (O_1096,N_29294,N_29361);
nand UO_1097 (O_1097,N_28835,N_28805);
xnor UO_1098 (O_1098,N_28837,N_28997);
and UO_1099 (O_1099,N_29675,N_28870);
nand UO_1100 (O_1100,N_29540,N_29330);
nand UO_1101 (O_1101,N_29075,N_28886);
xnor UO_1102 (O_1102,N_29301,N_29232);
and UO_1103 (O_1103,N_29866,N_29941);
nor UO_1104 (O_1104,N_28830,N_28956);
or UO_1105 (O_1105,N_29195,N_28940);
nand UO_1106 (O_1106,N_29416,N_29454);
or UO_1107 (O_1107,N_29331,N_29558);
or UO_1108 (O_1108,N_28895,N_29198);
nor UO_1109 (O_1109,N_29902,N_29640);
nor UO_1110 (O_1110,N_29240,N_29622);
and UO_1111 (O_1111,N_29604,N_29164);
nor UO_1112 (O_1112,N_28811,N_29277);
xnor UO_1113 (O_1113,N_29078,N_29725);
and UO_1114 (O_1114,N_29587,N_29550);
nor UO_1115 (O_1115,N_29003,N_29639);
and UO_1116 (O_1116,N_29222,N_29616);
and UO_1117 (O_1117,N_29306,N_29572);
xor UO_1118 (O_1118,N_29342,N_29028);
nor UO_1119 (O_1119,N_29874,N_29838);
nand UO_1120 (O_1120,N_29364,N_29766);
xnor UO_1121 (O_1121,N_29830,N_29773);
nand UO_1122 (O_1122,N_29246,N_29082);
xnor UO_1123 (O_1123,N_29880,N_29484);
and UO_1124 (O_1124,N_29665,N_28934);
nand UO_1125 (O_1125,N_29246,N_29874);
nor UO_1126 (O_1126,N_29849,N_29146);
nor UO_1127 (O_1127,N_29874,N_29456);
and UO_1128 (O_1128,N_29570,N_29372);
or UO_1129 (O_1129,N_28859,N_28824);
nor UO_1130 (O_1130,N_29879,N_29631);
xnor UO_1131 (O_1131,N_29929,N_29020);
nor UO_1132 (O_1132,N_28929,N_29172);
or UO_1133 (O_1133,N_29286,N_29156);
or UO_1134 (O_1134,N_28978,N_29260);
and UO_1135 (O_1135,N_29403,N_29673);
nor UO_1136 (O_1136,N_29865,N_29606);
or UO_1137 (O_1137,N_28939,N_28874);
xor UO_1138 (O_1138,N_29514,N_29445);
or UO_1139 (O_1139,N_29465,N_29082);
nor UO_1140 (O_1140,N_29371,N_29078);
xor UO_1141 (O_1141,N_29507,N_29563);
and UO_1142 (O_1142,N_29580,N_29328);
xnor UO_1143 (O_1143,N_29088,N_29730);
xnor UO_1144 (O_1144,N_29674,N_29949);
xor UO_1145 (O_1145,N_29937,N_29790);
nand UO_1146 (O_1146,N_28896,N_29809);
and UO_1147 (O_1147,N_29510,N_29416);
or UO_1148 (O_1148,N_28852,N_29137);
nand UO_1149 (O_1149,N_29108,N_29915);
nand UO_1150 (O_1150,N_29776,N_29030);
or UO_1151 (O_1151,N_29507,N_28955);
xnor UO_1152 (O_1152,N_29024,N_29629);
and UO_1153 (O_1153,N_29594,N_29830);
nand UO_1154 (O_1154,N_29579,N_29508);
nand UO_1155 (O_1155,N_29063,N_29111);
nand UO_1156 (O_1156,N_29944,N_29266);
or UO_1157 (O_1157,N_29481,N_29806);
nor UO_1158 (O_1158,N_29101,N_29517);
and UO_1159 (O_1159,N_29417,N_29987);
xor UO_1160 (O_1160,N_29953,N_29717);
and UO_1161 (O_1161,N_29087,N_29954);
nor UO_1162 (O_1162,N_29161,N_29082);
xor UO_1163 (O_1163,N_29734,N_29214);
and UO_1164 (O_1164,N_29662,N_29044);
xor UO_1165 (O_1165,N_29078,N_29564);
nand UO_1166 (O_1166,N_29131,N_28863);
or UO_1167 (O_1167,N_29942,N_29538);
xnor UO_1168 (O_1168,N_29650,N_29244);
nor UO_1169 (O_1169,N_29113,N_29084);
or UO_1170 (O_1170,N_29648,N_28929);
xnor UO_1171 (O_1171,N_28954,N_29217);
nor UO_1172 (O_1172,N_28852,N_29504);
nand UO_1173 (O_1173,N_28944,N_29079);
nand UO_1174 (O_1174,N_29251,N_28883);
or UO_1175 (O_1175,N_29624,N_29561);
nand UO_1176 (O_1176,N_29113,N_29603);
xor UO_1177 (O_1177,N_29373,N_29098);
nand UO_1178 (O_1178,N_29043,N_29977);
or UO_1179 (O_1179,N_28811,N_29070);
or UO_1180 (O_1180,N_29140,N_29234);
and UO_1181 (O_1181,N_29567,N_29218);
and UO_1182 (O_1182,N_29091,N_29498);
and UO_1183 (O_1183,N_29987,N_29548);
and UO_1184 (O_1184,N_28819,N_29978);
nor UO_1185 (O_1185,N_29865,N_29287);
nor UO_1186 (O_1186,N_29746,N_29140);
nor UO_1187 (O_1187,N_29779,N_29881);
nand UO_1188 (O_1188,N_28879,N_29969);
nor UO_1189 (O_1189,N_28901,N_29200);
and UO_1190 (O_1190,N_28864,N_29705);
and UO_1191 (O_1191,N_28885,N_29671);
and UO_1192 (O_1192,N_29977,N_29540);
or UO_1193 (O_1193,N_29397,N_29498);
nand UO_1194 (O_1194,N_29988,N_29690);
and UO_1195 (O_1195,N_29767,N_28848);
nand UO_1196 (O_1196,N_29063,N_28829);
nor UO_1197 (O_1197,N_29317,N_29988);
nor UO_1198 (O_1198,N_29338,N_29759);
nand UO_1199 (O_1199,N_29446,N_28803);
xnor UO_1200 (O_1200,N_29074,N_29899);
nor UO_1201 (O_1201,N_29216,N_29868);
nor UO_1202 (O_1202,N_29648,N_29635);
xor UO_1203 (O_1203,N_29640,N_29557);
nand UO_1204 (O_1204,N_29564,N_29293);
or UO_1205 (O_1205,N_29863,N_29189);
xor UO_1206 (O_1206,N_29421,N_29513);
nand UO_1207 (O_1207,N_29623,N_29915);
nand UO_1208 (O_1208,N_29018,N_29062);
nand UO_1209 (O_1209,N_29254,N_28857);
xor UO_1210 (O_1210,N_29834,N_29330);
and UO_1211 (O_1211,N_29464,N_28940);
xor UO_1212 (O_1212,N_28900,N_29528);
xnor UO_1213 (O_1213,N_29439,N_29102);
xor UO_1214 (O_1214,N_29292,N_29591);
xnor UO_1215 (O_1215,N_29567,N_29870);
nor UO_1216 (O_1216,N_29624,N_29081);
and UO_1217 (O_1217,N_29537,N_28831);
and UO_1218 (O_1218,N_29390,N_29831);
nor UO_1219 (O_1219,N_29210,N_29754);
or UO_1220 (O_1220,N_29169,N_29878);
or UO_1221 (O_1221,N_28986,N_29242);
nor UO_1222 (O_1222,N_29205,N_29492);
nor UO_1223 (O_1223,N_29715,N_28861);
or UO_1224 (O_1224,N_28997,N_29305);
nor UO_1225 (O_1225,N_29170,N_29420);
nor UO_1226 (O_1226,N_28914,N_29130);
nor UO_1227 (O_1227,N_29339,N_28866);
or UO_1228 (O_1228,N_29545,N_29492);
nor UO_1229 (O_1229,N_29142,N_29024);
xnor UO_1230 (O_1230,N_29725,N_29152);
or UO_1231 (O_1231,N_29030,N_28888);
nor UO_1232 (O_1232,N_29516,N_29828);
or UO_1233 (O_1233,N_29918,N_28906);
nand UO_1234 (O_1234,N_28825,N_29914);
and UO_1235 (O_1235,N_29563,N_28958);
nor UO_1236 (O_1236,N_29876,N_29010);
or UO_1237 (O_1237,N_29717,N_29674);
and UO_1238 (O_1238,N_29393,N_29183);
or UO_1239 (O_1239,N_29952,N_29488);
or UO_1240 (O_1240,N_29179,N_29448);
xnor UO_1241 (O_1241,N_29439,N_29062);
nand UO_1242 (O_1242,N_28810,N_29091);
xor UO_1243 (O_1243,N_29486,N_29116);
or UO_1244 (O_1244,N_29191,N_29011);
or UO_1245 (O_1245,N_29554,N_29365);
xnor UO_1246 (O_1246,N_29202,N_29292);
nand UO_1247 (O_1247,N_29831,N_29625);
nand UO_1248 (O_1248,N_28917,N_29767);
nand UO_1249 (O_1249,N_29849,N_29514);
nor UO_1250 (O_1250,N_29977,N_29687);
nand UO_1251 (O_1251,N_28962,N_29780);
xor UO_1252 (O_1252,N_29357,N_29482);
xnor UO_1253 (O_1253,N_29579,N_28853);
and UO_1254 (O_1254,N_29622,N_29856);
nor UO_1255 (O_1255,N_29159,N_29903);
nand UO_1256 (O_1256,N_29711,N_28986);
nor UO_1257 (O_1257,N_29432,N_29719);
xnor UO_1258 (O_1258,N_29712,N_29878);
xnor UO_1259 (O_1259,N_29129,N_28804);
nor UO_1260 (O_1260,N_28859,N_29607);
or UO_1261 (O_1261,N_29167,N_29718);
and UO_1262 (O_1262,N_29070,N_29536);
nand UO_1263 (O_1263,N_29667,N_29641);
xor UO_1264 (O_1264,N_29808,N_28894);
or UO_1265 (O_1265,N_29593,N_28815);
nand UO_1266 (O_1266,N_29107,N_29219);
and UO_1267 (O_1267,N_29417,N_29770);
and UO_1268 (O_1268,N_29097,N_29837);
and UO_1269 (O_1269,N_29293,N_29887);
nand UO_1270 (O_1270,N_29346,N_29059);
and UO_1271 (O_1271,N_29093,N_29392);
and UO_1272 (O_1272,N_28979,N_29194);
nand UO_1273 (O_1273,N_29160,N_29225);
or UO_1274 (O_1274,N_29171,N_29719);
xnor UO_1275 (O_1275,N_29777,N_29266);
and UO_1276 (O_1276,N_29254,N_28966);
or UO_1277 (O_1277,N_29895,N_29818);
nand UO_1278 (O_1278,N_28824,N_29366);
or UO_1279 (O_1279,N_29491,N_29249);
xnor UO_1280 (O_1280,N_28977,N_29742);
xnor UO_1281 (O_1281,N_29867,N_29643);
and UO_1282 (O_1282,N_29345,N_29592);
or UO_1283 (O_1283,N_29495,N_29829);
nand UO_1284 (O_1284,N_29967,N_29021);
and UO_1285 (O_1285,N_29148,N_29701);
nor UO_1286 (O_1286,N_29239,N_29240);
and UO_1287 (O_1287,N_29265,N_28892);
and UO_1288 (O_1288,N_29524,N_28992);
and UO_1289 (O_1289,N_29922,N_29231);
xnor UO_1290 (O_1290,N_28816,N_29774);
or UO_1291 (O_1291,N_29163,N_29958);
and UO_1292 (O_1292,N_29093,N_29520);
or UO_1293 (O_1293,N_29027,N_29864);
and UO_1294 (O_1294,N_29001,N_28963);
or UO_1295 (O_1295,N_29154,N_29603);
or UO_1296 (O_1296,N_29713,N_29145);
and UO_1297 (O_1297,N_28827,N_29480);
and UO_1298 (O_1298,N_28880,N_29225);
and UO_1299 (O_1299,N_29580,N_28979);
and UO_1300 (O_1300,N_29085,N_29303);
and UO_1301 (O_1301,N_29395,N_29263);
nor UO_1302 (O_1302,N_28966,N_29513);
nor UO_1303 (O_1303,N_28837,N_28985);
xnor UO_1304 (O_1304,N_29010,N_29472);
and UO_1305 (O_1305,N_29620,N_29750);
nand UO_1306 (O_1306,N_29995,N_29406);
nand UO_1307 (O_1307,N_29344,N_29368);
nand UO_1308 (O_1308,N_29310,N_28969);
nor UO_1309 (O_1309,N_29977,N_29722);
or UO_1310 (O_1310,N_29212,N_28931);
xnor UO_1311 (O_1311,N_29160,N_29156);
nor UO_1312 (O_1312,N_28846,N_29821);
xor UO_1313 (O_1313,N_29839,N_28902);
nand UO_1314 (O_1314,N_29623,N_29425);
or UO_1315 (O_1315,N_29428,N_28995);
nor UO_1316 (O_1316,N_29046,N_29693);
and UO_1317 (O_1317,N_29228,N_29741);
nor UO_1318 (O_1318,N_29575,N_29521);
xnor UO_1319 (O_1319,N_29207,N_29460);
or UO_1320 (O_1320,N_29538,N_29013);
xnor UO_1321 (O_1321,N_29985,N_28834);
and UO_1322 (O_1322,N_29661,N_29368);
nor UO_1323 (O_1323,N_29226,N_29662);
and UO_1324 (O_1324,N_28948,N_29632);
xnor UO_1325 (O_1325,N_29451,N_29018);
and UO_1326 (O_1326,N_29316,N_29156);
nor UO_1327 (O_1327,N_28911,N_28830);
and UO_1328 (O_1328,N_28900,N_29169);
nor UO_1329 (O_1329,N_29878,N_29735);
or UO_1330 (O_1330,N_29639,N_29318);
and UO_1331 (O_1331,N_29906,N_29140);
nand UO_1332 (O_1332,N_29579,N_29573);
nor UO_1333 (O_1333,N_29567,N_29997);
or UO_1334 (O_1334,N_28892,N_29974);
nor UO_1335 (O_1335,N_29219,N_29723);
xor UO_1336 (O_1336,N_29010,N_29866);
xnor UO_1337 (O_1337,N_29409,N_29586);
nor UO_1338 (O_1338,N_29563,N_29939);
nor UO_1339 (O_1339,N_29009,N_29246);
or UO_1340 (O_1340,N_28940,N_29566);
and UO_1341 (O_1341,N_29356,N_29662);
and UO_1342 (O_1342,N_29307,N_29495);
xor UO_1343 (O_1343,N_29623,N_29719);
and UO_1344 (O_1344,N_28950,N_28869);
nand UO_1345 (O_1345,N_29454,N_29874);
xor UO_1346 (O_1346,N_29756,N_29118);
or UO_1347 (O_1347,N_29915,N_29604);
xnor UO_1348 (O_1348,N_29274,N_29090);
or UO_1349 (O_1349,N_28989,N_29861);
nand UO_1350 (O_1350,N_29430,N_29335);
nand UO_1351 (O_1351,N_29006,N_29017);
or UO_1352 (O_1352,N_29877,N_29737);
or UO_1353 (O_1353,N_29994,N_29426);
or UO_1354 (O_1354,N_29958,N_29002);
xnor UO_1355 (O_1355,N_29901,N_29020);
or UO_1356 (O_1356,N_29525,N_28845);
nand UO_1357 (O_1357,N_28843,N_28994);
nor UO_1358 (O_1358,N_29502,N_28903);
nand UO_1359 (O_1359,N_28814,N_29000);
or UO_1360 (O_1360,N_29603,N_29240);
or UO_1361 (O_1361,N_29123,N_28902);
and UO_1362 (O_1362,N_29251,N_29961);
nor UO_1363 (O_1363,N_29129,N_29197);
or UO_1364 (O_1364,N_28937,N_29726);
or UO_1365 (O_1365,N_29587,N_28852);
nand UO_1366 (O_1366,N_29911,N_28839);
xor UO_1367 (O_1367,N_28830,N_29417);
and UO_1368 (O_1368,N_28890,N_29768);
and UO_1369 (O_1369,N_29755,N_29895);
and UO_1370 (O_1370,N_29268,N_29062);
nand UO_1371 (O_1371,N_29044,N_29160);
nand UO_1372 (O_1372,N_29051,N_29188);
nand UO_1373 (O_1373,N_29275,N_29504);
nor UO_1374 (O_1374,N_29905,N_29406);
and UO_1375 (O_1375,N_29306,N_29845);
or UO_1376 (O_1376,N_29474,N_29361);
nand UO_1377 (O_1377,N_28838,N_29846);
and UO_1378 (O_1378,N_29369,N_28890);
or UO_1379 (O_1379,N_29994,N_29921);
xnor UO_1380 (O_1380,N_29666,N_29804);
xnor UO_1381 (O_1381,N_29477,N_28905);
and UO_1382 (O_1382,N_29966,N_29434);
nor UO_1383 (O_1383,N_29395,N_29795);
xnor UO_1384 (O_1384,N_28968,N_29702);
xor UO_1385 (O_1385,N_29055,N_28914);
and UO_1386 (O_1386,N_28936,N_29443);
xnor UO_1387 (O_1387,N_29035,N_28877);
or UO_1388 (O_1388,N_29508,N_29264);
and UO_1389 (O_1389,N_28996,N_29388);
nand UO_1390 (O_1390,N_29602,N_29355);
nor UO_1391 (O_1391,N_29373,N_29820);
xnor UO_1392 (O_1392,N_29407,N_29598);
or UO_1393 (O_1393,N_28815,N_29475);
or UO_1394 (O_1394,N_29834,N_29236);
nand UO_1395 (O_1395,N_29723,N_29332);
xnor UO_1396 (O_1396,N_29171,N_29320);
xor UO_1397 (O_1397,N_29661,N_29154);
or UO_1398 (O_1398,N_29398,N_29840);
nand UO_1399 (O_1399,N_29267,N_29673);
nor UO_1400 (O_1400,N_29439,N_28814);
xnor UO_1401 (O_1401,N_29530,N_29933);
nor UO_1402 (O_1402,N_29934,N_29891);
nor UO_1403 (O_1403,N_28901,N_28816);
xor UO_1404 (O_1404,N_29726,N_29891);
nand UO_1405 (O_1405,N_29777,N_29739);
xor UO_1406 (O_1406,N_29157,N_28802);
xor UO_1407 (O_1407,N_29895,N_29252);
nor UO_1408 (O_1408,N_28947,N_29111);
nor UO_1409 (O_1409,N_28914,N_29053);
nand UO_1410 (O_1410,N_29930,N_28935);
nor UO_1411 (O_1411,N_29503,N_29462);
nand UO_1412 (O_1412,N_29701,N_28807);
nor UO_1413 (O_1413,N_29686,N_28957);
xor UO_1414 (O_1414,N_29097,N_29465);
xor UO_1415 (O_1415,N_29005,N_29156);
or UO_1416 (O_1416,N_29174,N_29682);
or UO_1417 (O_1417,N_28814,N_28843);
nor UO_1418 (O_1418,N_29919,N_29855);
and UO_1419 (O_1419,N_29872,N_29159);
nand UO_1420 (O_1420,N_28925,N_29103);
and UO_1421 (O_1421,N_29953,N_29306);
or UO_1422 (O_1422,N_29060,N_29576);
nand UO_1423 (O_1423,N_29410,N_29178);
nor UO_1424 (O_1424,N_28838,N_29300);
nor UO_1425 (O_1425,N_29651,N_28864);
nand UO_1426 (O_1426,N_29510,N_29089);
or UO_1427 (O_1427,N_29734,N_29733);
nor UO_1428 (O_1428,N_29992,N_29477);
nor UO_1429 (O_1429,N_29634,N_29555);
or UO_1430 (O_1430,N_29682,N_29298);
nand UO_1431 (O_1431,N_29293,N_29204);
or UO_1432 (O_1432,N_29900,N_29546);
xor UO_1433 (O_1433,N_29851,N_29678);
nand UO_1434 (O_1434,N_29560,N_29712);
nor UO_1435 (O_1435,N_29019,N_29763);
xnor UO_1436 (O_1436,N_29016,N_29862);
xnor UO_1437 (O_1437,N_28901,N_28890);
nand UO_1438 (O_1438,N_28988,N_29239);
xor UO_1439 (O_1439,N_29598,N_29792);
and UO_1440 (O_1440,N_29513,N_29662);
nor UO_1441 (O_1441,N_29534,N_29753);
or UO_1442 (O_1442,N_29697,N_29427);
and UO_1443 (O_1443,N_29105,N_29678);
and UO_1444 (O_1444,N_28855,N_28865);
nor UO_1445 (O_1445,N_29708,N_29556);
nor UO_1446 (O_1446,N_29638,N_28963);
and UO_1447 (O_1447,N_29699,N_29838);
xor UO_1448 (O_1448,N_29746,N_28838);
or UO_1449 (O_1449,N_29254,N_29240);
xnor UO_1450 (O_1450,N_29898,N_29895);
nand UO_1451 (O_1451,N_29361,N_29164);
nand UO_1452 (O_1452,N_29453,N_29013);
xnor UO_1453 (O_1453,N_29983,N_29616);
nor UO_1454 (O_1454,N_29461,N_29920);
nor UO_1455 (O_1455,N_29572,N_29999);
and UO_1456 (O_1456,N_28983,N_29256);
nand UO_1457 (O_1457,N_29655,N_29172);
nor UO_1458 (O_1458,N_29696,N_29289);
nand UO_1459 (O_1459,N_29215,N_28806);
nor UO_1460 (O_1460,N_29576,N_29164);
or UO_1461 (O_1461,N_28808,N_29543);
xnor UO_1462 (O_1462,N_29879,N_29227);
nor UO_1463 (O_1463,N_29038,N_28805);
nand UO_1464 (O_1464,N_29169,N_29503);
or UO_1465 (O_1465,N_29580,N_28926);
nand UO_1466 (O_1466,N_29788,N_29965);
xnor UO_1467 (O_1467,N_29220,N_29989);
and UO_1468 (O_1468,N_29373,N_29484);
nand UO_1469 (O_1469,N_28848,N_29185);
and UO_1470 (O_1470,N_29787,N_29763);
and UO_1471 (O_1471,N_29279,N_29867);
and UO_1472 (O_1472,N_28902,N_29396);
and UO_1473 (O_1473,N_28862,N_29545);
or UO_1474 (O_1474,N_29929,N_29492);
nand UO_1475 (O_1475,N_29766,N_29353);
xnor UO_1476 (O_1476,N_29031,N_29949);
xnor UO_1477 (O_1477,N_29946,N_29616);
nand UO_1478 (O_1478,N_29164,N_29831);
nor UO_1479 (O_1479,N_29195,N_29689);
and UO_1480 (O_1480,N_29621,N_29739);
nand UO_1481 (O_1481,N_29869,N_29412);
nor UO_1482 (O_1482,N_28942,N_29602);
nand UO_1483 (O_1483,N_29058,N_29255);
and UO_1484 (O_1484,N_29738,N_29651);
nor UO_1485 (O_1485,N_29439,N_28815);
nor UO_1486 (O_1486,N_29237,N_29608);
nand UO_1487 (O_1487,N_29150,N_28824);
nand UO_1488 (O_1488,N_29182,N_29515);
nand UO_1489 (O_1489,N_29100,N_29443);
nor UO_1490 (O_1490,N_29454,N_28898);
nand UO_1491 (O_1491,N_28909,N_29962);
nor UO_1492 (O_1492,N_29541,N_28852);
and UO_1493 (O_1493,N_29828,N_29208);
and UO_1494 (O_1494,N_29145,N_29179);
xnor UO_1495 (O_1495,N_29026,N_29016);
nor UO_1496 (O_1496,N_29150,N_29779);
and UO_1497 (O_1497,N_28990,N_29189);
xor UO_1498 (O_1498,N_29534,N_29274);
and UO_1499 (O_1499,N_29827,N_28846);
xor UO_1500 (O_1500,N_29526,N_29015);
xor UO_1501 (O_1501,N_28946,N_29022);
nand UO_1502 (O_1502,N_29898,N_29350);
and UO_1503 (O_1503,N_29664,N_29536);
and UO_1504 (O_1504,N_29849,N_29311);
and UO_1505 (O_1505,N_29007,N_29998);
nor UO_1506 (O_1506,N_29017,N_29000);
xnor UO_1507 (O_1507,N_29547,N_28937);
nand UO_1508 (O_1508,N_29183,N_29908);
nor UO_1509 (O_1509,N_29307,N_29648);
or UO_1510 (O_1510,N_29483,N_29611);
nand UO_1511 (O_1511,N_29038,N_28963);
nand UO_1512 (O_1512,N_28973,N_29338);
nand UO_1513 (O_1513,N_29503,N_29149);
xnor UO_1514 (O_1514,N_29104,N_29142);
xor UO_1515 (O_1515,N_29135,N_28881);
nor UO_1516 (O_1516,N_29033,N_29152);
or UO_1517 (O_1517,N_29274,N_29278);
nand UO_1518 (O_1518,N_29109,N_29431);
and UO_1519 (O_1519,N_29852,N_28912);
nand UO_1520 (O_1520,N_29141,N_29026);
or UO_1521 (O_1521,N_29965,N_29425);
and UO_1522 (O_1522,N_29841,N_29346);
nand UO_1523 (O_1523,N_29207,N_28849);
nand UO_1524 (O_1524,N_28861,N_29948);
nor UO_1525 (O_1525,N_29183,N_29485);
xnor UO_1526 (O_1526,N_29196,N_29763);
and UO_1527 (O_1527,N_29273,N_29868);
and UO_1528 (O_1528,N_28914,N_29735);
or UO_1529 (O_1529,N_29680,N_29071);
nand UO_1530 (O_1530,N_29786,N_29507);
or UO_1531 (O_1531,N_28833,N_29767);
xnor UO_1532 (O_1532,N_28853,N_29613);
and UO_1533 (O_1533,N_28825,N_29454);
and UO_1534 (O_1534,N_29740,N_29744);
nand UO_1535 (O_1535,N_29529,N_29783);
or UO_1536 (O_1536,N_29037,N_28995);
nor UO_1537 (O_1537,N_29253,N_29121);
xor UO_1538 (O_1538,N_29169,N_28929);
nand UO_1539 (O_1539,N_29523,N_29533);
xnor UO_1540 (O_1540,N_29840,N_29357);
or UO_1541 (O_1541,N_29040,N_29860);
xnor UO_1542 (O_1542,N_29313,N_29740);
xnor UO_1543 (O_1543,N_29343,N_29812);
xor UO_1544 (O_1544,N_29627,N_29574);
nand UO_1545 (O_1545,N_29975,N_29022);
xnor UO_1546 (O_1546,N_29620,N_28888);
xnor UO_1547 (O_1547,N_29701,N_29114);
and UO_1548 (O_1548,N_29750,N_29343);
nand UO_1549 (O_1549,N_29266,N_29984);
nor UO_1550 (O_1550,N_29907,N_28933);
nor UO_1551 (O_1551,N_29133,N_29159);
or UO_1552 (O_1552,N_29263,N_28947);
nand UO_1553 (O_1553,N_29680,N_29995);
xnor UO_1554 (O_1554,N_29529,N_28982);
xor UO_1555 (O_1555,N_29529,N_29823);
xnor UO_1556 (O_1556,N_28903,N_28911);
xnor UO_1557 (O_1557,N_29620,N_29888);
or UO_1558 (O_1558,N_29224,N_28895);
nor UO_1559 (O_1559,N_29716,N_29659);
and UO_1560 (O_1560,N_28902,N_29407);
and UO_1561 (O_1561,N_29545,N_29586);
and UO_1562 (O_1562,N_29352,N_29398);
and UO_1563 (O_1563,N_29730,N_29595);
xnor UO_1564 (O_1564,N_29019,N_29585);
or UO_1565 (O_1565,N_29420,N_29998);
xnor UO_1566 (O_1566,N_29257,N_29347);
nor UO_1567 (O_1567,N_29813,N_29438);
nand UO_1568 (O_1568,N_29622,N_28808);
and UO_1569 (O_1569,N_29658,N_29628);
and UO_1570 (O_1570,N_29956,N_29494);
nand UO_1571 (O_1571,N_29623,N_29042);
xor UO_1572 (O_1572,N_29433,N_29149);
nand UO_1573 (O_1573,N_29811,N_29720);
nand UO_1574 (O_1574,N_28827,N_29238);
nor UO_1575 (O_1575,N_29959,N_29739);
or UO_1576 (O_1576,N_29935,N_29804);
nor UO_1577 (O_1577,N_28930,N_28992);
nor UO_1578 (O_1578,N_29637,N_29189);
and UO_1579 (O_1579,N_29730,N_29545);
nand UO_1580 (O_1580,N_29427,N_28966);
nor UO_1581 (O_1581,N_29505,N_28824);
xor UO_1582 (O_1582,N_29977,N_29904);
or UO_1583 (O_1583,N_29638,N_28989);
nor UO_1584 (O_1584,N_29847,N_29162);
or UO_1585 (O_1585,N_29915,N_29988);
nand UO_1586 (O_1586,N_29608,N_28967);
nand UO_1587 (O_1587,N_29381,N_29059);
or UO_1588 (O_1588,N_28882,N_29447);
or UO_1589 (O_1589,N_29244,N_29170);
or UO_1590 (O_1590,N_29488,N_29789);
and UO_1591 (O_1591,N_29092,N_28860);
nor UO_1592 (O_1592,N_29963,N_29202);
nor UO_1593 (O_1593,N_29965,N_28874);
or UO_1594 (O_1594,N_28895,N_29374);
or UO_1595 (O_1595,N_29233,N_29330);
and UO_1596 (O_1596,N_28833,N_29278);
or UO_1597 (O_1597,N_29091,N_29906);
or UO_1598 (O_1598,N_29443,N_29868);
or UO_1599 (O_1599,N_29393,N_29632);
nor UO_1600 (O_1600,N_29715,N_29708);
xor UO_1601 (O_1601,N_29244,N_29131);
nand UO_1602 (O_1602,N_29554,N_28922);
nor UO_1603 (O_1603,N_29545,N_29828);
and UO_1604 (O_1604,N_29734,N_29131);
nand UO_1605 (O_1605,N_28808,N_29942);
or UO_1606 (O_1606,N_29184,N_29680);
xor UO_1607 (O_1607,N_29239,N_29634);
or UO_1608 (O_1608,N_29683,N_29418);
and UO_1609 (O_1609,N_29092,N_29791);
nor UO_1610 (O_1610,N_29956,N_29593);
nand UO_1611 (O_1611,N_28886,N_29767);
xnor UO_1612 (O_1612,N_29479,N_28815);
nor UO_1613 (O_1613,N_28986,N_29118);
nor UO_1614 (O_1614,N_29381,N_29439);
xnor UO_1615 (O_1615,N_28832,N_29438);
nand UO_1616 (O_1616,N_29397,N_29810);
nor UO_1617 (O_1617,N_29656,N_28883);
nand UO_1618 (O_1618,N_28963,N_29402);
and UO_1619 (O_1619,N_28835,N_29642);
or UO_1620 (O_1620,N_29206,N_29699);
or UO_1621 (O_1621,N_29787,N_29094);
or UO_1622 (O_1622,N_29044,N_28906);
and UO_1623 (O_1623,N_29499,N_29525);
nor UO_1624 (O_1624,N_29136,N_29672);
or UO_1625 (O_1625,N_29525,N_29771);
nor UO_1626 (O_1626,N_28814,N_29578);
nand UO_1627 (O_1627,N_29930,N_29419);
xor UO_1628 (O_1628,N_29471,N_29963);
nand UO_1629 (O_1629,N_29768,N_28827);
nand UO_1630 (O_1630,N_29951,N_28989);
or UO_1631 (O_1631,N_29103,N_28889);
nand UO_1632 (O_1632,N_29369,N_29270);
nor UO_1633 (O_1633,N_29839,N_29078);
and UO_1634 (O_1634,N_29585,N_29633);
xor UO_1635 (O_1635,N_29762,N_29624);
and UO_1636 (O_1636,N_29670,N_29792);
xor UO_1637 (O_1637,N_29617,N_29753);
xnor UO_1638 (O_1638,N_29467,N_29262);
and UO_1639 (O_1639,N_29722,N_28967);
and UO_1640 (O_1640,N_29137,N_29123);
nor UO_1641 (O_1641,N_29182,N_29952);
or UO_1642 (O_1642,N_28861,N_29549);
or UO_1643 (O_1643,N_29218,N_29467);
or UO_1644 (O_1644,N_29083,N_28846);
and UO_1645 (O_1645,N_28847,N_29766);
nand UO_1646 (O_1646,N_28965,N_29431);
nor UO_1647 (O_1647,N_29169,N_29702);
and UO_1648 (O_1648,N_29475,N_29635);
nand UO_1649 (O_1649,N_29323,N_28977);
and UO_1650 (O_1650,N_29810,N_29864);
nand UO_1651 (O_1651,N_28805,N_28924);
nor UO_1652 (O_1652,N_29127,N_29659);
or UO_1653 (O_1653,N_28830,N_29559);
nor UO_1654 (O_1654,N_28843,N_29739);
xor UO_1655 (O_1655,N_29535,N_29578);
nand UO_1656 (O_1656,N_28834,N_29935);
nor UO_1657 (O_1657,N_29751,N_29491);
xor UO_1658 (O_1658,N_28962,N_29596);
or UO_1659 (O_1659,N_29221,N_29749);
nand UO_1660 (O_1660,N_29462,N_29915);
and UO_1661 (O_1661,N_29879,N_29237);
xnor UO_1662 (O_1662,N_29822,N_28889);
or UO_1663 (O_1663,N_29833,N_28928);
xnor UO_1664 (O_1664,N_29788,N_28802);
nor UO_1665 (O_1665,N_29167,N_29876);
and UO_1666 (O_1666,N_29297,N_29906);
xnor UO_1667 (O_1667,N_29563,N_29887);
nor UO_1668 (O_1668,N_28867,N_29190);
or UO_1669 (O_1669,N_29873,N_29809);
and UO_1670 (O_1670,N_29751,N_29408);
xor UO_1671 (O_1671,N_29654,N_29662);
xnor UO_1672 (O_1672,N_29172,N_29219);
nor UO_1673 (O_1673,N_29394,N_29419);
xor UO_1674 (O_1674,N_29729,N_29578);
nand UO_1675 (O_1675,N_29652,N_28936);
or UO_1676 (O_1676,N_29804,N_29879);
or UO_1677 (O_1677,N_28819,N_28953);
nor UO_1678 (O_1678,N_29460,N_29227);
or UO_1679 (O_1679,N_29985,N_29278);
or UO_1680 (O_1680,N_29361,N_29435);
nand UO_1681 (O_1681,N_29923,N_29224);
xnor UO_1682 (O_1682,N_29644,N_29717);
or UO_1683 (O_1683,N_29670,N_29912);
nand UO_1684 (O_1684,N_29257,N_29062);
and UO_1685 (O_1685,N_29363,N_29319);
and UO_1686 (O_1686,N_29710,N_29364);
nor UO_1687 (O_1687,N_29161,N_29052);
or UO_1688 (O_1688,N_28845,N_29833);
xnor UO_1689 (O_1689,N_29191,N_29228);
xor UO_1690 (O_1690,N_29159,N_29198);
and UO_1691 (O_1691,N_28837,N_29904);
xnor UO_1692 (O_1692,N_29325,N_29794);
nor UO_1693 (O_1693,N_29516,N_28947);
nand UO_1694 (O_1694,N_29956,N_29578);
or UO_1695 (O_1695,N_29704,N_29573);
and UO_1696 (O_1696,N_28981,N_29963);
nor UO_1697 (O_1697,N_29324,N_29535);
nand UO_1698 (O_1698,N_29456,N_29135);
or UO_1699 (O_1699,N_29836,N_29049);
or UO_1700 (O_1700,N_29611,N_29336);
xnor UO_1701 (O_1701,N_29565,N_28871);
nor UO_1702 (O_1702,N_29945,N_29266);
or UO_1703 (O_1703,N_29464,N_29130);
nand UO_1704 (O_1704,N_28882,N_28810);
nor UO_1705 (O_1705,N_29906,N_29747);
and UO_1706 (O_1706,N_29985,N_29698);
or UO_1707 (O_1707,N_29914,N_29642);
and UO_1708 (O_1708,N_29502,N_29472);
nor UO_1709 (O_1709,N_29462,N_29839);
nand UO_1710 (O_1710,N_29298,N_29725);
and UO_1711 (O_1711,N_28975,N_29407);
and UO_1712 (O_1712,N_29898,N_28990);
or UO_1713 (O_1713,N_29056,N_28914);
or UO_1714 (O_1714,N_29197,N_29235);
xnor UO_1715 (O_1715,N_29460,N_29233);
or UO_1716 (O_1716,N_29212,N_29848);
or UO_1717 (O_1717,N_29394,N_29978);
or UO_1718 (O_1718,N_29352,N_29753);
nor UO_1719 (O_1719,N_29022,N_28986);
nand UO_1720 (O_1720,N_29607,N_29284);
or UO_1721 (O_1721,N_29096,N_29022);
and UO_1722 (O_1722,N_29389,N_29594);
and UO_1723 (O_1723,N_29710,N_29075);
nor UO_1724 (O_1724,N_29803,N_29201);
nor UO_1725 (O_1725,N_29191,N_28828);
or UO_1726 (O_1726,N_29567,N_29146);
nand UO_1727 (O_1727,N_29672,N_29932);
and UO_1728 (O_1728,N_29780,N_29943);
or UO_1729 (O_1729,N_29036,N_29564);
or UO_1730 (O_1730,N_29327,N_29883);
nand UO_1731 (O_1731,N_29785,N_29947);
xor UO_1732 (O_1732,N_29691,N_29955);
xnor UO_1733 (O_1733,N_29756,N_29816);
nor UO_1734 (O_1734,N_29642,N_29014);
or UO_1735 (O_1735,N_28907,N_29109);
xnor UO_1736 (O_1736,N_29629,N_28866);
nor UO_1737 (O_1737,N_29502,N_29930);
or UO_1738 (O_1738,N_29242,N_28903);
xor UO_1739 (O_1739,N_29583,N_29972);
xnor UO_1740 (O_1740,N_29952,N_29898);
nand UO_1741 (O_1741,N_29912,N_28935);
nor UO_1742 (O_1742,N_29322,N_29133);
or UO_1743 (O_1743,N_29870,N_29469);
xnor UO_1744 (O_1744,N_29242,N_29060);
and UO_1745 (O_1745,N_29186,N_28921);
or UO_1746 (O_1746,N_29242,N_29012);
nand UO_1747 (O_1747,N_29941,N_29057);
xor UO_1748 (O_1748,N_29461,N_29805);
nor UO_1749 (O_1749,N_29671,N_29612);
and UO_1750 (O_1750,N_28826,N_29523);
or UO_1751 (O_1751,N_28913,N_29264);
and UO_1752 (O_1752,N_29482,N_29011);
and UO_1753 (O_1753,N_29196,N_28834);
nor UO_1754 (O_1754,N_29304,N_29229);
nor UO_1755 (O_1755,N_29824,N_28901);
nor UO_1756 (O_1756,N_29606,N_28921);
nor UO_1757 (O_1757,N_29537,N_29372);
nor UO_1758 (O_1758,N_29521,N_29323);
nand UO_1759 (O_1759,N_29169,N_29237);
and UO_1760 (O_1760,N_29627,N_29864);
and UO_1761 (O_1761,N_28876,N_29081);
nand UO_1762 (O_1762,N_29202,N_29160);
nand UO_1763 (O_1763,N_28837,N_29836);
nor UO_1764 (O_1764,N_29100,N_29696);
or UO_1765 (O_1765,N_29925,N_29559);
nand UO_1766 (O_1766,N_28925,N_29025);
nor UO_1767 (O_1767,N_29904,N_29618);
nand UO_1768 (O_1768,N_29612,N_29018);
nor UO_1769 (O_1769,N_29176,N_29000);
nor UO_1770 (O_1770,N_29636,N_28936);
nand UO_1771 (O_1771,N_29666,N_29484);
and UO_1772 (O_1772,N_29961,N_28941);
nand UO_1773 (O_1773,N_29119,N_29729);
or UO_1774 (O_1774,N_29396,N_29678);
and UO_1775 (O_1775,N_29384,N_29929);
nor UO_1776 (O_1776,N_29574,N_29342);
nand UO_1777 (O_1777,N_28940,N_28931);
nand UO_1778 (O_1778,N_29955,N_29343);
nor UO_1779 (O_1779,N_29193,N_28808);
nand UO_1780 (O_1780,N_29008,N_29384);
and UO_1781 (O_1781,N_28820,N_29820);
or UO_1782 (O_1782,N_29451,N_29691);
nor UO_1783 (O_1783,N_29875,N_29861);
and UO_1784 (O_1784,N_29699,N_29497);
nand UO_1785 (O_1785,N_29161,N_29492);
xor UO_1786 (O_1786,N_29774,N_29176);
xnor UO_1787 (O_1787,N_29327,N_28809);
xor UO_1788 (O_1788,N_29086,N_29800);
or UO_1789 (O_1789,N_29504,N_29003);
nand UO_1790 (O_1790,N_28890,N_29545);
xor UO_1791 (O_1791,N_29807,N_29673);
and UO_1792 (O_1792,N_28878,N_29701);
xor UO_1793 (O_1793,N_29246,N_29477);
and UO_1794 (O_1794,N_29964,N_28853);
xnor UO_1795 (O_1795,N_28917,N_29000);
nor UO_1796 (O_1796,N_29587,N_29864);
nor UO_1797 (O_1797,N_29727,N_28915);
or UO_1798 (O_1798,N_29521,N_29001);
nand UO_1799 (O_1799,N_29908,N_29877);
xnor UO_1800 (O_1800,N_29454,N_28917);
nor UO_1801 (O_1801,N_29528,N_28835);
nand UO_1802 (O_1802,N_29416,N_29272);
and UO_1803 (O_1803,N_29712,N_29407);
or UO_1804 (O_1804,N_29433,N_29557);
nand UO_1805 (O_1805,N_28975,N_28979);
xnor UO_1806 (O_1806,N_29122,N_29832);
nor UO_1807 (O_1807,N_29823,N_29028);
xnor UO_1808 (O_1808,N_29997,N_28920);
nor UO_1809 (O_1809,N_29142,N_29232);
and UO_1810 (O_1810,N_29725,N_29468);
xor UO_1811 (O_1811,N_29652,N_29529);
nor UO_1812 (O_1812,N_28993,N_28984);
and UO_1813 (O_1813,N_29054,N_28979);
or UO_1814 (O_1814,N_29538,N_29754);
nor UO_1815 (O_1815,N_29720,N_29774);
or UO_1816 (O_1816,N_29131,N_29559);
or UO_1817 (O_1817,N_29212,N_28966);
nor UO_1818 (O_1818,N_29334,N_29708);
or UO_1819 (O_1819,N_28812,N_29147);
and UO_1820 (O_1820,N_28972,N_29632);
xnor UO_1821 (O_1821,N_29404,N_29805);
nor UO_1822 (O_1822,N_29148,N_29900);
or UO_1823 (O_1823,N_29842,N_29853);
nand UO_1824 (O_1824,N_29362,N_29975);
and UO_1825 (O_1825,N_29838,N_29370);
or UO_1826 (O_1826,N_29786,N_29985);
nand UO_1827 (O_1827,N_29860,N_28941);
nor UO_1828 (O_1828,N_29277,N_29932);
nor UO_1829 (O_1829,N_29739,N_28983);
nand UO_1830 (O_1830,N_29858,N_29633);
nand UO_1831 (O_1831,N_29906,N_29885);
and UO_1832 (O_1832,N_29226,N_29702);
nor UO_1833 (O_1833,N_29692,N_28880);
or UO_1834 (O_1834,N_29426,N_29050);
nor UO_1835 (O_1835,N_28955,N_29870);
and UO_1836 (O_1836,N_29918,N_29488);
nand UO_1837 (O_1837,N_28826,N_29248);
or UO_1838 (O_1838,N_29578,N_29055);
nand UO_1839 (O_1839,N_29470,N_29294);
nor UO_1840 (O_1840,N_29513,N_29094);
and UO_1841 (O_1841,N_29135,N_29685);
nor UO_1842 (O_1842,N_29414,N_29886);
nor UO_1843 (O_1843,N_29209,N_28962);
nand UO_1844 (O_1844,N_29100,N_29401);
and UO_1845 (O_1845,N_29960,N_29574);
nand UO_1846 (O_1846,N_29830,N_29567);
and UO_1847 (O_1847,N_29574,N_28971);
and UO_1848 (O_1848,N_29548,N_29723);
xor UO_1849 (O_1849,N_29100,N_29371);
xor UO_1850 (O_1850,N_29441,N_29779);
nand UO_1851 (O_1851,N_29720,N_29524);
or UO_1852 (O_1852,N_29327,N_29880);
nor UO_1853 (O_1853,N_29076,N_29677);
nor UO_1854 (O_1854,N_28970,N_29555);
nor UO_1855 (O_1855,N_28846,N_29716);
nand UO_1856 (O_1856,N_29096,N_29814);
nor UO_1857 (O_1857,N_29684,N_29239);
or UO_1858 (O_1858,N_28950,N_29958);
and UO_1859 (O_1859,N_29614,N_28934);
nor UO_1860 (O_1860,N_29778,N_29903);
or UO_1861 (O_1861,N_29017,N_29097);
nand UO_1862 (O_1862,N_29197,N_29417);
xor UO_1863 (O_1863,N_29396,N_29911);
and UO_1864 (O_1864,N_29138,N_29133);
xnor UO_1865 (O_1865,N_29041,N_29701);
and UO_1866 (O_1866,N_29465,N_29068);
or UO_1867 (O_1867,N_29957,N_29803);
and UO_1868 (O_1868,N_29969,N_29284);
nor UO_1869 (O_1869,N_29522,N_28891);
and UO_1870 (O_1870,N_28955,N_28996);
and UO_1871 (O_1871,N_28858,N_29539);
nand UO_1872 (O_1872,N_29312,N_28806);
nand UO_1873 (O_1873,N_28906,N_29765);
xnor UO_1874 (O_1874,N_29652,N_29759);
nand UO_1875 (O_1875,N_28965,N_29986);
nor UO_1876 (O_1876,N_28923,N_29357);
or UO_1877 (O_1877,N_28961,N_28967);
nand UO_1878 (O_1878,N_29349,N_29495);
or UO_1879 (O_1879,N_29611,N_29289);
xnor UO_1880 (O_1880,N_29294,N_29319);
xor UO_1881 (O_1881,N_29830,N_29356);
or UO_1882 (O_1882,N_29111,N_29833);
and UO_1883 (O_1883,N_28850,N_28963);
nand UO_1884 (O_1884,N_29468,N_29967);
nand UO_1885 (O_1885,N_29699,N_29728);
or UO_1886 (O_1886,N_29214,N_29668);
or UO_1887 (O_1887,N_29618,N_29657);
and UO_1888 (O_1888,N_29286,N_29009);
or UO_1889 (O_1889,N_29870,N_29260);
and UO_1890 (O_1890,N_29157,N_29245);
and UO_1891 (O_1891,N_29425,N_29845);
xor UO_1892 (O_1892,N_29443,N_29618);
xnor UO_1893 (O_1893,N_29046,N_29228);
and UO_1894 (O_1894,N_29462,N_29303);
nor UO_1895 (O_1895,N_29023,N_29670);
nand UO_1896 (O_1896,N_29145,N_29044);
nand UO_1897 (O_1897,N_29734,N_28947);
nor UO_1898 (O_1898,N_29992,N_29505);
and UO_1899 (O_1899,N_29494,N_29449);
xnor UO_1900 (O_1900,N_29885,N_29238);
nand UO_1901 (O_1901,N_29504,N_29909);
and UO_1902 (O_1902,N_29561,N_29778);
or UO_1903 (O_1903,N_28913,N_29496);
nand UO_1904 (O_1904,N_29373,N_29517);
xor UO_1905 (O_1905,N_29712,N_29745);
nand UO_1906 (O_1906,N_29342,N_29208);
or UO_1907 (O_1907,N_29585,N_29178);
nor UO_1908 (O_1908,N_29550,N_29363);
or UO_1909 (O_1909,N_29986,N_29555);
xor UO_1910 (O_1910,N_29357,N_29310);
or UO_1911 (O_1911,N_28877,N_29224);
xnor UO_1912 (O_1912,N_29818,N_29283);
or UO_1913 (O_1913,N_29315,N_28822);
nor UO_1914 (O_1914,N_28833,N_29194);
or UO_1915 (O_1915,N_29113,N_29593);
and UO_1916 (O_1916,N_29879,N_29577);
nor UO_1917 (O_1917,N_29151,N_28810);
nand UO_1918 (O_1918,N_29763,N_28932);
or UO_1919 (O_1919,N_29131,N_29857);
and UO_1920 (O_1920,N_29661,N_29659);
and UO_1921 (O_1921,N_29852,N_29343);
nand UO_1922 (O_1922,N_28800,N_28845);
nand UO_1923 (O_1923,N_29604,N_29379);
or UO_1924 (O_1924,N_29667,N_29155);
or UO_1925 (O_1925,N_29941,N_29203);
xnor UO_1926 (O_1926,N_29371,N_29578);
and UO_1927 (O_1927,N_29723,N_29555);
nand UO_1928 (O_1928,N_28898,N_29053);
nor UO_1929 (O_1929,N_29727,N_29619);
nor UO_1930 (O_1930,N_29900,N_29150);
or UO_1931 (O_1931,N_29245,N_29455);
nor UO_1932 (O_1932,N_29746,N_29598);
nor UO_1933 (O_1933,N_29575,N_29596);
xor UO_1934 (O_1934,N_29027,N_29776);
and UO_1935 (O_1935,N_28946,N_29210);
nor UO_1936 (O_1936,N_28951,N_29301);
and UO_1937 (O_1937,N_29192,N_29058);
nand UO_1938 (O_1938,N_29707,N_29626);
nand UO_1939 (O_1939,N_28954,N_29668);
and UO_1940 (O_1940,N_28935,N_29493);
xnor UO_1941 (O_1941,N_29397,N_29753);
or UO_1942 (O_1942,N_29149,N_29792);
nor UO_1943 (O_1943,N_29464,N_29364);
xor UO_1944 (O_1944,N_28991,N_29738);
nor UO_1945 (O_1945,N_29858,N_29687);
xnor UO_1946 (O_1946,N_29947,N_29669);
nand UO_1947 (O_1947,N_29031,N_29759);
xor UO_1948 (O_1948,N_28901,N_29519);
nor UO_1949 (O_1949,N_29225,N_29515);
and UO_1950 (O_1950,N_29167,N_29657);
xor UO_1951 (O_1951,N_29083,N_29340);
nand UO_1952 (O_1952,N_28974,N_28836);
nor UO_1953 (O_1953,N_29941,N_29830);
nor UO_1954 (O_1954,N_29684,N_29048);
nor UO_1955 (O_1955,N_29715,N_28857);
and UO_1956 (O_1956,N_29031,N_29677);
and UO_1957 (O_1957,N_29521,N_29943);
or UO_1958 (O_1958,N_28968,N_29281);
nor UO_1959 (O_1959,N_29782,N_29560);
and UO_1960 (O_1960,N_29317,N_28908);
nand UO_1961 (O_1961,N_29972,N_29816);
nand UO_1962 (O_1962,N_29127,N_29760);
or UO_1963 (O_1963,N_28856,N_29999);
and UO_1964 (O_1964,N_29370,N_29361);
nand UO_1965 (O_1965,N_28859,N_29731);
nor UO_1966 (O_1966,N_29505,N_29078);
and UO_1967 (O_1967,N_28905,N_29063);
or UO_1968 (O_1968,N_29016,N_29651);
or UO_1969 (O_1969,N_29897,N_28933);
and UO_1970 (O_1970,N_29880,N_29397);
xor UO_1971 (O_1971,N_29712,N_29255);
nor UO_1972 (O_1972,N_29187,N_29433);
nand UO_1973 (O_1973,N_28998,N_29563);
xnor UO_1974 (O_1974,N_29476,N_29666);
nor UO_1975 (O_1975,N_29018,N_29187);
and UO_1976 (O_1976,N_29472,N_29955);
nor UO_1977 (O_1977,N_29056,N_29347);
and UO_1978 (O_1978,N_29048,N_29520);
xor UO_1979 (O_1979,N_29505,N_29030);
or UO_1980 (O_1980,N_29525,N_29296);
xnor UO_1981 (O_1981,N_29734,N_29254);
and UO_1982 (O_1982,N_29094,N_29399);
xor UO_1983 (O_1983,N_29907,N_28887);
xnor UO_1984 (O_1984,N_29078,N_29534);
or UO_1985 (O_1985,N_29278,N_29309);
nor UO_1986 (O_1986,N_29645,N_28961);
nand UO_1987 (O_1987,N_29943,N_29833);
or UO_1988 (O_1988,N_29953,N_29463);
and UO_1989 (O_1989,N_29858,N_29449);
nor UO_1990 (O_1990,N_29707,N_29050);
or UO_1991 (O_1991,N_29103,N_29905);
xor UO_1992 (O_1992,N_29973,N_28861);
and UO_1993 (O_1993,N_29742,N_29762);
xnor UO_1994 (O_1994,N_29387,N_29301);
nand UO_1995 (O_1995,N_29653,N_28958);
nand UO_1996 (O_1996,N_29305,N_29555);
nor UO_1997 (O_1997,N_28960,N_29126);
nand UO_1998 (O_1998,N_29697,N_29371);
and UO_1999 (O_1999,N_29259,N_28835);
and UO_2000 (O_2000,N_29618,N_29499);
or UO_2001 (O_2001,N_29053,N_29881);
or UO_2002 (O_2002,N_28853,N_29599);
or UO_2003 (O_2003,N_29052,N_29389);
nand UO_2004 (O_2004,N_28962,N_28894);
or UO_2005 (O_2005,N_29430,N_29710);
and UO_2006 (O_2006,N_29693,N_29217);
or UO_2007 (O_2007,N_29427,N_29215);
and UO_2008 (O_2008,N_29954,N_29403);
and UO_2009 (O_2009,N_29096,N_29157);
and UO_2010 (O_2010,N_28847,N_29715);
xor UO_2011 (O_2011,N_29949,N_29581);
nor UO_2012 (O_2012,N_28997,N_29683);
and UO_2013 (O_2013,N_29964,N_29942);
nand UO_2014 (O_2014,N_29220,N_29200);
nor UO_2015 (O_2015,N_29603,N_29201);
nor UO_2016 (O_2016,N_29380,N_29056);
or UO_2017 (O_2017,N_29548,N_29623);
nand UO_2018 (O_2018,N_29879,N_29124);
nand UO_2019 (O_2019,N_29955,N_28809);
and UO_2020 (O_2020,N_29865,N_29760);
or UO_2021 (O_2021,N_29651,N_29941);
and UO_2022 (O_2022,N_29000,N_29706);
xor UO_2023 (O_2023,N_29668,N_29742);
and UO_2024 (O_2024,N_28841,N_29256);
nor UO_2025 (O_2025,N_29460,N_28812);
nor UO_2026 (O_2026,N_29025,N_28978);
xor UO_2027 (O_2027,N_29445,N_28822);
nor UO_2028 (O_2028,N_29082,N_28996);
nand UO_2029 (O_2029,N_29768,N_29292);
nor UO_2030 (O_2030,N_29008,N_29130);
xor UO_2031 (O_2031,N_29391,N_29325);
nand UO_2032 (O_2032,N_29227,N_29456);
nand UO_2033 (O_2033,N_28862,N_29799);
xor UO_2034 (O_2034,N_29089,N_28955);
nor UO_2035 (O_2035,N_29858,N_28890);
or UO_2036 (O_2036,N_28851,N_29528);
nor UO_2037 (O_2037,N_29763,N_29035);
or UO_2038 (O_2038,N_29286,N_29685);
or UO_2039 (O_2039,N_29632,N_29678);
nor UO_2040 (O_2040,N_28844,N_28845);
nand UO_2041 (O_2041,N_29154,N_29563);
nor UO_2042 (O_2042,N_29856,N_29304);
nand UO_2043 (O_2043,N_29377,N_28976);
and UO_2044 (O_2044,N_28820,N_29394);
and UO_2045 (O_2045,N_29257,N_29129);
xor UO_2046 (O_2046,N_29536,N_29326);
or UO_2047 (O_2047,N_29454,N_28935);
nand UO_2048 (O_2048,N_29529,N_29387);
xnor UO_2049 (O_2049,N_29699,N_29344);
or UO_2050 (O_2050,N_29192,N_28936);
xnor UO_2051 (O_2051,N_29981,N_29067);
or UO_2052 (O_2052,N_29092,N_29010);
nand UO_2053 (O_2053,N_29418,N_29643);
nand UO_2054 (O_2054,N_28888,N_29894);
or UO_2055 (O_2055,N_29408,N_29833);
xnor UO_2056 (O_2056,N_28989,N_29528);
and UO_2057 (O_2057,N_29611,N_28908);
nor UO_2058 (O_2058,N_29213,N_29179);
xor UO_2059 (O_2059,N_29723,N_29863);
nor UO_2060 (O_2060,N_29902,N_29580);
and UO_2061 (O_2061,N_29942,N_29256);
and UO_2062 (O_2062,N_29386,N_28947);
nand UO_2063 (O_2063,N_29751,N_29892);
or UO_2064 (O_2064,N_29565,N_29486);
xnor UO_2065 (O_2065,N_29618,N_29392);
xnor UO_2066 (O_2066,N_29821,N_29582);
nand UO_2067 (O_2067,N_29688,N_28930);
xor UO_2068 (O_2068,N_29685,N_28833);
or UO_2069 (O_2069,N_29630,N_28932);
nor UO_2070 (O_2070,N_29465,N_29219);
or UO_2071 (O_2071,N_29617,N_29733);
nor UO_2072 (O_2072,N_29409,N_29437);
and UO_2073 (O_2073,N_29602,N_29863);
xnor UO_2074 (O_2074,N_29352,N_29387);
nor UO_2075 (O_2075,N_29783,N_29959);
xor UO_2076 (O_2076,N_29552,N_29256);
nor UO_2077 (O_2077,N_29443,N_29386);
nand UO_2078 (O_2078,N_29267,N_29556);
nand UO_2079 (O_2079,N_29151,N_29297);
nand UO_2080 (O_2080,N_29958,N_28899);
xnor UO_2081 (O_2081,N_29650,N_29050);
nor UO_2082 (O_2082,N_29177,N_29297);
nand UO_2083 (O_2083,N_29063,N_29322);
xor UO_2084 (O_2084,N_29602,N_29706);
nor UO_2085 (O_2085,N_29930,N_29370);
nand UO_2086 (O_2086,N_29261,N_29288);
and UO_2087 (O_2087,N_29028,N_29058);
xnor UO_2088 (O_2088,N_29032,N_28956);
nor UO_2089 (O_2089,N_28892,N_28828);
nor UO_2090 (O_2090,N_29143,N_29339);
xnor UO_2091 (O_2091,N_29245,N_28809);
or UO_2092 (O_2092,N_29535,N_28988);
xor UO_2093 (O_2093,N_28832,N_29749);
nand UO_2094 (O_2094,N_29693,N_29343);
nand UO_2095 (O_2095,N_29497,N_29044);
and UO_2096 (O_2096,N_29849,N_28967);
or UO_2097 (O_2097,N_29260,N_29416);
or UO_2098 (O_2098,N_29144,N_29938);
nand UO_2099 (O_2099,N_29270,N_29474);
xnor UO_2100 (O_2100,N_29516,N_29793);
nor UO_2101 (O_2101,N_29971,N_29670);
nor UO_2102 (O_2102,N_28964,N_29629);
and UO_2103 (O_2103,N_28852,N_29455);
nor UO_2104 (O_2104,N_29686,N_29860);
nand UO_2105 (O_2105,N_29020,N_29241);
xnor UO_2106 (O_2106,N_29732,N_28816);
and UO_2107 (O_2107,N_28819,N_29118);
nand UO_2108 (O_2108,N_29100,N_29231);
xnor UO_2109 (O_2109,N_29334,N_29891);
xnor UO_2110 (O_2110,N_28986,N_28882);
and UO_2111 (O_2111,N_29023,N_29728);
nor UO_2112 (O_2112,N_28870,N_29221);
nor UO_2113 (O_2113,N_29228,N_28808);
nand UO_2114 (O_2114,N_29915,N_28855);
or UO_2115 (O_2115,N_29874,N_29008);
and UO_2116 (O_2116,N_29738,N_29784);
xor UO_2117 (O_2117,N_29531,N_28820);
or UO_2118 (O_2118,N_29877,N_28911);
nor UO_2119 (O_2119,N_29873,N_29293);
nor UO_2120 (O_2120,N_29727,N_29327);
and UO_2121 (O_2121,N_29295,N_29460);
nand UO_2122 (O_2122,N_29166,N_29453);
nand UO_2123 (O_2123,N_29787,N_28918);
nand UO_2124 (O_2124,N_28846,N_28929);
or UO_2125 (O_2125,N_29907,N_29760);
nor UO_2126 (O_2126,N_29557,N_29525);
and UO_2127 (O_2127,N_29433,N_29537);
and UO_2128 (O_2128,N_29451,N_29927);
or UO_2129 (O_2129,N_29817,N_29704);
xor UO_2130 (O_2130,N_28886,N_28930);
or UO_2131 (O_2131,N_28931,N_29853);
xnor UO_2132 (O_2132,N_28825,N_29303);
xor UO_2133 (O_2133,N_29120,N_29988);
nand UO_2134 (O_2134,N_28814,N_28842);
xor UO_2135 (O_2135,N_29626,N_28824);
or UO_2136 (O_2136,N_28845,N_29671);
nor UO_2137 (O_2137,N_28906,N_29661);
nand UO_2138 (O_2138,N_29271,N_29202);
or UO_2139 (O_2139,N_29674,N_29686);
and UO_2140 (O_2140,N_29730,N_28956);
or UO_2141 (O_2141,N_29584,N_29010);
or UO_2142 (O_2142,N_28965,N_28930);
xnor UO_2143 (O_2143,N_29606,N_29850);
or UO_2144 (O_2144,N_29475,N_29647);
or UO_2145 (O_2145,N_28913,N_29625);
or UO_2146 (O_2146,N_29542,N_29843);
xnor UO_2147 (O_2147,N_29650,N_29167);
and UO_2148 (O_2148,N_29576,N_29085);
and UO_2149 (O_2149,N_29150,N_29110);
or UO_2150 (O_2150,N_29493,N_28970);
xor UO_2151 (O_2151,N_29081,N_29783);
and UO_2152 (O_2152,N_29942,N_28857);
and UO_2153 (O_2153,N_29753,N_29612);
nor UO_2154 (O_2154,N_29253,N_29568);
and UO_2155 (O_2155,N_29322,N_29560);
or UO_2156 (O_2156,N_29676,N_28910);
nand UO_2157 (O_2157,N_29184,N_28950);
or UO_2158 (O_2158,N_29641,N_28886);
and UO_2159 (O_2159,N_29534,N_29447);
nor UO_2160 (O_2160,N_29036,N_28940);
xnor UO_2161 (O_2161,N_29431,N_29095);
or UO_2162 (O_2162,N_29208,N_29798);
nand UO_2163 (O_2163,N_29173,N_29082);
nand UO_2164 (O_2164,N_29814,N_29968);
nand UO_2165 (O_2165,N_29942,N_29460);
or UO_2166 (O_2166,N_29380,N_28862);
or UO_2167 (O_2167,N_29505,N_29196);
and UO_2168 (O_2168,N_29191,N_28866);
or UO_2169 (O_2169,N_29865,N_29234);
or UO_2170 (O_2170,N_29985,N_29970);
nor UO_2171 (O_2171,N_29589,N_29873);
nand UO_2172 (O_2172,N_29213,N_29880);
or UO_2173 (O_2173,N_28957,N_29255);
xnor UO_2174 (O_2174,N_29413,N_29047);
xnor UO_2175 (O_2175,N_29201,N_29760);
nand UO_2176 (O_2176,N_28850,N_29508);
nand UO_2177 (O_2177,N_29426,N_29035);
or UO_2178 (O_2178,N_29077,N_29881);
or UO_2179 (O_2179,N_29930,N_29018);
nand UO_2180 (O_2180,N_29785,N_29733);
nand UO_2181 (O_2181,N_29677,N_29283);
nor UO_2182 (O_2182,N_28967,N_29963);
and UO_2183 (O_2183,N_29195,N_29381);
or UO_2184 (O_2184,N_29559,N_29330);
or UO_2185 (O_2185,N_28822,N_29483);
and UO_2186 (O_2186,N_29823,N_29291);
xnor UO_2187 (O_2187,N_29020,N_29221);
nand UO_2188 (O_2188,N_29160,N_28993);
nand UO_2189 (O_2189,N_28938,N_29805);
or UO_2190 (O_2190,N_29209,N_29424);
and UO_2191 (O_2191,N_29119,N_29855);
or UO_2192 (O_2192,N_29697,N_29750);
and UO_2193 (O_2193,N_29633,N_28969);
nor UO_2194 (O_2194,N_29837,N_29829);
and UO_2195 (O_2195,N_29337,N_29788);
and UO_2196 (O_2196,N_28914,N_29005);
nand UO_2197 (O_2197,N_29356,N_29740);
xnor UO_2198 (O_2198,N_29964,N_29896);
and UO_2199 (O_2199,N_29299,N_29869);
or UO_2200 (O_2200,N_29595,N_29805);
xnor UO_2201 (O_2201,N_28858,N_29573);
and UO_2202 (O_2202,N_29145,N_29306);
nor UO_2203 (O_2203,N_29268,N_29409);
nand UO_2204 (O_2204,N_29833,N_29261);
xnor UO_2205 (O_2205,N_29735,N_28893);
and UO_2206 (O_2206,N_29059,N_29891);
or UO_2207 (O_2207,N_29376,N_29135);
or UO_2208 (O_2208,N_29151,N_29402);
or UO_2209 (O_2209,N_29502,N_29856);
nor UO_2210 (O_2210,N_28971,N_29460);
and UO_2211 (O_2211,N_29330,N_29456);
or UO_2212 (O_2212,N_28853,N_28813);
or UO_2213 (O_2213,N_29276,N_29789);
and UO_2214 (O_2214,N_28910,N_29577);
nor UO_2215 (O_2215,N_29680,N_29849);
nand UO_2216 (O_2216,N_28892,N_29790);
or UO_2217 (O_2217,N_29384,N_29156);
and UO_2218 (O_2218,N_29894,N_28821);
and UO_2219 (O_2219,N_29237,N_29519);
nand UO_2220 (O_2220,N_29659,N_29607);
xor UO_2221 (O_2221,N_29234,N_29156);
nor UO_2222 (O_2222,N_29318,N_29806);
nor UO_2223 (O_2223,N_28814,N_29348);
or UO_2224 (O_2224,N_29196,N_29281);
nor UO_2225 (O_2225,N_29489,N_29168);
nor UO_2226 (O_2226,N_29251,N_28983);
xor UO_2227 (O_2227,N_29756,N_29862);
or UO_2228 (O_2228,N_29376,N_29546);
and UO_2229 (O_2229,N_29788,N_28959);
or UO_2230 (O_2230,N_29095,N_29781);
nand UO_2231 (O_2231,N_29853,N_28810);
or UO_2232 (O_2232,N_29154,N_28853);
or UO_2233 (O_2233,N_29707,N_29794);
and UO_2234 (O_2234,N_29893,N_29116);
nor UO_2235 (O_2235,N_29301,N_29413);
and UO_2236 (O_2236,N_29626,N_28980);
and UO_2237 (O_2237,N_29984,N_29606);
and UO_2238 (O_2238,N_29114,N_29672);
xnor UO_2239 (O_2239,N_29741,N_29101);
and UO_2240 (O_2240,N_29541,N_28831);
and UO_2241 (O_2241,N_29127,N_29853);
and UO_2242 (O_2242,N_28868,N_29197);
nand UO_2243 (O_2243,N_28842,N_29661);
or UO_2244 (O_2244,N_28908,N_29064);
or UO_2245 (O_2245,N_29881,N_29554);
or UO_2246 (O_2246,N_28993,N_29125);
or UO_2247 (O_2247,N_29512,N_29664);
xnor UO_2248 (O_2248,N_29141,N_29226);
and UO_2249 (O_2249,N_29802,N_29943);
nor UO_2250 (O_2250,N_29357,N_28967);
nor UO_2251 (O_2251,N_29425,N_29878);
and UO_2252 (O_2252,N_29987,N_28884);
and UO_2253 (O_2253,N_29909,N_29452);
or UO_2254 (O_2254,N_28963,N_29773);
and UO_2255 (O_2255,N_29503,N_29953);
nor UO_2256 (O_2256,N_29577,N_28948);
nand UO_2257 (O_2257,N_29535,N_29065);
or UO_2258 (O_2258,N_29761,N_29488);
xor UO_2259 (O_2259,N_29711,N_29330);
or UO_2260 (O_2260,N_29818,N_29741);
or UO_2261 (O_2261,N_29544,N_29356);
nand UO_2262 (O_2262,N_29984,N_28851);
xnor UO_2263 (O_2263,N_28861,N_29237);
xnor UO_2264 (O_2264,N_29540,N_29585);
xor UO_2265 (O_2265,N_29542,N_29512);
or UO_2266 (O_2266,N_29399,N_28827);
nor UO_2267 (O_2267,N_29189,N_28900);
nor UO_2268 (O_2268,N_29814,N_29761);
nor UO_2269 (O_2269,N_29758,N_29790);
and UO_2270 (O_2270,N_29429,N_28894);
and UO_2271 (O_2271,N_29604,N_29264);
nand UO_2272 (O_2272,N_29127,N_29505);
nor UO_2273 (O_2273,N_29350,N_28839);
nand UO_2274 (O_2274,N_29744,N_29301);
nand UO_2275 (O_2275,N_29700,N_29340);
nand UO_2276 (O_2276,N_28902,N_29308);
xnor UO_2277 (O_2277,N_29263,N_28835);
xnor UO_2278 (O_2278,N_29199,N_29241);
and UO_2279 (O_2279,N_29667,N_29072);
xnor UO_2280 (O_2280,N_29675,N_29493);
xor UO_2281 (O_2281,N_29990,N_29530);
nor UO_2282 (O_2282,N_29694,N_28919);
xnor UO_2283 (O_2283,N_28952,N_29865);
or UO_2284 (O_2284,N_29026,N_29494);
nor UO_2285 (O_2285,N_29946,N_29032);
and UO_2286 (O_2286,N_29563,N_29921);
nor UO_2287 (O_2287,N_29480,N_29789);
nor UO_2288 (O_2288,N_29854,N_29648);
xnor UO_2289 (O_2289,N_29056,N_29272);
or UO_2290 (O_2290,N_29495,N_29581);
nor UO_2291 (O_2291,N_28960,N_28964);
xnor UO_2292 (O_2292,N_29527,N_29949);
xor UO_2293 (O_2293,N_29280,N_29655);
nor UO_2294 (O_2294,N_29809,N_29504);
xor UO_2295 (O_2295,N_29803,N_29050);
nand UO_2296 (O_2296,N_29022,N_28967);
or UO_2297 (O_2297,N_28804,N_29702);
nand UO_2298 (O_2298,N_29901,N_29681);
nor UO_2299 (O_2299,N_29147,N_29002);
xnor UO_2300 (O_2300,N_29620,N_28904);
nand UO_2301 (O_2301,N_29058,N_28894);
nand UO_2302 (O_2302,N_29730,N_29541);
or UO_2303 (O_2303,N_29449,N_29709);
nand UO_2304 (O_2304,N_29153,N_29473);
nor UO_2305 (O_2305,N_29641,N_29193);
and UO_2306 (O_2306,N_29598,N_29194);
xnor UO_2307 (O_2307,N_29312,N_29702);
and UO_2308 (O_2308,N_28957,N_28972);
nand UO_2309 (O_2309,N_29590,N_29444);
nand UO_2310 (O_2310,N_28961,N_29148);
nor UO_2311 (O_2311,N_29666,N_29413);
nor UO_2312 (O_2312,N_29570,N_29527);
xnor UO_2313 (O_2313,N_28856,N_29750);
or UO_2314 (O_2314,N_29881,N_28896);
xor UO_2315 (O_2315,N_29608,N_29684);
and UO_2316 (O_2316,N_29470,N_29996);
nor UO_2317 (O_2317,N_29450,N_29198);
xnor UO_2318 (O_2318,N_29427,N_29101);
xor UO_2319 (O_2319,N_29955,N_29338);
or UO_2320 (O_2320,N_28899,N_29105);
nand UO_2321 (O_2321,N_29520,N_29004);
nor UO_2322 (O_2322,N_29626,N_29541);
nor UO_2323 (O_2323,N_29716,N_29703);
nor UO_2324 (O_2324,N_29456,N_29716);
nand UO_2325 (O_2325,N_29300,N_29270);
nand UO_2326 (O_2326,N_29869,N_29822);
nand UO_2327 (O_2327,N_29266,N_29478);
or UO_2328 (O_2328,N_29163,N_29831);
nor UO_2329 (O_2329,N_29487,N_29620);
and UO_2330 (O_2330,N_29561,N_29443);
or UO_2331 (O_2331,N_29209,N_29723);
or UO_2332 (O_2332,N_29281,N_28935);
nor UO_2333 (O_2333,N_29110,N_29583);
nand UO_2334 (O_2334,N_29604,N_29657);
and UO_2335 (O_2335,N_29677,N_29681);
and UO_2336 (O_2336,N_29227,N_29185);
nand UO_2337 (O_2337,N_29950,N_29112);
nor UO_2338 (O_2338,N_29355,N_29901);
nor UO_2339 (O_2339,N_29253,N_29921);
and UO_2340 (O_2340,N_29873,N_28932);
xor UO_2341 (O_2341,N_29923,N_29976);
or UO_2342 (O_2342,N_29553,N_29132);
xor UO_2343 (O_2343,N_28802,N_29842);
or UO_2344 (O_2344,N_29117,N_28912);
or UO_2345 (O_2345,N_29010,N_29119);
nand UO_2346 (O_2346,N_28826,N_29379);
nor UO_2347 (O_2347,N_29504,N_29823);
nand UO_2348 (O_2348,N_29449,N_29889);
or UO_2349 (O_2349,N_29321,N_29482);
and UO_2350 (O_2350,N_29934,N_29767);
nor UO_2351 (O_2351,N_29826,N_28888);
or UO_2352 (O_2352,N_29166,N_29067);
or UO_2353 (O_2353,N_29220,N_29293);
and UO_2354 (O_2354,N_29505,N_28815);
or UO_2355 (O_2355,N_29480,N_29177);
nor UO_2356 (O_2356,N_29794,N_29295);
xnor UO_2357 (O_2357,N_29087,N_29193);
nand UO_2358 (O_2358,N_29614,N_29408);
nand UO_2359 (O_2359,N_29219,N_28849);
nand UO_2360 (O_2360,N_29244,N_29892);
xnor UO_2361 (O_2361,N_29693,N_29909);
nor UO_2362 (O_2362,N_28885,N_29887);
and UO_2363 (O_2363,N_29489,N_28934);
nor UO_2364 (O_2364,N_29712,N_29050);
and UO_2365 (O_2365,N_29236,N_28841);
and UO_2366 (O_2366,N_29881,N_28876);
or UO_2367 (O_2367,N_29363,N_29406);
nand UO_2368 (O_2368,N_29159,N_29631);
nand UO_2369 (O_2369,N_29582,N_29112);
nand UO_2370 (O_2370,N_29180,N_29938);
nor UO_2371 (O_2371,N_29770,N_28814);
nand UO_2372 (O_2372,N_29628,N_29971);
and UO_2373 (O_2373,N_29178,N_29841);
nand UO_2374 (O_2374,N_28849,N_29516);
or UO_2375 (O_2375,N_29444,N_29568);
xnor UO_2376 (O_2376,N_29185,N_29210);
or UO_2377 (O_2377,N_29736,N_29450);
or UO_2378 (O_2378,N_29585,N_29712);
nor UO_2379 (O_2379,N_29453,N_29062);
and UO_2380 (O_2380,N_29449,N_29365);
or UO_2381 (O_2381,N_29614,N_29558);
or UO_2382 (O_2382,N_29877,N_29777);
nor UO_2383 (O_2383,N_29755,N_29994);
xor UO_2384 (O_2384,N_29734,N_29476);
xnor UO_2385 (O_2385,N_29673,N_29903);
nor UO_2386 (O_2386,N_29403,N_29731);
nand UO_2387 (O_2387,N_28909,N_29076);
xnor UO_2388 (O_2388,N_29787,N_28929);
nor UO_2389 (O_2389,N_29114,N_29041);
nor UO_2390 (O_2390,N_28935,N_29906);
xnor UO_2391 (O_2391,N_29322,N_29598);
nand UO_2392 (O_2392,N_29108,N_28926);
or UO_2393 (O_2393,N_28969,N_29115);
nor UO_2394 (O_2394,N_28980,N_29235);
nor UO_2395 (O_2395,N_28978,N_29321);
nand UO_2396 (O_2396,N_28991,N_29893);
and UO_2397 (O_2397,N_29749,N_29660);
xor UO_2398 (O_2398,N_28893,N_29005);
or UO_2399 (O_2399,N_29443,N_29913);
nand UO_2400 (O_2400,N_29540,N_29438);
and UO_2401 (O_2401,N_29849,N_28972);
xor UO_2402 (O_2402,N_29014,N_29615);
and UO_2403 (O_2403,N_29508,N_29464);
xnor UO_2404 (O_2404,N_29777,N_29056);
or UO_2405 (O_2405,N_28882,N_28812);
xnor UO_2406 (O_2406,N_29718,N_29743);
and UO_2407 (O_2407,N_28941,N_29394);
or UO_2408 (O_2408,N_28973,N_29665);
and UO_2409 (O_2409,N_29654,N_29781);
xor UO_2410 (O_2410,N_29916,N_28925);
or UO_2411 (O_2411,N_29252,N_29859);
xor UO_2412 (O_2412,N_29623,N_28975);
xnor UO_2413 (O_2413,N_29588,N_29847);
nand UO_2414 (O_2414,N_29794,N_29321);
or UO_2415 (O_2415,N_28962,N_29632);
nor UO_2416 (O_2416,N_29446,N_29622);
xor UO_2417 (O_2417,N_29175,N_29575);
and UO_2418 (O_2418,N_29172,N_29876);
and UO_2419 (O_2419,N_29518,N_28874);
and UO_2420 (O_2420,N_29849,N_29381);
nand UO_2421 (O_2421,N_29730,N_28847);
nor UO_2422 (O_2422,N_29499,N_29428);
nand UO_2423 (O_2423,N_29585,N_29656);
nand UO_2424 (O_2424,N_29204,N_29464);
xor UO_2425 (O_2425,N_29484,N_29755);
nand UO_2426 (O_2426,N_28991,N_29673);
nand UO_2427 (O_2427,N_29498,N_29170);
and UO_2428 (O_2428,N_29268,N_28966);
nand UO_2429 (O_2429,N_29170,N_29243);
xnor UO_2430 (O_2430,N_29249,N_29664);
and UO_2431 (O_2431,N_28834,N_29175);
and UO_2432 (O_2432,N_29535,N_29254);
and UO_2433 (O_2433,N_29403,N_29485);
xnor UO_2434 (O_2434,N_29324,N_29893);
xor UO_2435 (O_2435,N_29214,N_29102);
nand UO_2436 (O_2436,N_29886,N_29502);
and UO_2437 (O_2437,N_29887,N_29446);
xor UO_2438 (O_2438,N_29645,N_29915);
and UO_2439 (O_2439,N_29536,N_29557);
or UO_2440 (O_2440,N_29967,N_29881);
nand UO_2441 (O_2441,N_29772,N_29799);
nand UO_2442 (O_2442,N_29520,N_28837);
nor UO_2443 (O_2443,N_29475,N_29330);
or UO_2444 (O_2444,N_29390,N_28868);
and UO_2445 (O_2445,N_28911,N_29367);
nand UO_2446 (O_2446,N_29917,N_29709);
nor UO_2447 (O_2447,N_28869,N_28859);
xnor UO_2448 (O_2448,N_29647,N_29454);
nand UO_2449 (O_2449,N_29965,N_29724);
or UO_2450 (O_2450,N_29281,N_29682);
or UO_2451 (O_2451,N_29242,N_29850);
xnor UO_2452 (O_2452,N_29427,N_29840);
nor UO_2453 (O_2453,N_29546,N_29033);
or UO_2454 (O_2454,N_29904,N_29343);
nand UO_2455 (O_2455,N_29477,N_29784);
nor UO_2456 (O_2456,N_28921,N_29496);
xnor UO_2457 (O_2457,N_29670,N_29787);
or UO_2458 (O_2458,N_29108,N_29169);
or UO_2459 (O_2459,N_28991,N_28987);
xnor UO_2460 (O_2460,N_28961,N_29904);
nor UO_2461 (O_2461,N_29216,N_28823);
nand UO_2462 (O_2462,N_29972,N_29699);
nand UO_2463 (O_2463,N_29749,N_29511);
xnor UO_2464 (O_2464,N_29616,N_29686);
or UO_2465 (O_2465,N_28915,N_29827);
nand UO_2466 (O_2466,N_29858,N_29855);
or UO_2467 (O_2467,N_28971,N_29733);
or UO_2468 (O_2468,N_29382,N_29580);
and UO_2469 (O_2469,N_29307,N_28829);
nor UO_2470 (O_2470,N_28855,N_29524);
nand UO_2471 (O_2471,N_29368,N_29649);
nand UO_2472 (O_2472,N_29468,N_29801);
and UO_2473 (O_2473,N_29595,N_28849);
and UO_2474 (O_2474,N_29012,N_29985);
nor UO_2475 (O_2475,N_29618,N_29468);
and UO_2476 (O_2476,N_29177,N_29970);
nand UO_2477 (O_2477,N_29565,N_29172);
nand UO_2478 (O_2478,N_29292,N_29145);
nor UO_2479 (O_2479,N_29852,N_29611);
and UO_2480 (O_2480,N_29696,N_29060);
and UO_2481 (O_2481,N_29356,N_29344);
or UO_2482 (O_2482,N_29928,N_28934);
nand UO_2483 (O_2483,N_29380,N_29587);
nand UO_2484 (O_2484,N_28905,N_29538);
xor UO_2485 (O_2485,N_29789,N_29013);
or UO_2486 (O_2486,N_29061,N_28807);
or UO_2487 (O_2487,N_29551,N_29226);
and UO_2488 (O_2488,N_29898,N_29727);
nor UO_2489 (O_2489,N_29310,N_29490);
nand UO_2490 (O_2490,N_29410,N_29237);
xnor UO_2491 (O_2491,N_29497,N_29933);
nand UO_2492 (O_2492,N_29122,N_29038);
nor UO_2493 (O_2493,N_29472,N_29741);
nand UO_2494 (O_2494,N_29765,N_29681);
nor UO_2495 (O_2495,N_29496,N_29768);
or UO_2496 (O_2496,N_29910,N_29353);
xor UO_2497 (O_2497,N_28990,N_29317);
nand UO_2498 (O_2498,N_29382,N_29425);
and UO_2499 (O_2499,N_29076,N_29092);
nand UO_2500 (O_2500,N_29209,N_29689);
nor UO_2501 (O_2501,N_29695,N_29989);
and UO_2502 (O_2502,N_29160,N_29653);
nor UO_2503 (O_2503,N_29698,N_28967);
xor UO_2504 (O_2504,N_29136,N_29883);
and UO_2505 (O_2505,N_29291,N_29922);
nand UO_2506 (O_2506,N_29572,N_28885);
xor UO_2507 (O_2507,N_29071,N_29039);
nor UO_2508 (O_2508,N_29829,N_29998);
nor UO_2509 (O_2509,N_29965,N_29656);
or UO_2510 (O_2510,N_29827,N_29953);
nand UO_2511 (O_2511,N_29754,N_29433);
nor UO_2512 (O_2512,N_29280,N_29250);
xor UO_2513 (O_2513,N_29298,N_29986);
or UO_2514 (O_2514,N_29130,N_28991);
and UO_2515 (O_2515,N_29058,N_29519);
or UO_2516 (O_2516,N_29437,N_29874);
xor UO_2517 (O_2517,N_29544,N_29001);
or UO_2518 (O_2518,N_29903,N_29206);
and UO_2519 (O_2519,N_29702,N_29965);
xnor UO_2520 (O_2520,N_29116,N_29802);
and UO_2521 (O_2521,N_29704,N_28905);
or UO_2522 (O_2522,N_29678,N_29026);
or UO_2523 (O_2523,N_29244,N_29982);
nand UO_2524 (O_2524,N_29555,N_29088);
nor UO_2525 (O_2525,N_29907,N_28925);
and UO_2526 (O_2526,N_29605,N_28873);
or UO_2527 (O_2527,N_29116,N_29868);
nand UO_2528 (O_2528,N_28982,N_29813);
nor UO_2529 (O_2529,N_28948,N_29021);
and UO_2530 (O_2530,N_29669,N_29278);
nor UO_2531 (O_2531,N_29917,N_29727);
xor UO_2532 (O_2532,N_29388,N_29060);
xnor UO_2533 (O_2533,N_29149,N_29576);
and UO_2534 (O_2534,N_29751,N_29901);
nor UO_2535 (O_2535,N_29312,N_29961);
or UO_2536 (O_2536,N_28979,N_28955);
and UO_2537 (O_2537,N_28951,N_29944);
xnor UO_2538 (O_2538,N_29823,N_29230);
nand UO_2539 (O_2539,N_29390,N_29290);
nor UO_2540 (O_2540,N_28848,N_29985);
and UO_2541 (O_2541,N_29710,N_29518);
and UO_2542 (O_2542,N_29730,N_29445);
xor UO_2543 (O_2543,N_29449,N_28861);
and UO_2544 (O_2544,N_29182,N_29277);
xnor UO_2545 (O_2545,N_28850,N_29147);
or UO_2546 (O_2546,N_29107,N_29134);
nor UO_2547 (O_2547,N_29707,N_29264);
nand UO_2548 (O_2548,N_29705,N_29992);
or UO_2549 (O_2549,N_29800,N_29187);
and UO_2550 (O_2550,N_29560,N_29617);
nand UO_2551 (O_2551,N_29715,N_29187);
and UO_2552 (O_2552,N_29103,N_29799);
xnor UO_2553 (O_2553,N_29208,N_28845);
xnor UO_2554 (O_2554,N_29729,N_29579);
nand UO_2555 (O_2555,N_29793,N_28914);
nand UO_2556 (O_2556,N_29361,N_29039);
and UO_2557 (O_2557,N_29378,N_29523);
xnor UO_2558 (O_2558,N_29564,N_29429);
nor UO_2559 (O_2559,N_29117,N_28998);
nor UO_2560 (O_2560,N_29873,N_29165);
and UO_2561 (O_2561,N_29057,N_28970);
and UO_2562 (O_2562,N_29639,N_29363);
xor UO_2563 (O_2563,N_29123,N_28866);
and UO_2564 (O_2564,N_29865,N_29410);
and UO_2565 (O_2565,N_29710,N_29387);
nand UO_2566 (O_2566,N_29526,N_29065);
or UO_2567 (O_2567,N_29956,N_29940);
or UO_2568 (O_2568,N_28823,N_29421);
nand UO_2569 (O_2569,N_29761,N_29022);
and UO_2570 (O_2570,N_29913,N_28876);
and UO_2571 (O_2571,N_29088,N_29132);
nand UO_2572 (O_2572,N_29310,N_29245);
xor UO_2573 (O_2573,N_29019,N_29055);
xnor UO_2574 (O_2574,N_29744,N_29715);
nor UO_2575 (O_2575,N_29435,N_29196);
xnor UO_2576 (O_2576,N_29665,N_29759);
and UO_2577 (O_2577,N_28911,N_29558);
xnor UO_2578 (O_2578,N_29488,N_29683);
and UO_2579 (O_2579,N_29761,N_29306);
nand UO_2580 (O_2580,N_29327,N_29119);
nand UO_2581 (O_2581,N_29532,N_29053);
or UO_2582 (O_2582,N_29319,N_29137);
xnor UO_2583 (O_2583,N_29015,N_28982);
and UO_2584 (O_2584,N_28894,N_29904);
or UO_2585 (O_2585,N_29116,N_29688);
and UO_2586 (O_2586,N_29108,N_28803);
and UO_2587 (O_2587,N_29677,N_29447);
or UO_2588 (O_2588,N_29710,N_29982);
nor UO_2589 (O_2589,N_29266,N_29706);
and UO_2590 (O_2590,N_29687,N_29400);
or UO_2591 (O_2591,N_29321,N_29277);
and UO_2592 (O_2592,N_29014,N_29071);
nand UO_2593 (O_2593,N_29566,N_29930);
and UO_2594 (O_2594,N_29226,N_29680);
nand UO_2595 (O_2595,N_29904,N_29278);
and UO_2596 (O_2596,N_29978,N_29184);
and UO_2597 (O_2597,N_29175,N_29012);
and UO_2598 (O_2598,N_29873,N_28976);
and UO_2599 (O_2599,N_29493,N_29109);
nor UO_2600 (O_2600,N_29153,N_29746);
xor UO_2601 (O_2601,N_29956,N_28912);
nor UO_2602 (O_2602,N_29984,N_29262);
nor UO_2603 (O_2603,N_29579,N_29997);
nor UO_2604 (O_2604,N_29282,N_29537);
or UO_2605 (O_2605,N_29390,N_29924);
or UO_2606 (O_2606,N_29013,N_29780);
and UO_2607 (O_2607,N_29180,N_28996);
nor UO_2608 (O_2608,N_29563,N_29104);
nor UO_2609 (O_2609,N_29597,N_29807);
or UO_2610 (O_2610,N_29105,N_29274);
xnor UO_2611 (O_2611,N_29239,N_28912);
nand UO_2612 (O_2612,N_29450,N_28979);
and UO_2613 (O_2613,N_29482,N_28944);
and UO_2614 (O_2614,N_28823,N_29334);
nor UO_2615 (O_2615,N_29613,N_29100);
nor UO_2616 (O_2616,N_28830,N_29668);
xnor UO_2617 (O_2617,N_29818,N_29415);
xor UO_2618 (O_2618,N_29480,N_29939);
nand UO_2619 (O_2619,N_29616,N_29567);
nor UO_2620 (O_2620,N_29876,N_28978);
nand UO_2621 (O_2621,N_29157,N_28943);
xor UO_2622 (O_2622,N_29785,N_28942);
and UO_2623 (O_2623,N_28988,N_29665);
and UO_2624 (O_2624,N_29926,N_29918);
and UO_2625 (O_2625,N_29678,N_29874);
or UO_2626 (O_2626,N_28938,N_28904);
and UO_2627 (O_2627,N_29795,N_29293);
and UO_2628 (O_2628,N_29180,N_29852);
xor UO_2629 (O_2629,N_29334,N_29740);
nor UO_2630 (O_2630,N_29337,N_29163);
nand UO_2631 (O_2631,N_29545,N_29656);
nor UO_2632 (O_2632,N_28802,N_29456);
and UO_2633 (O_2633,N_29448,N_29230);
nand UO_2634 (O_2634,N_28802,N_28971);
nand UO_2635 (O_2635,N_29499,N_29890);
or UO_2636 (O_2636,N_29497,N_29948);
xnor UO_2637 (O_2637,N_29195,N_29522);
nand UO_2638 (O_2638,N_29389,N_28864);
xnor UO_2639 (O_2639,N_29127,N_29272);
or UO_2640 (O_2640,N_29510,N_29392);
or UO_2641 (O_2641,N_29231,N_29923);
nor UO_2642 (O_2642,N_29742,N_29390);
nand UO_2643 (O_2643,N_29480,N_29661);
xor UO_2644 (O_2644,N_29314,N_29558);
nor UO_2645 (O_2645,N_29765,N_29285);
nor UO_2646 (O_2646,N_29564,N_29466);
xor UO_2647 (O_2647,N_29947,N_28913);
nand UO_2648 (O_2648,N_29656,N_29007);
and UO_2649 (O_2649,N_29782,N_29050);
nand UO_2650 (O_2650,N_29939,N_29196);
xnor UO_2651 (O_2651,N_29282,N_29325);
nand UO_2652 (O_2652,N_29478,N_29045);
or UO_2653 (O_2653,N_29775,N_29564);
xnor UO_2654 (O_2654,N_29675,N_29831);
xor UO_2655 (O_2655,N_29804,N_29158);
or UO_2656 (O_2656,N_29888,N_29801);
and UO_2657 (O_2657,N_29920,N_29478);
nand UO_2658 (O_2658,N_29281,N_29097);
or UO_2659 (O_2659,N_28821,N_29819);
xor UO_2660 (O_2660,N_29806,N_29488);
nand UO_2661 (O_2661,N_29411,N_28855);
xor UO_2662 (O_2662,N_29761,N_29948);
or UO_2663 (O_2663,N_29352,N_29242);
and UO_2664 (O_2664,N_28952,N_29986);
and UO_2665 (O_2665,N_28814,N_29703);
nor UO_2666 (O_2666,N_29957,N_29461);
and UO_2667 (O_2667,N_29741,N_29634);
or UO_2668 (O_2668,N_29979,N_29938);
nand UO_2669 (O_2669,N_29210,N_29654);
or UO_2670 (O_2670,N_29567,N_29788);
and UO_2671 (O_2671,N_29012,N_29363);
nand UO_2672 (O_2672,N_28917,N_29716);
xor UO_2673 (O_2673,N_29801,N_29578);
nor UO_2674 (O_2674,N_29956,N_29027);
nand UO_2675 (O_2675,N_29105,N_29754);
nand UO_2676 (O_2676,N_29833,N_29978);
xor UO_2677 (O_2677,N_29030,N_29127);
nand UO_2678 (O_2678,N_29353,N_29170);
and UO_2679 (O_2679,N_29589,N_28953);
xor UO_2680 (O_2680,N_29563,N_29923);
and UO_2681 (O_2681,N_29291,N_28958);
xnor UO_2682 (O_2682,N_29114,N_29716);
and UO_2683 (O_2683,N_29885,N_29428);
nand UO_2684 (O_2684,N_29581,N_29922);
or UO_2685 (O_2685,N_29469,N_29808);
xor UO_2686 (O_2686,N_29330,N_29211);
xnor UO_2687 (O_2687,N_29499,N_29663);
nand UO_2688 (O_2688,N_29657,N_29189);
xor UO_2689 (O_2689,N_29701,N_29299);
and UO_2690 (O_2690,N_29555,N_29000);
xnor UO_2691 (O_2691,N_28846,N_29059);
or UO_2692 (O_2692,N_29659,N_29016);
nand UO_2693 (O_2693,N_29259,N_29561);
and UO_2694 (O_2694,N_29640,N_29941);
and UO_2695 (O_2695,N_29298,N_29882);
or UO_2696 (O_2696,N_28980,N_29655);
nand UO_2697 (O_2697,N_29061,N_29930);
nor UO_2698 (O_2698,N_29595,N_29366);
nor UO_2699 (O_2699,N_29841,N_29922);
and UO_2700 (O_2700,N_29743,N_29435);
xnor UO_2701 (O_2701,N_28878,N_29039);
nand UO_2702 (O_2702,N_29247,N_29745);
nor UO_2703 (O_2703,N_29443,N_29521);
xnor UO_2704 (O_2704,N_29312,N_29307);
or UO_2705 (O_2705,N_29542,N_29736);
xnor UO_2706 (O_2706,N_29249,N_29425);
nor UO_2707 (O_2707,N_29311,N_29636);
nand UO_2708 (O_2708,N_28865,N_28983);
xor UO_2709 (O_2709,N_28853,N_29296);
nor UO_2710 (O_2710,N_29416,N_29599);
nor UO_2711 (O_2711,N_29129,N_29323);
nor UO_2712 (O_2712,N_29087,N_29559);
and UO_2713 (O_2713,N_29229,N_29173);
xor UO_2714 (O_2714,N_28883,N_29481);
xnor UO_2715 (O_2715,N_29930,N_29746);
and UO_2716 (O_2716,N_29704,N_29306);
xor UO_2717 (O_2717,N_29570,N_29718);
nand UO_2718 (O_2718,N_29634,N_29814);
nor UO_2719 (O_2719,N_29782,N_29965);
xnor UO_2720 (O_2720,N_29194,N_29533);
and UO_2721 (O_2721,N_29808,N_29682);
and UO_2722 (O_2722,N_28927,N_29569);
xor UO_2723 (O_2723,N_29625,N_29710);
or UO_2724 (O_2724,N_29644,N_29383);
nor UO_2725 (O_2725,N_29686,N_29167);
and UO_2726 (O_2726,N_29341,N_29266);
or UO_2727 (O_2727,N_29644,N_29123);
or UO_2728 (O_2728,N_29262,N_29142);
xor UO_2729 (O_2729,N_28802,N_29303);
and UO_2730 (O_2730,N_29019,N_29722);
and UO_2731 (O_2731,N_28959,N_29117);
or UO_2732 (O_2732,N_28833,N_29101);
and UO_2733 (O_2733,N_29824,N_29220);
or UO_2734 (O_2734,N_29686,N_29779);
nand UO_2735 (O_2735,N_29608,N_28827);
nand UO_2736 (O_2736,N_29387,N_29015);
or UO_2737 (O_2737,N_29015,N_29929);
or UO_2738 (O_2738,N_29663,N_29418);
or UO_2739 (O_2739,N_29885,N_29954);
nor UO_2740 (O_2740,N_29245,N_29499);
or UO_2741 (O_2741,N_29628,N_29860);
nor UO_2742 (O_2742,N_29671,N_29051);
nor UO_2743 (O_2743,N_29538,N_28823);
nand UO_2744 (O_2744,N_29574,N_29889);
and UO_2745 (O_2745,N_28997,N_29372);
or UO_2746 (O_2746,N_29263,N_29270);
and UO_2747 (O_2747,N_29706,N_29679);
nand UO_2748 (O_2748,N_29317,N_29797);
and UO_2749 (O_2749,N_29315,N_29378);
xor UO_2750 (O_2750,N_29828,N_29756);
xor UO_2751 (O_2751,N_29846,N_28904);
xor UO_2752 (O_2752,N_29158,N_29221);
nand UO_2753 (O_2753,N_29467,N_29181);
nor UO_2754 (O_2754,N_29082,N_29300);
or UO_2755 (O_2755,N_29137,N_29468);
xor UO_2756 (O_2756,N_29313,N_29683);
and UO_2757 (O_2757,N_29894,N_29113);
and UO_2758 (O_2758,N_28806,N_29807);
and UO_2759 (O_2759,N_29246,N_29538);
and UO_2760 (O_2760,N_29371,N_29906);
nand UO_2761 (O_2761,N_29098,N_29150);
nand UO_2762 (O_2762,N_28892,N_28815);
nand UO_2763 (O_2763,N_29992,N_29805);
xor UO_2764 (O_2764,N_29166,N_29248);
nand UO_2765 (O_2765,N_29183,N_29387);
and UO_2766 (O_2766,N_29830,N_28811);
nand UO_2767 (O_2767,N_29158,N_28943);
nor UO_2768 (O_2768,N_29818,N_28823);
and UO_2769 (O_2769,N_29797,N_29068);
xor UO_2770 (O_2770,N_28942,N_29580);
xor UO_2771 (O_2771,N_29159,N_29170);
nand UO_2772 (O_2772,N_29000,N_29762);
xnor UO_2773 (O_2773,N_29251,N_28953);
nor UO_2774 (O_2774,N_29384,N_29544);
nor UO_2775 (O_2775,N_29353,N_28854);
xnor UO_2776 (O_2776,N_28943,N_29801);
xnor UO_2777 (O_2777,N_29746,N_29631);
and UO_2778 (O_2778,N_29866,N_29949);
or UO_2779 (O_2779,N_29658,N_29215);
and UO_2780 (O_2780,N_29111,N_29669);
xnor UO_2781 (O_2781,N_29022,N_29464);
and UO_2782 (O_2782,N_28983,N_29751);
nor UO_2783 (O_2783,N_29735,N_29821);
nand UO_2784 (O_2784,N_29968,N_29048);
xnor UO_2785 (O_2785,N_29209,N_29618);
or UO_2786 (O_2786,N_29505,N_28975);
nand UO_2787 (O_2787,N_29304,N_29433);
and UO_2788 (O_2788,N_29861,N_29121);
and UO_2789 (O_2789,N_29568,N_29006);
nand UO_2790 (O_2790,N_29913,N_28998);
or UO_2791 (O_2791,N_29936,N_29262);
xnor UO_2792 (O_2792,N_29249,N_28966);
nor UO_2793 (O_2793,N_29047,N_29625);
or UO_2794 (O_2794,N_29517,N_29836);
nor UO_2795 (O_2795,N_29769,N_28847);
xnor UO_2796 (O_2796,N_29332,N_28995);
xor UO_2797 (O_2797,N_28889,N_28955);
xnor UO_2798 (O_2798,N_29518,N_29017);
nor UO_2799 (O_2799,N_29833,N_29856);
nand UO_2800 (O_2800,N_29635,N_29941);
xor UO_2801 (O_2801,N_29001,N_29012);
xnor UO_2802 (O_2802,N_29744,N_29510);
nand UO_2803 (O_2803,N_29179,N_29745);
and UO_2804 (O_2804,N_28852,N_29618);
or UO_2805 (O_2805,N_29933,N_29794);
nand UO_2806 (O_2806,N_29335,N_28832);
or UO_2807 (O_2807,N_28803,N_29233);
xnor UO_2808 (O_2808,N_29567,N_28894);
and UO_2809 (O_2809,N_29250,N_29464);
or UO_2810 (O_2810,N_29217,N_29144);
xnor UO_2811 (O_2811,N_29750,N_29250);
or UO_2812 (O_2812,N_29959,N_29253);
nor UO_2813 (O_2813,N_29387,N_29552);
and UO_2814 (O_2814,N_29693,N_28861);
and UO_2815 (O_2815,N_29235,N_28870);
or UO_2816 (O_2816,N_29047,N_29680);
or UO_2817 (O_2817,N_29096,N_29628);
xnor UO_2818 (O_2818,N_29501,N_29031);
or UO_2819 (O_2819,N_29099,N_29309);
and UO_2820 (O_2820,N_29927,N_29752);
nor UO_2821 (O_2821,N_28846,N_29659);
or UO_2822 (O_2822,N_29165,N_29439);
nor UO_2823 (O_2823,N_28872,N_29590);
nor UO_2824 (O_2824,N_29342,N_29024);
nand UO_2825 (O_2825,N_29079,N_29314);
and UO_2826 (O_2826,N_29022,N_29128);
and UO_2827 (O_2827,N_29618,N_29217);
or UO_2828 (O_2828,N_29640,N_29251);
or UO_2829 (O_2829,N_29147,N_29192);
or UO_2830 (O_2830,N_28806,N_29535);
or UO_2831 (O_2831,N_29124,N_29901);
nand UO_2832 (O_2832,N_29704,N_29644);
xor UO_2833 (O_2833,N_29318,N_29168);
xor UO_2834 (O_2834,N_28832,N_28808);
and UO_2835 (O_2835,N_29600,N_29390);
or UO_2836 (O_2836,N_28832,N_29574);
xor UO_2837 (O_2837,N_29677,N_29739);
xnor UO_2838 (O_2838,N_29527,N_29880);
xnor UO_2839 (O_2839,N_29078,N_29491);
or UO_2840 (O_2840,N_29819,N_29808);
nor UO_2841 (O_2841,N_29212,N_28802);
and UO_2842 (O_2842,N_29672,N_29188);
and UO_2843 (O_2843,N_29882,N_29431);
xnor UO_2844 (O_2844,N_29445,N_28932);
xnor UO_2845 (O_2845,N_28847,N_29216);
xnor UO_2846 (O_2846,N_28829,N_28826);
or UO_2847 (O_2847,N_29755,N_28938);
nor UO_2848 (O_2848,N_28954,N_29808);
nor UO_2849 (O_2849,N_29827,N_29443);
or UO_2850 (O_2850,N_29645,N_29238);
nand UO_2851 (O_2851,N_29930,N_29568);
or UO_2852 (O_2852,N_29547,N_29660);
xnor UO_2853 (O_2853,N_28840,N_28888);
xor UO_2854 (O_2854,N_28875,N_29924);
nand UO_2855 (O_2855,N_29105,N_28932);
or UO_2856 (O_2856,N_29631,N_29519);
or UO_2857 (O_2857,N_29220,N_29907);
nand UO_2858 (O_2858,N_29803,N_28907);
and UO_2859 (O_2859,N_29039,N_29310);
nor UO_2860 (O_2860,N_29658,N_29722);
or UO_2861 (O_2861,N_29471,N_29156);
or UO_2862 (O_2862,N_29334,N_29259);
and UO_2863 (O_2863,N_28994,N_29349);
xor UO_2864 (O_2864,N_29370,N_29932);
nor UO_2865 (O_2865,N_28834,N_29756);
nand UO_2866 (O_2866,N_29119,N_29120);
nand UO_2867 (O_2867,N_29778,N_28888);
nor UO_2868 (O_2868,N_29957,N_28836);
nor UO_2869 (O_2869,N_29796,N_29261);
nand UO_2870 (O_2870,N_28896,N_29841);
and UO_2871 (O_2871,N_29630,N_28897);
and UO_2872 (O_2872,N_29271,N_29106);
nor UO_2873 (O_2873,N_29023,N_29809);
nand UO_2874 (O_2874,N_29142,N_29187);
nand UO_2875 (O_2875,N_29197,N_29106);
and UO_2876 (O_2876,N_29323,N_28924);
nand UO_2877 (O_2877,N_29267,N_29654);
nand UO_2878 (O_2878,N_28856,N_29694);
nand UO_2879 (O_2879,N_29369,N_29435);
xor UO_2880 (O_2880,N_28809,N_29486);
or UO_2881 (O_2881,N_28911,N_29825);
xor UO_2882 (O_2882,N_29218,N_29555);
and UO_2883 (O_2883,N_28962,N_29407);
nand UO_2884 (O_2884,N_29279,N_29144);
xnor UO_2885 (O_2885,N_29818,N_29925);
nand UO_2886 (O_2886,N_28898,N_29867);
or UO_2887 (O_2887,N_29526,N_28835);
xnor UO_2888 (O_2888,N_28820,N_29172);
xor UO_2889 (O_2889,N_29606,N_29375);
nand UO_2890 (O_2890,N_29093,N_29564);
xnor UO_2891 (O_2891,N_29002,N_29227);
xnor UO_2892 (O_2892,N_28908,N_29493);
xnor UO_2893 (O_2893,N_29035,N_29452);
nand UO_2894 (O_2894,N_29386,N_29664);
xnor UO_2895 (O_2895,N_28869,N_29107);
nand UO_2896 (O_2896,N_28851,N_29193);
nor UO_2897 (O_2897,N_29510,N_29807);
or UO_2898 (O_2898,N_29697,N_29136);
and UO_2899 (O_2899,N_29155,N_29598);
or UO_2900 (O_2900,N_28951,N_29588);
nand UO_2901 (O_2901,N_29766,N_28840);
nor UO_2902 (O_2902,N_29525,N_29490);
and UO_2903 (O_2903,N_29517,N_29230);
and UO_2904 (O_2904,N_29747,N_29064);
or UO_2905 (O_2905,N_29780,N_29602);
nand UO_2906 (O_2906,N_29774,N_29483);
or UO_2907 (O_2907,N_29307,N_29971);
xnor UO_2908 (O_2908,N_29003,N_29068);
or UO_2909 (O_2909,N_28801,N_29277);
or UO_2910 (O_2910,N_29655,N_29295);
nor UO_2911 (O_2911,N_29706,N_29155);
and UO_2912 (O_2912,N_29196,N_29115);
xor UO_2913 (O_2913,N_28961,N_29725);
and UO_2914 (O_2914,N_29059,N_29226);
or UO_2915 (O_2915,N_29060,N_29027);
and UO_2916 (O_2916,N_29593,N_29780);
nand UO_2917 (O_2917,N_29022,N_28920);
and UO_2918 (O_2918,N_28894,N_29354);
nand UO_2919 (O_2919,N_29275,N_29119);
nand UO_2920 (O_2920,N_28884,N_29083);
xnor UO_2921 (O_2921,N_29512,N_29181);
nand UO_2922 (O_2922,N_29741,N_29896);
nor UO_2923 (O_2923,N_29046,N_29317);
or UO_2924 (O_2924,N_28831,N_28818);
xnor UO_2925 (O_2925,N_29005,N_29169);
and UO_2926 (O_2926,N_29282,N_28837);
and UO_2927 (O_2927,N_29692,N_29430);
and UO_2928 (O_2928,N_28951,N_28825);
nand UO_2929 (O_2929,N_29912,N_29546);
and UO_2930 (O_2930,N_29761,N_28947);
xor UO_2931 (O_2931,N_29814,N_29866);
nand UO_2932 (O_2932,N_29756,N_29609);
nor UO_2933 (O_2933,N_29533,N_29430);
nor UO_2934 (O_2934,N_29632,N_29122);
nor UO_2935 (O_2935,N_29577,N_29249);
and UO_2936 (O_2936,N_29168,N_29141);
nor UO_2937 (O_2937,N_29367,N_28979);
or UO_2938 (O_2938,N_28887,N_29310);
or UO_2939 (O_2939,N_29345,N_29788);
nand UO_2940 (O_2940,N_29700,N_29222);
nand UO_2941 (O_2941,N_29317,N_29744);
nor UO_2942 (O_2942,N_29861,N_29669);
xnor UO_2943 (O_2943,N_29540,N_29407);
or UO_2944 (O_2944,N_29360,N_29513);
xnor UO_2945 (O_2945,N_29190,N_28929);
nand UO_2946 (O_2946,N_29731,N_29490);
nand UO_2947 (O_2947,N_29719,N_29030);
and UO_2948 (O_2948,N_29333,N_29958);
nand UO_2949 (O_2949,N_29886,N_29255);
xnor UO_2950 (O_2950,N_29962,N_29213);
nand UO_2951 (O_2951,N_29837,N_29069);
or UO_2952 (O_2952,N_29834,N_28860);
nor UO_2953 (O_2953,N_29935,N_29585);
xor UO_2954 (O_2954,N_29673,N_29563);
nor UO_2955 (O_2955,N_29843,N_29393);
xor UO_2956 (O_2956,N_28834,N_29507);
or UO_2957 (O_2957,N_29402,N_29314);
and UO_2958 (O_2958,N_29041,N_29156);
xnor UO_2959 (O_2959,N_29244,N_29092);
or UO_2960 (O_2960,N_29173,N_29991);
nor UO_2961 (O_2961,N_29377,N_28803);
or UO_2962 (O_2962,N_29390,N_29492);
nor UO_2963 (O_2963,N_29353,N_29073);
or UO_2964 (O_2964,N_29153,N_29480);
or UO_2965 (O_2965,N_29243,N_29499);
nand UO_2966 (O_2966,N_29741,N_29631);
nor UO_2967 (O_2967,N_28946,N_28981);
xor UO_2968 (O_2968,N_29620,N_29989);
xor UO_2969 (O_2969,N_29595,N_29858);
and UO_2970 (O_2970,N_28993,N_29121);
nor UO_2971 (O_2971,N_29496,N_29630);
nand UO_2972 (O_2972,N_29459,N_29104);
nor UO_2973 (O_2973,N_28961,N_29854);
nand UO_2974 (O_2974,N_28907,N_29749);
and UO_2975 (O_2975,N_29547,N_29104);
and UO_2976 (O_2976,N_29741,N_29423);
or UO_2977 (O_2977,N_29393,N_29863);
nor UO_2978 (O_2978,N_29162,N_29253);
nor UO_2979 (O_2979,N_29549,N_29101);
nand UO_2980 (O_2980,N_29773,N_29815);
and UO_2981 (O_2981,N_29415,N_29931);
or UO_2982 (O_2982,N_28904,N_29908);
or UO_2983 (O_2983,N_29715,N_29934);
nand UO_2984 (O_2984,N_29931,N_29099);
xnor UO_2985 (O_2985,N_29843,N_29738);
and UO_2986 (O_2986,N_29913,N_29522);
and UO_2987 (O_2987,N_28964,N_28999);
nor UO_2988 (O_2988,N_28816,N_29632);
nand UO_2989 (O_2989,N_29046,N_28914);
and UO_2990 (O_2990,N_29871,N_29953);
and UO_2991 (O_2991,N_29910,N_29249);
xnor UO_2992 (O_2992,N_29486,N_28911);
nand UO_2993 (O_2993,N_29538,N_29639);
xor UO_2994 (O_2994,N_29825,N_29914);
and UO_2995 (O_2995,N_29889,N_29722);
nand UO_2996 (O_2996,N_29931,N_29784);
and UO_2997 (O_2997,N_29630,N_29060);
or UO_2998 (O_2998,N_29114,N_28967);
or UO_2999 (O_2999,N_29994,N_29715);
nand UO_3000 (O_3000,N_29850,N_29875);
or UO_3001 (O_3001,N_29905,N_29474);
and UO_3002 (O_3002,N_29505,N_29220);
nand UO_3003 (O_3003,N_29864,N_29173);
xor UO_3004 (O_3004,N_29745,N_29431);
xor UO_3005 (O_3005,N_29118,N_29244);
nor UO_3006 (O_3006,N_28929,N_29927);
nor UO_3007 (O_3007,N_29113,N_29147);
nand UO_3008 (O_3008,N_29001,N_29918);
nor UO_3009 (O_3009,N_29629,N_29054);
xor UO_3010 (O_3010,N_29440,N_28815);
or UO_3011 (O_3011,N_28881,N_28959);
xor UO_3012 (O_3012,N_28807,N_29766);
or UO_3013 (O_3013,N_29388,N_29633);
or UO_3014 (O_3014,N_29052,N_29333);
and UO_3015 (O_3015,N_29090,N_29425);
or UO_3016 (O_3016,N_29207,N_29640);
nor UO_3017 (O_3017,N_29018,N_29692);
or UO_3018 (O_3018,N_29643,N_28969);
xnor UO_3019 (O_3019,N_29172,N_29402);
and UO_3020 (O_3020,N_29982,N_29271);
or UO_3021 (O_3021,N_29041,N_29225);
and UO_3022 (O_3022,N_29248,N_29446);
or UO_3023 (O_3023,N_29883,N_29207);
or UO_3024 (O_3024,N_29678,N_29872);
or UO_3025 (O_3025,N_29431,N_29993);
nor UO_3026 (O_3026,N_28815,N_29468);
and UO_3027 (O_3027,N_28950,N_28928);
nand UO_3028 (O_3028,N_29554,N_29423);
nand UO_3029 (O_3029,N_29510,N_29219);
xor UO_3030 (O_3030,N_29992,N_29889);
and UO_3031 (O_3031,N_29308,N_29356);
xnor UO_3032 (O_3032,N_29140,N_29065);
xor UO_3033 (O_3033,N_29206,N_29956);
nor UO_3034 (O_3034,N_29368,N_29821);
nand UO_3035 (O_3035,N_29638,N_29104);
and UO_3036 (O_3036,N_29264,N_29377);
nand UO_3037 (O_3037,N_29290,N_29214);
or UO_3038 (O_3038,N_29912,N_29823);
nand UO_3039 (O_3039,N_29149,N_29811);
and UO_3040 (O_3040,N_29826,N_29016);
xor UO_3041 (O_3041,N_29293,N_29868);
nand UO_3042 (O_3042,N_29907,N_29977);
nand UO_3043 (O_3043,N_28930,N_29333);
or UO_3044 (O_3044,N_29210,N_29749);
xnor UO_3045 (O_3045,N_29153,N_29509);
or UO_3046 (O_3046,N_29633,N_29329);
or UO_3047 (O_3047,N_29577,N_29221);
or UO_3048 (O_3048,N_28918,N_29329);
nand UO_3049 (O_3049,N_28957,N_29121);
or UO_3050 (O_3050,N_29649,N_29324);
and UO_3051 (O_3051,N_29268,N_28858);
xor UO_3052 (O_3052,N_28924,N_29261);
xor UO_3053 (O_3053,N_29706,N_29976);
and UO_3054 (O_3054,N_29958,N_29030);
nor UO_3055 (O_3055,N_29681,N_28845);
and UO_3056 (O_3056,N_29948,N_29004);
xnor UO_3057 (O_3057,N_29151,N_29262);
xor UO_3058 (O_3058,N_29146,N_29800);
xor UO_3059 (O_3059,N_29461,N_29047);
nand UO_3060 (O_3060,N_29998,N_29424);
nor UO_3061 (O_3061,N_29348,N_29459);
or UO_3062 (O_3062,N_29211,N_29088);
xor UO_3063 (O_3063,N_29951,N_28848);
nor UO_3064 (O_3064,N_29264,N_29478);
nand UO_3065 (O_3065,N_29844,N_29167);
nor UO_3066 (O_3066,N_29582,N_28877);
nand UO_3067 (O_3067,N_29642,N_29016);
and UO_3068 (O_3068,N_28925,N_29897);
nor UO_3069 (O_3069,N_28817,N_29694);
xnor UO_3070 (O_3070,N_29883,N_29014);
nand UO_3071 (O_3071,N_29216,N_29391);
or UO_3072 (O_3072,N_29371,N_29820);
or UO_3073 (O_3073,N_29910,N_29089);
nand UO_3074 (O_3074,N_29632,N_29328);
or UO_3075 (O_3075,N_29029,N_29631);
nand UO_3076 (O_3076,N_29906,N_29835);
xnor UO_3077 (O_3077,N_28838,N_29665);
nor UO_3078 (O_3078,N_29877,N_28901);
or UO_3079 (O_3079,N_29054,N_29199);
and UO_3080 (O_3080,N_29233,N_29072);
or UO_3081 (O_3081,N_29400,N_28957);
nand UO_3082 (O_3082,N_29975,N_29836);
nand UO_3083 (O_3083,N_28957,N_29791);
nand UO_3084 (O_3084,N_29325,N_29554);
or UO_3085 (O_3085,N_28882,N_28818);
nand UO_3086 (O_3086,N_29992,N_29497);
nor UO_3087 (O_3087,N_29908,N_29074);
xnor UO_3088 (O_3088,N_28987,N_29872);
nor UO_3089 (O_3089,N_29970,N_29820);
xnor UO_3090 (O_3090,N_29296,N_29007);
nand UO_3091 (O_3091,N_29452,N_29513);
or UO_3092 (O_3092,N_29289,N_29697);
nor UO_3093 (O_3093,N_29939,N_29391);
xnor UO_3094 (O_3094,N_28902,N_29757);
nand UO_3095 (O_3095,N_29822,N_29785);
and UO_3096 (O_3096,N_29351,N_29518);
xnor UO_3097 (O_3097,N_29123,N_29753);
nand UO_3098 (O_3098,N_29286,N_29797);
nor UO_3099 (O_3099,N_29415,N_29845);
nand UO_3100 (O_3100,N_28850,N_28851);
or UO_3101 (O_3101,N_28964,N_29766);
nor UO_3102 (O_3102,N_29234,N_29070);
nor UO_3103 (O_3103,N_29651,N_29150);
and UO_3104 (O_3104,N_29179,N_28866);
or UO_3105 (O_3105,N_29342,N_29177);
nand UO_3106 (O_3106,N_29802,N_29028);
or UO_3107 (O_3107,N_29871,N_29005);
and UO_3108 (O_3108,N_29076,N_29297);
xor UO_3109 (O_3109,N_28901,N_28969);
or UO_3110 (O_3110,N_29248,N_29981);
xor UO_3111 (O_3111,N_29367,N_29078);
or UO_3112 (O_3112,N_28904,N_29956);
or UO_3113 (O_3113,N_29167,N_29013);
xnor UO_3114 (O_3114,N_29336,N_28973);
nand UO_3115 (O_3115,N_29524,N_29112);
nor UO_3116 (O_3116,N_28817,N_29776);
nor UO_3117 (O_3117,N_29082,N_29418);
nand UO_3118 (O_3118,N_29967,N_29169);
or UO_3119 (O_3119,N_29342,N_29445);
xnor UO_3120 (O_3120,N_28882,N_29629);
nand UO_3121 (O_3121,N_29733,N_29984);
and UO_3122 (O_3122,N_29164,N_29756);
or UO_3123 (O_3123,N_29392,N_29290);
xor UO_3124 (O_3124,N_29942,N_28957);
nor UO_3125 (O_3125,N_29794,N_29437);
xor UO_3126 (O_3126,N_29308,N_29015);
and UO_3127 (O_3127,N_29758,N_29915);
or UO_3128 (O_3128,N_29506,N_29798);
or UO_3129 (O_3129,N_29913,N_29313);
nand UO_3130 (O_3130,N_29756,N_29197);
xor UO_3131 (O_3131,N_29192,N_29649);
nand UO_3132 (O_3132,N_28889,N_28858);
nand UO_3133 (O_3133,N_29546,N_29366);
and UO_3134 (O_3134,N_29070,N_29730);
xor UO_3135 (O_3135,N_29569,N_29881);
xor UO_3136 (O_3136,N_29375,N_29814);
nand UO_3137 (O_3137,N_29299,N_29010);
and UO_3138 (O_3138,N_29308,N_29609);
or UO_3139 (O_3139,N_29466,N_29727);
xnor UO_3140 (O_3140,N_29166,N_29742);
nand UO_3141 (O_3141,N_29637,N_28999);
nand UO_3142 (O_3142,N_29613,N_29183);
and UO_3143 (O_3143,N_29502,N_29201);
nor UO_3144 (O_3144,N_29858,N_29262);
and UO_3145 (O_3145,N_29040,N_29634);
and UO_3146 (O_3146,N_29086,N_29712);
and UO_3147 (O_3147,N_29210,N_29423);
nand UO_3148 (O_3148,N_29332,N_29128);
and UO_3149 (O_3149,N_29737,N_28933);
xor UO_3150 (O_3150,N_28859,N_29592);
or UO_3151 (O_3151,N_29054,N_29293);
and UO_3152 (O_3152,N_29566,N_29734);
nand UO_3153 (O_3153,N_29870,N_29528);
nand UO_3154 (O_3154,N_28960,N_29900);
nor UO_3155 (O_3155,N_29080,N_29581);
or UO_3156 (O_3156,N_29708,N_29964);
or UO_3157 (O_3157,N_29330,N_29239);
nor UO_3158 (O_3158,N_29313,N_28881);
or UO_3159 (O_3159,N_29092,N_29388);
or UO_3160 (O_3160,N_29728,N_29031);
and UO_3161 (O_3161,N_29325,N_29899);
or UO_3162 (O_3162,N_29268,N_29235);
nand UO_3163 (O_3163,N_28948,N_28827);
or UO_3164 (O_3164,N_29343,N_29283);
nand UO_3165 (O_3165,N_29204,N_29236);
and UO_3166 (O_3166,N_28880,N_29607);
xor UO_3167 (O_3167,N_29267,N_29017);
nor UO_3168 (O_3168,N_29323,N_29389);
and UO_3169 (O_3169,N_29645,N_29715);
nand UO_3170 (O_3170,N_29595,N_29572);
nor UO_3171 (O_3171,N_29046,N_28853);
or UO_3172 (O_3172,N_29527,N_29183);
nor UO_3173 (O_3173,N_29511,N_28938);
nor UO_3174 (O_3174,N_29147,N_28878);
xnor UO_3175 (O_3175,N_29400,N_29234);
or UO_3176 (O_3176,N_28897,N_28876);
nor UO_3177 (O_3177,N_29179,N_29706);
nor UO_3178 (O_3178,N_29124,N_29028);
nor UO_3179 (O_3179,N_29908,N_28939);
nor UO_3180 (O_3180,N_29423,N_29342);
nand UO_3181 (O_3181,N_29256,N_29081);
nor UO_3182 (O_3182,N_29632,N_28987);
and UO_3183 (O_3183,N_29176,N_28851);
or UO_3184 (O_3184,N_29710,N_28958);
xnor UO_3185 (O_3185,N_29860,N_28999);
nor UO_3186 (O_3186,N_29483,N_29917);
or UO_3187 (O_3187,N_29304,N_29263);
and UO_3188 (O_3188,N_29671,N_29742);
nor UO_3189 (O_3189,N_29701,N_29231);
xor UO_3190 (O_3190,N_28971,N_29269);
and UO_3191 (O_3191,N_29111,N_29620);
nand UO_3192 (O_3192,N_29585,N_29489);
nand UO_3193 (O_3193,N_29436,N_29880);
xnor UO_3194 (O_3194,N_28994,N_29746);
or UO_3195 (O_3195,N_28889,N_29835);
nor UO_3196 (O_3196,N_29572,N_29141);
nor UO_3197 (O_3197,N_28915,N_28812);
and UO_3198 (O_3198,N_29633,N_29326);
xor UO_3199 (O_3199,N_29248,N_29000);
nor UO_3200 (O_3200,N_29208,N_29205);
or UO_3201 (O_3201,N_29802,N_29079);
and UO_3202 (O_3202,N_29942,N_28916);
or UO_3203 (O_3203,N_29897,N_29068);
xnor UO_3204 (O_3204,N_29354,N_29454);
and UO_3205 (O_3205,N_29389,N_29034);
nor UO_3206 (O_3206,N_29447,N_29422);
nand UO_3207 (O_3207,N_29222,N_29946);
or UO_3208 (O_3208,N_29454,N_29235);
or UO_3209 (O_3209,N_29730,N_29212);
and UO_3210 (O_3210,N_29021,N_28849);
xor UO_3211 (O_3211,N_29764,N_28862);
nor UO_3212 (O_3212,N_29075,N_29051);
nand UO_3213 (O_3213,N_29255,N_29958);
nand UO_3214 (O_3214,N_29218,N_29681);
or UO_3215 (O_3215,N_29532,N_29126);
or UO_3216 (O_3216,N_28999,N_29060);
nand UO_3217 (O_3217,N_28890,N_29381);
nand UO_3218 (O_3218,N_29009,N_29921);
nor UO_3219 (O_3219,N_29878,N_29603);
nand UO_3220 (O_3220,N_29660,N_28814);
nor UO_3221 (O_3221,N_29491,N_29436);
xnor UO_3222 (O_3222,N_29910,N_29937);
xnor UO_3223 (O_3223,N_29726,N_29463);
nand UO_3224 (O_3224,N_28940,N_29747);
xor UO_3225 (O_3225,N_29587,N_29708);
or UO_3226 (O_3226,N_29794,N_28995);
nand UO_3227 (O_3227,N_29015,N_28887);
and UO_3228 (O_3228,N_29713,N_29585);
and UO_3229 (O_3229,N_29501,N_29431);
nor UO_3230 (O_3230,N_29605,N_29462);
or UO_3231 (O_3231,N_29530,N_29447);
xnor UO_3232 (O_3232,N_29834,N_29379);
and UO_3233 (O_3233,N_29184,N_29233);
and UO_3234 (O_3234,N_29693,N_28812);
and UO_3235 (O_3235,N_29535,N_29332);
xnor UO_3236 (O_3236,N_29777,N_28933);
and UO_3237 (O_3237,N_28991,N_29334);
nor UO_3238 (O_3238,N_29659,N_28801);
and UO_3239 (O_3239,N_29665,N_29074);
or UO_3240 (O_3240,N_29432,N_29506);
and UO_3241 (O_3241,N_29990,N_29149);
nand UO_3242 (O_3242,N_29585,N_28883);
or UO_3243 (O_3243,N_28941,N_29889);
and UO_3244 (O_3244,N_28834,N_29222);
nor UO_3245 (O_3245,N_29169,N_29232);
xnor UO_3246 (O_3246,N_29965,N_29375);
xnor UO_3247 (O_3247,N_29290,N_29818);
nor UO_3248 (O_3248,N_29488,N_29089);
nor UO_3249 (O_3249,N_29147,N_29712);
or UO_3250 (O_3250,N_29592,N_29472);
nor UO_3251 (O_3251,N_28850,N_28872);
nand UO_3252 (O_3252,N_29758,N_29413);
and UO_3253 (O_3253,N_29890,N_29223);
xnor UO_3254 (O_3254,N_29299,N_29067);
nand UO_3255 (O_3255,N_29984,N_29981);
and UO_3256 (O_3256,N_29852,N_29443);
nand UO_3257 (O_3257,N_29061,N_29745);
xor UO_3258 (O_3258,N_28871,N_29111);
or UO_3259 (O_3259,N_29122,N_29610);
nand UO_3260 (O_3260,N_29594,N_29756);
nand UO_3261 (O_3261,N_28866,N_29104);
nor UO_3262 (O_3262,N_29795,N_29386);
xnor UO_3263 (O_3263,N_29387,N_29296);
xnor UO_3264 (O_3264,N_29820,N_29445);
nand UO_3265 (O_3265,N_29602,N_29376);
and UO_3266 (O_3266,N_28909,N_29247);
or UO_3267 (O_3267,N_29964,N_28819);
nand UO_3268 (O_3268,N_29242,N_28951);
nor UO_3269 (O_3269,N_29119,N_29453);
or UO_3270 (O_3270,N_29607,N_29430);
and UO_3271 (O_3271,N_29340,N_29857);
nand UO_3272 (O_3272,N_29446,N_28946);
xnor UO_3273 (O_3273,N_28995,N_29368);
nor UO_3274 (O_3274,N_29934,N_29303);
nor UO_3275 (O_3275,N_29200,N_29507);
or UO_3276 (O_3276,N_29074,N_29408);
and UO_3277 (O_3277,N_28871,N_29449);
and UO_3278 (O_3278,N_29238,N_29837);
xor UO_3279 (O_3279,N_29440,N_29413);
xor UO_3280 (O_3280,N_29030,N_28822);
nand UO_3281 (O_3281,N_29735,N_29690);
or UO_3282 (O_3282,N_29736,N_28975);
nor UO_3283 (O_3283,N_29854,N_29243);
and UO_3284 (O_3284,N_29273,N_29051);
or UO_3285 (O_3285,N_29720,N_29759);
nand UO_3286 (O_3286,N_29160,N_29115);
and UO_3287 (O_3287,N_29642,N_28892);
nor UO_3288 (O_3288,N_28930,N_29096);
nor UO_3289 (O_3289,N_29236,N_29852);
xor UO_3290 (O_3290,N_28948,N_29961);
and UO_3291 (O_3291,N_29799,N_29725);
or UO_3292 (O_3292,N_28945,N_29576);
nand UO_3293 (O_3293,N_29002,N_29153);
nand UO_3294 (O_3294,N_29501,N_29211);
or UO_3295 (O_3295,N_28950,N_29459);
or UO_3296 (O_3296,N_29901,N_28903);
and UO_3297 (O_3297,N_29555,N_28819);
or UO_3298 (O_3298,N_29009,N_29892);
nor UO_3299 (O_3299,N_29759,N_29188);
nor UO_3300 (O_3300,N_29323,N_29939);
nor UO_3301 (O_3301,N_29422,N_29875);
xnor UO_3302 (O_3302,N_29713,N_28970);
or UO_3303 (O_3303,N_29210,N_29183);
or UO_3304 (O_3304,N_28863,N_29594);
xor UO_3305 (O_3305,N_29797,N_29124);
nor UO_3306 (O_3306,N_29064,N_29439);
nand UO_3307 (O_3307,N_28876,N_29655);
xnor UO_3308 (O_3308,N_29543,N_29297);
or UO_3309 (O_3309,N_29005,N_29316);
and UO_3310 (O_3310,N_29521,N_29364);
xnor UO_3311 (O_3311,N_29357,N_29486);
nor UO_3312 (O_3312,N_28901,N_29094);
nor UO_3313 (O_3313,N_29392,N_28934);
and UO_3314 (O_3314,N_29430,N_29259);
or UO_3315 (O_3315,N_29553,N_29276);
and UO_3316 (O_3316,N_28967,N_29878);
and UO_3317 (O_3317,N_29746,N_28985);
xnor UO_3318 (O_3318,N_29639,N_29648);
nand UO_3319 (O_3319,N_29487,N_29893);
xor UO_3320 (O_3320,N_29673,N_29780);
nor UO_3321 (O_3321,N_29494,N_28963);
nor UO_3322 (O_3322,N_28919,N_29510);
nand UO_3323 (O_3323,N_29056,N_29116);
xor UO_3324 (O_3324,N_28808,N_29387);
and UO_3325 (O_3325,N_29214,N_28822);
and UO_3326 (O_3326,N_28921,N_29842);
xor UO_3327 (O_3327,N_29390,N_28956);
nand UO_3328 (O_3328,N_29753,N_28908);
xnor UO_3329 (O_3329,N_29822,N_28908);
and UO_3330 (O_3330,N_29225,N_29133);
or UO_3331 (O_3331,N_28997,N_29126);
and UO_3332 (O_3332,N_29690,N_29422);
nand UO_3333 (O_3333,N_29462,N_29851);
xnor UO_3334 (O_3334,N_29177,N_29571);
nor UO_3335 (O_3335,N_29998,N_29555);
or UO_3336 (O_3336,N_29676,N_28810);
xnor UO_3337 (O_3337,N_29603,N_28930);
xnor UO_3338 (O_3338,N_29049,N_29494);
or UO_3339 (O_3339,N_29420,N_29430);
or UO_3340 (O_3340,N_29115,N_29553);
xnor UO_3341 (O_3341,N_29169,N_29856);
or UO_3342 (O_3342,N_28806,N_29129);
and UO_3343 (O_3343,N_28990,N_29074);
or UO_3344 (O_3344,N_29293,N_29108);
nand UO_3345 (O_3345,N_29684,N_29371);
and UO_3346 (O_3346,N_29430,N_29656);
xnor UO_3347 (O_3347,N_29573,N_29937);
and UO_3348 (O_3348,N_29864,N_29856);
nand UO_3349 (O_3349,N_29830,N_28944);
and UO_3350 (O_3350,N_29453,N_29108);
nand UO_3351 (O_3351,N_29579,N_29359);
or UO_3352 (O_3352,N_29661,N_28975);
nand UO_3353 (O_3353,N_29112,N_29137);
and UO_3354 (O_3354,N_29207,N_29962);
nor UO_3355 (O_3355,N_28861,N_29003);
or UO_3356 (O_3356,N_29319,N_29528);
and UO_3357 (O_3357,N_28909,N_28845);
and UO_3358 (O_3358,N_28935,N_29986);
and UO_3359 (O_3359,N_29309,N_29422);
and UO_3360 (O_3360,N_29554,N_29798);
nand UO_3361 (O_3361,N_29597,N_29185);
nor UO_3362 (O_3362,N_29891,N_29220);
nand UO_3363 (O_3363,N_29473,N_29199);
or UO_3364 (O_3364,N_29412,N_29005);
nor UO_3365 (O_3365,N_29076,N_29938);
and UO_3366 (O_3366,N_29826,N_29597);
xnor UO_3367 (O_3367,N_28877,N_29789);
or UO_3368 (O_3368,N_29941,N_29768);
nor UO_3369 (O_3369,N_29673,N_29799);
nand UO_3370 (O_3370,N_29956,N_29714);
nor UO_3371 (O_3371,N_29755,N_29684);
or UO_3372 (O_3372,N_29116,N_29958);
nand UO_3373 (O_3373,N_28959,N_29298);
or UO_3374 (O_3374,N_29097,N_29242);
nor UO_3375 (O_3375,N_29277,N_29027);
and UO_3376 (O_3376,N_29350,N_29454);
nor UO_3377 (O_3377,N_29743,N_29745);
nor UO_3378 (O_3378,N_29394,N_29407);
nand UO_3379 (O_3379,N_29577,N_29020);
xnor UO_3380 (O_3380,N_29291,N_29582);
nand UO_3381 (O_3381,N_29521,N_29829);
or UO_3382 (O_3382,N_29471,N_29140);
nor UO_3383 (O_3383,N_28970,N_29667);
or UO_3384 (O_3384,N_29497,N_29579);
nor UO_3385 (O_3385,N_29796,N_29575);
xor UO_3386 (O_3386,N_29425,N_29112);
or UO_3387 (O_3387,N_29567,N_29220);
nand UO_3388 (O_3388,N_28958,N_29207);
and UO_3389 (O_3389,N_29929,N_29026);
nor UO_3390 (O_3390,N_29944,N_29635);
and UO_3391 (O_3391,N_29240,N_29506);
and UO_3392 (O_3392,N_29653,N_28940);
nand UO_3393 (O_3393,N_29419,N_29284);
xnor UO_3394 (O_3394,N_29333,N_29417);
nor UO_3395 (O_3395,N_29935,N_29682);
nand UO_3396 (O_3396,N_29331,N_29536);
nand UO_3397 (O_3397,N_29003,N_29908);
and UO_3398 (O_3398,N_29271,N_29707);
or UO_3399 (O_3399,N_29367,N_29109);
or UO_3400 (O_3400,N_29354,N_29630);
nand UO_3401 (O_3401,N_29871,N_29790);
and UO_3402 (O_3402,N_29325,N_29026);
nand UO_3403 (O_3403,N_29762,N_28802);
nand UO_3404 (O_3404,N_29032,N_28829);
nand UO_3405 (O_3405,N_29535,N_29630);
or UO_3406 (O_3406,N_29248,N_28819);
nand UO_3407 (O_3407,N_29112,N_29388);
nor UO_3408 (O_3408,N_29715,N_29622);
nor UO_3409 (O_3409,N_29317,N_28828);
and UO_3410 (O_3410,N_29079,N_29766);
and UO_3411 (O_3411,N_29635,N_28817);
or UO_3412 (O_3412,N_29000,N_29102);
nor UO_3413 (O_3413,N_28863,N_28828);
or UO_3414 (O_3414,N_28854,N_28826);
xnor UO_3415 (O_3415,N_28981,N_28806);
nor UO_3416 (O_3416,N_29344,N_29413);
nand UO_3417 (O_3417,N_29471,N_29632);
nor UO_3418 (O_3418,N_29743,N_29470);
nor UO_3419 (O_3419,N_29728,N_29805);
and UO_3420 (O_3420,N_29630,N_29539);
nand UO_3421 (O_3421,N_29005,N_29112);
nor UO_3422 (O_3422,N_29734,N_29679);
xnor UO_3423 (O_3423,N_29485,N_29054);
nor UO_3424 (O_3424,N_29084,N_29733);
nand UO_3425 (O_3425,N_29981,N_29682);
nor UO_3426 (O_3426,N_29630,N_29976);
xor UO_3427 (O_3427,N_29079,N_29358);
or UO_3428 (O_3428,N_28970,N_28883);
or UO_3429 (O_3429,N_29773,N_28996);
xor UO_3430 (O_3430,N_29421,N_29779);
or UO_3431 (O_3431,N_29221,N_29535);
xor UO_3432 (O_3432,N_29047,N_29477);
and UO_3433 (O_3433,N_29848,N_29864);
nor UO_3434 (O_3434,N_29198,N_28976);
or UO_3435 (O_3435,N_28847,N_29405);
xor UO_3436 (O_3436,N_29569,N_29066);
nor UO_3437 (O_3437,N_28803,N_28812);
or UO_3438 (O_3438,N_29534,N_29575);
xor UO_3439 (O_3439,N_29042,N_29945);
and UO_3440 (O_3440,N_29064,N_29216);
and UO_3441 (O_3441,N_29667,N_29095);
or UO_3442 (O_3442,N_29527,N_29412);
and UO_3443 (O_3443,N_28850,N_29191);
or UO_3444 (O_3444,N_28801,N_29690);
nand UO_3445 (O_3445,N_28933,N_29346);
or UO_3446 (O_3446,N_28972,N_29212);
xnor UO_3447 (O_3447,N_29898,N_29919);
xnor UO_3448 (O_3448,N_29720,N_29552);
or UO_3449 (O_3449,N_28848,N_28978);
xor UO_3450 (O_3450,N_29962,N_29572);
nor UO_3451 (O_3451,N_29270,N_28819);
xnor UO_3452 (O_3452,N_29291,N_29778);
nor UO_3453 (O_3453,N_29675,N_29502);
nor UO_3454 (O_3454,N_29110,N_29600);
or UO_3455 (O_3455,N_29298,N_29487);
and UO_3456 (O_3456,N_28907,N_29343);
nor UO_3457 (O_3457,N_29494,N_29166);
xnor UO_3458 (O_3458,N_29796,N_29272);
nand UO_3459 (O_3459,N_29624,N_28907);
and UO_3460 (O_3460,N_29537,N_29926);
nor UO_3461 (O_3461,N_29682,N_29599);
nand UO_3462 (O_3462,N_28943,N_29608);
and UO_3463 (O_3463,N_28850,N_29131);
nand UO_3464 (O_3464,N_29914,N_29841);
xnor UO_3465 (O_3465,N_29502,N_29154);
nand UO_3466 (O_3466,N_29052,N_28831);
and UO_3467 (O_3467,N_29600,N_29074);
nand UO_3468 (O_3468,N_29970,N_29240);
xnor UO_3469 (O_3469,N_28912,N_29618);
and UO_3470 (O_3470,N_29196,N_29687);
xor UO_3471 (O_3471,N_29754,N_29746);
nor UO_3472 (O_3472,N_29445,N_29694);
nand UO_3473 (O_3473,N_29787,N_29049);
xnor UO_3474 (O_3474,N_28826,N_29675);
xor UO_3475 (O_3475,N_29174,N_28850);
and UO_3476 (O_3476,N_29900,N_29807);
xnor UO_3477 (O_3477,N_29436,N_29239);
and UO_3478 (O_3478,N_28842,N_28820);
nand UO_3479 (O_3479,N_29664,N_29436);
nand UO_3480 (O_3480,N_29298,N_29545);
or UO_3481 (O_3481,N_29605,N_29219);
nor UO_3482 (O_3482,N_29252,N_29266);
nor UO_3483 (O_3483,N_29587,N_29502);
xor UO_3484 (O_3484,N_29795,N_28849);
xor UO_3485 (O_3485,N_29758,N_29611);
nor UO_3486 (O_3486,N_29561,N_28860);
or UO_3487 (O_3487,N_29218,N_29928);
nand UO_3488 (O_3488,N_28891,N_29177);
xor UO_3489 (O_3489,N_29810,N_28981);
nand UO_3490 (O_3490,N_29202,N_28885);
nand UO_3491 (O_3491,N_29592,N_29573);
xor UO_3492 (O_3492,N_28938,N_29918);
nor UO_3493 (O_3493,N_29798,N_29355);
and UO_3494 (O_3494,N_29934,N_29279);
xor UO_3495 (O_3495,N_29367,N_29402);
and UO_3496 (O_3496,N_29629,N_29796);
xnor UO_3497 (O_3497,N_29490,N_28894);
or UO_3498 (O_3498,N_29941,N_29820);
nor UO_3499 (O_3499,N_29916,N_29965);
endmodule