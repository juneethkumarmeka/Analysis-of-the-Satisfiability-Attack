module basic_750_5000_1000_50_levels_2xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_459,In_646);
xor U1 (N_1,In_297,In_303);
or U2 (N_2,In_249,In_526);
and U3 (N_3,In_189,In_117);
nor U4 (N_4,In_559,In_164);
xor U5 (N_5,In_748,In_229);
nor U6 (N_6,In_364,In_190);
or U7 (N_7,In_617,In_165);
nand U8 (N_8,In_736,In_603);
nor U9 (N_9,In_644,In_132);
or U10 (N_10,In_264,In_708);
and U11 (N_11,In_10,In_524);
or U12 (N_12,In_284,In_51);
nand U13 (N_13,In_329,In_719);
or U14 (N_14,In_104,In_40);
and U15 (N_15,In_697,In_607);
nand U16 (N_16,In_677,In_182);
and U17 (N_17,In_722,In_73);
and U18 (N_18,In_274,In_246);
nand U19 (N_19,In_270,In_342);
or U20 (N_20,In_674,In_409);
or U21 (N_21,In_56,In_354);
nand U22 (N_22,In_8,In_433);
and U23 (N_23,In_363,In_95);
xnor U24 (N_24,In_590,In_248);
nor U25 (N_25,In_3,In_474);
xnor U26 (N_26,In_346,In_703);
and U27 (N_27,In_322,In_691);
or U28 (N_28,In_578,In_536);
and U29 (N_29,In_285,In_694);
nor U30 (N_30,In_307,In_67);
nand U31 (N_31,In_667,In_592);
or U32 (N_32,In_493,In_375);
or U33 (N_33,In_49,In_563);
and U34 (N_34,In_54,In_201);
and U35 (N_35,In_567,In_114);
or U36 (N_36,In_729,In_406);
and U37 (N_37,In_373,In_370);
or U38 (N_38,In_398,In_64);
or U39 (N_39,In_324,In_239);
and U40 (N_40,In_580,In_53);
nor U41 (N_41,In_135,In_689);
or U42 (N_42,In_491,In_449);
and U43 (N_43,In_129,In_629);
and U44 (N_44,In_14,In_365);
xnor U45 (N_45,In_296,In_41);
nor U46 (N_46,In_352,In_514);
nor U47 (N_47,In_315,In_328);
and U48 (N_48,In_181,In_392);
nor U49 (N_49,In_210,In_118);
nor U50 (N_50,In_441,In_747);
nand U51 (N_51,In_388,In_573);
or U52 (N_52,In_456,In_528);
or U53 (N_53,In_331,In_338);
nor U54 (N_54,In_688,In_205);
nand U55 (N_55,In_253,In_26);
xnor U56 (N_56,In_620,In_684);
and U57 (N_57,In_636,In_275);
or U58 (N_58,In_653,In_657);
nand U59 (N_59,In_672,In_568);
nor U60 (N_60,In_626,In_213);
nor U61 (N_61,In_22,In_538);
or U62 (N_62,In_675,In_487);
xor U63 (N_63,In_749,In_659);
or U64 (N_64,In_485,In_432);
or U65 (N_65,In_278,In_161);
or U66 (N_66,In_318,In_531);
nand U67 (N_67,In_612,In_44);
or U68 (N_68,In_125,In_709);
or U69 (N_69,In_577,In_665);
and U70 (N_70,In_304,In_469);
or U71 (N_71,In_453,In_214);
nand U72 (N_72,In_168,In_103);
nor U73 (N_73,In_735,In_276);
and U74 (N_74,In_481,In_654);
nand U75 (N_75,In_316,In_402);
or U76 (N_76,In_596,In_72);
nor U77 (N_77,In_692,In_298);
nor U78 (N_78,In_426,In_455);
and U79 (N_79,In_77,In_394);
xnor U80 (N_80,In_357,In_130);
nor U81 (N_81,In_341,In_725);
nand U82 (N_82,In_250,In_687);
nand U83 (N_83,In_154,In_434);
nor U84 (N_84,In_685,In_579);
nor U85 (N_85,In_660,In_673);
nor U86 (N_86,In_334,In_272);
or U87 (N_87,In_34,In_25);
nor U88 (N_88,In_153,In_712);
and U89 (N_89,In_497,In_256);
and U90 (N_90,In_427,In_705);
nand U91 (N_91,In_302,In_18);
or U92 (N_92,In_242,In_415);
nor U93 (N_93,In_390,In_696);
and U94 (N_94,In_61,In_199);
nand U95 (N_95,In_289,In_216);
xnor U96 (N_96,In_68,In_174);
or U97 (N_97,In_737,In_45);
nand U98 (N_98,In_136,In_281);
nor U99 (N_99,In_327,In_698);
and U100 (N_100,In_221,In_88);
nand U101 (N_101,In_312,In_115);
and U102 (N_102,N_19,In_509);
and U103 (N_103,In_499,In_177);
or U104 (N_104,In_55,In_510);
nor U105 (N_105,In_668,In_58);
nor U106 (N_106,In_360,In_158);
xnor U107 (N_107,In_183,In_70);
or U108 (N_108,In_385,N_96);
xnor U109 (N_109,In_410,In_448);
nand U110 (N_110,In_128,In_635);
nor U111 (N_111,N_15,In_400);
and U112 (N_112,In_506,In_314);
nand U113 (N_113,In_423,In_741);
nor U114 (N_114,In_126,In_358);
or U115 (N_115,In_720,In_621);
or U116 (N_116,In_669,In_141);
or U117 (N_117,In_9,In_157);
or U118 (N_118,In_82,In_560);
nand U119 (N_119,In_389,In_288);
xor U120 (N_120,N_41,In_268);
or U121 (N_121,In_191,N_85);
or U122 (N_122,In_173,N_95);
nor U123 (N_123,In_471,In_238);
nand U124 (N_124,In_57,In_727);
or U125 (N_125,In_219,In_504);
nand U126 (N_126,In_149,In_206);
nand U127 (N_127,In_468,N_39);
or U128 (N_128,N_30,In_624);
nand U129 (N_129,In_446,In_255);
or U130 (N_130,In_147,In_156);
nand U131 (N_131,In_337,In_148);
nor U132 (N_132,N_89,N_40);
or U133 (N_133,In_562,In_107);
nor U134 (N_134,N_20,In_584);
nand U135 (N_135,In_37,In_355);
nand U136 (N_136,In_31,N_93);
and U137 (N_137,In_325,In_627);
and U138 (N_138,In_421,N_67);
nor U139 (N_139,N_9,In_185);
nand U140 (N_140,In_106,In_273);
nor U141 (N_141,In_671,In_267);
and U142 (N_142,In_16,In_525);
and U143 (N_143,In_172,In_111);
or U144 (N_144,In_378,In_211);
or U145 (N_145,In_376,In_645);
and U146 (N_146,In_412,In_439);
nand U147 (N_147,In_15,In_176);
or U148 (N_148,In_223,In_81);
xor U149 (N_149,In_466,In_305);
nor U150 (N_150,N_57,In_102);
and U151 (N_151,In_383,In_532);
nor U152 (N_152,N_90,In_723);
or U153 (N_153,In_39,In_245);
nor U154 (N_154,In_593,In_407);
nand U155 (N_155,In_680,N_59);
and U156 (N_156,In_230,In_699);
or U157 (N_157,N_16,In_43);
and U158 (N_158,In_399,In_537);
and U159 (N_159,In_226,N_97);
or U160 (N_160,N_68,In_279);
or U161 (N_161,In_236,N_14);
nand U162 (N_162,In_353,In_196);
xor U163 (N_163,In_333,In_171);
and U164 (N_164,In_343,In_556);
xor U165 (N_165,In_554,In_724);
or U166 (N_166,In_379,N_88);
and U167 (N_167,In_451,In_101);
nand U168 (N_168,N_53,In_489);
nor U169 (N_169,In_260,In_252);
or U170 (N_170,In_637,In_23);
or U171 (N_171,In_6,In_583);
nor U172 (N_172,In_571,In_293);
or U173 (N_173,In_743,In_21);
nor U174 (N_174,N_12,In_12);
or U175 (N_175,N_8,N_65);
nand U176 (N_176,N_74,In_552);
nand U177 (N_177,In_367,In_732);
nand U178 (N_178,In_251,In_257);
or U179 (N_179,In_184,In_283);
xor U180 (N_180,N_98,In_344);
or U181 (N_181,In_372,In_643);
or U182 (N_182,In_47,In_461);
and U183 (N_183,In_369,N_2);
nand U184 (N_184,In_35,N_33);
and U185 (N_185,In_7,N_47);
nand U186 (N_186,In_122,In_457);
nand U187 (N_187,In_160,In_244);
and U188 (N_188,N_4,N_81);
and U189 (N_189,In_235,In_622);
and U190 (N_190,In_262,In_17);
or U191 (N_191,In_475,In_124);
and U192 (N_192,In_616,N_91);
and U193 (N_193,In_734,In_11);
xnor U194 (N_194,In_710,In_505);
nand U195 (N_195,In_313,In_166);
nor U196 (N_196,In_65,In_589);
or U197 (N_197,In_60,N_78);
nor U198 (N_198,In_460,In_19);
nand U199 (N_199,In_359,In_588);
nor U200 (N_200,N_54,N_42);
and U201 (N_201,In_5,In_83);
nand U202 (N_202,N_119,In_619);
nand U203 (N_203,In_140,In_495);
and U204 (N_204,In_100,In_381);
and U205 (N_205,N_162,In_96);
nor U206 (N_206,In_85,In_512);
or U207 (N_207,N_172,N_189);
nor U208 (N_208,In_76,N_108);
and U209 (N_209,N_140,In_467);
or U210 (N_210,N_167,In_564);
and U211 (N_211,N_173,In_714);
and U212 (N_212,In_349,In_530);
nor U213 (N_213,In_179,N_154);
nor U214 (N_214,In_430,N_182);
nand U215 (N_215,In_84,In_695);
nor U216 (N_216,N_21,In_437);
or U217 (N_217,In_187,In_693);
or U218 (N_218,N_66,N_23);
nor U219 (N_219,In_701,In_387);
and U220 (N_220,In_112,In_48);
nor U221 (N_221,In_280,N_24);
or U222 (N_222,In_27,N_70);
xor U223 (N_223,In_292,In_527);
nand U224 (N_224,In_595,In_553);
and U225 (N_225,In_247,N_191);
nor U226 (N_226,N_158,In_608);
and U227 (N_227,In_610,N_87);
and U228 (N_228,In_744,In_348);
nor U229 (N_229,N_132,N_174);
or U230 (N_230,N_64,In_80);
nor U231 (N_231,N_60,In_92);
nand U232 (N_232,In_638,In_424);
nor U233 (N_233,In_465,In_306);
or U234 (N_234,N_55,In_193);
nand U235 (N_235,N_139,N_178);
or U236 (N_236,N_50,In_332);
or U237 (N_237,In_404,In_75);
nor U238 (N_238,In_641,In_265);
nand U239 (N_239,In_731,N_192);
and U240 (N_240,N_113,In_414);
or U241 (N_241,N_123,In_702);
and U242 (N_242,In_613,In_91);
nor U243 (N_243,In_566,In_428);
or U244 (N_244,In_301,In_97);
and U245 (N_245,In_79,N_197);
or U246 (N_246,In_66,In_138);
nor U247 (N_247,In_78,In_87);
nand U248 (N_248,In_50,In_29);
nor U249 (N_249,N_45,In_59);
nor U250 (N_250,In_632,N_159);
nor U251 (N_251,In_452,In_227);
nand U252 (N_252,In_263,In_438);
and U253 (N_253,In_520,In_686);
nand U254 (N_254,N_69,In_217);
and U255 (N_255,N_46,In_631);
nand U256 (N_256,In_224,N_177);
nand U257 (N_257,In_287,N_34);
nor U258 (N_258,N_143,N_22);
nor U259 (N_259,In_682,In_24);
nor U260 (N_260,N_99,N_166);
nand U261 (N_261,In_46,N_161);
nor U262 (N_262,In_71,N_104);
nand U263 (N_263,In_311,N_6);
and U264 (N_264,In_728,In_110);
and U265 (N_265,In_733,N_129);
nand U266 (N_266,N_138,In_462);
or U267 (N_267,N_29,In_561);
nand U268 (N_268,In_522,N_28);
and U269 (N_269,In_548,In_266);
nand U270 (N_270,In_642,In_715);
or U271 (N_271,N_36,In_557);
and U272 (N_272,N_196,In_175);
nand U273 (N_273,In_13,In_739);
and U274 (N_274,In_420,In_707);
or U275 (N_275,In_0,In_258);
nor U276 (N_276,In_33,In_625);
nand U277 (N_277,In_551,In_116);
or U278 (N_278,In_99,In_546);
nor U279 (N_279,N_115,In_678);
or U280 (N_280,In_194,In_347);
nand U281 (N_281,N_117,In_738);
or U282 (N_282,In_170,In_339);
or U283 (N_283,In_317,N_121);
or U284 (N_284,N_125,In_123);
nor U285 (N_285,N_185,N_71);
nand U286 (N_286,In_565,In_572);
or U287 (N_287,In_28,N_48);
and U288 (N_288,In_483,N_175);
xnor U289 (N_289,N_109,In_628);
or U290 (N_290,In_144,In_458);
or U291 (N_291,In_215,N_195);
nor U292 (N_292,In_146,In_52);
nor U293 (N_293,In_615,N_114);
nor U294 (N_294,In_105,N_112);
or U295 (N_295,N_151,In_134);
nor U296 (N_296,In_716,N_94);
or U297 (N_297,In_178,N_92);
and U298 (N_298,N_120,In_501);
nor U299 (N_299,N_26,N_61);
nand U300 (N_300,N_211,In_361);
or U301 (N_301,In_374,In_547);
or U302 (N_302,N_253,In_472);
or U303 (N_303,N_126,In_366);
nor U304 (N_304,In_609,In_648);
nand U305 (N_305,N_141,N_246);
xnor U306 (N_306,In_290,In_425);
or U307 (N_307,In_651,In_600);
nand U308 (N_308,In_517,In_198);
nand U309 (N_309,In_746,In_42);
nand U310 (N_310,In_323,N_13);
or U311 (N_311,In_188,N_106);
nor U312 (N_312,In_435,In_575);
nand U313 (N_313,In_454,N_221);
and U314 (N_314,N_5,N_200);
nor U315 (N_315,In_336,N_179);
or U316 (N_316,N_241,N_282);
and U317 (N_317,N_204,In_486);
and U318 (N_318,N_283,In_507);
or U319 (N_319,In_241,N_248);
and U320 (N_320,N_18,N_77);
nor U321 (N_321,In_220,N_226);
nor U322 (N_322,In_38,N_233);
and U323 (N_323,In_391,N_133);
or U324 (N_324,N_199,In_601);
nand U325 (N_325,N_203,N_270);
nand U326 (N_326,N_144,In_650);
nand U327 (N_327,In_192,In_320);
or U328 (N_328,N_205,In_259);
or U329 (N_329,N_231,N_86);
nor U330 (N_330,In_569,N_38);
nor U331 (N_331,In_291,N_100);
or U332 (N_332,In_422,N_103);
or U333 (N_333,N_296,In_2);
and U334 (N_334,In_606,In_647);
and U335 (N_335,In_145,In_585);
and U336 (N_336,In_431,N_152);
nor U337 (N_337,In_405,N_238);
and U338 (N_338,In_534,N_130);
nor U339 (N_339,N_214,In_277);
xnor U340 (N_340,N_116,N_142);
and U341 (N_341,In_202,N_237);
nor U342 (N_342,In_395,In_121);
xnor U343 (N_343,N_217,N_35);
nand U344 (N_344,In_535,In_598);
and U345 (N_345,In_150,In_479);
and U346 (N_346,N_150,N_193);
nor U347 (N_347,N_213,In_594);
nand U348 (N_348,N_273,In_113);
and U349 (N_349,In_62,N_7);
or U350 (N_350,N_279,In_418);
nand U351 (N_351,In_683,N_275);
nand U352 (N_352,In_208,In_614);
nor U353 (N_353,N_52,N_239);
and U354 (N_354,N_297,In_386);
or U355 (N_355,In_679,In_294);
and U356 (N_356,In_321,In_233);
nand U357 (N_357,In_232,In_740);
nand U358 (N_358,N_235,N_25);
or U359 (N_359,In_602,N_223);
and U360 (N_360,N_80,In_384);
nor U361 (N_361,In_429,N_146);
and U362 (N_362,In_652,In_162);
and U363 (N_363,In_502,In_203);
or U364 (N_364,In_351,In_704);
nor U365 (N_365,In_450,N_181);
or U366 (N_366,In_237,In_151);
nor U367 (N_367,N_222,N_194);
nand U368 (N_368,In_340,In_20);
or U369 (N_369,N_267,In_139);
nor U370 (N_370,N_274,In_717);
nor U371 (N_371,In_167,In_666);
or U372 (N_372,In_403,N_201);
or U373 (N_373,In_380,In_180);
or U374 (N_374,N_134,In_261);
and U375 (N_375,N_288,In_549);
and U376 (N_376,N_176,In_591);
nand U377 (N_377,In_243,N_298);
nor U378 (N_378,N_83,N_252);
and U379 (N_379,In_396,N_148);
nand U380 (N_380,In_271,N_276);
and U381 (N_381,In_36,N_281);
or U382 (N_382,In_498,In_543);
and U383 (N_383,In_401,In_131);
and U384 (N_384,In_300,In_195);
and U385 (N_385,In_670,N_230);
or U386 (N_386,In_4,N_157);
or U387 (N_387,In_408,In_478);
and U388 (N_388,N_245,N_17);
or U389 (N_389,N_266,In_663);
and U390 (N_390,In_254,N_198);
or U391 (N_391,In_119,In_661);
or U392 (N_392,N_206,In_599);
nand U393 (N_393,In_513,N_163);
xnor U394 (N_394,N_72,N_287);
nor U395 (N_395,In_204,In_633);
nand U396 (N_396,N_215,N_294);
or U397 (N_397,N_180,N_153);
or U398 (N_398,In_611,N_10);
nand U399 (N_399,N_11,N_299);
and U400 (N_400,In_545,N_155);
and U401 (N_401,N_271,In_93);
nand U402 (N_402,N_269,In_586);
nor U403 (N_403,N_372,N_236);
and U404 (N_404,In_269,In_681);
xor U405 (N_405,N_171,N_102);
nor U406 (N_406,In_368,N_122);
nand U407 (N_407,In_382,In_664);
nor U408 (N_408,N_316,N_327);
and U409 (N_409,N_347,N_396);
and U410 (N_410,N_389,In_89);
nand U411 (N_411,N_128,N_278);
nor U412 (N_412,In_477,N_188);
nand U413 (N_413,N_355,N_261);
and U414 (N_414,N_262,In_186);
or U415 (N_415,N_118,In_662);
and U416 (N_416,N_247,N_345);
nor U417 (N_417,N_292,In_496);
or U418 (N_418,N_349,N_111);
or U419 (N_419,N_361,N_331);
nor U420 (N_420,N_322,N_351);
nor U421 (N_421,N_376,In_444);
and U422 (N_422,N_326,N_310);
or U423 (N_423,In_464,In_605);
and U424 (N_424,In_630,In_533);
and U425 (N_425,In_445,In_350);
and U426 (N_426,N_391,N_308);
nor U427 (N_427,N_343,N_380);
or U428 (N_428,N_284,N_265);
nor U429 (N_429,In_209,N_381);
or U430 (N_430,In_443,N_263);
or U431 (N_431,N_306,N_369);
and U432 (N_432,N_346,N_320);
or U433 (N_433,In_529,In_94);
or U434 (N_434,In_745,N_318);
and U435 (N_435,In_713,N_0);
nand U436 (N_436,In_442,N_313);
or U437 (N_437,In_1,In_228);
nor U438 (N_438,In_623,In_480);
or U439 (N_439,In_676,N_232);
and U440 (N_440,In_523,N_377);
nand U441 (N_441,N_291,In_411);
or U442 (N_442,N_300,N_110);
and U443 (N_443,N_229,N_228);
or U444 (N_444,In_133,In_159);
and U445 (N_445,N_341,In_63);
or U446 (N_446,N_354,N_136);
or U447 (N_447,N_301,N_249);
or U448 (N_448,N_302,N_49);
and U449 (N_449,In_393,In_447);
nand U450 (N_450,N_368,N_290);
xor U451 (N_451,In_440,In_711);
or U452 (N_452,In_30,N_367);
nor U453 (N_453,In_511,N_286);
nor U454 (N_454,In_463,In_582);
and U455 (N_455,N_186,N_360);
nor U456 (N_456,N_319,In_212);
nor U457 (N_457,In_362,N_348);
and U458 (N_458,N_107,N_335);
nand U459 (N_459,In_730,N_309);
nand U460 (N_460,In_508,N_168);
nand U461 (N_461,In_234,N_105);
nand U462 (N_462,N_165,N_329);
nor U463 (N_463,In_299,In_518);
nor U464 (N_464,In_127,N_342);
nor U465 (N_465,N_295,In_492);
nand U466 (N_466,In_482,N_3);
nand U467 (N_467,N_73,In_516);
nand U468 (N_468,N_219,N_190);
nor U469 (N_469,In_690,In_155);
nor U470 (N_470,In_413,N_280);
nor U471 (N_471,In_587,In_706);
nor U472 (N_472,In_576,N_51);
and U473 (N_473,In_310,N_137);
nor U474 (N_474,In_503,N_220);
nor U475 (N_475,N_124,N_210);
xnor U476 (N_476,N_75,N_383);
or U477 (N_477,N_164,N_251);
or U478 (N_478,N_135,N_315);
or U479 (N_479,In_200,In_597);
or U480 (N_480,N_340,In_640);
or U481 (N_481,N_337,N_390);
nand U482 (N_482,In_143,N_386);
and U483 (N_483,N_258,N_37);
and U484 (N_484,N_359,In_604);
and U485 (N_485,In_488,N_240);
and U486 (N_486,N_255,N_339);
and U487 (N_487,In_335,In_541);
nand U488 (N_488,In_377,In_558);
nand U489 (N_489,In_86,N_285);
and U490 (N_490,In_581,In_417);
nand U491 (N_491,N_366,N_392);
nor U492 (N_492,In_225,N_388);
nor U493 (N_493,N_311,In_169);
or U494 (N_494,N_314,N_382);
nand U495 (N_495,N_32,N_272);
nor U496 (N_496,In_397,N_31);
nand U497 (N_497,N_208,In_718);
or U498 (N_498,In_319,N_330);
xnor U499 (N_499,In_419,N_324);
and U500 (N_500,N_387,N_234);
nor U501 (N_501,N_460,N_499);
nand U502 (N_502,N_452,N_437);
or U503 (N_503,N_356,N_187);
or U504 (N_504,In_550,N_491);
or U505 (N_505,N_259,N_464);
nor U506 (N_506,N_76,N_403);
nor U507 (N_507,N_471,N_477);
nor U508 (N_508,N_462,N_183);
nor U509 (N_509,In_282,N_394);
nor U510 (N_510,In_634,N_486);
or U511 (N_511,N_370,N_438);
nor U512 (N_512,N_225,In_473);
nor U513 (N_513,N_489,N_439);
nor U514 (N_514,In_618,N_469);
nor U515 (N_515,N_427,In_137);
nor U516 (N_516,N_227,N_257);
nor U517 (N_517,N_58,In_286);
nor U518 (N_518,N_467,N_454);
and U519 (N_519,N_304,N_364);
or U520 (N_520,N_357,N_393);
and U521 (N_521,In_90,N_451);
nand U522 (N_522,N_411,N_498);
nor U523 (N_523,N_317,N_293);
xnor U524 (N_524,N_307,N_435);
nor U525 (N_525,N_425,N_260);
and U526 (N_526,N_374,N_127);
nand U527 (N_527,In_726,In_542);
and U528 (N_528,N_432,In_570);
nor U529 (N_529,N_242,N_420);
and U530 (N_530,In_163,In_539);
and U531 (N_531,N_493,N_1);
and U532 (N_532,N_145,N_365);
nand U533 (N_533,N_268,N_422);
and U534 (N_534,In_544,N_218);
nor U535 (N_535,N_413,In_656);
nand U536 (N_536,N_475,N_43);
nor U537 (N_537,In_218,N_338);
or U538 (N_538,N_375,N_379);
and U539 (N_539,N_400,In_197);
or U540 (N_540,N_56,N_332);
nor U541 (N_541,N_484,N_428);
or U542 (N_542,In_152,N_494);
nand U543 (N_543,N_463,N_418);
nand U544 (N_544,N_79,In_655);
nor U545 (N_545,N_402,N_419);
nor U546 (N_546,N_373,In_519);
or U547 (N_547,N_256,N_449);
nand U548 (N_548,In_356,N_455);
nor U549 (N_549,N_264,N_434);
and U550 (N_550,N_82,N_212);
nor U551 (N_551,N_149,In_500);
nand U552 (N_552,N_344,N_352);
nand U553 (N_553,N_385,N_417);
or U554 (N_554,In_490,In_309);
nand U555 (N_555,N_414,N_416);
or U556 (N_556,In_371,N_336);
nand U557 (N_557,N_325,In_98);
nand U558 (N_558,N_453,N_209);
and U559 (N_559,N_458,N_488);
nor U560 (N_560,N_457,N_430);
nor U561 (N_561,In_484,N_131);
nor U562 (N_562,N_490,N_456);
nor U563 (N_563,N_481,N_443);
nand U564 (N_564,In_515,In_555);
xnor U565 (N_565,N_371,N_409);
and U566 (N_566,N_424,N_480);
or U567 (N_567,In_742,In_326);
nand U568 (N_568,N_429,N_224);
and U569 (N_569,N_412,N_436);
and U570 (N_570,N_470,N_479);
and U571 (N_571,In_308,N_243);
nor U572 (N_572,N_447,In_470);
and U573 (N_573,N_170,N_450);
nor U574 (N_574,N_353,N_358);
nor U575 (N_575,In_32,In_120);
and U576 (N_576,N_495,N_482);
and U577 (N_577,N_433,N_250);
nor U578 (N_578,N_277,In_74);
or U579 (N_579,N_63,N_431);
nand U580 (N_580,N_483,In_207);
nand U581 (N_581,N_444,N_334);
or U582 (N_582,N_384,In_721);
nand U583 (N_583,N_321,N_440);
nand U584 (N_584,N_378,N_207);
nand U585 (N_585,N_487,N_363);
nand U586 (N_586,N_350,N_305);
nor U587 (N_587,N_473,N_398);
nand U588 (N_588,N_147,In_540);
and U589 (N_589,In_436,N_303);
or U590 (N_590,N_406,N_492);
nor U591 (N_591,N_395,N_468);
and U592 (N_592,N_216,N_44);
or U593 (N_593,In_416,N_442);
and U594 (N_594,N_101,N_84);
nand U595 (N_595,N_423,In_658);
or U596 (N_596,N_497,N_408);
nand U597 (N_597,N_407,In_69);
and U598 (N_598,N_496,N_399);
and U599 (N_599,N_472,In_240);
nand U600 (N_600,N_564,N_156);
nor U601 (N_601,N_546,N_549);
nor U602 (N_602,N_536,N_244);
and U603 (N_603,N_555,N_571);
nand U604 (N_604,N_590,N_515);
xor U605 (N_605,In_574,N_542);
xnor U606 (N_606,N_563,N_511);
and U607 (N_607,N_476,N_593);
nor U608 (N_608,N_551,N_589);
nand U609 (N_609,N_531,N_538);
or U610 (N_610,N_574,N_27);
nor U611 (N_611,N_585,N_202);
xor U612 (N_612,N_508,N_459);
or U613 (N_613,N_501,N_500);
and U614 (N_614,N_333,In_222);
nand U615 (N_615,N_405,N_441);
and U616 (N_616,N_502,N_410);
or U617 (N_617,N_362,N_598);
nand U618 (N_618,N_62,N_583);
or U619 (N_619,N_503,N_510);
or U620 (N_620,N_597,N_596);
or U621 (N_621,N_506,N_576);
nand U622 (N_622,N_592,N_573);
nand U623 (N_623,N_528,N_530);
or U624 (N_624,In_142,In_330);
nand U625 (N_625,N_512,N_560);
nand U626 (N_626,N_540,N_523);
and U627 (N_627,N_594,N_513);
and U628 (N_628,N_577,N_586);
nor U629 (N_629,N_580,In_494);
xor U630 (N_630,N_565,N_547);
nand U631 (N_631,N_507,N_397);
nor U632 (N_632,N_567,N_529);
or U633 (N_633,N_527,N_505);
nor U634 (N_634,N_461,N_570);
and U635 (N_635,N_509,N_543);
nand U636 (N_636,N_552,N_595);
nor U637 (N_637,In_639,N_466);
nand U638 (N_638,N_520,In_345);
nor U639 (N_639,In_649,N_578);
or U640 (N_640,N_553,N_289);
and U641 (N_641,N_525,N_584);
or U642 (N_642,N_558,N_474);
and U643 (N_643,N_514,In_108);
nand U644 (N_644,N_537,N_478);
nor U645 (N_645,N_445,N_562);
and U646 (N_646,N_519,N_569);
nor U647 (N_647,N_517,N_404);
or U648 (N_648,N_485,N_591);
xnor U649 (N_649,N_581,In_521);
and U650 (N_650,N_579,N_522);
and U651 (N_651,N_328,N_524);
and U652 (N_652,N_254,N_534);
nand U653 (N_653,N_446,N_184);
and U654 (N_654,N_426,In_295);
xnor U655 (N_655,In_109,N_572);
nand U656 (N_656,In_700,N_312);
or U657 (N_657,N_575,N_539);
and U658 (N_658,N_401,N_544);
nor U659 (N_659,N_532,N_599);
nand U660 (N_660,N_516,N_556);
nand U661 (N_661,N_526,N_550);
nor U662 (N_662,N_541,N_533);
or U663 (N_663,N_587,N_548);
xnor U664 (N_664,N_588,N_465);
nor U665 (N_665,N_554,N_557);
nand U666 (N_666,N_421,N_169);
nor U667 (N_667,N_566,N_323);
nand U668 (N_668,N_545,N_561);
nand U669 (N_669,In_476,In_231);
or U670 (N_670,N_582,N_160);
nand U671 (N_671,N_535,N_568);
nand U672 (N_672,N_504,N_521);
and U673 (N_673,N_415,N_448);
and U674 (N_674,N_518,N_559);
and U675 (N_675,In_494,N_485);
nand U676 (N_676,N_585,N_546);
or U677 (N_677,N_590,N_474);
nand U678 (N_678,N_503,N_502);
and U679 (N_679,N_465,N_574);
nor U680 (N_680,N_466,N_543);
nand U681 (N_681,N_596,N_548);
or U682 (N_682,N_545,N_519);
nor U683 (N_683,In_639,N_550);
or U684 (N_684,N_554,N_551);
and U685 (N_685,N_521,In_521);
or U686 (N_686,N_574,N_579);
and U687 (N_687,In_222,N_62);
nor U688 (N_688,N_535,N_558);
and U689 (N_689,N_527,N_254);
nor U690 (N_690,N_529,N_596);
nand U691 (N_691,N_567,N_539);
nand U692 (N_692,N_513,N_579);
xnor U693 (N_693,N_578,N_596);
nor U694 (N_694,N_534,N_510);
or U695 (N_695,N_530,N_583);
or U696 (N_696,N_587,N_404);
nor U697 (N_697,N_524,In_521);
xor U698 (N_698,In_231,N_575);
and U699 (N_699,N_520,N_461);
and U700 (N_700,N_602,N_637);
nand U701 (N_701,N_650,N_629);
and U702 (N_702,N_679,N_625);
nor U703 (N_703,N_661,N_645);
and U704 (N_704,N_609,N_627);
nor U705 (N_705,N_657,N_655);
nor U706 (N_706,N_663,N_692);
nand U707 (N_707,N_611,N_667);
and U708 (N_708,N_668,N_605);
and U709 (N_709,N_684,N_606);
or U710 (N_710,N_699,N_672);
nor U711 (N_711,N_669,N_673);
or U712 (N_712,N_632,N_656);
and U713 (N_713,N_666,N_665);
nor U714 (N_714,N_610,N_630);
nor U715 (N_715,N_628,N_634);
nor U716 (N_716,N_643,N_674);
or U717 (N_717,N_604,N_618);
and U718 (N_718,N_659,N_608);
or U719 (N_719,N_614,N_664);
nor U720 (N_720,N_631,N_623);
or U721 (N_721,N_658,N_678);
and U722 (N_722,N_646,N_683);
or U723 (N_723,N_698,N_607);
nand U724 (N_724,N_603,N_621);
nor U725 (N_725,N_697,N_696);
and U726 (N_726,N_662,N_686);
or U727 (N_727,N_681,N_651);
and U728 (N_728,N_671,N_653);
or U729 (N_729,N_615,N_691);
nor U730 (N_730,N_641,N_654);
or U731 (N_731,N_693,N_617);
or U732 (N_732,N_670,N_633);
nand U733 (N_733,N_694,N_695);
or U734 (N_734,N_660,N_600);
nand U735 (N_735,N_613,N_644);
nor U736 (N_736,N_626,N_639);
or U737 (N_737,N_642,N_690);
nor U738 (N_738,N_635,N_619);
nand U739 (N_739,N_647,N_675);
or U740 (N_740,N_649,N_688);
and U741 (N_741,N_680,N_685);
or U742 (N_742,N_612,N_622);
nor U743 (N_743,N_620,N_640);
nor U744 (N_744,N_687,N_601);
or U745 (N_745,N_636,N_682);
and U746 (N_746,N_689,N_677);
nor U747 (N_747,N_652,N_648);
nor U748 (N_748,N_616,N_624);
or U749 (N_749,N_638,N_676);
nor U750 (N_750,N_644,N_618);
and U751 (N_751,N_697,N_648);
nor U752 (N_752,N_686,N_622);
nand U753 (N_753,N_651,N_631);
nor U754 (N_754,N_612,N_641);
and U755 (N_755,N_640,N_684);
or U756 (N_756,N_604,N_688);
nand U757 (N_757,N_677,N_629);
nor U758 (N_758,N_619,N_616);
nand U759 (N_759,N_615,N_620);
nor U760 (N_760,N_630,N_694);
nand U761 (N_761,N_686,N_617);
and U762 (N_762,N_657,N_624);
and U763 (N_763,N_642,N_670);
nand U764 (N_764,N_672,N_667);
xor U765 (N_765,N_668,N_696);
or U766 (N_766,N_612,N_682);
nor U767 (N_767,N_602,N_687);
and U768 (N_768,N_628,N_688);
or U769 (N_769,N_637,N_624);
or U770 (N_770,N_647,N_625);
xnor U771 (N_771,N_669,N_675);
nor U772 (N_772,N_623,N_648);
nand U773 (N_773,N_655,N_608);
nor U774 (N_774,N_699,N_693);
nand U775 (N_775,N_678,N_612);
nor U776 (N_776,N_681,N_644);
or U777 (N_777,N_650,N_683);
or U778 (N_778,N_610,N_694);
or U779 (N_779,N_666,N_681);
and U780 (N_780,N_695,N_629);
or U781 (N_781,N_678,N_693);
or U782 (N_782,N_633,N_671);
or U783 (N_783,N_615,N_611);
or U784 (N_784,N_629,N_684);
nor U785 (N_785,N_688,N_694);
or U786 (N_786,N_662,N_609);
and U787 (N_787,N_605,N_696);
nand U788 (N_788,N_698,N_616);
and U789 (N_789,N_642,N_637);
nor U790 (N_790,N_621,N_661);
or U791 (N_791,N_672,N_617);
or U792 (N_792,N_649,N_661);
or U793 (N_793,N_608,N_688);
or U794 (N_794,N_627,N_611);
or U795 (N_795,N_675,N_688);
nand U796 (N_796,N_656,N_619);
xor U797 (N_797,N_697,N_645);
or U798 (N_798,N_625,N_669);
or U799 (N_799,N_627,N_621);
or U800 (N_800,N_718,N_746);
nor U801 (N_801,N_776,N_708);
nor U802 (N_802,N_745,N_792);
and U803 (N_803,N_709,N_756);
nor U804 (N_804,N_759,N_700);
nand U805 (N_805,N_783,N_790);
or U806 (N_806,N_740,N_764);
or U807 (N_807,N_748,N_772);
nor U808 (N_808,N_777,N_744);
and U809 (N_809,N_780,N_755);
nand U810 (N_810,N_762,N_771);
nand U811 (N_811,N_795,N_785);
and U812 (N_812,N_722,N_714);
nand U813 (N_813,N_770,N_768);
nand U814 (N_814,N_774,N_702);
nor U815 (N_815,N_710,N_728);
nor U816 (N_816,N_742,N_712);
nor U817 (N_817,N_723,N_743);
and U818 (N_818,N_791,N_711);
nand U819 (N_819,N_765,N_719);
nor U820 (N_820,N_731,N_734);
nand U821 (N_821,N_757,N_775);
and U822 (N_822,N_736,N_766);
nand U823 (N_823,N_752,N_788);
nor U824 (N_824,N_758,N_721);
nor U825 (N_825,N_727,N_703);
or U826 (N_826,N_751,N_781);
nand U827 (N_827,N_707,N_761);
nor U828 (N_828,N_729,N_773);
nand U829 (N_829,N_705,N_701);
or U830 (N_830,N_778,N_716);
xor U831 (N_831,N_749,N_787);
nor U832 (N_832,N_706,N_767);
or U833 (N_833,N_720,N_799);
or U834 (N_834,N_763,N_733);
or U835 (N_835,N_779,N_753);
and U836 (N_836,N_713,N_735);
nand U837 (N_837,N_747,N_717);
nand U838 (N_838,N_704,N_798);
or U839 (N_839,N_796,N_741);
nand U840 (N_840,N_789,N_726);
and U841 (N_841,N_760,N_739);
nor U842 (N_842,N_732,N_737);
nor U843 (N_843,N_794,N_724);
or U844 (N_844,N_750,N_784);
and U845 (N_845,N_730,N_715);
nand U846 (N_846,N_769,N_725);
nor U847 (N_847,N_754,N_782);
and U848 (N_848,N_793,N_797);
nor U849 (N_849,N_738,N_786);
or U850 (N_850,N_769,N_794);
nor U851 (N_851,N_720,N_748);
or U852 (N_852,N_741,N_712);
nand U853 (N_853,N_741,N_771);
nor U854 (N_854,N_799,N_746);
or U855 (N_855,N_750,N_759);
or U856 (N_856,N_729,N_755);
nor U857 (N_857,N_775,N_765);
nor U858 (N_858,N_795,N_734);
xor U859 (N_859,N_716,N_771);
nand U860 (N_860,N_706,N_709);
nor U861 (N_861,N_764,N_786);
nand U862 (N_862,N_739,N_708);
or U863 (N_863,N_744,N_764);
or U864 (N_864,N_742,N_799);
or U865 (N_865,N_758,N_782);
or U866 (N_866,N_733,N_799);
nor U867 (N_867,N_707,N_726);
nor U868 (N_868,N_781,N_757);
nor U869 (N_869,N_794,N_712);
or U870 (N_870,N_734,N_721);
nor U871 (N_871,N_720,N_753);
and U872 (N_872,N_706,N_795);
or U873 (N_873,N_786,N_713);
nand U874 (N_874,N_750,N_755);
or U875 (N_875,N_700,N_771);
nand U876 (N_876,N_755,N_763);
nand U877 (N_877,N_712,N_757);
and U878 (N_878,N_722,N_751);
or U879 (N_879,N_770,N_736);
and U880 (N_880,N_782,N_762);
and U881 (N_881,N_767,N_777);
nor U882 (N_882,N_705,N_727);
and U883 (N_883,N_790,N_728);
xnor U884 (N_884,N_714,N_756);
or U885 (N_885,N_767,N_791);
and U886 (N_886,N_732,N_779);
nor U887 (N_887,N_781,N_729);
nor U888 (N_888,N_777,N_781);
nand U889 (N_889,N_738,N_793);
nor U890 (N_890,N_766,N_768);
nand U891 (N_891,N_764,N_768);
or U892 (N_892,N_756,N_778);
or U893 (N_893,N_732,N_703);
xor U894 (N_894,N_709,N_798);
nor U895 (N_895,N_749,N_735);
nand U896 (N_896,N_726,N_799);
nand U897 (N_897,N_771,N_795);
and U898 (N_898,N_761,N_734);
and U899 (N_899,N_735,N_721);
xor U900 (N_900,N_867,N_875);
nand U901 (N_901,N_887,N_822);
nand U902 (N_902,N_874,N_825);
nor U903 (N_903,N_892,N_808);
and U904 (N_904,N_800,N_894);
nor U905 (N_905,N_878,N_877);
or U906 (N_906,N_827,N_873);
nand U907 (N_907,N_841,N_820);
or U908 (N_908,N_809,N_835);
or U909 (N_909,N_858,N_834);
nor U910 (N_910,N_816,N_885);
nor U911 (N_911,N_831,N_859);
or U912 (N_912,N_861,N_828);
nand U913 (N_913,N_871,N_872);
or U914 (N_914,N_882,N_824);
or U915 (N_915,N_863,N_847);
and U916 (N_916,N_837,N_851);
or U917 (N_917,N_850,N_817);
nand U918 (N_918,N_854,N_832);
and U919 (N_919,N_826,N_853);
or U920 (N_920,N_844,N_899);
and U921 (N_921,N_807,N_889);
nand U922 (N_922,N_890,N_860);
nand U923 (N_923,N_866,N_865);
or U924 (N_924,N_893,N_840);
or U925 (N_925,N_838,N_836);
and U926 (N_926,N_842,N_843);
and U927 (N_927,N_833,N_830);
and U928 (N_928,N_849,N_857);
and U929 (N_929,N_898,N_888);
or U930 (N_930,N_879,N_805);
nor U931 (N_931,N_855,N_896);
and U932 (N_932,N_848,N_846);
and U933 (N_933,N_880,N_870);
and U934 (N_934,N_812,N_823);
nor U935 (N_935,N_814,N_862);
nor U936 (N_936,N_802,N_868);
nor U937 (N_937,N_891,N_884);
or U938 (N_938,N_818,N_801);
and U939 (N_939,N_821,N_829);
nor U940 (N_940,N_845,N_804);
or U941 (N_941,N_869,N_819);
nand U942 (N_942,N_856,N_864);
nand U943 (N_943,N_881,N_810);
nor U944 (N_944,N_813,N_806);
and U945 (N_945,N_811,N_803);
nor U946 (N_946,N_897,N_883);
nand U947 (N_947,N_876,N_852);
and U948 (N_948,N_815,N_886);
nand U949 (N_949,N_895,N_839);
nor U950 (N_950,N_885,N_890);
or U951 (N_951,N_812,N_867);
or U952 (N_952,N_811,N_868);
nor U953 (N_953,N_861,N_886);
nand U954 (N_954,N_869,N_823);
and U955 (N_955,N_805,N_838);
and U956 (N_956,N_839,N_825);
nor U957 (N_957,N_874,N_813);
nand U958 (N_958,N_813,N_884);
nor U959 (N_959,N_872,N_864);
or U960 (N_960,N_867,N_861);
or U961 (N_961,N_828,N_856);
and U962 (N_962,N_873,N_800);
nor U963 (N_963,N_815,N_821);
nand U964 (N_964,N_829,N_875);
or U965 (N_965,N_887,N_873);
and U966 (N_966,N_868,N_884);
nor U967 (N_967,N_805,N_835);
or U968 (N_968,N_817,N_889);
and U969 (N_969,N_860,N_817);
or U970 (N_970,N_815,N_833);
and U971 (N_971,N_824,N_873);
nand U972 (N_972,N_807,N_874);
nand U973 (N_973,N_828,N_848);
nand U974 (N_974,N_815,N_888);
and U975 (N_975,N_890,N_879);
xnor U976 (N_976,N_876,N_871);
nor U977 (N_977,N_888,N_821);
nand U978 (N_978,N_830,N_877);
nand U979 (N_979,N_817,N_803);
and U980 (N_980,N_881,N_816);
nor U981 (N_981,N_896,N_831);
nand U982 (N_982,N_863,N_835);
or U983 (N_983,N_847,N_874);
nor U984 (N_984,N_847,N_827);
or U985 (N_985,N_860,N_858);
and U986 (N_986,N_802,N_849);
or U987 (N_987,N_839,N_878);
nand U988 (N_988,N_803,N_805);
and U989 (N_989,N_825,N_850);
nand U990 (N_990,N_891,N_814);
or U991 (N_991,N_895,N_809);
nand U992 (N_992,N_859,N_857);
or U993 (N_993,N_848,N_822);
and U994 (N_994,N_887,N_856);
or U995 (N_995,N_840,N_819);
or U996 (N_996,N_897,N_894);
nand U997 (N_997,N_888,N_819);
nand U998 (N_998,N_811,N_831);
or U999 (N_999,N_826,N_801);
and U1000 (N_1000,N_937,N_950);
nor U1001 (N_1001,N_946,N_989);
nand U1002 (N_1002,N_949,N_917);
nor U1003 (N_1003,N_943,N_952);
nand U1004 (N_1004,N_931,N_904);
nor U1005 (N_1005,N_957,N_972);
nand U1006 (N_1006,N_969,N_920);
and U1007 (N_1007,N_945,N_901);
nand U1008 (N_1008,N_915,N_903);
or U1009 (N_1009,N_925,N_973);
nand U1010 (N_1010,N_999,N_916);
nor U1011 (N_1011,N_998,N_935);
nor U1012 (N_1012,N_909,N_960);
nor U1013 (N_1013,N_923,N_974);
nand U1014 (N_1014,N_968,N_911);
or U1015 (N_1015,N_985,N_979);
xnor U1016 (N_1016,N_933,N_956);
and U1017 (N_1017,N_992,N_994);
nand U1018 (N_1018,N_918,N_988);
nand U1019 (N_1019,N_930,N_947);
nor U1020 (N_1020,N_981,N_982);
and U1021 (N_1021,N_983,N_993);
nor U1022 (N_1022,N_914,N_936);
and U1023 (N_1023,N_921,N_951);
or U1024 (N_1024,N_906,N_941);
or U1025 (N_1025,N_959,N_964);
and U1026 (N_1026,N_978,N_996);
nor U1027 (N_1027,N_902,N_970);
nor U1028 (N_1028,N_984,N_962);
or U1029 (N_1029,N_910,N_991);
nor U1030 (N_1030,N_966,N_975);
nor U1031 (N_1031,N_928,N_905);
and U1032 (N_1032,N_944,N_940);
nor U1033 (N_1033,N_927,N_977);
or U1034 (N_1034,N_958,N_997);
xor U1035 (N_1035,N_990,N_961);
nand U1036 (N_1036,N_912,N_976);
nand U1037 (N_1037,N_922,N_900);
nand U1038 (N_1038,N_919,N_980);
or U1039 (N_1039,N_924,N_953);
or U1040 (N_1040,N_986,N_934);
nand U1041 (N_1041,N_965,N_987);
nand U1042 (N_1042,N_954,N_938);
xnor U1043 (N_1043,N_908,N_995);
nand U1044 (N_1044,N_948,N_913);
and U1045 (N_1045,N_939,N_971);
nand U1046 (N_1046,N_907,N_932);
or U1047 (N_1047,N_942,N_929);
nand U1048 (N_1048,N_967,N_926);
nand U1049 (N_1049,N_955,N_963);
nand U1050 (N_1050,N_907,N_908);
or U1051 (N_1051,N_967,N_973);
nor U1052 (N_1052,N_912,N_941);
xor U1053 (N_1053,N_945,N_940);
and U1054 (N_1054,N_979,N_984);
or U1055 (N_1055,N_917,N_901);
and U1056 (N_1056,N_947,N_994);
nor U1057 (N_1057,N_989,N_944);
or U1058 (N_1058,N_927,N_904);
nor U1059 (N_1059,N_978,N_981);
nor U1060 (N_1060,N_910,N_977);
or U1061 (N_1061,N_919,N_950);
nand U1062 (N_1062,N_995,N_945);
nor U1063 (N_1063,N_983,N_960);
nor U1064 (N_1064,N_957,N_965);
and U1065 (N_1065,N_959,N_906);
and U1066 (N_1066,N_974,N_917);
nand U1067 (N_1067,N_947,N_924);
nor U1068 (N_1068,N_980,N_963);
and U1069 (N_1069,N_913,N_976);
nor U1070 (N_1070,N_974,N_922);
nor U1071 (N_1071,N_946,N_981);
nor U1072 (N_1072,N_946,N_968);
nor U1073 (N_1073,N_937,N_927);
nor U1074 (N_1074,N_943,N_991);
and U1075 (N_1075,N_929,N_915);
and U1076 (N_1076,N_966,N_934);
nor U1077 (N_1077,N_933,N_984);
and U1078 (N_1078,N_940,N_914);
nor U1079 (N_1079,N_951,N_900);
nor U1080 (N_1080,N_990,N_954);
or U1081 (N_1081,N_945,N_904);
nand U1082 (N_1082,N_981,N_910);
or U1083 (N_1083,N_996,N_908);
nor U1084 (N_1084,N_995,N_931);
and U1085 (N_1085,N_935,N_989);
and U1086 (N_1086,N_935,N_985);
or U1087 (N_1087,N_960,N_993);
nor U1088 (N_1088,N_982,N_901);
nor U1089 (N_1089,N_931,N_900);
nand U1090 (N_1090,N_958,N_929);
or U1091 (N_1091,N_991,N_949);
nor U1092 (N_1092,N_983,N_906);
nand U1093 (N_1093,N_915,N_995);
and U1094 (N_1094,N_914,N_918);
and U1095 (N_1095,N_928,N_911);
nor U1096 (N_1096,N_975,N_916);
or U1097 (N_1097,N_914,N_974);
and U1098 (N_1098,N_918,N_987);
and U1099 (N_1099,N_939,N_907);
nand U1100 (N_1100,N_1041,N_1031);
and U1101 (N_1101,N_1016,N_1065);
and U1102 (N_1102,N_1023,N_1027);
or U1103 (N_1103,N_1095,N_1060);
or U1104 (N_1104,N_1034,N_1052);
and U1105 (N_1105,N_1040,N_1096);
nor U1106 (N_1106,N_1067,N_1097);
nor U1107 (N_1107,N_1066,N_1091);
nor U1108 (N_1108,N_1071,N_1010);
or U1109 (N_1109,N_1053,N_1044);
nand U1110 (N_1110,N_1004,N_1050);
or U1111 (N_1111,N_1076,N_1056);
or U1112 (N_1112,N_1001,N_1089);
or U1113 (N_1113,N_1064,N_1025);
and U1114 (N_1114,N_1092,N_1014);
or U1115 (N_1115,N_1030,N_1000);
nand U1116 (N_1116,N_1009,N_1012);
or U1117 (N_1117,N_1055,N_1072);
and U1118 (N_1118,N_1046,N_1094);
nor U1119 (N_1119,N_1007,N_1058);
or U1120 (N_1120,N_1086,N_1070);
nand U1121 (N_1121,N_1051,N_1083);
and U1122 (N_1122,N_1022,N_1063);
and U1123 (N_1123,N_1013,N_1049);
nand U1124 (N_1124,N_1087,N_1045);
nand U1125 (N_1125,N_1098,N_1077);
or U1126 (N_1126,N_1028,N_1061);
nand U1127 (N_1127,N_1036,N_1069);
nand U1128 (N_1128,N_1018,N_1024);
nand U1129 (N_1129,N_1059,N_1084);
nor U1130 (N_1130,N_1021,N_1035);
nor U1131 (N_1131,N_1090,N_1075);
or U1132 (N_1132,N_1099,N_1048);
nand U1133 (N_1133,N_1073,N_1029);
and U1134 (N_1134,N_1082,N_1088);
nand U1135 (N_1135,N_1037,N_1057);
or U1136 (N_1136,N_1006,N_1068);
nor U1137 (N_1137,N_1042,N_1080);
and U1138 (N_1138,N_1011,N_1062);
and U1139 (N_1139,N_1032,N_1093);
and U1140 (N_1140,N_1026,N_1039);
nor U1141 (N_1141,N_1043,N_1005);
or U1142 (N_1142,N_1074,N_1079);
nor U1143 (N_1143,N_1081,N_1002);
nand U1144 (N_1144,N_1038,N_1078);
nand U1145 (N_1145,N_1047,N_1019);
nor U1146 (N_1146,N_1008,N_1017);
nor U1147 (N_1147,N_1033,N_1020);
and U1148 (N_1148,N_1054,N_1003);
nor U1149 (N_1149,N_1085,N_1015);
or U1150 (N_1150,N_1019,N_1074);
or U1151 (N_1151,N_1008,N_1029);
and U1152 (N_1152,N_1095,N_1076);
or U1153 (N_1153,N_1087,N_1091);
and U1154 (N_1154,N_1002,N_1028);
xnor U1155 (N_1155,N_1003,N_1032);
xor U1156 (N_1156,N_1003,N_1023);
and U1157 (N_1157,N_1014,N_1097);
nand U1158 (N_1158,N_1008,N_1087);
nor U1159 (N_1159,N_1014,N_1083);
or U1160 (N_1160,N_1042,N_1064);
nor U1161 (N_1161,N_1037,N_1080);
nor U1162 (N_1162,N_1078,N_1042);
nand U1163 (N_1163,N_1073,N_1036);
and U1164 (N_1164,N_1014,N_1026);
or U1165 (N_1165,N_1008,N_1033);
nand U1166 (N_1166,N_1019,N_1092);
and U1167 (N_1167,N_1086,N_1002);
and U1168 (N_1168,N_1033,N_1001);
or U1169 (N_1169,N_1045,N_1060);
and U1170 (N_1170,N_1054,N_1060);
nor U1171 (N_1171,N_1065,N_1019);
and U1172 (N_1172,N_1005,N_1034);
and U1173 (N_1173,N_1064,N_1072);
and U1174 (N_1174,N_1092,N_1017);
or U1175 (N_1175,N_1065,N_1087);
and U1176 (N_1176,N_1082,N_1084);
or U1177 (N_1177,N_1024,N_1072);
nand U1178 (N_1178,N_1082,N_1093);
and U1179 (N_1179,N_1024,N_1048);
nor U1180 (N_1180,N_1091,N_1057);
nor U1181 (N_1181,N_1060,N_1055);
nand U1182 (N_1182,N_1001,N_1053);
nand U1183 (N_1183,N_1027,N_1063);
nand U1184 (N_1184,N_1021,N_1013);
and U1185 (N_1185,N_1068,N_1036);
nand U1186 (N_1186,N_1010,N_1098);
nand U1187 (N_1187,N_1092,N_1078);
nand U1188 (N_1188,N_1038,N_1041);
nand U1189 (N_1189,N_1013,N_1020);
or U1190 (N_1190,N_1087,N_1011);
or U1191 (N_1191,N_1093,N_1039);
and U1192 (N_1192,N_1029,N_1063);
nand U1193 (N_1193,N_1035,N_1023);
nand U1194 (N_1194,N_1025,N_1049);
nor U1195 (N_1195,N_1063,N_1033);
and U1196 (N_1196,N_1053,N_1028);
nor U1197 (N_1197,N_1046,N_1044);
and U1198 (N_1198,N_1067,N_1026);
nand U1199 (N_1199,N_1093,N_1001);
nor U1200 (N_1200,N_1194,N_1134);
nor U1201 (N_1201,N_1150,N_1117);
nand U1202 (N_1202,N_1190,N_1159);
xor U1203 (N_1203,N_1115,N_1149);
and U1204 (N_1204,N_1163,N_1131);
and U1205 (N_1205,N_1124,N_1184);
or U1206 (N_1206,N_1181,N_1105);
nand U1207 (N_1207,N_1172,N_1161);
nand U1208 (N_1208,N_1145,N_1192);
and U1209 (N_1209,N_1114,N_1162);
or U1210 (N_1210,N_1195,N_1197);
nand U1211 (N_1211,N_1170,N_1173);
nor U1212 (N_1212,N_1169,N_1136);
and U1213 (N_1213,N_1121,N_1156);
nor U1214 (N_1214,N_1113,N_1189);
or U1215 (N_1215,N_1130,N_1157);
nand U1216 (N_1216,N_1140,N_1106);
nand U1217 (N_1217,N_1100,N_1144);
nor U1218 (N_1218,N_1142,N_1186);
and U1219 (N_1219,N_1177,N_1110);
nor U1220 (N_1220,N_1178,N_1135);
xnor U1221 (N_1221,N_1122,N_1152);
or U1222 (N_1222,N_1193,N_1132);
nand U1223 (N_1223,N_1179,N_1166);
or U1224 (N_1224,N_1176,N_1183);
nor U1225 (N_1225,N_1147,N_1168);
nand U1226 (N_1226,N_1167,N_1141);
nor U1227 (N_1227,N_1127,N_1111);
nor U1228 (N_1228,N_1187,N_1188);
nor U1229 (N_1229,N_1175,N_1155);
xor U1230 (N_1230,N_1138,N_1120);
nand U1231 (N_1231,N_1185,N_1102);
nand U1232 (N_1232,N_1101,N_1108);
and U1233 (N_1233,N_1139,N_1182);
nor U1234 (N_1234,N_1196,N_1104);
or U1235 (N_1235,N_1112,N_1109);
and U1236 (N_1236,N_1123,N_1107);
or U1237 (N_1237,N_1133,N_1154);
or U1238 (N_1238,N_1153,N_1146);
and U1239 (N_1239,N_1128,N_1148);
nor U1240 (N_1240,N_1180,N_1116);
nand U1241 (N_1241,N_1198,N_1199);
and U1242 (N_1242,N_1174,N_1160);
nor U1243 (N_1243,N_1164,N_1191);
nor U1244 (N_1244,N_1129,N_1118);
nor U1245 (N_1245,N_1126,N_1103);
and U1246 (N_1246,N_1171,N_1119);
or U1247 (N_1247,N_1143,N_1151);
or U1248 (N_1248,N_1137,N_1158);
and U1249 (N_1249,N_1165,N_1125);
nand U1250 (N_1250,N_1140,N_1168);
nand U1251 (N_1251,N_1167,N_1194);
and U1252 (N_1252,N_1191,N_1131);
nand U1253 (N_1253,N_1120,N_1163);
or U1254 (N_1254,N_1109,N_1150);
nor U1255 (N_1255,N_1193,N_1156);
nand U1256 (N_1256,N_1177,N_1180);
or U1257 (N_1257,N_1127,N_1195);
nor U1258 (N_1258,N_1125,N_1162);
or U1259 (N_1259,N_1139,N_1116);
nand U1260 (N_1260,N_1107,N_1195);
nor U1261 (N_1261,N_1181,N_1153);
and U1262 (N_1262,N_1123,N_1118);
nor U1263 (N_1263,N_1171,N_1109);
or U1264 (N_1264,N_1147,N_1131);
or U1265 (N_1265,N_1186,N_1166);
and U1266 (N_1266,N_1170,N_1123);
and U1267 (N_1267,N_1120,N_1116);
nand U1268 (N_1268,N_1127,N_1115);
xor U1269 (N_1269,N_1114,N_1158);
xnor U1270 (N_1270,N_1171,N_1108);
and U1271 (N_1271,N_1193,N_1125);
nand U1272 (N_1272,N_1106,N_1109);
nor U1273 (N_1273,N_1161,N_1157);
nor U1274 (N_1274,N_1165,N_1157);
nand U1275 (N_1275,N_1133,N_1123);
nand U1276 (N_1276,N_1144,N_1110);
nand U1277 (N_1277,N_1160,N_1156);
and U1278 (N_1278,N_1159,N_1151);
or U1279 (N_1279,N_1129,N_1115);
nor U1280 (N_1280,N_1116,N_1187);
and U1281 (N_1281,N_1177,N_1144);
and U1282 (N_1282,N_1138,N_1141);
or U1283 (N_1283,N_1181,N_1177);
nand U1284 (N_1284,N_1127,N_1126);
or U1285 (N_1285,N_1157,N_1199);
nand U1286 (N_1286,N_1179,N_1103);
nor U1287 (N_1287,N_1152,N_1131);
xor U1288 (N_1288,N_1107,N_1140);
and U1289 (N_1289,N_1168,N_1104);
nor U1290 (N_1290,N_1188,N_1144);
and U1291 (N_1291,N_1102,N_1133);
and U1292 (N_1292,N_1140,N_1119);
nand U1293 (N_1293,N_1127,N_1169);
and U1294 (N_1294,N_1166,N_1187);
or U1295 (N_1295,N_1139,N_1174);
and U1296 (N_1296,N_1104,N_1130);
nor U1297 (N_1297,N_1123,N_1161);
and U1298 (N_1298,N_1111,N_1156);
nand U1299 (N_1299,N_1161,N_1142);
and U1300 (N_1300,N_1250,N_1294);
or U1301 (N_1301,N_1223,N_1241);
or U1302 (N_1302,N_1225,N_1236);
nor U1303 (N_1303,N_1292,N_1287);
nand U1304 (N_1304,N_1217,N_1263);
and U1305 (N_1305,N_1286,N_1260);
nor U1306 (N_1306,N_1298,N_1226);
and U1307 (N_1307,N_1230,N_1216);
and U1308 (N_1308,N_1276,N_1239);
and U1309 (N_1309,N_1272,N_1243);
and U1310 (N_1310,N_1252,N_1227);
or U1311 (N_1311,N_1270,N_1211);
xor U1312 (N_1312,N_1273,N_1283);
nor U1313 (N_1313,N_1258,N_1234);
or U1314 (N_1314,N_1289,N_1207);
nor U1315 (N_1315,N_1251,N_1267);
nor U1316 (N_1316,N_1209,N_1215);
nor U1317 (N_1317,N_1229,N_1256);
nand U1318 (N_1318,N_1237,N_1271);
nand U1319 (N_1319,N_1268,N_1224);
xor U1320 (N_1320,N_1240,N_1214);
and U1321 (N_1321,N_1293,N_1245);
nand U1322 (N_1322,N_1202,N_1206);
and U1323 (N_1323,N_1259,N_1295);
nor U1324 (N_1324,N_1218,N_1242);
and U1325 (N_1325,N_1232,N_1281);
or U1326 (N_1326,N_1269,N_1220);
and U1327 (N_1327,N_1222,N_1253);
xor U1328 (N_1328,N_1282,N_1262);
and U1329 (N_1329,N_1201,N_1291);
nand U1330 (N_1330,N_1257,N_1265);
and U1331 (N_1331,N_1244,N_1228);
or U1332 (N_1332,N_1279,N_1285);
nand U1333 (N_1333,N_1284,N_1219);
nand U1334 (N_1334,N_1212,N_1297);
nor U1335 (N_1335,N_1247,N_1213);
nand U1336 (N_1336,N_1254,N_1233);
and U1337 (N_1337,N_1278,N_1288);
or U1338 (N_1338,N_1296,N_1204);
nand U1339 (N_1339,N_1274,N_1249);
and U1340 (N_1340,N_1299,N_1200);
or U1341 (N_1341,N_1290,N_1235);
or U1342 (N_1342,N_1264,N_1208);
nand U1343 (N_1343,N_1246,N_1280);
and U1344 (N_1344,N_1261,N_1248);
or U1345 (N_1345,N_1221,N_1238);
nor U1346 (N_1346,N_1275,N_1231);
and U1347 (N_1347,N_1266,N_1277);
and U1348 (N_1348,N_1210,N_1203);
and U1349 (N_1349,N_1255,N_1205);
nor U1350 (N_1350,N_1248,N_1252);
nand U1351 (N_1351,N_1275,N_1251);
or U1352 (N_1352,N_1201,N_1219);
nor U1353 (N_1353,N_1201,N_1256);
nand U1354 (N_1354,N_1280,N_1271);
nor U1355 (N_1355,N_1229,N_1263);
nand U1356 (N_1356,N_1207,N_1262);
or U1357 (N_1357,N_1231,N_1207);
nor U1358 (N_1358,N_1286,N_1216);
nor U1359 (N_1359,N_1246,N_1222);
nor U1360 (N_1360,N_1233,N_1280);
and U1361 (N_1361,N_1255,N_1267);
nor U1362 (N_1362,N_1298,N_1272);
nand U1363 (N_1363,N_1260,N_1274);
and U1364 (N_1364,N_1244,N_1233);
or U1365 (N_1365,N_1279,N_1271);
nor U1366 (N_1366,N_1287,N_1255);
nor U1367 (N_1367,N_1287,N_1282);
nand U1368 (N_1368,N_1275,N_1210);
nor U1369 (N_1369,N_1206,N_1282);
nand U1370 (N_1370,N_1232,N_1259);
or U1371 (N_1371,N_1253,N_1275);
nand U1372 (N_1372,N_1268,N_1216);
and U1373 (N_1373,N_1238,N_1219);
or U1374 (N_1374,N_1222,N_1293);
or U1375 (N_1375,N_1211,N_1255);
or U1376 (N_1376,N_1231,N_1253);
nand U1377 (N_1377,N_1251,N_1265);
nor U1378 (N_1378,N_1292,N_1260);
and U1379 (N_1379,N_1221,N_1264);
nand U1380 (N_1380,N_1209,N_1281);
nor U1381 (N_1381,N_1295,N_1265);
nor U1382 (N_1382,N_1255,N_1285);
and U1383 (N_1383,N_1270,N_1218);
nand U1384 (N_1384,N_1248,N_1256);
and U1385 (N_1385,N_1283,N_1220);
and U1386 (N_1386,N_1266,N_1236);
nor U1387 (N_1387,N_1235,N_1285);
or U1388 (N_1388,N_1226,N_1204);
nand U1389 (N_1389,N_1222,N_1203);
and U1390 (N_1390,N_1289,N_1252);
and U1391 (N_1391,N_1219,N_1294);
and U1392 (N_1392,N_1259,N_1247);
and U1393 (N_1393,N_1259,N_1272);
and U1394 (N_1394,N_1298,N_1284);
and U1395 (N_1395,N_1226,N_1282);
nand U1396 (N_1396,N_1284,N_1271);
and U1397 (N_1397,N_1272,N_1220);
or U1398 (N_1398,N_1218,N_1284);
nand U1399 (N_1399,N_1260,N_1279);
xnor U1400 (N_1400,N_1364,N_1392);
nor U1401 (N_1401,N_1331,N_1341);
xnor U1402 (N_1402,N_1356,N_1375);
nand U1403 (N_1403,N_1393,N_1355);
or U1404 (N_1404,N_1316,N_1318);
or U1405 (N_1405,N_1329,N_1388);
and U1406 (N_1406,N_1308,N_1303);
and U1407 (N_1407,N_1377,N_1300);
xnor U1408 (N_1408,N_1362,N_1322);
nor U1409 (N_1409,N_1335,N_1357);
nor U1410 (N_1410,N_1383,N_1307);
and U1411 (N_1411,N_1397,N_1321);
nand U1412 (N_1412,N_1344,N_1311);
nand U1413 (N_1413,N_1302,N_1326);
nand U1414 (N_1414,N_1309,N_1334);
or U1415 (N_1415,N_1354,N_1378);
nand U1416 (N_1416,N_1337,N_1312);
nor U1417 (N_1417,N_1340,N_1310);
nand U1418 (N_1418,N_1374,N_1305);
or U1419 (N_1419,N_1315,N_1313);
nor U1420 (N_1420,N_1361,N_1359);
nor U1421 (N_1421,N_1330,N_1304);
nand U1422 (N_1422,N_1347,N_1346);
and U1423 (N_1423,N_1306,N_1390);
nor U1424 (N_1424,N_1399,N_1332);
and U1425 (N_1425,N_1342,N_1301);
nand U1426 (N_1426,N_1398,N_1319);
nor U1427 (N_1427,N_1353,N_1387);
nor U1428 (N_1428,N_1373,N_1360);
and U1429 (N_1429,N_1369,N_1317);
nand U1430 (N_1430,N_1395,N_1386);
and U1431 (N_1431,N_1382,N_1320);
or U1432 (N_1432,N_1384,N_1367);
and U1433 (N_1433,N_1339,N_1336);
and U1434 (N_1434,N_1325,N_1372);
nand U1435 (N_1435,N_1363,N_1371);
xnor U1436 (N_1436,N_1314,N_1391);
nor U1437 (N_1437,N_1396,N_1385);
or U1438 (N_1438,N_1389,N_1338);
and U1439 (N_1439,N_1352,N_1376);
nand U1440 (N_1440,N_1343,N_1370);
and U1441 (N_1441,N_1328,N_1368);
and U1442 (N_1442,N_1324,N_1327);
or U1443 (N_1443,N_1365,N_1345);
nand U1444 (N_1444,N_1379,N_1351);
nand U1445 (N_1445,N_1333,N_1348);
nand U1446 (N_1446,N_1380,N_1358);
or U1447 (N_1447,N_1366,N_1350);
and U1448 (N_1448,N_1381,N_1394);
nand U1449 (N_1449,N_1349,N_1323);
nand U1450 (N_1450,N_1358,N_1396);
nand U1451 (N_1451,N_1317,N_1316);
and U1452 (N_1452,N_1377,N_1334);
nor U1453 (N_1453,N_1339,N_1398);
or U1454 (N_1454,N_1372,N_1303);
nor U1455 (N_1455,N_1389,N_1309);
and U1456 (N_1456,N_1349,N_1329);
nand U1457 (N_1457,N_1346,N_1322);
and U1458 (N_1458,N_1343,N_1303);
or U1459 (N_1459,N_1319,N_1371);
or U1460 (N_1460,N_1398,N_1385);
or U1461 (N_1461,N_1379,N_1307);
nor U1462 (N_1462,N_1340,N_1352);
nand U1463 (N_1463,N_1349,N_1339);
nor U1464 (N_1464,N_1348,N_1341);
or U1465 (N_1465,N_1309,N_1332);
nor U1466 (N_1466,N_1390,N_1336);
nor U1467 (N_1467,N_1323,N_1315);
nand U1468 (N_1468,N_1334,N_1359);
nand U1469 (N_1469,N_1316,N_1345);
or U1470 (N_1470,N_1324,N_1300);
and U1471 (N_1471,N_1327,N_1337);
nand U1472 (N_1472,N_1393,N_1359);
or U1473 (N_1473,N_1364,N_1389);
nand U1474 (N_1474,N_1346,N_1315);
nand U1475 (N_1475,N_1310,N_1307);
nand U1476 (N_1476,N_1349,N_1388);
and U1477 (N_1477,N_1362,N_1391);
nand U1478 (N_1478,N_1332,N_1398);
and U1479 (N_1479,N_1399,N_1378);
or U1480 (N_1480,N_1386,N_1325);
or U1481 (N_1481,N_1399,N_1304);
nor U1482 (N_1482,N_1375,N_1303);
xnor U1483 (N_1483,N_1318,N_1315);
nand U1484 (N_1484,N_1323,N_1356);
nand U1485 (N_1485,N_1391,N_1346);
xnor U1486 (N_1486,N_1332,N_1393);
nor U1487 (N_1487,N_1397,N_1363);
nor U1488 (N_1488,N_1345,N_1379);
and U1489 (N_1489,N_1385,N_1334);
nand U1490 (N_1490,N_1387,N_1384);
and U1491 (N_1491,N_1374,N_1397);
and U1492 (N_1492,N_1319,N_1334);
and U1493 (N_1493,N_1326,N_1375);
and U1494 (N_1494,N_1377,N_1368);
nand U1495 (N_1495,N_1368,N_1336);
nor U1496 (N_1496,N_1376,N_1397);
and U1497 (N_1497,N_1324,N_1312);
nor U1498 (N_1498,N_1325,N_1352);
nand U1499 (N_1499,N_1341,N_1329);
nand U1500 (N_1500,N_1434,N_1437);
or U1501 (N_1501,N_1421,N_1435);
xor U1502 (N_1502,N_1476,N_1444);
nor U1503 (N_1503,N_1409,N_1432);
or U1504 (N_1504,N_1477,N_1469);
nand U1505 (N_1505,N_1486,N_1443);
nand U1506 (N_1506,N_1447,N_1403);
and U1507 (N_1507,N_1489,N_1466);
nor U1508 (N_1508,N_1484,N_1474);
nor U1509 (N_1509,N_1406,N_1415);
nand U1510 (N_1510,N_1423,N_1450);
or U1511 (N_1511,N_1488,N_1426);
xor U1512 (N_1512,N_1433,N_1405);
nand U1513 (N_1513,N_1408,N_1494);
nand U1514 (N_1514,N_1479,N_1496);
or U1515 (N_1515,N_1468,N_1464);
and U1516 (N_1516,N_1430,N_1429);
nor U1517 (N_1517,N_1472,N_1411);
and U1518 (N_1518,N_1407,N_1445);
nor U1519 (N_1519,N_1438,N_1401);
and U1520 (N_1520,N_1442,N_1424);
and U1521 (N_1521,N_1451,N_1465);
or U1522 (N_1522,N_1473,N_1498);
or U1523 (N_1523,N_1417,N_1495);
nand U1524 (N_1524,N_1436,N_1418);
nor U1525 (N_1525,N_1493,N_1462);
and U1526 (N_1526,N_1457,N_1459);
or U1527 (N_1527,N_1499,N_1454);
nand U1528 (N_1528,N_1414,N_1425);
nor U1529 (N_1529,N_1467,N_1458);
nand U1530 (N_1530,N_1448,N_1490);
and U1531 (N_1531,N_1419,N_1481);
and U1532 (N_1532,N_1400,N_1420);
or U1533 (N_1533,N_1410,N_1453);
nand U1534 (N_1534,N_1485,N_1404);
and U1535 (N_1535,N_1455,N_1446);
nand U1536 (N_1536,N_1412,N_1492);
nor U1537 (N_1537,N_1416,N_1471);
or U1538 (N_1538,N_1497,N_1456);
nor U1539 (N_1539,N_1431,N_1478);
nor U1540 (N_1540,N_1470,N_1452);
xnor U1541 (N_1541,N_1413,N_1428);
or U1542 (N_1542,N_1480,N_1449);
nor U1543 (N_1543,N_1402,N_1475);
nor U1544 (N_1544,N_1440,N_1483);
nor U1545 (N_1545,N_1422,N_1439);
or U1546 (N_1546,N_1463,N_1427);
and U1547 (N_1547,N_1441,N_1482);
or U1548 (N_1548,N_1460,N_1487);
and U1549 (N_1549,N_1461,N_1491);
and U1550 (N_1550,N_1412,N_1455);
or U1551 (N_1551,N_1488,N_1405);
or U1552 (N_1552,N_1424,N_1410);
nand U1553 (N_1553,N_1465,N_1490);
and U1554 (N_1554,N_1407,N_1430);
and U1555 (N_1555,N_1413,N_1436);
or U1556 (N_1556,N_1456,N_1401);
or U1557 (N_1557,N_1439,N_1460);
nor U1558 (N_1558,N_1465,N_1433);
nand U1559 (N_1559,N_1483,N_1474);
or U1560 (N_1560,N_1468,N_1444);
and U1561 (N_1561,N_1440,N_1443);
nor U1562 (N_1562,N_1448,N_1410);
or U1563 (N_1563,N_1469,N_1408);
nand U1564 (N_1564,N_1437,N_1411);
or U1565 (N_1565,N_1439,N_1493);
and U1566 (N_1566,N_1498,N_1461);
nor U1567 (N_1567,N_1421,N_1413);
or U1568 (N_1568,N_1423,N_1433);
and U1569 (N_1569,N_1490,N_1463);
nor U1570 (N_1570,N_1420,N_1498);
or U1571 (N_1571,N_1478,N_1402);
or U1572 (N_1572,N_1446,N_1478);
nor U1573 (N_1573,N_1426,N_1427);
nor U1574 (N_1574,N_1485,N_1470);
nand U1575 (N_1575,N_1498,N_1486);
nor U1576 (N_1576,N_1493,N_1495);
nor U1577 (N_1577,N_1465,N_1408);
nand U1578 (N_1578,N_1420,N_1478);
nor U1579 (N_1579,N_1474,N_1401);
or U1580 (N_1580,N_1437,N_1401);
nand U1581 (N_1581,N_1464,N_1409);
nor U1582 (N_1582,N_1432,N_1408);
or U1583 (N_1583,N_1427,N_1476);
nand U1584 (N_1584,N_1445,N_1444);
nor U1585 (N_1585,N_1492,N_1429);
or U1586 (N_1586,N_1413,N_1456);
nor U1587 (N_1587,N_1437,N_1441);
nor U1588 (N_1588,N_1479,N_1408);
nor U1589 (N_1589,N_1444,N_1481);
nor U1590 (N_1590,N_1447,N_1471);
and U1591 (N_1591,N_1473,N_1497);
nand U1592 (N_1592,N_1491,N_1438);
or U1593 (N_1593,N_1463,N_1493);
and U1594 (N_1594,N_1429,N_1481);
nand U1595 (N_1595,N_1450,N_1491);
and U1596 (N_1596,N_1432,N_1436);
and U1597 (N_1597,N_1448,N_1498);
nor U1598 (N_1598,N_1441,N_1415);
nor U1599 (N_1599,N_1471,N_1444);
and U1600 (N_1600,N_1591,N_1506);
or U1601 (N_1601,N_1585,N_1507);
nand U1602 (N_1602,N_1570,N_1594);
and U1603 (N_1603,N_1511,N_1552);
nor U1604 (N_1604,N_1522,N_1572);
and U1605 (N_1605,N_1538,N_1525);
and U1606 (N_1606,N_1505,N_1542);
and U1607 (N_1607,N_1564,N_1504);
and U1608 (N_1608,N_1568,N_1547);
nor U1609 (N_1609,N_1571,N_1579);
nor U1610 (N_1610,N_1595,N_1502);
nand U1611 (N_1611,N_1598,N_1597);
or U1612 (N_1612,N_1589,N_1532);
nand U1613 (N_1613,N_1583,N_1510);
and U1614 (N_1614,N_1576,N_1562);
nand U1615 (N_1615,N_1582,N_1531);
nand U1616 (N_1616,N_1596,N_1586);
and U1617 (N_1617,N_1527,N_1563);
and U1618 (N_1618,N_1518,N_1556);
or U1619 (N_1619,N_1534,N_1578);
nand U1620 (N_1620,N_1577,N_1548);
or U1621 (N_1621,N_1539,N_1573);
or U1622 (N_1622,N_1560,N_1565);
or U1623 (N_1623,N_1509,N_1537);
and U1624 (N_1624,N_1544,N_1584);
nand U1625 (N_1625,N_1540,N_1517);
nand U1626 (N_1626,N_1557,N_1528);
nand U1627 (N_1627,N_1574,N_1566);
and U1628 (N_1628,N_1529,N_1575);
or U1629 (N_1629,N_1545,N_1561);
nand U1630 (N_1630,N_1558,N_1519);
and U1631 (N_1631,N_1555,N_1536);
nand U1632 (N_1632,N_1567,N_1503);
nor U1633 (N_1633,N_1515,N_1530);
nor U1634 (N_1634,N_1513,N_1559);
nand U1635 (N_1635,N_1599,N_1535);
xnor U1636 (N_1636,N_1581,N_1541);
nor U1637 (N_1637,N_1512,N_1592);
nand U1638 (N_1638,N_1533,N_1587);
and U1639 (N_1639,N_1569,N_1520);
nand U1640 (N_1640,N_1546,N_1580);
nor U1641 (N_1641,N_1550,N_1514);
and U1642 (N_1642,N_1590,N_1516);
nor U1643 (N_1643,N_1593,N_1551);
and U1644 (N_1644,N_1543,N_1549);
nand U1645 (N_1645,N_1523,N_1526);
nor U1646 (N_1646,N_1521,N_1524);
nor U1647 (N_1647,N_1500,N_1508);
or U1648 (N_1648,N_1588,N_1501);
nor U1649 (N_1649,N_1553,N_1554);
nor U1650 (N_1650,N_1580,N_1579);
nand U1651 (N_1651,N_1558,N_1565);
or U1652 (N_1652,N_1554,N_1549);
nand U1653 (N_1653,N_1515,N_1518);
nor U1654 (N_1654,N_1556,N_1560);
nor U1655 (N_1655,N_1577,N_1545);
nor U1656 (N_1656,N_1543,N_1560);
nor U1657 (N_1657,N_1568,N_1566);
and U1658 (N_1658,N_1572,N_1506);
nor U1659 (N_1659,N_1575,N_1570);
nor U1660 (N_1660,N_1535,N_1566);
nor U1661 (N_1661,N_1543,N_1551);
or U1662 (N_1662,N_1517,N_1582);
and U1663 (N_1663,N_1547,N_1535);
or U1664 (N_1664,N_1519,N_1553);
nor U1665 (N_1665,N_1594,N_1581);
nor U1666 (N_1666,N_1558,N_1597);
nand U1667 (N_1667,N_1561,N_1543);
nor U1668 (N_1668,N_1512,N_1554);
and U1669 (N_1669,N_1555,N_1565);
nor U1670 (N_1670,N_1587,N_1541);
nor U1671 (N_1671,N_1502,N_1546);
and U1672 (N_1672,N_1583,N_1538);
nor U1673 (N_1673,N_1531,N_1506);
or U1674 (N_1674,N_1598,N_1523);
nand U1675 (N_1675,N_1585,N_1594);
and U1676 (N_1676,N_1525,N_1534);
xnor U1677 (N_1677,N_1561,N_1578);
nand U1678 (N_1678,N_1547,N_1593);
nor U1679 (N_1679,N_1597,N_1535);
and U1680 (N_1680,N_1548,N_1581);
and U1681 (N_1681,N_1594,N_1586);
or U1682 (N_1682,N_1529,N_1560);
and U1683 (N_1683,N_1541,N_1504);
or U1684 (N_1684,N_1577,N_1501);
or U1685 (N_1685,N_1534,N_1579);
nand U1686 (N_1686,N_1561,N_1515);
or U1687 (N_1687,N_1571,N_1521);
nand U1688 (N_1688,N_1547,N_1521);
nor U1689 (N_1689,N_1595,N_1556);
or U1690 (N_1690,N_1543,N_1584);
and U1691 (N_1691,N_1557,N_1565);
and U1692 (N_1692,N_1538,N_1550);
nor U1693 (N_1693,N_1513,N_1568);
and U1694 (N_1694,N_1597,N_1538);
nor U1695 (N_1695,N_1537,N_1589);
nor U1696 (N_1696,N_1544,N_1543);
nor U1697 (N_1697,N_1575,N_1510);
and U1698 (N_1698,N_1557,N_1554);
or U1699 (N_1699,N_1558,N_1595);
and U1700 (N_1700,N_1614,N_1605);
nor U1701 (N_1701,N_1649,N_1657);
or U1702 (N_1702,N_1618,N_1678);
nor U1703 (N_1703,N_1646,N_1694);
and U1704 (N_1704,N_1693,N_1659);
nand U1705 (N_1705,N_1683,N_1630);
and U1706 (N_1706,N_1635,N_1661);
nand U1707 (N_1707,N_1611,N_1626);
nand U1708 (N_1708,N_1653,N_1603);
nand U1709 (N_1709,N_1695,N_1625);
nor U1710 (N_1710,N_1606,N_1602);
or U1711 (N_1711,N_1638,N_1623);
nor U1712 (N_1712,N_1664,N_1641);
xnor U1713 (N_1713,N_1655,N_1667);
and U1714 (N_1714,N_1662,N_1680);
and U1715 (N_1715,N_1676,N_1650);
and U1716 (N_1716,N_1697,N_1688);
or U1717 (N_1717,N_1698,N_1636);
and U1718 (N_1718,N_1612,N_1682);
or U1719 (N_1719,N_1633,N_1604);
nand U1720 (N_1720,N_1613,N_1687);
and U1721 (N_1721,N_1620,N_1608);
nor U1722 (N_1722,N_1645,N_1651);
nand U1723 (N_1723,N_1684,N_1666);
and U1724 (N_1724,N_1690,N_1677);
nand U1725 (N_1725,N_1663,N_1669);
or U1726 (N_1726,N_1654,N_1627);
nor U1727 (N_1727,N_1643,N_1692);
nand U1728 (N_1728,N_1672,N_1689);
or U1729 (N_1729,N_1648,N_1632);
and U1730 (N_1730,N_1622,N_1699);
or U1731 (N_1731,N_1607,N_1674);
or U1732 (N_1732,N_1665,N_1670);
nor U1733 (N_1733,N_1629,N_1656);
nand U1734 (N_1734,N_1609,N_1610);
nor U1735 (N_1735,N_1685,N_1671);
or U1736 (N_1736,N_1647,N_1652);
nor U1737 (N_1737,N_1634,N_1660);
or U1738 (N_1738,N_1600,N_1624);
nand U1739 (N_1739,N_1617,N_1675);
nor U1740 (N_1740,N_1637,N_1619);
and U1741 (N_1741,N_1640,N_1696);
or U1742 (N_1742,N_1668,N_1644);
nand U1743 (N_1743,N_1615,N_1658);
and U1744 (N_1744,N_1642,N_1631);
nor U1745 (N_1745,N_1621,N_1679);
or U1746 (N_1746,N_1681,N_1616);
and U1747 (N_1747,N_1639,N_1673);
or U1748 (N_1748,N_1628,N_1691);
and U1749 (N_1749,N_1601,N_1686);
nand U1750 (N_1750,N_1650,N_1690);
nor U1751 (N_1751,N_1639,N_1674);
or U1752 (N_1752,N_1606,N_1633);
or U1753 (N_1753,N_1649,N_1651);
and U1754 (N_1754,N_1660,N_1620);
nand U1755 (N_1755,N_1626,N_1650);
nor U1756 (N_1756,N_1633,N_1628);
nand U1757 (N_1757,N_1663,N_1602);
or U1758 (N_1758,N_1680,N_1638);
or U1759 (N_1759,N_1650,N_1663);
nand U1760 (N_1760,N_1643,N_1696);
nor U1761 (N_1761,N_1691,N_1687);
nor U1762 (N_1762,N_1663,N_1649);
and U1763 (N_1763,N_1658,N_1692);
xnor U1764 (N_1764,N_1601,N_1662);
nand U1765 (N_1765,N_1679,N_1640);
or U1766 (N_1766,N_1665,N_1679);
and U1767 (N_1767,N_1690,N_1664);
or U1768 (N_1768,N_1676,N_1602);
and U1769 (N_1769,N_1685,N_1674);
nand U1770 (N_1770,N_1693,N_1649);
and U1771 (N_1771,N_1683,N_1672);
or U1772 (N_1772,N_1617,N_1669);
nand U1773 (N_1773,N_1624,N_1604);
nor U1774 (N_1774,N_1658,N_1677);
or U1775 (N_1775,N_1669,N_1628);
and U1776 (N_1776,N_1668,N_1696);
nor U1777 (N_1777,N_1655,N_1670);
or U1778 (N_1778,N_1660,N_1631);
or U1779 (N_1779,N_1671,N_1647);
or U1780 (N_1780,N_1653,N_1642);
xnor U1781 (N_1781,N_1686,N_1630);
and U1782 (N_1782,N_1647,N_1681);
or U1783 (N_1783,N_1612,N_1656);
and U1784 (N_1784,N_1687,N_1650);
nor U1785 (N_1785,N_1676,N_1618);
and U1786 (N_1786,N_1603,N_1681);
and U1787 (N_1787,N_1693,N_1602);
and U1788 (N_1788,N_1612,N_1642);
or U1789 (N_1789,N_1603,N_1674);
or U1790 (N_1790,N_1677,N_1630);
and U1791 (N_1791,N_1689,N_1659);
nand U1792 (N_1792,N_1613,N_1611);
and U1793 (N_1793,N_1626,N_1683);
or U1794 (N_1794,N_1644,N_1678);
nor U1795 (N_1795,N_1604,N_1625);
nand U1796 (N_1796,N_1680,N_1657);
nor U1797 (N_1797,N_1655,N_1688);
or U1798 (N_1798,N_1645,N_1663);
or U1799 (N_1799,N_1691,N_1672);
or U1800 (N_1800,N_1724,N_1791);
nand U1801 (N_1801,N_1787,N_1736);
nor U1802 (N_1802,N_1797,N_1762);
nor U1803 (N_1803,N_1709,N_1730);
nor U1804 (N_1804,N_1749,N_1788);
nand U1805 (N_1805,N_1772,N_1731);
and U1806 (N_1806,N_1777,N_1739);
nand U1807 (N_1807,N_1715,N_1775);
nand U1808 (N_1808,N_1751,N_1750);
and U1809 (N_1809,N_1774,N_1794);
or U1810 (N_1810,N_1726,N_1785);
nand U1811 (N_1811,N_1767,N_1765);
or U1812 (N_1812,N_1738,N_1752);
or U1813 (N_1813,N_1799,N_1746);
and U1814 (N_1814,N_1719,N_1756);
nand U1815 (N_1815,N_1790,N_1759);
nand U1816 (N_1816,N_1720,N_1761);
or U1817 (N_1817,N_1735,N_1722);
nand U1818 (N_1818,N_1773,N_1770);
nand U1819 (N_1819,N_1723,N_1796);
nand U1820 (N_1820,N_1795,N_1713);
nor U1821 (N_1821,N_1729,N_1703);
and U1822 (N_1822,N_1748,N_1728);
and U1823 (N_1823,N_1781,N_1742);
and U1824 (N_1824,N_1776,N_1793);
and U1825 (N_1825,N_1718,N_1786);
nor U1826 (N_1826,N_1792,N_1711);
or U1827 (N_1827,N_1733,N_1798);
and U1828 (N_1828,N_1783,N_1755);
and U1829 (N_1829,N_1725,N_1743);
nand U1830 (N_1830,N_1753,N_1778);
nand U1831 (N_1831,N_1766,N_1780);
or U1832 (N_1832,N_1701,N_1789);
and U1833 (N_1833,N_1763,N_1784);
or U1834 (N_1834,N_1744,N_1768);
nand U1835 (N_1835,N_1712,N_1740);
nor U1836 (N_1836,N_1721,N_1741);
and U1837 (N_1837,N_1705,N_1702);
nand U1838 (N_1838,N_1706,N_1734);
nand U1839 (N_1839,N_1747,N_1708);
xor U1840 (N_1840,N_1745,N_1707);
nand U1841 (N_1841,N_1782,N_1757);
and U1842 (N_1842,N_1716,N_1710);
and U1843 (N_1843,N_1737,N_1717);
and U1844 (N_1844,N_1754,N_1700);
nand U1845 (N_1845,N_1704,N_1732);
nor U1846 (N_1846,N_1727,N_1779);
and U1847 (N_1847,N_1771,N_1714);
nor U1848 (N_1848,N_1764,N_1758);
or U1849 (N_1849,N_1760,N_1769);
nor U1850 (N_1850,N_1748,N_1702);
and U1851 (N_1851,N_1781,N_1739);
nor U1852 (N_1852,N_1713,N_1758);
and U1853 (N_1853,N_1791,N_1794);
or U1854 (N_1854,N_1729,N_1700);
or U1855 (N_1855,N_1787,N_1785);
nand U1856 (N_1856,N_1770,N_1718);
nand U1857 (N_1857,N_1712,N_1778);
and U1858 (N_1858,N_1728,N_1783);
nor U1859 (N_1859,N_1734,N_1710);
or U1860 (N_1860,N_1787,N_1731);
and U1861 (N_1861,N_1725,N_1757);
nor U1862 (N_1862,N_1760,N_1785);
nand U1863 (N_1863,N_1755,N_1740);
or U1864 (N_1864,N_1741,N_1715);
nor U1865 (N_1865,N_1774,N_1714);
and U1866 (N_1866,N_1727,N_1721);
and U1867 (N_1867,N_1785,N_1715);
nand U1868 (N_1868,N_1781,N_1726);
and U1869 (N_1869,N_1728,N_1719);
nor U1870 (N_1870,N_1744,N_1793);
and U1871 (N_1871,N_1749,N_1723);
or U1872 (N_1872,N_1702,N_1792);
or U1873 (N_1873,N_1748,N_1749);
and U1874 (N_1874,N_1784,N_1755);
nand U1875 (N_1875,N_1745,N_1792);
nand U1876 (N_1876,N_1701,N_1773);
nor U1877 (N_1877,N_1788,N_1735);
nor U1878 (N_1878,N_1735,N_1738);
and U1879 (N_1879,N_1780,N_1708);
and U1880 (N_1880,N_1778,N_1782);
or U1881 (N_1881,N_1745,N_1702);
nand U1882 (N_1882,N_1765,N_1764);
nand U1883 (N_1883,N_1792,N_1769);
or U1884 (N_1884,N_1797,N_1703);
or U1885 (N_1885,N_1764,N_1783);
nand U1886 (N_1886,N_1762,N_1702);
and U1887 (N_1887,N_1787,N_1773);
nor U1888 (N_1888,N_1774,N_1708);
or U1889 (N_1889,N_1718,N_1738);
and U1890 (N_1890,N_1777,N_1727);
and U1891 (N_1891,N_1783,N_1710);
and U1892 (N_1892,N_1761,N_1743);
nand U1893 (N_1893,N_1750,N_1723);
nor U1894 (N_1894,N_1709,N_1777);
nand U1895 (N_1895,N_1749,N_1737);
and U1896 (N_1896,N_1729,N_1773);
and U1897 (N_1897,N_1769,N_1711);
nor U1898 (N_1898,N_1754,N_1737);
nand U1899 (N_1899,N_1704,N_1789);
or U1900 (N_1900,N_1866,N_1824);
and U1901 (N_1901,N_1892,N_1812);
or U1902 (N_1902,N_1810,N_1897);
and U1903 (N_1903,N_1895,N_1831);
and U1904 (N_1904,N_1829,N_1819);
and U1905 (N_1905,N_1885,N_1888);
and U1906 (N_1906,N_1849,N_1847);
or U1907 (N_1907,N_1863,N_1889);
nand U1908 (N_1908,N_1899,N_1877);
nand U1909 (N_1909,N_1893,N_1868);
and U1910 (N_1910,N_1805,N_1835);
nand U1911 (N_1911,N_1882,N_1858);
nor U1912 (N_1912,N_1871,N_1867);
or U1913 (N_1913,N_1878,N_1803);
or U1914 (N_1914,N_1883,N_1840);
and U1915 (N_1915,N_1813,N_1854);
nand U1916 (N_1916,N_1881,N_1860);
and U1917 (N_1917,N_1859,N_1875);
nand U1918 (N_1918,N_1839,N_1820);
or U1919 (N_1919,N_1815,N_1862);
nand U1920 (N_1920,N_1876,N_1822);
or U1921 (N_1921,N_1879,N_1865);
or U1922 (N_1922,N_1896,N_1830);
or U1923 (N_1923,N_1870,N_1845);
and U1924 (N_1924,N_1872,N_1821);
or U1925 (N_1925,N_1811,N_1848);
nand U1926 (N_1926,N_1836,N_1825);
or U1927 (N_1927,N_1886,N_1894);
or U1928 (N_1928,N_1828,N_1887);
or U1929 (N_1929,N_1891,N_1808);
xnor U1930 (N_1930,N_1841,N_1801);
nand U1931 (N_1931,N_1827,N_1818);
or U1932 (N_1932,N_1809,N_1817);
and U1933 (N_1933,N_1833,N_1834);
or U1934 (N_1934,N_1846,N_1898);
or U1935 (N_1935,N_1852,N_1806);
nor U1936 (N_1936,N_1843,N_1800);
or U1937 (N_1937,N_1857,N_1838);
or U1938 (N_1938,N_1850,N_1853);
nor U1939 (N_1939,N_1804,N_1807);
and U1940 (N_1940,N_1844,N_1855);
nor U1941 (N_1941,N_1890,N_1814);
nor U1942 (N_1942,N_1816,N_1826);
and U1943 (N_1943,N_1823,N_1884);
and U1944 (N_1944,N_1802,N_1873);
and U1945 (N_1945,N_1851,N_1856);
nor U1946 (N_1946,N_1842,N_1864);
and U1947 (N_1947,N_1861,N_1869);
and U1948 (N_1948,N_1880,N_1874);
or U1949 (N_1949,N_1832,N_1837);
and U1950 (N_1950,N_1817,N_1897);
nor U1951 (N_1951,N_1844,N_1820);
and U1952 (N_1952,N_1831,N_1847);
or U1953 (N_1953,N_1839,N_1824);
nor U1954 (N_1954,N_1898,N_1807);
nor U1955 (N_1955,N_1828,N_1847);
xor U1956 (N_1956,N_1850,N_1881);
and U1957 (N_1957,N_1899,N_1878);
or U1958 (N_1958,N_1842,N_1811);
and U1959 (N_1959,N_1896,N_1878);
nand U1960 (N_1960,N_1816,N_1837);
and U1961 (N_1961,N_1847,N_1805);
or U1962 (N_1962,N_1865,N_1897);
or U1963 (N_1963,N_1815,N_1800);
or U1964 (N_1964,N_1838,N_1848);
nand U1965 (N_1965,N_1802,N_1833);
or U1966 (N_1966,N_1846,N_1851);
nor U1967 (N_1967,N_1896,N_1881);
and U1968 (N_1968,N_1821,N_1831);
or U1969 (N_1969,N_1860,N_1893);
and U1970 (N_1970,N_1878,N_1870);
and U1971 (N_1971,N_1850,N_1889);
and U1972 (N_1972,N_1812,N_1883);
and U1973 (N_1973,N_1857,N_1867);
and U1974 (N_1974,N_1864,N_1874);
and U1975 (N_1975,N_1822,N_1896);
xor U1976 (N_1976,N_1899,N_1841);
nor U1977 (N_1977,N_1803,N_1850);
nand U1978 (N_1978,N_1826,N_1817);
nand U1979 (N_1979,N_1801,N_1868);
nand U1980 (N_1980,N_1850,N_1840);
nor U1981 (N_1981,N_1873,N_1888);
nand U1982 (N_1982,N_1811,N_1882);
xnor U1983 (N_1983,N_1832,N_1894);
nor U1984 (N_1984,N_1826,N_1824);
and U1985 (N_1985,N_1864,N_1878);
nor U1986 (N_1986,N_1852,N_1836);
xor U1987 (N_1987,N_1846,N_1868);
and U1988 (N_1988,N_1820,N_1800);
or U1989 (N_1989,N_1817,N_1819);
and U1990 (N_1990,N_1852,N_1891);
xor U1991 (N_1991,N_1871,N_1879);
nand U1992 (N_1992,N_1814,N_1886);
or U1993 (N_1993,N_1819,N_1827);
and U1994 (N_1994,N_1800,N_1894);
and U1995 (N_1995,N_1885,N_1872);
nor U1996 (N_1996,N_1825,N_1813);
nand U1997 (N_1997,N_1836,N_1887);
and U1998 (N_1998,N_1825,N_1847);
or U1999 (N_1999,N_1876,N_1851);
nand U2000 (N_2000,N_1909,N_1997);
nand U2001 (N_2001,N_1937,N_1965);
nor U2002 (N_2002,N_1935,N_1933);
or U2003 (N_2003,N_1946,N_1947);
or U2004 (N_2004,N_1994,N_1914);
nand U2005 (N_2005,N_1916,N_1989);
and U2006 (N_2006,N_1969,N_1966);
nand U2007 (N_2007,N_1918,N_1939);
nor U2008 (N_2008,N_1974,N_1982);
nor U2009 (N_2009,N_1949,N_1921);
nor U2010 (N_2010,N_1911,N_1905);
and U2011 (N_2011,N_1993,N_1951);
or U2012 (N_2012,N_1901,N_1922);
and U2013 (N_2013,N_1998,N_1996);
and U2014 (N_2014,N_1983,N_1971);
nand U2015 (N_2015,N_1931,N_1978);
or U2016 (N_2016,N_1912,N_1925);
and U2017 (N_2017,N_1957,N_1995);
or U2018 (N_2018,N_1924,N_1908);
and U2019 (N_2019,N_1975,N_1988);
or U2020 (N_2020,N_1900,N_1953);
or U2021 (N_2021,N_1906,N_1944);
or U2022 (N_2022,N_1992,N_1943);
nand U2023 (N_2023,N_1981,N_1929);
and U2024 (N_2024,N_1930,N_1938);
and U2025 (N_2025,N_1941,N_1904);
nor U2026 (N_2026,N_1903,N_1984);
nand U2027 (N_2027,N_1920,N_1963);
nand U2028 (N_2028,N_1932,N_1959);
nor U2029 (N_2029,N_1952,N_1910);
nor U2030 (N_2030,N_1923,N_1915);
nand U2031 (N_2031,N_1985,N_1934);
or U2032 (N_2032,N_1973,N_1987);
nand U2033 (N_2033,N_1926,N_1907);
or U2034 (N_2034,N_1956,N_1972);
nand U2035 (N_2035,N_1942,N_1948);
or U2036 (N_2036,N_1999,N_1990);
and U2037 (N_2037,N_1967,N_1902);
nand U2038 (N_2038,N_1958,N_1950);
nor U2039 (N_2039,N_1979,N_1960);
and U2040 (N_2040,N_1928,N_1964);
nand U2041 (N_2041,N_1970,N_1913);
or U2042 (N_2042,N_1968,N_1940);
nand U2043 (N_2043,N_1919,N_1962);
nand U2044 (N_2044,N_1986,N_1955);
nor U2045 (N_2045,N_1991,N_1961);
or U2046 (N_2046,N_1980,N_1976);
and U2047 (N_2047,N_1936,N_1927);
nor U2048 (N_2048,N_1945,N_1917);
and U2049 (N_2049,N_1954,N_1977);
nand U2050 (N_2050,N_1930,N_1918);
nand U2051 (N_2051,N_1900,N_1950);
or U2052 (N_2052,N_1949,N_1982);
xnor U2053 (N_2053,N_1948,N_1930);
and U2054 (N_2054,N_1916,N_1994);
nand U2055 (N_2055,N_1965,N_1903);
nand U2056 (N_2056,N_1935,N_1936);
nor U2057 (N_2057,N_1901,N_1918);
and U2058 (N_2058,N_1944,N_1981);
nor U2059 (N_2059,N_1952,N_1934);
and U2060 (N_2060,N_1912,N_1915);
nand U2061 (N_2061,N_1907,N_1976);
or U2062 (N_2062,N_1932,N_1993);
nand U2063 (N_2063,N_1924,N_1943);
nand U2064 (N_2064,N_1998,N_1916);
and U2065 (N_2065,N_1983,N_1910);
nand U2066 (N_2066,N_1959,N_1951);
and U2067 (N_2067,N_1916,N_1940);
or U2068 (N_2068,N_1991,N_1940);
or U2069 (N_2069,N_1922,N_1996);
or U2070 (N_2070,N_1999,N_1954);
nor U2071 (N_2071,N_1942,N_1905);
nor U2072 (N_2072,N_1987,N_1961);
nor U2073 (N_2073,N_1902,N_1964);
and U2074 (N_2074,N_1987,N_1918);
nand U2075 (N_2075,N_1997,N_1963);
nand U2076 (N_2076,N_1976,N_1914);
or U2077 (N_2077,N_1936,N_1983);
or U2078 (N_2078,N_1918,N_1950);
and U2079 (N_2079,N_1916,N_1942);
or U2080 (N_2080,N_1923,N_1971);
and U2081 (N_2081,N_1994,N_1980);
nand U2082 (N_2082,N_1968,N_1991);
nand U2083 (N_2083,N_1933,N_1945);
nand U2084 (N_2084,N_1936,N_1988);
or U2085 (N_2085,N_1940,N_1979);
nand U2086 (N_2086,N_1902,N_1991);
nand U2087 (N_2087,N_1961,N_1931);
nand U2088 (N_2088,N_1928,N_1936);
xnor U2089 (N_2089,N_1994,N_1991);
and U2090 (N_2090,N_1919,N_1933);
nand U2091 (N_2091,N_1960,N_1936);
and U2092 (N_2092,N_1961,N_1917);
or U2093 (N_2093,N_1990,N_1995);
nor U2094 (N_2094,N_1978,N_1939);
and U2095 (N_2095,N_1910,N_1959);
nor U2096 (N_2096,N_1988,N_1944);
nor U2097 (N_2097,N_1951,N_1995);
nor U2098 (N_2098,N_1950,N_1965);
xor U2099 (N_2099,N_1906,N_1995);
xnor U2100 (N_2100,N_2070,N_2044);
nor U2101 (N_2101,N_2069,N_2013);
or U2102 (N_2102,N_2036,N_2005);
and U2103 (N_2103,N_2067,N_2064);
nor U2104 (N_2104,N_2001,N_2055);
nand U2105 (N_2105,N_2084,N_2008);
nand U2106 (N_2106,N_2086,N_2078);
and U2107 (N_2107,N_2068,N_2030);
nand U2108 (N_2108,N_2077,N_2056);
nand U2109 (N_2109,N_2079,N_2090);
nand U2110 (N_2110,N_2071,N_2073);
or U2111 (N_2111,N_2065,N_2000);
nor U2112 (N_2112,N_2095,N_2096);
nand U2113 (N_2113,N_2029,N_2022);
and U2114 (N_2114,N_2066,N_2088);
nand U2115 (N_2115,N_2082,N_2033);
and U2116 (N_2116,N_2019,N_2031);
and U2117 (N_2117,N_2028,N_2007);
or U2118 (N_2118,N_2032,N_2010);
or U2119 (N_2119,N_2015,N_2012);
nand U2120 (N_2120,N_2061,N_2011);
or U2121 (N_2121,N_2023,N_2020);
nand U2122 (N_2122,N_2024,N_2051);
and U2123 (N_2123,N_2091,N_2076);
and U2124 (N_2124,N_2050,N_2060);
or U2125 (N_2125,N_2081,N_2087);
nor U2126 (N_2126,N_2062,N_2058);
and U2127 (N_2127,N_2049,N_2047);
and U2128 (N_2128,N_2080,N_2006);
and U2129 (N_2129,N_2097,N_2083);
nand U2130 (N_2130,N_2025,N_2027);
nand U2131 (N_2131,N_2052,N_2048);
and U2132 (N_2132,N_2098,N_2053);
nand U2133 (N_2133,N_2094,N_2009);
and U2134 (N_2134,N_2035,N_2043);
nor U2135 (N_2135,N_2002,N_2074);
or U2136 (N_2136,N_2004,N_2014);
or U2137 (N_2137,N_2003,N_2045);
or U2138 (N_2138,N_2034,N_2039);
and U2139 (N_2139,N_2026,N_2038);
or U2140 (N_2140,N_2072,N_2092);
and U2141 (N_2141,N_2063,N_2075);
and U2142 (N_2142,N_2042,N_2099);
nand U2143 (N_2143,N_2041,N_2089);
and U2144 (N_2144,N_2057,N_2059);
xnor U2145 (N_2145,N_2017,N_2046);
nor U2146 (N_2146,N_2085,N_2021);
nor U2147 (N_2147,N_2016,N_2018);
nand U2148 (N_2148,N_2040,N_2093);
nor U2149 (N_2149,N_2054,N_2037);
nand U2150 (N_2150,N_2033,N_2020);
or U2151 (N_2151,N_2029,N_2074);
nor U2152 (N_2152,N_2067,N_2091);
or U2153 (N_2153,N_2012,N_2003);
nand U2154 (N_2154,N_2013,N_2099);
nor U2155 (N_2155,N_2096,N_2022);
nand U2156 (N_2156,N_2013,N_2045);
nor U2157 (N_2157,N_2032,N_2025);
nor U2158 (N_2158,N_2056,N_2063);
nand U2159 (N_2159,N_2040,N_2010);
nor U2160 (N_2160,N_2066,N_2015);
nand U2161 (N_2161,N_2023,N_2036);
and U2162 (N_2162,N_2035,N_2008);
or U2163 (N_2163,N_2052,N_2017);
nand U2164 (N_2164,N_2059,N_2093);
nor U2165 (N_2165,N_2072,N_2021);
nand U2166 (N_2166,N_2049,N_2055);
or U2167 (N_2167,N_2070,N_2036);
nand U2168 (N_2168,N_2011,N_2075);
or U2169 (N_2169,N_2080,N_2064);
or U2170 (N_2170,N_2067,N_2055);
and U2171 (N_2171,N_2019,N_2006);
nand U2172 (N_2172,N_2072,N_2015);
nor U2173 (N_2173,N_2052,N_2026);
or U2174 (N_2174,N_2012,N_2062);
xnor U2175 (N_2175,N_2049,N_2067);
nand U2176 (N_2176,N_2066,N_2046);
and U2177 (N_2177,N_2038,N_2083);
nand U2178 (N_2178,N_2083,N_2061);
or U2179 (N_2179,N_2020,N_2074);
and U2180 (N_2180,N_2078,N_2002);
nor U2181 (N_2181,N_2035,N_2054);
and U2182 (N_2182,N_2098,N_2024);
and U2183 (N_2183,N_2022,N_2057);
or U2184 (N_2184,N_2004,N_2077);
nand U2185 (N_2185,N_2064,N_2087);
and U2186 (N_2186,N_2034,N_2095);
nand U2187 (N_2187,N_2064,N_2071);
nor U2188 (N_2188,N_2093,N_2018);
nor U2189 (N_2189,N_2077,N_2092);
nor U2190 (N_2190,N_2010,N_2099);
nor U2191 (N_2191,N_2008,N_2098);
nor U2192 (N_2192,N_2005,N_2037);
nor U2193 (N_2193,N_2089,N_2055);
or U2194 (N_2194,N_2068,N_2015);
and U2195 (N_2195,N_2067,N_2099);
nand U2196 (N_2196,N_2087,N_2040);
or U2197 (N_2197,N_2071,N_2043);
nand U2198 (N_2198,N_2019,N_2067);
or U2199 (N_2199,N_2089,N_2046);
and U2200 (N_2200,N_2131,N_2137);
or U2201 (N_2201,N_2194,N_2130);
nor U2202 (N_2202,N_2133,N_2189);
and U2203 (N_2203,N_2199,N_2147);
nand U2204 (N_2204,N_2121,N_2145);
nor U2205 (N_2205,N_2144,N_2168);
or U2206 (N_2206,N_2116,N_2174);
or U2207 (N_2207,N_2126,N_2105);
nand U2208 (N_2208,N_2141,N_2109);
or U2209 (N_2209,N_2110,N_2192);
and U2210 (N_2210,N_2124,N_2142);
and U2211 (N_2211,N_2106,N_2107);
or U2212 (N_2212,N_2167,N_2134);
xnor U2213 (N_2213,N_2112,N_2193);
nand U2214 (N_2214,N_2177,N_2103);
nand U2215 (N_2215,N_2195,N_2187);
nand U2216 (N_2216,N_2152,N_2161);
xnor U2217 (N_2217,N_2101,N_2169);
or U2218 (N_2218,N_2182,N_2188);
nor U2219 (N_2219,N_2191,N_2154);
nor U2220 (N_2220,N_2159,N_2151);
nor U2221 (N_2221,N_2128,N_2104);
and U2222 (N_2222,N_2111,N_2136);
nor U2223 (N_2223,N_2102,N_2171);
nand U2224 (N_2224,N_2186,N_2138);
nand U2225 (N_2225,N_2143,N_2160);
nand U2226 (N_2226,N_2178,N_2115);
xnor U2227 (N_2227,N_2162,N_2119);
and U2228 (N_2228,N_2158,N_2120);
and U2229 (N_2229,N_2164,N_2118);
and U2230 (N_2230,N_2175,N_2197);
and U2231 (N_2231,N_2148,N_2149);
or U2232 (N_2232,N_2163,N_2185);
or U2233 (N_2233,N_2114,N_2146);
and U2234 (N_2234,N_2184,N_2196);
and U2235 (N_2235,N_2179,N_2153);
nand U2236 (N_2236,N_2166,N_2156);
nor U2237 (N_2237,N_2123,N_2183);
nor U2238 (N_2238,N_2190,N_2122);
and U2239 (N_2239,N_2117,N_2129);
or U2240 (N_2240,N_2132,N_2181);
nand U2241 (N_2241,N_2127,N_2173);
nor U2242 (N_2242,N_2172,N_2100);
xnor U2243 (N_2243,N_2198,N_2108);
or U2244 (N_2244,N_2155,N_2150);
nand U2245 (N_2245,N_2113,N_2165);
and U2246 (N_2246,N_2140,N_2125);
nor U2247 (N_2247,N_2170,N_2139);
nor U2248 (N_2248,N_2176,N_2180);
nand U2249 (N_2249,N_2157,N_2135);
and U2250 (N_2250,N_2163,N_2192);
nor U2251 (N_2251,N_2194,N_2171);
or U2252 (N_2252,N_2101,N_2151);
nor U2253 (N_2253,N_2174,N_2155);
nor U2254 (N_2254,N_2161,N_2104);
or U2255 (N_2255,N_2170,N_2147);
nand U2256 (N_2256,N_2134,N_2155);
or U2257 (N_2257,N_2165,N_2104);
nor U2258 (N_2258,N_2165,N_2159);
and U2259 (N_2259,N_2154,N_2116);
nand U2260 (N_2260,N_2115,N_2180);
and U2261 (N_2261,N_2125,N_2102);
and U2262 (N_2262,N_2123,N_2180);
nor U2263 (N_2263,N_2158,N_2140);
nand U2264 (N_2264,N_2150,N_2112);
or U2265 (N_2265,N_2196,N_2199);
or U2266 (N_2266,N_2179,N_2137);
or U2267 (N_2267,N_2107,N_2178);
or U2268 (N_2268,N_2181,N_2147);
nor U2269 (N_2269,N_2100,N_2116);
or U2270 (N_2270,N_2118,N_2105);
nor U2271 (N_2271,N_2196,N_2108);
nand U2272 (N_2272,N_2172,N_2160);
nor U2273 (N_2273,N_2152,N_2166);
or U2274 (N_2274,N_2164,N_2183);
nor U2275 (N_2275,N_2161,N_2132);
or U2276 (N_2276,N_2103,N_2115);
or U2277 (N_2277,N_2103,N_2157);
nor U2278 (N_2278,N_2128,N_2193);
or U2279 (N_2279,N_2126,N_2154);
nor U2280 (N_2280,N_2152,N_2190);
or U2281 (N_2281,N_2121,N_2119);
nor U2282 (N_2282,N_2117,N_2141);
nand U2283 (N_2283,N_2113,N_2123);
or U2284 (N_2284,N_2175,N_2199);
nand U2285 (N_2285,N_2123,N_2187);
and U2286 (N_2286,N_2155,N_2106);
or U2287 (N_2287,N_2116,N_2110);
nor U2288 (N_2288,N_2147,N_2179);
nand U2289 (N_2289,N_2117,N_2176);
nand U2290 (N_2290,N_2192,N_2182);
and U2291 (N_2291,N_2117,N_2151);
and U2292 (N_2292,N_2188,N_2100);
and U2293 (N_2293,N_2109,N_2188);
or U2294 (N_2294,N_2199,N_2136);
nand U2295 (N_2295,N_2135,N_2192);
nand U2296 (N_2296,N_2133,N_2171);
and U2297 (N_2297,N_2117,N_2197);
nand U2298 (N_2298,N_2175,N_2116);
or U2299 (N_2299,N_2124,N_2132);
xnor U2300 (N_2300,N_2266,N_2275);
and U2301 (N_2301,N_2227,N_2267);
nand U2302 (N_2302,N_2278,N_2236);
or U2303 (N_2303,N_2244,N_2276);
nor U2304 (N_2304,N_2280,N_2265);
nand U2305 (N_2305,N_2230,N_2295);
and U2306 (N_2306,N_2260,N_2270);
and U2307 (N_2307,N_2291,N_2239);
nand U2308 (N_2308,N_2247,N_2256);
nand U2309 (N_2309,N_2282,N_2297);
xnor U2310 (N_2310,N_2219,N_2211);
and U2311 (N_2311,N_2246,N_2251);
and U2312 (N_2312,N_2279,N_2212);
and U2313 (N_2313,N_2294,N_2245);
and U2314 (N_2314,N_2252,N_2250);
or U2315 (N_2315,N_2223,N_2284);
and U2316 (N_2316,N_2285,N_2216);
and U2317 (N_2317,N_2209,N_2262);
or U2318 (N_2318,N_2237,N_2255);
or U2319 (N_2319,N_2273,N_2269);
or U2320 (N_2320,N_2253,N_2206);
and U2321 (N_2321,N_2298,N_2202);
nand U2322 (N_2322,N_2221,N_2268);
nor U2323 (N_2323,N_2296,N_2261);
nor U2324 (N_2324,N_2254,N_2203);
nand U2325 (N_2325,N_2241,N_2225);
or U2326 (N_2326,N_2213,N_2271);
xor U2327 (N_2327,N_2287,N_2242);
nor U2328 (N_2328,N_2231,N_2204);
nor U2329 (N_2329,N_2218,N_2283);
nand U2330 (N_2330,N_2288,N_2248);
and U2331 (N_2331,N_2200,N_2263);
or U2332 (N_2332,N_2201,N_2233);
nand U2333 (N_2333,N_2222,N_2220);
nand U2334 (N_2334,N_2293,N_2207);
nor U2335 (N_2335,N_2272,N_2274);
nand U2336 (N_2336,N_2214,N_2243);
nor U2337 (N_2337,N_2249,N_2264);
and U2338 (N_2338,N_2281,N_2226);
or U2339 (N_2339,N_2205,N_2277);
nor U2340 (N_2340,N_2259,N_2229);
or U2341 (N_2341,N_2234,N_2286);
and U2342 (N_2342,N_2217,N_2258);
or U2343 (N_2343,N_2289,N_2228);
nor U2344 (N_2344,N_2290,N_2208);
nand U2345 (N_2345,N_2292,N_2238);
xor U2346 (N_2346,N_2299,N_2232);
and U2347 (N_2347,N_2224,N_2210);
nor U2348 (N_2348,N_2240,N_2257);
nand U2349 (N_2349,N_2215,N_2235);
nor U2350 (N_2350,N_2280,N_2230);
or U2351 (N_2351,N_2201,N_2257);
or U2352 (N_2352,N_2208,N_2206);
or U2353 (N_2353,N_2248,N_2280);
and U2354 (N_2354,N_2234,N_2241);
xor U2355 (N_2355,N_2263,N_2205);
nand U2356 (N_2356,N_2265,N_2255);
and U2357 (N_2357,N_2266,N_2272);
and U2358 (N_2358,N_2225,N_2240);
nand U2359 (N_2359,N_2205,N_2214);
nor U2360 (N_2360,N_2257,N_2287);
and U2361 (N_2361,N_2228,N_2287);
and U2362 (N_2362,N_2283,N_2203);
nor U2363 (N_2363,N_2251,N_2288);
nor U2364 (N_2364,N_2241,N_2235);
xor U2365 (N_2365,N_2236,N_2232);
nor U2366 (N_2366,N_2268,N_2270);
nor U2367 (N_2367,N_2271,N_2276);
or U2368 (N_2368,N_2294,N_2282);
nor U2369 (N_2369,N_2242,N_2262);
nor U2370 (N_2370,N_2232,N_2218);
nand U2371 (N_2371,N_2242,N_2209);
xnor U2372 (N_2372,N_2269,N_2240);
nand U2373 (N_2373,N_2203,N_2290);
nor U2374 (N_2374,N_2288,N_2277);
or U2375 (N_2375,N_2207,N_2251);
nor U2376 (N_2376,N_2278,N_2267);
nand U2377 (N_2377,N_2228,N_2209);
or U2378 (N_2378,N_2224,N_2240);
or U2379 (N_2379,N_2211,N_2255);
nor U2380 (N_2380,N_2219,N_2250);
or U2381 (N_2381,N_2200,N_2223);
nand U2382 (N_2382,N_2207,N_2242);
nand U2383 (N_2383,N_2238,N_2203);
or U2384 (N_2384,N_2243,N_2232);
and U2385 (N_2385,N_2291,N_2247);
nor U2386 (N_2386,N_2266,N_2257);
nor U2387 (N_2387,N_2242,N_2294);
nor U2388 (N_2388,N_2238,N_2250);
nand U2389 (N_2389,N_2282,N_2217);
nor U2390 (N_2390,N_2272,N_2253);
nand U2391 (N_2391,N_2297,N_2296);
xor U2392 (N_2392,N_2266,N_2215);
and U2393 (N_2393,N_2284,N_2267);
or U2394 (N_2394,N_2203,N_2294);
nand U2395 (N_2395,N_2254,N_2200);
and U2396 (N_2396,N_2220,N_2216);
or U2397 (N_2397,N_2259,N_2263);
nor U2398 (N_2398,N_2275,N_2273);
and U2399 (N_2399,N_2283,N_2297);
or U2400 (N_2400,N_2331,N_2392);
nor U2401 (N_2401,N_2372,N_2349);
xor U2402 (N_2402,N_2321,N_2329);
nand U2403 (N_2403,N_2348,N_2328);
nor U2404 (N_2404,N_2373,N_2316);
or U2405 (N_2405,N_2394,N_2326);
and U2406 (N_2406,N_2374,N_2307);
or U2407 (N_2407,N_2376,N_2339);
and U2408 (N_2408,N_2335,N_2386);
and U2409 (N_2409,N_2300,N_2340);
and U2410 (N_2410,N_2365,N_2337);
or U2411 (N_2411,N_2342,N_2390);
and U2412 (N_2412,N_2370,N_2315);
or U2413 (N_2413,N_2338,N_2334);
or U2414 (N_2414,N_2378,N_2311);
nor U2415 (N_2415,N_2345,N_2343);
or U2416 (N_2416,N_2350,N_2356);
and U2417 (N_2417,N_2352,N_2319);
and U2418 (N_2418,N_2324,N_2333);
and U2419 (N_2419,N_2330,N_2367);
nor U2420 (N_2420,N_2308,N_2397);
nand U2421 (N_2421,N_2332,N_2369);
or U2422 (N_2422,N_2313,N_2325);
and U2423 (N_2423,N_2382,N_2317);
nor U2424 (N_2424,N_2381,N_2398);
or U2425 (N_2425,N_2346,N_2368);
and U2426 (N_2426,N_2357,N_2318);
nor U2427 (N_2427,N_2309,N_2385);
and U2428 (N_2428,N_2387,N_2379);
xor U2429 (N_2429,N_2351,N_2302);
or U2430 (N_2430,N_2312,N_2375);
nor U2431 (N_2431,N_2362,N_2380);
nor U2432 (N_2432,N_2305,N_2354);
or U2433 (N_2433,N_2344,N_2383);
nor U2434 (N_2434,N_2314,N_2358);
and U2435 (N_2435,N_2320,N_2389);
nand U2436 (N_2436,N_2322,N_2301);
nor U2437 (N_2437,N_2355,N_2323);
and U2438 (N_2438,N_2364,N_2341);
nand U2439 (N_2439,N_2310,N_2377);
and U2440 (N_2440,N_2306,N_2304);
and U2441 (N_2441,N_2303,N_2393);
nand U2442 (N_2442,N_2361,N_2395);
or U2443 (N_2443,N_2336,N_2399);
and U2444 (N_2444,N_2384,N_2396);
xnor U2445 (N_2445,N_2371,N_2360);
nand U2446 (N_2446,N_2363,N_2366);
nand U2447 (N_2447,N_2391,N_2327);
nand U2448 (N_2448,N_2359,N_2347);
nor U2449 (N_2449,N_2388,N_2353);
nor U2450 (N_2450,N_2339,N_2358);
and U2451 (N_2451,N_2315,N_2339);
or U2452 (N_2452,N_2381,N_2328);
nor U2453 (N_2453,N_2391,N_2331);
and U2454 (N_2454,N_2347,N_2330);
or U2455 (N_2455,N_2324,N_2365);
and U2456 (N_2456,N_2393,N_2397);
nor U2457 (N_2457,N_2318,N_2343);
and U2458 (N_2458,N_2352,N_2331);
and U2459 (N_2459,N_2358,N_2368);
nor U2460 (N_2460,N_2383,N_2334);
or U2461 (N_2461,N_2308,N_2354);
nand U2462 (N_2462,N_2389,N_2346);
xor U2463 (N_2463,N_2367,N_2350);
or U2464 (N_2464,N_2326,N_2304);
and U2465 (N_2465,N_2365,N_2316);
or U2466 (N_2466,N_2361,N_2388);
nor U2467 (N_2467,N_2300,N_2394);
and U2468 (N_2468,N_2379,N_2350);
or U2469 (N_2469,N_2364,N_2386);
or U2470 (N_2470,N_2320,N_2374);
nand U2471 (N_2471,N_2309,N_2365);
nor U2472 (N_2472,N_2329,N_2318);
nor U2473 (N_2473,N_2364,N_2321);
and U2474 (N_2474,N_2351,N_2308);
nor U2475 (N_2475,N_2394,N_2316);
nand U2476 (N_2476,N_2383,N_2319);
or U2477 (N_2477,N_2396,N_2353);
and U2478 (N_2478,N_2336,N_2308);
nor U2479 (N_2479,N_2390,N_2376);
or U2480 (N_2480,N_2360,N_2378);
nor U2481 (N_2481,N_2382,N_2393);
or U2482 (N_2482,N_2389,N_2317);
nor U2483 (N_2483,N_2335,N_2363);
and U2484 (N_2484,N_2380,N_2349);
nor U2485 (N_2485,N_2335,N_2327);
or U2486 (N_2486,N_2345,N_2302);
nor U2487 (N_2487,N_2300,N_2330);
and U2488 (N_2488,N_2315,N_2393);
or U2489 (N_2489,N_2393,N_2326);
nand U2490 (N_2490,N_2317,N_2311);
nor U2491 (N_2491,N_2363,N_2396);
and U2492 (N_2492,N_2306,N_2331);
or U2493 (N_2493,N_2309,N_2391);
or U2494 (N_2494,N_2380,N_2318);
nor U2495 (N_2495,N_2347,N_2367);
nor U2496 (N_2496,N_2341,N_2346);
and U2497 (N_2497,N_2326,N_2332);
nand U2498 (N_2498,N_2389,N_2329);
nor U2499 (N_2499,N_2312,N_2322);
xor U2500 (N_2500,N_2419,N_2421);
and U2501 (N_2501,N_2409,N_2454);
nand U2502 (N_2502,N_2438,N_2417);
and U2503 (N_2503,N_2443,N_2404);
nor U2504 (N_2504,N_2471,N_2477);
and U2505 (N_2505,N_2401,N_2455);
or U2506 (N_2506,N_2433,N_2484);
nor U2507 (N_2507,N_2446,N_2463);
nand U2508 (N_2508,N_2479,N_2457);
or U2509 (N_2509,N_2423,N_2440);
nor U2510 (N_2510,N_2428,N_2424);
or U2511 (N_2511,N_2422,N_2472);
nor U2512 (N_2512,N_2482,N_2447);
nand U2513 (N_2513,N_2449,N_2437);
nand U2514 (N_2514,N_2458,N_2451);
and U2515 (N_2515,N_2462,N_2431);
nor U2516 (N_2516,N_2441,N_2489);
nand U2517 (N_2517,N_2465,N_2429);
nand U2518 (N_2518,N_2402,N_2420);
nor U2519 (N_2519,N_2430,N_2445);
or U2520 (N_2520,N_2498,N_2450);
nor U2521 (N_2521,N_2411,N_2494);
nor U2522 (N_2522,N_2416,N_2407);
nand U2523 (N_2523,N_2478,N_2476);
nand U2524 (N_2524,N_2493,N_2453);
nand U2525 (N_2525,N_2499,N_2480);
nor U2526 (N_2526,N_2444,N_2403);
or U2527 (N_2527,N_2492,N_2406);
and U2528 (N_2528,N_2468,N_2464);
nand U2529 (N_2529,N_2436,N_2483);
nor U2530 (N_2530,N_2427,N_2466);
or U2531 (N_2531,N_2442,N_2408);
or U2532 (N_2532,N_2475,N_2481);
nand U2533 (N_2533,N_2469,N_2467);
nor U2534 (N_2534,N_2439,N_2488);
nand U2535 (N_2535,N_2414,N_2459);
and U2536 (N_2536,N_2410,N_2485);
nand U2537 (N_2537,N_2435,N_2461);
or U2538 (N_2538,N_2491,N_2495);
and U2539 (N_2539,N_2434,N_2412);
nand U2540 (N_2540,N_2452,N_2486);
nand U2541 (N_2541,N_2456,N_2474);
nor U2542 (N_2542,N_2413,N_2490);
or U2543 (N_2543,N_2448,N_2496);
nor U2544 (N_2544,N_2425,N_2400);
or U2545 (N_2545,N_2473,N_2426);
or U2546 (N_2546,N_2418,N_2432);
or U2547 (N_2547,N_2460,N_2415);
and U2548 (N_2548,N_2497,N_2405);
nor U2549 (N_2549,N_2470,N_2487);
nor U2550 (N_2550,N_2473,N_2480);
or U2551 (N_2551,N_2459,N_2408);
and U2552 (N_2552,N_2465,N_2414);
or U2553 (N_2553,N_2475,N_2434);
and U2554 (N_2554,N_2483,N_2423);
or U2555 (N_2555,N_2440,N_2455);
and U2556 (N_2556,N_2454,N_2414);
or U2557 (N_2557,N_2489,N_2451);
and U2558 (N_2558,N_2474,N_2412);
nor U2559 (N_2559,N_2436,N_2481);
and U2560 (N_2560,N_2437,N_2461);
nand U2561 (N_2561,N_2437,N_2466);
or U2562 (N_2562,N_2467,N_2415);
or U2563 (N_2563,N_2436,N_2439);
or U2564 (N_2564,N_2429,N_2443);
nand U2565 (N_2565,N_2422,N_2420);
nand U2566 (N_2566,N_2457,N_2420);
nand U2567 (N_2567,N_2496,N_2405);
nor U2568 (N_2568,N_2435,N_2463);
or U2569 (N_2569,N_2498,N_2403);
or U2570 (N_2570,N_2443,N_2428);
or U2571 (N_2571,N_2466,N_2426);
and U2572 (N_2572,N_2416,N_2438);
nor U2573 (N_2573,N_2465,N_2462);
nand U2574 (N_2574,N_2485,N_2422);
and U2575 (N_2575,N_2497,N_2487);
and U2576 (N_2576,N_2401,N_2464);
nand U2577 (N_2577,N_2439,N_2408);
and U2578 (N_2578,N_2424,N_2489);
nor U2579 (N_2579,N_2433,N_2453);
or U2580 (N_2580,N_2439,N_2487);
and U2581 (N_2581,N_2464,N_2470);
or U2582 (N_2582,N_2455,N_2472);
or U2583 (N_2583,N_2411,N_2417);
nand U2584 (N_2584,N_2449,N_2419);
nand U2585 (N_2585,N_2433,N_2472);
nand U2586 (N_2586,N_2474,N_2429);
and U2587 (N_2587,N_2478,N_2498);
and U2588 (N_2588,N_2488,N_2418);
nand U2589 (N_2589,N_2463,N_2487);
nand U2590 (N_2590,N_2405,N_2420);
and U2591 (N_2591,N_2456,N_2484);
nand U2592 (N_2592,N_2480,N_2471);
and U2593 (N_2593,N_2465,N_2447);
nand U2594 (N_2594,N_2476,N_2490);
or U2595 (N_2595,N_2406,N_2409);
nor U2596 (N_2596,N_2490,N_2491);
and U2597 (N_2597,N_2481,N_2446);
nor U2598 (N_2598,N_2415,N_2453);
nand U2599 (N_2599,N_2459,N_2431);
nand U2600 (N_2600,N_2596,N_2502);
nand U2601 (N_2601,N_2551,N_2556);
and U2602 (N_2602,N_2507,N_2524);
or U2603 (N_2603,N_2563,N_2565);
nand U2604 (N_2604,N_2567,N_2575);
xnor U2605 (N_2605,N_2521,N_2532);
or U2606 (N_2606,N_2553,N_2541);
nand U2607 (N_2607,N_2511,N_2539);
nand U2608 (N_2608,N_2585,N_2548);
nor U2609 (N_2609,N_2594,N_2529);
and U2610 (N_2610,N_2552,N_2543);
xnor U2611 (N_2611,N_2582,N_2508);
nand U2612 (N_2612,N_2591,N_2590);
and U2613 (N_2613,N_2522,N_2560);
or U2614 (N_2614,N_2527,N_2588);
and U2615 (N_2615,N_2569,N_2501);
or U2616 (N_2616,N_2534,N_2530);
nor U2617 (N_2617,N_2528,N_2577);
nand U2618 (N_2618,N_2513,N_2557);
and U2619 (N_2619,N_2549,N_2520);
nand U2620 (N_2620,N_2576,N_2525);
nand U2621 (N_2621,N_2566,N_2535);
nand U2622 (N_2622,N_2568,N_2559);
nand U2623 (N_2623,N_2504,N_2518);
nand U2624 (N_2624,N_2516,N_2538);
nand U2625 (N_2625,N_2579,N_2597);
nor U2626 (N_2626,N_2550,N_2546);
or U2627 (N_2627,N_2514,N_2533);
and U2628 (N_2628,N_2506,N_2571);
or U2629 (N_2629,N_2558,N_2505);
nor U2630 (N_2630,N_2572,N_2581);
nor U2631 (N_2631,N_2570,N_2580);
and U2632 (N_2632,N_2545,N_2500);
nor U2633 (N_2633,N_2584,N_2573);
nand U2634 (N_2634,N_2536,N_2595);
and U2635 (N_2635,N_2510,N_2554);
nand U2636 (N_2636,N_2574,N_2540);
xnor U2637 (N_2637,N_2537,N_2586);
or U2638 (N_2638,N_2587,N_2517);
nor U2639 (N_2639,N_2547,N_2589);
and U2640 (N_2640,N_2544,N_2578);
or U2641 (N_2641,N_2598,N_2599);
and U2642 (N_2642,N_2509,N_2512);
and U2643 (N_2643,N_2564,N_2526);
or U2644 (N_2644,N_2592,N_2503);
and U2645 (N_2645,N_2515,N_2593);
nand U2646 (N_2646,N_2523,N_2562);
nand U2647 (N_2647,N_2531,N_2519);
nand U2648 (N_2648,N_2555,N_2561);
and U2649 (N_2649,N_2542,N_2583);
and U2650 (N_2650,N_2520,N_2524);
nor U2651 (N_2651,N_2599,N_2557);
and U2652 (N_2652,N_2551,N_2536);
nor U2653 (N_2653,N_2516,N_2509);
nor U2654 (N_2654,N_2561,N_2578);
or U2655 (N_2655,N_2512,N_2597);
xor U2656 (N_2656,N_2550,N_2583);
or U2657 (N_2657,N_2515,N_2544);
or U2658 (N_2658,N_2532,N_2583);
and U2659 (N_2659,N_2563,N_2596);
and U2660 (N_2660,N_2598,N_2500);
nand U2661 (N_2661,N_2542,N_2523);
nor U2662 (N_2662,N_2565,N_2529);
or U2663 (N_2663,N_2539,N_2591);
nand U2664 (N_2664,N_2550,N_2508);
or U2665 (N_2665,N_2524,N_2577);
and U2666 (N_2666,N_2589,N_2527);
nor U2667 (N_2667,N_2551,N_2523);
xnor U2668 (N_2668,N_2537,N_2526);
or U2669 (N_2669,N_2532,N_2555);
or U2670 (N_2670,N_2589,N_2525);
and U2671 (N_2671,N_2579,N_2568);
and U2672 (N_2672,N_2514,N_2530);
nand U2673 (N_2673,N_2534,N_2525);
and U2674 (N_2674,N_2529,N_2579);
or U2675 (N_2675,N_2544,N_2534);
and U2676 (N_2676,N_2571,N_2566);
and U2677 (N_2677,N_2570,N_2510);
xor U2678 (N_2678,N_2507,N_2569);
nand U2679 (N_2679,N_2535,N_2512);
and U2680 (N_2680,N_2535,N_2565);
and U2681 (N_2681,N_2588,N_2552);
nand U2682 (N_2682,N_2597,N_2556);
nor U2683 (N_2683,N_2591,N_2599);
or U2684 (N_2684,N_2502,N_2595);
or U2685 (N_2685,N_2509,N_2510);
or U2686 (N_2686,N_2587,N_2505);
or U2687 (N_2687,N_2578,N_2585);
nand U2688 (N_2688,N_2506,N_2595);
nor U2689 (N_2689,N_2576,N_2573);
nand U2690 (N_2690,N_2538,N_2561);
nand U2691 (N_2691,N_2530,N_2598);
nor U2692 (N_2692,N_2551,N_2538);
and U2693 (N_2693,N_2563,N_2553);
and U2694 (N_2694,N_2599,N_2578);
nand U2695 (N_2695,N_2531,N_2532);
and U2696 (N_2696,N_2592,N_2596);
nand U2697 (N_2697,N_2570,N_2576);
nand U2698 (N_2698,N_2551,N_2505);
and U2699 (N_2699,N_2504,N_2538);
or U2700 (N_2700,N_2640,N_2677);
or U2701 (N_2701,N_2644,N_2620);
and U2702 (N_2702,N_2657,N_2632);
nor U2703 (N_2703,N_2633,N_2605);
or U2704 (N_2704,N_2694,N_2668);
nand U2705 (N_2705,N_2645,N_2651);
nor U2706 (N_2706,N_2616,N_2696);
and U2707 (N_2707,N_2661,N_2664);
or U2708 (N_2708,N_2681,N_2663);
and U2709 (N_2709,N_2623,N_2627);
or U2710 (N_2710,N_2660,N_2603);
or U2711 (N_2711,N_2695,N_2669);
xor U2712 (N_2712,N_2637,N_2631);
or U2713 (N_2713,N_2647,N_2646);
or U2714 (N_2714,N_2670,N_2693);
nor U2715 (N_2715,N_2641,N_2672);
nand U2716 (N_2716,N_2671,N_2684);
and U2717 (N_2717,N_2665,N_2679);
nand U2718 (N_2718,N_2636,N_2609);
and U2719 (N_2719,N_2662,N_2689);
nor U2720 (N_2720,N_2630,N_2692);
or U2721 (N_2721,N_2610,N_2654);
or U2722 (N_2722,N_2659,N_2678);
nand U2723 (N_2723,N_2622,N_2674);
nor U2724 (N_2724,N_2613,N_2650);
xnor U2725 (N_2725,N_2619,N_2638);
and U2726 (N_2726,N_2621,N_2600);
nor U2727 (N_2727,N_2691,N_2690);
xor U2728 (N_2728,N_2653,N_2655);
nor U2729 (N_2729,N_2652,N_2624);
nor U2730 (N_2730,N_2688,N_2625);
nand U2731 (N_2731,N_2687,N_2673);
nor U2732 (N_2732,N_2699,N_2626);
or U2733 (N_2733,N_2628,N_2614);
nor U2734 (N_2734,N_2604,N_2698);
nand U2735 (N_2735,N_2648,N_2602);
nor U2736 (N_2736,N_2615,N_2607);
or U2737 (N_2737,N_2601,N_2611);
or U2738 (N_2738,N_2682,N_2656);
and U2739 (N_2739,N_2618,N_2634);
and U2740 (N_2740,N_2658,N_2685);
nand U2741 (N_2741,N_2639,N_2635);
and U2742 (N_2742,N_2680,N_2617);
or U2743 (N_2743,N_2697,N_2612);
and U2744 (N_2744,N_2629,N_2683);
nand U2745 (N_2745,N_2606,N_2643);
and U2746 (N_2746,N_2686,N_2667);
nand U2747 (N_2747,N_2666,N_2675);
nand U2748 (N_2748,N_2676,N_2642);
nand U2749 (N_2749,N_2608,N_2649);
or U2750 (N_2750,N_2669,N_2684);
nor U2751 (N_2751,N_2650,N_2618);
or U2752 (N_2752,N_2650,N_2646);
or U2753 (N_2753,N_2638,N_2636);
or U2754 (N_2754,N_2688,N_2606);
nand U2755 (N_2755,N_2630,N_2625);
and U2756 (N_2756,N_2633,N_2668);
nor U2757 (N_2757,N_2667,N_2613);
nor U2758 (N_2758,N_2649,N_2646);
nor U2759 (N_2759,N_2670,N_2657);
nand U2760 (N_2760,N_2694,N_2623);
and U2761 (N_2761,N_2669,N_2605);
or U2762 (N_2762,N_2605,N_2650);
or U2763 (N_2763,N_2635,N_2659);
and U2764 (N_2764,N_2674,N_2691);
or U2765 (N_2765,N_2635,N_2699);
and U2766 (N_2766,N_2674,N_2685);
and U2767 (N_2767,N_2684,N_2612);
nor U2768 (N_2768,N_2618,N_2640);
or U2769 (N_2769,N_2602,N_2670);
and U2770 (N_2770,N_2611,N_2624);
nand U2771 (N_2771,N_2658,N_2621);
or U2772 (N_2772,N_2687,N_2618);
or U2773 (N_2773,N_2695,N_2639);
and U2774 (N_2774,N_2671,N_2694);
and U2775 (N_2775,N_2641,N_2689);
or U2776 (N_2776,N_2651,N_2687);
or U2777 (N_2777,N_2628,N_2676);
or U2778 (N_2778,N_2690,N_2627);
and U2779 (N_2779,N_2667,N_2690);
or U2780 (N_2780,N_2636,N_2604);
and U2781 (N_2781,N_2686,N_2668);
or U2782 (N_2782,N_2693,N_2615);
nand U2783 (N_2783,N_2658,N_2648);
or U2784 (N_2784,N_2688,N_2607);
nor U2785 (N_2785,N_2644,N_2641);
nor U2786 (N_2786,N_2658,N_2670);
nor U2787 (N_2787,N_2676,N_2691);
and U2788 (N_2788,N_2677,N_2687);
or U2789 (N_2789,N_2600,N_2636);
nand U2790 (N_2790,N_2614,N_2668);
xnor U2791 (N_2791,N_2690,N_2656);
nor U2792 (N_2792,N_2676,N_2661);
and U2793 (N_2793,N_2660,N_2659);
and U2794 (N_2794,N_2690,N_2635);
or U2795 (N_2795,N_2637,N_2663);
nand U2796 (N_2796,N_2640,N_2636);
nor U2797 (N_2797,N_2674,N_2665);
or U2798 (N_2798,N_2620,N_2631);
or U2799 (N_2799,N_2678,N_2611);
or U2800 (N_2800,N_2702,N_2723);
and U2801 (N_2801,N_2784,N_2767);
nand U2802 (N_2802,N_2758,N_2746);
or U2803 (N_2803,N_2745,N_2782);
nand U2804 (N_2804,N_2756,N_2726);
and U2805 (N_2805,N_2793,N_2717);
nand U2806 (N_2806,N_2787,N_2710);
nor U2807 (N_2807,N_2778,N_2741);
or U2808 (N_2808,N_2754,N_2714);
and U2809 (N_2809,N_2716,N_2736);
and U2810 (N_2810,N_2762,N_2797);
or U2811 (N_2811,N_2768,N_2753);
nand U2812 (N_2812,N_2776,N_2777);
or U2813 (N_2813,N_2712,N_2780);
and U2814 (N_2814,N_2747,N_2790);
xnor U2815 (N_2815,N_2720,N_2759);
nor U2816 (N_2816,N_2722,N_2740);
and U2817 (N_2817,N_2701,N_2738);
nand U2818 (N_2818,N_2750,N_2704);
nor U2819 (N_2819,N_2772,N_2715);
or U2820 (N_2820,N_2734,N_2774);
and U2821 (N_2821,N_2733,N_2771);
xor U2822 (N_2822,N_2770,N_2783);
nand U2823 (N_2823,N_2739,N_2728);
and U2824 (N_2824,N_2708,N_2765);
or U2825 (N_2825,N_2711,N_2725);
nor U2826 (N_2826,N_2737,N_2785);
or U2827 (N_2827,N_2732,N_2744);
nor U2828 (N_2828,N_2794,N_2709);
nand U2829 (N_2829,N_2703,N_2773);
nand U2830 (N_2830,N_2775,N_2791);
nor U2831 (N_2831,N_2727,N_2721);
nor U2832 (N_2832,N_2766,N_2718);
nor U2833 (N_2833,N_2757,N_2731);
nand U2834 (N_2834,N_2706,N_2760);
nor U2835 (N_2835,N_2799,N_2789);
nand U2836 (N_2836,N_2792,N_2764);
and U2837 (N_2837,N_2713,N_2724);
nor U2838 (N_2838,N_2749,N_2761);
nand U2839 (N_2839,N_2755,N_2730);
nor U2840 (N_2840,N_2795,N_2788);
and U2841 (N_2841,N_2742,N_2796);
nand U2842 (N_2842,N_2798,N_2735);
nand U2843 (N_2843,N_2700,N_2763);
or U2844 (N_2844,N_2769,N_2748);
nand U2845 (N_2845,N_2781,N_2743);
xnor U2846 (N_2846,N_2779,N_2707);
or U2847 (N_2847,N_2705,N_2751);
xor U2848 (N_2848,N_2786,N_2719);
or U2849 (N_2849,N_2729,N_2752);
nand U2850 (N_2850,N_2790,N_2744);
and U2851 (N_2851,N_2713,N_2797);
nor U2852 (N_2852,N_2732,N_2727);
and U2853 (N_2853,N_2787,N_2703);
nor U2854 (N_2854,N_2752,N_2703);
or U2855 (N_2855,N_2701,N_2724);
nor U2856 (N_2856,N_2785,N_2715);
nand U2857 (N_2857,N_2716,N_2756);
nand U2858 (N_2858,N_2745,N_2707);
and U2859 (N_2859,N_2765,N_2700);
nand U2860 (N_2860,N_2778,N_2735);
or U2861 (N_2861,N_2785,N_2738);
and U2862 (N_2862,N_2776,N_2702);
nor U2863 (N_2863,N_2763,N_2718);
nand U2864 (N_2864,N_2794,N_2701);
and U2865 (N_2865,N_2777,N_2739);
and U2866 (N_2866,N_2783,N_2718);
nand U2867 (N_2867,N_2739,N_2796);
nand U2868 (N_2868,N_2789,N_2740);
nor U2869 (N_2869,N_2713,N_2758);
and U2870 (N_2870,N_2773,N_2796);
and U2871 (N_2871,N_2793,N_2703);
nand U2872 (N_2872,N_2751,N_2734);
or U2873 (N_2873,N_2712,N_2770);
nand U2874 (N_2874,N_2787,N_2799);
or U2875 (N_2875,N_2798,N_2737);
nor U2876 (N_2876,N_2778,N_2712);
nand U2877 (N_2877,N_2779,N_2773);
nand U2878 (N_2878,N_2734,N_2792);
nand U2879 (N_2879,N_2751,N_2748);
nor U2880 (N_2880,N_2726,N_2781);
xor U2881 (N_2881,N_2761,N_2701);
and U2882 (N_2882,N_2734,N_2767);
xnor U2883 (N_2883,N_2706,N_2765);
xor U2884 (N_2884,N_2705,N_2727);
nand U2885 (N_2885,N_2700,N_2719);
nand U2886 (N_2886,N_2727,N_2704);
or U2887 (N_2887,N_2737,N_2772);
nor U2888 (N_2888,N_2740,N_2716);
nand U2889 (N_2889,N_2766,N_2749);
nor U2890 (N_2890,N_2705,N_2788);
or U2891 (N_2891,N_2793,N_2763);
or U2892 (N_2892,N_2707,N_2737);
and U2893 (N_2893,N_2733,N_2743);
nand U2894 (N_2894,N_2717,N_2708);
nand U2895 (N_2895,N_2729,N_2799);
nor U2896 (N_2896,N_2776,N_2797);
nand U2897 (N_2897,N_2753,N_2791);
or U2898 (N_2898,N_2795,N_2728);
and U2899 (N_2899,N_2753,N_2735);
or U2900 (N_2900,N_2802,N_2868);
or U2901 (N_2901,N_2814,N_2806);
nor U2902 (N_2902,N_2895,N_2896);
nand U2903 (N_2903,N_2834,N_2811);
or U2904 (N_2904,N_2870,N_2893);
and U2905 (N_2905,N_2862,N_2854);
and U2906 (N_2906,N_2844,N_2855);
or U2907 (N_2907,N_2848,N_2866);
and U2908 (N_2908,N_2884,N_2832);
or U2909 (N_2909,N_2851,N_2826);
and U2910 (N_2910,N_2841,N_2888);
nor U2911 (N_2911,N_2894,N_2804);
and U2912 (N_2912,N_2847,N_2873);
xnor U2913 (N_2913,N_2840,N_2885);
and U2914 (N_2914,N_2861,N_2805);
nor U2915 (N_2915,N_2838,N_2882);
nor U2916 (N_2916,N_2877,N_2881);
nor U2917 (N_2917,N_2842,N_2878);
or U2918 (N_2918,N_2883,N_2887);
and U2919 (N_2919,N_2818,N_2867);
or U2920 (N_2920,N_2869,N_2850);
and U2921 (N_2921,N_2810,N_2897);
and U2922 (N_2922,N_2807,N_2821);
nor U2923 (N_2923,N_2817,N_2865);
nand U2924 (N_2924,N_2803,N_2800);
or U2925 (N_2925,N_2809,N_2875);
and U2926 (N_2926,N_2899,N_2830);
nand U2927 (N_2927,N_2843,N_2836);
nor U2928 (N_2928,N_2859,N_2879);
nand U2929 (N_2929,N_2860,N_2828);
and U2930 (N_2930,N_2833,N_2822);
and U2931 (N_2931,N_2831,N_2872);
nand U2932 (N_2932,N_2824,N_2890);
or U2933 (N_2933,N_2845,N_2876);
nand U2934 (N_2934,N_2849,N_2858);
nand U2935 (N_2935,N_2863,N_2819);
or U2936 (N_2936,N_2837,N_2839);
nand U2937 (N_2937,N_2892,N_2816);
or U2938 (N_2938,N_2846,N_2815);
nor U2939 (N_2939,N_2880,N_2857);
nor U2940 (N_2940,N_2891,N_2808);
nor U2941 (N_2941,N_2827,N_2820);
or U2942 (N_2942,N_2852,N_2898);
nor U2943 (N_2943,N_2812,N_2825);
or U2944 (N_2944,N_2829,N_2813);
or U2945 (N_2945,N_2853,N_2889);
or U2946 (N_2946,N_2835,N_2874);
nor U2947 (N_2947,N_2823,N_2871);
and U2948 (N_2948,N_2886,N_2856);
xor U2949 (N_2949,N_2864,N_2801);
and U2950 (N_2950,N_2833,N_2878);
nor U2951 (N_2951,N_2839,N_2808);
nand U2952 (N_2952,N_2865,N_2814);
nand U2953 (N_2953,N_2873,N_2820);
nor U2954 (N_2954,N_2862,N_2824);
and U2955 (N_2955,N_2856,N_2848);
and U2956 (N_2956,N_2840,N_2877);
nor U2957 (N_2957,N_2874,N_2834);
nor U2958 (N_2958,N_2831,N_2826);
and U2959 (N_2959,N_2890,N_2886);
nor U2960 (N_2960,N_2882,N_2862);
and U2961 (N_2961,N_2879,N_2849);
nor U2962 (N_2962,N_2838,N_2857);
or U2963 (N_2963,N_2847,N_2806);
or U2964 (N_2964,N_2882,N_2839);
nor U2965 (N_2965,N_2835,N_2801);
and U2966 (N_2966,N_2851,N_2828);
or U2967 (N_2967,N_2866,N_2822);
nand U2968 (N_2968,N_2878,N_2860);
nand U2969 (N_2969,N_2862,N_2884);
or U2970 (N_2970,N_2867,N_2850);
and U2971 (N_2971,N_2816,N_2821);
or U2972 (N_2972,N_2858,N_2855);
and U2973 (N_2973,N_2888,N_2866);
or U2974 (N_2974,N_2834,N_2888);
and U2975 (N_2975,N_2876,N_2827);
nor U2976 (N_2976,N_2821,N_2872);
nor U2977 (N_2977,N_2892,N_2894);
and U2978 (N_2978,N_2872,N_2829);
nand U2979 (N_2979,N_2833,N_2876);
nor U2980 (N_2980,N_2821,N_2847);
or U2981 (N_2981,N_2824,N_2843);
and U2982 (N_2982,N_2803,N_2850);
or U2983 (N_2983,N_2843,N_2890);
or U2984 (N_2984,N_2801,N_2818);
nor U2985 (N_2985,N_2837,N_2806);
or U2986 (N_2986,N_2838,N_2856);
nor U2987 (N_2987,N_2894,N_2813);
nand U2988 (N_2988,N_2898,N_2889);
nand U2989 (N_2989,N_2883,N_2833);
or U2990 (N_2990,N_2890,N_2895);
and U2991 (N_2991,N_2875,N_2808);
nand U2992 (N_2992,N_2831,N_2850);
and U2993 (N_2993,N_2837,N_2844);
and U2994 (N_2994,N_2831,N_2861);
and U2995 (N_2995,N_2878,N_2820);
nand U2996 (N_2996,N_2828,N_2807);
or U2997 (N_2997,N_2879,N_2802);
or U2998 (N_2998,N_2800,N_2831);
nand U2999 (N_2999,N_2805,N_2844);
or U3000 (N_3000,N_2901,N_2949);
and U3001 (N_3001,N_2912,N_2936);
or U3002 (N_3002,N_2937,N_2938);
and U3003 (N_3003,N_2968,N_2954);
and U3004 (N_3004,N_2984,N_2999);
or U3005 (N_3005,N_2916,N_2928);
nand U3006 (N_3006,N_2959,N_2971);
xnor U3007 (N_3007,N_2989,N_2965);
nor U3008 (N_3008,N_2947,N_2978);
and U3009 (N_3009,N_2990,N_2941);
nor U3010 (N_3010,N_2986,N_2917);
or U3011 (N_3011,N_2956,N_2930);
nor U3012 (N_3012,N_2913,N_2943);
nand U3013 (N_3013,N_2988,N_2905);
and U3014 (N_3014,N_2994,N_2972);
and U3015 (N_3015,N_2922,N_2987);
or U3016 (N_3016,N_2977,N_2973);
nand U3017 (N_3017,N_2918,N_2952);
nand U3018 (N_3018,N_2921,N_2908);
xor U3019 (N_3019,N_2926,N_2942);
nand U3020 (N_3020,N_2967,N_2909);
and U3021 (N_3021,N_2945,N_2980);
and U3022 (N_3022,N_2933,N_2904);
nand U3023 (N_3023,N_2906,N_2931);
nand U3024 (N_3024,N_2914,N_2974);
nor U3025 (N_3025,N_2979,N_2970);
nand U3026 (N_3026,N_2934,N_2935);
and U3027 (N_3027,N_2950,N_2981);
and U3028 (N_3028,N_2940,N_2927);
nor U3029 (N_3029,N_2932,N_2946);
or U3030 (N_3030,N_2944,N_2923);
and U3031 (N_3031,N_2992,N_2996);
nor U3032 (N_3032,N_2920,N_2985);
nor U3033 (N_3033,N_2948,N_2958);
nand U3034 (N_3034,N_2966,N_2907);
nand U3035 (N_3035,N_2955,N_2957);
and U3036 (N_3036,N_2925,N_2997);
and U3037 (N_3037,N_2953,N_2919);
nand U3038 (N_3038,N_2976,N_2924);
or U3039 (N_3039,N_2963,N_2975);
nor U3040 (N_3040,N_2998,N_2951);
nand U3041 (N_3041,N_2910,N_2929);
or U3042 (N_3042,N_2900,N_2903);
or U3043 (N_3043,N_2991,N_2962);
or U3044 (N_3044,N_2993,N_2983);
nand U3045 (N_3045,N_2982,N_2969);
or U3046 (N_3046,N_2995,N_2911);
nor U3047 (N_3047,N_2964,N_2939);
and U3048 (N_3048,N_2902,N_2961);
nor U3049 (N_3049,N_2960,N_2915);
nand U3050 (N_3050,N_2959,N_2926);
and U3051 (N_3051,N_2934,N_2987);
and U3052 (N_3052,N_2901,N_2914);
xnor U3053 (N_3053,N_2934,N_2962);
nor U3054 (N_3054,N_2943,N_2921);
or U3055 (N_3055,N_2944,N_2942);
or U3056 (N_3056,N_2940,N_2918);
nor U3057 (N_3057,N_2943,N_2936);
or U3058 (N_3058,N_2941,N_2907);
and U3059 (N_3059,N_2907,N_2902);
or U3060 (N_3060,N_2936,N_2993);
or U3061 (N_3061,N_2919,N_2928);
and U3062 (N_3062,N_2972,N_2979);
nand U3063 (N_3063,N_2986,N_2930);
and U3064 (N_3064,N_2917,N_2958);
nand U3065 (N_3065,N_2934,N_2919);
nand U3066 (N_3066,N_2904,N_2931);
nand U3067 (N_3067,N_2950,N_2986);
nor U3068 (N_3068,N_2920,N_2908);
and U3069 (N_3069,N_2960,N_2912);
nor U3070 (N_3070,N_2988,N_2940);
nor U3071 (N_3071,N_2915,N_2953);
nand U3072 (N_3072,N_2933,N_2950);
and U3073 (N_3073,N_2996,N_2947);
and U3074 (N_3074,N_2952,N_2944);
and U3075 (N_3075,N_2968,N_2960);
nand U3076 (N_3076,N_2948,N_2935);
and U3077 (N_3077,N_2992,N_2932);
or U3078 (N_3078,N_2954,N_2922);
and U3079 (N_3079,N_2958,N_2904);
or U3080 (N_3080,N_2956,N_2909);
nor U3081 (N_3081,N_2921,N_2971);
or U3082 (N_3082,N_2942,N_2923);
or U3083 (N_3083,N_2932,N_2976);
and U3084 (N_3084,N_2962,N_2938);
nand U3085 (N_3085,N_2932,N_2974);
nor U3086 (N_3086,N_2925,N_2911);
and U3087 (N_3087,N_2984,N_2996);
or U3088 (N_3088,N_2907,N_2965);
nand U3089 (N_3089,N_2907,N_2919);
and U3090 (N_3090,N_2950,N_2931);
nand U3091 (N_3091,N_2921,N_2949);
and U3092 (N_3092,N_2934,N_2965);
or U3093 (N_3093,N_2961,N_2978);
and U3094 (N_3094,N_2916,N_2963);
or U3095 (N_3095,N_2906,N_2905);
nand U3096 (N_3096,N_2989,N_2925);
nor U3097 (N_3097,N_2900,N_2916);
or U3098 (N_3098,N_2912,N_2977);
and U3099 (N_3099,N_2961,N_2930);
and U3100 (N_3100,N_3044,N_3006);
nor U3101 (N_3101,N_3011,N_3097);
nor U3102 (N_3102,N_3007,N_3033);
nand U3103 (N_3103,N_3080,N_3028);
nor U3104 (N_3104,N_3096,N_3057);
and U3105 (N_3105,N_3027,N_3052);
nor U3106 (N_3106,N_3072,N_3039);
xnor U3107 (N_3107,N_3064,N_3099);
nand U3108 (N_3108,N_3075,N_3013);
nand U3109 (N_3109,N_3022,N_3067);
nor U3110 (N_3110,N_3016,N_3055);
nor U3111 (N_3111,N_3050,N_3062);
and U3112 (N_3112,N_3002,N_3046);
nor U3113 (N_3113,N_3078,N_3088);
xnor U3114 (N_3114,N_3043,N_3017);
or U3115 (N_3115,N_3070,N_3024);
and U3116 (N_3116,N_3003,N_3009);
or U3117 (N_3117,N_3071,N_3091);
or U3118 (N_3118,N_3041,N_3037);
and U3119 (N_3119,N_3093,N_3004);
and U3120 (N_3120,N_3074,N_3056);
and U3121 (N_3121,N_3098,N_3069);
nor U3122 (N_3122,N_3047,N_3077);
and U3123 (N_3123,N_3026,N_3029);
and U3124 (N_3124,N_3087,N_3094);
and U3125 (N_3125,N_3073,N_3015);
and U3126 (N_3126,N_3049,N_3048);
nor U3127 (N_3127,N_3060,N_3081);
nor U3128 (N_3128,N_3051,N_3066);
or U3129 (N_3129,N_3085,N_3019);
or U3130 (N_3130,N_3021,N_3086);
nand U3131 (N_3131,N_3076,N_3010);
or U3132 (N_3132,N_3092,N_3040);
or U3133 (N_3133,N_3023,N_3045);
xor U3134 (N_3134,N_3095,N_3084);
nor U3135 (N_3135,N_3031,N_3082);
and U3136 (N_3136,N_3053,N_3000);
or U3137 (N_3137,N_3065,N_3001);
and U3138 (N_3138,N_3083,N_3089);
or U3139 (N_3139,N_3036,N_3012);
nor U3140 (N_3140,N_3032,N_3018);
or U3141 (N_3141,N_3008,N_3061);
nand U3142 (N_3142,N_3068,N_3054);
or U3143 (N_3143,N_3034,N_3038);
nor U3144 (N_3144,N_3035,N_3020);
nand U3145 (N_3145,N_3063,N_3058);
nand U3146 (N_3146,N_3014,N_3079);
xnor U3147 (N_3147,N_3025,N_3005);
and U3148 (N_3148,N_3030,N_3042);
or U3149 (N_3149,N_3090,N_3059);
xnor U3150 (N_3150,N_3009,N_3091);
nand U3151 (N_3151,N_3023,N_3085);
nor U3152 (N_3152,N_3070,N_3017);
and U3153 (N_3153,N_3045,N_3000);
nor U3154 (N_3154,N_3097,N_3019);
and U3155 (N_3155,N_3091,N_3000);
nor U3156 (N_3156,N_3033,N_3040);
and U3157 (N_3157,N_3036,N_3089);
nand U3158 (N_3158,N_3044,N_3011);
nand U3159 (N_3159,N_3016,N_3025);
xnor U3160 (N_3160,N_3000,N_3086);
nand U3161 (N_3161,N_3004,N_3075);
nor U3162 (N_3162,N_3072,N_3027);
and U3163 (N_3163,N_3043,N_3062);
or U3164 (N_3164,N_3014,N_3074);
nand U3165 (N_3165,N_3033,N_3084);
nand U3166 (N_3166,N_3045,N_3086);
nand U3167 (N_3167,N_3043,N_3071);
or U3168 (N_3168,N_3021,N_3019);
nor U3169 (N_3169,N_3084,N_3020);
and U3170 (N_3170,N_3013,N_3036);
and U3171 (N_3171,N_3073,N_3021);
or U3172 (N_3172,N_3006,N_3016);
nand U3173 (N_3173,N_3003,N_3081);
nand U3174 (N_3174,N_3077,N_3019);
or U3175 (N_3175,N_3076,N_3050);
or U3176 (N_3176,N_3013,N_3022);
or U3177 (N_3177,N_3003,N_3055);
nand U3178 (N_3178,N_3009,N_3012);
nor U3179 (N_3179,N_3099,N_3063);
or U3180 (N_3180,N_3016,N_3050);
nor U3181 (N_3181,N_3015,N_3061);
or U3182 (N_3182,N_3074,N_3071);
xnor U3183 (N_3183,N_3049,N_3014);
or U3184 (N_3184,N_3076,N_3019);
and U3185 (N_3185,N_3061,N_3078);
and U3186 (N_3186,N_3068,N_3072);
or U3187 (N_3187,N_3035,N_3009);
or U3188 (N_3188,N_3035,N_3068);
nand U3189 (N_3189,N_3072,N_3088);
nor U3190 (N_3190,N_3050,N_3032);
and U3191 (N_3191,N_3099,N_3084);
or U3192 (N_3192,N_3098,N_3024);
and U3193 (N_3193,N_3044,N_3014);
or U3194 (N_3194,N_3040,N_3032);
nor U3195 (N_3195,N_3050,N_3059);
xnor U3196 (N_3196,N_3083,N_3076);
and U3197 (N_3197,N_3030,N_3058);
nand U3198 (N_3198,N_3002,N_3071);
and U3199 (N_3199,N_3008,N_3057);
or U3200 (N_3200,N_3121,N_3127);
nor U3201 (N_3201,N_3193,N_3174);
nor U3202 (N_3202,N_3170,N_3154);
nor U3203 (N_3203,N_3119,N_3130);
nor U3204 (N_3204,N_3166,N_3195);
nor U3205 (N_3205,N_3146,N_3109);
or U3206 (N_3206,N_3138,N_3155);
or U3207 (N_3207,N_3197,N_3135);
and U3208 (N_3208,N_3117,N_3157);
nor U3209 (N_3209,N_3176,N_3141);
or U3210 (N_3210,N_3111,N_3198);
nand U3211 (N_3211,N_3100,N_3162);
and U3212 (N_3212,N_3124,N_3129);
nand U3213 (N_3213,N_3115,N_3196);
and U3214 (N_3214,N_3131,N_3172);
and U3215 (N_3215,N_3142,N_3188);
nand U3216 (N_3216,N_3156,N_3153);
nand U3217 (N_3217,N_3181,N_3136);
and U3218 (N_3218,N_3110,N_3180);
nor U3219 (N_3219,N_3160,N_3186);
nand U3220 (N_3220,N_3158,N_3149);
and U3221 (N_3221,N_3161,N_3137);
nand U3222 (N_3222,N_3125,N_3101);
or U3223 (N_3223,N_3116,N_3183);
or U3224 (N_3224,N_3102,N_3106);
or U3225 (N_3225,N_3167,N_3192);
nand U3226 (N_3226,N_3194,N_3190);
and U3227 (N_3227,N_3163,N_3189);
or U3228 (N_3228,N_3151,N_3126);
nor U3229 (N_3229,N_3148,N_3144);
or U3230 (N_3230,N_3199,N_3187);
or U3231 (N_3231,N_3128,N_3139);
or U3232 (N_3232,N_3118,N_3152);
nor U3233 (N_3233,N_3143,N_3175);
nor U3234 (N_3234,N_3140,N_3177);
or U3235 (N_3235,N_3173,N_3104);
and U3236 (N_3236,N_3191,N_3132);
or U3237 (N_3237,N_3134,N_3108);
xnor U3238 (N_3238,N_3184,N_3107);
nand U3239 (N_3239,N_3123,N_3105);
or U3240 (N_3240,N_3185,N_3114);
nand U3241 (N_3241,N_3122,N_3133);
xnor U3242 (N_3242,N_3112,N_3164);
nand U3243 (N_3243,N_3150,N_3159);
and U3244 (N_3244,N_3113,N_3168);
and U3245 (N_3245,N_3182,N_3147);
and U3246 (N_3246,N_3145,N_3169);
nor U3247 (N_3247,N_3120,N_3179);
or U3248 (N_3248,N_3171,N_3165);
and U3249 (N_3249,N_3103,N_3178);
nand U3250 (N_3250,N_3159,N_3119);
nor U3251 (N_3251,N_3123,N_3155);
nand U3252 (N_3252,N_3180,N_3137);
and U3253 (N_3253,N_3101,N_3102);
nand U3254 (N_3254,N_3137,N_3101);
and U3255 (N_3255,N_3167,N_3157);
and U3256 (N_3256,N_3160,N_3145);
and U3257 (N_3257,N_3100,N_3150);
and U3258 (N_3258,N_3141,N_3158);
or U3259 (N_3259,N_3132,N_3145);
or U3260 (N_3260,N_3181,N_3133);
nand U3261 (N_3261,N_3123,N_3138);
and U3262 (N_3262,N_3185,N_3128);
nand U3263 (N_3263,N_3190,N_3186);
nand U3264 (N_3264,N_3176,N_3108);
and U3265 (N_3265,N_3141,N_3196);
nor U3266 (N_3266,N_3169,N_3167);
or U3267 (N_3267,N_3174,N_3165);
or U3268 (N_3268,N_3128,N_3169);
or U3269 (N_3269,N_3198,N_3168);
or U3270 (N_3270,N_3142,N_3137);
and U3271 (N_3271,N_3108,N_3129);
and U3272 (N_3272,N_3109,N_3126);
and U3273 (N_3273,N_3115,N_3112);
nand U3274 (N_3274,N_3170,N_3187);
nor U3275 (N_3275,N_3104,N_3184);
and U3276 (N_3276,N_3149,N_3175);
and U3277 (N_3277,N_3119,N_3120);
or U3278 (N_3278,N_3197,N_3116);
nand U3279 (N_3279,N_3177,N_3101);
nand U3280 (N_3280,N_3128,N_3187);
nor U3281 (N_3281,N_3129,N_3183);
or U3282 (N_3282,N_3137,N_3135);
nor U3283 (N_3283,N_3166,N_3128);
nor U3284 (N_3284,N_3187,N_3132);
or U3285 (N_3285,N_3167,N_3165);
nand U3286 (N_3286,N_3158,N_3162);
nor U3287 (N_3287,N_3111,N_3108);
or U3288 (N_3288,N_3165,N_3199);
or U3289 (N_3289,N_3141,N_3133);
nor U3290 (N_3290,N_3114,N_3112);
or U3291 (N_3291,N_3115,N_3188);
or U3292 (N_3292,N_3182,N_3112);
or U3293 (N_3293,N_3153,N_3152);
or U3294 (N_3294,N_3103,N_3172);
nand U3295 (N_3295,N_3155,N_3114);
or U3296 (N_3296,N_3103,N_3110);
or U3297 (N_3297,N_3121,N_3160);
nor U3298 (N_3298,N_3160,N_3183);
nor U3299 (N_3299,N_3170,N_3102);
or U3300 (N_3300,N_3278,N_3263);
or U3301 (N_3301,N_3266,N_3290);
nor U3302 (N_3302,N_3218,N_3294);
xor U3303 (N_3303,N_3234,N_3297);
and U3304 (N_3304,N_3286,N_3272);
and U3305 (N_3305,N_3284,N_3221);
and U3306 (N_3306,N_3257,N_3204);
or U3307 (N_3307,N_3250,N_3212);
nand U3308 (N_3308,N_3267,N_3219);
or U3309 (N_3309,N_3271,N_3265);
nor U3310 (N_3310,N_3223,N_3280);
nand U3311 (N_3311,N_3296,N_3251);
nand U3312 (N_3312,N_3207,N_3247);
and U3313 (N_3313,N_3229,N_3225);
and U3314 (N_3314,N_3269,N_3201);
and U3315 (N_3315,N_3228,N_3246);
or U3316 (N_3316,N_3240,N_3277);
nand U3317 (N_3317,N_3262,N_3282);
or U3318 (N_3318,N_3205,N_3235);
or U3319 (N_3319,N_3222,N_3275);
or U3320 (N_3320,N_3230,N_3249);
and U3321 (N_3321,N_3208,N_3299);
or U3322 (N_3322,N_3264,N_3211);
and U3323 (N_3323,N_3231,N_3253);
and U3324 (N_3324,N_3281,N_3291);
nor U3325 (N_3325,N_3270,N_3226);
or U3326 (N_3326,N_3283,N_3213);
nor U3327 (N_3327,N_3239,N_3243);
nor U3328 (N_3328,N_3217,N_3214);
xor U3329 (N_3329,N_3289,N_3227);
and U3330 (N_3330,N_3287,N_3224);
nand U3331 (N_3331,N_3274,N_3242);
or U3332 (N_3332,N_3209,N_3295);
or U3333 (N_3333,N_3202,N_3260);
nand U3334 (N_3334,N_3279,N_3210);
nor U3335 (N_3335,N_3236,N_3256);
nor U3336 (N_3336,N_3293,N_3268);
and U3337 (N_3337,N_3292,N_3200);
nand U3338 (N_3338,N_3220,N_3232);
or U3339 (N_3339,N_3261,N_3233);
or U3340 (N_3340,N_3259,N_3298);
nand U3341 (N_3341,N_3254,N_3248);
and U3342 (N_3342,N_3276,N_3288);
nor U3343 (N_3343,N_3203,N_3216);
nor U3344 (N_3344,N_3206,N_3258);
nand U3345 (N_3345,N_3285,N_3244);
nor U3346 (N_3346,N_3273,N_3238);
and U3347 (N_3347,N_3252,N_3245);
and U3348 (N_3348,N_3241,N_3237);
nor U3349 (N_3349,N_3215,N_3255);
nor U3350 (N_3350,N_3210,N_3212);
nor U3351 (N_3351,N_3280,N_3272);
and U3352 (N_3352,N_3236,N_3252);
or U3353 (N_3353,N_3223,N_3281);
or U3354 (N_3354,N_3226,N_3289);
or U3355 (N_3355,N_3213,N_3264);
and U3356 (N_3356,N_3287,N_3202);
and U3357 (N_3357,N_3231,N_3202);
nor U3358 (N_3358,N_3241,N_3207);
nand U3359 (N_3359,N_3207,N_3217);
nor U3360 (N_3360,N_3297,N_3293);
nand U3361 (N_3361,N_3286,N_3239);
xnor U3362 (N_3362,N_3226,N_3256);
or U3363 (N_3363,N_3222,N_3242);
or U3364 (N_3364,N_3259,N_3263);
nor U3365 (N_3365,N_3296,N_3285);
nand U3366 (N_3366,N_3226,N_3261);
nand U3367 (N_3367,N_3288,N_3228);
and U3368 (N_3368,N_3293,N_3229);
nand U3369 (N_3369,N_3201,N_3240);
or U3370 (N_3370,N_3247,N_3219);
xnor U3371 (N_3371,N_3229,N_3291);
nand U3372 (N_3372,N_3204,N_3272);
nand U3373 (N_3373,N_3243,N_3204);
nand U3374 (N_3374,N_3250,N_3229);
nand U3375 (N_3375,N_3236,N_3244);
nor U3376 (N_3376,N_3218,N_3269);
nor U3377 (N_3377,N_3215,N_3293);
nand U3378 (N_3378,N_3278,N_3238);
nor U3379 (N_3379,N_3224,N_3275);
and U3380 (N_3380,N_3236,N_3257);
nor U3381 (N_3381,N_3281,N_3261);
nor U3382 (N_3382,N_3262,N_3211);
nor U3383 (N_3383,N_3271,N_3292);
xor U3384 (N_3384,N_3292,N_3287);
nor U3385 (N_3385,N_3286,N_3289);
or U3386 (N_3386,N_3208,N_3233);
nand U3387 (N_3387,N_3202,N_3296);
or U3388 (N_3388,N_3214,N_3229);
or U3389 (N_3389,N_3248,N_3286);
nor U3390 (N_3390,N_3249,N_3257);
nand U3391 (N_3391,N_3233,N_3292);
and U3392 (N_3392,N_3206,N_3269);
xor U3393 (N_3393,N_3270,N_3245);
nor U3394 (N_3394,N_3275,N_3260);
nand U3395 (N_3395,N_3269,N_3235);
nor U3396 (N_3396,N_3256,N_3231);
or U3397 (N_3397,N_3226,N_3201);
nor U3398 (N_3398,N_3285,N_3238);
and U3399 (N_3399,N_3293,N_3213);
xor U3400 (N_3400,N_3357,N_3343);
and U3401 (N_3401,N_3342,N_3334);
nor U3402 (N_3402,N_3373,N_3396);
and U3403 (N_3403,N_3330,N_3375);
and U3404 (N_3404,N_3335,N_3322);
nor U3405 (N_3405,N_3369,N_3350);
nand U3406 (N_3406,N_3388,N_3344);
nand U3407 (N_3407,N_3362,N_3301);
nor U3408 (N_3408,N_3337,N_3393);
and U3409 (N_3409,N_3329,N_3313);
and U3410 (N_3410,N_3399,N_3332);
nand U3411 (N_3411,N_3338,N_3394);
nor U3412 (N_3412,N_3326,N_3345);
or U3413 (N_3413,N_3351,N_3360);
nand U3414 (N_3414,N_3398,N_3300);
nor U3415 (N_3415,N_3327,N_3309);
and U3416 (N_3416,N_3307,N_3349);
nand U3417 (N_3417,N_3325,N_3318);
and U3418 (N_3418,N_3353,N_3386);
and U3419 (N_3419,N_3379,N_3319);
nor U3420 (N_3420,N_3364,N_3363);
nor U3421 (N_3421,N_3374,N_3387);
nand U3422 (N_3422,N_3352,N_3312);
and U3423 (N_3423,N_3308,N_3358);
nand U3424 (N_3424,N_3392,N_3302);
or U3425 (N_3425,N_3310,N_3315);
and U3426 (N_3426,N_3391,N_3361);
or U3427 (N_3427,N_3306,N_3382);
nand U3428 (N_3428,N_3368,N_3377);
or U3429 (N_3429,N_3381,N_3316);
nor U3430 (N_3430,N_3346,N_3339);
nor U3431 (N_3431,N_3372,N_3378);
or U3432 (N_3432,N_3367,N_3376);
nor U3433 (N_3433,N_3366,N_3321);
nor U3434 (N_3434,N_3348,N_3311);
nand U3435 (N_3435,N_3384,N_3390);
nand U3436 (N_3436,N_3324,N_3320);
and U3437 (N_3437,N_3389,N_3305);
xor U3438 (N_3438,N_3304,N_3355);
and U3439 (N_3439,N_3347,N_3340);
nor U3440 (N_3440,N_3380,N_3356);
and U3441 (N_3441,N_3385,N_3333);
nor U3442 (N_3442,N_3314,N_3323);
nor U3443 (N_3443,N_3354,N_3370);
and U3444 (N_3444,N_3397,N_3341);
nand U3445 (N_3445,N_3365,N_3359);
or U3446 (N_3446,N_3328,N_3317);
nor U3447 (N_3447,N_3336,N_3395);
nand U3448 (N_3448,N_3303,N_3383);
or U3449 (N_3449,N_3371,N_3331);
or U3450 (N_3450,N_3349,N_3369);
or U3451 (N_3451,N_3345,N_3340);
and U3452 (N_3452,N_3332,N_3368);
nor U3453 (N_3453,N_3389,N_3316);
and U3454 (N_3454,N_3312,N_3361);
and U3455 (N_3455,N_3384,N_3332);
nand U3456 (N_3456,N_3312,N_3319);
nor U3457 (N_3457,N_3380,N_3384);
nor U3458 (N_3458,N_3324,N_3360);
nor U3459 (N_3459,N_3322,N_3350);
and U3460 (N_3460,N_3344,N_3342);
and U3461 (N_3461,N_3314,N_3320);
and U3462 (N_3462,N_3348,N_3301);
nand U3463 (N_3463,N_3320,N_3399);
and U3464 (N_3464,N_3389,N_3391);
or U3465 (N_3465,N_3342,N_3319);
xnor U3466 (N_3466,N_3370,N_3338);
and U3467 (N_3467,N_3351,N_3376);
and U3468 (N_3468,N_3373,N_3365);
or U3469 (N_3469,N_3399,N_3395);
or U3470 (N_3470,N_3394,N_3346);
nor U3471 (N_3471,N_3382,N_3319);
and U3472 (N_3472,N_3317,N_3365);
nor U3473 (N_3473,N_3366,N_3352);
and U3474 (N_3474,N_3307,N_3390);
nor U3475 (N_3475,N_3321,N_3389);
and U3476 (N_3476,N_3373,N_3314);
nor U3477 (N_3477,N_3314,N_3307);
nor U3478 (N_3478,N_3363,N_3311);
nand U3479 (N_3479,N_3363,N_3314);
and U3480 (N_3480,N_3322,N_3394);
nand U3481 (N_3481,N_3355,N_3389);
nand U3482 (N_3482,N_3394,N_3365);
or U3483 (N_3483,N_3397,N_3337);
or U3484 (N_3484,N_3322,N_3315);
and U3485 (N_3485,N_3305,N_3379);
nand U3486 (N_3486,N_3325,N_3357);
nand U3487 (N_3487,N_3326,N_3340);
or U3488 (N_3488,N_3398,N_3388);
nor U3489 (N_3489,N_3396,N_3342);
or U3490 (N_3490,N_3366,N_3305);
or U3491 (N_3491,N_3359,N_3337);
or U3492 (N_3492,N_3382,N_3376);
or U3493 (N_3493,N_3350,N_3391);
or U3494 (N_3494,N_3323,N_3362);
or U3495 (N_3495,N_3313,N_3340);
and U3496 (N_3496,N_3307,N_3311);
and U3497 (N_3497,N_3378,N_3390);
or U3498 (N_3498,N_3317,N_3358);
nor U3499 (N_3499,N_3336,N_3330);
or U3500 (N_3500,N_3411,N_3487);
or U3501 (N_3501,N_3449,N_3407);
or U3502 (N_3502,N_3431,N_3496);
or U3503 (N_3503,N_3475,N_3457);
and U3504 (N_3504,N_3438,N_3460);
or U3505 (N_3505,N_3479,N_3406);
or U3506 (N_3506,N_3466,N_3491);
and U3507 (N_3507,N_3470,N_3417);
nand U3508 (N_3508,N_3430,N_3456);
nand U3509 (N_3509,N_3462,N_3489);
nor U3510 (N_3510,N_3464,N_3469);
nor U3511 (N_3511,N_3420,N_3476);
and U3512 (N_3512,N_3415,N_3447);
and U3513 (N_3513,N_3459,N_3481);
nand U3514 (N_3514,N_3403,N_3497);
nand U3515 (N_3515,N_3477,N_3445);
or U3516 (N_3516,N_3482,N_3452);
or U3517 (N_3517,N_3483,N_3427);
and U3518 (N_3518,N_3422,N_3488);
nand U3519 (N_3519,N_3424,N_3421);
or U3520 (N_3520,N_3448,N_3473);
and U3521 (N_3521,N_3468,N_3499);
nand U3522 (N_3522,N_3437,N_3478);
and U3523 (N_3523,N_3401,N_3418);
nand U3524 (N_3524,N_3455,N_3409);
or U3525 (N_3525,N_3404,N_3495);
or U3526 (N_3526,N_3485,N_3463);
or U3527 (N_3527,N_3480,N_3454);
and U3528 (N_3528,N_3474,N_3414);
or U3529 (N_3529,N_3435,N_3451);
or U3530 (N_3530,N_3472,N_3402);
and U3531 (N_3531,N_3432,N_3441);
and U3532 (N_3532,N_3494,N_3410);
xnor U3533 (N_3533,N_3498,N_3484);
and U3534 (N_3534,N_3458,N_3446);
nand U3535 (N_3535,N_3433,N_3442);
nand U3536 (N_3536,N_3416,N_3440);
nor U3537 (N_3537,N_3400,N_3493);
nand U3538 (N_3538,N_3486,N_3444);
nand U3539 (N_3539,N_3419,N_3492);
and U3540 (N_3540,N_3412,N_3436);
and U3541 (N_3541,N_3467,N_3439);
nor U3542 (N_3542,N_3434,N_3426);
nand U3543 (N_3543,N_3461,N_3465);
and U3544 (N_3544,N_3443,N_3413);
and U3545 (N_3545,N_3453,N_3425);
nand U3546 (N_3546,N_3405,N_3428);
and U3547 (N_3547,N_3471,N_3490);
or U3548 (N_3548,N_3429,N_3450);
xor U3549 (N_3549,N_3423,N_3408);
or U3550 (N_3550,N_3472,N_3465);
and U3551 (N_3551,N_3439,N_3485);
xnor U3552 (N_3552,N_3462,N_3481);
and U3553 (N_3553,N_3408,N_3411);
nor U3554 (N_3554,N_3423,N_3446);
nor U3555 (N_3555,N_3403,N_3437);
nand U3556 (N_3556,N_3409,N_3446);
or U3557 (N_3557,N_3437,N_3491);
or U3558 (N_3558,N_3400,N_3466);
nor U3559 (N_3559,N_3461,N_3430);
nand U3560 (N_3560,N_3403,N_3412);
xnor U3561 (N_3561,N_3421,N_3488);
nor U3562 (N_3562,N_3413,N_3410);
nand U3563 (N_3563,N_3454,N_3498);
nor U3564 (N_3564,N_3401,N_3403);
or U3565 (N_3565,N_3403,N_3478);
nor U3566 (N_3566,N_3490,N_3424);
nand U3567 (N_3567,N_3404,N_3484);
nor U3568 (N_3568,N_3435,N_3490);
or U3569 (N_3569,N_3438,N_3413);
or U3570 (N_3570,N_3434,N_3473);
or U3571 (N_3571,N_3498,N_3451);
nor U3572 (N_3572,N_3497,N_3434);
nor U3573 (N_3573,N_3403,N_3480);
nand U3574 (N_3574,N_3433,N_3469);
nor U3575 (N_3575,N_3497,N_3452);
nand U3576 (N_3576,N_3486,N_3448);
or U3577 (N_3577,N_3472,N_3459);
and U3578 (N_3578,N_3483,N_3456);
or U3579 (N_3579,N_3485,N_3475);
or U3580 (N_3580,N_3432,N_3468);
nand U3581 (N_3581,N_3459,N_3428);
xor U3582 (N_3582,N_3481,N_3455);
and U3583 (N_3583,N_3432,N_3497);
or U3584 (N_3584,N_3492,N_3425);
nor U3585 (N_3585,N_3463,N_3457);
or U3586 (N_3586,N_3404,N_3416);
nor U3587 (N_3587,N_3441,N_3445);
and U3588 (N_3588,N_3459,N_3471);
nand U3589 (N_3589,N_3406,N_3486);
and U3590 (N_3590,N_3455,N_3472);
and U3591 (N_3591,N_3475,N_3411);
nand U3592 (N_3592,N_3468,N_3405);
xnor U3593 (N_3593,N_3433,N_3467);
or U3594 (N_3594,N_3481,N_3493);
nor U3595 (N_3595,N_3476,N_3459);
and U3596 (N_3596,N_3471,N_3477);
or U3597 (N_3597,N_3454,N_3476);
nor U3598 (N_3598,N_3419,N_3430);
and U3599 (N_3599,N_3446,N_3400);
and U3600 (N_3600,N_3557,N_3518);
or U3601 (N_3601,N_3566,N_3539);
and U3602 (N_3602,N_3591,N_3550);
or U3603 (N_3603,N_3593,N_3582);
nor U3604 (N_3604,N_3524,N_3534);
nor U3605 (N_3605,N_3573,N_3594);
xor U3606 (N_3606,N_3576,N_3597);
nand U3607 (N_3607,N_3537,N_3586);
and U3608 (N_3608,N_3584,N_3533);
or U3609 (N_3609,N_3567,N_3569);
nand U3610 (N_3610,N_3509,N_3555);
or U3611 (N_3611,N_3577,N_3513);
nor U3612 (N_3612,N_3504,N_3536);
nand U3613 (N_3613,N_3511,N_3562);
or U3614 (N_3614,N_3581,N_3587);
nor U3615 (N_3615,N_3549,N_3522);
nand U3616 (N_3616,N_3547,N_3568);
nor U3617 (N_3617,N_3519,N_3579);
nor U3618 (N_3618,N_3528,N_3502);
nor U3619 (N_3619,N_3538,N_3510);
and U3620 (N_3620,N_3515,N_3505);
nor U3621 (N_3621,N_3598,N_3572);
nor U3622 (N_3622,N_3517,N_3527);
nor U3623 (N_3623,N_3560,N_3585);
or U3624 (N_3624,N_3595,N_3552);
nand U3625 (N_3625,N_3545,N_3574);
nand U3626 (N_3626,N_3529,N_3503);
or U3627 (N_3627,N_3575,N_3516);
nand U3628 (N_3628,N_3563,N_3551);
nand U3629 (N_3629,N_3558,N_3506);
nand U3630 (N_3630,N_3570,N_3531);
and U3631 (N_3631,N_3520,N_3530);
nor U3632 (N_3632,N_3500,N_3565);
or U3633 (N_3633,N_3512,N_3590);
nand U3634 (N_3634,N_3507,N_3501);
xor U3635 (N_3635,N_3589,N_3540);
and U3636 (N_3636,N_3541,N_3571);
nor U3637 (N_3637,N_3588,N_3542);
or U3638 (N_3638,N_3561,N_3544);
nand U3639 (N_3639,N_3508,N_3554);
or U3640 (N_3640,N_3548,N_3583);
and U3641 (N_3641,N_3526,N_3578);
xor U3642 (N_3642,N_3580,N_3556);
and U3643 (N_3643,N_3514,N_3546);
nor U3644 (N_3644,N_3564,N_3523);
or U3645 (N_3645,N_3592,N_3599);
or U3646 (N_3646,N_3596,N_3553);
nand U3647 (N_3647,N_3525,N_3559);
nor U3648 (N_3648,N_3521,N_3532);
or U3649 (N_3649,N_3543,N_3535);
and U3650 (N_3650,N_3528,N_3571);
or U3651 (N_3651,N_3533,N_3500);
xnor U3652 (N_3652,N_3518,N_3587);
and U3653 (N_3653,N_3589,N_3534);
xnor U3654 (N_3654,N_3526,N_3521);
xor U3655 (N_3655,N_3518,N_3528);
or U3656 (N_3656,N_3595,N_3572);
and U3657 (N_3657,N_3506,N_3543);
nand U3658 (N_3658,N_3555,N_3534);
nor U3659 (N_3659,N_3538,N_3543);
nor U3660 (N_3660,N_3507,N_3539);
and U3661 (N_3661,N_3526,N_3540);
or U3662 (N_3662,N_3544,N_3583);
or U3663 (N_3663,N_3505,N_3543);
and U3664 (N_3664,N_3574,N_3528);
nand U3665 (N_3665,N_3574,N_3526);
and U3666 (N_3666,N_3565,N_3521);
or U3667 (N_3667,N_3557,N_3565);
or U3668 (N_3668,N_3525,N_3566);
nand U3669 (N_3669,N_3526,N_3506);
and U3670 (N_3670,N_3521,N_3515);
nand U3671 (N_3671,N_3527,N_3570);
nor U3672 (N_3672,N_3582,N_3508);
nand U3673 (N_3673,N_3527,N_3519);
or U3674 (N_3674,N_3576,N_3556);
or U3675 (N_3675,N_3514,N_3519);
and U3676 (N_3676,N_3594,N_3563);
nor U3677 (N_3677,N_3547,N_3531);
and U3678 (N_3678,N_3555,N_3561);
and U3679 (N_3679,N_3594,N_3592);
nor U3680 (N_3680,N_3509,N_3518);
and U3681 (N_3681,N_3553,N_3507);
nand U3682 (N_3682,N_3511,N_3525);
nor U3683 (N_3683,N_3503,N_3525);
nor U3684 (N_3684,N_3500,N_3527);
or U3685 (N_3685,N_3523,N_3574);
nand U3686 (N_3686,N_3596,N_3580);
or U3687 (N_3687,N_3500,N_3545);
nand U3688 (N_3688,N_3540,N_3513);
nand U3689 (N_3689,N_3549,N_3530);
or U3690 (N_3690,N_3517,N_3518);
nand U3691 (N_3691,N_3535,N_3588);
nand U3692 (N_3692,N_3549,N_3513);
or U3693 (N_3693,N_3552,N_3583);
xnor U3694 (N_3694,N_3549,N_3543);
and U3695 (N_3695,N_3576,N_3535);
or U3696 (N_3696,N_3531,N_3541);
nand U3697 (N_3697,N_3506,N_3565);
nand U3698 (N_3698,N_3509,N_3558);
or U3699 (N_3699,N_3534,N_3532);
nor U3700 (N_3700,N_3655,N_3611);
nand U3701 (N_3701,N_3665,N_3613);
nand U3702 (N_3702,N_3685,N_3643);
or U3703 (N_3703,N_3689,N_3674);
and U3704 (N_3704,N_3607,N_3624);
nor U3705 (N_3705,N_3666,N_3630);
and U3706 (N_3706,N_3697,N_3602);
or U3707 (N_3707,N_3647,N_3629);
and U3708 (N_3708,N_3652,N_3688);
and U3709 (N_3709,N_3653,N_3641);
and U3710 (N_3710,N_3619,N_3632);
nor U3711 (N_3711,N_3622,N_3606);
or U3712 (N_3712,N_3642,N_3663);
and U3713 (N_3713,N_3637,N_3693);
and U3714 (N_3714,N_3644,N_3683);
xnor U3715 (N_3715,N_3603,N_3692);
or U3716 (N_3716,N_3612,N_3654);
nand U3717 (N_3717,N_3691,N_3680);
or U3718 (N_3718,N_3673,N_3660);
nand U3719 (N_3719,N_3690,N_3640);
and U3720 (N_3720,N_3626,N_3684);
and U3721 (N_3721,N_3604,N_3651);
or U3722 (N_3722,N_3656,N_3618);
nor U3723 (N_3723,N_3670,N_3625);
nor U3724 (N_3724,N_3600,N_3676);
or U3725 (N_3725,N_3698,N_3672);
or U3726 (N_3726,N_3609,N_3650);
nand U3727 (N_3727,N_3636,N_3679);
or U3728 (N_3728,N_3635,N_3648);
nand U3729 (N_3729,N_3617,N_3687);
or U3730 (N_3730,N_3633,N_3645);
nor U3731 (N_3731,N_3694,N_3627);
or U3732 (N_3732,N_3662,N_3659);
nand U3733 (N_3733,N_3658,N_3682);
and U3734 (N_3734,N_3649,N_3615);
nor U3735 (N_3735,N_3668,N_3699);
nor U3736 (N_3736,N_3661,N_3634);
nand U3737 (N_3737,N_3608,N_3686);
nor U3738 (N_3738,N_3621,N_3657);
and U3739 (N_3739,N_3628,N_3675);
xor U3740 (N_3740,N_3695,N_3664);
nor U3741 (N_3741,N_3677,N_3623);
or U3742 (N_3742,N_3614,N_3669);
nor U3743 (N_3743,N_3605,N_3696);
nand U3744 (N_3744,N_3646,N_3616);
nand U3745 (N_3745,N_3620,N_3631);
nor U3746 (N_3746,N_3667,N_3638);
and U3747 (N_3747,N_3671,N_3610);
or U3748 (N_3748,N_3639,N_3681);
or U3749 (N_3749,N_3678,N_3601);
nand U3750 (N_3750,N_3681,N_3695);
nand U3751 (N_3751,N_3695,N_3671);
or U3752 (N_3752,N_3626,N_3677);
nor U3753 (N_3753,N_3660,N_3691);
xnor U3754 (N_3754,N_3678,N_3633);
nor U3755 (N_3755,N_3605,N_3670);
and U3756 (N_3756,N_3668,N_3685);
or U3757 (N_3757,N_3640,N_3696);
nor U3758 (N_3758,N_3670,N_3653);
nand U3759 (N_3759,N_3692,N_3668);
or U3760 (N_3760,N_3618,N_3606);
and U3761 (N_3761,N_3682,N_3689);
or U3762 (N_3762,N_3699,N_3629);
nand U3763 (N_3763,N_3613,N_3670);
xnor U3764 (N_3764,N_3627,N_3679);
nor U3765 (N_3765,N_3643,N_3630);
nand U3766 (N_3766,N_3619,N_3688);
or U3767 (N_3767,N_3648,N_3682);
nor U3768 (N_3768,N_3666,N_3684);
nand U3769 (N_3769,N_3651,N_3689);
nor U3770 (N_3770,N_3651,N_3665);
and U3771 (N_3771,N_3666,N_3622);
and U3772 (N_3772,N_3692,N_3628);
and U3773 (N_3773,N_3611,N_3656);
nand U3774 (N_3774,N_3659,N_3624);
or U3775 (N_3775,N_3653,N_3660);
or U3776 (N_3776,N_3637,N_3669);
nor U3777 (N_3777,N_3659,N_3675);
and U3778 (N_3778,N_3640,N_3654);
nand U3779 (N_3779,N_3620,N_3658);
or U3780 (N_3780,N_3625,N_3644);
nor U3781 (N_3781,N_3641,N_3603);
nand U3782 (N_3782,N_3603,N_3670);
or U3783 (N_3783,N_3669,N_3643);
nor U3784 (N_3784,N_3649,N_3692);
or U3785 (N_3785,N_3650,N_3653);
and U3786 (N_3786,N_3617,N_3682);
nor U3787 (N_3787,N_3660,N_3605);
nor U3788 (N_3788,N_3612,N_3698);
nor U3789 (N_3789,N_3603,N_3676);
nand U3790 (N_3790,N_3692,N_3640);
and U3791 (N_3791,N_3604,N_3636);
nor U3792 (N_3792,N_3631,N_3647);
or U3793 (N_3793,N_3686,N_3606);
nand U3794 (N_3794,N_3631,N_3625);
or U3795 (N_3795,N_3636,N_3634);
nand U3796 (N_3796,N_3647,N_3627);
nand U3797 (N_3797,N_3675,N_3696);
or U3798 (N_3798,N_3633,N_3666);
or U3799 (N_3799,N_3666,N_3654);
nor U3800 (N_3800,N_3741,N_3791);
or U3801 (N_3801,N_3776,N_3746);
nand U3802 (N_3802,N_3757,N_3780);
or U3803 (N_3803,N_3785,N_3793);
or U3804 (N_3804,N_3759,N_3766);
and U3805 (N_3805,N_3720,N_3765);
nor U3806 (N_3806,N_3792,N_3799);
and U3807 (N_3807,N_3768,N_3713);
or U3808 (N_3808,N_3762,N_3706);
and U3809 (N_3809,N_3775,N_3754);
nor U3810 (N_3810,N_3726,N_3772);
and U3811 (N_3811,N_3728,N_3731);
nand U3812 (N_3812,N_3712,N_3761);
or U3813 (N_3813,N_3755,N_3794);
nand U3814 (N_3814,N_3718,N_3704);
or U3815 (N_3815,N_3739,N_3778);
nand U3816 (N_3816,N_3700,N_3748);
and U3817 (N_3817,N_3771,N_3716);
nand U3818 (N_3818,N_3742,N_3796);
or U3819 (N_3819,N_3790,N_3737);
nand U3820 (N_3820,N_3786,N_3744);
nor U3821 (N_3821,N_3701,N_3747);
and U3822 (N_3822,N_3727,N_3784);
and U3823 (N_3823,N_3715,N_3730);
and U3824 (N_3824,N_3735,N_3783);
or U3825 (N_3825,N_3752,N_3724);
nand U3826 (N_3826,N_3702,N_3769);
nand U3827 (N_3827,N_3773,N_3732);
nand U3828 (N_3828,N_3764,N_3750);
nand U3829 (N_3829,N_3745,N_3711);
or U3830 (N_3830,N_3710,N_3709);
or U3831 (N_3831,N_3777,N_3703);
nor U3832 (N_3832,N_3714,N_3722);
xor U3833 (N_3833,N_3743,N_3787);
and U3834 (N_3834,N_3749,N_3779);
or U3835 (N_3835,N_3767,N_3798);
or U3836 (N_3836,N_3795,N_3733);
and U3837 (N_3837,N_3721,N_3736);
nand U3838 (N_3838,N_3753,N_3797);
or U3839 (N_3839,N_3729,N_3763);
nor U3840 (N_3840,N_3758,N_3717);
and U3841 (N_3841,N_3734,N_3782);
nor U3842 (N_3842,N_3725,N_3788);
or U3843 (N_3843,N_3751,N_3760);
nand U3844 (N_3844,N_3740,N_3781);
and U3845 (N_3845,N_3723,N_3789);
or U3846 (N_3846,N_3770,N_3705);
nor U3847 (N_3847,N_3756,N_3738);
or U3848 (N_3848,N_3708,N_3707);
nor U3849 (N_3849,N_3774,N_3719);
xor U3850 (N_3850,N_3798,N_3725);
or U3851 (N_3851,N_3702,N_3739);
xnor U3852 (N_3852,N_3754,N_3799);
nor U3853 (N_3853,N_3726,N_3771);
and U3854 (N_3854,N_3776,N_3782);
and U3855 (N_3855,N_3733,N_3771);
or U3856 (N_3856,N_3748,N_3745);
and U3857 (N_3857,N_3726,N_3759);
nand U3858 (N_3858,N_3719,N_3733);
nor U3859 (N_3859,N_3707,N_3788);
and U3860 (N_3860,N_3754,N_3763);
or U3861 (N_3861,N_3798,N_3705);
and U3862 (N_3862,N_3766,N_3782);
nand U3863 (N_3863,N_3780,N_3771);
nor U3864 (N_3864,N_3746,N_3716);
or U3865 (N_3865,N_3765,N_3786);
nand U3866 (N_3866,N_3769,N_3772);
and U3867 (N_3867,N_3705,N_3788);
nor U3868 (N_3868,N_3783,N_3780);
xnor U3869 (N_3869,N_3736,N_3774);
and U3870 (N_3870,N_3705,N_3739);
or U3871 (N_3871,N_3721,N_3735);
xor U3872 (N_3872,N_3707,N_3790);
and U3873 (N_3873,N_3740,N_3786);
nor U3874 (N_3874,N_3721,N_3781);
nor U3875 (N_3875,N_3704,N_3770);
nor U3876 (N_3876,N_3788,N_3779);
or U3877 (N_3877,N_3705,N_3715);
and U3878 (N_3878,N_3716,N_3769);
nand U3879 (N_3879,N_3739,N_3720);
or U3880 (N_3880,N_3716,N_3777);
and U3881 (N_3881,N_3708,N_3739);
and U3882 (N_3882,N_3758,N_3724);
or U3883 (N_3883,N_3757,N_3717);
and U3884 (N_3884,N_3783,N_3777);
or U3885 (N_3885,N_3722,N_3701);
nor U3886 (N_3886,N_3764,N_3727);
nor U3887 (N_3887,N_3780,N_3749);
nand U3888 (N_3888,N_3711,N_3707);
nor U3889 (N_3889,N_3752,N_3740);
nand U3890 (N_3890,N_3742,N_3728);
or U3891 (N_3891,N_3725,N_3746);
or U3892 (N_3892,N_3738,N_3732);
nor U3893 (N_3893,N_3752,N_3793);
xnor U3894 (N_3894,N_3740,N_3767);
nand U3895 (N_3895,N_3705,N_3777);
nor U3896 (N_3896,N_3793,N_3722);
nor U3897 (N_3897,N_3780,N_3750);
or U3898 (N_3898,N_3790,N_3772);
and U3899 (N_3899,N_3774,N_3712);
nand U3900 (N_3900,N_3807,N_3850);
nor U3901 (N_3901,N_3846,N_3878);
xnor U3902 (N_3902,N_3854,N_3837);
nand U3903 (N_3903,N_3864,N_3826);
and U3904 (N_3904,N_3832,N_3882);
and U3905 (N_3905,N_3816,N_3872);
nor U3906 (N_3906,N_3802,N_3842);
nand U3907 (N_3907,N_3843,N_3862);
nand U3908 (N_3908,N_3830,N_3890);
and U3909 (N_3909,N_3818,N_3841);
and U3910 (N_3910,N_3800,N_3883);
and U3911 (N_3911,N_3803,N_3819);
nor U3912 (N_3912,N_3861,N_3860);
nand U3913 (N_3913,N_3899,N_3814);
and U3914 (N_3914,N_3879,N_3829);
or U3915 (N_3915,N_3884,N_3891);
nand U3916 (N_3916,N_3893,N_3871);
nor U3917 (N_3917,N_3885,N_3853);
and U3918 (N_3918,N_3876,N_3895);
nand U3919 (N_3919,N_3867,N_3805);
nand U3920 (N_3920,N_3809,N_3849);
nor U3921 (N_3921,N_3851,N_3886);
and U3922 (N_3922,N_3855,N_3844);
nor U3923 (N_3923,N_3875,N_3823);
or U3924 (N_3924,N_3866,N_3827);
or U3925 (N_3925,N_3859,N_3894);
or U3926 (N_3926,N_3856,N_3847);
nand U3927 (N_3927,N_3887,N_3820);
nor U3928 (N_3928,N_3801,N_3865);
and U3929 (N_3929,N_3881,N_3812);
nand U3930 (N_3930,N_3840,N_3833);
nand U3931 (N_3931,N_3821,N_3868);
nor U3932 (N_3932,N_3835,N_3870);
nand U3933 (N_3933,N_3845,N_3880);
nand U3934 (N_3934,N_3858,N_3811);
or U3935 (N_3935,N_3808,N_3806);
nor U3936 (N_3936,N_3834,N_3825);
nor U3937 (N_3937,N_3813,N_3831);
or U3938 (N_3938,N_3863,N_3848);
nand U3939 (N_3939,N_3836,N_3817);
nor U3940 (N_3940,N_3839,N_3869);
or U3941 (N_3941,N_3877,N_3824);
nand U3942 (N_3942,N_3873,N_3828);
or U3943 (N_3943,N_3898,N_3852);
nand U3944 (N_3944,N_3897,N_3804);
nor U3945 (N_3945,N_3810,N_3822);
nand U3946 (N_3946,N_3896,N_3892);
and U3947 (N_3947,N_3857,N_3838);
nand U3948 (N_3948,N_3815,N_3888);
nor U3949 (N_3949,N_3889,N_3874);
nand U3950 (N_3950,N_3815,N_3891);
nor U3951 (N_3951,N_3873,N_3860);
nor U3952 (N_3952,N_3875,N_3836);
nand U3953 (N_3953,N_3858,N_3842);
and U3954 (N_3954,N_3836,N_3893);
nand U3955 (N_3955,N_3857,N_3861);
nand U3956 (N_3956,N_3866,N_3847);
and U3957 (N_3957,N_3824,N_3849);
or U3958 (N_3958,N_3899,N_3805);
nand U3959 (N_3959,N_3804,N_3872);
xnor U3960 (N_3960,N_3868,N_3831);
nand U3961 (N_3961,N_3880,N_3868);
nor U3962 (N_3962,N_3894,N_3847);
nor U3963 (N_3963,N_3830,N_3827);
and U3964 (N_3964,N_3894,N_3834);
nor U3965 (N_3965,N_3857,N_3843);
and U3966 (N_3966,N_3825,N_3869);
or U3967 (N_3967,N_3819,N_3875);
nand U3968 (N_3968,N_3860,N_3882);
and U3969 (N_3969,N_3816,N_3835);
nor U3970 (N_3970,N_3859,N_3885);
nand U3971 (N_3971,N_3874,N_3822);
or U3972 (N_3972,N_3859,N_3823);
nand U3973 (N_3973,N_3813,N_3817);
nor U3974 (N_3974,N_3816,N_3866);
and U3975 (N_3975,N_3801,N_3877);
nand U3976 (N_3976,N_3807,N_3877);
and U3977 (N_3977,N_3826,N_3816);
nor U3978 (N_3978,N_3860,N_3887);
and U3979 (N_3979,N_3815,N_3889);
or U3980 (N_3980,N_3846,N_3850);
nor U3981 (N_3981,N_3875,N_3814);
and U3982 (N_3982,N_3841,N_3829);
nand U3983 (N_3983,N_3899,N_3850);
nand U3984 (N_3984,N_3814,N_3829);
xnor U3985 (N_3985,N_3854,N_3897);
or U3986 (N_3986,N_3862,N_3885);
and U3987 (N_3987,N_3875,N_3884);
or U3988 (N_3988,N_3811,N_3882);
nor U3989 (N_3989,N_3896,N_3862);
or U3990 (N_3990,N_3891,N_3883);
nor U3991 (N_3991,N_3826,N_3869);
nor U3992 (N_3992,N_3837,N_3817);
and U3993 (N_3993,N_3836,N_3843);
and U3994 (N_3994,N_3813,N_3819);
nor U3995 (N_3995,N_3870,N_3859);
nand U3996 (N_3996,N_3857,N_3816);
nand U3997 (N_3997,N_3831,N_3884);
nand U3998 (N_3998,N_3865,N_3869);
nor U3999 (N_3999,N_3818,N_3800);
nor U4000 (N_4000,N_3918,N_3911);
xnor U4001 (N_4001,N_3930,N_3981);
nor U4002 (N_4002,N_3990,N_3970);
nand U4003 (N_4003,N_3914,N_3982);
and U4004 (N_4004,N_3905,N_3935);
nand U4005 (N_4005,N_3973,N_3975);
and U4006 (N_4006,N_3902,N_3932);
xor U4007 (N_4007,N_3972,N_3934);
and U4008 (N_4008,N_3931,N_3910);
nor U4009 (N_4009,N_3995,N_3950);
nand U4010 (N_4010,N_3998,N_3985);
nor U4011 (N_4011,N_3925,N_3923);
and U4012 (N_4012,N_3957,N_3958);
nand U4013 (N_4013,N_3920,N_3922);
nand U4014 (N_4014,N_3913,N_3983);
or U4015 (N_4015,N_3954,N_3936);
and U4016 (N_4016,N_3939,N_3933);
or U4017 (N_4017,N_3976,N_3959);
nand U4018 (N_4018,N_3900,N_3997);
nor U4019 (N_4019,N_3961,N_3974);
nor U4020 (N_4020,N_3915,N_3901);
xnor U4021 (N_4021,N_3952,N_3989);
nor U4022 (N_4022,N_3907,N_3908);
nand U4023 (N_4023,N_3948,N_3945);
nand U4024 (N_4024,N_3946,N_3926);
and U4025 (N_4025,N_3979,N_3964);
nand U4026 (N_4026,N_3924,N_3978);
nor U4027 (N_4027,N_3969,N_3992);
nor U4028 (N_4028,N_3944,N_3971);
or U4029 (N_4029,N_3965,N_3993);
or U4030 (N_4030,N_3919,N_3916);
nand U4031 (N_4031,N_3951,N_3904);
or U4032 (N_4032,N_3962,N_3968);
nand U4033 (N_4033,N_3940,N_3938);
or U4034 (N_4034,N_3955,N_3980);
or U4035 (N_4035,N_3949,N_3999);
nor U4036 (N_4036,N_3953,N_3917);
nand U4037 (N_4037,N_3909,N_3986);
and U4038 (N_4038,N_3960,N_3977);
and U4039 (N_4039,N_3927,N_3988);
nor U4040 (N_4040,N_3921,N_3996);
or U4041 (N_4041,N_3906,N_3963);
and U4042 (N_4042,N_3991,N_3956);
or U4043 (N_4043,N_3937,N_3912);
or U4044 (N_4044,N_3987,N_3941);
or U4045 (N_4045,N_3966,N_3928);
or U4046 (N_4046,N_3929,N_3967);
or U4047 (N_4047,N_3903,N_3984);
and U4048 (N_4048,N_3947,N_3943);
nand U4049 (N_4049,N_3942,N_3994);
nor U4050 (N_4050,N_3946,N_3971);
nand U4051 (N_4051,N_3971,N_3909);
nor U4052 (N_4052,N_3972,N_3973);
nand U4053 (N_4053,N_3963,N_3903);
and U4054 (N_4054,N_3982,N_3918);
nor U4055 (N_4055,N_3956,N_3982);
nand U4056 (N_4056,N_3983,N_3991);
or U4057 (N_4057,N_3989,N_3964);
nand U4058 (N_4058,N_3976,N_3905);
nor U4059 (N_4059,N_3986,N_3994);
nor U4060 (N_4060,N_3941,N_3993);
or U4061 (N_4061,N_3932,N_3935);
nor U4062 (N_4062,N_3920,N_3936);
nor U4063 (N_4063,N_3991,N_3900);
nand U4064 (N_4064,N_3907,N_3985);
nand U4065 (N_4065,N_3937,N_3908);
or U4066 (N_4066,N_3980,N_3923);
and U4067 (N_4067,N_3905,N_3995);
nand U4068 (N_4068,N_3900,N_3977);
and U4069 (N_4069,N_3979,N_3950);
and U4070 (N_4070,N_3988,N_3938);
or U4071 (N_4071,N_3978,N_3988);
and U4072 (N_4072,N_3983,N_3952);
nor U4073 (N_4073,N_3975,N_3998);
nand U4074 (N_4074,N_3912,N_3963);
nand U4075 (N_4075,N_3994,N_3945);
nor U4076 (N_4076,N_3988,N_3976);
nand U4077 (N_4077,N_3964,N_3901);
and U4078 (N_4078,N_3999,N_3935);
and U4079 (N_4079,N_3972,N_3949);
or U4080 (N_4080,N_3948,N_3923);
and U4081 (N_4081,N_3987,N_3984);
nor U4082 (N_4082,N_3941,N_3999);
nand U4083 (N_4083,N_3956,N_3955);
nand U4084 (N_4084,N_3932,N_3982);
nand U4085 (N_4085,N_3961,N_3971);
nor U4086 (N_4086,N_3904,N_3949);
nand U4087 (N_4087,N_3916,N_3912);
nor U4088 (N_4088,N_3910,N_3953);
and U4089 (N_4089,N_3954,N_3955);
and U4090 (N_4090,N_3917,N_3933);
or U4091 (N_4091,N_3960,N_3917);
and U4092 (N_4092,N_3943,N_3988);
and U4093 (N_4093,N_3921,N_3909);
or U4094 (N_4094,N_3917,N_3926);
and U4095 (N_4095,N_3981,N_3937);
and U4096 (N_4096,N_3967,N_3959);
and U4097 (N_4097,N_3987,N_3959);
and U4098 (N_4098,N_3972,N_3918);
or U4099 (N_4099,N_3965,N_3967);
nand U4100 (N_4100,N_4040,N_4093);
or U4101 (N_4101,N_4052,N_4066);
or U4102 (N_4102,N_4073,N_4071);
nand U4103 (N_4103,N_4046,N_4023);
nor U4104 (N_4104,N_4090,N_4053);
nor U4105 (N_4105,N_4038,N_4014);
or U4106 (N_4106,N_4056,N_4069);
nor U4107 (N_4107,N_4029,N_4003);
or U4108 (N_4108,N_4076,N_4041);
nor U4109 (N_4109,N_4062,N_4086);
and U4110 (N_4110,N_4009,N_4010);
and U4111 (N_4111,N_4055,N_4022);
and U4112 (N_4112,N_4048,N_4008);
and U4113 (N_4113,N_4002,N_4015);
and U4114 (N_4114,N_4001,N_4005);
and U4115 (N_4115,N_4063,N_4039);
nor U4116 (N_4116,N_4070,N_4077);
nor U4117 (N_4117,N_4037,N_4017);
and U4118 (N_4118,N_4047,N_4020);
xor U4119 (N_4119,N_4024,N_4072);
nand U4120 (N_4120,N_4075,N_4049);
nor U4121 (N_4121,N_4012,N_4030);
and U4122 (N_4122,N_4021,N_4064);
xor U4123 (N_4123,N_4054,N_4057);
and U4124 (N_4124,N_4016,N_4067);
and U4125 (N_4125,N_4081,N_4096);
or U4126 (N_4126,N_4036,N_4099);
or U4127 (N_4127,N_4044,N_4061);
and U4128 (N_4128,N_4098,N_4051);
and U4129 (N_4129,N_4042,N_4043);
nand U4130 (N_4130,N_4013,N_4019);
nand U4131 (N_4131,N_4089,N_4034);
xor U4132 (N_4132,N_4027,N_4079);
nor U4133 (N_4133,N_4088,N_4065);
and U4134 (N_4134,N_4060,N_4035);
or U4135 (N_4135,N_4080,N_4006);
and U4136 (N_4136,N_4094,N_4082);
nand U4137 (N_4137,N_4026,N_4059);
or U4138 (N_4138,N_4031,N_4025);
nand U4139 (N_4139,N_4095,N_4028);
or U4140 (N_4140,N_4084,N_4032);
nor U4141 (N_4141,N_4068,N_4091);
nand U4142 (N_4142,N_4074,N_4050);
and U4143 (N_4143,N_4033,N_4000);
nand U4144 (N_4144,N_4018,N_4083);
and U4145 (N_4145,N_4097,N_4045);
nor U4146 (N_4146,N_4011,N_4004);
and U4147 (N_4147,N_4007,N_4078);
or U4148 (N_4148,N_4092,N_4087);
or U4149 (N_4149,N_4085,N_4058);
and U4150 (N_4150,N_4009,N_4039);
xnor U4151 (N_4151,N_4060,N_4022);
or U4152 (N_4152,N_4010,N_4089);
nand U4153 (N_4153,N_4030,N_4003);
or U4154 (N_4154,N_4055,N_4042);
or U4155 (N_4155,N_4075,N_4044);
or U4156 (N_4156,N_4033,N_4087);
or U4157 (N_4157,N_4096,N_4061);
nor U4158 (N_4158,N_4083,N_4071);
or U4159 (N_4159,N_4038,N_4080);
or U4160 (N_4160,N_4015,N_4035);
or U4161 (N_4161,N_4080,N_4068);
and U4162 (N_4162,N_4017,N_4064);
and U4163 (N_4163,N_4016,N_4008);
nand U4164 (N_4164,N_4038,N_4033);
nor U4165 (N_4165,N_4038,N_4070);
nand U4166 (N_4166,N_4054,N_4008);
or U4167 (N_4167,N_4022,N_4039);
or U4168 (N_4168,N_4000,N_4020);
nand U4169 (N_4169,N_4012,N_4043);
or U4170 (N_4170,N_4021,N_4080);
nor U4171 (N_4171,N_4082,N_4057);
xnor U4172 (N_4172,N_4068,N_4095);
nand U4173 (N_4173,N_4022,N_4083);
or U4174 (N_4174,N_4042,N_4077);
or U4175 (N_4175,N_4059,N_4018);
nor U4176 (N_4176,N_4049,N_4063);
nor U4177 (N_4177,N_4042,N_4050);
nor U4178 (N_4178,N_4065,N_4091);
nor U4179 (N_4179,N_4072,N_4029);
and U4180 (N_4180,N_4098,N_4032);
or U4181 (N_4181,N_4058,N_4012);
or U4182 (N_4182,N_4061,N_4064);
and U4183 (N_4183,N_4031,N_4043);
and U4184 (N_4184,N_4070,N_4074);
nor U4185 (N_4185,N_4022,N_4077);
or U4186 (N_4186,N_4001,N_4097);
and U4187 (N_4187,N_4052,N_4017);
or U4188 (N_4188,N_4081,N_4097);
and U4189 (N_4189,N_4072,N_4004);
and U4190 (N_4190,N_4017,N_4018);
or U4191 (N_4191,N_4040,N_4089);
nand U4192 (N_4192,N_4026,N_4039);
or U4193 (N_4193,N_4044,N_4085);
nand U4194 (N_4194,N_4094,N_4056);
and U4195 (N_4195,N_4010,N_4019);
nor U4196 (N_4196,N_4013,N_4009);
nand U4197 (N_4197,N_4028,N_4057);
nor U4198 (N_4198,N_4018,N_4028);
nor U4199 (N_4199,N_4039,N_4034);
or U4200 (N_4200,N_4169,N_4147);
nand U4201 (N_4201,N_4131,N_4181);
nor U4202 (N_4202,N_4106,N_4178);
and U4203 (N_4203,N_4197,N_4188);
xnor U4204 (N_4204,N_4149,N_4150);
and U4205 (N_4205,N_4133,N_4153);
nor U4206 (N_4206,N_4179,N_4192);
nand U4207 (N_4207,N_4164,N_4154);
nor U4208 (N_4208,N_4165,N_4196);
nand U4209 (N_4209,N_4142,N_4171);
nand U4210 (N_4210,N_4114,N_4173);
and U4211 (N_4211,N_4140,N_4117);
xor U4212 (N_4212,N_4107,N_4199);
and U4213 (N_4213,N_4110,N_4104);
and U4214 (N_4214,N_4146,N_4198);
nor U4215 (N_4215,N_4136,N_4183);
nor U4216 (N_4216,N_4134,N_4162);
and U4217 (N_4217,N_4159,N_4151);
and U4218 (N_4218,N_4130,N_4176);
or U4219 (N_4219,N_4109,N_4184);
nor U4220 (N_4220,N_4124,N_4121);
or U4221 (N_4221,N_4128,N_4115);
or U4222 (N_4222,N_4119,N_4158);
nand U4223 (N_4223,N_4108,N_4135);
nand U4224 (N_4224,N_4141,N_4143);
nand U4225 (N_4225,N_4116,N_4191);
or U4226 (N_4226,N_4144,N_4170);
nand U4227 (N_4227,N_4102,N_4195);
or U4228 (N_4228,N_4139,N_4182);
nor U4229 (N_4229,N_4156,N_4100);
and U4230 (N_4230,N_4137,N_4145);
and U4231 (N_4231,N_4163,N_4155);
nand U4232 (N_4232,N_4148,N_4129);
nor U4233 (N_4233,N_4193,N_4185);
nor U4234 (N_4234,N_4123,N_4132);
and U4235 (N_4235,N_4167,N_4186);
nand U4236 (N_4236,N_4161,N_4103);
and U4237 (N_4237,N_4112,N_4180);
or U4238 (N_4238,N_4152,N_4111);
and U4239 (N_4239,N_4172,N_4190);
and U4240 (N_4240,N_4105,N_4127);
nand U4241 (N_4241,N_4118,N_4125);
nand U4242 (N_4242,N_4174,N_4175);
and U4243 (N_4243,N_4177,N_4189);
and U4244 (N_4244,N_4101,N_4138);
nor U4245 (N_4245,N_4160,N_4120);
nor U4246 (N_4246,N_4157,N_4126);
or U4247 (N_4247,N_4166,N_4122);
or U4248 (N_4248,N_4113,N_4168);
or U4249 (N_4249,N_4187,N_4194);
and U4250 (N_4250,N_4156,N_4109);
and U4251 (N_4251,N_4199,N_4138);
nor U4252 (N_4252,N_4170,N_4161);
nand U4253 (N_4253,N_4187,N_4198);
nor U4254 (N_4254,N_4129,N_4106);
or U4255 (N_4255,N_4126,N_4152);
and U4256 (N_4256,N_4154,N_4156);
xnor U4257 (N_4257,N_4115,N_4143);
nand U4258 (N_4258,N_4148,N_4167);
or U4259 (N_4259,N_4173,N_4186);
and U4260 (N_4260,N_4116,N_4137);
or U4261 (N_4261,N_4131,N_4172);
nor U4262 (N_4262,N_4192,N_4170);
nor U4263 (N_4263,N_4167,N_4118);
and U4264 (N_4264,N_4101,N_4175);
or U4265 (N_4265,N_4180,N_4121);
or U4266 (N_4266,N_4134,N_4168);
nand U4267 (N_4267,N_4195,N_4144);
nor U4268 (N_4268,N_4199,N_4148);
nor U4269 (N_4269,N_4123,N_4174);
nand U4270 (N_4270,N_4132,N_4137);
and U4271 (N_4271,N_4152,N_4108);
nand U4272 (N_4272,N_4117,N_4122);
and U4273 (N_4273,N_4192,N_4152);
nor U4274 (N_4274,N_4148,N_4116);
nand U4275 (N_4275,N_4115,N_4145);
nor U4276 (N_4276,N_4117,N_4183);
and U4277 (N_4277,N_4118,N_4142);
and U4278 (N_4278,N_4175,N_4162);
and U4279 (N_4279,N_4119,N_4137);
or U4280 (N_4280,N_4175,N_4186);
nor U4281 (N_4281,N_4117,N_4139);
or U4282 (N_4282,N_4146,N_4140);
nor U4283 (N_4283,N_4143,N_4178);
nor U4284 (N_4284,N_4143,N_4109);
nand U4285 (N_4285,N_4129,N_4157);
nand U4286 (N_4286,N_4170,N_4118);
nor U4287 (N_4287,N_4100,N_4182);
nor U4288 (N_4288,N_4159,N_4134);
or U4289 (N_4289,N_4103,N_4157);
or U4290 (N_4290,N_4194,N_4152);
nand U4291 (N_4291,N_4127,N_4139);
and U4292 (N_4292,N_4110,N_4154);
nand U4293 (N_4293,N_4133,N_4169);
or U4294 (N_4294,N_4167,N_4195);
nor U4295 (N_4295,N_4194,N_4100);
and U4296 (N_4296,N_4138,N_4126);
nand U4297 (N_4297,N_4188,N_4199);
nand U4298 (N_4298,N_4144,N_4167);
nand U4299 (N_4299,N_4153,N_4188);
and U4300 (N_4300,N_4227,N_4269);
and U4301 (N_4301,N_4206,N_4288);
nand U4302 (N_4302,N_4281,N_4221);
nor U4303 (N_4303,N_4202,N_4267);
nor U4304 (N_4304,N_4296,N_4223);
and U4305 (N_4305,N_4253,N_4271);
and U4306 (N_4306,N_4239,N_4265);
nand U4307 (N_4307,N_4278,N_4252);
or U4308 (N_4308,N_4220,N_4273);
or U4309 (N_4309,N_4216,N_4204);
or U4310 (N_4310,N_4236,N_4240);
and U4311 (N_4311,N_4270,N_4233);
and U4312 (N_4312,N_4285,N_4277);
and U4313 (N_4313,N_4209,N_4243);
and U4314 (N_4314,N_4222,N_4207);
and U4315 (N_4315,N_4213,N_4257);
and U4316 (N_4316,N_4231,N_4200);
and U4317 (N_4317,N_4228,N_4266);
nor U4318 (N_4318,N_4234,N_4298);
and U4319 (N_4319,N_4217,N_4259);
nor U4320 (N_4320,N_4274,N_4290);
nor U4321 (N_4321,N_4294,N_4201);
xor U4322 (N_4322,N_4255,N_4275);
and U4323 (N_4323,N_4284,N_4247);
and U4324 (N_4324,N_4235,N_4250);
nor U4325 (N_4325,N_4293,N_4276);
nor U4326 (N_4326,N_4242,N_4289);
or U4327 (N_4327,N_4268,N_4219);
xor U4328 (N_4328,N_4226,N_4264);
nor U4329 (N_4329,N_4272,N_4212);
or U4330 (N_4330,N_4232,N_4299);
and U4331 (N_4331,N_4297,N_4210);
and U4332 (N_4332,N_4229,N_4291);
nor U4333 (N_4333,N_4237,N_4287);
and U4334 (N_4334,N_4279,N_4224);
and U4335 (N_4335,N_4214,N_4292);
nand U4336 (N_4336,N_4225,N_4286);
nand U4337 (N_4337,N_4215,N_4263);
nor U4338 (N_4338,N_4254,N_4249);
or U4339 (N_4339,N_4258,N_4248);
nor U4340 (N_4340,N_4260,N_4218);
nor U4341 (N_4341,N_4280,N_4211);
nand U4342 (N_4342,N_4205,N_4241);
nor U4343 (N_4343,N_4295,N_4245);
nor U4344 (N_4344,N_4246,N_4244);
or U4345 (N_4345,N_4261,N_4283);
or U4346 (N_4346,N_4282,N_4230);
xor U4347 (N_4347,N_4238,N_4203);
or U4348 (N_4348,N_4208,N_4262);
or U4349 (N_4349,N_4251,N_4256);
and U4350 (N_4350,N_4229,N_4211);
nand U4351 (N_4351,N_4244,N_4211);
nand U4352 (N_4352,N_4237,N_4259);
nand U4353 (N_4353,N_4240,N_4241);
nand U4354 (N_4354,N_4259,N_4265);
or U4355 (N_4355,N_4270,N_4260);
nand U4356 (N_4356,N_4281,N_4204);
or U4357 (N_4357,N_4268,N_4295);
nand U4358 (N_4358,N_4296,N_4228);
xnor U4359 (N_4359,N_4216,N_4247);
or U4360 (N_4360,N_4278,N_4253);
or U4361 (N_4361,N_4268,N_4262);
nor U4362 (N_4362,N_4277,N_4226);
nand U4363 (N_4363,N_4226,N_4201);
nand U4364 (N_4364,N_4278,N_4237);
nand U4365 (N_4365,N_4229,N_4216);
xor U4366 (N_4366,N_4249,N_4216);
nand U4367 (N_4367,N_4249,N_4250);
and U4368 (N_4368,N_4209,N_4266);
or U4369 (N_4369,N_4253,N_4273);
or U4370 (N_4370,N_4268,N_4227);
nand U4371 (N_4371,N_4283,N_4218);
and U4372 (N_4372,N_4262,N_4299);
and U4373 (N_4373,N_4271,N_4297);
and U4374 (N_4374,N_4291,N_4212);
nand U4375 (N_4375,N_4295,N_4251);
or U4376 (N_4376,N_4289,N_4215);
nor U4377 (N_4377,N_4239,N_4219);
nor U4378 (N_4378,N_4277,N_4214);
xnor U4379 (N_4379,N_4265,N_4209);
nor U4380 (N_4380,N_4201,N_4238);
nand U4381 (N_4381,N_4241,N_4211);
nand U4382 (N_4382,N_4208,N_4236);
nand U4383 (N_4383,N_4293,N_4288);
nor U4384 (N_4384,N_4232,N_4268);
and U4385 (N_4385,N_4289,N_4253);
or U4386 (N_4386,N_4200,N_4286);
nand U4387 (N_4387,N_4290,N_4254);
or U4388 (N_4388,N_4271,N_4269);
nor U4389 (N_4389,N_4284,N_4282);
nand U4390 (N_4390,N_4261,N_4250);
and U4391 (N_4391,N_4281,N_4226);
nand U4392 (N_4392,N_4211,N_4297);
xnor U4393 (N_4393,N_4240,N_4261);
or U4394 (N_4394,N_4278,N_4283);
or U4395 (N_4395,N_4267,N_4298);
or U4396 (N_4396,N_4240,N_4204);
and U4397 (N_4397,N_4258,N_4282);
xor U4398 (N_4398,N_4295,N_4267);
or U4399 (N_4399,N_4282,N_4227);
or U4400 (N_4400,N_4357,N_4326);
and U4401 (N_4401,N_4308,N_4321);
or U4402 (N_4402,N_4358,N_4328);
nand U4403 (N_4403,N_4397,N_4349);
or U4404 (N_4404,N_4355,N_4341);
nand U4405 (N_4405,N_4320,N_4359);
or U4406 (N_4406,N_4324,N_4390);
and U4407 (N_4407,N_4368,N_4374);
nand U4408 (N_4408,N_4330,N_4337);
nand U4409 (N_4409,N_4301,N_4360);
or U4410 (N_4410,N_4365,N_4392);
or U4411 (N_4411,N_4316,N_4396);
or U4412 (N_4412,N_4312,N_4347);
and U4413 (N_4413,N_4344,N_4303);
or U4414 (N_4414,N_4319,N_4313);
and U4415 (N_4415,N_4348,N_4354);
or U4416 (N_4416,N_4352,N_4332);
and U4417 (N_4417,N_4329,N_4309);
nor U4418 (N_4418,N_4371,N_4399);
nor U4419 (N_4419,N_4336,N_4323);
nand U4420 (N_4420,N_4388,N_4381);
nand U4421 (N_4421,N_4318,N_4373);
or U4422 (N_4422,N_4379,N_4331);
or U4423 (N_4423,N_4366,N_4395);
nand U4424 (N_4424,N_4361,N_4302);
and U4425 (N_4425,N_4300,N_4322);
nand U4426 (N_4426,N_4377,N_4315);
and U4427 (N_4427,N_4380,N_4398);
nor U4428 (N_4428,N_4353,N_4370);
or U4429 (N_4429,N_4369,N_4306);
nand U4430 (N_4430,N_4317,N_4351);
or U4431 (N_4431,N_4376,N_4334);
nand U4432 (N_4432,N_4372,N_4333);
and U4433 (N_4433,N_4384,N_4375);
nor U4434 (N_4434,N_4304,N_4342);
nand U4435 (N_4435,N_4356,N_4394);
nand U4436 (N_4436,N_4378,N_4346);
and U4437 (N_4437,N_4314,N_4382);
or U4438 (N_4438,N_4386,N_4364);
nor U4439 (N_4439,N_4367,N_4305);
xnor U4440 (N_4440,N_4310,N_4338);
and U4441 (N_4441,N_4335,N_4325);
nor U4442 (N_4442,N_4363,N_4385);
and U4443 (N_4443,N_4391,N_4327);
and U4444 (N_4444,N_4389,N_4343);
and U4445 (N_4445,N_4311,N_4383);
and U4446 (N_4446,N_4387,N_4307);
nand U4447 (N_4447,N_4345,N_4339);
and U4448 (N_4448,N_4362,N_4340);
nor U4449 (N_4449,N_4393,N_4350);
and U4450 (N_4450,N_4311,N_4398);
or U4451 (N_4451,N_4371,N_4340);
nor U4452 (N_4452,N_4316,N_4388);
or U4453 (N_4453,N_4315,N_4352);
or U4454 (N_4454,N_4361,N_4313);
and U4455 (N_4455,N_4365,N_4389);
nor U4456 (N_4456,N_4302,N_4385);
nor U4457 (N_4457,N_4314,N_4374);
nand U4458 (N_4458,N_4309,N_4375);
or U4459 (N_4459,N_4390,N_4351);
or U4460 (N_4460,N_4369,N_4312);
and U4461 (N_4461,N_4361,N_4392);
xor U4462 (N_4462,N_4337,N_4359);
and U4463 (N_4463,N_4331,N_4334);
nand U4464 (N_4464,N_4337,N_4377);
nand U4465 (N_4465,N_4363,N_4309);
and U4466 (N_4466,N_4385,N_4318);
nor U4467 (N_4467,N_4321,N_4345);
nor U4468 (N_4468,N_4340,N_4389);
or U4469 (N_4469,N_4311,N_4301);
nor U4470 (N_4470,N_4393,N_4355);
and U4471 (N_4471,N_4321,N_4355);
or U4472 (N_4472,N_4330,N_4361);
nand U4473 (N_4473,N_4338,N_4359);
or U4474 (N_4474,N_4368,N_4339);
or U4475 (N_4475,N_4339,N_4393);
and U4476 (N_4476,N_4368,N_4388);
and U4477 (N_4477,N_4391,N_4336);
and U4478 (N_4478,N_4361,N_4337);
nor U4479 (N_4479,N_4301,N_4357);
or U4480 (N_4480,N_4389,N_4330);
nor U4481 (N_4481,N_4360,N_4368);
nand U4482 (N_4482,N_4311,N_4305);
or U4483 (N_4483,N_4380,N_4373);
nand U4484 (N_4484,N_4303,N_4385);
nand U4485 (N_4485,N_4396,N_4398);
nor U4486 (N_4486,N_4312,N_4308);
and U4487 (N_4487,N_4322,N_4343);
nand U4488 (N_4488,N_4313,N_4312);
nor U4489 (N_4489,N_4372,N_4362);
nor U4490 (N_4490,N_4376,N_4328);
or U4491 (N_4491,N_4319,N_4378);
nand U4492 (N_4492,N_4393,N_4301);
nor U4493 (N_4493,N_4335,N_4383);
or U4494 (N_4494,N_4302,N_4382);
nand U4495 (N_4495,N_4337,N_4345);
and U4496 (N_4496,N_4391,N_4366);
nor U4497 (N_4497,N_4393,N_4352);
or U4498 (N_4498,N_4371,N_4327);
nand U4499 (N_4499,N_4337,N_4375);
and U4500 (N_4500,N_4400,N_4486);
and U4501 (N_4501,N_4441,N_4411);
and U4502 (N_4502,N_4448,N_4439);
and U4503 (N_4503,N_4407,N_4481);
nand U4504 (N_4504,N_4424,N_4416);
or U4505 (N_4505,N_4467,N_4432);
nand U4506 (N_4506,N_4446,N_4456);
nor U4507 (N_4507,N_4468,N_4488);
nor U4508 (N_4508,N_4415,N_4443);
or U4509 (N_4509,N_4451,N_4427);
nand U4510 (N_4510,N_4401,N_4408);
and U4511 (N_4511,N_4466,N_4460);
nor U4512 (N_4512,N_4483,N_4413);
or U4513 (N_4513,N_4462,N_4428);
nand U4514 (N_4514,N_4426,N_4435);
or U4515 (N_4515,N_4499,N_4492);
xor U4516 (N_4516,N_4497,N_4459);
nand U4517 (N_4517,N_4417,N_4404);
nor U4518 (N_4518,N_4493,N_4473);
and U4519 (N_4519,N_4457,N_4423);
or U4520 (N_4520,N_4494,N_4490);
and U4521 (N_4521,N_4429,N_4447);
or U4522 (N_4522,N_4498,N_4496);
nor U4523 (N_4523,N_4461,N_4470);
xor U4524 (N_4524,N_4484,N_4440);
or U4525 (N_4525,N_4458,N_4438);
nor U4526 (N_4526,N_4479,N_4478);
and U4527 (N_4527,N_4454,N_4422);
or U4528 (N_4528,N_4482,N_4465);
and U4529 (N_4529,N_4410,N_4449);
xor U4530 (N_4530,N_4476,N_4434);
or U4531 (N_4531,N_4444,N_4491);
and U4532 (N_4532,N_4433,N_4477);
or U4533 (N_4533,N_4412,N_4431);
nor U4534 (N_4534,N_4437,N_4430);
nor U4535 (N_4535,N_4487,N_4474);
nor U4536 (N_4536,N_4419,N_4420);
nand U4537 (N_4537,N_4414,N_4469);
or U4538 (N_4538,N_4442,N_4418);
nor U4539 (N_4539,N_4485,N_4489);
nand U4540 (N_4540,N_4421,N_4403);
nor U4541 (N_4541,N_4475,N_4463);
nand U4542 (N_4542,N_4406,N_4471);
or U4543 (N_4543,N_4464,N_4453);
or U4544 (N_4544,N_4495,N_4452);
nor U4545 (N_4545,N_4480,N_4436);
or U4546 (N_4546,N_4425,N_4405);
xor U4547 (N_4547,N_4409,N_4472);
nor U4548 (N_4548,N_4455,N_4450);
or U4549 (N_4549,N_4402,N_4445);
nor U4550 (N_4550,N_4456,N_4431);
nand U4551 (N_4551,N_4428,N_4497);
or U4552 (N_4552,N_4432,N_4449);
or U4553 (N_4553,N_4484,N_4427);
and U4554 (N_4554,N_4455,N_4494);
and U4555 (N_4555,N_4493,N_4418);
and U4556 (N_4556,N_4407,N_4429);
or U4557 (N_4557,N_4400,N_4407);
and U4558 (N_4558,N_4451,N_4433);
xnor U4559 (N_4559,N_4442,N_4496);
and U4560 (N_4560,N_4413,N_4450);
and U4561 (N_4561,N_4401,N_4466);
nand U4562 (N_4562,N_4461,N_4413);
nor U4563 (N_4563,N_4400,N_4498);
nand U4564 (N_4564,N_4482,N_4425);
nand U4565 (N_4565,N_4418,N_4497);
and U4566 (N_4566,N_4413,N_4442);
and U4567 (N_4567,N_4452,N_4474);
or U4568 (N_4568,N_4461,N_4468);
nand U4569 (N_4569,N_4485,N_4435);
or U4570 (N_4570,N_4473,N_4471);
and U4571 (N_4571,N_4437,N_4405);
nor U4572 (N_4572,N_4435,N_4491);
xor U4573 (N_4573,N_4407,N_4435);
or U4574 (N_4574,N_4466,N_4475);
nand U4575 (N_4575,N_4440,N_4481);
and U4576 (N_4576,N_4432,N_4469);
nor U4577 (N_4577,N_4424,N_4455);
or U4578 (N_4578,N_4406,N_4475);
xor U4579 (N_4579,N_4408,N_4429);
nand U4580 (N_4580,N_4484,N_4435);
or U4581 (N_4581,N_4472,N_4470);
nor U4582 (N_4582,N_4454,N_4493);
or U4583 (N_4583,N_4464,N_4416);
and U4584 (N_4584,N_4429,N_4485);
or U4585 (N_4585,N_4438,N_4498);
and U4586 (N_4586,N_4420,N_4499);
nor U4587 (N_4587,N_4474,N_4475);
and U4588 (N_4588,N_4481,N_4459);
or U4589 (N_4589,N_4414,N_4466);
and U4590 (N_4590,N_4488,N_4453);
nand U4591 (N_4591,N_4479,N_4410);
and U4592 (N_4592,N_4448,N_4475);
nor U4593 (N_4593,N_4457,N_4452);
nor U4594 (N_4594,N_4464,N_4460);
or U4595 (N_4595,N_4448,N_4460);
nor U4596 (N_4596,N_4475,N_4433);
and U4597 (N_4597,N_4424,N_4482);
nor U4598 (N_4598,N_4478,N_4423);
nand U4599 (N_4599,N_4491,N_4436);
xor U4600 (N_4600,N_4506,N_4591);
nand U4601 (N_4601,N_4583,N_4530);
nand U4602 (N_4602,N_4540,N_4502);
nor U4603 (N_4603,N_4545,N_4590);
nor U4604 (N_4604,N_4539,N_4543);
nor U4605 (N_4605,N_4531,N_4579);
xnor U4606 (N_4606,N_4598,N_4524);
and U4607 (N_4607,N_4589,N_4554);
nand U4608 (N_4608,N_4534,N_4525);
nand U4609 (N_4609,N_4535,N_4552);
nor U4610 (N_4610,N_4510,N_4527);
nor U4611 (N_4611,N_4551,N_4520);
nand U4612 (N_4612,N_4567,N_4526);
nor U4613 (N_4613,N_4599,N_4562);
or U4614 (N_4614,N_4528,N_4582);
nand U4615 (N_4615,N_4558,N_4574);
and U4616 (N_4616,N_4503,N_4593);
nand U4617 (N_4617,N_4594,N_4577);
nand U4618 (N_4618,N_4521,N_4553);
xnor U4619 (N_4619,N_4519,N_4573);
nand U4620 (N_4620,N_4513,N_4565);
nor U4621 (N_4621,N_4536,N_4585);
nand U4622 (N_4622,N_4550,N_4570);
and U4623 (N_4623,N_4507,N_4548);
nand U4624 (N_4624,N_4508,N_4597);
or U4625 (N_4625,N_4557,N_4563);
nand U4626 (N_4626,N_4547,N_4511);
xor U4627 (N_4627,N_4549,N_4501);
xor U4628 (N_4628,N_4556,N_4564);
and U4629 (N_4629,N_4587,N_4537);
nand U4630 (N_4630,N_4571,N_4514);
and U4631 (N_4631,N_4505,N_4575);
nor U4632 (N_4632,N_4578,N_4588);
or U4633 (N_4633,N_4566,N_4584);
and U4634 (N_4634,N_4572,N_4561);
nor U4635 (N_4635,N_4569,N_4560);
and U4636 (N_4636,N_4586,N_4529);
or U4637 (N_4637,N_4580,N_4518);
xor U4638 (N_4638,N_4533,N_4576);
or U4639 (N_4639,N_4542,N_4541);
nor U4640 (N_4640,N_4500,N_4546);
nand U4641 (N_4641,N_4555,N_4568);
nand U4642 (N_4642,N_4596,N_4516);
xor U4643 (N_4643,N_4532,N_4504);
and U4644 (N_4644,N_4515,N_4595);
and U4645 (N_4645,N_4559,N_4544);
and U4646 (N_4646,N_4592,N_4509);
and U4647 (N_4647,N_4522,N_4538);
or U4648 (N_4648,N_4517,N_4512);
and U4649 (N_4649,N_4523,N_4581);
nand U4650 (N_4650,N_4503,N_4562);
xnor U4651 (N_4651,N_4553,N_4505);
or U4652 (N_4652,N_4511,N_4522);
nor U4653 (N_4653,N_4559,N_4569);
or U4654 (N_4654,N_4518,N_4595);
nor U4655 (N_4655,N_4558,N_4592);
nor U4656 (N_4656,N_4559,N_4598);
nand U4657 (N_4657,N_4556,N_4516);
xnor U4658 (N_4658,N_4525,N_4559);
or U4659 (N_4659,N_4537,N_4524);
nand U4660 (N_4660,N_4596,N_4574);
and U4661 (N_4661,N_4556,N_4536);
and U4662 (N_4662,N_4520,N_4578);
and U4663 (N_4663,N_4591,N_4568);
xnor U4664 (N_4664,N_4559,N_4585);
and U4665 (N_4665,N_4544,N_4556);
or U4666 (N_4666,N_4539,N_4589);
or U4667 (N_4667,N_4550,N_4540);
or U4668 (N_4668,N_4563,N_4533);
nand U4669 (N_4669,N_4570,N_4567);
nor U4670 (N_4670,N_4591,N_4530);
nor U4671 (N_4671,N_4589,N_4599);
nor U4672 (N_4672,N_4507,N_4523);
or U4673 (N_4673,N_4589,N_4565);
and U4674 (N_4674,N_4557,N_4555);
or U4675 (N_4675,N_4567,N_4572);
xnor U4676 (N_4676,N_4547,N_4509);
or U4677 (N_4677,N_4509,N_4541);
nand U4678 (N_4678,N_4584,N_4546);
nand U4679 (N_4679,N_4562,N_4546);
or U4680 (N_4680,N_4541,N_4508);
or U4681 (N_4681,N_4513,N_4503);
nor U4682 (N_4682,N_4508,N_4580);
nand U4683 (N_4683,N_4551,N_4585);
and U4684 (N_4684,N_4560,N_4518);
or U4685 (N_4685,N_4536,N_4500);
nor U4686 (N_4686,N_4564,N_4577);
nand U4687 (N_4687,N_4586,N_4510);
nor U4688 (N_4688,N_4518,N_4503);
xor U4689 (N_4689,N_4576,N_4503);
or U4690 (N_4690,N_4595,N_4516);
and U4691 (N_4691,N_4569,N_4543);
or U4692 (N_4692,N_4539,N_4553);
nand U4693 (N_4693,N_4574,N_4519);
or U4694 (N_4694,N_4513,N_4575);
or U4695 (N_4695,N_4551,N_4558);
nand U4696 (N_4696,N_4550,N_4531);
nand U4697 (N_4697,N_4538,N_4515);
or U4698 (N_4698,N_4529,N_4531);
or U4699 (N_4699,N_4560,N_4567);
and U4700 (N_4700,N_4648,N_4644);
nor U4701 (N_4701,N_4616,N_4647);
nor U4702 (N_4702,N_4641,N_4623);
or U4703 (N_4703,N_4687,N_4668);
and U4704 (N_4704,N_4629,N_4696);
or U4705 (N_4705,N_4626,N_4652);
nor U4706 (N_4706,N_4637,N_4628);
or U4707 (N_4707,N_4638,N_4615);
nand U4708 (N_4708,N_4610,N_4646);
or U4709 (N_4709,N_4600,N_4620);
or U4710 (N_4710,N_4653,N_4667);
and U4711 (N_4711,N_4654,N_4657);
and U4712 (N_4712,N_4606,N_4672);
nor U4713 (N_4713,N_4660,N_4614);
and U4714 (N_4714,N_4692,N_4686);
or U4715 (N_4715,N_4642,N_4697);
nor U4716 (N_4716,N_4619,N_4608);
nor U4717 (N_4717,N_4694,N_4607);
nand U4718 (N_4718,N_4604,N_4664);
or U4719 (N_4719,N_4679,N_4680);
nor U4720 (N_4720,N_4681,N_4689);
and U4721 (N_4721,N_4601,N_4633);
nor U4722 (N_4722,N_4693,N_4675);
and U4723 (N_4723,N_4656,N_4632);
or U4724 (N_4724,N_4695,N_4645);
nor U4725 (N_4725,N_4682,N_4662);
nor U4726 (N_4726,N_4661,N_4613);
nand U4727 (N_4727,N_4627,N_4677);
or U4728 (N_4728,N_4678,N_4636);
nor U4729 (N_4729,N_4665,N_4618);
and U4730 (N_4730,N_4649,N_4666);
nand U4731 (N_4731,N_4691,N_4658);
nand U4732 (N_4732,N_4617,N_4625);
and U4733 (N_4733,N_4651,N_4685);
xor U4734 (N_4734,N_4688,N_4684);
and U4735 (N_4735,N_4622,N_4624);
nand U4736 (N_4736,N_4609,N_4640);
nand U4737 (N_4737,N_4630,N_4643);
or U4738 (N_4738,N_4655,N_4650);
xor U4739 (N_4739,N_4635,N_4683);
nor U4740 (N_4740,N_4690,N_4631);
nand U4741 (N_4741,N_4602,N_4670);
or U4742 (N_4742,N_4639,N_4698);
nor U4743 (N_4743,N_4674,N_4605);
and U4744 (N_4744,N_4611,N_4673);
nor U4745 (N_4745,N_4659,N_4669);
and U4746 (N_4746,N_4671,N_4612);
or U4747 (N_4747,N_4603,N_4663);
or U4748 (N_4748,N_4621,N_4699);
and U4749 (N_4749,N_4676,N_4634);
nor U4750 (N_4750,N_4697,N_4670);
nand U4751 (N_4751,N_4622,N_4614);
xnor U4752 (N_4752,N_4647,N_4691);
nand U4753 (N_4753,N_4666,N_4623);
or U4754 (N_4754,N_4653,N_4662);
and U4755 (N_4755,N_4664,N_4655);
or U4756 (N_4756,N_4659,N_4601);
nor U4757 (N_4757,N_4607,N_4677);
or U4758 (N_4758,N_4660,N_4687);
nor U4759 (N_4759,N_4664,N_4690);
nor U4760 (N_4760,N_4659,N_4620);
nor U4761 (N_4761,N_4655,N_4682);
or U4762 (N_4762,N_4669,N_4618);
or U4763 (N_4763,N_4612,N_4620);
nand U4764 (N_4764,N_4682,N_4642);
or U4765 (N_4765,N_4656,N_4603);
nand U4766 (N_4766,N_4671,N_4660);
or U4767 (N_4767,N_4629,N_4603);
nand U4768 (N_4768,N_4667,N_4617);
and U4769 (N_4769,N_4627,N_4679);
or U4770 (N_4770,N_4687,N_4691);
nand U4771 (N_4771,N_4698,N_4603);
and U4772 (N_4772,N_4692,N_4697);
and U4773 (N_4773,N_4619,N_4688);
nand U4774 (N_4774,N_4684,N_4617);
nand U4775 (N_4775,N_4608,N_4642);
nor U4776 (N_4776,N_4627,N_4629);
or U4777 (N_4777,N_4627,N_4683);
and U4778 (N_4778,N_4699,N_4656);
nor U4779 (N_4779,N_4603,N_4606);
or U4780 (N_4780,N_4682,N_4647);
nor U4781 (N_4781,N_4618,N_4625);
and U4782 (N_4782,N_4634,N_4604);
nor U4783 (N_4783,N_4640,N_4661);
nand U4784 (N_4784,N_4664,N_4678);
nand U4785 (N_4785,N_4672,N_4633);
or U4786 (N_4786,N_4693,N_4671);
or U4787 (N_4787,N_4651,N_4648);
nor U4788 (N_4788,N_4669,N_4613);
and U4789 (N_4789,N_4655,N_4672);
nor U4790 (N_4790,N_4637,N_4677);
or U4791 (N_4791,N_4630,N_4647);
nor U4792 (N_4792,N_4645,N_4671);
or U4793 (N_4793,N_4681,N_4628);
nor U4794 (N_4794,N_4663,N_4614);
nor U4795 (N_4795,N_4630,N_4661);
nor U4796 (N_4796,N_4697,N_4601);
nand U4797 (N_4797,N_4652,N_4619);
or U4798 (N_4798,N_4658,N_4651);
nand U4799 (N_4799,N_4661,N_4632);
or U4800 (N_4800,N_4751,N_4740);
and U4801 (N_4801,N_4772,N_4715);
and U4802 (N_4802,N_4789,N_4744);
nor U4803 (N_4803,N_4756,N_4734);
nand U4804 (N_4804,N_4735,N_4764);
nand U4805 (N_4805,N_4749,N_4785);
nor U4806 (N_4806,N_4758,N_4717);
and U4807 (N_4807,N_4729,N_4709);
nor U4808 (N_4808,N_4700,N_4760);
and U4809 (N_4809,N_4798,N_4712);
or U4810 (N_4810,N_4786,N_4790);
nor U4811 (N_4811,N_4723,N_4728);
and U4812 (N_4812,N_4788,N_4784);
nor U4813 (N_4813,N_4707,N_4776);
xor U4814 (N_4814,N_4799,N_4763);
or U4815 (N_4815,N_4741,N_4701);
and U4816 (N_4816,N_4752,N_4710);
xor U4817 (N_4817,N_4721,N_4738);
or U4818 (N_4818,N_4725,N_4711);
nor U4819 (N_4819,N_4783,N_4742);
nor U4820 (N_4820,N_4761,N_4743);
and U4821 (N_4821,N_4718,N_4765);
or U4822 (N_4822,N_4705,N_4755);
nand U4823 (N_4823,N_4708,N_4753);
nand U4824 (N_4824,N_4793,N_4766);
or U4825 (N_4825,N_4754,N_4792);
nand U4826 (N_4826,N_4716,N_4770);
nor U4827 (N_4827,N_4722,N_4778);
nand U4828 (N_4828,N_4724,N_4732);
nand U4829 (N_4829,N_4791,N_4787);
and U4830 (N_4830,N_4703,N_4794);
nand U4831 (N_4831,N_4714,N_4777);
nand U4832 (N_4832,N_4713,N_4737);
and U4833 (N_4833,N_4773,N_4733);
nor U4834 (N_4834,N_4750,N_4747);
nand U4835 (N_4835,N_4731,N_4762);
nor U4836 (N_4836,N_4782,N_4727);
nand U4837 (N_4837,N_4774,N_4736);
nand U4838 (N_4838,N_4795,N_4771);
and U4839 (N_4839,N_4726,N_4781);
nand U4840 (N_4840,N_4779,N_4757);
and U4841 (N_4841,N_4768,N_4759);
nor U4842 (N_4842,N_4704,N_4780);
and U4843 (N_4843,N_4796,N_4748);
or U4844 (N_4844,N_4719,N_4797);
or U4845 (N_4845,N_4775,N_4720);
and U4846 (N_4846,N_4746,N_4745);
and U4847 (N_4847,N_4739,N_4769);
and U4848 (N_4848,N_4702,N_4730);
and U4849 (N_4849,N_4706,N_4767);
or U4850 (N_4850,N_4743,N_4780);
nand U4851 (N_4851,N_4708,N_4752);
nand U4852 (N_4852,N_4794,N_4723);
and U4853 (N_4853,N_4747,N_4703);
or U4854 (N_4854,N_4778,N_4792);
nor U4855 (N_4855,N_4769,N_4711);
or U4856 (N_4856,N_4706,N_4781);
or U4857 (N_4857,N_4791,N_4740);
nor U4858 (N_4858,N_4701,N_4784);
nor U4859 (N_4859,N_4799,N_4748);
nor U4860 (N_4860,N_4762,N_4724);
and U4861 (N_4861,N_4757,N_4710);
nand U4862 (N_4862,N_4708,N_4793);
nor U4863 (N_4863,N_4704,N_4795);
or U4864 (N_4864,N_4765,N_4773);
and U4865 (N_4865,N_4751,N_4712);
or U4866 (N_4866,N_4732,N_4799);
xnor U4867 (N_4867,N_4775,N_4791);
nand U4868 (N_4868,N_4797,N_4750);
and U4869 (N_4869,N_4770,N_4769);
and U4870 (N_4870,N_4716,N_4765);
and U4871 (N_4871,N_4717,N_4735);
nand U4872 (N_4872,N_4789,N_4735);
nor U4873 (N_4873,N_4792,N_4726);
nand U4874 (N_4874,N_4738,N_4743);
nand U4875 (N_4875,N_4779,N_4758);
and U4876 (N_4876,N_4740,N_4745);
nor U4877 (N_4877,N_4736,N_4767);
or U4878 (N_4878,N_4776,N_4720);
nand U4879 (N_4879,N_4728,N_4781);
and U4880 (N_4880,N_4772,N_4775);
and U4881 (N_4881,N_4724,N_4766);
nor U4882 (N_4882,N_4790,N_4795);
and U4883 (N_4883,N_4773,N_4722);
and U4884 (N_4884,N_4739,N_4797);
nand U4885 (N_4885,N_4772,N_4709);
or U4886 (N_4886,N_4720,N_4730);
nand U4887 (N_4887,N_4732,N_4793);
nand U4888 (N_4888,N_4778,N_4795);
or U4889 (N_4889,N_4782,N_4771);
or U4890 (N_4890,N_4739,N_4718);
and U4891 (N_4891,N_4793,N_4745);
or U4892 (N_4892,N_4756,N_4778);
and U4893 (N_4893,N_4792,N_4795);
nor U4894 (N_4894,N_4766,N_4722);
or U4895 (N_4895,N_4704,N_4755);
nor U4896 (N_4896,N_4798,N_4779);
nand U4897 (N_4897,N_4780,N_4784);
nand U4898 (N_4898,N_4752,N_4788);
nand U4899 (N_4899,N_4702,N_4780);
and U4900 (N_4900,N_4839,N_4864);
nand U4901 (N_4901,N_4898,N_4804);
and U4902 (N_4902,N_4896,N_4833);
and U4903 (N_4903,N_4815,N_4892);
and U4904 (N_4904,N_4811,N_4840);
nor U4905 (N_4905,N_4865,N_4825);
and U4906 (N_4906,N_4843,N_4879);
or U4907 (N_4907,N_4818,N_4871);
or U4908 (N_4908,N_4822,N_4841);
and U4909 (N_4909,N_4828,N_4893);
or U4910 (N_4910,N_4881,N_4860);
or U4911 (N_4911,N_4829,N_4854);
and U4912 (N_4912,N_4848,N_4886);
nor U4913 (N_4913,N_4890,N_4847);
or U4914 (N_4914,N_4810,N_4888);
nor U4915 (N_4915,N_4866,N_4801);
or U4916 (N_4916,N_4883,N_4884);
nand U4917 (N_4917,N_4856,N_4846);
or U4918 (N_4918,N_4823,N_4838);
xor U4919 (N_4919,N_4869,N_4874);
or U4920 (N_4920,N_4835,N_4813);
nor U4921 (N_4921,N_4859,N_4819);
nand U4922 (N_4922,N_4891,N_4895);
or U4923 (N_4923,N_4873,N_4803);
and U4924 (N_4924,N_4831,N_4816);
or U4925 (N_4925,N_4844,N_4867);
and U4926 (N_4926,N_4832,N_4876);
or U4927 (N_4927,N_4849,N_4870);
nor U4928 (N_4928,N_4889,N_4855);
xor U4929 (N_4929,N_4836,N_4830);
nand U4930 (N_4930,N_4897,N_4880);
or U4931 (N_4931,N_4807,N_4894);
nand U4932 (N_4932,N_4845,N_4887);
nand U4933 (N_4933,N_4800,N_4885);
or U4934 (N_4934,N_4899,N_4802);
or U4935 (N_4935,N_4826,N_4878);
nand U4936 (N_4936,N_4820,N_4857);
nor U4937 (N_4937,N_4805,N_4824);
and U4938 (N_4938,N_4850,N_4875);
nor U4939 (N_4939,N_4863,N_4834);
and U4940 (N_4940,N_4817,N_4877);
nand U4941 (N_4941,N_4851,N_4858);
or U4942 (N_4942,N_4852,N_4842);
and U4943 (N_4943,N_4812,N_4868);
nand U4944 (N_4944,N_4861,N_4821);
or U4945 (N_4945,N_4862,N_4827);
and U4946 (N_4946,N_4853,N_4837);
nor U4947 (N_4947,N_4882,N_4808);
nand U4948 (N_4948,N_4814,N_4809);
nor U4949 (N_4949,N_4872,N_4806);
or U4950 (N_4950,N_4803,N_4880);
nand U4951 (N_4951,N_4859,N_4896);
or U4952 (N_4952,N_4885,N_4832);
or U4953 (N_4953,N_4854,N_4817);
nor U4954 (N_4954,N_4898,N_4842);
or U4955 (N_4955,N_4859,N_4857);
or U4956 (N_4956,N_4818,N_4841);
nand U4957 (N_4957,N_4828,N_4855);
nand U4958 (N_4958,N_4825,N_4885);
nand U4959 (N_4959,N_4806,N_4824);
nand U4960 (N_4960,N_4825,N_4802);
and U4961 (N_4961,N_4832,N_4869);
and U4962 (N_4962,N_4841,N_4880);
or U4963 (N_4963,N_4819,N_4824);
and U4964 (N_4964,N_4816,N_4844);
nor U4965 (N_4965,N_4845,N_4867);
nor U4966 (N_4966,N_4853,N_4805);
nor U4967 (N_4967,N_4891,N_4873);
nor U4968 (N_4968,N_4875,N_4878);
nor U4969 (N_4969,N_4811,N_4894);
nand U4970 (N_4970,N_4884,N_4877);
nor U4971 (N_4971,N_4897,N_4895);
xnor U4972 (N_4972,N_4830,N_4813);
nand U4973 (N_4973,N_4872,N_4837);
nand U4974 (N_4974,N_4869,N_4807);
and U4975 (N_4975,N_4819,N_4805);
nor U4976 (N_4976,N_4869,N_4889);
and U4977 (N_4977,N_4832,N_4878);
nand U4978 (N_4978,N_4875,N_4893);
nand U4979 (N_4979,N_4836,N_4868);
nand U4980 (N_4980,N_4890,N_4882);
or U4981 (N_4981,N_4864,N_4855);
or U4982 (N_4982,N_4889,N_4805);
and U4983 (N_4983,N_4810,N_4804);
nand U4984 (N_4984,N_4851,N_4841);
or U4985 (N_4985,N_4802,N_4856);
nor U4986 (N_4986,N_4892,N_4890);
and U4987 (N_4987,N_4814,N_4803);
or U4988 (N_4988,N_4898,N_4893);
xnor U4989 (N_4989,N_4853,N_4871);
nand U4990 (N_4990,N_4875,N_4887);
nor U4991 (N_4991,N_4899,N_4807);
or U4992 (N_4992,N_4892,N_4851);
xnor U4993 (N_4993,N_4829,N_4848);
and U4994 (N_4994,N_4835,N_4832);
xor U4995 (N_4995,N_4895,N_4875);
nor U4996 (N_4996,N_4879,N_4889);
or U4997 (N_4997,N_4815,N_4860);
and U4998 (N_4998,N_4896,N_4846);
or U4999 (N_4999,N_4845,N_4882);
and UO_0 (O_0,N_4959,N_4988);
nand UO_1 (O_1,N_4998,N_4960);
or UO_2 (O_2,N_4964,N_4987);
or UO_3 (O_3,N_4949,N_4996);
nor UO_4 (O_4,N_4989,N_4900);
nor UO_5 (O_5,N_4983,N_4945);
nand UO_6 (O_6,N_4923,N_4934);
nand UO_7 (O_7,N_4980,N_4997);
and UO_8 (O_8,N_4995,N_4990);
nor UO_9 (O_9,N_4924,N_4971);
and UO_10 (O_10,N_4912,N_4955);
nand UO_11 (O_11,N_4985,N_4919);
nor UO_12 (O_12,N_4941,N_4931);
nor UO_13 (O_13,N_4940,N_4921);
and UO_14 (O_14,N_4975,N_4984);
and UO_15 (O_15,N_4942,N_4993);
and UO_16 (O_16,N_4968,N_4939);
nand UO_17 (O_17,N_4927,N_4992);
nand UO_18 (O_18,N_4925,N_4906);
nor UO_19 (O_19,N_4963,N_4946);
nor UO_20 (O_20,N_4937,N_4977);
or UO_21 (O_21,N_4933,N_4928);
nor UO_22 (O_22,N_4974,N_4994);
nand UO_23 (O_23,N_4972,N_4967);
nand UO_24 (O_24,N_4978,N_4999);
nand UO_25 (O_25,N_4961,N_4904);
nand UO_26 (O_26,N_4944,N_4991);
and UO_27 (O_27,N_4910,N_4929);
nand UO_28 (O_28,N_4905,N_4950);
nand UO_29 (O_29,N_4966,N_4951);
nand UO_30 (O_30,N_4920,N_4947);
or UO_31 (O_31,N_4953,N_4957);
nand UO_32 (O_32,N_4901,N_4982);
nand UO_33 (O_33,N_4918,N_4943);
nor UO_34 (O_34,N_4962,N_4916);
nand UO_35 (O_35,N_4902,N_4970);
or UO_36 (O_36,N_4903,N_4958);
nor UO_37 (O_37,N_4915,N_4979);
xnor UO_38 (O_38,N_4917,N_4936);
nand UO_39 (O_39,N_4969,N_4954);
xnor UO_40 (O_40,N_4926,N_4911);
nand UO_41 (O_41,N_4976,N_4922);
nand UO_42 (O_42,N_4952,N_4938);
nor UO_43 (O_43,N_4930,N_4956);
or UO_44 (O_44,N_4935,N_4986);
or UO_45 (O_45,N_4981,N_4907);
and UO_46 (O_46,N_4948,N_4932);
and UO_47 (O_47,N_4914,N_4908);
nor UO_48 (O_48,N_4965,N_4973);
or UO_49 (O_49,N_4913,N_4909);
nand UO_50 (O_50,N_4961,N_4990);
nand UO_51 (O_51,N_4930,N_4915);
and UO_52 (O_52,N_4949,N_4913);
nor UO_53 (O_53,N_4986,N_4977);
or UO_54 (O_54,N_4947,N_4949);
and UO_55 (O_55,N_4934,N_4986);
nand UO_56 (O_56,N_4913,N_4932);
and UO_57 (O_57,N_4968,N_4911);
or UO_58 (O_58,N_4924,N_4969);
nor UO_59 (O_59,N_4930,N_4924);
or UO_60 (O_60,N_4907,N_4992);
nand UO_61 (O_61,N_4986,N_4959);
xnor UO_62 (O_62,N_4971,N_4965);
nand UO_63 (O_63,N_4960,N_4955);
or UO_64 (O_64,N_4962,N_4911);
nand UO_65 (O_65,N_4938,N_4925);
or UO_66 (O_66,N_4979,N_4917);
and UO_67 (O_67,N_4961,N_4932);
nor UO_68 (O_68,N_4929,N_4940);
and UO_69 (O_69,N_4912,N_4948);
or UO_70 (O_70,N_4968,N_4900);
or UO_71 (O_71,N_4972,N_4986);
and UO_72 (O_72,N_4919,N_4901);
nand UO_73 (O_73,N_4933,N_4961);
nor UO_74 (O_74,N_4952,N_4932);
xnor UO_75 (O_75,N_4999,N_4945);
nand UO_76 (O_76,N_4913,N_4910);
nor UO_77 (O_77,N_4910,N_4988);
nand UO_78 (O_78,N_4957,N_4925);
and UO_79 (O_79,N_4915,N_4932);
nand UO_80 (O_80,N_4910,N_4938);
or UO_81 (O_81,N_4992,N_4906);
nand UO_82 (O_82,N_4942,N_4916);
nand UO_83 (O_83,N_4931,N_4980);
or UO_84 (O_84,N_4936,N_4983);
and UO_85 (O_85,N_4908,N_4955);
or UO_86 (O_86,N_4952,N_4925);
and UO_87 (O_87,N_4926,N_4937);
nor UO_88 (O_88,N_4981,N_4910);
xnor UO_89 (O_89,N_4969,N_4903);
and UO_90 (O_90,N_4994,N_4927);
or UO_91 (O_91,N_4941,N_4952);
and UO_92 (O_92,N_4968,N_4989);
or UO_93 (O_93,N_4982,N_4938);
nor UO_94 (O_94,N_4986,N_4924);
or UO_95 (O_95,N_4924,N_4932);
nor UO_96 (O_96,N_4909,N_4971);
and UO_97 (O_97,N_4970,N_4953);
or UO_98 (O_98,N_4981,N_4968);
and UO_99 (O_99,N_4974,N_4940);
xnor UO_100 (O_100,N_4964,N_4915);
and UO_101 (O_101,N_4986,N_4956);
and UO_102 (O_102,N_4986,N_4971);
or UO_103 (O_103,N_4994,N_4967);
nor UO_104 (O_104,N_4928,N_4963);
or UO_105 (O_105,N_4946,N_4952);
and UO_106 (O_106,N_4986,N_4908);
nor UO_107 (O_107,N_4960,N_4925);
nand UO_108 (O_108,N_4932,N_4945);
or UO_109 (O_109,N_4992,N_4954);
nor UO_110 (O_110,N_4951,N_4976);
nor UO_111 (O_111,N_4905,N_4908);
nor UO_112 (O_112,N_4908,N_4971);
nand UO_113 (O_113,N_4924,N_4984);
nor UO_114 (O_114,N_4956,N_4987);
or UO_115 (O_115,N_4976,N_4956);
nor UO_116 (O_116,N_4991,N_4912);
or UO_117 (O_117,N_4929,N_4941);
or UO_118 (O_118,N_4925,N_4920);
nand UO_119 (O_119,N_4921,N_4934);
xnor UO_120 (O_120,N_4948,N_4914);
or UO_121 (O_121,N_4923,N_4918);
nand UO_122 (O_122,N_4961,N_4997);
nand UO_123 (O_123,N_4955,N_4947);
and UO_124 (O_124,N_4924,N_4917);
and UO_125 (O_125,N_4957,N_4999);
or UO_126 (O_126,N_4987,N_4993);
nand UO_127 (O_127,N_4918,N_4982);
nand UO_128 (O_128,N_4916,N_4937);
and UO_129 (O_129,N_4964,N_4953);
or UO_130 (O_130,N_4950,N_4954);
nor UO_131 (O_131,N_4906,N_4964);
nor UO_132 (O_132,N_4914,N_4916);
nor UO_133 (O_133,N_4923,N_4982);
and UO_134 (O_134,N_4976,N_4907);
nand UO_135 (O_135,N_4958,N_4937);
nand UO_136 (O_136,N_4901,N_4959);
or UO_137 (O_137,N_4930,N_4974);
and UO_138 (O_138,N_4954,N_4967);
nor UO_139 (O_139,N_4997,N_4932);
or UO_140 (O_140,N_4994,N_4931);
nor UO_141 (O_141,N_4905,N_4961);
or UO_142 (O_142,N_4967,N_4970);
nor UO_143 (O_143,N_4983,N_4972);
nor UO_144 (O_144,N_4990,N_4936);
and UO_145 (O_145,N_4962,N_4978);
nor UO_146 (O_146,N_4967,N_4932);
or UO_147 (O_147,N_4907,N_4975);
and UO_148 (O_148,N_4961,N_4988);
or UO_149 (O_149,N_4995,N_4923);
nand UO_150 (O_150,N_4958,N_4946);
or UO_151 (O_151,N_4947,N_4985);
and UO_152 (O_152,N_4967,N_4983);
nor UO_153 (O_153,N_4968,N_4950);
nor UO_154 (O_154,N_4999,N_4991);
or UO_155 (O_155,N_4908,N_4929);
nor UO_156 (O_156,N_4904,N_4919);
and UO_157 (O_157,N_4997,N_4986);
nor UO_158 (O_158,N_4923,N_4962);
nand UO_159 (O_159,N_4971,N_4976);
xnor UO_160 (O_160,N_4960,N_4910);
or UO_161 (O_161,N_4920,N_4906);
nand UO_162 (O_162,N_4916,N_4966);
nand UO_163 (O_163,N_4900,N_4950);
nor UO_164 (O_164,N_4960,N_4952);
or UO_165 (O_165,N_4921,N_4981);
or UO_166 (O_166,N_4904,N_4941);
nor UO_167 (O_167,N_4923,N_4926);
and UO_168 (O_168,N_4965,N_4927);
nand UO_169 (O_169,N_4973,N_4971);
and UO_170 (O_170,N_4934,N_4969);
nand UO_171 (O_171,N_4998,N_4968);
and UO_172 (O_172,N_4923,N_4904);
nor UO_173 (O_173,N_4971,N_4907);
or UO_174 (O_174,N_4918,N_4973);
nand UO_175 (O_175,N_4903,N_4970);
or UO_176 (O_176,N_4925,N_4998);
nor UO_177 (O_177,N_4900,N_4909);
and UO_178 (O_178,N_4973,N_4998);
nand UO_179 (O_179,N_4909,N_4960);
or UO_180 (O_180,N_4977,N_4903);
or UO_181 (O_181,N_4920,N_4971);
or UO_182 (O_182,N_4948,N_4993);
or UO_183 (O_183,N_4937,N_4934);
nand UO_184 (O_184,N_4925,N_4918);
nand UO_185 (O_185,N_4965,N_4997);
nand UO_186 (O_186,N_4993,N_4922);
and UO_187 (O_187,N_4980,N_4933);
nand UO_188 (O_188,N_4999,N_4932);
nand UO_189 (O_189,N_4990,N_4976);
nor UO_190 (O_190,N_4943,N_4977);
or UO_191 (O_191,N_4949,N_4934);
or UO_192 (O_192,N_4918,N_4942);
nand UO_193 (O_193,N_4946,N_4959);
or UO_194 (O_194,N_4980,N_4928);
nand UO_195 (O_195,N_4938,N_4994);
and UO_196 (O_196,N_4986,N_4999);
and UO_197 (O_197,N_4990,N_4937);
and UO_198 (O_198,N_4998,N_4945);
nor UO_199 (O_199,N_4944,N_4976);
and UO_200 (O_200,N_4925,N_4989);
and UO_201 (O_201,N_4974,N_4969);
or UO_202 (O_202,N_4950,N_4926);
nand UO_203 (O_203,N_4912,N_4958);
and UO_204 (O_204,N_4916,N_4971);
nand UO_205 (O_205,N_4909,N_4951);
and UO_206 (O_206,N_4988,N_4931);
nand UO_207 (O_207,N_4978,N_4917);
and UO_208 (O_208,N_4960,N_4951);
or UO_209 (O_209,N_4952,N_4959);
or UO_210 (O_210,N_4974,N_4924);
xnor UO_211 (O_211,N_4955,N_4981);
or UO_212 (O_212,N_4901,N_4974);
or UO_213 (O_213,N_4926,N_4922);
nand UO_214 (O_214,N_4992,N_4994);
and UO_215 (O_215,N_4992,N_4956);
nand UO_216 (O_216,N_4907,N_4915);
or UO_217 (O_217,N_4971,N_4930);
and UO_218 (O_218,N_4976,N_4913);
and UO_219 (O_219,N_4988,N_4900);
or UO_220 (O_220,N_4985,N_4967);
or UO_221 (O_221,N_4902,N_4963);
nand UO_222 (O_222,N_4988,N_4956);
or UO_223 (O_223,N_4991,N_4981);
and UO_224 (O_224,N_4990,N_4948);
and UO_225 (O_225,N_4913,N_4940);
or UO_226 (O_226,N_4937,N_4905);
and UO_227 (O_227,N_4984,N_4932);
and UO_228 (O_228,N_4927,N_4987);
nand UO_229 (O_229,N_4906,N_4933);
or UO_230 (O_230,N_4993,N_4905);
nand UO_231 (O_231,N_4931,N_4996);
and UO_232 (O_232,N_4908,N_4927);
nor UO_233 (O_233,N_4907,N_4906);
nor UO_234 (O_234,N_4925,N_4980);
or UO_235 (O_235,N_4990,N_4932);
nand UO_236 (O_236,N_4991,N_4934);
or UO_237 (O_237,N_4993,N_4970);
or UO_238 (O_238,N_4920,N_4960);
nand UO_239 (O_239,N_4919,N_4989);
and UO_240 (O_240,N_4980,N_4915);
nand UO_241 (O_241,N_4918,N_4940);
and UO_242 (O_242,N_4974,N_4961);
or UO_243 (O_243,N_4909,N_4916);
xnor UO_244 (O_244,N_4925,N_4955);
nor UO_245 (O_245,N_4904,N_4915);
nor UO_246 (O_246,N_4907,N_4928);
nor UO_247 (O_247,N_4948,N_4974);
nand UO_248 (O_248,N_4922,N_4985);
and UO_249 (O_249,N_4969,N_4986);
nor UO_250 (O_250,N_4992,N_4977);
or UO_251 (O_251,N_4921,N_4945);
and UO_252 (O_252,N_4962,N_4958);
nand UO_253 (O_253,N_4983,N_4918);
nand UO_254 (O_254,N_4921,N_4974);
or UO_255 (O_255,N_4963,N_4908);
nor UO_256 (O_256,N_4973,N_4919);
nor UO_257 (O_257,N_4926,N_4928);
and UO_258 (O_258,N_4937,N_4918);
nand UO_259 (O_259,N_4910,N_4953);
and UO_260 (O_260,N_4949,N_4989);
or UO_261 (O_261,N_4964,N_4934);
nor UO_262 (O_262,N_4902,N_4946);
nand UO_263 (O_263,N_4984,N_4942);
or UO_264 (O_264,N_4957,N_4900);
or UO_265 (O_265,N_4946,N_4950);
or UO_266 (O_266,N_4950,N_4944);
or UO_267 (O_267,N_4908,N_4918);
and UO_268 (O_268,N_4984,N_4944);
nand UO_269 (O_269,N_4957,N_4965);
or UO_270 (O_270,N_4956,N_4983);
or UO_271 (O_271,N_4940,N_4926);
nor UO_272 (O_272,N_4953,N_4904);
nor UO_273 (O_273,N_4932,N_4939);
nor UO_274 (O_274,N_4930,N_4960);
nor UO_275 (O_275,N_4952,N_4957);
and UO_276 (O_276,N_4924,N_4903);
or UO_277 (O_277,N_4980,N_4929);
nand UO_278 (O_278,N_4988,N_4990);
nand UO_279 (O_279,N_4943,N_4911);
or UO_280 (O_280,N_4912,N_4920);
or UO_281 (O_281,N_4981,N_4943);
or UO_282 (O_282,N_4949,N_4988);
or UO_283 (O_283,N_4934,N_4936);
nand UO_284 (O_284,N_4993,N_4902);
and UO_285 (O_285,N_4948,N_4966);
or UO_286 (O_286,N_4909,N_4999);
or UO_287 (O_287,N_4914,N_4912);
or UO_288 (O_288,N_4906,N_4919);
or UO_289 (O_289,N_4922,N_4967);
nor UO_290 (O_290,N_4943,N_4935);
or UO_291 (O_291,N_4904,N_4964);
or UO_292 (O_292,N_4965,N_4995);
or UO_293 (O_293,N_4964,N_4996);
nand UO_294 (O_294,N_4908,N_4924);
and UO_295 (O_295,N_4996,N_4902);
nand UO_296 (O_296,N_4935,N_4992);
or UO_297 (O_297,N_4978,N_4915);
or UO_298 (O_298,N_4982,N_4964);
nor UO_299 (O_299,N_4930,N_4927);
or UO_300 (O_300,N_4945,N_4973);
or UO_301 (O_301,N_4935,N_4914);
nand UO_302 (O_302,N_4916,N_4920);
nand UO_303 (O_303,N_4912,N_4909);
nor UO_304 (O_304,N_4948,N_4978);
or UO_305 (O_305,N_4987,N_4913);
nor UO_306 (O_306,N_4978,N_4907);
and UO_307 (O_307,N_4937,N_4906);
or UO_308 (O_308,N_4967,N_4957);
and UO_309 (O_309,N_4981,N_4986);
nand UO_310 (O_310,N_4957,N_4915);
nand UO_311 (O_311,N_4984,N_4922);
nor UO_312 (O_312,N_4976,N_4986);
nor UO_313 (O_313,N_4936,N_4903);
and UO_314 (O_314,N_4913,N_4943);
nor UO_315 (O_315,N_4946,N_4999);
and UO_316 (O_316,N_4982,N_4972);
nand UO_317 (O_317,N_4998,N_4947);
nor UO_318 (O_318,N_4978,N_4927);
or UO_319 (O_319,N_4924,N_4934);
nand UO_320 (O_320,N_4958,N_4947);
and UO_321 (O_321,N_4991,N_4947);
nor UO_322 (O_322,N_4962,N_4976);
nor UO_323 (O_323,N_4927,N_4929);
nand UO_324 (O_324,N_4927,N_4997);
nor UO_325 (O_325,N_4981,N_4918);
nor UO_326 (O_326,N_4980,N_4943);
or UO_327 (O_327,N_4932,N_4902);
nand UO_328 (O_328,N_4960,N_4990);
or UO_329 (O_329,N_4913,N_4992);
and UO_330 (O_330,N_4963,N_4972);
nor UO_331 (O_331,N_4958,N_4981);
nand UO_332 (O_332,N_4963,N_4933);
nand UO_333 (O_333,N_4993,N_4960);
or UO_334 (O_334,N_4985,N_4982);
and UO_335 (O_335,N_4949,N_4943);
and UO_336 (O_336,N_4990,N_4962);
nand UO_337 (O_337,N_4982,N_4925);
or UO_338 (O_338,N_4912,N_4921);
nand UO_339 (O_339,N_4962,N_4939);
nor UO_340 (O_340,N_4918,N_4997);
nor UO_341 (O_341,N_4924,N_4939);
nand UO_342 (O_342,N_4954,N_4990);
or UO_343 (O_343,N_4905,N_4973);
and UO_344 (O_344,N_4997,N_4920);
or UO_345 (O_345,N_4953,N_4927);
nand UO_346 (O_346,N_4930,N_4998);
nor UO_347 (O_347,N_4930,N_4961);
nand UO_348 (O_348,N_4909,N_4936);
nand UO_349 (O_349,N_4904,N_4963);
nand UO_350 (O_350,N_4938,N_4903);
or UO_351 (O_351,N_4931,N_4973);
and UO_352 (O_352,N_4944,N_4959);
nand UO_353 (O_353,N_4968,N_4949);
nor UO_354 (O_354,N_4906,N_4934);
and UO_355 (O_355,N_4947,N_4990);
nor UO_356 (O_356,N_4960,N_4966);
and UO_357 (O_357,N_4932,N_4987);
and UO_358 (O_358,N_4972,N_4975);
or UO_359 (O_359,N_4971,N_4922);
or UO_360 (O_360,N_4924,N_4931);
and UO_361 (O_361,N_4917,N_4905);
and UO_362 (O_362,N_4972,N_4947);
and UO_363 (O_363,N_4968,N_4919);
nor UO_364 (O_364,N_4952,N_4908);
nand UO_365 (O_365,N_4900,N_4967);
or UO_366 (O_366,N_4917,N_4980);
xor UO_367 (O_367,N_4992,N_4937);
nor UO_368 (O_368,N_4941,N_4932);
nor UO_369 (O_369,N_4925,N_4996);
or UO_370 (O_370,N_4934,N_4987);
nand UO_371 (O_371,N_4952,N_4976);
nand UO_372 (O_372,N_4950,N_4979);
and UO_373 (O_373,N_4960,N_4988);
nor UO_374 (O_374,N_4934,N_4997);
nor UO_375 (O_375,N_4953,N_4986);
or UO_376 (O_376,N_4934,N_4988);
nor UO_377 (O_377,N_4988,N_4968);
nand UO_378 (O_378,N_4970,N_4992);
nor UO_379 (O_379,N_4980,N_4979);
or UO_380 (O_380,N_4954,N_4921);
nand UO_381 (O_381,N_4931,N_4962);
nor UO_382 (O_382,N_4943,N_4919);
or UO_383 (O_383,N_4942,N_4931);
or UO_384 (O_384,N_4968,N_4941);
or UO_385 (O_385,N_4904,N_4922);
nor UO_386 (O_386,N_4986,N_4968);
nand UO_387 (O_387,N_4953,N_4994);
nand UO_388 (O_388,N_4970,N_4968);
and UO_389 (O_389,N_4936,N_4952);
and UO_390 (O_390,N_4963,N_4968);
and UO_391 (O_391,N_4975,N_4923);
or UO_392 (O_392,N_4929,N_4974);
and UO_393 (O_393,N_4913,N_4930);
or UO_394 (O_394,N_4957,N_4968);
nand UO_395 (O_395,N_4901,N_4942);
and UO_396 (O_396,N_4969,N_4904);
nor UO_397 (O_397,N_4982,N_4975);
or UO_398 (O_398,N_4948,N_4986);
nor UO_399 (O_399,N_4957,N_4949);
nand UO_400 (O_400,N_4969,N_4988);
or UO_401 (O_401,N_4933,N_4990);
or UO_402 (O_402,N_4921,N_4957);
or UO_403 (O_403,N_4904,N_4974);
nand UO_404 (O_404,N_4970,N_4971);
and UO_405 (O_405,N_4925,N_4968);
and UO_406 (O_406,N_4958,N_4931);
nor UO_407 (O_407,N_4981,N_4900);
nor UO_408 (O_408,N_4950,N_4929);
or UO_409 (O_409,N_4931,N_4952);
and UO_410 (O_410,N_4952,N_4973);
nor UO_411 (O_411,N_4996,N_4952);
or UO_412 (O_412,N_4909,N_4945);
nor UO_413 (O_413,N_4983,N_4958);
nor UO_414 (O_414,N_4971,N_4993);
or UO_415 (O_415,N_4920,N_4963);
and UO_416 (O_416,N_4980,N_4978);
nor UO_417 (O_417,N_4945,N_4919);
nand UO_418 (O_418,N_4902,N_4903);
nand UO_419 (O_419,N_4969,N_4962);
and UO_420 (O_420,N_4935,N_4991);
nand UO_421 (O_421,N_4979,N_4922);
xnor UO_422 (O_422,N_4974,N_4954);
nor UO_423 (O_423,N_4955,N_4986);
nor UO_424 (O_424,N_4991,N_4975);
and UO_425 (O_425,N_4988,N_4924);
and UO_426 (O_426,N_4955,N_4995);
or UO_427 (O_427,N_4912,N_4956);
and UO_428 (O_428,N_4917,N_4973);
and UO_429 (O_429,N_4918,N_4948);
nor UO_430 (O_430,N_4956,N_4950);
or UO_431 (O_431,N_4922,N_4994);
or UO_432 (O_432,N_4928,N_4904);
and UO_433 (O_433,N_4997,N_4941);
or UO_434 (O_434,N_4949,N_4927);
or UO_435 (O_435,N_4952,N_4972);
nand UO_436 (O_436,N_4962,N_4932);
nand UO_437 (O_437,N_4985,N_4974);
nand UO_438 (O_438,N_4974,N_4946);
and UO_439 (O_439,N_4927,N_4984);
and UO_440 (O_440,N_4998,N_4926);
nand UO_441 (O_441,N_4997,N_4944);
nor UO_442 (O_442,N_4967,N_4901);
nand UO_443 (O_443,N_4926,N_4933);
xor UO_444 (O_444,N_4996,N_4968);
or UO_445 (O_445,N_4933,N_4909);
or UO_446 (O_446,N_4932,N_4982);
and UO_447 (O_447,N_4909,N_4914);
or UO_448 (O_448,N_4971,N_4992);
nand UO_449 (O_449,N_4965,N_4937);
nand UO_450 (O_450,N_4964,N_4954);
or UO_451 (O_451,N_4914,N_4913);
nor UO_452 (O_452,N_4992,N_4941);
or UO_453 (O_453,N_4915,N_4909);
and UO_454 (O_454,N_4972,N_4913);
or UO_455 (O_455,N_4945,N_4978);
and UO_456 (O_456,N_4950,N_4990);
and UO_457 (O_457,N_4904,N_4905);
nor UO_458 (O_458,N_4974,N_4922);
and UO_459 (O_459,N_4903,N_4916);
and UO_460 (O_460,N_4929,N_4934);
nand UO_461 (O_461,N_4904,N_4926);
nor UO_462 (O_462,N_4913,N_4964);
nand UO_463 (O_463,N_4913,N_4951);
or UO_464 (O_464,N_4932,N_4960);
nor UO_465 (O_465,N_4950,N_4914);
and UO_466 (O_466,N_4925,N_4958);
or UO_467 (O_467,N_4903,N_4959);
nand UO_468 (O_468,N_4985,N_4910);
and UO_469 (O_469,N_4941,N_4955);
nand UO_470 (O_470,N_4964,N_4942);
or UO_471 (O_471,N_4996,N_4961);
nand UO_472 (O_472,N_4982,N_4928);
and UO_473 (O_473,N_4949,N_4901);
nor UO_474 (O_474,N_4902,N_4960);
nor UO_475 (O_475,N_4983,N_4902);
xnor UO_476 (O_476,N_4995,N_4924);
nand UO_477 (O_477,N_4974,N_4931);
or UO_478 (O_478,N_4990,N_4996);
or UO_479 (O_479,N_4988,N_4954);
and UO_480 (O_480,N_4957,N_4923);
and UO_481 (O_481,N_4951,N_4987);
nor UO_482 (O_482,N_4949,N_4967);
nand UO_483 (O_483,N_4958,N_4949);
nor UO_484 (O_484,N_4919,N_4972);
nand UO_485 (O_485,N_4906,N_4979);
and UO_486 (O_486,N_4914,N_4953);
and UO_487 (O_487,N_4912,N_4917);
nor UO_488 (O_488,N_4960,N_4931);
or UO_489 (O_489,N_4991,N_4932);
and UO_490 (O_490,N_4930,N_4911);
or UO_491 (O_491,N_4930,N_4916);
or UO_492 (O_492,N_4930,N_4910);
nand UO_493 (O_493,N_4960,N_4908);
nor UO_494 (O_494,N_4969,N_4943);
or UO_495 (O_495,N_4975,N_4965);
or UO_496 (O_496,N_4987,N_4971);
or UO_497 (O_497,N_4910,N_4909);
or UO_498 (O_498,N_4923,N_4929);
nand UO_499 (O_499,N_4937,N_4911);
or UO_500 (O_500,N_4965,N_4932);
nor UO_501 (O_501,N_4994,N_4991);
nand UO_502 (O_502,N_4908,N_4900);
nor UO_503 (O_503,N_4953,N_4908);
nor UO_504 (O_504,N_4913,N_4998);
and UO_505 (O_505,N_4971,N_4925);
nand UO_506 (O_506,N_4937,N_4930);
or UO_507 (O_507,N_4986,N_4991);
or UO_508 (O_508,N_4902,N_4994);
nand UO_509 (O_509,N_4976,N_4981);
and UO_510 (O_510,N_4965,N_4956);
nor UO_511 (O_511,N_4903,N_4904);
nand UO_512 (O_512,N_4964,N_4952);
nor UO_513 (O_513,N_4919,N_4980);
nand UO_514 (O_514,N_4993,N_4947);
nand UO_515 (O_515,N_4944,N_4975);
nor UO_516 (O_516,N_4971,N_4994);
or UO_517 (O_517,N_4934,N_4960);
and UO_518 (O_518,N_4908,N_4992);
or UO_519 (O_519,N_4934,N_4925);
and UO_520 (O_520,N_4968,N_4954);
and UO_521 (O_521,N_4991,N_4937);
and UO_522 (O_522,N_4940,N_4946);
nor UO_523 (O_523,N_4911,N_4981);
xor UO_524 (O_524,N_4939,N_4955);
and UO_525 (O_525,N_4998,N_4972);
or UO_526 (O_526,N_4937,N_4954);
nand UO_527 (O_527,N_4919,N_4946);
nand UO_528 (O_528,N_4923,N_4954);
or UO_529 (O_529,N_4919,N_4912);
and UO_530 (O_530,N_4905,N_4922);
nor UO_531 (O_531,N_4940,N_4954);
and UO_532 (O_532,N_4988,N_4994);
nand UO_533 (O_533,N_4957,N_4908);
and UO_534 (O_534,N_4932,N_4933);
nor UO_535 (O_535,N_4902,N_4931);
nand UO_536 (O_536,N_4925,N_4963);
nand UO_537 (O_537,N_4940,N_4998);
nand UO_538 (O_538,N_4996,N_4991);
nor UO_539 (O_539,N_4993,N_4976);
and UO_540 (O_540,N_4913,N_4922);
nand UO_541 (O_541,N_4938,N_4996);
or UO_542 (O_542,N_4996,N_4997);
and UO_543 (O_543,N_4973,N_4970);
or UO_544 (O_544,N_4947,N_4968);
nand UO_545 (O_545,N_4916,N_4981);
or UO_546 (O_546,N_4955,N_4918);
or UO_547 (O_547,N_4986,N_4944);
or UO_548 (O_548,N_4932,N_4950);
nand UO_549 (O_549,N_4973,N_4920);
and UO_550 (O_550,N_4927,N_4922);
nor UO_551 (O_551,N_4941,N_4975);
nand UO_552 (O_552,N_4908,N_4968);
nand UO_553 (O_553,N_4989,N_4922);
nor UO_554 (O_554,N_4946,N_4920);
nand UO_555 (O_555,N_4958,N_4999);
nand UO_556 (O_556,N_4989,N_4902);
nor UO_557 (O_557,N_4905,N_4929);
and UO_558 (O_558,N_4958,N_4972);
nand UO_559 (O_559,N_4960,N_4924);
nor UO_560 (O_560,N_4998,N_4931);
nand UO_561 (O_561,N_4942,N_4940);
nand UO_562 (O_562,N_4971,N_4969);
nand UO_563 (O_563,N_4964,N_4957);
or UO_564 (O_564,N_4954,N_4953);
nor UO_565 (O_565,N_4985,N_4905);
and UO_566 (O_566,N_4961,N_4916);
nor UO_567 (O_567,N_4937,N_4910);
and UO_568 (O_568,N_4925,N_4944);
nand UO_569 (O_569,N_4978,N_4931);
nand UO_570 (O_570,N_4958,N_4990);
and UO_571 (O_571,N_4974,N_4902);
or UO_572 (O_572,N_4931,N_4970);
or UO_573 (O_573,N_4973,N_4962);
or UO_574 (O_574,N_4913,N_4945);
nand UO_575 (O_575,N_4932,N_4944);
or UO_576 (O_576,N_4904,N_4967);
and UO_577 (O_577,N_4994,N_4960);
nand UO_578 (O_578,N_4922,N_4940);
nand UO_579 (O_579,N_4923,N_4946);
nand UO_580 (O_580,N_4900,N_4951);
nor UO_581 (O_581,N_4977,N_4913);
and UO_582 (O_582,N_4916,N_4946);
and UO_583 (O_583,N_4919,N_4967);
nand UO_584 (O_584,N_4976,N_4996);
and UO_585 (O_585,N_4998,N_4904);
or UO_586 (O_586,N_4915,N_4925);
and UO_587 (O_587,N_4905,N_4933);
and UO_588 (O_588,N_4944,N_4987);
nor UO_589 (O_589,N_4936,N_4925);
nand UO_590 (O_590,N_4916,N_4968);
nor UO_591 (O_591,N_4905,N_4964);
nor UO_592 (O_592,N_4944,N_4923);
nor UO_593 (O_593,N_4958,N_4950);
nand UO_594 (O_594,N_4992,N_4979);
nor UO_595 (O_595,N_4967,N_4999);
nor UO_596 (O_596,N_4945,N_4972);
nand UO_597 (O_597,N_4957,N_4947);
nor UO_598 (O_598,N_4999,N_4903);
xor UO_599 (O_599,N_4901,N_4945);
nand UO_600 (O_600,N_4972,N_4918);
and UO_601 (O_601,N_4941,N_4915);
and UO_602 (O_602,N_4986,N_4947);
and UO_603 (O_603,N_4990,N_4931);
nand UO_604 (O_604,N_4906,N_4922);
and UO_605 (O_605,N_4942,N_4960);
nor UO_606 (O_606,N_4969,N_4991);
nor UO_607 (O_607,N_4941,N_4935);
or UO_608 (O_608,N_4985,N_4965);
nand UO_609 (O_609,N_4923,N_4986);
nand UO_610 (O_610,N_4960,N_4974);
nor UO_611 (O_611,N_4955,N_4957);
nor UO_612 (O_612,N_4929,N_4957);
or UO_613 (O_613,N_4997,N_4978);
nor UO_614 (O_614,N_4977,N_4905);
and UO_615 (O_615,N_4966,N_4965);
or UO_616 (O_616,N_4907,N_4991);
nor UO_617 (O_617,N_4901,N_4944);
nand UO_618 (O_618,N_4997,N_4900);
or UO_619 (O_619,N_4932,N_4900);
and UO_620 (O_620,N_4946,N_4996);
or UO_621 (O_621,N_4946,N_4900);
nor UO_622 (O_622,N_4908,N_4907);
nor UO_623 (O_623,N_4924,N_4954);
or UO_624 (O_624,N_4992,N_4958);
xnor UO_625 (O_625,N_4936,N_4949);
or UO_626 (O_626,N_4961,N_4993);
and UO_627 (O_627,N_4932,N_4935);
or UO_628 (O_628,N_4909,N_4937);
nor UO_629 (O_629,N_4949,N_4933);
or UO_630 (O_630,N_4993,N_4933);
nor UO_631 (O_631,N_4943,N_4903);
nor UO_632 (O_632,N_4914,N_4900);
or UO_633 (O_633,N_4916,N_4982);
or UO_634 (O_634,N_4965,N_4944);
and UO_635 (O_635,N_4902,N_4962);
or UO_636 (O_636,N_4900,N_4992);
or UO_637 (O_637,N_4985,N_4997);
nand UO_638 (O_638,N_4951,N_4992);
and UO_639 (O_639,N_4951,N_4945);
or UO_640 (O_640,N_4983,N_4949);
xor UO_641 (O_641,N_4997,N_4975);
and UO_642 (O_642,N_4947,N_4915);
and UO_643 (O_643,N_4933,N_4958);
or UO_644 (O_644,N_4964,N_4903);
nand UO_645 (O_645,N_4963,N_4903);
and UO_646 (O_646,N_4964,N_4971);
and UO_647 (O_647,N_4953,N_4968);
or UO_648 (O_648,N_4940,N_4902);
or UO_649 (O_649,N_4925,N_4973);
and UO_650 (O_650,N_4975,N_4903);
and UO_651 (O_651,N_4945,N_4917);
or UO_652 (O_652,N_4973,N_4991);
and UO_653 (O_653,N_4912,N_4908);
nor UO_654 (O_654,N_4952,N_4929);
nor UO_655 (O_655,N_4975,N_4904);
and UO_656 (O_656,N_4972,N_4910);
or UO_657 (O_657,N_4924,N_4973);
nor UO_658 (O_658,N_4938,N_4945);
nand UO_659 (O_659,N_4978,N_4908);
or UO_660 (O_660,N_4978,N_4966);
nor UO_661 (O_661,N_4952,N_4913);
nand UO_662 (O_662,N_4945,N_4950);
nor UO_663 (O_663,N_4990,N_4927);
nor UO_664 (O_664,N_4945,N_4971);
and UO_665 (O_665,N_4905,N_4921);
nand UO_666 (O_666,N_4958,N_4945);
and UO_667 (O_667,N_4985,N_4913);
or UO_668 (O_668,N_4914,N_4925);
nor UO_669 (O_669,N_4909,N_4955);
nor UO_670 (O_670,N_4940,N_4947);
and UO_671 (O_671,N_4975,N_4936);
nor UO_672 (O_672,N_4915,N_4905);
nor UO_673 (O_673,N_4923,N_4941);
and UO_674 (O_674,N_4901,N_4972);
nand UO_675 (O_675,N_4932,N_4925);
nor UO_676 (O_676,N_4950,N_4915);
nand UO_677 (O_677,N_4966,N_4969);
nand UO_678 (O_678,N_4953,N_4929);
xnor UO_679 (O_679,N_4914,N_4941);
nor UO_680 (O_680,N_4929,N_4994);
nor UO_681 (O_681,N_4922,N_4957);
nor UO_682 (O_682,N_4988,N_4911);
or UO_683 (O_683,N_4913,N_4954);
and UO_684 (O_684,N_4906,N_4932);
or UO_685 (O_685,N_4993,N_4932);
nor UO_686 (O_686,N_4984,N_4983);
or UO_687 (O_687,N_4957,N_4934);
nor UO_688 (O_688,N_4996,N_4943);
or UO_689 (O_689,N_4913,N_4905);
nand UO_690 (O_690,N_4928,N_4975);
nand UO_691 (O_691,N_4946,N_4991);
and UO_692 (O_692,N_4963,N_4953);
nor UO_693 (O_693,N_4964,N_4976);
nor UO_694 (O_694,N_4970,N_4991);
or UO_695 (O_695,N_4960,N_4992);
nor UO_696 (O_696,N_4979,N_4907);
and UO_697 (O_697,N_4959,N_4989);
and UO_698 (O_698,N_4965,N_4951);
nor UO_699 (O_699,N_4956,N_4915);
or UO_700 (O_700,N_4957,N_4920);
nand UO_701 (O_701,N_4916,N_4906);
or UO_702 (O_702,N_4998,N_4919);
and UO_703 (O_703,N_4951,N_4928);
and UO_704 (O_704,N_4996,N_4922);
or UO_705 (O_705,N_4935,N_4977);
nor UO_706 (O_706,N_4981,N_4925);
or UO_707 (O_707,N_4980,N_4911);
or UO_708 (O_708,N_4905,N_4927);
nor UO_709 (O_709,N_4943,N_4967);
nor UO_710 (O_710,N_4978,N_4979);
nor UO_711 (O_711,N_4921,N_4969);
and UO_712 (O_712,N_4955,N_4940);
nor UO_713 (O_713,N_4911,N_4965);
or UO_714 (O_714,N_4991,N_4909);
xnor UO_715 (O_715,N_4933,N_4997);
or UO_716 (O_716,N_4916,N_4949);
nor UO_717 (O_717,N_4936,N_4948);
xnor UO_718 (O_718,N_4991,N_4917);
or UO_719 (O_719,N_4991,N_4901);
nand UO_720 (O_720,N_4927,N_4901);
and UO_721 (O_721,N_4951,N_4944);
or UO_722 (O_722,N_4964,N_4922);
and UO_723 (O_723,N_4967,N_4923);
nor UO_724 (O_724,N_4963,N_4966);
nand UO_725 (O_725,N_4950,N_4904);
and UO_726 (O_726,N_4986,N_4915);
nand UO_727 (O_727,N_4908,N_4991);
nand UO_728 (O_728,N_4945,N_4947);
nand UO_729 (O_729,N_4940,N_4906);
nor UO_730 (O_730,N_4927,N_4950);
nand UO_731 (O_731,N_4975,N_4994);
nor UO_732 (O_732,N_4900,N_4977);
nand UO_733 (O_733,N_4980,N_4975);
nand UO_734 (O_734,N_4950,N_4910);
nand UO_735 (O_735,N_4970,N_4930);
or UO_736 (O_736,N_4989,N_4908);
nor UO_737 (O_737,N_4972,N_4900);
nand UO_738 (O_738,N_4976,N_4940);
nor UO_739 (O_739,N_4973,N_4900);
or UO_740 (O_740,N_4950,N_4919);
and UO_741 (O_741,N_4954,N_4947);
nor UO_742 (O_742,N_4911,N_4936);
and UO_743 (O_743,N_4956,N_4946);
or UO_744 (O_744,N_4978,N_4900);
and UO_745 (O_745,N_4992,N_4919);
nand UO_746 (O_746,N_4988,N_4904);
nor UO_747 (O_747,N_4990,N_4900);
or UO_748 (O_748,N_4988,N_4915);
or UO_749 (O_749,N_4904,N_4997);
nand UO_750 (O_750,N_4929,N_4991);
and UO_751 (O_751,N_4920,N_4952);
nor UO_752 (O_752,N_4904,N_4912);
nor UO_753 (O_753,N_4929,N_4996);
nor UO_754 (O_754,N_4984,N_4968);
nor UO_755 (O_755,N_4908,N_4993);
nor UO_756 (O_756,N_4968,N_4937);
or UO_757 (O_757,N_4918,N_4954);
nor UO_758 (O_758,N_4927,N_4944);
xnor UO_759 (O_759,N_4982,N_4980);
or UO_760 (O_760,N_4996,N_4959);
nor UO_761 (O_761,N_4971,N_4936);
nand UO_762 (O_762,N_4921,N_4917);
nand UO_763 (O_763,N_4944,N_4908);
nor UO_764 (O_764,N_4960,N_4945);
nand UO_765 (O_765,N_4907,N_4902);
or UO_766 (O_766,N_4900,N_4937);
or UO_767 (O_767,N_4976,N_4912);
nor UO_768 (O_768,N_4997,N_4913);
and UO_769 (O_769,N_4981,N_4941);
nand UO_770 (O_770,N_4971,N_4984);
xor UO_771 (O_771,N_4931,N_4959);
and UO_772 (O_772,N_4955,N_4984);
and UO_773 (O_773,N_4930,N_4925);
nor UO_774 (O_774,N_4933,N_4902);
nor UO_775 (O_775,N_4915,N_4971);
nand UO_776 (O_776,N_4952,N_4977);
nor UO_777 (O_777,N_4933,N_4945);
nand UO_778 (O_778,N_4994,N_4958);
or UO_779 (O_779,N_4955,N_4994);
nand UO_780 (O_780,N_4927,N_4989);
and UO_781 (O_781,N_4916,N_4990);
nor UO_782 (O_782,N_4911,N_4902);
nand UO_783 (O_783,N_4984,N_4960);
and UO_784 (O_784,N_4965,N_4933);
and UO_785 (O_785,N_4974,N_4993);
nor UO_786 (O_786,N_4973,N_4953);
nor UO_787 (O_787,N_4978,N_4984);
and UO_788 (O_788,N_4988,N_4997);
nor UO_789 (O_789,N_4956,N_4963);
and UO_790 (O_790,N_4901,N_4914);
xor UO_791 (O_791,N_4921,N_4922);
or UO_792 (O_792,N_4907,N_4984);
nand UO_793 (O_793,N_4925,N_4927);
nand UO_794 (O_794,N_4983,N_4944);
nand UO_795 (O_795,N_4974,N_4982);
and UO_796 (O_796,N_4995,N_4999);
nor UO_797 (O_797,N_4975,N_4946);
nor UO_798 (O_798,N_4902,N_4929);
nand UO_799 (O_799,N_4936,N_4961);
or UO_800 (O_800,N_4902,N_4979);
or UO_801 (O_801,N_4960,N_4999);
nor UO_802 (O_802,N_4955,N_4977);
nand UO_803 (O_803,N_4991,N_4983);
nand UO_804 (O_804,N_4937,N_4919);
and UO_805 (O_805,N_4937,N_4976);
or UO_806 (O_806,N_4945,N_4979);
or UO_807 (O_807,N_4941,N_4976);
nand UO_808 (O_808,N_4936,N_4995);
and UO_809 (O_809,N_4956,N_4999);
and UO_810 (O_810,N_4940,N_4981);
nand UO_811 (O_811,N_4999,N_4914);
or UO_812 (O_812,N_4926,N_4907);
and UO_813 (O_813,N_4979,N_4984);
or UO_814 (O_814,N_4988,N_4967);
nor UO_815 (O_815,N_4914,N_4989);
nand UO_816 (O_816,N_4901,N_4978);
nor UO_817 (O_817,N_4939,N_4980);
and UO_818 (O_818,N_4935,N_4939);
nand UO_819 (O_819,N_4920,N_4984);
and UO_820 (O_820,N_4962,N_4934);
nand UO_821 (O_821,N_4928,N_4971);
nand UO_822 (O_822,N_4982,N_4903);
or UO_823 (O_823,N_4940,N_4948);
nand UO_824 (O_824,N_4942,N_4909);
or UO_825 (O_825,N_4980,N_4949);
or UO_826 (O_826,N_4933,N_4951);
or UO_827 (O_827,N_4951,N_4982);
nand UO_828 (O_828,N_4953,N_4961);
and UO_829 (O_829,N_4910,N_4942);
nor UO_830 (O_830,N_4950,N_4969);
nor UO_831 (O_831,N_4935,N_4995);
nand UO_832 (O_832,N_4996,N_4975);
nand UO_833 (O_833,N_4959,N_4983);
nand UO_834 (O_834,N_4997,N_4919);
or UO_835 (O_835,N_4987,N_4978);
or UO_836 (O_836,N_4908,N_4985);
and UO_837 (O_837,N_4905,N_4984);
or UO_838 (O_838,N_4937,N_4964);
and UO_839 (O_839,N_4967,N_4910);
nand UO_840 (O_840,N_4985,N_4918);
nor UO_841 (O_841,N_4984,N_4981);
xnor UO_842 (O_842,N_4952,N_4975);
nor UO_843 (O_843,N_4960,N_4971);
and UO_844 (O_844,N_4945,N_4970);
or UO_845 (O_845,N_4967,N_4998);
and UO_846 (O_846,N_4941,N_4969);
nand UO_847 (O_847,N_4950,N_4935);
nor UO_848 (O_848,N_4993,N_4996);
nand UO_849 (O_849,N_4987,N_4911);
nand UO_850 (O_850,N_4948,N_4968);
or UO_851 (O_851,N_4971,N_4927);
and UO_852 (O_852,N_4904,N_4962);
nand UO_853 (O_853,N_4964,N_4958);
or UO_854 (O_854,N_4953,N_4939);
nand UO_855 (O_855,N_4910,N_4934);
nor UO_856 (O_856,N_4963,N_4916);
and UO_857 (O_857,N_4930,N_4923);
or UO_858 (O_858,N_4950,N_4984);
and UO_859 (O_859,N_4910,N_4926);
nand UO_860 (O_860,N_4987,N_4954);
nand UO_861 (O_861,N_4922,N_4981);
and UO_862 (O_862,N_4956,N_4949);
or UO_863 (O_863,N_4960,N_4962);
nor UO_864 (O_864,N_4949,N_4921);
and UO_865 (O_865,N_4935,N_4989);
and UO_866 (O_866,N_4957,N_4911);
and UO_867 (O_867,N_4962,N_4957);
and UO_868 (O_868,N_4921,N_4939);
or UO_869 (O_869,N_4946,N_4981);
nor UO_870 (O_870,N_4927,N_4904);
and UO_871 (O_871,N_4957,N_4979);
or UO_872 (O_872,N_4924,N_4993);
nand UO_873 (O_873,N_4971,N_4948);
or UO_874 (O_874,N_4973,N_4908);
or UO_875 (O_875,N_4911,N_4916);
nor UO_876 (O_876,N_4995,N_4931);
and UO_877 (O_877,N_4925,N_4941);
or UO_878 (O_878,N_4952,N_4933);
nand UO_879 (O_879,N_4975,N_4926);
and UO_880 (O_880,N_4970,N_4908);
and UO_881 (O_881,N_4947,N_4914);
nor UO_882 (O_882,N_4900,N_4952);
nand UO_883 (O_883,N_4948,N_4916);
nor UO_884 (O_884,N_4967,N_4980);
and UO_885 (O_885,N_4902,N_4914);
or UO_886 (O_886,N_4945,N_4985);
xor UO_887 (O_887,N_4966,N_4912);
or UO_888 (O_888,N_4937,N_4972);
and UO_889 (O_889,N_4915,N_4933);
or UO_890 (O_890,N_4910,N_4947);
and UO_891 (O_891,N_4998,N_4974);
nand UO_892 (O_892,N_4976,N_4972);
or UO_893 (O_893,N_4905,N_4912);
or UO_894 (O_894,N_4926,N_4935);
nand UO_895 (O_895,N_4962,N_4994);
and UO_896 (O_896,N_4933,N_4959);
or UO_897 (O_897,N_4960,N_4980);
nand UO_898 (O_898,N_4915,N_4968);
nor UO_899 (O_899,N_4950,N_4987);
and UO_900 (O_900,N_4900,N_4904);
or UO_901 (O_901,N_4913,N_4993);
and UO_902 (O_902,N_4999,N_4934);
or UO_903 (O_903,N_4963,N_4992);
nand UO_904 (O_904,N_4985,N_4995);
or UO_905 (O_905,N_4978,N_4955);
and UO_906 (O_906,N_4997,N_4969);
nor UO_907 (O_907,N_4998,N_4966);
nor UO_908 (O_908,N_4984,N_4969);
and UO_909 (O_909,N_4922,N_4918);
and UO_910 (O_910,N_4933,N_4919);
nand UO_911 (O_911,N_4979,N_4905);
or UO_912 (O_912,N_4975,N_4958);
and UO_913 (O_913,N_4988,N_4966);
or UO_914 (O_914,N_4916,N_4910);
nor UO_915 (O_915,N_4946,N_4925);
nor UO_916 (O_916,N_4931,N_4929);
and UO_917 (O_917,N_4920,N_4993);
nand UO_918 (O_918,N_4915,N_4924);
or UO_919 (O_919,N_4901,N_4957);
nor UO_920 (O_920,N_4951,N_4948);
nor UO_921 (O_921,N_4932,N_4958);
nor UO_922 (O_922,N_4924,N_4996);
nand UO_923 (O_923,N_4907,N_4913);
nor UO_924 (O_924,N_4950,N_4970);
and UO_925 (O_925,N_4923,N_4952);
or UO_926 (O_926,N_4917,N_4929);
or UO_927 (O_927,N_4947,N_4999);
and UO_928 (O_928,N_4962,N_4988);
nand UO_929 (O_929,N_4950,N_4913);
xor UO_930 (O_930,N_4944,N_4907);
and UO_931 (O_931,N_4961,N_4948);
nor UO_932 (O_932,N_4918,N_4938);
nor UO_933 (O_933,N_4996,N_4988);
or UO_934 (O_934,N_4934,N_4976);
and UO_935 (O_935,N_4946,N_4906);
and UO_936 (O_936,N_4977,N_4982);
and UO_937 (O_937,N_4905,N_4903);
and UO_938 (O_938,N_4955,N_4900);
nand UO_939 (O_939,N_4969,N_4963);
nor UO_940 (O_940,N_4920,N_4932);
and UO_941 (O_941,N_4934,N_4980);
nand UO_942 (O_942,N_4935,N_4951);
nor UO_943 (O_943,N_4953,N_4998);
nor UO_944 (O_944,N_4947,N_4932);
nand UO_945 (O_945,N_4984,N_4991);
nand UO_946 (O_946,N_4940,N_4941);
and UO_947 (O_947,N_4924,N_4978);
and UO_948 (O_948,N_4914,N_4920);
nor UO_949 (O_949,N_4977,N_4968);
and UO_950 (O_950,N_4980,N_4958);
and UO_951 (O_951,N_4991,N_4993);
nand UO_952 (O_952,N_4941,N_4948);
nor UO_953 (O_953,N_4905,N_4924);
nor UO_954 (O_954,N_4955,N_4983);
nor UO_955 (O_955,N_4922,N_4911);
or UO_956 (O_956,N_4970,N_4952);
nand UO_957 (O_957,N_4954,N_4916);
or UO_958 (O_958,N_4936,N_4920);
nand UO_959 (O_959,N_4967,N_4973);
nor UO_960 (O_960,N_4950,N_4930);
or UO_961 (O_961,N_4939,N_4971);
nor UO_962 (O_962,N_4946,N_4983);
nand UO_963 (O_963,N_4918,N_4931);
or UO_964 (O_964,N_4959,N_4947);
or UO_965 (O_965,N_4935,N_4921);
nand UO_966 (O_966,N_4922,N_4999);
and UO_967 (O_967,N_4931,N_4948);
xor UO_968 (O_968,N_4967,N_4931);
nor UO_969 (O_969,N_4933,N_4954);
nor UO_970 (O_970,N_4964,N_4920);
nor UO_971 (O_971,N_4971,N_4931);
nand UO_972 (O_972,N_4974,N_4933);
and UO_973 (O_973,N_4936,N_4951);
and UO_974 (O_974,N_4991,N_4911);
nor UO_975 (O_975,N_4974,N_4970);
and UO_976 (O_976,N_4948,N_4956);
or UO_977 (O_977,N_4911,N_4905);
xor UO_978 (O_978,N_4905,N_4925);
nor UO_979 (O_979,N_4955,N_4928);
nor UO_980 (O_980,N_4922,N_4928);
xor UO_981 (O_981,N_4983,N_4971);
nand UO_982 (O_982,N_4953,N_4924);
or UO_983 (O_983,N_4913,N_4939);
nor UO_984 (O_984,N_4911,N_4998);
nor UO_985 (O_985,N_4974,N_4949);
or UO_986 (O_986,N_4949,N_4932);
and UO_987 (O_987,N_4946,N_4964);
nand UO_988 (O_988,N_4950,N_4931);
or UO_989 (O_989,N_4966,N_4950);
and UO_990 (O_990,N_4980,N_4923);
or UO_991 (O_991,N_4962,N_4946);
xor UO_992 (O_992,N_4999,N_4983);
or UO_993 (O_993,N_4998,N_4933);
nor UO_994 (O_994,N_4908,N_4902);
or UO_995 (O_995,N_4976,N_4987);
xnor UO_996 (O_996,N_4964,N_4919);
nor UO_997 (O_997,N_4905,N_4936);
nor UO_998 (O_998,N_4927,N_4972);
nor UO_999 (O_999,N_4977,N_4995);
endmodule