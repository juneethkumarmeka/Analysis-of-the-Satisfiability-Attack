module basic_2500_25000_3000_20_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
and U0 (N_0,In_1167,In_962);
nand U1 (N_1,In_825,In_657);
or U2 (N_2,In_484,In_1085);
nand U3 (N_3,In_997,In_1092);
nor U4 (N_4,In_2115,In_1969);
xnor U5 (N_5,In_1105,In_1359);
or U6 (N_6,In_2245,In_476);
xor U7 (N_7,In_1975,In_1494);
nand U8 (N_8,In_1889,In_1285);
nor U9 (N_9,In_134,In_805);
and U10 (N_10,In_1340,In_937);
or U11 (N_11,In_192,In_274);
xor U12 (N_12,In_1112,In_2278);
nor U13 (N_13,In_866,In_1010);
xnor U14 (N_14,In_640,In_773);
nor U15 (N_15,In_2369,In_517);
or U16 (N_16,In_1307,In_79);
nand U17 (N_17,In_2061,In_322);
nand U18 (N_18,In_1472,In_2094);
nand U19 (N_19,In_1398,In_1294);
xnor U20 (N_20,In_1028,In_1148);
nand U21 (N_21,In_2430,In_1577);
and U22 (N_22,In_463,In_404);
xor U23 (N_23,In_1566,In_1266);
nor U24 (N_24,In_1888,In_2335);
xor U25 (N_25,In_802,In_454);
xor U26 (N_26,In_102,In_1449);
and U27 (N_27,In_2065,In_2029);
xor U28 (N_28,In_2285,In_277);
nor U29 (N_29,In_1676,In_818);
nand U30 (N_30,In_2219,In_2379);
or U31 (N_31,In_191,In_612);
and U32 (N_32,In_392,In_219);
or U33 (N_33,In_2046,In_1200);
nand U34 (N_34,In_1293,In_1925);
xor U35 (N_35,In_1065,In_296);
xnor U36 (N_36,In_1048,In_2414);
xnor U37 (N_37,In_336,In_590);
nand U38 (N_38,In_1938,In_1988);
nor U39 (N_39,In_1662,In_1612);
nand U40 (N_40,In_493,In_508);
and U41 (N_41,In_433,In_1042);
nor U42 (N_42,In_1950,In_376);
or U43 (N_43,In_173,In_679);
xnor U44 (N_44,In_418,In_2121);
xnor U45 (N_45,In_967,In_2069);
or U46 (N_46,In_1180,In_1927);
nor U47 (N_47,In_2087,In_1502);
nor U48 (N_48,In_490,In_437);
nor U49 (N_49,In_1102,In_1273);
and U50 (N_50,In_1729,In_45);
or U51 (N_51,In_609,In_1191);
or U52 (N_52,In_1891,In_1773);
nand U53 (N_53,In_1739,In_1688);
nand U54 (N_54,In_1617,In_1344);
or U55 (N_55,In_1986,In_1335);
xor U56 (N_56,In_2328,In_2075);
xnor U57 (N_57,In_1257,In_1972);
nor U58 (N_58,In_2008,In_2176);
xnor U59 (N_59,In_248,In_2330);
or U60 (N_60,In_1334,In_1245);
and U61 (N_61,In_2064,In_42);
and U62 (N_62,In_390,In_668);
or U63 (N_63,In_152,In_2169);
nand U64 (N_64,In_1051,In_511);
nand U65 (N_65,In_177,In_592);
nor U66 (N_66,In_228,In_25);
xor U67 (N_67,In_214,In_1527);
or U68 (N_68,In_602,In_1208);
xnor U69 (N_69,In_681,In_330);
nand U70 (N_70,In_798,In_350);
and U71 (N_71,In_1815,In_1685);
and U72 (N_72,In_408,In_1901);
nand U73 (N_73,In_1223,In_243);
nand U74 (N_74,In_2036,In_557);
nand U75 (N_75,In_2256,In_1415);
nor U76 (N_76,In_844,In_477);
and U77 (N_77,In_1757,In_975);
or U78 (N_78,In_1535,In_647);
or U79 (N_79,In_287,In_67);
nor U80 (N_80,In_982,In_2054);
and U81 (N_81,In_648,In_231);
nand U82 (N_82,In_817,In_1263);
nand U83 (N_83,In_1680,In_1402);
nor U84 (N_84,In_1802,In_136);
nor U85 (N_85,In_986,In_1130);
nor U86 (N_86,In_1118,In_1342);
nor U87 (N_87,In_1162,In_1567);
and U88 (N_88,In_1633,In_553);
nand U89 (N_89,In_1880,In_2186);
and U90 (N_90,In_2324,In_2400);
or U91 (N_91,In_1934,In_1176);
nand U92 (N_92,In_512,In_2487);
or U93 (N_93,In_2048,In_1740);
or U94 (N_94,In_1545,In_1380);
xor U95 (N_95,In_298,In_1337);
nand U96 (N_96,In_1262,In_1411);
or U97 (N_97,In_1893,In_1900);
or U98 (N_98,In_1957,In_1390);
and U99 (N_99,In_789,In_1247);
or U100 (N_100,In_217,In_721);
nor U101 (N_101,In_1997,In_394);
and U102 (N_102,In_1844,In_1106);
xnor U103 (N_103,In_1687,In_2150);
nand U104 (N_104,In_930,In_444);
nand U105 (N_105,In_1447,In_1722);
and U106 (N_106,In_529,In_251);
and U107 (N_107,In_2000,In_2091);
and U108 (N_108,In_1603,In_854);
nand U109 (N_109,In_1470,In_2331);
or U110 (N_110,In_522,In_22);
nand U111 (N_111,In_1933,In_288);
nor U112 (N_112,In_429,In_329);
nand U113 (N_113,In_342,In_1939);
nor U114 (N_114,In_128,In_1872);
nand U115 (N_115,In_2337,In_951);
nand U116 (N_116,In_398,In_2103);
and U117 (N_117,In_201,In_2031);
and U118 (N_118,In_1296,In_486);
or U119 (N_119,In_331,In_283);
xnor U120 (N_120,In_513,In_725);
or U121 (N_121,In_1562,In_893);
xnor U122 (N_122,In_1735,In_1797);
and U123 (N_123,In_880,In_1446);
xnor U124 (N_124,In_1227,In_1963);
and U125 (N_125,In_1890,In_1543);
or U126 (N_126,In_138,In_510);
nor U127 (N_127,In_1994,In_2300);
nor U128 (N_128,In_1279,In_1357);
xnor U129 (N_129,In_1462,In_2154);
nand U130 (N_130,In_1752,In_302);
xnor U131 (N_131,In_850,In_2021);
and U132 (N_132,In_2153,In_103);
nand U133 (N_133,In_1322,In_1333);
or U134 (N_134,In_621,In_348);
and U135 (N_135,In_1749,In_940);
or U136 (N_136,In_1116,In_2211);
nor U137 (N_137,In_2173,In_865);
nor U138 (N_138,In_717,In_868);
and U139 (N_139,In_1374,In_1941);
nor U140 (N_140,In_713,In_2005);
nand U141 (N_141,In_1239,In_5);
and U142 (N_142,In_1049,In_110);
nand U143 (N_143,In_1730,In_2033);
and U144 (N_144,In_2267,In_2015);
and U145 (N_145,In_1177,In_1706);
or U146 (N_146,In_2417,In_1012);
xnor U147 (N_147,In_1626,In_1634);
nand U148 (N_148,In_838,In_2477);
xnor U149 (N_149,In_642,In_2009);
nand U150 (N_150,In_1817,In_1153);
or U151 (N_151,In_597,In_821);
xnor U152 (N_152,In_846,In_605);
xor U153 (N_153,In_1955,In_1666);
xor U154 (N_154,In_263,In_1859);
nand U155 (N_155,In_1766,In_1134);
nand U156 (N_156,In_87,In_1576);
xnor U157 (N_157,In_935,In_1769);
nor U158 (N_158,In_917,In_858);
xnor U159 (N_159,In_1828,In_2078);
nor U160 (N_160,In_816,In_895);
xor U161 (N_161,In_2360,In_2393);
nor U162 (N_162,In_699,In_1647);
and U163 (N_163,In_1811,In_1942);
nand U164 (N_164,In_595,In_1231);
and U165 (N_165,In_2212,In_677);
nor U166 (N_166,In_536,In_1723);
xor U167 (N_167,In_181,In_1038);
or U168 (N_168,In_255,In_2081);
nor U169 (N_169,In_1354,In_1305);
and U170 (N_170,In_2019,In_669);
nand U171 (N_171,In_2411,In_1765);
xnor U172 (N_172,In_1993,In_2207);
xnor U173 (N_173,In_1186,In_807);
nor U174 (N_174,In_730,In_1318);
nor U175 (N_175,In_2436,In_1675);
nand U176 (N_176,In_772,In_1520);
nor U177 (N_177,In_2425,In_2114);
and U178 (N_178,In_803,In_631);
xnor U179 (N_179,In_505,In_2308);
xor U180 (N_180,In_1921,In_548);
or U181 (N_181,In_460,In_1211);
xnor U182 (N_182,In_2066,In_1024);
nand U183 (N_183,In_443,In_1556);
xor U184 (N_184,In_2011,In_1001);
and U185 (N_185,In_445,In_2101);
nor U186 (N_186,In_1631,In_666);
xor U187 (N_187,In_1873,In_89);
xor U188 (N_188,In_1281,In_1373);
or U189 (N_189,In_545,In_1426);
xnor U190 (N_190,In_1850,In_913);
and U191 (N_191,In_912,In_1516);
or U192 (N_192,In_161,In_746);
and U193 (N_193,In_2344,In_11);
nor U194 (N_194,In_1827,In_886);
nor U195 (N_195,In_2292,In_422);
nor U196 (N_196,In_869,In_726);
and U197 (N_197,In_2349,In_1259);
and U198 (N_198,In_573,In_2467);
or U199 (N_199,In_2225,In_1151);
xnor U200 (N_200,In_981,In_171);
or U201 (N_201,In_1220,In_2437);
nand U202 (N_202,In_313,In_574);
nor U203 (N_203,In_1958,In_569);
xor U204 (N_204,In_964,In_2110);
nand U205 (N_205,In_963,In_897);
or U206 (N_206,In_1463,In_987);
nand U207 (N_207,In_2144,In_83);
and U208 (N_208,In_2161,In_1824);
nor U209 (N_209,In_1096,In_831);
nand U210 (N_210,In_1254,In_1272);
and U211 (N_211,In_1141,In_1442);
and U212 (N_212,In_1212,In_386);
nor U213 (N_213,In_2096,In_253);
xnor U214 (N_214,In_372,In_1338);
or U215 (N_215,In_1104,In_18);
nor U216 (N_216,In_1636,In_1756);
and U217 (N_217,In_1393,In_48);
or U218 (N_218,In_2276,In_76);
nand U219 (N_219,In_1816,In_2403);
and U220 (N_220,In_377,In_1388);
nand U221 (N_221,In_1260,In_949);
or U222 (N_222,In_1860,In_1173);
or U223 (N_223,In_1922,In_1488);
nor U224 (N_224,In_114,In_1629);
nand U225 (N_225,In_141,In_523);
nand U226 (N_226,In_97,In_1882);
nor U227 (N_227,In_1268,In_1965);
or U228 (N_228,In_1299,In_2018);
xor U229 (N_229,In_1836,In_1763);
or U230 (N_230,In_1871,In_169);
or U231 (N_231,In_1482,In_1786);
nand U232 (N_232,In_2220,In_1286);
xor U233 (N_233,In_1733,In_2465);
and U234 (N_234,In_2269,In_1109);
nand U235 (N_235,In_636,In_1269);
nor U236 (N_236,In_945,In_1495);
or U237 (N_237,In_1854,In_2104);
nand U238 (N_238,In_1724,In_380);
nor U239 (N_239,In_1005,In_1421);
or U240 (N_240,In_1264,In_604);
nor U241 (N_241,In_2304,In_2310);
or U242 (N_242,In_627,In_2298);
nand U243 (N_243,In_1652,In_914);
and U244 (N_244,In_1140,In_349);
and U245 (N_245,In_1003,In_93);
or U246 (N_246,In_402,In_994);
nand U247 (N_247,In_225,In_485);
nand U248 (N_248,In_1774,In_2357);
nand U249 (N_249,In_2387,In_310);
and U250 (N_250,In_1485,In_2301);
xor U251 (N_251,In_665,In_20);
nand U252 (N_252,In_2440,In_800);
and U253 (N_253,In_2463,In_2395);
nand U254 (N_254,In_2258,In_759);
nand U255 (N_255,In_2312,In_279);
and U256 (N_256,In_1098,In_29);
nor U257 (N_257,In_1758,In_521);
nor U258 (N_258,In_345,In_1677);
or U259 (N_259,In_2442,In_591);
and U260 (N_260,In_1613,In_1297);
nor U261 (N_261,In_1360,In_927);
nor U262 (N_262,In_203,In_983);
xor U263 (N_263,In_689,In_1404);
xnor U264 (N_264,In_1182,In_306);
nor U265 (N_265,In_1420,In_760);
or U266 (N_266,In_535,In_2406);
nand U267 (N_267,In_1233,In_1940);
nor U268 (N_268,In_776,In_1914);
nand U269 (N_269,In_1445,In_256);
and U270 (N_270,In_224,In_1280);
nor U271 (N_271,In_2082,In_43);
nand U272 (N_272,In_791,In_147);
and U273 (N_273,In_2012,In_2486);
xor U274 (N_274,In_881,In_1776);
nor U275 (N_275,In_1812,In_1936);
xnor U276 (N_276,In_1413,In_2025);
xnor U277 (N_277,In_1499,In_27);
nor U278 (N_278,In_2108,In_1466);
and U279 (N_279,In_1129,In_1163);
xnor U280 (N_280,In_2364,In_1632);
nand U281 (N_281,In_1863,In_252);
or U282 (N_282,In_526,In_2419);
or U283 (N_283,In_2255,In_2452);
and U284 (N_284,In_455,In_614);
xnor U285 (N_285,In_496,In_0);
nand U286 (N_286,In_1084,In_2228);
nor U287 (N_287,In_840,In_124);
xor U288 (N_288,In_2164,In_1255);
nor U289 (N_289,In_448,In_1935);
or U290 (N_290,In_2028,In_2356);
and U291 (N_291,In_635,In_696);
and U292 (N_292,In_2351,In_2183);
nand U293 (N_293,In_1584,In_921);
xor U294 (N_294,In_1309,In_2290);
and U295 (N_295,In_1371,In_2429);
or U296 (N_296,In_1581,In_49);
nor U297 (N_297,In_140,In_1206);
nand U298 (N_298,In_206,In_775);
and U299 (N_299,In_26,In_1833);
and U300 (N_300,In_544,In_2178);
or U301 (N_301,In_2171,In_797);
or U302 (N_302,In_1923,In_1968);
nor U303 (N_303,In_2151,In_780);
and U304 (N_304,In_1287,In_1616);
and U305 (N_305,In_339,In_2197);
and U306 (N_306,In_1989,In_946);
nand U307 (N_307,In_2149,In_2318);
xor U308 (N_308,In_2187,In_1928);
and U309 (N_309,In_497,In_1573);
nor U310 (N_310,In_1668,In_1987);
and U311 (N_311,In_616,In_450);
nand U312 (N_312,In_2405,In_1205);
or U313 (N_313,In_2490,In_1887);
nand U314 (N_314,In_1468,In_487);
or U315 (N_315,In_1131,In_728);
nand U316 (N_316,In_471,In_947);
or U317 (N_317,In_2205,In_1588);
and U318 (N_318,In_1667,In_1951);
nand U319 (N_319,In_673,In_1378);
or U320 (N_320,In_2136,In_1214);
or U321 (N_321,In_1423,In_989);
or U322 (N_322,In_1326,In_462);
xor U323 (N_323,In_1031,In_1156);
xnor U324 (N_324,In_1295,In_853);
or U325 (N_325,In_318,In_808);
and U326 (N_326,In_1501,In_388);
xor U327 (N_327,In_13,In_561);
nand U328 (N_328,In_290,In_1181);
nand U329 (N_329,In_1138,In_499);
and U330 (N_330,In_1553,In_1672);
and U331 (N_331,In_323,In_516);
xor U332 (N_332,In_2232,In_745);
nand U333 (N_333,In_570,In_1356);
and U334 (N_334,In_1114,In_1355);
nor U335 (N_335,In_195,In_1582);
nand U336 (N_336,In_1209,In_1029);
or U337 (N_337,In_515,In_1215);
nor U338 (N_338,In_1438,In_271);
xor U339 (N_339,In_506,In_1103);
nand U340 (N_340,In_953,In_1228);
or U341 (N_341,In_828,In_1315);
nor U342 (N_342,In_2063,In_1074);
nand U343 (N_343,In_2489,In_2476);
nor U344 (N_344,In_1731,In_729);
xnor U345 (N_345,In_509,In_1699);
nor U346 (N_346,In_2263,In_183);
xnor U347 (N_347,In_1018,In_1546);
and U348 (N_348,In_2257,In_382);
xnor U349 (N_349,In_643,In_149);
xor U350 (N_350,In_2127,In_1391);
nand U351 (N_351,In_1199,In_1319);
and U352 (N_352,In_1312,In_1119);
nand U353 (N_353,In_1243,In_324);
or U354 (N_354,In_1169,In_2239);
xor U355 (N_355,In_1658,In_240);
xor U356 (N_356,In_1583,In_559);
xnor U357 (N_357,In_142,In_1060);
or U358 (N_358,In_2479,In_2168);
and U359 (N_359,In_2472,In_2170);
nor U360 (N_360,In_78,In_1819);
xor U361 (N_361,In_885,In_552);
nor U362 (N_362,In_174,In_738);
nor U363 (N_363,In_424,In_2462);
or U364 (N_364,In_2010,In_1068);
or U365 (N_365,In_98,In_2359);
xnor U366 (N_366,In_1977,In_1165);
or U367 (N_367,In_1943,In_1023);
nand U368 (N_368,In_2448,In_2071);
nand U369 (N_369,In_267,In_107);
or U370 (N_370,In_2043,In_2459);
nor U371 (N_371,In_1409,In_985);
xnor U372 (N_372,In_756,In_2342);
or U373 (N_373,In_675,In_835);
xor U374 (N_374,In_539,In_1548);
nor U375 (N_375,In_1659,In_1784);
nor U376 (N_376,In_46,In_420);
xor U377 (N_377,In_346,In_1715);
nor U378 (N_378,In_2293,In_855);
nor U379 (N_379,In_1241,In_1352);
xor U380 (N_380,In_974,In_2446);
xnor U381 (N_381,In_626,In_2279);
nand U382 (N_382,In_1753,In_2370);
nor U383 (N_383,In_1006,In_1793);
and U384 (N_384,In_1078,In_1747);
and U385 (N_385,In_1099,In_481);
xnor U386 (N_386,In_576,In_1483);
xnor U387 (N_387,In_1275,In_734);
or U388 (N_388,In_75,In_1175);
and U389 (N_389,In_2248,In_1072);
xor U390 (N_390,In_1086,In_623);
xor U391 (N_391,In_1184,In_1477);
and U392 (N_392,In_2365,In_784);
xor U393 (N_393,In_1304,In_309);
nor U394 (N_394,In_1133,In_1419);
xor U395 (N_395,In_754,In_1585);
xnor U396 (N_396,In_2264,In_2402);
and U397 (N_397,In_1610,In_90);
and U398 (N_398,In_413,In_1121);
xnor U399 (N_399,In_1213,In_2280);
and U400 (N_400,In_761,In_2152);
nand U401 (N_401,In_2399,In_1792);
and U402 (N_402,In_1804,In_145);
and U403 (N_403,In_1909,In_888);
nor U404 (N_404,In_379,In_1606);
nand U405 (N_405,In_439,In_572);
and U406 (N_406,In_118,In_1755);
xor U407 (N_407,In_2034,In_286);
and U408 (N_408,In_1403,In_1320);
xnor U409 (N_409,In_1575,In_2496);
xnor U410 (N_410,In_2193,In_1796);
nor U411 (N_411,In_1471,In_64);
nand U412 (N_412,In_1517,In_827);
or U413 (N_413,In_1400,In_347);
and U414 (N_414,In_1240,In_1506);
nand U415 (N_415,In_1427,In_1826);
nor U416 (N_416,In_861,In_2195);
or U417 (N_417,In_524,In_1912);
nand U418 (N_418,In_2072,In_2247);
or U419 (N_419,In_2003,In_1999);
xnor U420 (N_420,In_712,In_1703);
and U421 (N_421,In_527,In_676);
nor U422 (N_422,In_495,In_193);
xnor U423 (N_423,In_1253,In_1478);
or U424 (N_424,In_2123,In_958);
nand U425 (N_425,In_1429,In_1679);
nor U426 (N_426,In_2179,In_826);
or U427 (N_427,In_580,In_362);
and U428 (N_428,In_541,In_1136);
nand U429 (N_429,In_1370,In_272);
nand U430 (N_430,In_1978,In_1539);
or U431 (N_431,In_239,In_2460);
and U432 (N_432,In_132,In_2286);
nor U433 (N_433,In_1041,In_334);
nor U434 (N_434,In_1061,In_1020);
nand U435 (N_435,In_2068,In_1578);
or U436 (N_436,In_633,In_859);
nand U437 (N_437,In_1823,In_2391);
or U438 (N_438,In_2233,In_2322);
nor U439 (N_439,In_979,In_1852);
xnor U440 (N_440,In_2394,In_211);
nor U441 (N_441,In_2478,In_582);
nor U442 (N_442,In_2013,In_1298);
nand U443 (N_443,In_66,In_1772);
and U444 (N_444,In_2456,In_624);
nor U445 (N_445,In_500,In_992);
and U446 (N_446,In_900,In_2373);
or U447 (N_447,In_2026,In_915);
xor U448 (N_448,In_2491,In_765);
or U449 (N_449,In_664,In_1079);
nand U450 (N_450,In_1845,In_1377);
nand U451 (N_451,In_998,In_2319);
xnor U452 (N_452,In_1709,In_1290);
or U453 (N_453,In_1011,In_2231);
or U454 (N_454,In_877,In_144);
nand U455 (N_455,In_2354,In_1700);
or U456 (N_456,In_355,In_189);
or U457 (N_457,In_758,In_94);
or U458 (N_458,In_2027,In_1097);
nand U459 (N_459,In_902,In_1368);
and U460 (N_460,In_2014,In_993);
xor U461 (N_461,In_2067,In_2044);
nand U462 (N_462,In_33,In_2332);
or U463 (N_463,In_889,In_1066);
and U464 (N_464,In_325,In_442);
and U465 (N_465,In_864,In_1242);
xor U466 (N_466,In_1707,In_158);
and U467 (N_467,In_1032,In_670);
and U468 (N_468,In_957,In_710);
nand U469 (N_469,In_718,In_2201);
or U470 (N_470,In_397,In_1408);
or U471 (N_471,In_179,In_432);
nor U472 (N_472,In_1638,In_787);
or U473 (N_473,In_366,In_2133);
or U474 (N_474,In_2481,In_1996);
nor U475 (N_475,In_1743,In_96);
or U476 (N_476,In_1788,In_1910);
or U477 (N_477,In_823,In_1952);
xor U478 (N_478,In_2397,In_2346);
xnor U479 (N_479,In_790,In_1046);
xnor U480 (N_480,In_1568,In_1196);
nand U481 (N_481,In_467,In_1056);
and U482 (N_482,In_1248,In_1705);
nor U483 (N_483,In_237,In_1649);
nand U484 (N_484,In_1554,In_2077);
or U485 (N_485,In_1453,In_1226);
and U486 (N_486,In_724,In_954);
and U487 (N_487,In_1837,In_2106);
nand U488 (N_488,In_554,In_116);
xnor U489 (N_489,In_6,In_2485);
nor U490 (N_490,In_538,In_2381);
nor U491 (N_491,In_839,In_1441);
xor U492 (N_492,In_1512,In_1475);
nand U493 (N_493,In_518,In_1440);
and U494 (N_494,In_2102,In_2494);
nand U495 (N_495,In_690,In_2158);
nand U496 (N_496,In_1748,In_973);
nand U497 (N_497,In_632,In_1655);
or U498 (N_498,In_2085,In_73);
nand U499 (N_499,In_753,In_2499);
xnor U500 (N_500,In_655,In_1916);
nor U501 (N_501,In_999,In_1076);
nand U502 (N_502,In_1644,In_1713);
and U503 (N_503,In_2283,In_601);
or U504 (N_504,In_369,In_371);
nand U505 (N_505,In_740,In_2140);
or U506 (N_506,In_1971,In_2238);
nand U507 (N_507,In_1684,In_587);
xor U508 (N_508,In_737,In_1761);
nand U509 (N_509,In_1580,In_1113);
xnor U510 (N_510,In_1235,In_1372);
nor U511 (N_511,In_378,In_232);
nand U512 (N_512,In_1050,In_768);
nor U513 (N_513,In_2086,In_1981);
or U514 (N_514,In_1591,In_438);
nand U515 (N_515,In_153,In_2118);
nor U516 (N_516,In_1452,In_414);
nor U517 (N_517,In_2469,In_340);
or U518 (N_518,In_2262,In_550);
and U519 (N_519,In_1124,In_1611);
nand U520 (N_520,In_2362,In_164);
nand U521 (N_521,In_1407,In_783);
and U522 (N_522,In_2252,In_2441);
and U523 (N_523,In_1976,In_971);
nand U524 (N_524,In_697,In_1203);
nor U525 (N_525,In_319,In_1164);
nand U526 (N_526,In_333,In_777);
or U527 (N_527,In_568,In_1974);
nor U528 (N_528,In_1270,In_901);
nor U529 (N_529,In_1528,In_2311);
nor U530 (N_530,In_1428,In_99);
nand U531 (N_531,In_1911,In_1267);
or U532 (N_532,In_2297,In_2431);
or U533 (N_533,In_464,In_1155);
or U534 (N_534,In_1665,In_1460);
nor U535 (N_535,In_1806,In_411);
xor U536 (N_536,In_199,In_395);
xnor U537 (N_537,In_1330,In_1696);
nand U538 (N_538,In_215,In_2229);
nor U539 (N_539,In_2303,In_1868);
xor U540 (N_540,In_1216,In_1853);
or U541 (N_541,In_786,In_1329);
nand U542 (N_542,In_899,In_8);
xor U543 (N_543,In_950,In_1188);
or U544 (N_544,In_2306,In_1597);
and U545 (N_545,In_1217,In_412);
nand U546 (N_546,In_2145,In_1857);
nor U547 (N_547,In_2353,In_1710);
nor U548 (N_548,In_2343,In_1201);
or U549 (N_549,In_1434,In_61);
nor U550 (N_550,In_2017,In_824);
or U551 (N_551,In_533,In_292);
xor U552 (N_552,In_498,In_2032);
and U553 (N_553,In_703,In_752);
or U554 (N_554,In_1656,In_1646);
nand U555 (N_555,In_1848,In_260);
nand U556 (N_556,In_1077,In_1834);
or U557 (N_557,In_714,In_663);
or U558 (N_558,In_3,In_1654);
nand U559 (N_559,In_238,In_1664);
and U560 (N_560,In_608,In_1465);
nand U561 (N_561,In_1641,In_617);
nor U562 (N_562,In_36,In_151);
nand U563 (N_563,In_1132,In_1682);
nor U564 (N_564,In_1094,In_704);
nand U565 (N_565,In_794,In_31);
nor U566 (N_566,In_1949,In_425);
nor U567 (N_567,In_91,In_1689);
or U568 (N_568,In_1946,In_700);
and U569 (N_569,In_1779,In_312);
and U570 (N_570,In_1410,In_135);
nand U571 (N_571,In_363,In_2157);
nor U572 (N_572,In_875,In_354);
xnor U573 (N_573,In_2454,In_53);
and U574 (N_574,In_1302,In_2202);
nand U575 (N_575,In_919,In_2422);
or U576 (N_576,In_600,In_299);
or U577 (N_577,In_1067,In_2272);
nor U578 (N_578,In_870,In_1498);
and U579 (N_579,In_1932,In_1607);
xnor U580 (N_580,In_190,In_2338);
or U581 (N_581,In_2056,In_2246);
nand U582 (N_582,In_1448,In_1300);
or U583 (N_583,In_1146,In_1628);
nand U584 (N_584,In_130,In_549);
or U585 (N_585,In_127,In_2438);
nor U586 (N_586,In_2492,In_261);
nand U587 (N_587,In_1288,In_692);
xnor U588 (N_588,In_1547,In_2389);
xor U589 (N_589,In_126,In_2461);
nor U590 (N_590,In_2165,In_1847);
or U591 (N_591,In_204,In_1904);
xor U592 (N_592,In_16,In_1081);
or U593 (N_593,In_848,In_646);
or U594 (N_594,In_1635,In_2270);
nor U595 (N_595,In_1657,In_1021);
nand U596 (N_596,In_2327,In_131);
nand U597 (N_597,In_1271,In_44);
and U598 (N_598,In_1202,In_1849);
and U599 (N_599,In_332,In_2385);
xor U600 (N_600,In_2007,In_56);
and U601 (N_601,In_1365,In_2471);
and U602 (N_602,In_1425,In_2458);
nor U603 (N_603,In_531,In_565);
nand U604 (N_604,In_1159,In_1336);
nand U605 (N_605,In_2146,In_1918);
nand U606 (N_606,In_1039,In_2497);
nor U607 (N_607,In_81,In_1725);
nor U608 (N_608,In_766,In_2420);
xnor U609 (N_609,In_980,In_811);
and U610 (N_610,In_2206,In_685);
or U611 (N_611,In_1992,In_28);
nor U612 (N_612,In_2234,In_2407);
nor U613 (N_613,In_80,In_1533);
xor U614 (N_614,In_571,In_2244);
xnor U615 (N_615,In_2392,In_291);
nor U616 (N_616,In_1306,In_1037);
nand U617 (N_617,In_1135,In_2413);
and U618 (N_618,In_1497,In_1358);
nand U619 (N_619,In_810,In_1444);
or U620 (N_620,In_1630,In_820);
nor U621 (N_621,In_555,In_1439);
and U622 (N_622,In_1224,In_1839);
or U623 (N_623,In_918,In_133);
or U624 (N_624,In_747,In_2271);
or U625 (N_625,In_1161,In_2177);
or U626 (N_626,In_165,In_1734);
nor U627 (N_627,In_1956,In_57);
and U628 (N_628,In_2375,In_1139);
and U629 (N_629,In_1947,In_1120);
xnor U630 (N_630,In_2049,In_482);
and U631 (N_631,In_814,In_262);
and U632 (N_632,In_1171,In_1572);
nor U633 (N_633,In_1571,In_733);
xnor U634 (N_634,In_2453,In_1317);
xor U635 (N_635,In_1750,In_2210);
nand U636 (N_636,In_2167,In_1781);
nand U637 (N_637,In_652,In_406);
nand U638 (N_638,In_942,In_583);
and U639 (N_639,In_1147,In_436);
and U640 (N_640,In_47,In_1621);
and U641 (N_641,In_273,In_1876);
nor U642 (N_642,In_441,In_593);
or U643 (N_643,In_658,In_1970);
nand U644 (N_644,In_1830,In_1714);
nor U645 (N_645,In_1973,In_1948);
and U646 (N_646,In_2289,In_154);
or U647 (N_647,In_212,In_567);
or U648 (N_648,In_1461,In_1708);
and U649 (N_649,In_1258,In_852);
xnor U650 (N_650,In_2449,In_1898);
xnor U651 (N_651,In_830,In_1350);
nor U652 (N_652,In_4,In_680);
or U653 (N_653,In_739,In_661);
xor U654 (N_654,In_2129,In_1033);
nand U655 (N_655,In_300,In_1515);
or U656 (N_656,In_847,In_2367);
nand U657 (N_657,In_72,In_2409);
nor U658 (N_658,In_1157,In_1126);
xor U659 (N_659,In_85,In_494);
or U660 (N_660,In_387,In_2339);
or U661 (N_661,In_749,In_30);
nand U662 (N_662,In_588,In_1745);
and U663 (N_663,In_1651,In_819);
nor U664 (N_664,In_916,In_584);
or U665 (N_665,In_1732,In_105);
and U666 (N_666,In_1767,In_2138);
or U667 (N_667,In_12,In_1013);
nor U668 (N_668,In_2198,In_1813);
xnor U669 (N_669,In_220,In_837);
nand U670 (N_670,In_483,In_2250);
xnor U671 (N_671,In_2268,In_1154);
and U672 (N_672,In_2281,In_295);
and U673 (N_673,In_2122,In_2057);
and U674 (N_674,In_1283,In_108);
nand U675 (N_675,In_182,In_1917);
xnor U676 (N_676,In_480,In_1587);
xor U677 (N_677,In_822,In_1906);
xnor U678 (N_678,In_1540,In_2288);
xor U679 (N_679,In_2296,In_1505);
and U680 (N_680,In_2004,In_1924);
xor U681 (N_681,In_528,In_1491);
xnor U682 (N_682,In_1091,In_2390);
nand U683 (N_683,In_1100,In_1985);
nor U684 (N_684,In_929,In_1406);
xor U685 (N_685,In_735,In_1351);
nor U686 (N_686,In_2191,In_1111);
nand U687 (N_687,In_1907,In_702);
and U688 (N_688,In_389,In_546);
xor U689 (N_689,In_51,In_688);
and U690 (N_690,In_1381,In_2041);
xor U691 (N_691,In_70,In_1504);
xnor U692 (N_692,In_1375,In_1292);
and U693 (N_693,In_2240,In_218);
or U694 (N_694,In_71,In_1596);
or U695 (N_695,In_1101,In_1387);
or U696 (N_696,In_1799,In_2180);
nor U697 (N_697,In_1158,In_1814);
xnor U698 (N_698,In_2204,In_2060);
and U699 (N_699,In_1702,In_1087);
or U700 (N_700,In_265,In_1526);
nor U701 (N_701,In_208,In_955);
and U702 (N_702,In_1168,In_1608);
nand U703 (N_703,In_1323,In_654);
nor U704 (N_704,In_146,In_2445);
xor U705 (N_705,In_2251,In_1875);
nand U706 (N_706,In_1726,In_2483);
xnor U707 (N_707,In_769,In_1277);
nor U708 (N_708,In_1308,In_1467);
xor U709 (N_709,In_360,In_1489);
and U710 (N_710,In_1744,In_328);
or U711 (N_711,In_1598,In_1451);
nand U712 (N_712,In_1301,In_2433);
xor U713 (N_713,In_542,In_23);
and U714 (N_714,In_1251,In_234);
or U715 (N_715,In_101,In_1062);
or U716 (N_716,In_876,In_1313);
or U717 (N_717,In_1246,In_2474);
and U718 (N_718,In_1149,In_1238);
xor U719 (N_719,In_194,In_1059);
xor U720 (N_720,In_1794,In_1623);
xor U721 (N_721,In_1574,In_1443);
and U722 (N_722,In_1325,In_1007);
nand U723 (N_723,In_867,In_948);
and U724 (N_724,In_829,In_1265);
xnor U725 (N_725,In_566,In_629);
or U726 (N_726,In_2037,In_1660);
xor U727 (N_727,In_10,In_1341);
or U728 (N_728,In_1110,In_1291);
or U729 (N_729,In_1673,In_17);
or U730 (N_730,In_1361,In_249);
or U731 (N_731,In_368,In_2484);
and U732 (N_732,In_743,In_358);
or U733 (N_733,In_970,In_2361);
nor U734 (N_734,In_1829,In_1604);
or U735 (N_735,In_2113,In_2073);
nand U736 (N_736,In_1383,In_401);
and U737 (N_737,In_1095,In_1962);
xnor U738 (N_738,In_1386,In_672);
nand U739 (N_739,In_474,In_1117);
nor U740 (N_740,In_2287,In_229);
xor U741 (N_741,In_2218,In_579);
nand U742 (N_742,In_1069,In_375);
nor U743 (N_743,In_430,In_2098);
nor U744 (N_744,In_1864,In_2295);
nand U745 (N_745,In_137,In_1751);
nor U746 (N_746,In_1579,In_393);
and U747 (N_747,In_1521,In_1492);
nor U748 (N_748,In_956,In_671);
or U749 (N_749,In_62,In_1401);
xnor U750 (N_750,In_2428,In_1532);
xor U751 (N_751,In_452,In_1855);
nor U752 (N_752,In_2473,In_1884);
and U753 (N_753,In_143,In_2495);
and U754 (N_754,In_1982,In_695);
nor U755 (N_755,In_1160,In_155);
or U756 (N_756,In_1524,In_1174);
nor U757 (N_757,In_407,In_1818);
or U758 (N_758,In_431,In_180);
nand U759 (N_759,In_645,In_1920);
nand U760 (N_760,In_1937,In_1686);
nand U761 (N_761,In_197,In_501);
xor U762 (N_762,In_2030,In_2355);
xor U763 (N_763,In_1044,In_2137);
nand U764 (N_764,In_532,In_38);
nor U765 (N_765,In_578,In_245);
and U766 (N_766,In_1002,In_293);
or U767 (N_767,In_1599,In_911);
and U768 (N_768,In_1785,In_1841);
or U769 (N_769,In_1053,In_1822);
nand U770 (N_770,In_2230,In_1648);
and U771 (N_771,In_1289,In_2119);
nor U772 (N_772,In_938,In_1261);
nor U773 (N_773,In_1552,In_1192);
nand U774 (N_774,In_1047,In_788);
xor U775 (N_775,In_316,In_941);
and U776 (N_776,In_1719,In_281);
nand U777 (N_777,In_1697,In_1727);
or U778 (N_778,In_589,In_732);
xnor U779 (N_779,In_2336,In_175);
nand U780 (N_780,In_2421,In_1503);
nor U781 (N_781,In_491,In_2388);
xor U782 (N_782,In_32,In_399);
nand U783 (N_783,In_2498,In_157);
or U784 (N_784,In_320,In_2090);
xnor U785 (N_785,In_1026,In_2190);
nor U786 (N_786,In_2383,In_1954);
xnor U787 (N_787,In_2147,In_1027);
nor U788 (N_788,In_230,In_1570);
nand U789 (N_789,In_966,In_119);
and U790 (N_790,In_1040,In_1913);
nor U791 (N_791,In_2265,In_1800);
xnor U792 (N_792,In_851,In_1509);
xor U793 (N_793,In_1881,In_596);
xor U794 (N_794,In_650,In_2475);
nor U795 (N_795,In_34,In_1754);
and U796 (N_796,In_1883,In_284);
nor U797 (N_797,In_1627,In_326);
nand U798 (N_798,In_479,In_129);
nor U799 (N_799,In_1197,In_1366);
nor U800 (N_800,In_1590,In_236);
and U801 (N_801,In_2224,In_1518);
nor U802 (N_802,In_1225,In_1244);
nand U803 (N_803,In_1979,In_720);
xnor U804 (N_804,In_2384,In_356);
and U805 (N_805,In_1432,In_1557);
and U806 (N_806,In_1045,In_1866);
xnor U807 (N_807,In_1137,In_1362);
nand U808 (N_808,In_2059,In_473);
xnor U809 (N_809,In_610,In_2099);
xnor U810 (N_810,In_556,In_659);
and U811 (N_811,In_2047,In_841);
xor U812 (N_812,In_2334,In_2074);
or U813 (N_813,In_1430,In_1534);
xnor U814 (N_814,In_2016,In_2447);
and U815 (N_815,In_1959,In_2022);
nor U816 (N_816,In_453,In_1178);
or U817 (N_817,In_514,In_2092);
xor U818 (N_818,In_1960,In_742);
xnor U819 (N_819,In_684,In_415);
nand U820 (N_820,In_1624,In_2404);
xnor U821 (N_821,In_1219,In_184);
xnor U822 (N_822,In_1369,In_1693);
and U823 (N_823,In_613,In_1983);
or U824 (N_824,In_2038,In_2274);
nor U825 (N_825,In_1455,In_932);
xnor U826 (N_826,In_715,In_1967);
and U827 (N_827,In_2439,In_2345);
nand U828 (N_828,In_2325,In_122);
or U829 (N_829,In_2235,In_634);
nand U830 (N_830,In_907,In_1284);
xor U831 (N_831,In_1310,In_1125);
nand U832 (N_832,In_314,In_1510);
xnor U833 (N_833,In_2222,In_492);
xor U834 (N_834,In_812,In_125);
nand U835 (N_835,In_2209,In_1303);
xnor U836 (N_836,In_871,In_667);
xnor U837 (N_837,In_1321,In_470);
xor U838 (N_838,In_1569,In_1183);
xnor U839 (N_839,In_2199,In_2480);
and U840 (N_840,In_2307,In_1842);
nor U841 (N_841,In_1674,In_2208);
nor U842 (N_842,In_843,In_303);
xor U843 (N_843,In_435,In_308);
or U844 (N_844,In_410,In_285);
and U845 (N_845,In_475,In_988);
and U846 (N_846,In_1778,In_1550);
nand U847 (N_847,In_1807,In_123);
xnor U848 (N_848,In_707,In_1746);
xnor U849 (N_849,In_1276,In_2236);
and U850 (N_850,In_1064,In_2);
nor U851 (N_851,In_365,In_266);
and U852 (N_852,In_2214,In_931);
nand U853 (N_853,In_196,In_1484);
and U854 (N_854,In_1343,In_1456);
nand U855 (N_855,In_781,In_920);
nand U856 (N_856,In_1500,In_1090);
nand U857 (N_857,In_586,In_391);
or U858 (N_858,In_898,In_1523);
nand U859 (N_859,In_221,In_774);
or U860 (N_860,In_2084,In_1538);
nand U861 (N_861,In_504,In_1998);
and U862 (N_862,In_2001,In_2468);
and U863 (N_863,In_1650,In_1143);
xnor U864 (N_864,In_115,In_706);
or U865 (N_865,In_1052,In_1514);
nand U866 (N_866,In_2120,In_644);
or U867 (N_867,In_423,In_2377);
or U868 (N_868,In_1663,In_405);
nand U869 (N_869,In_383,In_925);
xor U870 (N_870,In_1549,In_1128);
nand U871 (N_871,In_2398,In_489);
xor U872 (N_872,In_205,In_936);
and U873 (N_873,In_1770,In_1622);
or U874 (N_874,In_1966,In_1704);
xor U875 (N_875,In_1782,In_560);
xnor U876 (N_876,In_187,In_166);
and U877 (N_877,In_202,In_2051);
and U878 (N_878,In_618,In_619);
and U879 (N_879,In_857,In_2450);
nor U880 (N_880,In_40,In_1737);
nand U881 (N_881,In_1145,In_2444);
xor U882 (N_882,In_1716,In_1594);
nand U883 (N_883,In_2079,In_1327);
or U884 (N_884,In_1022,In_694);
nand U885 (N_885,In_1809,In_2163);
xor U886 (N_886,In_163,In_2174);
and U887 (N_887,In_1152,In_534);
nor U888 (N_888,In_63,In_1783);
or U889 (N_889,In_2159,In_344);
nand U890 (N_890,In_186,In_693);
nand U891 (N_891,In_804,In_1414);
nor U892 (N_892,In_1437,In_834);
xor U893 (N_893,In_1670,In_748);
and U894 (N_894,In_2316,In_2020);
or U895 (N_895,In_2347,In_1496);
nor U896 (N_896,In_335,In_2401);
xor U897 (N_897,In_785,In_2260);
nand U898 (N_898,In_2097,In_1348);
nor U899 (N_899,In_370,In_2216);
and U900 (N_900,In_488,In_2155);
nor U901 (N_901,In_351,In_2006);
nand U902 (N_902,In_990,In_1363);
xor U903 (N_903,In_1412,In_562);
xor U904 (N_904,In_2058,In_1314);
and U905 (N_905,In_577,In_1195);
and U906 (N_906,In_311,In_530);
xor U907 (N_907,In_2243,In_611);
and U908 (N_908,In_1980,In_2432);
and U909 (N_909,In_1563,In_244);
xnor U910 (N_910,In_836,In_2415);
and U911 (N_911,In_1190,In_1278);
xor U912 (N_912,In_537,In_995);
and U913 (N_913,In_2217,In_2314);
and U914 (N_914,In_1185,In_74);
nand U915 (N_915,In_1108,In_69);
and U916 (N_916,In_1479,In_606);
nand U917 (N_917,In_943,In_939);
nand U918 (N_918,In_2434,In_1058);
and U919 (N_919,In_519,In_1895);
xnor U920 (N_920,In_68,In_1930);
and U921 (N_921,In_1431,In_168);
or U922 (N_922,In_1142,In_1625);
nor U923 (N_923,In_965,In_1832);
xnor U924 (N_924,In_628,In_1331);
xnor U925 (N_925,In_873,In_419);
xor U926 (N_926,In_417,In_1459);
nand U927 (N_927,In_361,In_1602);
xor U928 (N_928,In_1530,In_792);
nand U929 (N_929,In_905,In_19);
or U930 (N_930,In_1903,In_2125);
nor U931 (N_931,In_104,In_1944);
and U932 (N_932,In_1678,In_2052);
nor U933 (N_933,In_160,In_317);
nor U934 (N_934,In_1820,In_1671);
or U935 (N_935,In_2372,In_1620);
nor U936 (N_936,In_162,In_246);
nor U937 (N_937,In_1905,In_1529);
xnor U938 (N_938,In_1874,In_2143);
xnor U939 (N_939,In_1127,In_1464);
nor U940 (N_940,In_357,In_1742);
nand U941 (N_941,In_353,In_856);
nand U942 (N_942,In_1862,In_2302);
nor U943 (N_943,In_1869,In_416);
xnor U944 (N_944,In_2242,In_1892);
nand U945 (N_945,In_2408,In_1249);
nand U946 (N_946,In_2466,In_1179);
nor U947 (N_947,In_1218,In_615);
nand U948 (N_948,In_890,In_2317);
nand U949 (N_949,In_1964,In_2215);
xor U950 (N_950,In_117,In_223);
or U951 (N_951,In_1795,In_109);
xor U952 (N_952,In_959,In_233);
nor U953 (N_953,In_1718,In_1861);
nand U954 (N_954,In_1899,In_1669);
nor U955 (N_955,In_282,In_2277);
or U956 (N_956,In_1394,In_796);
or U957 (N_957,In_1055,In_2350);
nand U958 (N_958,In_594,In_1640);
xnor U959 (N_959,In_637,In_1843);
xor U960 (N_960,In_926,In_39);
or U961 (N_961,In_969,In_1712);
xor U962 (N_962,In_209,In_686);
xnor U963 (N_963,In_2112,In_2053);
nor U964 (N_964,In_1711,In_2380);
xor U965 (N_965,In_2294,In_1870);
xor U966 (N_966,In_1115,In_1399);
nand U967 (N_967,In_7,In_1172);
nor U968 (N_968,In_2132,In_1803);
and U969 (N_969,In_258,In_884);
nand U970 (N_970,In_2291,In_649);
nor U971 (N_971,In_440,In_226);
nand U972 (N_972,In_305,In_396);
and U973 (N_973,In_1274,In_1653);
or U974 (N_974,In_2203,In_1063);
nand U975 (N_975,In_58,In_2135);
or U976 (N_976,In_575,In_367);
xor U977 (N_977,In_167,In_1777);
xnor U978 (N_978,In_465,In_466);
nor U979 (N_979,In_674,In_1555);
or U980 (N_980,In_1436,In_2089);
and U981 (N_981,In_1609,In_148);
and U982 (N_982,In_2376,In_1416);
xnor U983 (N_983,In_1821,In_928);
or U984 (N_984,In_2130,In_2435);
or U985 (N_985,In_1511,In_2320);
or U986 (N_986,In_2416,In_923);
nand U987 (N_987,In_1878,In_1389);
xnor U988 (N_988,In_1222,In_849);
and U989 (N_989,In_1519,In_2366);
or U990 (N_990,In_1564,In_1690);
nand U991 (N_991,In_120,In_178);
and U992 (N_992,In_2266,In_1558);
or U993 (N_993,In_1486,In_35);
or U994 (N_994,In_52,In_1030);
or U995 (N_995,In_1728,In_2455);
and U996 (N_996,In_1695,In_247);
xor U997 (N_997,In_620,In_1537);
nor U998 (N_998,In_1897,In_2426);
nand U999 (N_999,In_543,In_540);
nand U1000 (N_1000,In_1990,In_2134);
nand U1001 (N_1001,In_1995,In_1741);
or U1002 (N_1002,In_1886,In_1639);
nor U1003 (N_1003,In_892,In_687);
xor U1004 (N_1004,In_1614,In_1595);
and U1005 (N_1005,In_2457,In_1392);
nor U1006 (N_1006,In_1454,In_276);
and U1007 (N_1007,In_2083,In_978);
or U1008 (N_1008,In_1825,In_2396);
or U1009 (N_1009,In_1984,In_1771);
or U1010 (N_1010,In_996,In_1122);
nor U1011 (N_1011,In_159,In_2427);
nor U1012 (N_1012,In_1229,In_1643);
xor U1013 (N_1013,In_1513,In_1234);
xnor U1014 (N_1014,In_2088,In_2382);
or U1015 (N_1015,In_2358,In_9);
nor U1016 (N_1016,In_458,In_933);
xnor U1017 (N_1017,In_1736,In_50);
and U1018 (N_1018,In_1250,In_1107);
nand U1019 (N_1019,In_1170,In_1379);
nor U1020 (N_1020,In_1931,In_656);
or U1021 (N_1021,In_2340,In_2378);
nand U1022 (N_1022,In_1282,In_2482);
and U1023 (N_1023,In_2148,In_2363);
xor U1024 (N_1024,In_1457,In_1542);
xnor U1025 (N_1025,In_1721,In_421);
and U1026 (N_1026,In_741,In_2035);
xor U1027 (N_1027,In_625,In_968);
xor U1028 (N_1028,In_832,In_213);
or U1029 (N_1029,In_2323,In_156);
nand U1030 (N_1030,In_1014,In_960);
and U1031 (N_1031,In_1490,In_1692);
nand U1032 (N_1032,In_972,In_86);
xor U1033 (N_1033,In_2200,In_1762);
and U1034 (N_1034,In_385,In_1384);
nand U1035 (N_1035,In_2128,In_558);
or U1036 (N_1036,In_2412,In_449);
xnor U1037 (N_1037,In_1808,In_1618);
and U1038 (N_1038,In_2055,In_1541);
or U1039 (N_1039,In_2175,In_2172);
nor U1040 (N_1040,In_2282,In_1458);
or U1041 (N_1041,In_1480,In_1561);
and U1042 (N_1042,In_210,In_1805);
nor U1043 (N_1043,In_1953,In_879);
nand U1044 (N_1044,In_1150,In_660);
or U1045 (N_1045,In_139,In_771);
nor U1046 (N_1046,In_1789,In_1780);
xnor U1047 (N_1047,In_198,In_1586);
nor U1048 (N_1048,In_2237,In_307);
xor U1049 (N_1049,In_1089,In_944);
nand U1050 (N_1050,In_37,In_1004);
nor U1051 (N_1051,In_84,In_250);
or U1052 (N_1052,In_21,In_563);
nor U1053 (N_1053,In_150,In_1544);
nand U1054 (N_1054,In_1661,In_2424);
or U1055 (N_1055,In_1424,In_908);
xnor U1056 (N_1056,In_1787,In_341);
xnor U1057 (N_1057,In_170,In_472);
nand U1058 (N_1058,In_1592,In_2194);
xnor U1059 (N_1059,In_268,In_2464);
and U1060 (N_1060,In_1720,In_1000);
and U1061 (N_1061,In_581,In_121);
and U1062 (N_1062,In_1417,In_2488);
and U1063 (N_1063,In_1810,In_1194);
nand U1064 (N_1064,In_1851,In_1189);
or U1065 (N_1065,In_2002,In_1450);
and U1066 (N_1066,In_1252,In_903);
and U1067 (N_1067,In_374,In_2249);
and U1068 (N_1068,In_1036,In_641);
xor U1069 (N_1069,In_1493,In_95);
and U1070 (N_1070,In_289,In_722);
nand U1071 (N_1071,In_779,In_241);
nor U1072 (N_1072,In_2253,In_1054);
nand U1073 (N_1073,In_2124,In_384);
xor U1074 (N_1074,In_427,In_1698);
nand U1075 (N_1075,In_185,In_1025);
nand U1076 (N_1076,In_2241,In_2076);
nor U1077 (N_1077,In_736,In_2418);
xor U1078 (N_1078,In_961,In_1637);
xnor U1079 (N_1079,In_984,In_507);
nand U1080 (N_1080,In_2107,In_2126);
xor U1081 (N_1081,In_1311,In_1798);
and U1082 (N_1082,In_709,In_1896);
nand U1083 (N_1083,In_2299,In_2141);
or U1084 (N_1084,In_842,In_106);
xnor U1085 (N_1085,In_1166,In_1198);
nand U1086 (N_1086,In_1043,In_1071);
xor U1087 (N_1087,In_2341,In_478);
xnor U1088 (N_1088,In_269,In_904);
or U1089 (N_1089,In_343,In_60);
nand U1090 (N_1090,In_2080,In_1082);
and U1091 (N_1091,In_1681,In_216);
or U1092 (N_1092,In_952,In_1057);
or U1093 (N_1093,In_2100,In_1316);
or U1094 (N_1094,In_2156,In_862);
and U1095 (N_1095,In_2045,In_653);
and U1096 (N_1096,In_564,In_359);
or U1097 (N_1097,In_41,In_751);
nand U1098 (N_1098,In_793,In_188);
xnor U1099 (N_1099,In_1902,In_2470);
xor U1100 (N_1100,In_2254,In_1070);
nor U1101 (N_1101,In_1418,In_711);
nand U1102 (N_1102,In_922,In_15);
nor U1103 (N_1103,In_259,In_82);
xor U1104 (N_1104,In_1345,In_801);
nand U1105 (N_1105,In_1193,In_200);
nor U1106 (N_1106,In_764,In_400);
and U1107 (N_1107,In_352,In_744);
or U1108 (N_1108,In_2093,In_906);
xor U1109 (N_1109,In_1256,In_731);
nor U1110 (N_1110,In_2309,In_1221);
nor U1111 (N_1111,In_1487,In_1885);
and U1112 (N_1112,In_1605,In_1367);
nand U1113 (N_1113,In_2184,In_698);
or U1114 (N_1114,In_1867,In_1422);
or U1115 (N_1115,In_2329,In_882);
or U1116 (N_1116,In_770,In_1790);
or U1117 (N_1117,In_1376,In_1531);
nor U1118 (N_1118,In_2443,In_1207);
and U1119 (N_1119,In_469,In_1144);
nand U1120 (N_1120,In_2227,In_172);
nand U1121 (N_1121,In_2023,In_1522);
nand U1122 (N_1122,In_878,In_2062);
nor U1123 (N_1123,In_1801,In_705);
and U1124 (N_1124,In_1019,In_778);
nor U1125 (N_1125,In_1775,In_1615);
nor U1126 (N_1126,In_599,In_1017);
nand U1127 (N_1127,In_428,In_1009);
or U1128 (N_1128,In_2352,In_991);
xnor U1129 (N_1129,In_1332,In_403);
xor U1130 (N_1130,In_1691,In_54);
xor U1131 (N_1131,In_2042,In_1397);
and U1132 (N_1132,In_2105,In_1476);
and U1133 (N_1133,In_1589,In_457);
nand U1134 (N_1134,In_1991,In_1768);
or U1135 (N_1135,In_662,In_1645);
xnor U1136 (N_1136,In_1349,In_2024);
nand U1137 (N_1137,In_691,In_2386);
xor U1138 (N_1138,In_207,In_1237);
nor U1139 (N_1139,In_639,In_1879);
and U1140 (N_1140,In_2259,In_845);
nor U1141 (N_1141,In_1565,In_782);
xnor U1142 (N_1142,In_315,In_321);
or U1143 (N_1143,In_92,In_2305);
and U1144 (N_1144,In_2131,In_2321);
nand U1145 (N_1145,In_910,In_24);
nor U1146 (N_1146,In_459,In_909);
nand U1147 (N_1147,In_264,In_327);
nor U1148 (N_1148,In_2182,In_1339);
nor U1149 (N_1149,In_833,In_2192);
nand U1150 (N_1150,In_2070,In_270);
or U1151 (N_1151,In_1123,In_887);
xor U1152 (N_1152,In_1395,In_1187);
or U1153 (N_1153,In_1877,In_1694);
and U1154 (N_1154,In_2226,In_304);
or U1155 (N_1155,In_294,In_1945);
nand U1156 (N_1156,In_2095,In_278);
and U1157 (N_1157,In_1908,In_2451);
nand U1158 (N_1158,In_1559,In_750);
nand U1159 (N_1159,In_2313,In_2116);
xnor U1160 (N_1160,In_2284,In_1232);
nor U1161 (N_1161,In_1915,In_1525);
nor U1162 (N_1162,In_520,In_1894);
xnor U1163 (N_1163,In_860,In_55);
xor U1164 (N_1164,In_1601,In_1008);
or U1165 (N_1165,In_1385,In_585);
nand U1166 (N_1166,In_1347,In_1396);
nor U1167 (N_1167,In_1034,In_2261);
nand U1168 (N_1168,In_1961,In_176);
nor U1169 (N_1169,In_2275,In_2166);
xor U1170 (N_1170,In_275,In_1717);
nor U1171 (N_1171,In_603,In_280);
or U1172 (N_1172,In_682,In_2326);
nand U1173 (N_1173,In_1600,In_1015);
nor U1174 (N_1174,In_2221,In_874);
xnor U1175 (N_1175,In_1328,In_607);
or U1176 (N_1176,In_1619,In_806);
nor U1177 (N_1177,In_65,In_502);
or U1178 (N_1178,In_2213,In_254);
and U1179 (N_1179,In_1856,In_891);
nand U1180 (N_1180,In_1593,In_1080);
nand U1181 (N_1181,In_1835,In_1364);
xor U1182 (N_1182,In_451,In_622);
and U1183 (N_1183,In_2189,In_2111);
and U1184 (N_1184,In_2040,In_434);
nor U1185 (N_1185,In_1831,In_883);
nand U1186 (N_1186,In_795,In_373);
nand U1187 (N_1187,In_2188,In_683);
nor U1188 (N_1188,In_77,In_723);
or U1189 (N_1189,In_767,In_716);
nand U1190 (N_1190,In_381,In_1738);
or U1191 (N_1191,In_1642,In_1701);
nor U1192 (N_1192,In_461,In_2142);
nand U1193 (N_1193,In_301,In_651);
xor U1194 (N_1194,In_1353,In_762);
xor U1195 (N_1195,In_409,In_88);
or U1196 (N_1196,In_1210,In_719);
and U1197 (N_1197,In_338,In_2185);
nand U1198 (N_1198,In_2223,In_934);
nand U1199 (N_1199,In_2181,In_1474);
and U1200 (N_1200,In_364,In_1858);
or U1201 (N_1201,In_1507,In_297);
nand U1202 (N_1202,In_1536,In_2039);
or U1203 (N_1203,In_456,In_1865);
or U1204 (N_1204,In_1230,In_227);
and U1205 (N_1205,In_2315,In_896);
xor U1206 (N_1206,In_872,In_242);
or U1207 (N_1207,In_1035,In_1560);
or U1208 (N_1208,In_446,In_1929);
nand U1209 (N_1209,In_14,In_1838);
or U1210 (N_1210,In_2493,In_547);
or U1211 (N_1211,In_1840,In_863);
xnor U1212 (N_1212,In_1324,In_257);
or U1213 (N_1213,In_1,In_1083);
or U1214 (N_1214,In_708,In_503);
nand U1215 (N_1215,In_1791,In_447);
and U1216 (N_1216,In_100,In_113);
xor U1217 (N_1217,In_1473,In_809);
or U1218 (N_1218,In_1846,In_1093);
and U1219 (N_1219,In_1764,In_630);
and U1220 (N_1220,In_1435,In_1551);
nand U1221 (N_1221,In_1469,In_222);
or U1222 (N_1222,In_701,In_799);
nand U1223 (N_1223,In_976,In_2050);
nand U1224 (N_1224,In_2368,In_1346);
xor U1225 (N_1225,In_678,In_1433);
nor U1226 (N_1226,In_551,In_2160);
xnor U1227 (N_1227,In_235,In_2109);
xnor U1228 (N_1228,In_2139,In_2410);
nor U1229 (N_1229,In_1760,In_924);
xor U1230 (N_1230,In_727,In_1073);
or U1231 (N_1231,In_2273,In_2117);
nand U1232 (N_1232,In_1016,In_1919);
xnor U1233 (N_1233,In_598,In_1405);
nor U1234 (N_1234,In_1926,In_337);
xor U1235 (N_1235,In_755,In_1236);
nand U1236 (N_1236,In_2374,In_1382);
or U1237 (N_1237,In_763,In_468);
nand U1238 (N_1238,In_977,In_2162);
or U1239 (N_1239,In_1759,In_111);
xor U1240 (N_1240,In_815,In_1204);
or U1241 (N_1241,In_1075,In_2371);
or U1242 (N_1242,In_1481,In_59);
or U1243 (N_1243,In_2348,In_1088);
nor U1244 (N_1244,In_525,In_757);
nand U1245 (N_1245,In_894,In_2423);
and U1246 (N_1246,In_813,In_638);
nand U1247 (N_1247,In_2333,In_112);
nand U1248 (N_1248,In_1508,In_1683);
or U1249 (N_1249,In_2196,In_426);
nand U1250 (N_1250,N_844,N_596);
and U1251 (N_1251,N_851,N_285);
nand U1252 (N_1252,N_979,N_337);
and U1253 (N_1253,N_45,N_738);
and U1254 (N_1254,N_144,N_1058);
nor U1255 (N_1255,N_730,N_968);
nor U1256 (N_1256,N_804,N_971);
nor U1257 (N_1257,N_1066,N_231);
and U1258 (N_1258,N_834,N_761);
and U1259 (N_1259,N_956,N_422);
nor U1260 (N_1260,N_1211,N_710);
and U1261 (N_1261,N_982,N_725);
nor U1262 (N_1262,N_600,N_94);
or U1263 (N_1263,N_9,N_443);
nor U1264 (N_1264,N_862,N_856);
nand U1265 (N_1265,N_469,N_809);
nand U1266 (N_1266,N_161,N_107);
xnor U1267 (N_1267,N_184,N_437);
and U1268 (N_1268,N_825,N_670);
or U1269 (N_1269,N_141,N_133);
and U1270 (N_1270,N_256,N_789);
nand U1271 (N_1271,N_120,N_272);
and U1272 (N_1272,N_666,N_1247);
nand U1273 (N_1273,N_1244,N_1231);
nor U1274 (N_1274,N_420,N_924);
nand U1275 (N_1275,N_233,N_440);
and U1276 (N_1276,N_375,N_876);
nor U1277 (N_1277,N_798,N_1176);
and U1278 (N_1278,N_215,N_214);
or U1279 (N_1279,N_707,N_52);
nand U1280 (N_1280,N_362,N_1097);
or U1281 (N_1281,N_152,N_753);
nor U1282 (N_1282,N_77,N_728);
and U1283 (N_1283,N_486,N_498);
nor U1284 (N_1284,N_413,N_99);
nor U1285 (N_1285,N_65,N_897);
nor U1286 (N_1286,N_354,N_183);
nor U1287 (N_1287,N_574,N_790);
or U1288 (N_1288,N_145,N_988);
nor U1289 (N_1289,N_867,N_903);
nor U1290 (N_1290,N_833,N_742);
nor U1291 (N_1291,N_985,N_506);
nor U1292 (N_1292,N_129,N_279);
nand U1293 (N_1293,N_431,N_868);
or U1294 (N_1294,N_368,N_1132);
xor U1295 (N_1295,N_509,N_986);
or U1296 (N_1296,N_296,N_394);
nand U1297 (N_1297,N_808,N_628);
xor U1298 (N_1298,N_745,N_276);
and U1299 (N_1299,N_308,N_114);
nor U1300 (N_1300,N_1119,N_896);
and U1301 (N_1301,N_1127,N_150);
or U1302 (N_1302,N_73,N_775);
or U1303 (N_1303,N_1174,N_474);
and U1304 (N_1304,N_686,N_992);
xor U1305 (N_1305,N_14,N_1234);
xor U1306 (N_1306,N_603,N_189);
or U1307 (N_1307,N_983,N_1002);
nand U1308 (N_1308,N_417,N_275);
xor U1309 (N_1309,N_583,N_1131);
nor U1310 (N_1310,N_581,N_1001);
nor U1311 (N_1311,N_698,N_1167);
xor U1312 (N_1312,N_1050,N_1102);
or U1313 (N_1313,N_1226,N_427);
nor U1314 (N_1314,N_945,N_799);
xnor U1315 (N_1315,N_301,N_955);
nor U1316 (N_1316,N_453,N_902);
or U1317 (N_1317,N_60,N_619);
nand U1318 (N_1318,N_485,N_489);
or U1319 (N_1319,N_1191,N_1116);
nor U1320 (N_1320,N_58,N_1246);
or U1321 (N_1321,N_1206,N_932);
and U1322 (N_1322,N_432,N_180);
or U1323 (N_1323,N_614,N_1183);
xnor U1324 (N_1324,N_282,N_126);
nand U1325 (N_1325,N_363,N_51);
or U1326 (N_1326,N_845,N_930);
and U1327 (N_1327,N_1089,N_1194);
nor U1328 (N_1328,N_885,N_714);
nor U1329 (N_1329,N_158,N_43);
xor U1330 (N_1330,N_1181,N_942);
nand U1331 (N_1331,N_605,N_861);
or U1332 (N_1332,N_401,N_931);
and U1333 (N_1333,N_267,N_732);
nor U1334 (N_1334,N_33,N_482);
nor U1335 (N_1335,N_447,N_195);
and U1336 (N_1336,N_578,N_801);
xor U1337 (N_1337,N_1180,N_733);
or U1338 (N_1338,N_936,N_1038);
nor U1339 (N_1339,N_226,N_492);
xnor U1340 (N_1340,N_83,N_879);
or U1341 (N_1341,N_390,N_335);
xnor U1342 (N_1342,N_944,N_984);
xor U1343 (N_1343,N_53,N_1138);
and U1344 (N_1344,N_253,N_981);
nor U1345 (N_1345,N_850,N_1228);
nor U1346 (N_1346,N_365,N_777);
nor U1347 (N_1347,N_963,N_330);
and U1348 (N_1348,N_539,N_220);
nor U1349 (N_1349,N_22,N_371);
xnor U1350 (N_1350,N_199,N_576);
nor U1351 (N_1351,N_779,N_1200);
nand U1352 (N_1352,N_84,N_379);
or U1353 (N_1353,N_917,N_1120);
and U1354 (N_1354,N_1039,N_56);
nand U1355 (N_1355,N_1125,N_1158);
nor U1356 (N_1356,N_892,N_46);
nand U1357 (N_1357,N_591,N_828);
xnor U1358 (N_1358,N_452,N_642);
xnor U1359 (N_1359,N_1151,N_617);
and U1360 (N_1360,N_722,N_1145);
nor U1361 (N_1361,N_697,N_211);
nand U1362 (N_1362,N_747,N_127);
nor U1363 (N_1363,N_108,N_797);
or U1364 (N_1364,N_1031,N_25);
or U1365 (N_1365,N_677,N_78);
nand U1366 (N_1366,N_806,N_197);
nor U1367 (N_1367,N_28,N_621);
or U1368 (N_1368,N_611,N_556);
and U1369 (N_1369,N_771,N_768);
and U1370 (N_1370,N_519,N_194);
nand U1371 (N_1371,N_185,N_555);
nor U1372 (N_1372,N_822,N_19);
and U1373 (N_1373,N_957,N_655);
and U1374 (N_1374,N_1065,N_160);
and U1375 (N_1375,N_863,N_991);
nand U1376 (N_1376,N_919,N_445);
nand U1377 (N_1377,N_265,N_159);
nand U1378 (N_1378,N_193,N_644);
nand U1379 (N_1379,N_1047,N_1087);
xor U1380 (N_1380,N_649,N_1043);
or U1381 (N_1381,N_675,N_706);
xnor U1382 (N_1382,N_709,N_1);
nand U1383 (N_1383,N_468,N_172);
xnor U1384 (N_1384,N_130,N_291);
nor U1385 (N_1385,N_813,N_1041);
nand U1386 (N_1386,N_374,N_181);
nor U1387 (N_1387,N_1018,N_1239);
xnor U1388 (N_1388,N_584,N_1232);
xnor U1389 (N_1389,N_1150,N_313);
or U1390 (N_1390,N_50,N_575);
nand U1391 (N_1391,N_71,N_1074);
nor U1392 (N_1392,N_695,N_380);
nor U1393 (N_1393,N_29,N_1019);
nand U1394 (N_1394,N_13,N_470);
nand U1395 (N_1395,N_893,N_859);
nand U1396 (N_1396,N_937,N_1040);
or U1397 (N_1397,N_438,N_638);
and U1398 (N_1398,N_1084,N_200);
nand U1399 (N_1399,N_1243,N_399);
or U1400 (N_1400,N_100,N_724);
nand U1401 (N_1401,N_997,N_1063);
nor U1402 (N_1402,N_103,N_418);
xor U1403 (N_1403,N_969,N_723);
and U1404 (N_1404,N_585,N_40);
and U1405 (N_1405,N_582,N_1190);
nor U1406 (N_1406,N_832,N_965);
nor U1407 (N_1407,N_461,N_30);
nor U1408 (N_1408,N_849,N_643);
and U1409 (N_1409,N_397,N_1135);
or U1410 (N_1410,N_577,N_98);
nand U1411 (N_1411,N_967,N_668);
xnor U1412 (N_1412,N_310,N_1219);
xnor U1413 (N_1413,N_1143,N_1179);
nor U1414 (N_1414,N_623,N_484);
and U1415 (N_1415,N_93,N_978);
xnor U1416 (N_1416,N_549,N_1113);
xnor U1417 (N_1417,N_987,N_400);
nand U1418 (N_1418,N_1128,N_1153);
nand U1419 (N_1419,N_280,N_398);
and U1420 (N_1420,N_412,N_650);
or U1421 (N_1421,N_713,N_63);
or U1422 (N_1422,N_1025,N_304);
nor U1423 (N_1423,N_536,N_866);
nand U1424 (N_1424,N_186,N_780);
xor U1425 (N_1425,N_444,N_744);
nor U1426 (N_1426,N_494,N_217);
nand U1427 (N_1427,N_535,N_680);
nand U1428 (N_1428,N_388,N_823);
nand U1429 (N_1429,N_915,N_880);
and U1430 (N_1430,N_387,N_659);
or U1431 (N_1431,N_615,N_735);
or U1432 (N_1432,N_1091,N_1157);
xnor U1433 (N_1433,N_403,N_1221);
nand U1434 (N_1434,N_531,N_772);
and U1435 (N_1435,N_188,N_1007);
or U1436 (N_1436,N_109,N_731);
nor U1437 (N_1437,N_175,N_673);
and U1438 (N_1438,N_297,N_602);
nor U1439 (N_1439,N_1136,N_318);
and U1440 (N_1440,N_760,N_222);
xor U1441 (N_1441,N_110,N_64);
nand U1442 (N_1442,N_456,N_176);
and U1443 (N_1443,N_292,N_3);
xor U1444 (N_1444,N_588,N_190);
nor U1445 (N_1445,N_571,N_993);
and U1446 (N_1446,N_756,N_700);
xor U1447 (N_1447,N_852,N_933);
xor U1448 (N_1448,N_202,N_38);
nor U1449 (N_1449,N_87,N_566);
nand U1450 (N_1450,N_68,N_701);
xor U1451 (N_1451,N_816,N_947);
nand U1452 (N_1452,N_1098,N_951);
nor U1453 (N_1453,N_1148,N_192);
and U1454 (N_1454,N_630,N_505);
or U1455 (N_1455,N_1201,N_562);
nand U1456 (N_1456,N_4,N_708);
or U1457 (N_1457,N_946,N_620);
nor U1458 (N_1458,N_1024,N_629);
or U1459 (N_1459,N_384,N_281);
and U1460 (N_1460,N_736,N_1093);
xor U1461 (N_1461,N_994,N_6);
xor U1462 (N_1462,N_163,N_977);
nor U1463 (N_1463,N_1053,N_721);
and U1464 (N_1464,N_689,N_858);
nor U1465 (N_1465,N_1035,N_392);
nand U1466 (N_1466,N_943,N_830);
and U1467 (N_1467,N_634,N_563);
or U1468 (N_1468,N_962,N_36);
nand U1469 (N_1469,N_196,N_106);
nor U1470 (N_1470,N_569,N_321);
or U1471 (N_1471,N_803,N_322);
or U1472 (N_1472,N_476,N_1071);
nor U1473 (N_1473,N_836,N_587);
or U1474 (N_1474,N_914,N_69);
nor U1475 (N_1475,N_212,N_1139);
nor U1476 (N_1476,N_317,N_323);
nand U1477 (N_1477,N_610,N_1107);
nor U1478 (N_1478,N_776,N_1077);
xnor U1479 (N_1479,N_1223,N_86);
xnor U1480 (N_1480,N_794,N_57);
and U1481 (N_1481,N_27,N_204);
nand U1482 (N_1482,N_511,N_157);
nand U1483 (N_1483,N_1195,N_299);
nor U1484 (N_1484,N_24,N_295);
xnor U1485 (N_1485,N_7,N_210);
or U1486 (N_1486,N_277,N_309);
and U1487 (N_1487,N_910,N_67);
xor U1488 (N_1488,N_402,N_409);
xor U1489 (N_1489,N_781,N_178);
nor U1490 (N_1490,N_653,N_840);
xor U1491 (N_1491,N_1202,N_283);
nand U1492 (N_1492,N_793,N_118);
nor U1493 (N_1493,N_284,N_847);
nor U1494 (N_1494,N_91,N_1215);
nand U1495 (N_1495,N_201,N_759);
and U1496 (N_1496,N_572,N_594);
or U1497 (N_1497,N_164,N_395);
xnor U1498 (N_1498,N_678,N_1070);
and U1499 (N_1499,N_11,N_522);
xnor U1500 (N_1500,N_922,N_815);
nand U1501 (N_1501,N_989,N_970);
or U1502 (N_1502,N_589,N_261);
and U1503 (N_1503,N_1173,N_934);
xnor U1504 (N_1504,N_82,N_829);
xnor U1505 (N_1505,N_1214,N_10);
xor U1506 (N_1506,N_458,N_351);
xnor U1507 (N_1507,N_601,N_302);
nor U1508 (N_1508,N_726,N_260);
nor U1509 (N_1509,N_757,N_1100);
and U1510 (N_1510,N_900,N_631);
xnor U1511 (N_1511,N_1187,N_853);
nand U1512 (N_1512,N_1154,N_891);
or U1513 (N_1513,N_676,N_618);
xor U1514 (N_1514,N_553,N_606);
and U1515 (N_1515,N_208,N_609);
nor U1516 (N_1516,N_1204,N_1069);
and U1517 (N_1517,N_382,N_389);
and U1518 (N_1518,N_1152,N_1017);
and U1519 (N_1519,N_533,N_952);
xor U1520 (N_1520,N_1014,N_499);
xor U1521 (N_1521,N_1122,N_908);
or U1522 (N_1522,N_143,N_1111);
xor U1523 (N_1523,N_1164,N_766);
nor U1524 (N_1524,N_405,N_258);
nor U1525 (N_1525,N_406,N_765);
or U1526 (N_1526,N_839,N_96);
or U1527 (N_1527,N_593,N_912);
nand U1528 (N_1528,N_521,N_205);
nand U1529 (N_1529,N_1196,N_213);
xnor U1530 (N_1530,N_439,N_819);
or U1531 (N_1531,N_672,N_1171);
and U1532 (N_1532,N_1210,N_331);
and U1533 (N_1533,N_913,N_39);
nand U1534 (N_1534,N_247,N_479);
nor U1535 (N_1535,N_121,N_428);
xnor U1536 (N_1536,N_637,N_1170);
xor U1537 (N_1537,N_383,N_1012);
or U1538 (N_1538,N_122,N_911);
or U1539 (N_1539,N_895,N_269);
nand U1540 (N_1540,N_316,N_1052);
xor U1541 (N_1541,N_287,N_541);
xor U1542 (N_1542,N_264,N_864);
xor U1543 (N_1543,N_300,N_907);
or U1544 (N_1544,N_1189,N_1048);
and U1545 (N_1545,N_537,N_72);
nand U1546 (N_1546,N_293,N_349);
or U1547 (N_1547,N_92,N_918);
or U1548 (N_1548,N_203,N_407);
nand U1549 (N_1549,N_361,N_750);
or U1550 (N_1550,N_855,N_831);
or U1551 (N_1551,N_921,N_570);
nor U1552 (N_1552,N_1126,N_117);
xnor U1553 (N_1553,N_254,N_294);
or U1554 (N_1554,N_481,N_230);
and U1555 (N_1555,N_385,N_54);
nand U1556 (N_1556,N_1178,N_1155);
nor U1557 (N_1557,N_906,N_705);
nand U1558 (N_1558,N_740,N_232);
or U1559 (N_1559,N_70,N_1220);
nand U1560 (N_1560,N_421,N_436);
or U1561 (N_1561,N_333,N_691);
nor U1562 (N_1562,N_755,N_179);
and U1563 (N_1563,N_717,N_37);
and U1564 (N_1564,N_661,N_329);
nor U1565 (N_1565,N_315,N_1099);
and U1566 (N_1566,N_378,N_353);
nor U1567 (N_1567,N_339,N_20);
and U1568 (N_1568,N_838,N_560);
or U1569 (N_1569,N_328,N_464);
nand U1570 (N_1570,N_42,N_888);
or U1571 (N_1571,N_534,N_105);
nor U1572 (N_1572,N_21,N_1163);
nand U1573 (N_1573,N_66,N_1227);
nor U1574 (N_1574,N_111,N_312);
nand U1575 (N_1575,N_507,N_552);
nor U1576 (N_1576,N_920,N_263);
nand U1577 (N_1577,N_927,N_1217);
or U1578 (N_1578,N_658,N_1209);
nand U1579 (N_1579,N_1090,N_251);
nor U1580 (N_1580,N_154,N_237);
nor U1581 (N_1581,N_1238,N_55);
and U1582 (N_1582,N_640,N_234);
nor U1583 (N_1583,N_460,N_718);
nor U1584 (N_1584,N_207,N_990);
and U1585 (N_1585,N_85,N_338);
nand U1586 (N_1586,N_1064,N_727);
nand U1587 (N_1587,N_169,N_404);
or U1588 (N_1588,N_741,N_125);
nand U1589 (N_1589,N_953,N_767);
or U1590 (N_1590,N_639,N_662);
nor U1591 (N_1591,N_580,N_925);
or U1592 (N_1592,N_567,N_1059);
and U1593 (N_1593,N_340,N_651);
xor U1594 (N_1594,N_1051,N_115);
nand U1595 (N_1595,N_31,N_1199);
nor U1596 (N_1596,N_414,N_450);
or U1597 (N_1597,N_423,N_1000);
and U1598 (N_1598,N_140,N_504);
and U1599 (N_1599,N_1081,N_811);
or U1600 (N_1600,N_457,N_787);
nand U1601 (N_1601,N_1029,N_748);
nor U1602 (N_1602,N_929,N_1108);
or U1603 (N_1603,N_871,N_788);
xor U1604 (N_1604,N_754,N_424);
or U1605 (N_1605,N_1022,N_465);
or U1606 (N_1606,N_478,N_88);
nand U1607 (N_1607,N_762,N_451);
nand U1608 (N_1608,N_1055,N_289);
nor U1609 (N_1609,N_664,N_1142);
nor U1610 (N_1610,N_848,N_616);
nand U1611 (N_1611,N_346,N_683);
or U1612 (N_1612,N_667,N_802);
or U1613 (N_1613,N_512,N_648);
or U1614 (N_1614,N_1061,N_818);
and U1615 (N_1615,N_669,N_645);
or U1616 (N_1616,N_235,N_660);
nand U1617 (N_1617,N_495,N_826);
or U1618 (N_1618,N_1208,N_1233);
nand U1619 (N_1619,N_182,N_49);
nor U1620 (N_1620,N_228,N_34);
and U1621 (N_1621,N_327,N_123);
xor U1622 (N_1622,N_1198,N_391);
or U1623 (N_1623,N_370,N_5);
xor U1624 (N_1624,N_995,N_475);
and U1625 (N_1625,N_147,N_598);
nand U1626 (N_1626,N_998,N_627);
xor U1627 (N_1627,N_48,N_262);
nor U1628 (N_1628,N_311,N_320);
nor U1629 (N_1629,N_1121,N_32);
and U1630 (N_1630,N_530,N_518);
and U1631 (N_1631,N_545,N_2);
nand U1632 (N_1632,N_959,N_1249);
nand U1633 (N_1633,N_646,N_796);
nand U1634 (N_1634,N_490,N_752);
nand U1635 (N_1635,N_131,N_1182);
and U1636 (N_1636,N_690,N_124);
nand U1637 (N_1637,N_1188,N_1205);
nand U1638 (N_1638,N_835,N_102);
nand U1639 (N_1639,N_255,N_1235);
and U1640 (N_1640,N_101,N_434);
nor U1641 (N_1641,N_1023,N_791);
and U1642 (N_1642,N_948,N_1129);
xor U1643 (N_1643,N_411,N_1060);
or U1644 (N_1644,N_949,N_687);
or U1645 (N_1645,N_156,N_347);
or U1646 (N_1646,N_62,N_113);
or U1647 (N_1647,N_41,N_358);
and U1648 (N_1648,N_1149,N_558);
or U1649 (N_1649,N_1082,N_1118);
xor U1650 (N_1650,N_692,N_274);
nor U1651 (N_1651,N_15,N_1095);
and U1652 (N_1652,N_1075,N_1030);
or U1653 (N_1653,N_865,N_454);
and U1654 (N_1654,N_1216,N_18);
nand U1655 (N_1655,N_1165,N_366);
or U1656 (N_1656,N_462,N_116);
or U1657 (N_1657,N_128,N_905);
or U1658 (N_1658,N_441,N_245);
xnor U1659 (N_1659,N_568,N_973);
or U1660 (N_1660,N_286,N_1088);
nor U1661 (N_1661,N_682,N_273);
and U1662 (N_1662,N_97,N_332);
nor U1663 (N_1663,N_225,N_1230);
or U1664 (N_1664,N_1192,N_95);
xnor U1665 (N_1665,N_278,N_1146);
or U1666 (N_1666,N_1123,N_90);
xor U1667 (N_1667,N_786,N_153);
and U1668 (N_1668,N_857,N_16);
nor U1669 (N_1669,N_820,N_1013);
and U1670 (N_1670,N_1057,N_854);
nor U1671 (N_1671,N_1026,N_257);
nand U1672 (N_1672,N_307,N_216);
xnor U1673 (N_1673,N_579,N_1044);
and U1674 (N_1674,N_1101,N_633);
xnor U1675 (N_1675,N_890,N_1166);
nor U1676 (N_1676,N_306,N_44);
nand U1677 (N_1677,N_972,N_954);
nand U1678 (N_1678,N_334,N_1197);
or U1679 (N_1679,N_266,N_1067);
and U1680 (N_1680,N_142,N_641);
and U1681 (N_1681,N_699,N_842);
or U1682 (N_1682,N_1159,N_1032);
nor U1683 (N_1683,N_860,N_980);
or U1684 (N_1684,N_246,N_626);
nand U1685 (N_1685,N_817,N_500);
xor U1686 (N_1686,N_149,N_1237);
nor U1687 (N_1687,N_80,N_875);
nor U1688 (N_1688,N_344,N_843);
nand U1689 (N_1689,N_372,N_416);
nand U1690 (N_1690,N_846,N_357);
nand U1691 (N_1691,N_1072,N_74);
and U1692 (N_1692,N_155,N_719);
and U1693 (N_1693,N_716,N_694);
or U1694 (N_1694,N_1076,N_119);
and U1695 (N_1695,N_523,N_1086);
or U1696 (N_1696,N_1046,N_559);
and U1697 (N_1697,N_1124,N_1103);
or U1698 (N_1698,N_47,N_1218);
nor U1699 (N_1699,N_151,N_684);
or U1700 (N_1700,N_1240,N_501);
nand U1701 (N_1701,N_961,N_206);
or U1702 (N_1702,N_1222,N_1169);
or U1703 (N_1703,N_976,N_1094);
or U1704 (N_1704,N_174,N_674);
nor U1705 (N_1705,N_227,N_1003);
or U1706 (N_1706,N_1045,N_527);
and U1707 (N_1707,N_764,N_1110);
and U1708 (N_1708,N_590,N_342);
and U1709 (N_1709,N_104,N_209);
nand U1710 (N_1710,N_841,N_1049);
nor U1711 (N_1711,N_904,N_784);
or U1712 (N_1712,N_502,N_314);
and U1713 (N_1713,N_599,N_1134);
xnor U1714 (N_1714,N_785,N_75);
and U1715 (N_1715,N_137,N_635);
nor U1716 (N_1716,N_729,N_1009);
nand U1717 (N_1717,N_548,N_168);
nand U1718 (N_1718,N_426,N_887);
or U1719 (N_1719,N_1005,N_878);
or U1720 (N_1720,N_173,N_1109);
nor U1721 (N_1721,N_165,N_711);
or U1722 (N_1722,N_517,N_187);
xnor U1723 (N_1723,N_268,N_61);
and U1724 (N_1724,N_369,N_430);
xnor U1725 (N_1725,N_1115,N_319);
or U1726 (N_1726,N_221,N_758);
nor U1727 (N_1727,N_138,N_167);
and U1728 (N_1728,N_244,N_1008);
xnor U1729 (N_1729,N_270,N_23);
xnor U1730 (N_1730,N_715,N_1034);
nor U1731 (N_1731,N_1042,N_0);
or U1732 (N_1732,N_442,N_837);
xnor U1733 (N_1733,N_547,N_751);
or U1734 (N_1734,N_26,N_783);
xnor U1735 (N_1735,N_551,N_496);
nand U1736 (N_1736,N_488,N_433);
and U1737 (N_1737,N_681,N_1172);
or U1738 (N_1738,N_364,N_1011);
or U1739 (N_1739,N_882,N_177);
nand U1740 (N_1740,N_359,N_219);
or U1741 (N_1741,N_557,N_1248);
nand U1742 (N_1742,N_1016,N_466);
or U1743 (N_1743,N_877,N_1033);
nand U1744 (N_1744,N_810,N_455);
xor U1745 (N_1745,N_248,N_1079);
nand U1746 (N_1746,N_770,N_367);
and U1747 (N_1747,N_493,N_529);
or U1748 (N_1748,N_162,N_345);
nor U1749 (N_1749,N_812,N_79);
or U1750 (N_1750,N_132,N_516);
nor U1751 (N_1751,N_769,N_480);
nor U1752 (N_1752,N_543,N_1130);
or U1753 (N_1753,N_393,N_238);
xnor U1754 (N_1754,N_693,N_1080);
xor U1755 (N_1755,N_1015,N_170);
and U1756 (N_1756,N_821,N_1245);
xnor U1757 (N_1757,N_1156,N_1068);
nor U1758 (N_1758,N_869,N_540);
xor U1759 (N_1759,N_89,N_1213);
xnor U1760 (N_1760,N_1027,N_1137);
nor U1761 (N_1761,N_1085,N_824);
nand U1762 (N_1762,N_1140,N_613);
and U1763 (N_1763,N_1203,N_355);
and U1764 (N_1764,N_795,N_1117);
or U1765 (N_1765,N_958,N_415);
or U1766 (N_1766,N_224,N_737);
nor U1767 (N_1767,N_1004,N_352);
nand U1768 (N_1768,N_446,N_792);
and U1769 (N_1769,N_1078,N_497);
nand U1770 (N_1770,N_1073,N_419);
and U1771 (N_1771,N_685,N_625);
xnor U1772 (N_1772,N_305,N_463);
nor U1773 (N_1773,N_704,N_325);
or U1774 (N_1774,N_940,N_647);
nor U1775 (N_1775,N_1186,N_889);
and U1776 (N_1776,N_1177,N_377);
or U1777 (N_1777,N_901,N_898);
nor U1778 (N_1778,N_435,N_514);
or U1779 (N_1779,N_449,N_76);
xor U1780 (N_1780,N_1021,N_146);
nand U1781 (N_1781,N_503,N_926);
and U1782 (N_1782,N_348,N_81);
xnor U1783 (N_1783,N_805,N_586);
nand U1784 (N_1784,N_243,N_1056);
nand U1785 (N_1785,N_1193,N_612);
nand U1786 (N_1786,N_554,N_564);
and U1787 (N_1787,N_881,N_1062);
nand U1788 (N_1788,N_671,N_1006);
or U1789 (N_1789,N_356,N_939);
nand U1790 (N_1790,N_595,N_712);
and U1791 (N_1791,N_739,N_565);
xnor U1792 (N_1792,N_1092,N_782);
or U1793 (N_1793,N_326,N_343);
nor U1794 (N_1794,N_526,N_1184);
nor U1795 (N_1795,N_872,N_975);
or U1796 (N_1796,N_999,N_1141);
xor U1797 (N_1797,N_259,N_960);
and U1798 (N_1798,N_923,N_1144);
nand U1799 (N_1799,N_886,N_654);
nor U1800 (N_1800,N_171,N_198);
or U1801 (N_1801,N_35,N_703);
xnor U1802 (N_1802,N_636,N_242);
or U1803 (N_1803,N_1207,N_800);
xnor U1804 (N_1804,N_1241,N_410);
xor U1805 (N_1805,N_396,N_477);
and U1806 (N_1806,N_1175,N_239);
or U1807 (N_1807,N_622,N_532);
nor U1808 (N_1808,N_1104,N_1133);
or U1809 (N_1809,N_112,N_544);
and U1810 (N_1810,N_223,N_139);
and U1811 (N_1811,N_899,N_166);
or U1812 (N_1812,N_241,N_1147);
nand U1813 (N_1813,N_657,N_763);
nand U1814 (N_1814,N_1185,N_966);
nand U1815 (N_1815,N_538,N_12);
nand U1816 (N_1816,N_607,N_240);
and U1817 (N_1817,N_136,N_592);
nand U1818 (N_1818,N_546,N_928);
or U1819 (N_1819,N_665,N_679);
xnor U1820 (N_1820,N_483,N_360);
or U1821 (N_1821,N_1160,N_191);
nand U1822 (N_1822,N_373,N_1020);
nor U1823 (N_1823,N_884,N_1168);
or U1824 (N_1824,N_814,N_303);
and U1825 (N_1825,N_1112,N_425);
and U1826 (N_1826,N_941,N_624);
xor U1827 (N_1827,N_873,N_17);
or U1828 (N_1828,N_778,N_938);
nor U1829 (N_1829,N_1054,N_218);
xnor U1830 (N_1830,N_1242,N_827);
and U1831 (N_1831,N_696,N_59);
or U1832 (N_1832,N_1236,N_608);
xor U1833 (N_1833,N_459,N_510);
nor U1834 (N_1834,N_429,N_1161);
nand U1835 (N_1835,N_471,N_148);
xnor U1836 (N_1836,N_1010,N_894);
or U1837 (N_1837,N_1028,N_376);
xnor U1838 (N_1838,N_996,N_491);
nor U1839 (N_1839,N_964,N_573);
and U1840 (N_1840,N_473,N_1212);
or U1841 (N_1841,N_298,N_513);
nor U1842 (N_1842,N_1225,N_870);
and U1843 (N_1843,N_909,N_448);
nand U1844 (N_1844,N_702,N_386);
or U1845 (N_1845,N_746,N_1162);
and U1846 (N_1846,N_652,N_935);
and U1847 (N_1847,N_229,N_974);
xor U1848 (N_1848,N_542,N_1229);
and U1849 (N_1849,N_874,N_663);
nand U1850 (N_1850,N_774,N_688);
nand U1851 (N_1851,N_250,N_135);
and U1852 (N_1852,N_271,N_1037);
or U1853 (N_1853,N_515,N_773);
nor U1854 (N_1854,N_604,N_290);
or U1855 (N_1855,N_249,N_467);
nand U1856 (N_1856,N_550,N_632);
xor U1857 (N_1857,N_1096,N_324);
nand U1858 (N_1858,N_528,N_341);
or U1859 (N_1859,N_508,N_252);
xor U1860 (N_1860,N_734,N_1105);
nand U1861 (N_1861,N_656,N_1036);
nand U1862 (N_1862,N_807,N_1114);
nand U1863 (N_1863,N_8,N_336);
nor U1864 (N_1864,N_134,N_288);
xor U1865 (N_1865,N_720,N_561);
nor U1866 (N_1866,N_1106,N_350);
nor U1867 (N_1867,N_883,N_525);
and U1868 (N_1868,N_1224,N_520);
xor U1869 (N_1869,N_524,N_749);
xor U1870 (N_1870,N_743,N_950);
or U1871 (N_1871,N_381,N_472);
nand U1872 (N_1872,N_487,N_1083);
nor U1873 (N_1873,N_236,N_408);
and U1874 (N_1874,N_916,N_597);
and U1875 (N_1875,N_63,N_1238);
xor U1876 (N_1876,N_412,N_111);
nor U1877 (N_1877,N_1039,N_305);
nor U1878 (N_1878,N_362,N_327);
nand U1879 (N_1879,N_570,N_563);
or U1880 (N_1880,N_783,N_459);
and U1881 (N_1881,N_756,N_169);
and U1882 (N_1882,N_886,N_1154);
nor U1883 (N_1883,N_641,N_1077);
and U1884 (N_1884,N_1221,N_1000);
nand U1885 (N_1885,N_974,N_1136);
and U1886 (N_1886,N_490,N_468);
xor U1887 (N_1887,N_1188,N_181);
or U1888 (N_1888,N_542,N_1063);
nor U1889 (N_1889,N_882,N_612);
nand U1890 (N_1890,N_672,N_19);
nand U1891 (N_1891,N_518,N_614);
and U1892 (N_1892,N_846,N_11);
nand U1893 (N_1893,N_960,N_745);
and U1894 (N_1894,N_762,N_865);
and U1895 (N_1895,N_1077,N_1069);
and U1896 (N_1896,N_777,N_527);
and U1897 (N_1897,N_904,N_1114);
nor U1898 (N_1898,N_644,N_615);
and U1899 (N_1899,N_190,N_1183);
nor U1900 (N_1900,N_865,N_1143);
nand U1901 (N_1901,N_1161,N_56);
and U1902 (N_1902,N_787,N_169);
nor U1903 (N_1903,N_1171,N_947);
nand U1904 (N_1904,N_293,N_866);
xnor U1905 (N_1905,N_1244,N_1201);
or U1906 (N_1906,N_447,N_165);
and U1907 (N_1907,N_680,N_526);
xor U1908 (N_1908,N_511,N_1188);
nand U1909 (N_1909,N_657,N_864);
nor U1910 (N_1910,N_225,N_601);
nor U1911 (N_1911,N_321,N_843);
xor U1912 (N_1912,N_1246,N_757);
nand U1913 (N_1913,N_1248,N_35);
nor U1914 (N_1914,N_235,N_66);
or U1915 (N_1915,N_425,N_92);
and U1916 (N_1916,N_1052,N_915);
nor U1917 (N_1917,N_729,N_1024);
xor U1918 (N_1918,N_861,N_476);
nand U1919 (N_1919,N_929,N_799);
nand U1920 (N_1920,N_489,N_1190);
nand U1921 (N_1921,N_1201,N_938);
or U1922 (N_1922,N_1002,N_785);
nor U1923 (N_1923,N_171,N_1153);
nand U1924 (N_1924,N_724,N_940);
and U1925 (N_1925,N_812,N_1089);
and U1926 (N_1926,N_809,N_127);
and U1927 (N_1927,N_347,N_213);
nand U1928 (N_1928,N_636,N_621);
nand U1929 (N_1929,N_61,N_770);
or U1930 (N_1930,N_788,N_1085);
nand U1931 (N_1931,N_398,N_475);
xor U1932 (N_1932,N_986,N_606);
xor U1933 (N_1933,N_436,N_810);
nand U1934 (N_1934,N_1062,N_183);
nor U1935 (N_1935,N_761,N_41);
or U1936 (N_1936,N_1242,N_998);
nor U1937 (N_1937,N_222,N_861);
xnor U1938 (N_1938,N_814,N_447);
nand U1939 (N_1939,N_1205,N_758);
nor U1940 (N_1940,N_175,N_340);
or U1941 (N_1941,N_1183,N_362);
xnor U1942 (N_1942,N_989,N_1246);
xor U1943 (N_1943,N_566,N_925);
nor U1944 (N_1944,N_428,N_724);
nand U1945 (N_1945,N_1227,N_1105);
or U1946 (N_1946,N_880,N_1247);
and U1947 (N_1947,N_301,N_1096);
nand U1948 (N_1948,N_1081,N_271);
nor U1949 (N_1949,N_1066,N_438);
or U1950 (N_1950,N_750,N_512);
nor U1951 (N_1951,N_279,N_658);
and U1952 (N_1952,N_543,N_1213);
and U1953 (N_1953,N_940,N_562);
and U1954 (N_1954,N_607,N_1219);
xnor U1955 (N_1955,N_77,N_1144);
and U1956 (N_1956,N_191,N_214);
xnor U1957 (N_1957,N_643,N_693);
xor U1958 (N_1958,N_595,N_1050);
xor U1959 (N_1959,N_960,N_829);
nor U1960 (N_1960,N_23,N_397);
nor U1961 (N_1961,N_441,N_1106);
xor U1962 (N_1962,N_503,N_750);
xor U1963 (N_1963,N_974,N_730);
or U1964 (N_1964,N_630,N_1221);
nand U1965 (N_1965,N_1113,N_843);
xor U1966 (N_1966,N_666,N_850);
and U1967 (N_1967,N_1113,N_619);
nor U1968 (N_1968,N_1094,N_537);
xnor U1969 (N_1969,N_533,N_896);
nand U1970 (N_1970,N_368,N_971);
xor U1971 (N_1971,N_906,N_912);
or U1972 (N_1972,N_615,N_260);
nand U1973 (N_1973,N_1191,N_77);
nand U1974 (N_1974,N_944,N_521);
nor U1975 (N_1975,N_727,N_364);
xor U1976 (N_1976,N_1033,N_398);
nand U1977 (N_1977,N_296,N_1163);
nand U1978 (N_1978,N_1191,N_123);
or U1979 (N_1979,N_336,N_470);
nor U1980 (N_1980,N_558,N_965);
and U1981 (N_1981,N_641,N_961);
nand U1982 (N_1982,N_708,N_966);
and U1983 (N_1983,N_1226,N_72);
nand U1984 (N_1984,N_44,N_1199);
xor U1985 (N_1985,N_1182,N_477);
nand U1986 (N_1986,N_866,N_997);
and U1987 (N_1987,N_279,N_972);
nor U1988 (N_1988,N_951,N_735);
and U1989 (N_1989,N_142,N_216);
nor U1990 (N_1990,N_146,N_886);
nand U1991 (N_1991,N_832,N_490);
xnor U1992 (N_1992,N_640,N_1002);
nand U1993 (N_1993,N_546,N_679);
nor U1994 (N_1994,N_971,N_364);
or U1995 (N_1995,N_775,N_1078);
xnor U1996 (N_1996,N_568,N_1000);
nand U1997 (N_1997,N_700,N_896);
nand U1998 (N_1998,N_1105,N_516);
or U1999 (N_1999,N_1185,N_1236);
or U2000 (N_2000,N_180,N_807);
nand U2001 (N_2001,N_53,N_667);
or U2002 (N_2002,N_431,N_162);
nand U2003 (N_2003,N_1046,N_969);
nor U2004 (N_2004,N_346,N_299);
and U2005 (N_2005,N_1093,N_500);
xor U2006 (N_2006,N_650,N_390);
nand U2007 (N_2007,N_584,N_705);
nand U2008 (N_2008,N_778,N_438);
nand U2009 (N_2009,N_1062,N_644);
nand U2010 (N_2010,N_313,N_352);
nor U2011 (N_2011,N_394,N_751);
or U2012 (N_2012,N_662,N_443);
nor U2013 (N_2013,N_131,N_648);
xnor U2014 (N_2014,N_743,N_568);
xnor U2015 (N_2015,N_438,N_279);
nand U2016 (N_2016,N_1046,N_616);
and U2017 (N_2017,N_649,N_1239);
xor U2018 (N_2018,N_1127,N_1020);
xnor U2019 (N_2019,N_384,N_317);
nand U2020 (N_2020,N_747,N_1038);
or U2021 (N_2021,N_345,N_1198);
nand U2022 (N_2022,N_658,N_443);
or U2023 (N_2023,N_527,N_314);
or U2024 (N_2024,N_519,N_986);
xnor U2025 (N_2025,N_458,N_479);
and U2026 (N_2026,N_247,N_17);
and U2027 (N_2027,N_946,N_693);
nand U2028 (N_2028,N_321,N_123);
nor U2029 (N_2029,N_783,N_693);
or U2030 (N_2030,N_1115,N_278);
or U2031 (N_2031,N_543,N_87);
or U2032 (N_2032,N_986,N_442);
nor U2033 (N_2033,N_615,N_147);
xnor U2034 (N_2034,N_1037,N_1222);
nor U2035 (N_2035,N_148,N_550);
and U2036 (N_2036,N_497,N_1035);
xor U2037 (N_2037,N_508,N_414);
or U2038 (N_2038,N_1142,N_1061);
nand U2039 (N_2039,N_1166,N_93);
and U2040 (N_2040,N_445,N_656);
and U2041 (N_2041,N_577,N_907);
nor U2042 (N_2042,N_1174,N_1129);
xor U2043 (N_2043,N_1174,N_819);
or U2044 (N_2044,N_1183,N_807);
and U2045 (N_2045,N_1239,N_377);
xor U2046 (N_2046,N_370,N_1208);
nand U2047 (N_2047,N_124,N_28);
nand U2048 (N_2048,N_760,N_355);
nand U2049 (N_2049,N_1112,N_103);
and U2050 (N_2050,N_995,N_1190);
and U2051 (N_2051,N_35,N_54);
and U2052 (N_2052,N_438,N_28);
or U2053 (N_2053,N_566,N_1192);
nor U2054 (N_2054,N_342,N_558);
nor U2055 (N_2055,N_1092,N_1012);
nor U2056 (N_2056,N_366,N_828);
xor U2057 (N_2057,N_225,N_607);
nor U2058 (N_2058,N_154,N_382);
and U2059 (N_2059,N_1168,N_588);
or U2060 (N_2060,N_1202,N_139);
and U2061 (N_2061,N_153,N_352);
and U2062 (N_2062,N_1145,N_49);
and U2063 (N_2063,N_1097,N_684);
xnor U2064 (N_2064,N_145,N_894);
nand U2065 (N_2065,N_771,N_25);
nor U2066 (N_2066,N_1227,N_517);
nor U2067 (N_2067,N_817,N_0);
or U2068 (N_2068,N_957,N_809);
or U2069 (N_2069,N_788,N_173);
or U2070 (N_2070,N_539,N_279);
and U2071 (N_2071,N_666,N_547);
nor U2072 (N_2072,N_1174,N_223);
and U2073 (N_2073,N_741,N_185);
nand U2074 (N_2074,N_1011,N_752);
nand U2075 (N_2075,N_403,N_684);
xor U2076 (N_2076,N_1006,N_812);
xor U2077 (N_2077,N_157,N_1140);
nor U2078 (N_2078,N_494,N_5);
or U2079 (N_2079,N_172,N_657);
xor U2080 (N_2080,N_1227,N_76);
or U2081 (N_2081,N_820,N_542);
xnor U2082 (N_2082,N_1154,N_938);
xor U2083 (N_2083,N_1220,N_322);
or U2084 (N_2084,N_1073,N_964);
or U2085 (N_2085,N_801,N_402);
and U2086 (N_2086,N_559,N_279);
nor U2087 (N_2087,N_155,N_280);
nor U2088 (N_2088,N_278,N_1003);
nand U2089 (N_2089,N_567,N_261);
nor U2090 (N_2090,N_944,N_211);
or U2091 (N_2091,N_413,N_640);
nor U2092 (N_2092,N_669,N_658);
and U2093 (N_2093,N_1213,N_66);
or U2094 (N_2094,N_75,N_110);
and U2095 (N_2095,N_846,N_463);
and U2096 (N_2096,N_427,N_489);
nor U2097 (N_2097,N_779,N_292);
nand U2098 (N_2098,N_994,N_864);
nand U2099 (N_2099,N_604,N_407);
or U2100 (N_2100,N_610,N_686);
and U2101 (N_2101,N_40,N_891);
or U2102 (N_2102,N_326,N_103);
or U2103 (N_2103,N_227,N_460);
or U2104 (N_2104,N_216,N_1088);
nor U2105 (N_2105,N_614,N_96);
nand U2106 (N_2106,N_994,N_118);
and U2107 (N_2107,N_113,N_1090);
xnor U2108 (N_2108,N_199,N_573);
nand U2109 (N_2109,N_1052,N_184);
or U2110 (N_2110,N_207,N_1213);
xor U2111 (N_2111,N_299,N_399);
nor U2112 (N_2112,N_406,N_59);
or U2113 (N_2113,N_1093,N_769);
or U2114 (N_2114,N_57,N_235);
nand U2115 (N_2115,N_662,N_189);
and U2116 (N_2116,N_644,N_858);
xor U2117 (N_2117,N_483,N_230);
nor U2118 (N_2118,N_635,N_657);
xor U2119 (N_2119,N_232,N_1076);
xor U2120 (N_2120,N_708,N_79);
or U2121 (N_2121,N_1006,N_1005);
nor U2122 (N_2122,N_292,N_1089);
xnor U2123 (N_2123,N_1042,N_1117);
or U2124 (N_2124,N_203,N_1124);
xnor U2125 (N_2125,N_86,N_937);
or U2126 (N_2126,N_1063,N_866);
or U2127 (N_2127,N_23,N_132);
or U2128 (N_2128,N_752,N_72);
or U2129 (N_2129,N_302,N_826);
and U2130 (N_2130,N_205,N_694);
nand U2131 (N_2131,N_135,N_1055);
or U2132 (N_2132,N_77,N_810);
or U2133 (N_2133,N_811,N_1040);
nor U2134 (N_2134,N_406,N_688);
or U2135 (N_2135,N_717,N_1037);
or U2136 (N_2136,N_826,N_824);
nand U2137 (N_2137,N_982,N_1008);
nor U2138 (N_2138,N_370,N_745);
xor U2139 (N_2139,N_1054,N_42);
and U2140 (N_2140,N_850,N_1045);
or U2141 (N_2141,N_665,N_289);
nor U2142 (N_2142,N_1179,N_1165);
or U2143 (N_2143,N_456,N_339);
nor U2144 (N_2144,N_969,N_1118);
nor U2145 (N_2145,N_929,N_668);
nor U2146 (N_2146,N_1080,N_1031);
and U2147 (N_2147,N_746,N_701);
or U2148 (N_2148,N_37,N_285);
nand U2149 (N_2149,N_1144,N_435);
or U2150 (N_2150,N_313,N_424);
and U2151 (N_2151,N_59,N_894);
nor U2152 (N_2152,N_774,N_709);
and U2153 (N_2153,N_780,N_1030);
nor U2154 (N_2154,N_336,N_1028);
nand U2155 (N_2155,N_341,N_991);
nand U2156 (N_2156,N_285,N_25);
nor U2157 (N_2157,N_694,N_543);
xor U2158 (N_2158,N_948,N_584);
nand U2159 (N_2159,N_966,N_607);
or U2160 (N_2160,N_313,N_884);
or U2161 (N_2161,N_41,N_1090);
or U2162 (N_2162,N_1110,N_21);
or U2163 (N_2163,N_358,N_953);
xnor U2164 (N_2164,N_679,N_611);
or U2165 (N_2165,N_751,N_955);
and U2166 (N_2166,N_956,N_688);
and U2167 (N_2167,N_339,N_668);
and U2168 (N_2168,N_1064,N_14);
nand U2169 (N_2169,N_869,N_528);
or U2170 (N_2170,N_198,N_399);
nand U2171 (N_2171,N_68,N_362);
or U2172 (N_2172,N_1085,N_517);
or U2173 (N_2173,N_1020,N_752);
and U2174 (N_2174,N_795,N_61);
nand U2175 (N_2175,N_1220,N_165);
nor U2176 (N_2176,N_910,N_182);
and U2177 (N_2177,N_56,N_244);
nand U2178 (N_2178,N_259,N_93);
nand U2179 (N_2179,N_424,N_1190);
nand U2180 (N_2180,N_55,N_720);
nor U2181 (N_2181,N_115,N_517);
and U2182 (N_2182,N_1244,N_391);
nand U2183 (N_2183,N_210,N_1055);
or U2184 (N_2184,N_346,N_104);
or U2185 (N_2185,N_1067,N_1004);
nand U2186 (N_2186,N_307,N_46);
xnor U2187 (N_2187,N_543,N_378);
nor U2188 (N_2188,N_620,N_575);
nand U2189 (N_2189,N_1108,N_9);
and U2190 (N_2190,N_346,N_309);
or U2191 (N_2191,N_1039,N_326);
nand U2192 (N_2192,N_774,N_649);
xor U2193 (N_2193,N_280,N_1018);
xor U2194 (N_2194,N_598,N_447);
and U2195 (N_2195,N_868,N_190);
nor U2196 (N_2196,N_225,N_411);
or U2197 (N_2197,N_395,N_255);
and U2198 (N_2198,N_1163,N_979);
or U2199 (N_2199,N_666,N_887);
nor U2200 (N_2200,N_1088,N_462);
nor U2201 (N_2201,N_125,N_6);
and U2202 (N_2202,N_380,N_290);
xor U2203 (N_2203,N_617,N_914);
nor U2204 (N_2204,N_122,N_1075);
xor U2205 (N_2205,N_418,N_581);
nor U2206 (N_2206,N_1063,N_91);
nand U2207 (N_2207,N_227,N_394);
nand U2208 (N_2208,N_405,N_219);
and U2209 (N_2209,N_934,N_946);
or U2210 (N_2210,N_1011,N_650);
and U2211 (N_2211,N_516,N_31);
xor U2212 (N_2212,N_741,N_406);
or U2213 (N_2213,N_198,N_485);
or U2214 (N_2214,N_104,N_900);
nor U2215 (N_2215,N_632,N_12);
nand U2216 (N_2216,N_649,N_1117);
nand U2217 (N_2217,N_185,N_418);
xor U2218 (N_2218,N_517,N_1040);
xor U2219 (N_2219,N_1040,N_783);
nand U2220 (N_2220,N_1071,N_1024);
or U2221 (N_2221,N_691,N_1216);
and U2222 (N_2222,N_1040,N_649);
or U2223 (N_2223,N_163,N_1184);
and U2224 (N_2224,N_23,N_461);
nand U2225 (N_2225,N_1108,N_292);
and U2226 (N_2226,N_351,N_212);
nor U2227 (N_2227,N_572,N_1137);
or U2228 (N_2228,N_128,N_916);
or U2229 (N_2229,N_730,N_237);
nor U2230 (N_2230,N_344,N_789);
and U2231 (N_2231,N_84,N_310);
xnor U2232 (N_2232,N_1218,N_667);
and U2233 (N_2233,N_340,N_270);
xor U2234 (N_2234,N_1115,N_643);
or U2235 (N_2235,N_386,N_1068);
nand U2236 (N_2236,N_793,N_182);
or U2237 (N_2237,N_42,N_1176);
nor U2238 (N_2238,N_280,N_278);
and U2239 (N_2239,N_684,N_10);
and U2240 (N_2240,N_126,N_634);
or U2241 (N_2241,N_60,N_776);
nand U2242 (N_2242,N_689,N_772);
nand U2243 (N_2243,N_897,N_829);
or U2244 (N_2244,N_321,N_527);
and U2245 (N_2245,N_967,N_834);
or U2246 (N_2246,N_5,N_727);
or U2247 (N_2247,N_569,N_731);
xnor U2248 (N_2248,N_150,N_921);
and U2249 (N_2249,N_537,N_522);
nor U2250 (N_2250,N_284,N_127);
or U2251 (N_2251,N_120,N_500);
nor U2252 (N_2252,N_546,N_1022);
nor U2253 (N_2253,N_1064,N_227);
xor U2254 (N_2254,N_72,N_1122);
xnor U2255 (N_2255,N_149,N_1134);
nor U2256 (N_2256,N_320,N_323);
or U2257 (N_2257,N_243,N_1026);
or U2258 (N_2258,N_100,N_1173);
nand U2259 (N_2259,N_727,N_558);
and U2260 (N_2260,N_1247,N_643);
xnor U2261 (N_2261,N_1040,N_677);
xor U2262 (N_2262,N_469,N_249);
xor U2263 (N_2263,N_755,N_1095);
nor U2264 (N_2264,N_727,N_602);
or U2265 (N_2265,N_1115,N_112);
xor U2266 (N_2266,N_67,N_332);
xnor U2267 (N_2267,N_1013,N_922);
nand U2268 (N_2268,N_1039,N_352);
and U2269 (N_2269,N_536,N_887);
or U2270 (N_2270,N_183,N_34);
nand U2271 (N_2271,N_914,N_97);
and U2272 (N_2272,N_372,N_255);
or U2273 (N_2273,N_189,N_469);
and U2274 (N_2274,N_4,N_781);
or U2275 (N_2275,N_858,N_1112);
and U2276 (N_2276,N_684,N_969);
nor U2277 (N_2277,N_1233,N_374);
nor U2278 (N_2278,N_480,N_12);
or U2279 (N_2279,N_929,N_293);
nand U2280 (N_2280,N_658,N_1177);
and U2281 (N_2281,N_506,N_473);
nor U2282 (N_2282,N_689,N_230);
nor U2283 (N_2283,N_518,N_157);
nand U2284 (N_2284,N_1171,N_62);
xor U2285 (N_2285,N_319,N_41);
and U2286 (N_2286,N_181,N_407);
nor U2287 (N_2287,N_461,N_699);
nor U2288 (N_2288,N_849,N_718);
nand U2289 (N_2289,N_224,N_332);
or U2290 (N_2290,N_439,N_207);
nand U2291 (N_2291,N_73,N_1060);
nor U2292 (N_2292,N_468,N_316);
xnor U2293 (N_2293,N_644,N_1140);
or U2294 (N_2294,N_692,N_245);
or U2295 (N_2295,N_802,N_548);
nand U2296 (N_2296,N_1209,N_640);
or U2297 (N_2297,N_85,N_1242);
or U2298 (N_2298,N_643,N_1118);
nor U2299 (N_2299,N_576,N_1133);
xnor U2300 (N_2300,N_572,N_549);
nor U2301 (N_2301,N_355,N_603);
xor U2302 (N_2302,N_1153,N_1154);
nand U2303 (N_2303,N_91,N_98);
xor U2304 (N_2304,N_217,N_998);
xor U2305 (N_2305,N_976,N_745);
nor U2306 (N_2306,N_337,N_347);
nor U2307 (N_2307,N_1208,N_890);
xor U2308 (N_2308,N_1108,N_766);
and U2309 (N_2309,N_1149,N_130);
xnor U2310 (N_2310,N_779,N_611);
xnor U2311 (N_2311,N_914,N_58);
nand U2312 (N_2312,N_784,N_655);
or U2313 (N_2313,N_1229,N_109);
and U2314 (N_2314,N_1,N_666);
nor U2315 (N_2315,N_1011,N_904);
nand U2316 (N_2316,N_1038,N_828);
or U2317 (N_2317,N_1068,N_1083);
nand U2318 (N_2318,N_295,N_14);
and U2319 (N_2319,N_927,N_1051);
nand U2320 (N_2320,N_147,N_1121);
nand U2321 (N_2321,N_637,N_373);
xnor U2322 (N_2322,N_677,N_436);
xnor U2323 (N_2323,N_162,N_859);
or U2324 (N_2324,N_1153,N_947);
nand U2325 (N_2325,N_701,N_845);
nor U2326 (N_2326,N_408,N_410);
nand U2327 (N_2327,N_784,N_900);
or U2328 (N_2328,N_204,N_1154);
xor U2329 (N_2329,N_1141,N_264);
and U2330 (N_2330,N_450,N_790);
nor U2331 (N_2331,N_487,N_714);
nand U2332 (N_2332,N_93,N_125);
nor U2333 (N_2333,N_610,N_764);
nor U2334 (N_2334,N_569,N_1220);
nand U2335 (N_2335,N_1111,N_13);
nand U2336 (N_2336,N_1231,N_838);
nand U2337 (N_2337,N_987,N_473);
or U2338 (N_2338,N_846,N_1053);
nand U2339 (N_2339,N_241,N_98);
or U2340 (N_2340,N_1217,N_780);
and U2341 (N_2341,N_1110,N_220);
nor U2342 (N_2342,N_410,N_948);
and U2343 (N_2343,N_576,N_872);
nor U2344 (N_2344,N_383,N_352);
nand U2345 (N_2345,N_243,N_641);
or U2346 (N_2346,N_1064,N_952);
nor U2347 (N_2347,N_936,N_450);
xnor U2348 (N_2348,N_400,N_784);
nor U2349 (N_2349,N_792,N_36);
nor U2350 (N_2350,N_592,N_264);
nand U2351 (N_2351,N_191,N_1046);
and U2352 (N_2352,N_946,N_55);
and U2353 (N_2353,N_711,N_1121);
or U2354 (N_2354,N_280,N_1152);
nand U2355 (N_2355,N_551,N_1207);
nand U2356 (N_2356,N_1141,N_639);
or U2357 (N_2357,N_457,N_1033);
nor U2358 (N_2358,N_832,N_210);
nor U2359 (N_2359,N_38,N_910);
nor U2360 (N_2360,N_11,N_259);
or U2361 (N_2361,N_105,N_501);
xnor U2362 (N_2362,N_690,N_1161);
nor U2363 (N_2363,N_706,N_819);
xnor U2364 (N_2364,N_189,N_910);
or U2365 (N_2365,N_1091,N_141);
or U2366 (N_2366,N_350,N_262);
and U2367 (N_2367,N_964,N_44);
and U2368 (N_2368,N_659,N_249);
nor U2369 (N_2369,N_404,N_1001);
and U2370 (N_2370,N_307,N_505);
nand U2371 (N_2371,N_987,N_825);
xnor U2372 (N_2372,N_951,N_1070);
and U2373 (N_2373,N_890,N_792);
or U2374 (N_2374,N_869,N_1037);
and U2375 (N_2375,N_207,N_383);
nand U2376 (N_2376,N_272,N_820);
and U2377 (N_2377,N_549,N_556);
nand U2378 (N_2378,N_247,N_637);
nor U2379 (N_2379,N_1002,N_1023);
nand U2380 (N_2380,N_1083,N_322);
or U2381 (N_2381,N_861,N_1108);
xnor U2382 (N_2382,N_230,N_312);
nand U2383 (N_2383,N_876,N_46);
nor U2384 (N_2384,N_1039,N_230);
nand U2385 (N_2385,N_864,N_389);
or U2386 (N_2386,N_1222,N_776);
or U2387 (N_2387,N_191,N_1090);
xnor U2388 (N_2388,N_195,N_994);
or U2389 (N_2389,N_443,N_955);
nand U2390 (N_2390,N_183,N_691);
nor U2391 (N_2391,N_6,N_510);
and U2392 (N_2392,N_689,N_496);
nand U2393 (N_2393,N_47,N_69);
nand U2394 (N_2394,N_610,N_238);
or U2395 (N_2395,N_1061,N_89);
nor U2396 (N_2396,N_579,N_905);
and U2397 (N_2397,N_551,N_297);
nor U2398 (N_2398,N_191,N_607);
or U2399 (N_2399,N_777,N_744);
or U2400 (N_2400,N_1146,N_442);
and U2401 (N_2401,N_677,N_984);
nand U2402 (N_2402,N_1007,N_17);
nand U2403 (N_2403,N_1028,N_191);
xnor U2404 (N_2404,N_1170,N_584);
nand U2405 (N_2405,N_711,N_114);
nor U2406 (N_2406,N_1233,N_795);
and U2407 (N_2407,N_275,N_951);
or U2408 (N_2408,N_428,N_89);
or U2409 (N_2409,N_370,N_579);
nand U2410 (N_2410,N_1231,N_481);
or U2411 (N_2411,N_282,N_454);
nor U2412 (N_2412,N_549,N_1235);
nand U2413 (N_2413,N_429,N_412);
xor U2414 (N_2414,N_416,N_64);
and U2415 (N_2415,N_1225,N_460);
nand U2416 (N_2416,N_539,N_698);
xor U2417 (N_2417,N_744,N_979);
or U2418 (N_2418,N_534,N_67);
and U2419 (N_2419,N_205,N_217);
nor U2420 (N_2420,N_395,N_676);
or U2421 (N_2421,N_678,N_1232);
and U2422 (N_2422,N_245,N_470);
nand U2423 (N_2423,N_350,N_1246);
nor U2424 (N_2424,N_604,N_1015);
or U2425 (N_2425,N_653,N_1143);
or U2426 (N_2426,N_828,N_1210);
or U2427 (N_2427,N_54,N_771);
or U2428 (N_2428,N_1160,N_1239);
and U2429 (N_2429,N_252,N_627);
nor U2430 (N_2430,N_1128,N_1104);
xor U2431 (N_2431,N_530,N_846);
nand U2432 (N_2432,N_194,N_379);
nand U2433 (N_2433,N_347,N_173);
and U2434 (N_2434,N_854,N_893);
xor U2435 (N_2435,N_518,N_489);
or U2436 (N_2436,N_1219,N_964);
xnor U2437 (N_2437,N_129,N_1190);
xnor U2438 (N_2438,N_117,N_1234);
nand U2439 (N_2439,N_578,N_297);
xor U2440 (N_2440,N_408,N_427);
and U2441 (N_2441,N_777,N_510);
nor U2442 (N_2442,N_722,N_93);
xor U2443 (N_2443,N_1125,N_1219);
or U2444 (N_2444,N_88,N_960);
nand U2445 (N_2445,N_498,N_1089);
nand U2446 (N_2446,N_805,N_577);
or U2447 (N_2447,N_221,N_54);
nand U2448 (N_2448,N_626,N_1125);
xor U2449 (N_2449,N_803,N_122);
xor U2450 (N_2450,N_910,N_1027);
nor U2451 (N_2451,N_422,N_1016);
and U2452 (N_2452,N_40,N_745);
nor U2453 (N_2453,N_36,N_1221);
and U2454 (N_2454,N_938,N_1177);
xor U2455 (N_2455,N_216,N_1050);
nand U2456 (N_2456,N_728,N_379);
nand U2457 (N_2457,N_721,N_730);
xnor U2458 (N_2458,N_896,N_623);
and U2459 (N_2459,N_141,N_428);
or U2460 (N_2460,N_255,N_503);
xnor U2461 (N_2461,N_848,N_493);
xnor U2462 (N_2462,N_868,N_134);
and U2463 (N_2463,N_663,N_1011);
nor U2464 (N_2464,N_480,N_501);
xnor U2465 (N_2465,N_735,N_371);
or U2466 (N_2466,N_466,N_688);
nand U2467 (N_2467,N_555,N_1114);
xnor U2468 (N_2468,N_121,N_579);
or U2469 (N_2469,N_445,N_28);
xnor U2470 (N_2470,N_1085,N_834);
nand U2471 (N_2471,N_730,N_1018);
or U2472 (N_2472,N_292,N_503);
and U2473 (N_2473,N_485,N_1230);
xor U2474 (N_2474,N_396,N_39);
or U2475 (N_2475,N_441,N_961);
and U2476 (N_2476,N_528,N_105);
and U2477 (N_2477,N_1035,N_478);
nand U2478 (N_2478,N_830,N_988);
and U2479 (N_2479,N_618,N_24);
xor U2480 (N_2480,N_1223,N_1123);
and U2481 (N_2481,N_375,N_432);
xnor U2482 (N_2482,N_288,N_406);
or U2483 (N_2483,N_686,N_101);
nand U2484 (N_2484,N_30,N_835);
nand U2485 (N_2485,N_696,N_967);
nand U2486 (N_2486,N_225,N_880);
and U2487 (N_2487,N_1215,N_490);
nand U2488 (N_2488,N_1233,N_840);
xnor U2489 (N_2489,N_827,N_919);
and U2490 (N_2490,N_914,N_323);
and U2491 (N_2491,N_349,N_9);
nor U2492 (N_2492,N_172,N_1087);
and U2493 (N_2493,N_382,N_749);
and U2494 (N_2494,N_846,N_801);
or U2495 (N_2495,N_972,N_814);
xnor U2496 (N_2496,N_783,N_376);
and U2497 (N_2497,N_122,N_573);
or U2498 (N_2498,N_279,N_528);
or U2499 (N_2499,N_574,N_20);
nor U2500 (N_2500,N_2017,N_1734);
xnor U2501 (N_2501,N_2161,N_2210);
nand U2502 (N_2502,N_1407,N_1963);
nand U2503 (N_2503,N_1566,N_2290);
nand U2504 (N_2504,N_1985,N_1532);
nor U2505 (N_2505,N_1468,N_1719);
or U2506 (N_2506,N_2132,N_2299);
nand U2507 (N_2507,N_1531,N_2120);
nand U2508 (N_2508,N_2312,N_1630);
or U2509 (N_2509,N_2007,N_1945);
nand U2510 (N_2510,N_1815,N_1336);
and U2511 (N_2511,N_1955,N_1415);
nand U2512 (N_2512,N_1895,N_1497);
and U2513 (N_2513,N_1387,N_2242);
nand U2514 (N_2514,N_1359,N_1943);
xor U2515 (N_2515,N_2183,N_1932);
nor U2516 (N_2516,N_2480,N_1363);
or U2517 (N_2517,N_1279,N_1297);
nand U2518 (N_2518,N_2412,N_1831);
or U2519 (N_2519,N_1644,N_1420);
xnor U2520 (N_2520,N_1461,N_1647);
and U2521 (N_2521,N_2366,N_1830);
nor U2522 (N_2522,N_1499,N_1633);
nor U2523 (N_2523,N_1349,N_1796);
or U2524 (N_2524,N_1341,N_2225);
nor U2525 (N_2525,N_2282,N_1813);
and U2526 (N_2526,N_1929,N_1556);
nand U2527 (N_2527,N_1626,N_2350);
nor U2528 (N_2528,N_1487,N_1944);
xor U2529 (N_2529,N_1718,N_2354);
and U2530 (N_2530,N_2451,N_2306);
or U2531 (N_2531,N_1896,N_2001);
xnor U2532 (N_2532,N_2437,N_2089);
xor U2533 (N_2533,N_1334,N_1933);
and U2534 (N_2534,N_2420,N_2086);
and U2535 (N_2535,N_1786,N_1738);
xnor U2536 (N_2536,N_1400,N_1260);
and U2537 (N_2537,N_2313,N_1322);
nand U2538 (N_2538,N_1370,N_2202);
nor U2539 (N_2539,N_1956,N_2296);
xor U2540 (N_2540,N_1864,N_2044);
and U2541 (N_2541,N_1386,N_2198);
and U2542 (N_2542,N_2331,N_1755);
or U2543 (N_2543,N_1635,N_2353);
nand U2544 (N_2544,N_1439,N_1263);
nor U2545 (N_2545,N_1975,N_2476);
nand U2546 (N_2546,N_2150,N_1754);
xnor U2547 (N_2547,N_1617,N_1666);
and U2548 (N_2548,N_2492,N_1654);
nand U2549 (N_2549,N_1305,N_2160);
xnor U2550 (N_2550,N_2119,N_2337);
nor U2551 (N_2551,N_2378,N_1332);
xor U2552 (N_2552,N_2240,N_2320);
and U2553 (N_2553,N_2146,N_2038);
xor U2554 (N_2554,N_1506,N_1558);
and U2555 (N_2555,N_1707,N_1920);
nand U2556 (N_2556,N_2030,N_2416);
xor U2557 (N_2557,N_1315,N_2372);
xnor U2558 (N_2558,N_1538,N_2403);
nor U2559 (N_2559,N_1458,N_1989);
or U2560 (N_2560,N_1312,N_1525);
xnor U2561 (N_2561,N_1803,N_1394);
nand U2562 (N_2562,N_1509,N_1431);
nand U2563 (N_2563,N_2167,N_1671);
nand U2564 (N_2564,N_2301,N_2228);
xor U2565 (N_2565,N_1588,N_1587);
nand U2566 (N_2566,N_1980,N_1595);
nand U2567 (N_2567,N_1730,N_1395);
or U2568 (N_2568,N_1379,N_1836);
and U2569 (N_2569,N_2303,N_2112);
nor U2570 (N_2570,N_2346,N_2367);
and U2571 (N_2571,N_1899,N_1521);
and U2572 (N_2572,N_2274,N_1947);
xnor U2573 (N_2573,N_2383,N_1294);
nor U2574 (N_2574,N_1560,N_2386);
xor U2575 (N_2575,N_1578,N_1976);
and U2576 (N_2576,N_2364,N_1612);
nand U2577 (N_2577,N_2052,N_1576);
xnor U2578 (N_2578,N_1575,N_2011);
nor U2579 (N_2579,N_1902,N_1492);
nand U2580 (N_2580,N_2307,N_1690);
nand U2581 (N_2581,N_2490,N_2427);
nor U2582 (N_2582,N_1256,N_2070);
nor U2583 (N_2583,N_2211,N_2236);
nor U2584 (N_2584,N_1467,N_2063);
nor U2585 (N_2585,N_1358,N_2128);
xnor U2586 (N_2586,N_2100,N_1473);
nor U2587 (N_2587,N_1314,N_1463);
nand U2588 (N_2588,N_2181,N_2401);
or U2589 (N_2589,N_1516,N_1378);
nor U2590 (N_2590,N_1990,N_2201);
xor U2591 (N_2591,N_2477,N_1539);
xnor U2592 (N_2592,N_2148,N_2145);
or U2593 (N_2593,N_2158,N_2238);
and U2594 (N_2594,N_2288,N_1562);
nand U2595 (N_2595,N_1392,N_2334);
or U2596 (N_2596,N_1591,N_2064);
xor U2597 (N_2597,N_2104,N_1605);
nand U2598 (N_2598,N_2097,N_2159);
or U2599 (N_2599,N_2212,N_1554);
or U2600 (N_2600,N_1888,N_1632);
nand U2601 (N_2601,N_1892,N_1816);
or U2602 (N_2602,N_1807,N_1780);
nor U2603 (N_2603,N_1916,N_2003);
xor U2604 (N_2604,N_1958,N_2096);
nor U2605 (N_2605,N_2072,N_1446);
nand U2606 (N_2606,N_1478,N_1289);
and U2607 (N_2607,N_1475,N_1393);
and U2608 (N_2608,N_1965,N_1277);
and U2609 (N_2609,N_1999,N_1427);
nand U2610 (N_2610,N_2495,N_1657);
or U2611 (N_2611,N_1858,N_2464);
and U2612 (N_2612,N_1802,N_1700);
or U2613 (N_2613,N_1327,N_2435);
xnor U2614 (N_2614,N_1917,N_2314);
nor U2615 (N_2615,N_1482,N_2116);
nor U2616 (N_2616,N_1979,N_1897);
nor U2617 (N_2617,N_1447,N_1798);
and U2618 (N_2618,N_2419,N_1889);
xnor U2619 (N_2619,N_1418,N_1847);
and U2620 (N_2620,N_1883,N_1424);
and U2621 (N_2621,N_1275,N_1953);
or U2622 (N_2622,N_1867,N_1855);
nor U2623 (N_2623,N_2027,N_1469);
nor U2624 (N_2624,N_2342,N_2393);
nor U2625 (N_2625,N_1293,N_2259);
and U2626 (N_2626,N_2074,N_2231);
nor U2627 (N_2627,N_2448,N_2170);
nor U2628 (N_2628,N_1949,N_2139);
xnor U2629 (N_2629,N_1749,N_2115);
nand U2630 (N_2630,N_2178,N_1586);
xor U2631 (N_2631,N_1561,N_2041);
nand U2632 (N_2632,N_1390,N_1269);
or U2633 (N_2633,N_1715,N_2287);
nand U2634 (N_2634,N_1419,N_1503);
and U2635 (N_2635,N_1744,N_2180);
or U2636 (N_2636,N_1930,N_1601);
xnor U2637 (N_2637,N_1573,N_2388);
nor U2638 (N_2638,N_1951,N_2262);
nor U2639 (N_2639,N_1887,N_1721);
nand U2640 (N_2640,N_2234,N_2226);
xor U2641 (N_2641,N_2018,N_2237);
and U2642 (N_2642,N_2136,N_2363);
or U2643 (N_2643,N_2034,N_1907);
and U2644 (N_2644,N_1423,N_2162);
or U2645 (N_2645,N_2200,N_2157);
nor U2646 (N_2646,N_2468,N_1880);
or U2647 (N_2647,N_1437,N_1849);
nor U2648 (N_2648,N_1912,N_1267);
and U2649 (N_2649,N_2394,N_2058);
nor U2650 (N_2650,N_1522,N_2143);
or U2651 (N_2651,N_2075,N_1675);
nand U2652 (N_2652,N_1316,N_1321);
xor U2653 (N_2653,N_1670,N_1607);
nor U2654 (N_2654,N_2369,N_1430);
xnor U2655 (N_2655,N_2449,N_1662);
nand U2656 (N_2656,N_1510,N_1723);
xor U2657 (N_2657,N_2377,N_2293);
and U2658 (N_2658,N_1585,N_1898);
or U2659 (N_2659,N_2281,N_1594);
and U2660 (N_2660,N_1391,N_2359);
nor U2661 (N_2661,N_1760,N_1524);
nor U2662 (N_2662,N_2121,N_2032);
nor U2663 (N_2663,N_1608,N_1704);
nand U2664 (N_2664,N_2418,N_1567);
or U2665 (N_2665,N_2182,N_2429);
xor U2666 (N_2666,N_2219,N_1735);
and U2667 (N_2667,N_1822,N_2279);
nand U2668 (N_2668,N_1967,N_1517);
or U2669 (N_2669,N_1346,N_1329);
nand U2670 (N_2670,N_1384,N_1716);
xor U2671 (N_2671,N_1500,N_1784);
and U2672 (N_2672,N_2229,N_2475);
or U2673 (N_2673,N_1637,N_1402);
xor U2674 (N_2674,N_1770,N_2043);
and U2675 (N_2675,N_1481,N_1834);
and U2676 (N_2676,N_2375,N_1992);
or U2677 (N_2677,N_2414,N_2322);
and U2678 (N_2678,N_2406,N_1863);
or U2679 (N_2679,N_2076,N_1298);
or U2680 (N_2680,N_1540,N_2494);
xor U2681 (N_2681,N_1776,N_2409);
nor U2682 (N_2682,N_1493,N_1536);
nand U2683 (N_2683,N_1927,N_1713);
or U2684 (N_2684,N_2190,N_1441);
nor U2685 (N_2685,N_2214,N_1766);
and U2686 (N_2686,N_2209,N_1812);
nor U2687 (N_2687,N_1619,N_1331);
xor U2688 (N_2688,N_2188,N_2381);
xnor U2689 (N_2689,N_1788,N_2048);
and U2690 (N_2690,N_1753,N_1765);
nor U2691 (N_2691,N_1310,N_2250);
nand U2692 (N_2692,N_1655,N_2125);
or U2693 (N_2693,N_2166,N_2151);
nor U2694 (N_2694,N_1380,N_1382);
xor U2695 (N_2695,N_2263,N_1860);
or U2696 (N_2696,N_1518,N_2141);
nor U2697 (N_2697,N_1258,N_2439);
and U2698 (N_2698,N_2223,N_2498);
nor U2699 (N_2699,N_1679,N_1599);
xor U2700 (N_2700,N_2488,N_2149);
nand U2701 (N_2701,N_2261,N_1904);
nand U2702 (N_2702,N_2071,N_2248);
and U2703 (N_2703,N_1443,N_2297);
and U2704 (N_2704,N_1593,N_2402);
or U2705 (N_2705,N_1253,N_1708);
or U2706 (N_2706,N_2020,N_2272);
nand U2707 (N_2707,N_2473,N_1792);
nor U2708 (N_2708,N_2187,N_1981);
and U2709 (N_2709,N_1729,N_2257);
or U2710 (N_2710,N_2298,N_2118);
nor U2711 (N_2711,N_1737,N_1577);
nand U2712 (N_2712,N_1598,N_1620);
nor U2713 (N_2713,N_1941,N_1782);
and U2714 (N_2714,N_1757,N_2305);
xor U2715 (N_2715,N_2332,N_1429);
xnor U2716 (N_2716,N_1820,N_1262);
xor U2717 (N_2717,N_1832,N_2054);
or U2718 (N_2718,N_1922,N_2442);
and U2719 (N_2719,N_1411,N_2487);
or U2720 (N_2720,N_2105,N_1891);
and U2721 (N_2721,N_1672,N_1703);
xor U2722 (N_2722,N_1374,N_2436);
xor U2723 (N_2723,N_1628,N_1271);
xnor U2724 (N_2724,N_2036,N_1938);
or U2725 (N_2725,N_1991,N_2454);
xor U2726 (N_2726,N_1848,N_1507);
or U2727 (N_2727,N_1701,N_2028);
and U2728 (N_2728,N_1465,N_1270);
nor U2729 (N_2729,N_2450,N_2341);
nand U2730 (N_2730,N_1604,N_1692);
xor U2731 (N_2731,N_2164,N_1736);
xor U2732 (N_2732,N_1972,N_2068);
or U2733 (N_2733,N_1344,N_2351);
or U2734 (N_2734,N_2222,N_1348);
nand U2735 (N_2735,N_1772,N_1661);
and U2736 (N_2736,N_1324,N_1552);
or U2737 (N_2737,N_2380,N_2042);
nand U2738 (N_2738,N_2343,N_1557);
or U2739 (N_2739,N_2285,N_1885);
nand U2740 (N_2740,N_1789,N_1569);
and U2741 (N_2741,N_2224,N_1347);
nand U2742 (N_2742,N_2333,N_1853);
and U2743 (N_2743,N_1290,N_2280);
or U2744 (N_2744,N_1523,N_1438);
xnor U2745 (N_2745,N_2066,N_2186);
xor U2746 (N_2746,N_1320,N_1828);
nor U2747 (N_2747,N_1921,N_2194);
or U2748 (N_2748,N_2452,N_1457);
and U2749 (N_2749,N_2047,N_2005);
or U2750 (N_2750,N_2455,N_1574);
nand U2751 (N_2751,N_2284,N_1629);
and U2752 (N_2752,N_2103,N_2156);
xnor U2753 (N_2753,N_2138,N_1937);
xor U2754 (N_2754,N_1988,N_1319);
and U2755 (N_2755,N_1352,N_2445);
and U2756 (N_2756,N_1696,N_2065);
nand U2757 (N_2757,N_1292,N_1873);
or U2758 (N_2758,N_1611,N_1652);
nand U2759 (N_2759,N_2217,N_1440);
and U2760 (N_2760,N_1971,N_2362);
nor U2761 (N_2761,N_1372,N_1846);
and U2762 (N_2762,N_1309,N_1551);
nand U2763 (N_2763,N_2407,N_1442);
and U2764 (N_2764,N_1251,N_1445);
and U2765 (N_2765,N_1706,N_2056);
nand U2766 (N_2766,N_1412,N_1903);
nor U2767 (N_2767,N_1535,N_2241);
nor U2768 (N_2768,N_1449,N_1702);
xor U2769 (N_2769,N_2046,N_1859);
nor U2770 (N_2770,N_1714,N_2215);
xnor U2771 (N_2771,N_1997,N_1781);
xnor U2772 (N_2772,N_1642,N_1810);
xor U2773 (N_2773,N_1356,N_1383);
xnor U2774 (N_2774,N_1422,N_1919);
nor U2775 (N_2775,N_1682,N_1732);
xnor U2776 (N_2776,N_2277,N_2268);
nand U2777 (N_2777,N_2176,N_1417);
or U2778 (N_2778,N_1805,N_2049);
nor U2779 (N_2779,N_2447,N_2078);
nor U2780 (N_2780,N_2286,N_2338);
nand U2781 (N_2781,N_1600,N_1814);
xnor U2782 (N_2782,N_1528,N_2318);
nor U2783 (N_2783,N_1763,N_1908);
xnor U2784 (N_2784,N_1693,N_2428);
nor U2785 (N_2785,N_1264,N_1301);
xor U2786 (N_2786,N_2483,N_1544);
xor U2787 (N_2787,N_1345,N_1491);
and U2788 (N_2788,N_1866,N_1350);
xor U2789 (N_2789,N_1366,N_2400);
and U2790 (N_2790,N_1527,N_1425);
nand U2791 (N_2791,N_1257,N_2039);
nor U2792 (N_2792,N_2317,N_1857);
or U2793 (N_2793,N_1874,N_1748);
xor U2794 (N_2794,N_1893,N_2023);
nor U2795 (N_2795,N_1308,N_1502);
or U2796 (N_2796,N_1845,N_1373);
nand U2797 (N_2797,N_2300,N_1284);
or U2798 (N_2798,N_1288,N_2191);
and U2799 (N_2799,N_1926,N_1399);
and U2800 (N_2800,N_1658,N_2422);
and U2801 (N_2801,N_2360,N_2197);
xnor U2802 (N_2802,N_1960,N_1759);
xnor U2803 (N_2803,N_2084,N_1689);
nand U2804 (N_2804,N_1747,N_2291);
nand U2805 (N_2805,N_2459,N_2395);
nor U2806 (N_2806,N_2127,N_1984);
nand U2807 (N_2807,N_2079,N_2432);
nor U2808 (N_2808,N_2472,N_1854);
nand U2809 (N_2809,N_2385,N_1389);
or U2810 (N_2810,N_1793,N_1526);
or U2811 (N_2811,N_2059,N_1335);
nor U2812 (N_2812,N_1592,N_2329);
xnor U2813 (N_2813,N_2361,N_1767);
nand U2814 (N_2814,N_2462,N_1490);
xnor U2815 (N_2815,N_1621,N_1444);
or U2816 (N_2816,N_1645,N_1838);
nand U2817 (N_2817,N_1882,N_1259);
nor U2818 (N_2818,N_2232,N_2324);
nor U2819 (N_2819,N_1973,N_1750);
xor U2820 (N_2820,N_1910,N_2499);
nor U2821 (N_2821,N_2405,N_1978);
and U2822 (N_2822,N_1787,N_1278);
nor U2823 (N_2823,N_1683,N_1280);
and U2824 (N_2824,N_1504,N_1638);
and U2825 (N_2825,N_1993,N_2153);
nor U2826 (N_2826,N_1306,N_2463);
and U2827 (N_2827,N_2008,N_2133);
xor U2828 (N_2828,N_1827,N_1687);
or U2829 (N_2829,N_2208,N_2321);
nor U2830 (N_2830,N_2294,N_1362);
or U2831 (N_2831,N_1841,N_2340);
nand U2832 (N_2832,N_1911,N_2255);
nor U2833 (N_2833,N_2345,N_1549);
and U2834 (N_2834,N_2423,N_1553);
and U2835 (N_2835,N_2175,N_1901);
xnor U2836 (N_2836,N_1641,N_2376);
xor U2837 (N_2837,N_1695,N_1783);
and U2838 (N_2838,N_1634,N_2374);
nand U2839 (N_2839,N_1741,N_1285);
nand U2840 (N_2840,N_1817,N_2037);
nand U2841 (N_2841,N_1940,N_1886);
nor U2842 (N_2842,N_1686,N_2328);
and U2843 (N_2843,N_2022,N_1307);
and U2844 (N_2844,N_1291,N_1618);
and U2845 (N_2845,N_1584,N_1564);
or U2846 (N_2846,N_2264,N_1785);
xor U2847 (N_2847,N_1808,N_1339);
or U2848 (N_2848,N_2135,N_1505);
or U2849 (N_2849,N_1954,N_2252);
xnor U2850 (N_2850,N_2040,N_1819);
or U2851 (N_2851,N_2355,N_2457);
or U2852 (N_2852,N_2016,N_2051);
nor U2853 (N_2853,N_1323,N_2174);
nand U2854 (N_2854,N_1751,N_1795);
and U2855 (N_2855,N_1453,N_1764);
xnor U2856 (N_2856,N_1923,N_2387);
xnor U2857 (N_2857,N_1746,N_2357);
nand U2858 (N_2858,N_2276,N_2273);
or U2859 (N_2859,N_1571,N_2478);
nand U2860 (N_2860,N_1381,N_1818);
nand U2861 (N_2861,N_1408,N_1663);
xnor U2862 (N_2862,N_1833,N_2216);
or U2863 (N_2863,N_2370,N_1649);
or U2864 (N_2864,N_2077,N_1733);
and U2865 (N_2865,N_2292,N_2247);
nor U2866 (N_2866,N_2244,N_1724);
xnor U2867 (N_2867,N_1840,N_2249);
or U2868 (N_2868,N_2129,N_2055);
and U2869 (N_2869,N_1881,N_1337);
nand U2870 (N_2870,N_1711,N_1274);
nor U2871 (N_2871,N_1851,N_1451);
and U2872 (N_2872,N_1842,N_2243);
nand U2873 (N_2873,N_2443,N_1712);
nor U2874 (N_2874,N_1579,N_1537);
nand U2875 (N_2875,N_1868,N_1799);
or U2876 (N_2876,N_1403,N_2140);
or U2877 (N_2877,N_2196,N_2348);
xnor U2878 (N_2878,N_2399,N_1416);
xor U2879 (N_2879,N_2122,N_2061);
or U2880 (N_2880,N_1821,N_1801);
and U2881 (N_2881,N_1761,N_2397);
xor U2882 (N_2882,N_1313,N_2347);
nor U2883 (N_2883,N_1287,N_1962);
or U2884 (N_2884,N_2456,N_2114);
or U2885 (N_2885,N_1928,N_1625);
or U2886 (N_2886,N_2053,N_1806);
nand U2887 (N_2887,N_2080,N_2304);
nor U2888 (N_2888,N_2382,N_1961);
xor U2889 (N_2889,N_2009,N_2349);
nor U2890 (N_2890,N_2458,N_2339);
and U2891 (N_2891,N_2021,N_1627);
xor U2892 (N_2892,N_1368,N_2431);
nor U2893 (N_2893,N_1771,N_2426);
or U2894 (N_2894,N_2206,N_2497);
and U2895 (N_2895,N_1325,N_2109);
or U2896 (N_2896,N_1508,N_2352);
nand U2897 (N_2897,N_1470,N_1850);
xor U2898 (N_2898,N_1534,N_2254);
nand U2899 (N_2899,N_2470,N_2316);
nor U2900 (N_2900,N_2134,N_1778);
or U2901 (N_2901,N_1565,N_2467);
xor U2902 (N_2902,N_2466,N_1823);
nor U2903 (N_2903,N_1317,N_1603);
xor U2904 (N_2904,N_1303,N_2315);
xnor U2905 (N_2905,N_1583,N_1773);
nand U2906 (N_2906,N_2433,N_1681);
nand U2907 (N_2907,N_1791,N_1631);
xor U2908 (N_2908,N_2270,N_1436);
or U2909 (N_2909,N_1871,N_1360);
nor U2910 (N_2910,N_1677,N_2368);
nand U2911 (N_2911,N_1698,N_1915);
or U2912 (N_2912,N_2269,N_1742);
or U2913 (N_2913,N_1466,N_2087);
xnor U2914 (N_2914,N_1472,N_1354);
nand U2915 (N_2915,N_2227,N_1296);
or U2916 (N_2916,N_1498,N_2025);
and U2917 (N_2917,N_1974,N_1343);
and U2918 (N_2918,N_1283,N_1530);
xor U2919 (N_2919,N_1648,N_1435);
nor U2920 (N_2920,N_1533,N_2496);
nor U2921 (N_2921,N_1454,N_2192);
nand U2922 (N_2922,N_1281,N_1340);
nand U2923 (N_2923,N_2108,N_1685);
nor U2924 (N_2924,N_2373,N_1676);
nor U2925 (N_2925,N_1636,N_2163);
xnor U2926 (N_2926,N_1501,N_1456);
or U2927 (N_2927,N_1865,N_2311);
and U2928 (N_2928,N_1769,N_1639);
or U2929 (N_2929,N_1462,N_1512);
nand U2930 (N_2930,N_2471,N_1694);
nor U2931 (N_2931,N_2171,N_1646);
xnor U2932 (N_2932,N_2092,N_1450);
xor U2933 (N_2933,N_1779,N_1998);
nor U2934 (N_2934,N_2205,N_1936);
nor U2935 (N_2935,N_2266,N_2195);
nand U2936 (N_2936,N_1946,N_1656);
nand U2937 (N_2937,N_1286,N_1545);
nor U2938 (N_2938,N_1884,N_1924);
xor U2939 (N_2939,N_2033,N_1826);
xor U2940 (N_2940,N_1514,N_1688);
and U2941 (N_2941,N_2213,N_2189);
nor U2942 (N_2942,N_1909,N_1367);
xor U2943 (N_2943,N_2168,N_2410);
nor U2944 (N_2944,N_2002,N_2265);
or U2945 (N_2945,N_2081,N_1768);
nor U2946 (N_2946,N_2278,N_1837);
nor U2947 (N_2947,N_1326,N_1311);
nor U2948 (N_2948,N_1756,N_1318);
and U2949 (N_2949,N_2204,N_2062);
or U2950 (N_2950,N_2123,N_1875);
xor U2951 (N_2951,N_1397,N_1674);
and U2952 (N_2952,N_1797,N_2358);
nor U2953 (N_2953,N_2094,N_1330);
or U2954 (N_2954,N_1844,N_1484);
xnor U2955 (N_2955,N_1968,N_2221);
and U2956 (N_2956,N_1494,N_1935);
nand U2957 (N_2957,N_2404,N_2179);
xor U2958 (N_2958,N_2106,N_2110);
or U2959 (N_2959,N_2199,N_1252);
or U2960 (N_2960,N_1485,N_2099);
nor U2961 (N_2961,N_2283,N_1809);
or U2962 (N_2962,N_2117,N_2260);
nand U2963 (N_2963,N_1572,N_2067);
or U2964 (N_2964,N_2111,N_1404);
nor U2965 (N_2965,N_2060,N_1869);
xor U2966 (N_2966,N_2126,N_1550);
nor U2967 (N_2967,N_1861,N_2319);
and U2968 (N_2968,N_2245,N_1464);
xor U2969 (N_2969,N_2218,N_1273);
or U2970 (N_2970,N_1614,N_2327);
xor U2971 (N_2971,N_1775,N_1459);
xor U2972 (N_2972,N_1942,N_1268);
and U2973 (N_2973,N_1299,N_1890);
nand U2974 (N_2974,N_1710,N_1665);
nand U2975 (N_2975,N_2230,N_1650);
nor U2976 (N_2976,N_2091,N_1667);
nor U2977 (N_2977,N_2408,N_2050);
nand U2978 (N_2978,N_1913,N_1987);
nand U2979 (N_2979,N_1905,N_1622);
or U2980 (N_2980,N_2107,N_1364);
and U2981 (N_2981,N_2469,N_1396);
nand U2982 (N_2982,N_1255,N_1669);
xnor U2983 (N_2983,N_1762,N_1406);
nor U2984 (N_2984,N_1964,N_2251);
and U2985 (N_2985,N_2485,N_1640);
or U2986 (N_2986,N_2093,N_2295);
or U2987 (N_2987,N_1388,N_1409);
xnor U2988 (N_2988,N_2391,N_2203);
xnor U2989 (N_2989,N_1800,N_1410);
or U2990 (N_2990,N_2323,N_2131);
nor U2991 (N_2991,N_2130,N_1982);
nor U2992 (N_2992,N_1477,N_1659);
or U2993 (N_2993,N_2491,N_1699);
nand U2994 (N_2994,N_1250,N_2102);
xnor U2995 (N_2995,N_1966,N_1835);
or U2996 (N_2996,N_1957,N_2172);
and U2997 (N_2997,N_1486,N_2253);
and U2998 (N_2998,N_1948,N_2256);
xnor U2999 (N_2999,N_2460,N_1474);
and U3000 (N_3000,N_1731,N_2124);
or U3001 (N_3001,N_1720,N_1994);
xnor U3002 (N_3002,N_1697,N_1254);
xnor U3003 (N_3003,N_1265,N_2177);
nand U3004 (N_3004,N_2101,N_2024);
and U3005 (N_3005,N_1375,N_2029);
or U3006 (N_3006,N_1931,N_1589);
or U3007 (N_3007,N_2233,N_1745);
nand U3008 (N_3008,N_1266,N_2098);
nand U3009 (N_3009,N_1684,N_1488);
nor U3010 (N_3010,N_1369,N_1548);
and U3011 (N_3011,N_1328,N_1597);
and U3012 (N_3012,N_2239,N_2258);
nor U3013 (N_3013,N_1624,N_2390);
xor U3014 (N_3014,N_2275,N_1261);
nand U3015 (N_3015,N_2235,N_2085);
xnor U3016 (N_3016,N_1879,N_1555);
and U3017 (N_3017,N_1804,N_1602);
and U3018 (N_3018,N_1609,N_1398);
nor U3019 (N_3019,N_2424,N_2169);
nand U3020 (N_3020,N_2095,N_1479);
and U3021 (N_3021,N_2438,N_1727);
and U3022 (N_3022,N_1483,N_2010);
xnor U3023 (N_3023,N_1623,N_1722);
or U3024 (N_3024,N_1547,N_1872);
xor U3025 (N_3025,N_1570,N_1758);
xnor U3026 (N_3026,N_2484,N_1705);
and U3027 (N_3027,N_2310,N_2326);
nor U3028 (N_3028,N_2035,N_1680);
xor U3029 (N_3029,N_1489,N_2246);
xor U3030 (N_3030,N_2271,N_1743);
and U3031 (N_3031,N_1914,N_1426);
and U3032 (N_3032,N_2482,N_1668);
nor U3033 (N_3033,N_1900,N_2302);
and U3034 (N_3034,N_1673,N_2365);
nor U3035 (N_3035,N_1546,N_1433);
or U3036 (N_3036,N_2481,N_1434);
xor U3037 (N_3037,N_1272,N_1333);
or U3038 (N_3038,N_1471,N_1351);
nand U3039 (N_3039,N_2015,N_1582);
xor U3040 (N_3040,N_2031,N_1774);
xnor U3041 (N_3041,N_2461,N_1728);
and U3042 (N_3042,N_2486,N_1581);
nor U3043 (N_3043,N_2113,N_1342);
and U3044 (N_3044,N_1495,N_1939);
nand U3045 (N_3045,N_1460,N_2384);
nor U3046 (N_3046,N_2014,N_2413);
nand U3047 (N_3047,N_2434,N_1413);
or U3048 (N_3048,N_1996,N_1829);
and U3049 (N_3049,N_2207,N_1643);
xnor U3050 (N_3050,N_1543,N_1925);
nor U3051 (N_3051,N_2069,N_1452);
and U3052 (N_3052,N_2088,N_1876);
and U3053 (N_3053,N_1357,N_2082);
nand U3054 (N_3054,N_1476,N_2417);
xor U3055 (N_3055,N_1519,N_2440);
or U3056 (N_3056,N_2444,N_2019);
or U3057 (N_3057,N_1455,N_2430);
and U3058 (N_3058,N_1338,N_1295);
nor U3059 (N_3059,N_2344,N_1983);
and U3060 (N_3060,N_2453,N_1302);
xnor U3061 (N_3061,N_1590,N_2441);
or U3062 (N_3062,N_2013,N_2155);
nand U3063 (N_3063,N_2083,N_2446);
nand U3064 (N_3064,N_2396,N_1365);
nand U3065 (N_3065,N_2185,N_1709);
and U3066 (N_3066,N_2411,N_2308);
nand U3067 (N_3067,N_1353,N_2371);
or U3068 (N_3068,N_1513,N_2389);
nand U3069 (N_3069,N_2026,N_1870);
nor U3070 (N_3070,N_2220,N_2073);
and U3071 (N_3071,N_1995,N_1480);
or U3072 (N_3072,N_2090,N_1934);
and U3073 (N_3073,N_1520,N_1496);
nor U3074 (N_3074,N_2336,N_1421);
and U3075 (N_3075,N_1276,N_2465);
xor U3076 (N_3076,N_1664,N_1660);
xor U3077 (N_3077,N_1856,N_2325);
nor U3078 (N_3078,N_1653,N_2045);
nor U3079 (N_3079,N_2415,N_1511);
nor U3080 (N_3080,N_1790,N_1613);
xnor U3081 (N_3081,N_2398,N_2012);
nor U3082 (N_3082,N_1878,N_1825);
nand U3083 (N_3083,N_1950,N_1739);
nor U3084 (N_3084,N_2137,N_1282);
or U3085 (N_3085,N_2154,N_1559);
nor U3086 (N_3086,N_1852,N_1824);
nor U3087 (N_3087,N_1371,N_2335);
nor U3088 (N_3088,N_1777,N_1969);
and U3089 (N_3089,N_2193,N_1952);
and U3090 (N_3090,N_1616,N_2289);
xor U3091 (N_3091,N_1678,N_2489);
xor U3092 (N_3092,N_2165,N_1894);
nor U3093 (N_3093,N_2142,N_1906);
and U3094 (N_3094,N_1839,N_1300);
and U3095 (N_3095,N_1568,N_1615);
and U3096 (N_3096,N_1606,N_2184);
nor U3097 (N_3097,N_1959,N_1432);
or U3098 (N_3098,N_1918,N_2425);
nand U3099 (N_3099,N_2152,N_2006);
and U3100 (N_3100,N_1405,N_1752);
and U3101 (N_3101,N_2144,N_1448);
and U3102 (N_3102,N_1877,N_1304);
nor U3103 (N_3103,N_1414,N_1542);
or U3104 (N_3104,N_1811,N_2421);
and U3105 (N_3105,N_1376,N_1377);
nand U3106 (N_3106,N_2392,N_1725);
xnor U3107 (N_3107,N_1717,N_2004);
and U3108 (N_3108,N_2057,N_1977);
nand U3109 (N_3109,N_1610,N_1361);
xor U3110 (N_3110,N_2000,N_2493);
nor U3111 (N_3111,N_2309,N_1794);
xnor U3112 (N_3112,N_2147,N_1691);
nor U3113 (N_3113,N_1651,N_1970);
nor U3114 (N_3114,N_1843,N_2173);
or U3115 (N_3115,N_1580,N_1385);
and U3116 (N_3116,N_1355,N_2479);
nand U3117 (N_3117,N_1563,N_1862);
and U3118 (N_3118,N_2330,N_1726);
or U3119 (N_3119,N_1515,N_1428);
xnor U3120 (N_3120,N_2379,N_1596);
or U3121 (N_3121,N_1541,N_2267);
nand U3122 (N_3122,N_1529,N_1986);
nand U3123 (N_3123,N_1401,N_1740);
nand U3124 (N_3124,N_2474,N_2356);
nor U3125 (N_3125,N_1284,N_2303);
nor U3126 (N_3126,N_1735,N_2047);
or U3127 (N_3127,N_2265,N_1757);
or U3128 (N_3128,N_2215,N_1730);
and U3129 (N_3129,N_1309,N_2293);
or U3130 (N_3130,N_2186,N_1784);
and U3131 (N_3131,N_2156,N_1304);
nand U3132 (N_3132,N_2417,N_1807);
nor U3133 (N_3133,N_1470,N_1809);
nand U3134 (N_3134,N_2400,N_1780);
nor U3135 (N_3135,N_1317,N_1753);
nor U3136 (N_3136,N_1304,N_1965);
nand U3137 (N_3137,N_2281,N_1277);
nand U3138 (N_3138,N_2348,N_1473);
or U3139 (N_3139,N_1760,N_1640);
nand U3140 (N_3140,N_1267,N_1266);
nor U3141 (N_3141,N_1294,N_1532);
and U3142 (N_3142,N_1930,N_1337);
and U3143 (N_3143,N_2103,N_1807);
nor U3144 (N_3144,N_1463,N_1299);
nand U3145 (N_3145,N_1643,N_1357);
nor U3146 (N_3146,N_2088,N_1672);
nor U3147 (N_3147,N_1861,N_2240);
and U3148 (N_3148,N_2475,N_1606);
xor U3149 (N_3149,N_1319,N_2107);
nand U3150 (N_3150,N_1675,N_2310);
nand U3151 (N_3151,N_1671,N_2093);
or U3152 (N_3152,N_2330,N_1716);
or U3153 (N_3153,N_2498,N_2284);
nor U3154 (N_3154,N_2357,N_2014);
nor U3155 (N_3155,N_2245,N_1768);
xnor U3156 (N_3156,N_2446,N_1270);
nand U3157 (N_3157,N_2436,N_1447);
and U3158 (N_3158,N_2220,N_2122);
nor U3159 (N_3159,N_2459,N_1499);
or U3160 (N_3160,N_2215,N_2199);
or U3161 (N_3161,N_1325,N_1377);
or U3162 (N_3162,N_1884,N_1728);
and U3163 (N_3163,N_2380,N_2354);
xor U3164 (N_3164,N_1978,N_1992);
or U3165 (N_3165,N_2439,N_2231);
and U3166 (N_3166,N_1803,N_2021);
nor U3167 (N_3167,N_2049,N_1992);
nand U3168 (N_3168,N_1441,N_2005);
xor U3169 (N_3169,N_2294,N_2317);
nor U3170 (N_3170,N_1510,N_1854);
xor U3171 (N_3171,N_1646,N_2378);
nand U3172 (N_3172,N_2179,N_1386);
xor U3173 (N_3173,N_1743,N_1906);
and U3174 (N_3174,N_1886,N_1313);
or U3175 (N_3175,N_1665,N_1528);
and U3176 (N_3176,N_1470,N_1927);
nand U3177 (N_3177,N_1945,N_1857);
xnor U3178 (N_3178,N_1809,N_2173);
and U3179 (N_3179,N_2150,N_2021);
xor U3180 (N_3180,N_2481,N_1494);
or U3181 (N_3181,N_1570,N_2102);
and U3182 (N_3182,N_1354,N_1646);
nand U3183 (N_3183,N_1990,N_1813);
xnor U3184 (N_3184,N_2394,N_1277);
nor U3185 (N_3185,N_2202,N_1748);
and U3186 (N_3186,N_2314,N_2035);
nand U3187 (N_3187,N_2211,N_1860);
nor U3188 (N_3188,N_1541,N_2333);
xor U3189 (N_3189,N_1384,N_2116);
xnor U3190 (N_3190,N_1273,N_1731);
and U3191 (N_3191,N_2498,N_2461);
and U3192 (N_3192,N_1251,N_1463);
or U3193 (N_3193,N_2453,N_1276);
nand U3194 (N_3194,N_1920,N_1691);
xor U3195 (N_3195,N_1965,N_2471);
xnor U3196 (N_3196,N_1887,N_1251);
xor U3197 (N_3197,N_1665,N_2074);
nand U3198 (N_3198,N_1994,N_1703);
nor U3199 (N_3199,N_1658,N_1670);
xnor U3200 (N_3200,N_1399,N_2110);
nand U3201 (N_3201,N_1965,N_1901);
nor U3202 (N_3202,N_1949,N_2244);
or U3203 (N_3203,N_1373,N_2183);
nor U3204 (N_3204,N_1872,N_1943);
nor U3205 (N_3205,N_1260,N_1407);
nor U3206 (N_3206,N_1643,N_1499);
nand U3207 (N_3207,N_1350,N_2166);
nand U3208 (N_3208,N_2039,N_2136);
xor U3209 (N_3209,N_1577,N_1931);
xor U3210 (N_3210,N_1370,N_1550);
nand U3211 (N_3211,N_1364,N_1919);
nand U3212 (N_3212,N_2358,N_2031);
or U3213 (N_3213,N_2287,N_2492);
nand U3214 (N_3214,N_2037,N_2429);
or U3215 (N_3215,N_2413,N_1699);
and U3216 (N_3216,N_1994,N_2462);
nand U3217 (N_3217,N_1589,N_2116);
or U3218 (N_3218,N_2322,N_2155);
xnor U3219 (N_3219,N_1704,N_1528);
and U3220 (N_3220,N_2088,N_2428);
xnor U3221 (N_3221,N_1730,N_1770);
and U3222 (N_3222,N_1520,N_2205);
or U3223 (N_3223,N_2354,N_2253);
nand U3224 (N_3224,N_1603,N_1737);
xor U3225 (N_3225,N_1859,N_2298);
and U3226 (N_3226,N_2211,N_1775);
and U3227 (N_3227,N_1527,N_2134);
xnor U3228 (N_3228,N_2051,N_1258);
nor U3229 (N_3229,N_1782,N_1666);
nand U3230 (N_3230,N_2449,N_1340);
nand U3231 (N_3231,N_1483,N_1662);
xnor U3232 (N_3232,N_2468,N_2360);
nor U3233 (N_3233,N_1377,N_2349);
nor U3234 (N_3234,N_2113,N_1422);
nand U3235 (N_3235,N_1515,N_1722);
nand U3236 (N_3236,N_2435,N_2141);
or U3237 (N_3237,N_1640,N_2326);
or U3238 (N_3238,N_1499,N_2227);
nand U3239 (N_3239,N_1934,N_2237);
nor U3240 (N_3240,N_2152,N_2074);
nand U3241 (N_3241,N_2482,N_1716);
nor U3242 (N_3242,N_1886,N_2269);
nand U3243 (N_3243,N_1913,N_1574);
nand U3244 (N_3244,N_2016,N_1510);
and U3245 (N_3245,N_2187,N_2164);
nor U3246 (N_3246,N_1692,N_1789);
nand U3247 (N_3247,N_1723,N_2467);
xor U3248 (N_3248,N_1887,N_1419);
nor U3249 (N_3249,N_2252,N_1931);
and U3250 (N_3250,N_1565,N_1752);
nand U3251 (N_3251,N_2496,N_1979);
xnor U3252 (N_3252,N_1462,N_2194);
and U3253 (N_3253,N_1568,N_2492);
or U3254 (N_3254,N_1809,N_1317);
nand U3255 (N_3255,N_2059,N_2090);
and U3256 (N_3256,N_1391,N_1729);
or U3257 (N_3257,N_1557,N_1342);
and U3258 (N_3258,N_2278,N_2493);
or U3259 (N_3259,N_2407,N_1850);
nand U3260 (N_3260,N_2382,N_2243);
and U3261 (N_3261,N_1453,N_1889);
nand U3262 (N_3262,N_2446,N_2334);
xnor U3263 (N_3263,N_1599,N_1788);
nor U3264 (N_3264,N_1696,N_1488);
or U3265 (N_3265,N_2014,N_1921);
nand U3266 (N_3266,N_2400,N_1472);
or U3267 (N_3267,N_2296,N_2111);
and U3268 (N_3268,N_2350,N_1668);
xnor U3269 (N_3269,N_1937,N_2289);
nand U3270 (N_3270,N_1281,N_1730);
xor U3271 (N_3271,N_2397,N_1446);
nor U3272 (N_3272,N_2145,N_2341);
nor U3273 (N_3273,N_2284,N_1338);
nand U3274 (N_3274,N_1889,N_1757);
and U3275 (N_3275,N_1761,N_2424);
xor U3276 (N_3276,N_2187,N_1928);
and U3277 (N_3277,N_1278,N_1751);
nand U3278 (N_3278,N_2206,N_1555);
and U3279 (N_3279,N_1507,N_1617);
nand U3280 (N_3280,N_1343,N_2324);
xor U3281 (N_3281,N_1329,N_2232);
xnor U3282 (N_3282,N_2491,N_1495);
and U3283 (N_3283,N_2092,N_1272);
nand U3284 (N_3284,N_1289,N_1861);
and U3285 (N_3285,N_2018,N_1328);
or U3286 (N_3286,N_2321,N_1705);
nor U3287 (N_3287,N_2077,N_1842);
or U3288 (N_3288,N_1557,N_2086);
nor U3289 (N_3289,N_1911,N_1459);
nor U3290 (N_3290,N_1954,N_1803);
nor U3291 (N_3291,N_1485,N_2276);
xor U3292 (N_3292,N_1327,N_2158);
and U3293 (N_3293,N_1636,N_1889);
and U3294 (N_3294,N_2362,N_1552);
and U3295 (N_3295,N_1313,N_1599);
xnor U3296 (N_3296,N_2407,N_1635);
nand U3297 (N_3297,N_2321,N_1829);
and U3298 (N_3298,N_1721,N_1741);
and U3299 (N_3299,N_1442,N_1566);
or U3300 (N_3300,N_1593,N_2354);
nor U3301 (N_3301,N_2308,N_2146);
and U3302 (N_3302,N_2494,N_1421);
nor U3303 (N_3303,N_2460,N_1757);
nand U3304 (N_3304,N_1803,N_2300);
nor U3305 (N_3305,N_2432,N_2151);
and U3306 (N_3306,N_1297,N_1481);
nor U3307 (N_3307,N_1696,N_2221);
nor U3308 (N_3308,N_2358,N_1737);
or U3309 (N_3309,N_2152,N_1803);
and U3310 (N_3310,N_1470,N_1966);
nor U3311 (N_3311,N_2444,N_1635);
or U3312 (N_3312,N_1939,N_2154);
and U3313 (N_3313,N_1315,N_2167);
and U3314 (N_3314,N_1965,N_2212);
xnor U3315 (N_3315,N_1488,N_2368);
and U3316 (N_3316,N_2416,N_1998);
nor U3317 (N_3317,N_2448,N_1913);
nand U3318 (N_3318,N_1335,N_1972);
or U3319 (N_3319,N_2218,N_1389);
or U3320 (N_3320,N_1396,N_2162);
or U3321 (N_3321,N_1858,N_1457);
nand U3322 (N_3322,N_1505,N_1486);
nand U3323 (N_3323,N_2438,N_2491);
and U3324 (N_3324,N_1837,N_2436);
or U3325 (N_3325,N_1340,N_1490);
and U3326 (N_3326,N_1963,N_1793);
and U3327 (N_3327,N_2032,N_2297);
xor U3328 (N_3328,N_1495,N_2433);
nand U3329 (N_3329,N_2030,N_2124);
nand U3330 (N_3330,N_2044,N_1751);
nor U3331 (N_3331,N_2038,N_1448);
xor U3332 (N_3332,N_2489,N_1392);
xnor U3333 (N_3333,N_1693,N_2459);
nand U3334 (N_3334,N_2393,N_1833);
nor U3335 (N_3335,N_2223,N_1844);
or U3336 (N_3336,N_1487,N_1803);
nand U3337 (N_3337,N_1643,N_2465);
xor U3338 (N_3338,N_1844,N_1763);
and U3339 (N_3339,N_2017,N_1488);
xnor U3340 (N_3340,N_2241,N_2162);
xor U3341 (N_3341,N_2177,N_2281);
or U3342 (N_3342,N_2029,N_1969);
and U3343 (N_3343,N_1748,N_1612);
and U3344 (N_3344,N_1986,N_1310);
or U3345 (N_3345,N_1405,N_2479);
nand U3346 (N_3346,N_2436,N_2021);
xor U3347 (N_3347,N_2153,N_2192);
xor U3348 (N_3348,N_1514,N_1947);
and U3349 (N_3349,N_1456,N_1286);
or U3350 (N_3350,N_1943,N_1515);
xor U3351 (N_3351,N_1475,N_1523);
and U3352 (N_3352,N_2434,N_1469);
nor U3353 (N_3353,N_1814,N_1963);
or U3354 (N_3354,N_2227,N_1904);
and U3355 (N_3355,N_1737,N_2444);
nand U3356 (N_3356,N_1867,N_1470);
nor U3357 (N_3357,N_2000,N_1782);
nand U3358 (N_3358,N_2400,N_1656);
and U3359 (N_3359,N_1275,N_1323);
nor U3360 (N_3360,N_1530,N_1483);
and U3361 (N_3361,N_2377,N_2460);
nor U3362 (N_3362,N_1321,N_2089);
nand U3363 (N_3363,N_2445,N_1324);
nand U3364 (N_3364,N_2269,N_1652);
nor U3365 (N_3365,N_2341,N_2197);
xnor U3366 (N_3366,N_1643,N_1407);
and U3367 (N_3367,N_1501,N_1766);
nand U3368 (N_3368,N_1673,N_1918);
xnor U3369 (N_3369,N_2008,N_1964);
and U3370 (N_3370,N_2309,N_1503);
nor U3371 (N_3371,N_2323,N_1457);
or U3372 (N_3372,N_1558,N_1682);
nand U3373 (N_3373,N_2400,N_1985);
nand U3374 (N_3374,N_2090,N_2335);
xor U3375 (N_3375,N_1360,N_1852);
or U3376 (N_3376,N_1875,N_1489);
xor U3377 (N_3377,N_2097,N_1819);
or U3378 (N_3378,N_1593,N_2287);
or U3379 (N_3379,N_1273,N_1816);
nand U3380 (N_3380,N_1404,N_2206);
nor U3381 (N_3381,N_2136,N_2256);
or U3382 (N_3382,N_1524,N_1868);
and U3383 (N_3383,N_1451,N_2090);
and U3384 (N_3384,N_2166,N_2149);
or U3385 (N_3385,N_1817,N_2227);
xor U3386 (N_3386,N_2089,N_2401);
xnor U3387 (N_3387,N_2102,N_1372);
and U3388 (N_3388,N_1438,N_2063);
xnor U3389 (N_3389,N_1696,N_1715);
nor U3390 (N_3390,N_1946,N_2264);
xnor U3391 (N_3391,N_1273,N_1388);
or U3392 (N_3392,N_2450,N_1871);
xnor U3393 (N_3393,N_2365,N_1613);
and U3394 (N_3394,N_2032,N_1267);
and U3395 (N_3395,N_1443,N_1269);
and U3396 (N_3396,N_2263,N_1580);
nor U3397 (N_3397,N_2074,N_1619);
and U3398 (N_3398,N_2353,N_1322);
and U3399 (N_3399,N_2318,N_2339);
xnor U3400 (N_3400,N_1411,N_1756);
or U3401 (N_3401,N_2294,N_2325);
or U3402 (N_3402,N_1354,N_1942);
nand U3403 (N_3403,N_1721,N_2137);
nor U3404 (N_3404,N_1426,N_1594);
xor U3405 (N_3405,N_2266,N_2446);
xnor U3406 (N_3406,N_1438,N_1633);
or U3407 (N_3407,N_1905,N_1556);
nand U3408 (N_3408,N_1521,N_2151);
xnor U3409 (N_3409,N_1881,N_1662);
and U3410 (N_3410,N_2102,N_1638);
xor U3411 (N_3411,N_1440,N_1645);
nor U3412 (N_3412,N_2445,N_2274);
nand U3413 (N_3413,N_2153,N_1649);
and U3414 (N_3414,N_1953,N_2096);
and U3415 (N_3415,N_2022,N_2070);
and U3416 (N_3416,N_2048,N_1968);
and U3417 (N_3417,N_2078,N_1648);
and U3418 (N_3418,N_2399,N_1533);
nor U3419 (N_3419,N_1684,N_1370);
nand U3420 (N_3420,N_1589,N_1617);
nor U3421 (N_3421,N_2488,N_2189);
nand U3422 (N_3422,N_1358,N_2258);
and U3423 (N_3423,N_2104,N_1827);
xor U3424 (N_3424,N_2219,N_2025);
nand U3425 (N_3425,N_2151,N_2025);
xnor U3426 (N_3426,N_2442,N_1985);
nand U3427 (N_3427,N_2036,N_1571);
and U3428 (N_3428,N_1731,N_1475);
or U3429 (N_3429,N_2104,N_2323);
and U3430 (N_3430,N_1420,N_1999);
nor U3431 (N_3431,N_2256,N_2117);
nor U3432 (N_3432,N_1946,N_2302);
and U3433 (N_3433,N_2115,N_1426);
nand U3434 (N_3434,N_2449,N_1565);
xor U3435 (N_3435,N_1908,N_1264);
xnor U3436 (N_3436,N_2448,N_2185);
or U3437 (N_3437,N_1504,N_1706);
nor U3438 (N_3438,N_1405,N_1940);
or U3439 (N_3439,N_1663,N_1929);
nor U3440 (N_3440,N_1944,N_1995);
nor U3441 (N_3441,N_2097,N_2357);
nand U3442 (N_3442,N_1932,N_2449);
and U3443 (N_3443,N_2423,N_1858);
nor U3444 (N_3444,N_2422,N_1771);
nand U3445 (N_3445,N_1393,N_2319);
or U3446 (N_3446,N_1594,N_1641);
nor U3447 (N_3447,N_2293,N_1672);
xnor U3448 (N_3448,N_1680,N_2406);
xnor U3449 (N_3449,N_1583,N_1759);
xnor U3450 (N_3450,N_2120,N_2374);
and U3451 (N_3451,N_1684,N_1787);
or U3452 (N_3452,N_1756,N_2323);
xnor U3453 (N_3453,N_2352,N_1869);
or U3454 (N_3454,N_2224,N_1403);
and U3455 (N_3455,N_2451,N_1953);
xnor U3456 (N_3456,N_1290,N_2050);
nand U3457 (N_3457,N_1293,N_2002);
nor U3458 (N_3458,N_1903,N_1618);
or U3459 (N_3459,N_1693,N_1409);
xor U3460 (N_3460,N_1909,N_2271);
nand U3461 (N_3461,N_1817,N_1496);
xor U3462 (N_3462,N_2464,N_2228);
xnor U3463 (N_3463,N_2043,N_1373);
nand U3464 (N_3464,N_1585,N_1849);
nand U3465 (N_3465,N_1804,N_2085);
nand U3466 (N_3466,N_2261,N_1543);
or U3467 (N_3467,N_1830,N_2310);
or U3468 (N_3468,N_2476,N_1631);
and U3469 (N_3469,N_2416,N_1323);
nor U3470 (N_3470,N_2274,N_1255);
nor U3471 (N_3471,N_1621,N_2155);
and U3472 (N_3472,N_2360,N_1805);
and U3473 (N_3473,N_1280,N_1569);
and U3474 (N_3474,N_1837,N_2301);
xnor U3475 (N_3475,N_1289,N_1716);
or U3476 (N_3476,N_2097,N_1287);
or U3477 (N_3477,N_1653,N_2004);
or U3478 (N_3478,N_1378,N_2167);
nor U3479 (N_3479,N_1947,N_1489);
nor U3480 (N_3480,N_1709,N_2455);
xnor U3481 (N_3481,N_2495,N_2072);
nand U3482 (N_3482,N_2315,N_1982);
nor U3483 (N_3483,N_2492,N_2023);
and U3484 (N_3484,N_1541,N_1809);
nand U3485 (N_3485,N_2297,N_2486);
and U3486 (N_3486,N_1449,N_2298);
nor U3487 (N_3487,N_1540,N_2135);
or U3488 (N_3488,N_1691,N_2297);
nand U3489 (N_3489,N_1541,N_2138);
nor U3490 (N_3490,N_1361,N_2158);
xnor U3491 (N_3491,N_2135,N_1479);
nor U3492 (N_3492,N_2019,N_2120);
nand U3493 (N_3493,N_1365,N_1268);
and U3494 (N_3494,N_1966,N_1688);
and U3495 (N_3495,N_1284,N_1705);
nand U3496 (N_3496,N_1924,N_1473);
and U3497 (N_3497,N_2475,N_1671);
or U3498 (N_3498,N_2046,N_2395);
and U3499 (N_3499,N_1255,N_1366);
nand U3500 (N_3500,N_2460,N_1363);
nand U3501 (N_3501,N_1880,N_1361);
nand U3502 (N_3502,N_2482,N_1502);
or U3503 (N_3503,N_1475,N_2454);
xor U3504 (N_3504,N_2407,N_1486);
xor U3505 (N_3505,N_1266,N_1535);
nor U3506 (N_3506,N_1825,N_2428);
or U3507 (N_3507,N_1453,N_1427);
and U3508 (N_3508,N_1800,N_1522);
and U3509 (N_3509,N_2460,N_1558);
nand U3510 (N_3510,N_1389,N_2372);
nor U3511 (N_3511,N_1660,N_1479);
nor U3512 (N_3512,N_2364,N_1696);
nand U3513 (N_3513,N_2420,N_1974);
xnor U3514 (N_3514,N_1367,N_2129);
nor U3515 (N_3515,N_1798,N_2040);
nor U3516 (N_3516,N_2466,N_2277);
nand U3517 (N_3517,N_1573,N_1537);
and U3518 (N_3518,N_1500,N_1597);
or U3519 (N_3519,N_1253,N_1977);
nor U3520 (N_3520,N_2428,N_1332);
or U3521 (N_3521,N_1726,N_2080);
or U3522 (N_3522,N_1677,N_1512);
or U3523 (N_3523,N_1624,N_1352);
nor U3524 (N_3524,N_1853,N_1710);
and U3525 (N_3525,N_2052,N_1622);
xor U3526 (N_3526,N_1395,N_1738);
xnor U3527 (N_3527,N_1443,N_2198);
xor U3528 (N_3528,N_1981,N_1973);
nor U3529 (N_3529,N_1515,N_2436);
xor U3530 (N_3530,N_1436,N_1528);
nand U3531 (N_3531,N_1595,N_2442);
or U3532 (N_3532,N_1810,N_2391);
or U3533 (N_3533,N_1252,N_2012);
nor U3534 (N_3534,N_2142,N_1354);
or U3535 (N_3535,N_1991,N_1827);
xor U3536 (N_3536,N_1276,N_1464);
and U3537 (N_3537,N_1633,N_2300);
nor U3538 (N_3538,N_1337,N_2158);
or U3539 (N_3539,N_2008,N_1750);
or U3540 (N_3540,N_1565,N_1413);
nand U3541 (N_3541,N_1743,N_1566);
and U3542 (N_3542,N_1596,N_1341);
or U3543 (N_3543,N_1917,N_1653);
nor U3544 (N_3544,N_1645,N_1368);
nand U3545 (N_3545,N_1717,N_2333);
nor U3546 (N_3546,N_2078,N_1524);
xnor U3547 (N_3547,N_1575,N_1665);
and U3548 (N_3548,N_1960,N_2250);
and U3549 (N_3549,N_1651,N_1523);
nor U3550 (N_3550,N_1897,N_2069);
xor U3551 (N_3551,N_2372,N_1594);
nor U3552 (N_3552,N_1795,N_1880);
or U3553 (N_3553,N_2047,N_1261);
xnor U3554 (N_3554,N_1358,N_2157);
and U3555 (N_3555,N_2405,N_1517);
or U3556 (N_3556,N_1870,N_2131);
and U3557 (N_3557,N_2287,N_1595);
or U3558 (N_3558,N_1861,N_1725);
nor U3559 (N_3559,N_2254,N_1873);
xor U3560 (N_3560,N_1465,N_2320);
xor U3561 (N_3561,N_1815,N_2314);
or U3562 (N_3562,N_2492,N_1763);
xor U3563 (N_3563,N_1949,N_1469);
xor U3564 (N_3564,N_2083,N_2332);
and U3565 (N_3565,N_1705,N_1648);
nor U3566 (N_3566,N_2223,N_1941);
and U3567 (N_3567,N_1787,N_1753);
nand U3568 (N_3568,N_1777,N_2161);
or U3569 (N_3569,N_2381,N_1377);
nor U3570 (N_3570,N_1359,N_1400);
or U3571 (N_3571,N_2119,N_1262);
and U3572 (N_3572,N_1628,N_1293);
nand U3573 (N_3573,N_2020,N_2058);
nand U3574 (N_3574,N_2319,N_2099);
and U3575 (N_3575,N_1630,N_2245);
or U3576 (N_3576,N_2070,N_2097);
nor U3577 (N_3577,N_1737,N_2130);
and U3578 (N_3578,N_1581,N_2272);
nor U3579 (N_3579,N_1756,N_1785);
nor U3580 (N_3580,N_1886,N_1432);
nand U3581 (N_3581,N_2485,N_1846);
and U3582 (N_3582,N_1446,N_1984);
nand U3583 (N_3583,N_1585,N_1668);
and U3584 (N_3584,N_1426,N_2347);
nand U3585 (N_3585,N_1971,N_2385);
or U3586 (N_3586,N_1854,N_1432);
and U3587 (N_3587,N_1706,N_2491);
or U3588 (N_3588,N_1972,N_1621);
nand U3589 (N_3589,N_1288,N_2332);
and U3590 (N_3590,N_1726,N_2052);
and U3591 (N_3591,N_2447,N_2038);
and U3592 (N_3592,N_1265,N_2327);
nand U3593 (N_3593,N_2107,N_1287);
or U3594 (N_3594,N_1533,N_2056);
and U3595 (N_3595,N_2338,N_1649);
and U3596 (N_3596,N_1731,N_2298);
and U3597 (N_3597,N_2478,N_1367);
nor U3598 (N_3598,N_1464,N_2335);
and U3599 (N_3599,N_1724,N_2342);
xor U3600 (N_3600,N_1809,N_2335);
or U3601 (N_3601,N_2490,N_1368);
nand U3602 (N_3602,N_2468,N_1811);
and U3603 (N_3603,N_1573,N_1606);
or U3604 (N_3604,N_2439,N_2056);
or U3605 (N_3605,N_2307,N_2093);
nand U3606 (N_3606,N_1285,N_1428);
nor U3607 (N_3607,N_1379,N_2452);
nand U3608 (N_3608,N_2107,N_2254);
nand U3609 (N_3609,N_1534,N_1863);
nor U3610 (N_3610,N_2412,N_2328);
xnor U3611 (N_3611,N_1575,N_1442);
nor U3612 (N_3612,N_1698,N_2029);
nor U3613 (N_3613,N_2338,N_1971);
nand U3614 (N_3614,N_2227,N_1900);
or U3615 (N_3615,N_1961,N_2148);
or U3616 (N_3616,N_1599,N_1928);
xor U3617 (N_3617,N_1629,N_1637);
nor U3618 (N_3618,N_1783,N_1574);
and U3619 (N_3619,N_2080,N_1615);
xor U3620 (N_3620,N_1713,N_1597);
and U3621 (N_3621,N_1821,N_1980);
nor U3622 (N_3622,N_1577,N_2210);
and U3623 (N_3623,N_1354,N_2226);
xor U3624 (N_3624,N_1726,N_1670);
nor U3625 (N_3625,N_1822,N_2174);
xor U3626 (N_3626,N_1509,N_2167);
xnor U3627 (N_3627,N_2050,N_1400);
nor U3628 (N_3628,N_1740,N_2163);
nor U3629 (N_3629,N_1276,N_1542);
or U3630 (N_3630,N_1398,N_2286);
or U3631 (N_3631,N_1627,N_1366);
and U3632 (N_3632,N_1352,N_1589);
xor U3633 (N_3633,N_1993,N_1479);
and U3634 (N_3634,N_1661,N_1485);
or U3635 (N_3635,N_1487,N_1817);
nor U3636 (N_3636,N_1547,N_2012);
xor U3637 (N_3637,N_2268,N_2311);
xnor U3638 (N_3638,N_2001,N_1663);
nor U3639 (N_3639,N_1338,N_1319);
xnor U3640 (N_3640,N_2296,N_2484);
xnor U3641 (N_3641,N_2383,N_1352);
nand U3642 (N_3642,N_1284,N_1993);
and U3643 (N_3643,N_1446,N_1749);
or U3644 (N_3644,N_2174,N_1664);
nor U3645 (N_3645,N_1653,N_1459);
and U3646 (N_3646,N_2208,N_2190);
nor U3647 (N_3647,N_2236,N_1485);
and U3648 (N_3648,N_1318,N_1747);
nor U3649 (N_3649,N_2460,N_1815);
and U3650 (N_3650,N_1967,N_1674);
nand U3651 (N_3651,N_1652,N_1299);
and U3652 (N_3652,N_1664,N_1412);
nand U3653 (N_3653,N_1404,N_1713);
or U3654 (N_3654,N_1854,N_1921);
nor U3655 (N_3655,N_1529,N_1850);
and U3656 (N_3656,N_1731,N_2470);
xor U3657 (N_3657,N_2493,N_1381);
and U3658 (N_3658,N_1728,N_2261);
nand U3659 (N_3659,N_1609,N_2267);
and U3660 (N_3660,N_2493,N_1358);
xnor U3661 (N_3661,N_2323,N_1630);
xnor U3662 (N_3662,N_2469,N_2108);
xnor U3663 (N_3663,N_1517,N_1807);
xor U3664 (N_3664,N_1493,N_2292);
nand U3665 (N_3665,N_2419,N_1381);
or U3666 (N_3666,N_1860,N_2243);
nand U3667 (N_3667,N_1962,N_2042);
or U3668 (N_3668,N_1312,N_1487);
or U3669 (N_3669,N_2466,N_1657);
xnor U3670 (N_3670,N_2184,N_1415);
nand U3671 (N_3671,N_2063,N_1502);
nor U3672 (N_3672,N_2108,N_1528);
xor U3673 (N_3673,N_2483,N_1447);
nor U3674 (N_3674,N_2498,N_1669);
nor U3675 (N_3675,N_2006,N_1345);
or U3676 (N_3676,N_2047,N_2203);
or U3677 (N_3677,N_2262,N_2099);
and U3678 (N_3678,N_1662,N_1844);
and U3679 (N_3679,N_1541,N_1642);
or U3680 (N_3680,N_1574,N_1393);
nand U3681 (N_3681,N_2272,N_1401);
or U3682 (N_3682,N_1479,N_1967);
nand U3683 (N_3683,N_2058,N_1815);
nand U3684 (N_3684,N_1563,N_1925);
xnor U3685 (N_3685,N_2089,N_2086);
nand U3686 (N_3686,N_2311,N_1519);
and U3687 (N_3687,N_1498,N_2333);
and U3688 (N_3688,N_1293,N_1701);
or U3689 (N_3689,N_1920,N_1560);
nand U3690 (N_3690,N_2101,N_1386);
or U3691 (N_3691,N_1314,N_1739);
or U3692 (N_3692,N_1890,N_2267);
xor U3693 (N_3693,N_1906,N_1299);
nor U3694 (N_3694,N_2442,N_1484);
or U3695 (N_3695,N_2191,N_2250);
nand U3696 (N_3696,N_1497,N_1395);
nand U3697 (N_3697,N_2102,N_2087);
nor U3698 (N_3698,N_1324,N_2312);
nand U3699 (N_3699,N_1364,N_1842);
nor U3700 (N_3700,N_2287,N_2183);
and U3701 (N_3701,N_1691,N_2086);
nand U3702 (N_3702,N_2220,N_2137);
or U3703 (N_3703,N_1540,N_2354);
nor U3704 (N_3704,N_2189,N_1898);
nand U3705 (N_3705,N_1961,N_1587);
nand U3706 (N_3706,N_1673,N_1969);
xnor U3707 (N_3707,N_1359,N_1899);
or U3708 (N_3708,N_2384,N_1305);
nor U3709 (N_3709,N_1362,N_2164);
or U3710 (N_3710,N_2056,N_2051);
xor U3711 (N_3711,N_1800,N_1755);
and U3712 (N_3712,N_1679,N_1524);
or U3713 (N_3713,N_1688,N_1528);
nor U3714 (N_3714,N_1271,N_2262);
nor U3715 (N_3715,N_2103,N_1673);
and U3716 (N_3716,N_1488,N_2376);
nor U3717 (N_3717,N_1574,N_1519);
xor U3718 (N_3718,N_2465,N_2459);
nor U3719 (N_3719,N_1532,N_2463);
xnor U3720 (N_3720,N_1809,N_2019);
nand U3721 (N_3721,N_1481,N_1870);
or U3722 (N_3722,N_1765,N_2220);
or U3723 (N_3723,N_2410,N_1682);
nand U3724 (N_3724,N_1353,N_2075);
xnor U3725 (N_3725,N_1467,N_2032);
nand U3726 (N_3726,N_2330,N_2194);
xor U3727 (N_3727,N_1725,N_1627);
nor U3728 (N_3728,N_2091,N_1883);
or U3729 (N_3729,N_2203,N_1888);
nand U3730 (N_3730,N_1700,N_2208);
nand U3731 (N_3731,N_2362,N_1588);
or U3732 (N_3732,N_1489,N_1468);
xor U3733 (N_3733,N_2349,N_2405);
and U3734 (N_3734,N_2327,N_1323);
xor U3735 (N_3735,N_1781,N_2161);
or U3736 (N_3736,N_1456,N_1548);
nor U3737 (N_3737,N_1551,N_1321);
nor U3738 (N_3738,N_1762,N_1391);
xnor U3739 (N_3739,N_2267,N_2149);
and U3740 (N_3740,N_1511,N_1502);
and U3741 (N_3741,N_1765,N_1692);
and U3742 (N_3742,N_1739,N_1764);
and U3743 (N_3743,N_2477,N_1628);
and U3744 (N_3744,N_1360,N_2235);
nor U3745 (N_3745,N_1677,N_1907);
or U3746 (N_3746,N_1325,N_2098);
or U3747 (N_3747,N_1625,N_1431);
nand U3748 (N_3748,N_1324,N_1305);
nand U3749 (N_3749,N_2144,N_2458);
xnor U3750 (N_3750,N_3674,N_2660);
and U3751 (N_3751,N_3435,N_2849);
and U3752 (N_3752,N_3685,N_2977);
nand U3753 (N_3753,N_2595,N_3360);
nand U3754 (N_3754,N_3651,N_3513);
xnor U3755 (N_3755,N_3111,N_3305);
nor U3756 (N_3756,N_3638,N_3377);
and U3757 (N_3757,N_3576,N_3125);
nand U3758 (N_3758,N_3494,N_2714);
xnor U3759 (N_3759,N_2774,N_2853);
nand U3760 (N_3760,N_2568,N_3598);
nor U3761 (N_3761,N_3668,N_3337);
xor U3762 (N_3762,N_3283,N_2709);
nand U3763 (N_3763,N_2866,N_2762);
or U3764 (N_3764,N_3041,N_2725);
and U3765 (N_3765,N_3112,N_3147);
and U3766 (N_3766,N_2563,N_3397);
nand U3767 (N_3767,N_3467,N_3134);
nor U3768 (N_3768,N_2843,N_2678);
and U3769 (N_3769,N_2847,N_2918);
and U3770 (N_3770,N_3298,N_3722);
or U3771 (N_3771,N_3120,N_2839);
nand U3772 (N_3772,N_2515,N_3471);
and U3773 (N_3773,N_3060,N_2674);
xnor U3774 (N_3774,N_2684,N_3252);
or U3775 (N_3775,N_3587,N_3361);
nor U3776 (N_3776,N_2830,N_3192);
xor U3777 (N_3777,N_2666,N_3569);
or U3778 (N_3778,N_2689,N_3392);
nor U3779 (N_3779,N_3284,N_2601);
nor U3780 (N_3780,N_2727,N_3364);
nor U3781 (N_3781,N_2531,N_2698);
or U3782 (N_3782,N_2731,N_2621);
and U3783 (N_3783,N_3222,N_2676);
nand U3784 (N_3784,N_3512,N_3458);
nand U3785 (N_3785,N_3716,N_3052);
nor U3786 (N_3786,N_2672,N_3531);
nand U3787 (N_3787,N_3537,N_3078);
xor U3788 (N_3788,N_3621,N_3406);
nand U3789 (N_3789,N_2862,N_3708);
nand U3790 (N_3790,N_3426,N_3143);
or U3791 (N_3791,N_3221,N_3092);
or U3792 (N_3792,N_3415,N_3084);
xnor U3793 (N_3793,N_3737,N_3522);
xnor U3794 (N_3794,N_3170,N_3289);
xor U3795 (N_3795,N_3367,N_3282);
xor U3796 (N_3796,N_2708,N_3586);
or U3797 (N_3797,N_3131,N_2986);
nor U3798 (N_3798,N_3195,N_3212);
nor U3799 (N_3799,N_2651,N_3074);
or U3800 (N_3800,N_2985,N_2603);
nand U3801 (N_3801,N_2873,N_2939);
or U3802 (N_3802,N_2613,N_3332);
and U3803 (N_3803,N_3632,N_3343);
xor U3804 (N_3804,N_3623,N_3509);
or U3805 (N_3805,N_3323,N_2569);
nand U3806 (N_3806,N_3382,N_3101);
or U3807 (N_3807,N_3521,N_3163);
nor U3808 (N_3808,N_3354,N_2822);
nor U3809 (N_3809,N_3327,N_3519);
nor U3810 (N_3810,N_2771,N_3404);
or U3811 (N_3811,N_2649,N_2742);
xnor U3812 (N_3812,N_3613,N_3579);
xnor U3813 (N_3813,N_3302,N_3237);
nand U3814 (N_3814,N_3504,N_2823);
nand U3815 (N_3815,N_3183,N_2671);
xnor U3816 (N_3816,N_2863,N_2722);
xnor U3817 (N_3817,N_2712,N_3691);
or U3818 (N_3818,N_3194,N_2753);
or U3819 (N_3819,N_2883,N_3244);
nor U3820 (N_3820,N_2658,N_3176);
or U3821 (N_3821,N_2574,N_3622);
xnor U3822 (N_3822,N_2735,N_3083);
nor U3823 (N_3823,N_3507,N_2656);
and U3824 (N_3824,N_3725,N_3312);
nor U3825 (N_3825,N_2917,N_3380);
xnor U3826 (N_3826,N_2590,N_3081);
nand U3827 (N_3827,N_2903,N_3420);
nand U3828 (N_3828,N_3270,N_3217);
nor U3829 (N_3829,N_3259,N_2836);
xnor U3830 (N_3830,N_2667,N_3291);
nor U3831 (N_3831,N_3501,N_2895);
nor U3832 (N_3832,N_2987,N_3310);
xnor U3833 (N_3833,N_3581,N_3373);
nor U3834 (N_3834,N_2891,N_3738);
nor U3835 (N_3835,N_3491,N_2653);
nand U3836 (N_3836,N_2793,N_3311);
xnor U3837 (N_3837,N_3599,N_2537);
and U3838 (N_3838,N_3269,N_2910);
nand U3839 (N_3839,N_3432,N_3096);
nand U3840 (N_3840,N_3144,N_3091);
xnor U3841 (N_3841,N_2788,N_3550);
xnor U3842 (N_3842,N_2796,N_3324);
nand U3843 (N_3843,N_2690,N_3330);
xnor U3844 (N_3844,N_3247,N_2705);
and U3845 (N_3845,N_2506,N_3308);
xor U3846 (N_3846,N_2966,N_3662);
and U3847 (N_3847,N_3139,N_2805);
and U3848 (N_3848,N_2645,N_3505);
nand U3849 (N_3849,N_3022,N_3715);
nor U3850 (N_3850,N_3487,N_3107);
xnor U3851 (N_3851,N_3309,N_3255);
nand U3852 (N_3852,N_3490,N_2553);
and U3853 (N_3853,N_2756,N_2973);
or U3854 (N_3854,N_3655,N_3293);
nor U3855 (N_3855,N_2661,N_3079);
nand U3856 (N_3856,N_2813,N_2535);
nand U3857 (N_3857,N_3077,N_3428);
nor U3858 (N_3858,N_3606,N_2975);
xor U3859 (N_3859,N_2600,N_3369);
nand U3860 (N_3860,N_3429,N_3085);
nor U3861 (N_3861,N_2767,N_3439);
xor U3862 (N_3862,N_3719,N_2730);
or U3863 (N_3863,N_3117,N_2953);
nand U3864 (N_3864,N_3390,N_3640);
nand U3865 (N_3865,N_2933,N_3393);
xnor U3866 (N_3866,N_2854,N_3158);
nand U3867 (N_3867,N_2631,N_2625);
and U3868 (N_3868,N_2510,N_2532);
nand U3869 (N_3869,N_3648,N_2720);
or U3870 (N_3870,N_3704,N_2865);
xnor U3871 (N_3871,N_2913,N_2588);
nand U3872 (N_3872,N_2525,N_2773);
nand U3873 (N_3873,N_2809,N_2996);
nor U3874 (N_3874,N_2812,N_2707);
nor U3875 (N_3875,N_2834,N_3645);
and U3876 (N_3876,N_2925,N_2587);
xnor U3877 (N_3877,N_3724,N_2875);
nand U3878 (N_3878,N_3307,N_2626);
nor U3879 (N_3879,N_3503,N_2501);
nand U3880 (N_3880,N_2604,N_2940);
xor U3881 (N_3881,N_2633,N_2923);
or U3882 (N_3882,N_3488,N_3625);
or U3883 (N_3883,N_2580,N_3654);
nor U3884 (N_3884,N_2792,N_2696);
xnor U3885 (N_3885,N_3510,N_3065);
nor U3886 (N_3886,N_2824,N_3043);
or U3887 (N_3887,N_3669,N_2900);
or U3888 (N_3888,N_3478,N_2745);
and U3889 (N_3889,N_3624,N_2963);
nor U3890 (N_3890,N_2710,N_3229);
nand U3891 (N_3891,N_3464,N_3299);
xor U3892 (N_3892,N_2964,N_3126);
or U3893 (N_3893,N_2775,N_2544);
nor U3894 (N_3894,N_3495,N_2572);
nand U3895 (N_3895,N_3303,N_2747);
or U3896 (N_3896,N_3591,N_3383);
and U3897 (N_3897,N_3540,N_3474);
and U3898 (N_3898,N_2789,N_3355);
and U3899 (N_3899,N_2970,N_2648);
or U3900 (N_3900,N_3167,N_3518);
nor U3901 (N_3901,N_3408,N_3683);
xnor U3902 (N_3902,N_3658,N_3571);
and U3903 (N_3903,N_3054,N_2871);
or U3904 (N_3904,N_2691,N_3376);
nand U3905 (N_3905,N_2508,N_2785);
and U3906 (N_3906,N_3580,N_3027);
or U3907 (N_3907,N_3350,N_2548);
and U3908 (N_3908,N_3690,N_3209);
xnor U3909 (N_3909,N_3066,N_3525);
nand U3910 (N_3910,N_3527,N_2882);
or U3911 (N_3911,N_3560,N_2706);
nand U3912 (N_3912,N_3447,N_3430);
and U3913 (N_3913,N_3403,N_2579);
xor U3914 (N_3914,N_2784,N_3193);
nand U3915 (N_3915,N_2962,N_2791);
and U3916 (N_3916,N_2860,N_2993);
nand U3917 (N_3917,N_3739,N_3391);
and U3918 (N_3918,N_2619,N_3394);
nand U3919 (N_3919,N_3486,N_2960);
xor U3920 (N_3920,N_2934,N_2602);
nor U3921 (N_3921,N_3075,N_3089);
nand U3922 (N_3922,N_3335,N_3529);
and U3923 (N_3923,N_3206,N_3196);
or U3924 (N_3924,N_3040,N_3438);
xnor U3925 (N_3925,N_3263,N_3733);
nand U3926 (N_3926,N_2897,N_2904);
nand U3927 (N_3927,N_2827,N_3100);
nor U3928 (N_3928,N_2555,N_3127);
nor U3929 (N_3929,N_3694,N_3460);
nor U3930 (N_3930,N_3031,N_2754);
nor U3931 (N_3931,N_3549,N_2598);
nor U3932 (N_3932,N_2743,N_2867);
nor U3933 (N_3933,N_3204,N_2577);
nand U3934 (N_3934,N_2591,N_2641);
or U3935 (N_3935,N_2978,N_2635);
or U3936 (N_3936,N_3233,N_2726);
nand U3937 (N_3937,N_3646,N_2787);
xnor U3938 (N_3938,N_2810,N_3681);
or U3939 (N_3939,N_2562,N_3703);
or U3940 (N_3940,N_3628,N_3747);
nor U3941 (N_3941,N_3046,N_3427);
nor U3942 (N_3942,N_2552,N_2816);
xor U3943 (N_3943,N_3370,N_3697);
or U3944 (N_3944,N_3250,N_3542);
and U3945 (N_3945,N_3556,N_2772);
or U3946 (N_3946,N_2794,N_2589);
nand U3947 (N_3947,N_3215,N_3320);
or U3948 (N_3948,N_2502,N_2768);
nand U3949 (N_3949,N_3496,N_3558);
and U3950 (N_3950,N_3457,N_3459);
nor U3951 (N_3951,N_2540,N_3258);
and U3952 (N_3952,N_3168,N_3082);
and U3953 (N_3953,N_3614,N_2517);
or U3954 (N_3954,N_2680,N_3468);
nor U3955 (N_3955,N_3326,N_3076);
xnor U3956 (N_3956,N_3453,N_2814);
or U3957 (N_3957,N_2738,N_2734);
nand U3958 (N_3958,N_2677,N_2872);
nand U3959 (N_3959,N_3200,N_3275);
and U3960 (N_3960,N_3469,N_3484);
xor U3961 (N_3961,N_2838,N_2636);
and U3962 (N_3962,N_3174,N_3064);
nand U3963 (N_3963,N_2869,N_2575);
xnor U3964 (N_3964,N_3345,N_3223);
and U3965 (N_3965,N_3595,N_3421);
and U3966 (N_3966,N_3620,N_3541);
xor U3967 (N_3967,N_3665,N_3166);
nor U3968 (N_3968,N_3021,N_2521);
and U3969 (N_3969,N_3678,N_2956);
nor U3970 (N_3970,N_3189,N_3635);
and U3971 (N_3971,N_2640,N_3449);
and U3972 (N_3972,N_3677,N_2536);
or U3973 (N_3973,N_2549,N_3265);
nand U3974 (N_3974,N_3007,N_2647);
nor U3975 (N_3975,N_3561,N_3175);
nand U3976 (N_3976,N_3604,N_2711);
nor U3977 (N_3977,N_3615,N_3012);
and U3978 (N_3978,N_3729,N_2652);
nand U3979 (N_3979,N_2991,N_3389);
nor U3980 (N_3980,N_3372,N_3379);
nor U3981 (N_3981,N_2976,N_2766);
and U3982 (N_3982,N_3524,N_2650);
nand U3983 (N_3983,N_2682,N_3019);
nand U3984 (N_3984,N_3619,N_3673);
xnor U3985 (N_3985,N_3042,N_2947);
or U3986 (N_3986,N_3161,N_2831);
xor U3987 (N_3987,N_2717,N_2783);
nand U3988 (N_3988,N_3115,N_2622);
nand U3989 (N_3989,N_2924,N_3543);
nand U3990 (N_3990,N_3441,N_2874);
nor U3991 (N_3991,N_3319,N_2686);
xnor U3992 (N_3992,N_3515,N_3349);
nand U3993 (N_3993,N_3262,N_3545);
nor U3994 (N_3994,N_3000,N_2921);
nand U3995 (N_3995,N_3231,N_2550);
xor U3996 (N_3996,N_3631,N_2505);
nor U3997 (N_3997,N_3274,N_3108);
and U3998 (N_3998,N_3741,N_2718);
nand U3999 (N_3999,N_3295,N_3506);
nand U4000 (N_4000,N_3557,N_2643);
or U4001 (N_4001,N_3664,N_3347);
nand U4002 (N_4002,N_3016,N_3154);
or U4003 (N_4003,N_2967,N_2901);
nor U4004 (N_4004,N_3051,N_3172);
or U4005 (N_4005,N_3136,N_3607);
xor U4006 (N_4006,N_3718,N_3080);
nand U4007 (N_4007,N_2832,N_2545);
or U4008 (N_4008,N_2994,N_3009);
xor U4009 (N_4009,N_3698,N_2530);
nor U4010 (N_4010,N_2606,N_2906);
or U4011 (N_4011,N_2868,N_2770);
and U4012 (N_4012,N_3516,N_2581);
nand U4013 (N_4013,N_3570,N_3709);
nor U4014 (N_4014,N_2748,N_2632);
and U4015 (N_4015,N_3732,N_2551);
and U4016 (N_4016,N_3058,N_2703);
nor U4017 (N_4017,N_3687,N_3436);
nand U4018 (N_4018,N_2559,N_3735);
and U4019 (N_4019,N_2937,N_3601);
nand U4020 (N_4020,N_3734,N_2802);
xor U4021 (N_4021,N_3353,N_2943);
xnor U4022 (N_4022,N_2858,N_2915);
nor U4023 (N_4023,N_3329,N_3650);
and U4024 (N_4024,N_3339,N_2841);
xor U4025 (N_4025,N_3700,N_2905);
nand U4026 (N_4026,N_2929,N_2571);
xnor U4027 (N_4027,N_3135,N_3608);
or U4028 (N_4028,N_2842,N_3358);
or U4029 (N_4029,N_3220,N_2765);
and U4030 (N_4030,N_3742,N_2700);
and U4031 (N_4031,N_2657,N_2739);
nor U4032 (N_4032,N_2557,N_3014);
nor U4033 (N_4033,N_3029,N_3564);
or U4034 (N_4034,N_3644,N_3670);
or U4035 (N_4035,N_3264,N_3036);
nor U4036 (N_4036,N_2538,N_3417);
and U4037 (N_4037,N_3479,N_3407);
or U4038 (N_4038,N_3256,N_2926);
or U4039 (N_4039,N_3248,N_3304);
nor U4040 (N_4040,N_3184,N_3149);
or U4041 (N_4041,N_2744,N_2879);
nand U4042 (N_4042,N_3371,N_2578);
xnor U4043 (N_4043,N_2899,N_3726);
xor U4044 (N_4044,N_3554,N_3642);
xor U4045 (N_4045,N_3536,N_3517);
nand U4046 (N_4046,N_2611,N_3097);
nor U4047 (N_4047,N_2694,N_2896);
nor U4048 (N_4048,N_3203,N_3321);
xnor U4049 (N_4049,N_3705,N_2751);
nand U4050 (N_4050,N_2629,N_2804);
nor U4051 (N_4051,N_3093,N_3113);
xnor U4052 (N_4052,N_2527,N_3348);
or U4053 (N_4053,N_3476,N_3450);
and U4054 (N_4054,N_3497,N_3008);
or U4055 (N_4055,N_2570,N_3446);
xor U4056 (N_4056,N_3612,N_3099);
xnor U4057 (N_4057,N_3400,N_3443);
xor U4058 (N_4058,N_3466,N_3288);
nor U4059 (N_4059,N_2876,N_2932);
xor U4060 (N_4060,N_3359,N_3649);
or U4061 (N_4061,N_3573,N_3226);
xnor U4062 (N_4062,N_2945,N_3205);
nor U4063 (N_4063,N_2980,N_3338);
xnor U4064 (N_4064,N_3475,N_2669);
nand U4065 (N_4065,N_3328,N_2884);
and U4066 (N_4066,N_2961,N_3013);
nor U4067 (N_4067,N_3489,N_2630);
xnor U4068 (N_4068,N_3603,N_3260);
nor U4069 (N_4069,N_3656,N_2586);
nor U4070 (N_4070,N_2807,N_2803);
xnor U4071 (N_4071,N_2662,N_2995);
xnor U4072 (N_4072,N_3562,N_2668);
nor U4073 (N_4073,N_3552,N_2776);
and U4074 (N_4074,N_3300,N_3480);
xor U4075 (N_4075,N_2779,N_2886);
or U4076 (N_4076,N_3234,N_3045);
and U4077 (N_4077,N_3728,N_3218);
and U4078 (N_4078,N_2971,N_2997);
and U4079 (N_4079,N_3362,N_2642);
nor U4080 (N_4080,N_3254,N_3721);
xor U4081 (N_4081,N_2732,N_3210);
and U4082 (N_4082,N_3104,N_2584);
nand U4083 (N_4083,N_3508,N_2713);
nand U4084 (N_4084,N_3130,N_3098);
and U4085 (N_4085,N_3156,N_3633);
or U4086 (N_4086,N_2808,N_3006);
nor U4087 (N_4087,N_3740,N_3088);
or U4088 (N_4088,N_2881,N_3179);
nor U4089 (N_4089,N_3609,N_3266);
or U4090 (N_4090,N_2935,N_3267);
nor U4091 (N_4091,N_3588,N_2931);
and U4092 (N_4092,N_2780,N_3368);
and U4093 (N_4093,N_2981,N_3463);
and U4094 (N_4094,N_2972,N_2556);
or U4095 (N_4095,N_3731,N_2692);
and U4096 (N_4096,N_3546,N_2654);
or U4097 (N_4097,N_3346,N_2543);
and U4098 (N_4098,N_3675,N_3555);
nor U4099 (N_4099,N_3461,N_2582);
nand U4100 (N_4100,N_2952,N_2646);
nand U4101 (N_4101,N_3211,N_3015);
and U4102 (N_4102,N_3138,N_3511);
xnor U4103 (N_4103,N_2982,N_3301);
nor U4104 (N_4104,N_2704,N_3157);
and U4105 (N_4105,N_3273,N_3693);
or U4106 (N_4106,N_2944,N_3087);
nand U4107 (N_4107,N_3745,N_2844);
or U4108 (N_4108,N_3230,N_2907);
or U4109 (N_4109,N_3069,N_3431);
nand U4110 (N_4110,N_3336,N_3243);
and U4111 (N_4111,N_2781,N_3473);
nor U4112 (N_4112,N_2815,N_3657);
or U4113 (N_4113,N_3412,N_3122);
or U4114 (N_4114,N_2968,N_3224);
or U4115 (N_4115,N_3162,N_3095);
and U4116 (N_4116,N_3035,N_2818);
and U4117 (N_4117,N_2512,N_3018);
or U4118 (N_4118,N_2992,N_2833);
xnor U4119 (N_4119,N_2511,N_3239);
nand U4120 (N_4120,N_3410,N_3433);
nand U4121 (N_4121,N_3315,N_3180);
nand U4122 (N_4122,N_2679,N_2859);
or U4123 (N_4123,N_3748,N_3137);
nor U4124 (N_4124,N_3434,N_2909);
or U4125 (N_4125,N_2688,N_2988);
nand U4126 (N_4126,N_3148,N_2524);
nand U4127 (N_4127,N_3232,N_2507);
and U4128 (N_4128,N_3236,N_3145);
xnor U4129 (N_4129,N_2889,N_3197);
nor U4130 (N_4130,N_2723,N_3672);
and U4131 (N_4131,N_3198,N_3245);
or U4132 (N_4132,N_3689,N_3589);
xnor U4133 (N_4133,N_3749,N_3228);
and U4134 (N_4134,N_2801,N_2520);
nor U4135 (N_4135,N_3584,N_3544);
or U4136 (N_4136,N_2673,N_2761);
nor U4137 (N_4137,N_3056,N_2855);
or U4138 (N_4138,N_3566,N_2795);
nor U4139 (N_4139,N_3444,N_3574);
or U4140 (N_4140,N_3271,N_3318);
xor U4141 (N_4141,N_3024,N_3647);
nor U4142 (N_4142,N_3707,N_2541);
and U4143 (N_4143,N_3044,N_3050);
or U4144 (N_4144,N_3695,N_3702);
or U4145 (N_4145,N_3068,N_2954);
and U4146 (N_4146,N_3538,N_3272);
nor U4147 (N_4147,N_3374,N_3711);
nand U4148 (N_4148,N_3568,N_3238);
xnor U4149 (N_4149,N_2638,N_3004);
and U4150 (N_4150,N_3061,N_3032);
and U4151 (N_4151,N_2983,N_2529);
and U4152 (N_4152,N_3578,N_2659);
nor U4153 (N_4153,N_3306,N_2979);
xor U4154 (N_4154,N_3661,N_2701);
nor U4155 (N_4155,N_3292,N_3381);
xor U4156 (N_4156,N_3634,N_2885);
or U4157 (N_4157,N_2573,N_3639);
nor U4158 (N_4158,N_3023,N_2644);
and U4159 (N_4159,N_3090,N_3616);
xor U4160 (N_4160,N_2503,N_3548);
nor U4161 (N_4161,N_3641,N_2856);
or U4162 (N_4162,N_2914,N_2697);
xnor U4163 (N_4163,N_3261,N_3325);
and U4164 (N_4164,N_3164,N_2655);
and U4165 (N_4165,N_3499,N_3001);
nand U4166 (N_4166,N_3626,N_2628);
and U4167 (N_4167,N_2817,N_2615);
and U4168 (N_4168,N_3413,N_3398);
and U4169 (N_4169,N_3280,N_2514);
xnor U4170 (N_4170,N_2695,N_2504);
nand U4171 (N_4171,N_2702,N_3534);
xor U4172 (N_4172,N_2685,N_3340);
and U4173 (N_4173,N_3106,N_3297);
and U4174 (N_4174,N_3186,N_3409);
nor U4175 (N_4175,N_3020,N_2806);
nor U4176 (N_4176,N_2821,N_2533);
nand U4177 (N_4177,N_2811,N_2547);
nor U4178 (N_4178,N_2612,N_3590);
nand U4179 (N_4179,N_3208,N_2893);
and U4180 (N_4180,N_3153,N_3314);
nand U4181 (N_4181,N_3105,N_3713);
nand U4182 (N_4182,N_3442,N_2759);
nor U4183 (N_4183,N_3744,N_3257);
xor U4184 (N_4184,N_2820,N_3202);
xor U4185 (N_4185,N_3706,N_3627);
nor U4186 (N_4186,N_3701,N_2825);
and U4187 (N_4187,N_3313,N_3492);
or U4188 (N_4188,N_3034,N_2764);
nor U4189 (N_4189,N_3684,N_2758);
nor U4190 (N_4190,N_3386,N_3414);
nor U4191 (N_4191,N_3481,N_3063);
nand U4192 (N_4192,N_3214,N_2597);
nand U4193 (N_4193,N_3454,N_2786);
or U4194 (N_4194,N_2888,N_3227);
nor U4195 (N_4195,N_3010,N_2675);
or U4196 (N_4196,N_2737,N_2887);
and U4197 (N_4197,N_3276,N_2528);
or U4198 (N_4198,N_2599,N_3026);
nor U4199 (N_4199,N_2741,N_3567);
or U4200 (N_4200,N_3643,N_2769);
nand U4201 (N_4201,N_2681,N_3539);
nor U4202 (N_4202,N_2878,N_2782);
xor U4203 (N_4203,N_3720,N_3387);
xor U4204 (N_4204,N_3660,N_3151);
and U4205 (N_4205,N_3388,N_3671);
nand U4206 (N_4206,N_3177,N_3094);
or U4207 (N_4207,N_2850,N_2687);
and U4208 (N_4208,N_3178,N_2938);
xor U4209 (N_4209,N_3611,N_3652);
and U4210 (N_4210,N_3416,N_3493);
or U4211 (N_4211,N_3047,N_3352);
nand U4212 (N_4212,N_3746,N_3235);
or U4213 (N_4213,N_3344,N_3422);
nor U4214 (N_4214,N_3563,N_3448);
and U4215 (N_4215,N_3577,N_2920);
or U4216 (N_4216,N_3712,N_2852);
nand U4217 (N_4217,N_3470,N_3455);
or U4218 (N_4218,N_2663,N_2800);
nor U4219 (N_4219,N_3680,N_3067);
or U4220 (N_4220,N_2519,N_2592);
nand U4221 (N_4221,N_2620,N_3532);
and U4222 (N_4222,N_3028,N_2513);
or U4223 (N_4223,N_3666,N_2951);
xor U4224 (N_4224,N_3251,N_2639);
nand U4225 (N_4225,N_3249,N_2919);
nand U4226 (N_4226,N_2627,N_3618);
nor U4227 (N_4227,N_3437,N_3341);
xnor U4228 (N_4228,N_3378,N_3600);
nand U4229 (N_4229,N_3073,N_3395);
nand U4230 (N_4230,N_2716,N_3278);
nor U4231 (N_4231,N_2797,N_2567);
and U4232 (N_4232,N_3692,N_3456);
nand U4233 (N_4233,N_2728,N_2936);
and U4234 (N_4234,N_3225,N_3190);
nand U4235 (N_4235,N_2892,N_3216);
or U4236 (N_4236,N_3401,N_3294);
nand U4237 (N_4237,N_3357,N_3743);
nor U4238 (N_4238,N_2683,N_3502);
nor U4239 (N_4239,N_2605,N_2583);
nand U4240 (N_4240,N_3285,N_2509);
xnor U4241 (N_4241,N_2607,N_3002);
and U4242 (N_4242,N_2616,N_2777);
nor U4243 (N_4243,N_3559,N_3005);
or U4244 (N_4244,N_2526,N_3688);
and U4245 (N_4245,N_2984,N_3356);
and U4246 (N_4246,N_3485,N_3116);
nand U4247 (N_4247,N_3637,N_3366);
xor U4248 (N_4248,N_3482,N_3605);
xnor U4249 (N_4249,N_3201,N_3452);
or U4250 (N_4250,N_3551,N_3363);
nand U4251 (N_4251,N_2958,N_3679);
xor U4252 (N_4252,N_2916,N_2826);
nor U4253 (N_4253,N_3425,N_3440);
nor U4254 (N_4254,N_2927,N_3317);
nor U4255 (N_4255,N_2594,N_3057);
nand U4256 (N_4256,N_3523,N_2928);
or U4257 (N_4257,N_3402,N_3017);
nand U4258 (N_4258,N_3171,N_3062);
xnor U4259 (N_4259,N_2848,N_3121);
xnor U4260 (N_4260,N_2665,N_3472);
nand U4261 (N_4261,N_2864,N_2908);
and U4262 (N_4262,N_2790,N_3533);
xnor U4263 (N_4263,N_2546,N_2560);
nand U4264 (N_4264,N_3636,N_3119);
or U4265 (N_4265,N_3181,N_2752);
xnor U4266 (N_4266,N_3253,N_2624);
nand U4267 (N_4267,N_2840,N_3142);
and U4268 (N_4268,N_3055,N_2990);
or U4269 (N_4269,N_2949,N_2554);
or U4270 (N_4270,N_2558,N_2942);
and U4271 (N_4271,N_3160,N_2999);
xnor U4272 (N_4272,N_2890,N_3037);
nand U4273 (N_4273,N_3268,N_3146);
nor U4274 (N_4274,N_3128,N_2846);
nand U4275 (N_4275,N_3039,N_3240);
nor U4276 (N_4276,N_3241,N_2617);
or U4277 (N_4277,N_2749,N_3290);
xnor U4278 (N_4278,N_3699,N_3059);
nand U4279 (N_4279,N_3025,N_2946);
and U4280 (N_4280,N_3405,N_2637);
or U4281 (N_4281,N_2880,N_3424);
or U4282 (N_4282,N_3477,N_3445);
and U4283 (N_4283,N_3583,N_3281);
nor U4284 (N_4284,N_3110,N_2835);
nor U4285 (N_4285,N_3682,N_2596);
nand U4286 (N_4286,N_3331,N_2912);
xnor U4287 (N_4287,N_2757,N_3686);
xnor U4288 (N_4288,N_3498,N_3030);
nand U4289 (N_4289,N_3322,N_3246);
or U4290 (N_4290,N_3053,N_3411);
nand U4291 (N_4291,N_3048,N_2715);
or U4292 (N_4292,N_3334,N_2719);
nor U4293 (N_4293,N_2564,N_2778);
nand U4294 (N_4294,N_2957,N_2736);
and U4295 (N_4295,N_3535,N_3730);
nor U4296 (N_4296,N_2950,N_3483);
nor U4297 (N_4297,N_3597,N_2941);
and U4298 (N_4298,N_2837,N_2500);
nand U4299 (N_4299,N_2798,N_3736);
nor U4300 (N_4300,N_3242,N_3103);
and U4301 (N_4301,N_3173,N_2516);
nor U4302 (N_4302,N_2699,N_3592);
and U4303 (N_4303,N_2565,N_3528);
nand U4304 (N_4304,N_2542,N_3629);
nand U4305 (N_4305,N_2634,N_3582);
xor U4306 (N_4306,N_2861,N_2877);
or U4307 (N_4307,N_2763,N_3526);
and U4308 (N_4308,N_3109,N_2755);
nand U4309 (N_4309,N_2955,N_3114);
nand U4310 (N_4310,N_3710,N_2539);
or U4311 (N_4311,N_2609,N_3132);
and U4312 (N_4312,N_3617,N_3165);
xor U4313 (N_4313,N_3553,N_3500);
xnor U4314 (N_4314,N_3033,N_2911);
or U4315 (N_4315,N_2828,N_3071);
or U4316 (N_4316,N_2989,N_3602);
or U4317 (N_4317,N_3011,N_3219);
xor U4318 (N_4318,N_2898,N_3199);
and U4319 (N_4319,N_3396,N_3049);
or U4320 (N_4320,N_2610,N_2566);
nor U4321 (N_4321,N_2534,N_3714);
xnor U4322 (N_4322,N_3610,N_2670);
or U4323 (N_4323,N_3572,N_2894);
and U4324 (N_4324,N_2959,N_2522);
nor U4325 (N_4325,N_3169,N_2746);
or U4326 (N_4326,N_2724,N_3723);
and U4327 (N_4327,N_3659,N_2576);
and U4328 (N_4328,N_3086,N_3585);
nor U4329 (N_4329,N_3277,N_2585);
nand U4330 (N_4330,N_3279,N_3696);
nor U4331 (N_4331,N_2614,N_3565);
or U4332 (N_4332,N_2851,N_2729);
nand U4333 (N_4333,N_3333,N_3123);
xnor U4334 (N_4334,N_3418,N_2930);
nand U4335 (N_4335,N_3520,N_2799);
nor U4336 (N_4336,N_3102,N_2922);
xor U4337 (N_4337,N_2948,N_2664);
nor U4338 (N_4338,N_2857,N_2740);
xnor U4339 (N_4339,N_2998,N_3072);
and U4340 (N_4340,N_3187,N_3593);
and U4341 (N_4341,N_3653,N_3419);
nor U4342 (N_4342,N_3375,N_3185);
nor U4343 (N_4343,N_3451,N_3594);
xor U4344 (N_4344,N_2965,N_3399);
and U4345 (N_4345,N_3667,N_3596);
nand U4346 (N_4346,N_3038,N_3129);
or U4347 (N_4347,N_2518,N_3286);
or U4348 (N_4348,N_3150,N_3630);
nand U4349 (N_4349,N_2969,N_2819);
nor U4350 (N_4350,N_3727,N_2623);
nor U4351 (N_4351,N_3365,N_3159);
and U4352 (N_4352,N_3124,N_3003);
and U4353 (N_4353,N_2845,N_3070);
nor U4354 (N_4354,N_3140,N_2523);
nor U4355 (N_4355,N_3207,N_2608);
xor U4356 (N_4356,N_3717,N_2561);
nand U4357 (N_4357,N_3530,N_3547);
and U4358 (N_4358,N_3287,N_3342);
xnor U4359 (N_4359,N_3188,N_3118);
and U4360 (N_4360,N_3465,N_2750);
and U4361 (N_4361,N_3385,N_3182);
and U4362 (N_4362,N_3213,N_2721);
xnor U4363 (N_4363,N_3514,N_3133);
xor U4364 (N_4364,N_3191,N_3152);
and U4365 (N_4365,N_3155,N_3316);
xnor U4366 (N_4366,N_3462,N_2902);
xnor U4367 (N_4367,N_2760,N_3351);
and U4368 (N_4368,N_3141,N_3663);
nor U4369 (N_4369,N_2593,N_3296);
or U4370 (N_4370,N_2733,N_3384);
and U4371 (N_4371,N_2618,N_3423);
nand U4372 (N_4372,N_3575,N_2974);
nand U4373 (N_4373,N_2870,N_3676);
nor U4374 (N_4374,N_2829,N_2693);
nor U4375 (N_4375,N_3097,N_2577);
or U4376 (N_4376,N_3422,N_2519);
nand U4377 (N_4377,N_3097,N_2899);
or U4378 (N_4378,N_3569,N_3083);
nor U4379 (N_4379,N_2846,N_3616);
or U4380 (N_4380,N_3696,N_3244);
xor U4381 (N_4381,N_3378,N_2678);
xnor U4382 (N_4382,N_2743,N_3247);
nor U4383 (N_4383,N_3629,N_3486);
or U4384 (N_4384,N_3084,N_2615);
and U4385 (N_4385,N_3641,N_3072);
nand U4386 (N_4386,N_3209,N_3688);
nor U4387 (N_4387,N_3483,N_3636);
or U4388 (N_4388,N_3061,N_3020);
xor U4389 (N_4389,N_3000,N_3221);
xor U4390 (N_4390,N_3317,N_3492);
or U4391 (N_4391,N_3371,N_3622);
nor U4392 (N_4392,N_3340,N_3165);
nand U4393 (N_4393,N_2655,N_2575);
and U4394 (N_4394,N_3336,N_3444);
or U4395 (N_4395,N_2683,N_3464);
nor U4396 (N_4396,N_2881,N_3206);
and U4397 (N_4397,N_3726,N_3224);
and U4398 (N_4398,N_3625,N_3627);
and U4399 (N_4399,N_3409,N_2908);
and U4400 (N_4400,N_3106,N_3636);
nand U4401 (N_4401,N_3622,N_2704);
and U4402 (N_4402,N_2990,N_3665);
or U4403 (N_4403,N_3395,N_3119);
and U4404 (N_4404,N_3633,N_3741);
nand U4405 (N_4405,N_2662,N_2675);
nor U4406 (N_4406,N_2634,N_3211);
nor U4407 (N_4407,N_3234,N_3745);
and U4408 (N_4408,N_2617,N_3053);
nand U4409 (N_4409,N_3633,N_2611);
nand U4410 (N_4410,N_2539,N_3174);
or U4411 (N_4411,N_3337,N_3232);
nor U4412 (N_4412,N_3153,N_2781);
xor U4413 (N_4413,N_3120,N_3114);
nor U4414 (N_4414,N_3275,N_2600);
nand U4415 (N_4415,N_3616,N_3434);
nor U4416 (N_4416,N_3521,N_3631);
and U4417 (N_4417,N_2513,N_2985);
or U4418 (N_4418,N_3496,N_3722);
xnor U4419 (N_4419,N_2628,N_3548);
or U4420 (N_4420,N_3605,N_3653);
and U4421 (N_4421,N_3365,N_3718);
or U4422 (N_4422,N_3172,N_2575);
or U4423 (N_4423,N_3360,N_3579);
nor U4424 (N_4424,N_3275,N_2655);
xor U4425 (N_4425,N_3379,N_3142);
and U4426 (N_4426,N_3609,N_2808);
nand U4427 (N_4427,N_3162,N_2763);
nand U4428 (N_4428,N_2948,N_3655);
nand U4429 (N_4429,N_3284,N_2748);
or U4430 (N_4430,N_3719,N_2936);
nor U4431 (N_4431,N_2543,N_3200);
xor U4432 (N_4432,N_3291,N_3597);
nand U4433 (N_4433,N_2728,N_3643);
and U4434 (N_4434,N_3742,N_3719);
xnor U4435 (N_4435,N_3010,N_2566);
or U4436 (N_4436,N_3329,N_3224);
xor U4437 (N_4437,N_3413,N_2594);
xor U4438 (N_4438,N_2649,N_3192);
nor U4439 (N_4439,N_2762,N_2530);
xnor U4440 (N_4440,N_3067,N_3165);
or U4441 (N_4441,N_3284,N_3350);
or U4442 (N_4442,N_3003,N_3075);
and U4443 (N_4443,N_2906,N_2741);
xor U4444 (N_4444,N_3646,N_3246);
xor U4445 (N_4445,N_3451,N_2562);
or U4446 (N_4446,N_2700,N_3548);
nand U4447 (N_4447,N_3614,N_3173);
nor U4448 (N_4448,N_2662,N_2775);
xor U4449 (N_4449,N_2980,N_3150);
xor U4450 (N_4450,N_2861,N_3427);
or U4451 (N_4451,N_3682,N_3158);
nand U4452 (N_4452,N_3090,N_3331);
and U4453 (N_4453,N_3251,N_2811);
nand U4454 (N_4454,N_3116,N_2591);
nand U4455 (N_4455,N_3505,N_3742);
and U4456 (N_4456,N_2932,N_3735);
nand U4457 (N_4457,N_2706,N_3296);
nand U4458 (N_4458,N_3669,N_3423);
xor U4459 (N_4459,N_3419,N_3025);
or U4460 (N_4460,N_3611,N_3297);
nor U4461 (N_4461,N_3380,N_3419);
xnor U4462 (N_4462,N_3230,N_3441);
nor U4463 (N_4463,N_2571,N_2812);
xnor U4464 (N_4464,N_2571,N_2809);
and U4465 (N_4465,N_3031,N_3667);
or U4466 (N_4466,N_2958,N_2846);
nor U4467 (N_4467,N_3082,N_2870);
and U4468 (N_4468,N_2931,N_2678);
nor U4469 (N_4469,N_2509,N_2982);
nand U4470 (N_4470,N_2758,N_2818);
and U4471 (N_4471,N_3351,N_3396);
xor U4472 (N_4472,N_3096,N_3040);
xnor U4473 (N_4473,N_2795,N_2866);
xor U4474 (N_4474,N_3692,N_2540);
or U4475 (N_4475,N_3330,N_2638);
nor U4476 (N_4476,N_3416,N_2578);
nor U4477 (N_4477,N_3121,N_2751);
and U4478 (N_4478,N_2628,N_3520);
nor U4479 (N_4479,N_2510,N_2695);
nand U4480 (N_4480,N_2562,N_3036);
xnor U4481 (N_4481,N_3114,N_2510);
nand U4482 (N_4482,N_2883,N_2625);
or U4483 (N_4483,N_2525,N_2784);
nand U4484 (N_4484,N_3037,N_3583);
or U4485 (N_4485,N_3692,N_2909);
nor U4486 (N_4486,N_3399,N_2519);
nor U4487 (N_4487,N_3161,N_2533);
nor U4488 (N_4488,N_2871,N_3253);
and U4489 (N_4489,N_3681,N_3557);
nor U4490 (N_4490,N_3639,N_3688);
nand U4491 (N_4491,N_2999,N_3027);
nor U4492 (N_4492,N_3510,N_2766);
xor U4493 (N_4493,N_3407,N_2936);
nor U4494 (N_4494,N_2627,N_2908);
or U4495 (N_4495,N_3427,N_3231);
nor U4496 (N_4496,N_3317,N_3140);
or U4497 (N_4497,N_3227,N_2531);
and U4498 (N_4498,N_3197,N_2783);
or U4499 (N_4499,N_3500,N_3624);
xor U4500 (N_4500,N_2677,N_3129);
nor U4501 (N_4501,N_3617,N_3235);
and U4502 (N_4502,N_3241,N_3233);
nor U4503 (N_4503,N_3292,N_3241);
and U4504 (N_4504,N_3729,N_3147);
nor U4505 (N_4505,N_2904,N_3562);
and U4506 (N_4506,N_3618,N_2995);
nand U4507 (N_4507,N_2618,N_3347);
nand U4508 (N_4508,N_3690,N_3541);
xnor U4509 (N_4509,N_3322,N_2883);
and U4510 (N_4510,N_2751,N_3591);
xnor U4511 (N_4511,N_2878,N_3122);
or U4512 (N_4512,N_3635,N_2516);
or U4513 (N_4513,N_3043,N_3188);
xor U4514 (N_4514,N_3141,N_2513);
or U4515 (N_4515,N_2801,N_3594);
nor U4516 (N_4516,N_3157,N_3428);
nand U4517 (N_4517,N_2974,N_3365);
nor U4518 (N_4518,N_2917,N_2975);
xor U4519 (N_4519,N_3076,N_3161);
nand U4520 (N_4520,N_2677,N_2735);
xor U4521 (N_4521,N_3605,N_3679);
nand U4522 (N_4522,N_2558,N_3668);
nor U4523 (N_4523,N_2716,N_3585);
or U4524 (N_4524,N_2848,N_2721);
and U4525 (N_4525,N_2930,N_3307);
nor U4526 (N_4526,N_3560,N_3670);
and U4527 (N_4527,N_3150,N_2566);
and U4528 (N_4528,N_2721,N_2711);
xnor U4529 (N_4529,N_3216,N_3224);
or U4530 (N_4530,N_3636,N_2575);
nor U4531 (N_4531,N_2660,N_2695);
xor U4532 (N_4532,N_3018,N_2801);
and U4533 (N_4533,N_3610,N_3612);
or U4534 (N_4534,N_3682,N_2718);
nor U4535 (N_4535,N_3572,N_3251);
or U4536 (N_4536,N_2642,N_3514);
nor U4537 (N_4537,N_3055,N_3343);
nand U4538 (N_4538,N_3576,N_3039);
and U4539 (N_4539,N_2593,N_3116);
nor U4540 (N_4540,N_3698,N_3053);
nand U4541 (N_4541,N_3565,N_3084);
xnor U4542 (N_4542,N_3492,N_2984);
nor U4543 (N_4543,N_3359,N_3038);
nor U4544 (N_4544,N_3073,N_3149);
nor U4545 (N_4545,N_3014,N_3144);
nand U4546 (N_4546,N_3508,N_3482);
and U4547 (N_4547,N_3414,N_3307);
nor U4548 (N_4548,N_3338,N_3502);
or U4549 (N_4549,N_3074,N_2733);
nor U4550 (N_4550,N_3469,N_2782);
or U4551 (N_4551,N_3183,N_2654);
nand U4552 (N_4552,N_3585,N_3386);
nand U4553 (N_4553,N_3038,N_3087);
and U4554 (N_4554,N_2925,N_3597);
and U4555 (N_4555,N_3648,N_3069);
or U4556 (N_4556,N_3173,N_3295);
xnor U4557 (N_4557,N_3176,N_3529);
nor U4558 (N_4558,N_3514,N_3298);
xnor U4559 (N_4559,N_2826,N_3610);
and U4560 (N_4560,N_2885,N_3147);
or U4561 (N_4561,N_2979,N_2658);
and U4562 (N_4562,N_2682,N_3346);
xor U4563 (N_4563,N_3397,N_3720);
nor U4564 (N_4564,N_2505,N_2661);
nand U4565 (N_4565,N_2712,N_2737);
xnor U4566 (N_4566,N_3741,N_3187);
or U4567 (N_4567,N_3172,N_2656);
xor U4568 (N_4568,N_3702,N_3419);
xnor U4569 (N_4569,N_2853,N_2917);
nand U4570 (N_4570,N_2505,N_2600);
and U4571 (N_4571,N_2650,N_3348);
nor U4572 (N_4572,N_2746,N_3524);
nor U4573 (N_4573,N_3190,N_2858);
nor U4574 (N_4574,N_3672,N_2831);
nor U4575 (N_4575,N_3048,N_3207);
or U4576 (N_4576,N_2754,N_2627);
xnor U4577 (N_4577,N_3523,N_2672);
nand U4578 (N_4578,N_3614,N_2708);
or U4579 (N_4579,N_3610,N_2806);
xnor U4580 (N_4580,N_3725,N_2727);
nor U4581 (N_4581,N_2918,N_2879);
or U4582 (N_4582,N_2922,N_2903);
nand U4583 (N_4583,N_3363,N_2712);
or U4584 (N_4584,N_2752,N_3462);
nor U4585 (N_4585,N_3554,N_3401);
nand U4586 (N_4586,N_3729,N_2817);
xor U4587 (N_4587,N_3481,N_2553);
and U4588 (N_4588,N_2533,N_2735);
xor U4589 (N_4589,N_2714,N_3544);
xnor U4590 (N_4590,N_3467,N_2700);
or U4591 (N_4591,N_3007,N_3100);
or U4592 (N_4592,N_2571,N_3357);
or U4593 (N_4593,N_3231,N_2641);
nand U4594 (N_4594,N_3048,N_3663);
xor U4595 (N_4595,N_2754,N_2865);
xor U4596 (N_4596,N_2618,N_3279);
xor U4597 (N_4597,N_3084,N_3037);
or U4598 (N_4598,N_3523,N_2763);
nor U4599 (N_4599,N_3353,N_3528);
nand U4600 (N_4600,N_3300,N_3079);
and U4601 (N_4601,N_2634,N_2978);
or U4602 (N_4602,N_2768,N_2967);
nor U4603 (N_4603,N_3655,N_2725);
nor U4604 (N_4604,N_3113,N_2862);
and U4605 (N_4605,N_3314,N_3258);
xnor U4606 (N_4606,N_2988,N_3397);
nand U4607 (N_4607,N_3200,N_2856);
and U4608 (N_4608,N_2950,N_3622);
xnor U4609 (N_4609,N_3450,N_2666);
nand U4610 (N_4610,N_3308,N_3239);
and U4611 (N_4611,N_3731,N_3435);
or U4612 (N_4612,N_3608,N_3658);
nor U4613 (N_4613,N_2620,N_2978);
and U4614 (N_4614,N_2852,N_3070);
xnor U4615 (N_4615,N_2791,N_3167);
or U4616 (N_4616,N_3714,N_2798);
or U4617 (N_4617,N_3026,N_3124);
nor U4618 (N_4618,N_3042,N_3724);
or U4619 (N_4619,N_2889,N_3449);
nand U4620 (N_4620,N_3348,N_3242);
and U4621 (N_4621,N_3540,N_2699);
or U4622 (N_4622,N_3066,N_2865);
nand U4623 (N_4623,N_3313,N_3320);
xnor U4624 (N_4624,N_3637,N_3028);
nor U4625 (N_4625,N_3005,N_3007);
or U4626 (N_4626,N_2817,N_2885);
nand U4627 (N_4627,N_3107,N_3410);
nand U4628 (N_4628,N_3360,N_2813);
xor U4629 (N_4629,N_2783,N_2977);
nor U4630 (N_4630,N_2838,N_2947);
and U4631 (N_4631,N_2638,N_2790);
xor U4632 (N_4632,N_2792,N_2740);
xor U4633 (N_4633,N_3737,N_2760);
xnor U4634 (N_4634,N_2974,N_2842);
and U4635 (N_4635,N_3061,N_3491);
or U4636 (N_4636,N_3110,N_3065);
or U4637 (N_4637,N_2956,N_2595);
xor U4638 (N_4638,N_3215,N_2840);
nand U4639 (N_4639,N_3200,N_3387);
or U4640 (N_4640,N_2816,N_3265);
nand U4641 (N_4641,N_3174,N_2500);
and U4642 (N_4642,N_2657,N_3336);
nand U4643 (N_4643,N_3196,N_3722);
nand U4644 (N_4644,N_3723,N_3466);
xnor U4645 (N_4645,N_2740,N_3050);
or U4646 (N_4646,N_3517,N_3749);
nand U4647 (N_4647,N_3296,N_2738);
or U4648 (N_4648,N_3509,N_2574);
xnor U4649 (N_4649,N_3530,N_3475);
nand U4650 (N_4650,N_3697,N_3593);
xnor U4651 (N_4651,N_2590,N_3721);
xnor U4652 (N_4652,N_2834,N_3358);
or U4653 (N_4653,N_3373,N_3447);
or U4654 (N_4654,N_3341,N_3302);
nand U4655 (N_4655,N_3528,N_3697);
nand U4656 (N_4656,N_3004,N_3334);
and U4657 (N_4657,N_2992,N_2838);
and U4658 (N_4658,N_3592,N_3234);
xnor U4659 (N_4659,N_3200,N_2608);
and U4660 (N_4660,N_3206,N_2549);
nor U4661 (N_4661,N_3081,N_3184);
nand U4662 (N_4662,N_2759,N_3104);
nand U4663 (N_4663,N_3016,N_3245);
and U4664 (N_4664,N_2633,N_2986);
or U4665 (N_4665,N_2523,N_3714);
and U4666 (N_4666,N_3172,N_2823);
xor U4667 (N_4667,N_3233,N_3727);
and U4668 (N_4668,N_2838,N_2602);
nand U4669 (N_4669,N_2920,N_3003);
or U4670 (N_4670,N_3606,N_3031);
nand U4671 (N_4671,N_3714,N_2968);
xnor U4672 (N_4672,N_2748,N_3371);
nor U4673 (N_4673,N_2749,N_3564);
nor U4674 (N_4674,N_2819,N_2519);
nand U4675 (N_4675,N_3603,N_3049);
xnor U4676 (N_4676,N_3411,N_2693);
or U4677 (N_4677,N_3408,N_2907);
and U4678 (N_4678,N_3296,N_3131);
xnor U4679 (N_4679,N_3733,N_3331);
xor U4680 (N_4680,N_3472,N_2569);
and U4681 (N_4681,N_3658,N_3505);
xor U4682 (N_4682,N_3232,N_3389);
nand U4683 (N_4683,N_2946,N_3622);
nand U4684 (N_4684,N_3296,N_3034);
nor U4685 (N_4685,N_3721,N_3691);
nand U4686 (N_4686,N_3189,N_2666);
or U4687 (N_4687,N_3334,N_2661);
xor U4688 (N_4688,N_3124,N_3156);
or U4689 (N_4689,N_2508,N_3122);
or U4690 (N_4690,N_3236,N_3377);
and U4691 (N_4691,N_3112,N_3208);
xnor U4692 (N_4692,N_2697,N_3233);
nor U4693 (N_4693,N_3338,N_3400);
nor U4694 (N_4694,N_2939,N_3320);
or U4695 (N_4695,N_2832,N_3159);
nand U4696 (N_4696,N_3532,N_2716);
xor U4697 (N_4697,N_2925,N_3359);
and U4698 (N_4698,N_3194,N_3519);
nor U4699 (N_4699,N_3326,N_3137);
nand U4700 (N_4700,N_3261,N_3078);
nand U4701 (N_4701,N_2527,N_3374);
nand U4702 (N_4702,N_3121,N_3533);
xor U4703 (N_4703,N_2884,N_2726);
or U4704 (N_4704,N_2516,N_2860);
nor U4705 (N_4705,N_3155,N_3598);
xor U4706 (N_4706,N_3369,N_3065);
xnor U4707 (N_4707,N_2658,N_3546);
nand U4708 (N_4708,N_3123,N_3713);
nand U4709 (N_4709,N_2726,N_3541);
and U4710 (N_4710,N_3261,N_3339);
nor U4711 (N_4711,N_3005,N_3575);
or U4712 (N_4712,N_3073,N_2795);
xnor U4713 (N_4713,N_2755,N_2748);
nor U4714 (N_4714,N_3321,N_3094);
or U4715 (N_4715,N_3293,N_2518);
nor U4716 (N_4716,N_2980,N_2659);
or U4717 (N_4717,N_2955,N_2502);
nand U4718 (N_4718,N_3095,N_2580);
and U4719 (N_4719,N_3442,N_2617);
and U4720 (N_4720,N_3093,N_3703);
xnor U4721 (N_4721,N_2558,N_2737);
xor U4722 (N_4722,N_3157,N_3188);
and U4723 (N_4723,N_3287,N_3541);
xnor U4724 (N_4724,N_2951,N_3743);
or U4725 (N_4725,N_2641,N_3167);
xnor U4726 (N_4726,N_3343,N_3050);
nand U4727 (N_4727,N_2529,N_3585);
nand U4728 (N_4728,N_2789,N_2640);
nand U4729 (N_4729,N_3169,N_3170);
nor U4730 (N_4730,N_2975,N_3171);
nor U4731 (N_4731,N_3153,N_2856);
and U4732 (N_4732,N_3188,N_3417);
and U4733 (N_4733,N_2541,N_3495);
nor U4734 (N_4734,N_3234,N_3091);
xnor U4735 (N_4735,N_2742,N_3641);
nand U4736 (N_4736,N_3380,N_3548);
xor U4737 (N_4737,N_3530,N_2744);
nor U4738 (N_4738,N_3393,N_3159);
xor U4739 (N_4739,N_3668,N_2537);
or U4740 (N_4740,N_3170,N_2985);
and U4741 (N_4741,N_2762,N_3265);
xor U4742 (N_4742,N_3242,N_2950);
xor U4743 (N_4743,N_3370,N_2809);
xor U4744 (N_4744,N_3447,N_3076);
or U4745 (N_4745,N_2664,N_3528);
and U4746 (N_4746,N_3248,N_3586);
nand U4747 (N_4747,N_2726,N_3606);
and U4748 (N_4748,N_2563,N_3704);
nand U4749 (N_4749,N_2732,N_3230);
nor U4750 (N_4750,N_2913,N_3473);
or U4751 (N_4751,N_2577,N_3268);
and U4752 (N_4752,N_2856,N_3096);
and U4753 (N_4753,N_3505,N_2552);
and U4754 (N_4754,N_3426,N_3374);
or U4755 (N_4755,N_3283,N_2636);
nor U4756 (N_4756,N_3020,N_3402);
xnor U4757 (N_4757,N_3374,N_3608);
nor U4758 (N_4758,N_3422,N_3179);
xor U4759 (N_4759,N_3658,N_3556);
nor U4760 (N_4760,N_2613,N_3143);
xor U4761 (N_4761,N_3688,N_3310);
or U4762 (N_4762,N_3501,N_3338);
and U4763 (N_4763,N_2986,N_3311);
nand U4764 (N_4764,N_3034,N_2625);
nand U4765 (N_4765,N_3195,N_3516);
xnor U4766 (N_4766,N_3236,N_3213);
nor U4767 (N_4767,N_3589,N_2838);
or U4768 (N_4768,N_3225,N_3140);
nor U4769 (N_4769,N_3373,N_2737);
and U4770 (N_4770,N_3543,N_2820);
nand U4771 (N_4771,N_3106,N_2876);
or U4772 (N_4772,N_2728,N_3640);
nor U4773 (N_4773,N_3233,N_3109);
nand U4774 (N_4774,N_2530,N_3332);
or U4775 (N_4775,N_2924,N_2862);
nor U4776 (N_4776,N_2869,N_3506);
nor U4777 (N_4777,N_2538,N_2558);
nor U4778 (N_4778,N_2568,N_3620);
or U4779 (N_4779,N_3163,N_3404);
nor U4780 (N_4780,N_2992,N_2991);
and U4781 (N_4781,N_2964,N_3710);
or U4782 (N_4782,N_3308,N_3557);
or U4783 (N_4783,N_3222,N_3440);
and U4784 (N_4784,N_2529,N_2844);
nor U4785 (N_4785,N_2516,N_2850);
or U4786 (N_4786,N_3612,N_2718);
nand U4787 (N_4787,N_2750,N_3671);
or U4788 (N_4788,N_3658,N_3309);
nor U4789 (N_4789,N_3243,N_2867);
xnor U4790 (N_4790,N_3316,N_3325);
nor U4791 (N_4791,N_2774,N_2608);
nor U4792 (N_4792,N_2681,N_3272);
nand U4793 (N_4793,N_3495,N_3426);
nand U4794 (N_4794,N_2926,N_3539);
or U4795 (N_4795,N_2555,N_3151);
nand U4796 (N_4796,N_3071,N_2883);
and U4797 (N_4797,N_2728,N_3715);
or U4798 (N_4798,N_3625,N_3250);
xor U4799 (N_4799,N_3189,N_2619);
xnor U4800 (N_4800,N_2867,N_2681);
xor U4801 (N_4801,N_3003,N_2911);
nand U4802 (N_4802,N_2599,N_3461);
nor U4803 (N_4803,N_2701,N_2511);
xnor U4804 (N_4804,N_2504,N_2517);
and U4805 (N_4805,N_2600,N_2995);
or U4806 (N_4806,N_2917,N_3524);
xnor U4807 (N_4807,N_3719,N_3187);
or U4808 (N_4808,N_2572,N_2949);
xnor U4809 (N_4809,N_3522,N_2907);
xor U4810 (N_4810,N_2654,N_2640);
nor U4811 (N_4811,N_3693,N_3652);
xnor U4812 (N_4812,N_3700,N_2938);
or U4813 (N_4813,N_2617,N_3534);
xnor U4814 (N_4814,N_2932,N_2815);
and U4815 (N_4815,N_2996,N_3304);
nand U4816 (N_4816,N_3368,N_3537);
and U4817 (N_4817,N_3220,N_3100);
nand U4818 (N_4818,N_3440,N_3362);
nand U4819 (N_4819,N_3533,N_3614);
or U4820 (N_4820,N_3416,N_3298);
nor U4821 (N_4821,N_2733,N_2546);
or U4822 (N_4822,N_2836,N_2628);
and U4823 (N_4823,N_3335,N_3357);
nor U4824 (N_4824,N_3017,N_2979);
and U4825 (N_4825,N_3617,N_3285);
xnor U4826 (N_4826,N_3257,N_3156);
nor U4827 (N_4827,N_2875,N_3294);
xor U4828 (N_4828,N_2905,N_3407);
nor U4829 (N_4829,N_3051,N_3155);
xnor U4830 (N_4830,N_3197,N_3688);
nor U4831 (N_4831,N_3443,N_2751);
nand U4832 (N_4832,N_2540,N_3368);
nand U4833 (N_4833,N_3210,N_3611);
nand U4834 (N_4834,N_3361,N_3584);
and U4835 (N_4835,N_3194,N_2957);
nor U4836 (N_4836,N_3334,N_3376);
or U4837 (N_4837,N_2539,N_3687);
xnor U4838 (N_4838,N_2838,N_3463);
nand U4839 (N_4839,N_2570,N_3727);
nor U4840 (N_4840,N_3524,N_3369);
nor U4841 (N_4841,N_3127,N_3227);
and U4842 (N_4842,N_3647,N_3734);
and U4843 (N_4843,N_2881,N_2628);
xnor U4844 (N_4844,N_3301,N_3199);
nand U4845 (N_4845,N_3242,N_2721);
xor U4846 (N_4846,N_2803,N_3476);
or U4847 (N_4847,N_3625,N_2667);
xor U4848 (N_4848,N_3422,N_3162);
nor U4849 (N_4849,N_3368,N_2563);
xnor U4850 (N_4850,N_3283,N_3693);
nand U4851 (N_4851,N_3003,N_3535);
and U4852 (N_4852,N_3525,N_3254);
xnor U4853 (N_4853,N_3190,N_3184);
and U4854 (N_4854,N_3268,N_3677);
or U4855 (N_4855,N_3674,N_2799);
nor U4856 (N_4856,N_3198,N_2915);
nor U4857 (N_4857,N_3427,N_3060);
nand U4858 (N_4858,N_3000,N_3580);
nor U4859 (N_4859,N_3598,N_3617);
nor U4860 (N_4860,N_3495,N_3346);
and U4861 (N_4861,N_3519,N_2591);
nor U4862 (N_4862,N_3729,N_3667);
and U4863 (N_4863,N_3695,N_3433);
or U4864 (N_4864,N_2651,N_2984);
nand U4865 (N_4865,N_2687,N_2700);
and U4866 (N_4866,N_3267,N_2681);
nand U4867 (N_4867,N_3063,N_2779);
xor U4868 (N_4868,N_2747,N_2862);
nand U4869 (N_4869,N_3392,N_3520);
nand U4870 (N_4870,N_2867,N_2538);
nor U4871 (N_4871,N_3457,N_3506);
xnor U4872 (N_4872,N_3625,N_2609);
and U4873 (N_4873,N_3115,N_3207);
nand U4874 (N_4874,N_3103,N_3386);
and U4875 (N_4875,N_2529,N_3710);
nor U4876 (N_4876,N_3102,N_3206);
xor U4877 (N_4877,N_3566,N_2792);
and U4878 (N_4878,N_3710,N_3732);
xnor U4879 (N_4879,N_3350,N_3244);
or U4880 (N_4880,N_3154,N_3353);
and U4881 (N_4881,N_3538,N_3516);
and U4882 (N_4882,N_3555,N_3371);
xor U4883 (N_4883,N_2698,N_3541);
or U4884 (N_4884,N_3089,N_3144);
or U4885 (N_4885,N_2809,N_2928);
or U4886 (N_4886,N_2999,N_2592);
nand U4887 (N_4887,N_3694,N_3402);
or U4888 (N_4888,N_2507,N_3493);
or U4889 (N_4889,N_2797,N_3580);
xor U4890 (N_4890,N_2565,N_3578);
or U4891 (N_4891,N_2592,N_3314);
nor U4892 (N_4892,N_2748,N_3181);
nand U4893 (N_4893,N_2834,N_2843);
and U4894 (N_4894,N_3158,N_3037);
nand U4895 (N_4895,N_2885,N_3669);
nor U4896 (N_4896,N_2935,N_3151);
nor U4897 (N_4897,N_3544,N_3404);
nand U4898 (N_4898,N_3250,N_3515);
nor U4899 (N_4899,N_2898,N_3510);
xnor U4900 (N_4900,N_2859,N_2755);
or U4901 (N_4901,N_2864,N_3174);
nor U4902 (N_4902,N_2868,N_3414);
nor U4903 (N_4903,N_2665,N_2633);
or U4904 (N_4904,N_2685,N_2551);
or U4905 (N_4905,N_2901,N_3747);
xnor U4906 (N_4906,N_3745,N_3529);
nor U4907 (N_4907,N_3313,N_2612);
xor U4908 (N_4908,N_2785,N_3095);
or U4909 (N_4909,N_3016,N_3134);
nand U4910 (N_4910,N_2917,N_2519);
xnor U4911 (N_4911,N_2566,N_3359);
xnor U4912 (N_4912,N_3703,N_3235);
xnor U4913 (N_4913,N_3247,N_3043);
xnor U4914 (N_4914,N_3206,N_3115);
nor U4915 (N_4915,N_3599,N_3036);
xor U4916 (N_4916,N_2675,N_3070);
or U4917 (N_4917,N_3552,N_3421);
and U4918 (N_4918,N_3600,N_2587);
xnor U4919 (N_4919,N_2668,N_3633);
nor U4920 (N_4920,N_3111,N_3194);
xor U4921 (N_4921,N_2937,N_2864);
or U4922 (N_4922,N_2999,N_3168);
nand U4923 (N_4923,N_3172,N_3748);
nand U4924 (N_4924,N_3642,N_3001);
and U4925 (N_4925,N_2508,N_3679);
xor U4926 (N_4926,N_2568,N_2793);
xor U4927 (N_4927,N_3047,N_2599);
xor U4928 (N_4928,N_2724,N_3561);
nor U4929 (N_4929,N_2855,N_2858);
nor U4930 (N_4930,N_2594,N_2610);
nor U4931 (N_4931,N_3357,N_3504);
nor U4932 (N_4932,N_3436,N_3215);
and U4933 (N_4933,N_2576,N_2867);
nand U4934 (N_4934,N_3032,N_2520);
nor U4935 (N_4935,N_2978,N_3227);
nand U4936 (N_4936,N_2715,N_2703);
nand U4937 (N_4937,N_3626,N_3354);
xor U4938 (N_4938,N_3567,N_3350);
xor U4939 (N_4939,N_3373,N_2820);
and U4940 (N_4940,N_2540,N_3385);
or U4941 (N_4941,N_3199,N_3612);
nand U4942 (N_4942,N_3556,N_2964);
nor U4943 (N_4943,N_2898,N_3651);
or U4944 (N_4944,N_3222,N_3392);
xnor U4945 (N_4945,N_3558,N_3306);
xor U4946 (N_4946,N_3147,N_3437);
xnor U4947 (N_4947,N_3433,N_2695);
nor U4948 (N_4948,N_3342,N_2721);
or U4949 (N_4949,N_3529,N_3682);
nor U4950 (N_4950,N_3178,N_3174);
and U4951 (N_4951,N_3477,N_3293);
or U4952 (N_4952,N_3564,N_2962);
and U4953 (N_4953,N_2582,N_3434);
and U4954 (N_4954,N_2893,N_3007);
or U4955 (N_4955,N_2709,N_3190);
nor U4956 (N_4956,N_3605,N_3254);
and U4957 (N_4957,N_2537,N_3525);
and U4958 (N_4958,N_3564,N_3251);
and U4959 (N_4959,N_3064,N_2587);
xnor U4960 (N_4960,N_2529,N_3110);
and U4961 (N_4961,N_2791,N_2533);
and U4962 (N_4962,N_2820,N_2536);
or U4963 (N_4963,N_2814,N_2533);
and U4964 (N_4964,N_3424,N_3277);
or U4965 (N_4965,N_3474,N_2506);
xor U4966 (N_4966,N_2537,N_3413);
nor U4967 (N_4967,N_3187,N_3066);
xnor U4968 (N_4968,N_3509,N_3096);
and U4969 (N_4969,N_3485,N_2547);
xor U4970 (N_4970,N_3180,N_3488);
nand U4971 (N_4971,N_3662,N_3489);
and U4972 (N_4972,N_3454,N_2669);
and U4973 (N_4973,N_2800,N_3537);
nor U4974 (N_4974,N_3171,N_3161);
or U4975 (N_4975,N_3620,N_2545);
and U4976 (N_4976,N_3308,N_3690);
nand U4977 (N_4977,N_3167,N_3341);
xnor U4978 (N_4978,N_2500,N_3327);
nor U4979 (N_4979,N_2680,N_2819);
xnor U4980 (N_4980,N_3021,N_2580);
nor U4981 (N_4981,N_3017,N_2761);
nand U4982 (N_4982,N_3496,N_3594);
nand U4983 (N_4983,N_2516,N_2947);
xnor U4984 (N_4984,N_3207,N_3598);
and U4985 (N_4985,N_3735,N_2912);
xnor U4986 (N_4986,N_3179,N_3492);
nand U4987 (N_4987,N_2829,N_2985);
nand U4988 (N_4988,N_2741,N_3506);
nand U4989 (N_4989,N_3655,N_2524);
and U4990 (N_4990,N_3659,N_3623);
nor U4991 (N_4991,N_2576,N_3693);
nand U4992 (N_4992,N_2780,N_3517);
nor U4993 (N_4993,N_3342,N_3723);
nand U4994 (N_4994,N_2836,N_2809);
xnor U4995 (N_4995,N_3237,N_2882);
nor U4996 (N_4996,N_2738,N_3202);
nor U4997 (N_4997,N_2866,N_2703);
nor U4998 (N_4998,N_2939,N_3692);
or U4999 (N_4999,N_2819,N_3388);
xor U5000 (N_5000,N_4029,N_3821);
xor U5001 (N_5001,N_4848,N_4605);
xnor U5002 (N_5002,N_4425,N_4583);
nand U5003 (N_5003,N_4638,N_4150);
nor U5004 (N_5004,N_4538,N_4164);
xnor U5005 (N_5005,N_4646,N_3929);
nor U5006 (N_5006,N_4759,N_4714);
or U5007 (N_5007,N_3818,N_4544);
nor U5008 (N_5008,N_4828,N_4230);
or U5009 (N_5009,N_3993,N_4069);
nor U5010 (N_5010,N_4672,N_4701);
nor U5011 (N_5011,N_4811,N_4500);
xor U5012 (N_5012,N_4876,N_4224);
and U5013 (N_5013,N_4409,N_4878);
or U5014 (N_5014,N_4383,N_4089);
xnor U5015 (N_5015,N_3908,N_4915);
nor U5016 (N_5016,N_4123,N_4570);
nor U5017 (N_5017,N_3927,N_3878);
and U5018 (N_5018,N_4242,N_4100);
or U5019 (N_5019,N_4328,N_4971);
xnor U5020 (N_5020,N_4795,N_4613);
and U5021 (N_5021,N_4340,N_4929);
nand U5022 (N_5022,N_4703,N_4105);
and U5023 (N_5023,N_4159,N_3970);
xnor U5024 (N_5024,N_3763,N_4593);
xnor U5025 (N_5025,N_4639,N_4839);
or U5026 (N_5026,N_3989,N_4663);
and U5027 (N_5027,N_3795,N_3883);
and U5028 (N_5028,N_4477,N_4749);
nand U5029 (N_5029,N_4531,N_4245);
xor U5030 (N_5030,N_3897,N_3779);
xnor U5031 (N_5031,N_4888,N_4945);
nand U5032 (N_5032,N_3930,N_4832);
xnor U5033 (N_5033,N_4063,N_4191);
nor U5034 (N_5034,N_4794,N_3774);
nor U5035 (N_5035,N_4960,N_3754);
nand U5036 (N_5036,N_4038,N_4655);
and U5037 (N_5037,N_3903,N_4112);
xnor U5038 (N_5038,N_4446,N_4621);
nand U5039 (N_5039,N_4428,N_4412);
and U5040 (N_5040,N_4943,N_4420);
nor U5041 (N_5041,N_4536,N_4445);
nand U5042 (N_5042,N_4900,N_3856);
nor U5043 (N_5043,N_4724,N_4156);
xor U5044 (N_5044,N_4297,N_4339);
or U5045 (N_5045,N_4979,N_4028);
nand U5046 (N_5046,N_4232,N_4264);
xor U5047 (N_5047,N_3782,N_4567);
and U5048 (N_5048,N_4873,N_4343);
nor U5049 (N_5049,N_4585,N_4345);
nor U5050 (N_5050,N_3750,N_4935);
nor U5051 (N_5051,N_4278,N_3951);
xnor U5052 (N_5052,N_4248,N_4186);
nand U5053 (N_5053,N_4001,N_4424);
nor U5054 (N_5054,N_4463,N_4306);
and U5055 (N_5055,N_4141,N_4901);
nand U5056 (N_5056,N_3974,N_4921);
nand U5057 (N_5057,N_4511,N_4842);
nand U5058 (N_5058,N_3952,N_4664);
nand U5059 (N_5059,N_4059,N_4775);
nor U5060 (N_5060,N_3934,N_3855);
or U5061 (N_5061,N_4235,N_4279);
nor U5062 (N_5062,N_4195,N_4354);
xor U5063 (N_5063,N_4801,N_3937);
nor U5064 (N_5064,N_4421,N_4524);
nand U5065 (N_5065,N_4007,N_4754);
xnor U5066 (N_5066,N_4146,N_4498);
nand U5067 (N_5067,N_4892,N_3914);
and U5068 (N_5068,N_4198,N_4697);
nand U5069 (N_5069,N_3881,N_4725);
xnor U5070 (N_5070,N_3938,N_4514);
and U5071 (N_5071,N_4379,N_3815);
or U5072 (N_5072,N_4018,N_3838);
nand U5073 (N_5073,N_4416,N_4782);
xnor U5074 (N_5074,N_4133,N_3783);
or U5075 (N_5075,N_4101,N_3979);
nor U5076 (N_5076,N_4118,N_4912);
and U5077 (N_5077,N_4678,N_3862);
nand U5078 (N_5078,N_4776,N_3891);
nor U5079 (N_5079,N_3922,N_3955);
xor U5080 (N_5080,N_4800,N_3845);
nand U5081 (N_5081,N_4826,N_4317);
nor U5082 (N_5082,N_4721,N_4061);
and U5083 (N_5083,N_4978,N_4617);
or U5084 (N_5084,N_4153,N_4868);
nand U5085 (N_5085,N_3960,N_4924);
nand U5086 (N_5086,N_4373,N_4351);
xnor U5087 (N_5087,N_4809,N_3958);
nand U5088 (N_5088,N_4958,N_4523);
nor U5089 (N_5089,N_4481,N_3947);
or U5090 (N_5090,N_4253,N_4624);
nand U5091 (N_5091,N_4115,N_4913);
nor U5092 (N_5092,N_4905,N_4108);
xor U5093 (N_5093,N_4649,N_4837);
or U5094 (N_5094,N_4576,N_4925);
and U5095 (N_5095,N_3765,N_4393);
nor U5096 (N_5096,N_4472,N_4067);
and U5097 (N_5097,N_4094,N_4685);
nor U5098 (N_5098,N_3785,N_4142);
nor U5099 (N_5099,N_4331,N_4267);
and U5100 (N_5100,N_4933,N_4045);
nor U5101 (N_5101,N_4798,N_3893);
and U5102 (N_5102,N_4777,N_4289);
nand U5103 (N_5103,N_4489,N_4551);
nor U5104 (N_5104,N_4200,N_3842);
xor U5105 (N_5105,N_4429,N_4990);
and U5106 (N_5106,N_4037,N_4993);
or U5107 (N_5107,N_4590,N_4095);
and U5108 (N_5108,N_4450,N_4569);
nand U5109 (N_5109,N_3847,N_4326);
xnor U5110 (N_5110,N_4715,N_4601);
and U5111 (N_5111,N_4092,N_4308);
and U5112 (N_5112,N_4930,N_4881);
nand U5113 (N_5113,N_4952,N_4185);
nor U5114 (N_5114,N_4290,N_3953);
or U5115 (N_5115,N_4596,N_4134);
xnor U5116 (N_5116,N_4020,N_4342);
nand U5117 (N_5117,N_3778,N_4987);
or U5118 (N_5118,N_3997,N_4507);
and U5119 (N_5119,N_3840,N_4581);
nor U5120 (N_5120,N_4997,N_4772);
xnor U5121 (N_5121,N_4559,N_4967);
nor U5122 (N_5122,N_4882,N_4937);
nand U5123 (N_5123,N_4822,N_4447);
nor U5124 (N_5124,N_3852,N_4865);
xor U5125 (N_5125,N_3931,N_3836);
nor U5126 (N_5126,N_4275,N_3933);
or U5127 (N_5127,N_3844,N_4367);
and U5128 (N_5128,N_4918,N_3764);
xnor U5129 (N_5129,N_4385,N_4456);
and U5130 (N_5130,N_3851,N_4615);
xor U5131 (N_5131,N_4680,N_4517);
and U5132 (N_5132,N_4293,N_3888);
nor U5133 (N_5133,N_4418,N_4009);
nand U5134 (N_5134,N_3944,N_4064);
and U5135 (N_5135,N_4212,N_4144);
nand U5136 (N_5136,N_4135,N_4914);
xor U5137 (N_5137,N_4642,N_4969);
nor U5138 (N_5138,N_4690,N_4155);
xnor U5139 (N_5139,N_4422,N_4553);
xor U5140 (N_5140,N_4196,N_4610);
nand U5141 (N_5141,N_4575,N_4874);
xnor U5142 (N_5142,N_4047,N_3866);
nand U5143 (N_5143,N_4183,N_3793);
or U5144 (N_5144,N_4369,N_4039);
or U5145 (N_5145,N_3973,N_4437);
nor U5146 (N_5146,N_3825,N_3936);
or U5147 (N_5147,N_3971,N_4512);
nor U5148 (N_5148,N_4558,N_4072);
nor U5149 (N_5149,N_4903,N_3757);
or U5150 (N_5150,N_4928,N_4194);
nand U5151 (N_5151,N_4075,N_4883);
nand U5152 (N_5152,N_3926,N_4533);
and U5153 (N_5153,N_4923,N_4199);
or U5154 (N_5154,N_4658,N_4390);
and U5155 (N_5155,N_4495,N_4218);
nor U5156 (N_5156,N_4549,N_3808);
or U5157 (N_5157,N_4854,N_4484);
or U5158 (N_5158,N_4864,N_4675);
nand U5159 (N_5159,N_4268,N_3776);
and U5160 (N_5160,N_4215,N_4619);
or U5161 (N_5161,N_3849,N_4137);
and U5162 (N_5162,N_4830,N_4124);
nand U5163 (N_5163,N_4051,N_4845);
and U5164 (N_5164,N_3963,N_4886);
and U5165 (N_5165,N_4666,N_4143);
and U5166 (N_5166,N_4396,N_4490);
or U5167 (N_5167,N_4614,N_4788);
nand U5168 (N_5168,N_4950,N_4626);
nor U5169 (N_5169,N_4019,N_4050);
nand U5170 (N_5170,N_4181,N_4085);
xor U5171 (N_5171,N_4850,N_3804);
xor U5172 (N_5172,N_4184,N_4947);
or U5173 (N_5173,N_3874,N_4258);
and U5174 (N_5174,N_4313,N_4844);
or U5175 (N_5175,N_3915,N_4126);
nor U5176 (N_5176,N_4255,N_4648);
or U5177 (N_5177,N_4399,N_3964);
and U5178 (N_5178,N_4073,N_4131);
nor U5179 (N_5179,N_3880,N_4766);
or U5180 (N_5180,N_4595,N_4470);
nor U5181 (N_5181,N_4748,N_3811);
nor U5182 (N_5182,N_4168,N_4352);
and U5183 (N_5183,N_3819,N_4249);
and U5184 (N_5184,N_4834,N_3954);
and U5185 (N_5185,N_3853,N_4309);
or U5186 (N_5186,N_4426,N_4008);
nand U5187 (N_5187,N_4751,N_4350);
xor U5188 (N_5188,N_4014,N_3787);
or U5189 (N_5189,N_4079,N_4908);
nor U5190 (N_5190,N_4529,N_4154);
and U5191 (N_5191,N_4157,N_3900);
and U5192 (N_5192,N_4525,N_4985);
or U5193 (N_5193,N_4962,N_4315);
xor U5194 (N_5194,N_4836,N_4314);
nor U5195 (N_5195,N_4843,N_4359);
and U5196 (N_5196,N_4756,N_3932);
or U5197 (N_5197,N_4656,N_4467);
nand U5198 (N_5198,N_3906,N_4841);
nor U5199 (N_5199,N_4374,N_4734);
nand U5200 (N_5200,N_3886,N_4474);
or U5201 (N_5201,N_3940,N_4528);
or U5202 (N_5202,N_4120,N_4025);
or U5203 (N_5203,N_4884,N_4210);
xnor U5204 (N_5204,N_4068,N_3758);
nor U5205 (N_5205,N_3755,N_4922);
and U5206 (N_5206,N_4849,N_4452);
nor U5207 (N_5207,N_4145,N_3983);
or U5208 (N_5208,N_4032,N_4438);
and U5209 (N_5209,N_4002,N_4332);
nor U5210 (N_5210,N_4860,N_3846);
xnor U5211 (N_5211,N_4622,N_4139);
xnor U5212 (N_5212,N_4125,N_4407);
nand U5213 (N_5213,N_4493,N_3981);
xnor U5214 (N_5214,N_4080,N_4877);
or U5215 (N_5215,N_4335,N_4228);
or U5216 (N_5216,N_3773,N_4793);
nor U5217 (N_5217,N_4743,N_4503);
xor U5218 (N_5218,N_4562,N_4401);
nand U5219 (N_5219,N_4982,N_4941);
and U5220 (N_5220,N_4720,N_4270);
and U5221 (N_5221,N_4440,N_3820);
and U5222 (N_5222,N_4833,N_4682);
and U5223 (N_5223,N_4329,N_4377);
nand U5224 (N_5224,N_4885,N_4838);
xnor U5225 (N_5225,N_4643,N_4341);
nor U5226 (N_5226,N_4592,N_4178);
nor U5227 (N_5227,N_4276,N_4594);
or U5228 (N_5228,N_3797,N_4226);
nor U5229 (N_5229,N_4879,N_4565);
nor U5230 (N_5230,N_4630,N_4203);
nand U5231 (N_5231,N_4414,N_4735);
nor U5232 (N_5232,N_4781,N_4482);
and U5233 (N_5233,N_4227,N_3884);
or U5234 (N_5234,N_3885,N_4867);
nand U5235 (N_5235,N_4010,N_4955);
or U5236 (N_5236,N_4820,N_4504);
nor U5237 (N_5237,N_3943,N_4205);
and U5238 (N_5238,N_3859,N_4322);
and U5239 (N_5239,N_4024,N_4087);
or U5240 (N_5240,N_4677,N_4713);
xor U5241 (N_5241,N_4805,N_4448);
or U5242 (N_5242,N_4034,N_4102);
xor U5243 (N_5243,N_4780,N_4855);
or U5244 (N_5244,N_4628,N_4556);
nand U5245 (N_5245,N_4706,N_4093);
and U5246 (N_5246,N_3772,N_4380);
xnor U5247 (N_5247,N_4975,N_3871);
or U5248 (N_5248,N_4505,N_3796);
and U5249 (N_5249,N_3876,N_4816);
or U5250 (N_5250,N_3999,N_4548);
xnor U5251 (N_5251,N_4304,N_4866);
nand U5252 (N_5252,N_4497,N_4693);
nor U5253 (N_5253,N_4113,N_4944);
xor U5254 (N_5254,N_4716,N_4634);
or U5255 (N_5255,N_4111,N_4213);
and U5256 (N_5256,N_3869,N_4819);
and U5257 (N_5257,N_4174,N_3830);
nor U5258 (N_5258,N_4904,N_4081);
nor U5259 (N_5259,N_4598,N_4449);
or U5260 (N_5260,N_4737,N_4861);
xor U5261 (N_5261,N_4998,N_4209);
nor U5262 (N_5262,N_4708,N_4689);
nor U5263 (N_5263,N_4763,N_4220);
nor U5264 (N_5264,N_3972,N_4208);
or U5265 (N_5265,N_4166,N_4435);
and U5266 (N_5266,N_4451,N_4729);
or U5267 (N_5267,N_4269,N_4964);
nor U5268 (N_5268,N_4023,N_3872);
nor U5269 (N_5269,N_4618,N_4831);
xnor U5270 (N_5270,N_4056,N_4821);
xnor U5271 (N_5271,N_4983,N_4476);
or U5272 (N_5272,N_4288,N_4015);
or U5273 (N_5273,N_4283,N_3810);
and U5274 (N_5274,N_4543,N_3998);
xor U5275 (N_5275,N_4600,N_4717);
or U5276 (N_5276,N_4263,N_3913);
nor U5277 (N_5277,N_4004,N_3889);
or U5278 (N_5278,N_4325,N_4286);
xor U5279 (N_5279,N_4176,N_4773);
and U5280 (N_5280,N_3780,N_4035);
nor U5281 (N_5281,N_4302,N_4303);
xnor U5282 (N_5282,N_4177,N_3994);
nand U5283 (N_5283,N_4358,N_4494);
xor U5284 (N_5284,N_4732,N_4243);
nor U5285 (N_5285,N_4650,N_4254);
or U5286 (N_5286,N_4956,N_3831);
nor U5287 (N_5287,N_4563,N_4858);
nor U5288 (N_5288,N_4285,N_4250);
xor U5289 (N_5289,N_4132,N_4239);
or U5290 (N_5290,N_4058,N_4271);
nand U5291 (N_5291,N_4740,N_4457);
xor U5292 (N_5292,N_4674,N_4665);
xnor U5293 (N_5293,N_4934,N_3865);
or U5294 (N_5294,N_4316,N_4392);
or U5295 (N_5295,N_4916,N_4103);
nor U5296 (N_5296,N_4608,N_3801);
or U5297 (N_5297,N_4728,N_4106);
or U5298 (N_5298,N_3867,N_3752);
nor U5299 (N_5299,N_4217,N_3833);
and U5300 (N_5300,N_4152,N_4588);
nand U5301 (N_5301,N_4455,N_3995);
and U5302 (N_5302,N_4652,N_3759);
nand U5303 (N_5303,N_4413,N_3996);
xor U5304 (N_5304,N_4077,N_4757);
and U5305 (N_5305,N_4410,N_4187);
nand U5306 (N_5306,N_4491,N_4550);
and U5307 (N_5307,N_4246,N_4627);
nor U5308 (N_5308,N_4486,N_4233);
nand U5309 (N_5309,N_3760,N_4284);
nand U5310 (N_5310,N_3991,N_4546);
nor U5311 (N_5311,N_4324,N_4587);
or U5312 (N_5312,N_4366,N_4963);
nand U5313 (N_5313,N_4078,N_4554);
xnor U5314 (N_5314,N_4829,N_4890);
and U5315 (N_5315,N_4043,N_4033);
nand U5316 (N_5316,N_4835,N_4696);
nand U5317 (N_5317,N_4599,N_4496);
nand U5318 (N_5318,N_4607,N_4620);
nor U5319 (N_5319,N_3761,N_4459);
nor U5320 (N_5320,N_4936,N_4259);
xor U5321 (N_5321,N_3968,N_4616);
nor U5322 (N_5322,N_4862,N_3977);
nor U5323 (N_5323,N_4948,N_3980);
xnor U5324 (N_5324,N_4999,N_4747);
xnor U5325 (N_5325,N_4182,N_3806);
and U5326 (N_5326,N_3792,N_4110);
and U5327 (N_5327,N_4347,N_4261);
xnor U5328 (N_5328,N_3984,N_4011);
xor U5329 (N_5329,N_3918,N_4119);
xor U5330 (N_5330,N_4355,N_3766);
xor U5331 (N_5331,N_3959,N_4973);
nand U5332 (N_5332,N_3789,N_4764);
nand U5333 (N_5333,N_4792,N_4898);
nand U5334 (N_5334,N_4247,N_4510);
xor U5335 (N_5335,N_3920,N_4623);
or U5336 (N_5336,N_4417,N_4856);
or U5337 (N_5337,N_4995,N_3912);
xor U5338 (N_5338,N_4785,N_4122);
nand U5339 (N_5339,N_4003,N_4175);
nor U5340 (N_5340,N_4786,N_4647);
xnor U5341 (N_5341,N_3800,N_4021);
and U5342 (N_5342,N_3767,N_4752);
nor U5343 (N_5343,N_4635,N_4953);
nand U5344 (N_5344,N_4461,N_3910);
nand U5345 (N_5345,N_4318,N_4116);
or U5346 (N_5346,N_4625,N_3911);
and U5347 (N_5347,N_4606,N_4698);
or U5348 (N_5348,N_4117,N_4815);
or U5349 (N_5349,N_4349,N_4274);
nand U5350 (N_5350,N_4827,N_4282);
nor U5351 (N_5351,N_3805,N_4799);
nor U5352 (N_5352,N_3894,N_3877);
and U5353 (N_5353,N_4571,N_3860);
xor U5354 (N_5354,N_4280,N_4522);
and U5355 (N_5355,N_3899,N_4502);
or U5356 (N_5356,N_4298,N_4530);
xor U5357 (N_5357,N_4761,N_4755);
nand U5358 (N_5358,N_4863,N_4244);
nor U5359 (N_5359,N_3822,N_4667);
and U5360 (N_5360,N_4668,N_4204);
and U5361 (N_5361,N_4741,N_4169);
xnor U5362 (N_5362,N_4013,N_4853);
and U5363 (N_5363,N_4984,N_4202);
nand U5364 (N_5364,N_4372,N_4659);
xor U5365 (N_5365,N_4669,N_4657);
xor U5366 (N_5366,N_4951,N_4796);
nand U5367 (N_5367,N_4026,N_4423);
nor U5368 (N_5368,N_3837,N_4684);
and U5369 (N_5369,N_4044,N_4336);
xor U5370 (N_5370,N_4338,N_4814);
and U5371 (N_5371,N_4609,N_4825);
nor U5372 (N_5372,N_4564,N_4171);
nand U5373 (N_5373,N_4419,N_4323);
xnor U5374 (N_5374,N_4758,N_4201);
nand U5375 (N_5375,N_4480,N_3924);
or U5376 (N_5376,N_4362,N_4506);
xnor U5377 (N_5377,N_4824,N_4695);
nor U5378 (N_5378,N_4234,N_4926);
and U5379 (N_5379,N_4574,N_4478);
and U5380 (N_5380,N_4189,N_4170);
and U5381 (N_5381,N_4031,N_4443);
xor U5382 (N_5382,N_4726,N_3902);
nor U5383 (N_5383,N_4810,N_3875);
or U5384 (N_5384,N_3948,N_3904);
nor U5385 (N_5385,N_3816,N_4236);
nor U5386 (N_5386,N_3803,N_4356);
xor U5387 (N_5387,N_4920,N_3919);
or U5388 (N_5388,N_4965,N_4840);
xnor U5389 (N_5389,N_4636,N_4197);
xor U5390 (N_5390,N_3957,N_4292);
or U5391 (N_5391,N_4750,N_4561);
nand U5392 (N_5392,N_3978,N_4968);
xor U5393 (N_5393,N_4083,N_4214);
nand U5394 (N_5394,N_4365,N_4744);
nand U5395 (N_5395,N_3975,N_4687);
nor U5396 (N_5396,N_4991,N_4730);
and U5397 (N_5397,N_3791,N_4770);
nor U5398 (N_5398,N_4910,N_3807);
nand U5399 (N_5399,N_3892,N_4055);
and U5400 (N_5400,N_4167,N_4296);
nor U5401 (N_5401,N_3835,N_4295);
xnor U5402 (N_5402,N_4468,N_4252);
nand U5403 (N_5403,N_4787,N_4513);
xnor U5404 (N_5404,N_4376,N_4791);
or U5405 (N_5405,N_4071,N_4560);
and U5406 (N_5406,N_4719,N_4797);
xor U5407 (N_5407,N_3857,N_4225);
nand U5408 (N_5408,N_4464,N_3923);
xnor U5409 (N_5409,N_4231,N_4475);
or U5410 (N_5410,N_4453,N_3850);
nor U5411 (N_5411,N_4699,N_4221);
nor U5412 (N_5412,N_4516,N_3770);
and U5413 (N_5413,N_3990,N_4291);
nor U5414 (N_5414,N_4109,N_4989);
nor U5415 (N_5415,N_4789,N_4662);
nor U5416 (N_5416,N_4959,N_4439);
nand U5417 (N_5417,N_4394,N_4483);
or U5418 (N_5418,N_4813,N_4573);
nor U5419 (N_5419,N_3864,N_3828);
nor U5420 (N_5420,N_3824,N_4760);
nand U5421 (N_5421,N_4006,N_4723);
nor U5422 (N_5422,N_4397,N_4753);
nor U5423 (N_5423,N_4547,N_4084);
and U5424 (N_5424,N_4344,N_4391);
or U5425 (N_5425,N_4320,N_4378);
nor U5426 (N_5426,N_4521,N_3949);
and U5427 (N_5427,N_4140,N_4400);
and U5428 (N_5428,N_3916,N_4603);
nand U5429 (N_5429,N_4686,N_4771);
or U5430 (N_5430,N_4906,N_4992);
nor U5431 (N_5431,N_4337,N_4532);
nand U5432 (N_5432,N_4192,N_4705);
and U5433 (N_5433,N_4460,N_4710);
and U5434 (N_5434,N_4193,N_4188);
xor U5435 (N_5435,N_4368,N_3898);
or U5436 (N_5436,N_4974,N_4762);
nor U5437 (N_5437,N_4148,N_4917);
and U5438 (N_5438,N_4712,N_4300);
and U5439 (N_5439,N_4847,N_4746);
xor U5440 (N_5440,N_4179,N_3873);
and U5441 (N_5441,N_4147,N_3917);
and U5442 (N_5442,N_4542,N_3939);
xor U5443 (N_5443,N_3802,N_4823);
nand U5444 (N_5444,N_4088,N_4541);
xnor U5445 (N_5445,N_3905,N_4333);
nor U5446 (N_5446,N_4207,N_4977);
or U5447 (N_5447,N_4645,N_4555);
or U5448 (N_5448,N_4954,N_4257);
and U5449 (N_5449,N_4671,N_4784);
and U5450 (N_5450,N_4818,N_3987);
nor U5451 (N_5451,N_4641,N_4961);
and U5452 (N_5452,N_4806,N_4889);
nand U5453 (N_5453,N_4582,N_4136);
xnor U5454 (N_5454,N_3775,N_3879);
nand U5455 (N_5455,N_4896,N_4299);
nor U5456 (N_5456,N_4897,N_4405);
xnor U5457 (N_5457,N_4540,N_4082);
and U5458 (N_5458,N_3928,N_3992);
nand U5459 (N_5459,N_4661,N_4017);
nor U5460 (N_5460,N_4005,N_3858);
and U5461 (N_5461,N_4653,N_4138);
xor U5462 (N_5462,N_4887,N_4099);
or U5463 (N_5463,N_3985,N_4273);
nand U5464 (N_5464,N_4731,N_3896);
or U5465 (N_5465,N_4996,N_4857);
or U5466 (N_5466,N_4287,N_4769);
or U5467 (N_5467,N_4040,N_4488);
xnor U5468 (N_5468,N_3966,N_4940);
or U5469 (N_5469,N_3781,N_4492);
nor U5470 (N_5470,N_4229,N_4894);
nand U5471 (N_5471,N_4096,N_4382);
or U5472 (N_5472,N_4441,N_4223);
nand U5473 (N_5473,N_4812,N_4363);
and U5474 (N_5474,N_4660,N_4846);
nor U5475 (N_5475,N_4222,N_3788);
nand U5476 (N_5476,N_4375,N_4370);
or U5477 (N_5477,N_3756,N_4537);
nor U5478 (N_5478,N_4281,N_4074);
xnor U5479 (N_5479,N_4535,N_4048);
or U5480 (N_5480,N_3909,N_4870);
nand U5481 (N_5481,N_4691,N_4869);
xnor U5482 (N_5482,N_4909,N_4027);
or U5483 (N_5483,N_3823,N_4980);
nand U5484 (N_5484,N_4577,N_4736);
nor U5485 (N_5485,N_4219,N_4041);
nor U5486 (N_5486,N_4568,N_4128);
and U5487 (N_5487,N_4462,N_4742);
nor U5488 (N_5488,N_4062,N_4104);
or U5489 (N_5489,N_3925,N_4859);
nand U5490 (N_5490,N_3946,N_4745);
nand U5491 (N_5491,N_4129,N_4049);
or U5492 (N_5492,N_4321,N_3812);
and U5493 (N_5493,N_4972,N_4262);
nand U5494 (N_5494,N_4465,N_4091);
nand U5495 (N_5495,N_4802,N_4557);
nor U5496 (N_5496,N_3769,N_4427);
nand U5497 (N_5497,N_4260,N_4121);
nor U5498 (N_5498,N_4957,N_4022);
xnor U5499 (N_5499,N_4411,N_4519);
or U5500 (N_5500,N_4683,N_4534);
nand U5501 (N_5501,N_4265,N_4808);
and U5502 (N_5502,N_4127,N_4479);
or U5503 (N_5503,N_3848,N_3976);
or U5504 (N_5504,N_4206,N_4790);
and U5505 (N_5505,N_4432,N_3895);
and U5506 (N_5506,N_4579,N_4310);
xnor U5507 (N_5507,N_3786,N_3814);
nor U5508 (N_5508,N_4589,N_4938);
or U5509 (N_5509,N_3907,N_4016);
and U5510 (N_5510,N_4807,N_4591);
nand U5511 (N_5511,N_4458,N_3882);
and U5512 (N_5512,N_4162,N_4895);
and U5513 (N_5513,N_3942,N_4942);
xnor U5514 (N_5514,N_4305,N_4702);
xor U5515 (N_5515,N_4767,N_4046);
or U5516 (N_5516,N_4240,N_4090);
xor U5517 (N_5517,N_4629,N_4611);
nor U5518 (N_5518,N_3870,N_4163);
and U5519 (N_5519,N_3961,N_3941);
and U5520 (N_5520,N_4803,N_4631);
or U5521 (N_5521,N_4097,N_4161);
and U5522 (N_5522,N_4241,N_4670);
nor U5523 (N_5523,N_4173,N_3982);
nor U5524 (N_5524,N_4509,N_3826);
and U5525 (N_5525,N_4733,N_4681);
or U5526 (N_5526,N_4692,N_4395);
or U5527 (N_5527,N_4386,N_4487);
and U5528 (N_5528,N_3887,N_4976);
nor U5529 (N_5529,N_4707,N_4433);
nor U5530 (N_5530,N_4779,N_4473);
nor U5531 (N_5531,N_4907,N_4700);
xnor U5532 (N_5532,N_4552,N_4272);
nor U5533 (N_5533,N_4216,N_4256);
nor U5534 (N_5534,N_3794,N_4604);
and U5535 (N_5535,N_4277,N_4353);
and U5536 (N_5536,N_4387,N_4893);
xor U5537 (N_5537,N_4526,N_4632);
nand U5538 (N_5538,N_4768,N_4651);
nand U5539 (N_5539,N_3841,N_4539);
nor U5540 (N_5540,N_3751,N_4981);
xor U5541 (N_5541,N_4398,N_4899);
and U5542 (N_5542,N_4566,N_4949);
or U5543 (N_5543,N_4676,N_3829);
nand U5544 (N_5544,N_4633,N_4644);
or U5545 (N_5545,N_4190,N_4722);
or U5546 (N_5546,N_4107,N_4070);
nor U5547 (N_5547,N_4436,N_4030);
xnor U5548 (N_5548,N_3901,N_3753);
or U5549 (N_5549,N_4381,N_4515);
and U5550 (N_5550,N_4311,N_4580);
xnor U5551 (N_5551,N_4151,N_3921);
nand U5552 (N_5552,N_4527,N_4872);
nor U5553 (N_5553,N_4442,N_4679);
nand U5554 (N_5554,N_4266,N_3950);
xnor U5555 (N_5555,N_4389,N_4334);
or U5556 (N_5556,N_4709,N_3965);
nand U5557 (N_5557,N_3861,N_4165);
nand U5558 (N_5558,N_4966,N_4348);
or U5559 (N_5559,N_3771,N_4932);
or U5560 (N_5560,N_4149,N_4817);
or U5561 (N_5561,N_4919,N_4361);
nor U5562 (N_5562,N_4158,N_4727);
and U5563 (N_5563,N_4012,N_4346);
nor U5564 (N_5564,N_4371,N_4042);
and U5565 (N_5565,N_4520,N_4431);
and U5566 (N_5566,N_4301,N_4430);
xnor U5567 (N_5567,N_4319,N_3868);
xnor U5568 (N_5568,N_4086,N_4406);
xnor U5569 (N_5569,N_4052,N_4673);
or U5570 (N_5570,N_4130,N_4388);
xnor U5571 (N_5571,N_4931,N_4804);
or U5572 (N_5572,N_4852,N_4880);
or U5573 (N_5573,N_4602,N_4499);
nand U5574 (N_5574,N_4307,N_3969);
nand U5575 (N_5575,N_4454,N_3843);
and U5576 (N_5576,N_4783,N_3967);
or U5577 (N_5577,N_4471,N_3863);
xnor U5578 (N_5578,N_4584,N_3839);
and U5579 (N_5579,N_4739,N_4180);
xor U5580 (N_5580,N_3834,N_4988);
or U5581 (N_5581,N_4778,N_4053);
or U5582 (N_5582,N_4970,N_4036);
xnor U5583 (N_5583,N_4384,N_4911);
nor U5584 (N_5584,N_3809,N_3790);
nor U5585 (N_5585,N_3827,N_4612);
and U5586 (N_5586,N_3817,N_4637);
nor U5587 (N_5587,N_4408,N_4060);
and U5588 (N_5588,N_4545,N_4054);
nand U5589 (N_5589,N_4572,N_3956);
and U5590 (N_5590,N_4000,N_4237);
or U5591 (N_5591,N_4444,N_4211);
nand U5592 (N_5592,N_3799,N_4327);
or U5593 (N_5593,N_4114,N_4597);
or U5594 (N_5594,N_4485,N_4312);
nor U5595 (N_5595,N_4774,N_3890);
xnor U5596 (N_5596,N_4688,N_4994);
nand U5597 (N_5597,N_4902,N_4694);
xor U5598 (N_5598,N_3935,N_4466);
or U5599 (N_5599,N_4294,N_3798);
nor U5600 (N_5600,N_4927,N_3813);
nand U5601 (N_5601,N_3962,N_4939);
nor U5602 (N_5602,N_4065,N_4330);
nand U5603 (N_5603,N_3986,N_4875);
nand U5604 (N_5604,N_4586,N_4402);
nor U5605 (N_5605,N_3854,N_4160);
xor U5606 (N_5606,N_4738,N_3777);
nand U5607 (N_5607,N_4434,N_4654);
xnor U5608 (N_5608,N_3784,N_4518);
and U5609 (N_5609,N_4578,N_4704);
xor U5610 (N_5610,N_4946,N_4404);
or U5611 (N_5611,N_4891,N_4238);
xor U5612 (N_5612,N_4357,N_3768);
nor U5613 (N_5613,N_4469,N_4508);
nor U5614 (N_5614,N_4172,N_3988);
or U5615 (N_5615,N_4098,N_4765);
nand U5616 (N_5616,N_4364,N_4711);
nand U5617 (N_5617,N_4640,N_4057);
and U5618 (N_5618,N_4501,N_3945);
nor U5619 (N_5619,N_4718,N_4415);
or U5620 (N_5620,N_4851,N_4360);
nor U5621 (N_5621,N_3762,N_4066);
xor U5622 (N_5622,N_4403,N_4251);
nor U5623 (N_5623,N_4076,N_3832);
nor U5624 (N_5624,N_4871,N_4986);
nor U5625 (N_5625,N_4741,N_4062);
nor U5626 (N_5626,N_4476,N_3788);
nand U5627 (N_5627,N_4604,N_3938);
and U5628 (N_5628,N_3893,N_4823);
xor U5629 (N_5629,N_4216,N_4289);
nand U5630 (N_5630,N_4853,N_4059);
or U5631 (N_5631,N_4941,N_4678);
nand U5632 (N_5632,N_4640,N_4441);
and U5633 (N_5633,N_4997,N_4125);
xor U5634 (N_5634,N_4450,N_4927);
nor U5635 (N_5635,N_3947,N_4915);
or U5636 (N_5636,N_4617,N_4092);
or U5637 (N_5637,N_3864,N_4924);
nor U5638 (N_5638,N_4428,N_4369);
or U5639 (N_5639,N_4024,N_4567);
or U5640 (N_5640,N_4033,N_3835);
nor U5641 (N_5641,N_4483,N_4251);
or U5642 (N_5642,N_3919,N_4917);
or U5643 (N_5643,N_4821,N_4268);
nor U5644 (N_5644,N_4743,N_4466);
nand U5645 (N_5645,N_4387,N_4021);
nor U5646 (N_5646,N_3758,N_4919);
or U5647 (N_5647,N_4483,N_4954);
xor U5648 (N_5648,N_3853,N_4195);
xor U5649 (N_5649,N_4607,N_4729);
and U5650 (N_5650,N_4535,N_3941);
and U5651 (N_5651,N_3893,N_4759);
xnor U5652 (N_5652,N_4602,N_4188);
nand U5653 (N_5653,N_4025,N_4209);
and U5654 (N_5654,N_4534,N_4315);
or U5655 (N_5655,N_4921,N_3917);
nor U5656 (N_5656,N_3974,N_4256);
or U5657 (N_5657,N_4344,N_4139);
or U5658 (N_5658,N_4465,N_4167);
nand U5659 (N_5659,N_4104,N_4792);
nand U5660 (N_5660,N_3955,N_4273);
nor U5661 (N_5661,N_4483,N_4652);
or U5662 (N_5662,N_3871,N_4862);
and U5663 (N_5663,N_4999,N_4169);
or U5664 (N_5664,N_4272,N_4101);
and U5665 (N_5665,N_4167,N_4694);
xnor U5666 (N_5666,N_4055,N_3872);
xor U5667 (N_5667,N_4938,N_4064);
or U5668 (N_5668,N_3984,N_4856);
nand U5669 (N_5669,N_3942,N_4795);
or U5670 (N_5670,N_3755,N_4385);
xor U5671 (N_5671,N_4382,N_3824);
nand U5672 (N_5672,N_4174,N_4980);
or U5673 (N_5673,N_4408,N_4588);
and U5674 (N_5674,N_4003,N_4461);
nand U5675 (N_5675,N_4419,N_3887);
nand U5676 (N_5676,N_3984,N_3912);
xnor U5677 (N_5677,N_4611,N_4795);
nor U5678 (N_5678,N_3760,N_3751);
or U5679 (N_5679,N_3941,N_4376);
and U5680 (N_5680,N_4267,N_3960);
or U5681 (N_5681,N_4223,N_4072);
xnor U5682 (N_5682,N_4871,N_3877);
and U5683 (N_5683,N_3942,N_4446);
nor U5684 (N_5684,N_4776,N_4031);
nor U5685 (N_5685,N_4802,N_4233);
and U5686 (N_5686,N_4565,N_3781);
nand U5687 (N_5687,N_4051,N_3959);
and U5688 (N_5688,N_4764,N_4755);
or U5689 (N_5689,N_4471,N_4224);
xnor U5690 (N_5690,N_4347,N_3792);
nor U5691 (N_5691,N_3978,N_4263);
nor U5692 (N_5692,N_4323,N_4431);
or U5693 (N_5693,N_4330,N_4416);
xor U5694 (N_5694,N_4421,N_3973);
or U5695 (N_5695,N_4360,N_3906);
xor U5696 (N_5696,N_3812,N_4898);
xnor U5697 (N_5697,N_4675,N_3832);
or U5698 (N_5698,N_3948,N_4318);
and U5699 (N_5699,N_4422,N_4018);
nand U5700 (N_5700,N_4935,N_4695);
or U5701 (N_5701,N_4191,N_4269);
and U5702 (N_5702,N_3875,N_3774);
nand U5703 (N_5703,N_4839,N_4161);
xnor U5704 (N_5704,N_4812,N_4333);
nor U5705 (N_5705,N_4210,N_4892);
or U5706 (N_5706,N_4792,N_4202);
xnor U5707 (N_5707,N_4782,N_3923);
and U5708 (N_5708,N_3996,N_4246);
or U5709 (N_5709,N_3956,N_4591);
nand U5710 (N_5710,N_4704,N_4031);
or U5711 (N_5711,N_4140,N_4830);
and U5712 (N_5712,N_4552,N_3934);
xor U5713 (N_5713,N_4432,N_4272);
nor U5714 (N_5714,N_4732,N_4088);
nor U5715 (N_5715,N_4193,N_4443);
and U5716 (N_5716,N_4081,N_4893);
or U5717 (N_5717,N_4117,N_4679);
nor U5718 (N_5718,N_4688,N_3774);
or U5719 (N_5719,N_4879,N_4469);
or U5720 (N_5720,N_4746,N_4218);
and U5721 (N_5721,N_4741,N_4273);
nor U5722 (N_5722,N_4097,N_3838);
and U5723 (N_5723,N_4551,N_4630);
xnor U5724 (N_5724,N_4842,N_4452);
and U5725 (N_5725,N_4676,N_4060);
or U5726 (N_5726,N_4953,N_4122);
or U5727 (N_5727,N_4691,N_4419);
or U5728 (N_5728,N_3908,N_4043);
nor U5729 (N_5729,N_3827,N_4486);
nand U5730 (N_5730,N_4454,N_4940);
xor U5731 (N_5731,N_3991,N_4238);
nor U5732 (N_5732,N_3788,N_4164);
xor U5733 (N_5733,N_4884,N_3813);
and U5734 (N_5734,N_4070,N_3990);
xor U5735 (N_5735,N_4105,N_4443);
nand U5736 (N_5736,N_4849,N_3758);
nor U5737 (N_5737,N_4661,N_4881);
nor U5738 (N_5738,N_4408,N_4771);
nor U5739 (N_5739,N_4180,N_4916);
xnor U5740 (N_5740,N_4686,N_3974);
xor U5741 (N_5741,N_4729,N_4816);
nand U5742 (N_5742,N_4643,N_4939);
nor U5743 (N_5743,N_4224,N_4472);
xnor U5744 (N_5744,N_4110,N_4473);
or U5745 (N_5745,N_3864,N_4397);
nand U5746 (N_5746,N_4061,N_3864);
xor U5747 (N_5747,N_4596,N_3998);
nand U5748 (N_5748,N_3988,N_4921);
xnor U5749 (N_5749,N_4010,N_4013);
or U5750 (N_5750,N_4888,N_4179);
nand U5751 (N_5751,N_4913,N_4316);
and U5752 (N_5752,N_4122,N_4916);
xnor U5753 (N_5753,N_4238,N_4023);
nand U5754 (N_5754,N_4312,N_4284);
xor U5755 (N_5755,N_4777,N_4839);
nor U5756 (N_5756,N_4059,N_4604);
and U5757 (N_5757,N_4609,N_4178);
nor U5758 (N_5758,N_4947,N_4758);
nand U5759 (N_5759,N_3916,N_3781);
xnor U5760 (N_5760,N_3937,N_4311);
xor U5761 (N_5761,N_4154,N_4185);
nor U5762 (N_5762,N_4613,N_4212);
and U5763 (N_5763,N_4460,N_4797);
nor U5764 (N_5764,N_4289,N_4797);
nand U5765 (N_5765,N_3971,N_4952);
or U5766 (N_5766,N_4163,N_3755);
and U5767 (N_5767,N_4770,N_3755);
xor U5768 (N_5768,N_4699,N_4607);
or U5769 (N_5769,N_3764,N_3970);
xor U5770 (N_5770,N_4166,N_3885);
or U5771 (N_5771,N_3979,N_4236);
nand U5772 (N_5772,N_4002,N_4762);
xor U5773 (N_5773,N_4934,N_4228);
nand U5774 (N_5774,N_3773,N_4835);
or U5775 (N_5775,N_4546,N_4470);
and U5776 (N_5776,N_4090,N_4943);
and U5777 (N_5777,N_4335,N_4013);
nor U5778 (N_5778,N_4415,N_4609);
nor U5779 (N_5779,N_4864,N_3906);
and U5780 (N_5780,N_4986,N_4506);
nor U5781 (N_5781,N_4845,N_4768);
and U5782 (N_5782,N_4698,N_3812);
and U5783 (N_5783,N_4640,N_4687);
nand U5784 (N_5784,N_4976,N_3910);
xor U5785 (N_5785,N_3947,N_3851);
and U5786 (N_5786,N_4416,N_4643);
or U5787 (N_5787,N_4278,N_4543);
or U5788 (N_5788,N_4068,N_4683);
and U5789 (N_5789,N_4368,N_4301);
and U5790 (N_5790,N_4633,N_4710);
or U5791 (N_5791,N_4483,N_3760);
and U5792 (N_5792,N_4576,N_4358);
nand U5793 (N_5793,N_4287,N_3783);
and U5794 (N_5794,N_4946,N_3908);
xnor U5795 (N_5795,N_4566,N_4930);
or U5796 (N_5796,N_4979,N_4790);
xnor U5797 (N_5797,N_4897,N_4085);
nor U5798 (N_5798,N_4705,N_4258);
nor U5799 (N_5799,N_4320,N_4991);
and U5800 (N_5800,N_3911,N_3924);
xor U5801 (N_5801,N_4026,N_4413);
nand U5802 (N_5802,N_4276,N_4843);
nand U5803 (N_5803,N_4603,N_4723);
or U5804 (N_5804,N_4042,N_4381);
and U5805 (N_5805,N_4265,N_4128);
nor U5806 (N_5806,N_4983,N_4974);
nor U5807 (N_5807,N_3973,N_4775);
nand U5808 (N_5808,N_4788,N_4623);
xor U5809 (N_5809,N_3876,N_4924);
nor U5810 (N_5810,N_4274,N_3959);
xnor U5811 (N_5811,N_4724,N_4888);
nor U5812 (N_5812,N_4088,N_4256);
xor U5813 (N_5813,N_4734,N_4587);
nand U5814 (N_5814,N_4441,N_4410);
nand U5815 (N_5815,N_4927,N_4299);
nor U5816 (N_5816,N_3971,N_4007);
or U5817 (N_5817,N_4858,N_4639);
or U5818 (N_5818,N_4257,N_4560);
xnor U5819 (N_5819,N_4899,N_4121);
nand U5820 (N_5820,N_4844,N_4010);
or U5821 (N_5821,N_4805,N_4288);
and U5822 (N_5822,N_4542,N_4909);
nand U5823 (N_5823,N_4888,N_4631);
nor U5824 (N_5824,N_4172,N_4594);
or U5825 (N_5825,N_4192,N_4072);
and U5826 (N_5826,N_4732,N_4993);
xnor U5827 (N_5827,N_4395,N_4637);
xnor U5828 (N_5828,N_4511,N_4886);
xor U5829 (N_5829,N_3997,N_4443);
and U5830 (N_5830,N_4586,N_4727);
xor U5831 (N_5831,N_4392,N_4535);
or U5832 (N_5832,N_4032,N_4830);
nand U5833 (N_5833,N_4390,N_4677);
xnor U5834 (N_5834,N_4694,N_4123);
nand U5835 (N_5835,N_4570,N_4883);
nand U5836 (N_5836,N_3981,N_4175);
or U5837 (N_5837,N_4203,N_4615);
nor U5838 (N_5838,N_3834,N_4020);
or U5839 (N_5839,N_3973,N_4128);
or U5840 (N_5840,N_3755,N_4358);
and U5841 (N_5841,N_4744,N_4055);
or U5842 (N_5842,N_4880,N_3751);
xnor U5843 (N_5843,N_3985,N_4588);
or U5844 (N_5844,N_4525,N_4911);
and U5845 (N_5845,N_4778,N_4759);
or U5846 (N_5846,N_4896,N_4173);
and U5847 (N_5847,N_4862,N_3802);
nor U5848 (N_5848,N_4464,N_4627);
or U5849 (N_5849,N_3766,N_4438);
nor U5850 (N_5850,N_4805,N_4454);
nor U5851 (N_5851,N_4697,N_4068);
or U5852 (N_5852,N_4632,N_4515);
nand U5853 (N_5853,N_4841,N_4965);
nor U5854 (N_5854,N_3853,N_3884);
nor U5855 (N_5855,N_4967,N_4592);
nand U5856 (N_5856,N_3889,N_4177);
nor U5857 (N_5857,N_4599,N_3764);
or U5858 (N_5858,N_4465,N_4090);
and U5859 (N_5859,N_4350,N_3952);
nor U5860 (N_5860,N_4310,N_4364);
xor U5861 (N_5861,N_4506,N_3895);
and U5862 (N_5862,N_4462,N_4702);
and U5863 (N_5863,N_3995,N_4802);
nor U5864 (N_5864,N_3759,N_3954);
nor U5865 (N_5865,N_3968,N_4015);
nand U5866 (N_5866,N_4321,N_4366);
xnor U5867 (N_5867,N_4743,N_4906);
and U5868 (N_5868,N_4213,N_4952);
xor U5869 (N_5869,N_3960,N_3901);
nor U5870 (N_5870,N_4396,N_3781);
and U5871 (N_5871,N_4872,N_4492);
nand U5872 (N_5872,N_4859,N_4032);
or U5873 (N_5873,N_3812,N_4827);
and U5874 (N_5874,N_4522,N_4913);
nor U5875 (N_5875,N_3859,N_4104);
or U5876 (N_5876,N_4191,N_4238);
and U5877 (N_5877,N_3970,N_4926);
xnor U5878 (N_5878,N_3960,N_4565);
xor U5879 (N_5879,N_4031,N_4877);
nor U5880 (N_5880,N_4344,N_4717);
nor U5881 (N_5881,N_4712,N_4653);
nor U5882 (N_5882,N_4900,N_3766);
nand U5883 (N_5883,N_4432,N_4640);
xor U5884 (N_5884,N_4557,N_3787);
nor U5885 (N_5885,N_4609,N_4845);
and U5886 (N_5886,N_4628,N_3862);
xnor U5887 (N_5887,N_4149,N_4209);
nor U5888 (N_5888,N_4658,N_4760);
nand U5889 (N_5889,N_4019,N_3886);
and U5890 (N_5890,N_4624,N_3948);
xor U5891 (N_5891,N_4588,N_4749);
nand U5892 (N_5892,N_4815,N_4326);
or U5893 (N_5893,N_4997,N_4669);
xor U5894 (N_5894,N_4016,N_4766);
xor U5895 (N_5895,N_4327,N_4086);
nand U5896 (N_5896,N_4314,N_4608);
nor U5897 (N_5897,N_3997,N_4619);
nor U5898 (N_5898,N_4461,N_4356);
xor U5899 (N_5899,N_4726,N_3988);
and U5900 (N_5900,N_4006,N_4799);
nand U5901 (N_5901,N_4915,N_4989);
nor U5902 (N_5902,N_4938,N_3973);
nor U5903 (N_5903,N_3831,N_4328);
and U5904 (N_5904,N_3901,N_4293);
xor U5905 (N_5905,N_4513,N_3975);
xor U5906 (N_5906,N_4148,N_4228);
nor U5907 (N_5907,N_4246,N_3908);
nor U5908 (N_5908,N_4644,N_4300);
or U5909 (N_5909,N_3901,N_4296);
or U5910 (N_5910,N_4104,N_4949);
nand U5911 (N_5911,N_4132,N_3922);
xnor U5912 (N_5912,N_3979,N_4871);
nand U5913 (N_5913,N_4952,N_3863);
and U5914 (N_5914,N_4518,N_4974);
nor U5915 (N_5915,N_4704,N_4916);
nand U5916 (N_5916,N_4600,N_4991);
nor U5917 (N_5917,N_4037,N_4223);
and U5918 (N_5918,N_4238,N_4583);
nand U5919 (N_5919,N_3835,N_3979);
xor U5920 (N_5920,N_4174,N_4062);
xnor U5921 (N_5921,N_4616,N_4910);
nor U5922 (N_5922,N_4753,N_4441);
nor U5923 (N_5923,N_4549,N_3761);
nor U5924 (N_5924,N_3950,N_4222);
xnor U5925 (N_5925,N_4330,N_4157);
or U5926 (N_5926,N_4813,N_4894);
xor U5927 (N_5927,N_4763,N_3988);
nor U5928 (N_5928,N_3877,N_4528);
nor U5929 (N_5929,N_4644,N_4741);
or U5930 (N_5930,N_3906,N_4730);
xor U5931 (N_5931,N_4664,N_3976);
and U5932 (N_5932,N_4264,N_3922);
or U5933 (N_5933,N_3889,N_3925);
xnor U5934 (N_5934,N_4019,N_4941);
xor U5935 (N_5935,N_4023,N_4781);
and U5936 (N_5936,N_4938,N_3835);
nor U5937 (N_5937,N_4068,N_4021);
and U5938 (N_5938,N_4043,N_4905);
and U5939 (N_5939,N_4671,N_4403);
nand U5940 (N_5940,N_4623,N_4649);
nand U5941 (N_5941,N_4438,N_4247);
xnor U5942 (N_5942,N_4837,N_4072);
nand U5943 (N_5943,N_4756,N_3884);
nor U5944 (N_5944,N_4623,N_4292);
xnor U5945 (N_5945,N_4723,N_4141);
or U5946 (N_5946,N_4598,N_4665);
and U5947 (N_5947,N_4163,N_4931);
nor U5948 (N_5948,N_4152,N_3888);
and U5949 (N_5949,N_4117,N_3976);
or U5950 (N_5950,N_4331,N_3983);
xnor U5951 (N_5951,N_4986,N_3938);
and U5952 (N_5952,N_4393,N_4767);
or U5953 (N_5953,N_4741,N_4235);
xnor U5954 (N_5954,N_4579,N_3888);
nand U5955 (N_5955,N_4217,N_3764);
and U5956 (N_5956,N_4456,N_4748);
nor U5957 (N_5957,N_4752,N_4480);
or U5958 (N_5958,N_4460,N_3818);
or U5959 (N_5959,N_4227,N_4996);
or U5960 (N_5960,N_4615,N_4542);
and U5961 (N_5961,N_4579,N_4572);
nand U5962 (N_5962,N_3780,N_4945);
and U5963 (N_5963,N_3794,N_4627);
xnor U5964 (N_5964,N_3786,N_4049);
nor U5965 (N_5965,N_4463,N_4001);
nand U5966 (N_5966,N_3982,N_4238);
or U5967 (N_5967,N_4082,N_4339);
and U5968 (N_5968,N_3757,N_4251);
or U5969 (N_5969,N_3814,N_4048);
and U5970 (N_5970,N_4904,N_4717);
xor U5971 (N_5971,N_4787,N_4487);
xnor U5972 (N_5972,N_4797,N_4812);
nand U5973 (N_5973,N_4723,N_4548);
nand U5974 (N_5974,N_4613,N_4279);
or U5975 (N_5975,N_4878,N_4647);
or U5976 (N_5976,N_4830,N_4909);
xor U5977 (N_5977,N_4032,N_3764);
xnor U5978 (N_5978,N_3910,N_4543);
or U5979 (N_5979,N_4751,N_4333);
nor U5980 (N_5980,N_4647,N_4806);
nor U5981 (N_5981,N_4278,N_4108);
xnor U5982 (N_5982,N_4859,N_4843);
nor U5983 (N_5983,N_3920,N_4683);
or U5984 (N_5984,N_4662,N_3866);
nand U5985 (N_5985,N_4779,N_4705);
and U5986 (N_5986,N_3770,N_3974);
xnor U5987 (N_5987,N_4600,N_4800);
nor U5988 (N_5988,N_4146,N_4480);
nor U5989 (N_5989,N_4797,N_4870);
xor U5990 (N_5990,N_4980,N_4290);
nand U5991 (N_5991,N_4110,N_4271);
xor U5992 (N_5992,N_3917,N_4344);
xnor U5993 (N_5993,N_3827,N_4916);
and U5994 (N_5994,N_4573,N_4153);
xnor U5995 (N_5995,N_4083,N_3812);
nand U5996 (N_5996,N_3759,N_4135);
xnor U5997 (N_5997,N_4992,N_4807);
nor U5998 (N_5998,N_3839,N_3790);
or U5999 (N_5999,N_4056,N_4137);
or U6000 (N_6000,N_3766,N_4931);
and U6001 (N_6001,N_4173,N_4534);
nand U6002 (N_6002,N_4302,N_4533);
nand U6003 (N_6003,N_4150,N_4599);
xnor U6004 (N_6004,N_3926,N_4937);
xnor U6005 (N_6005,N_4455,N_4784);
or U6006 (N_6006,N_4428,N_4836);
nand U6007 (N_6007,N_4198,N_4291);
or U6008 (N_6008,N_4454,N_4814);
xnor U6009 (N_6009,N_4472,N_3767);
nand U6010 (N_6010,N_4859,N_4252);
or U6011 (N_6011,N_4717,N_4839);
xnor U6012 (N_6012,N_4174,N_4409);
xnor U6013 (N_6013,N_4826,N_4945);
and U6014 (N_6014,N_3939,N_4470);
xnor U6015 (N_6015,N_4461,N_4518);
nand U6016 (N_6016,N_4369,N_4873);
nand U6017 (N_6017,N_4123,N_4145);
xnor U6018 (N_6018,N_3908,N_4045);
or U6019 (N_6019,N_4813,N_3761);
or U6020 (N_6020,N_4252,N_4813);
xnor U6021 (N_6021,N_4974,N_4754);
nor U6022 (N_6022,N_3911,N_4174);
and U6023 (N_6023,N_4757,N_4905);
and U6024 (N_6024,N_3962,N_3815);
nand U6025 (N_6025,N_4986,N_3902);
nand U6026 (N_6026,N_3833,N_4513);
nor U6027 (N_6027,N_4565,N_4110);
and U6028 (N_6028,N_4725,N_4290);
or U6029 (N_6029,N_4554,N_4347);
nand U6030 (N_6030,N_4027,N_4882);
and U6031 (N_6031,N_4351,N_4239);
nand U6032 (N_6032,N_4130,N_4520);
nand U6033 (N_6033,N_3761,N_4078);
xor U6034 (N_6034,N_3793,N_4976);
nand U6035 (N_6035,N_4992,N_4805);
nor U6036 (N_6036,N_3804,N_4985);
or U6037 (N_6037,N_3892,N_3863);
and U6038 (N_6038,N_4152,N_4860);
nor U6039 (N_6039,N_4774,N_4347);
nand U6040 (N_6040,N_4164,N_4046);
or U6041 (N_6041,N_3840,N_4422);
xor U6042 (N_6042,N_3805,N_4385);
and U6043 (N_6043,N_4180,N_4687);
nor U6044 (N_6044,N_4503,N_3755);
or U6045 (N_6045,N_4036,N_4717);
or U6046 (N_6046,N_4599,N_4452);
nand U6047 (N_6047,N_4412,N_4685);
xor U6048 (N_6048,N_3870,N_4476);
nand U6049 (N_6049,N_4565,N_4939);
or U6050 (N_6050,N_3897,N_4470);
nor U6051 (N_6051,N_4053,N_4012);
xor U6052 (N_6052,N_4164,N_4363);
nor U6053 (N_6053,N_4193,N_4080);
nor U6054 (N_6054,N_4190,N_4576);
xnor U6055 (N_6055,N_4644,N_4298);
xor U6056 (N_6056,N_3765,N_4266);
xnor U6057 (N_6057,N_3937,N_4386);
nand U6058 (N_6058,N_3941,N_4684);
or U6059 (N_6059,N_3962,N_4678);
nand U6060 (N_6060,N_3883,N_3852);
xor U6061 (N_6061,N_4624,N_4270);
and U6062 (N_6062,N_4577,N_3837);
or U6063 (N_6063,N_4724,N_3843);
and U6064 (N_6064,N_4943,N_4789);
nor U6065 (N_6065,N_4642,N_4132);
and U6066 (N_6066,N_4767,N_4471);
xnor U6067 (N_6067,N_4018,N_4336);
nand U6068 (N_6068,N_3984,N_4245);
or U6069 (N_6069,N_4483,N_4265);
nor U6070 (N_6070,N_4182,N_4528);
and U6071 (N_6071,N_3818,N_3954);
nor U6072 (N_6072,N_4208,N_4979);
xnor U6073 (N_6073,N_4260,N_4481);
xor U6074 (N_6074,N_4649,N_4275);
xor U6075 (N_6075,N_4918,N_4717);
nand U6076 (N_6076,N_4121,N_3965);
nor U6077 (N_6077,N_3866,N_3839);
xnor U6078 (N_6078,N_3779,N_4490);
or U6079 (N_6079,N_3862,N_3979);
and U6080 (N_6080,N_4934,N_4672);
nand U6081 (N_6081,N_4379,N_4372);
xnor U6082 (N_6082,N_4017,N_4631);
xor U6083 (N_6083,N_4442,N_3987);
nor U6084 (N_6084,N_4679,N_4189);
nand U6085 (N_6085,N_4258,N_4778);
and U6086 (N_6086,N_4314,N_3908);
or U6087 (N_6087,N_4936,N_4225);
xor U6088 (N_6088,N_3906,N_4651);
nand U6089 (N_6089,N_4445,N_4050);
or U6090 (N_6090,N_4413,N_3829);
nand U6091 (N_6091,N_4589,N_4670);
or U6092 (N_6092,N_3982,N_3941);
nand U6093 (N_6093,N_4256,N_4928);
nor U6094 (N_6094,N_4877,N_4168);
nand U6095 (N_6095,N_4854,N_4062);
and U6096 (N_6096,N_3881,N_3996);
nor U6097 (N_6097,N_4143,N_4581);
nand U6098 (N_6098,N_4475,N_4618);
nor U6099 (N_6099,N_4672,N_3993);
nor U6100 (N_6100,N_4371,N_4575);
and U6101 (N_6101,N_4332,N_4348);
nand U6102 (N_6102,N_4899,N_3791);
nor U6103 (N_6103,N_4833,N_4342);
xor U6104 (N_6104,N_4108,N_4653);
nand U6105 (N_6105,N_4315,N_4374);
nand U6106 (N_6106,N_3853,N_4152);
nand U6107 (N_6107,N_4753,N_4160);
nand U6108 (N_6108,N_4968,N_4131);
or U6109 (N_6109,N_3886,N_4927);
nor U6110 (N_6110,N_4735,N_4809);
or U6111 (N_6111,N_4735,N_4759);
nor U6112 (N_6112,N_4575,N_4618);
nand U6113 (N_6113,N_4947,N_4301);
nand U6114 (N_6114,N_4205,N_4266);
nor U6115 (N_6115,N_4158,N_4216);
and U6116 (N_6116,N_4987,N_4434);
xnor U6117 (N_6117,N_4138,N_4401);
or U6118 (N_6118,N_3778,N_3810);
or U6119 (N_6119,N_3865,N_4331);
nor U6120 (N_6120,N_4658,N_4599);
and U6121 (N_6121,N_4537,N_4277);
nand U6122 (N_6122,N_4054,N_4650);
xor U6123 (N_6123,N_4623,N_4850);
and U6124 (N_6124,N_4363,N_4406);
xor U6125 (N_6125,N_4128,N_4277);
xnor U6126 (N_6126,N_4323,N_4788);
xnor U6127 (N_6127,N_4004,N_4253);
and U6128 (N_6128,N_4738,N_4602);
xnor U6129 (N_6129,N_3893,N_3937);
nor U6130 (N_6130,N_4599,N_3894);
nor U6131 (N_6131,N_4170,N_4662);
nor U6132 (N_6132,N_4257,N_4816);
or U6133 (N_6133,N_4253,N_3954);
nand U6134 (N_6134,N_4881,N_3992);
xor U6135 (N_6135,N_4432,N_4853);
nor U6136 (N_6136,N_4732,N_4695);
xnor U6137 (N_6137,N_3784,N_4475);
and U6138 (N_6138,N_4090,N_4625);
xor U6139 (N_6139,N_4998,N_4514);
nand U6140 (N_6140,N_4806,N_4491);
nand U6141 (N_6141,N_4229,N_4807);
and U6142 (N_6142,N_4907,N_4820);
xnor U6143 (N_6143,N_4284,N_3808);
or U6144 (N_6144,N_4668,N_4447);
or U6145 (N_6145,N_4996,N_4232);
xnor U6146 (N_6146,N_4429,N_4301);
xnor U6147 (N_6147,N_4953,N_4134);
xnor U6148 (N_6148,N_4549,N_4810);
and U6149 (N_6149,N_4008,N_3923);
nand U6150 (N_6150,N_3801,N_4313);
and U6151 (N_6151,N_4661,N_4949);
or U6152 (N_6152,N_4313,N_3853);
xnor U6153 (N_6153,N_4704,N_4712);
xnor U6154 (N_6154,N_3800,N_4565);
xnor U6155 (N_6155,N_4468,N_4792);
nand U6156 (N_6156,N_4366,N_4424);
and U6157 (N_6157,N_4703,N_4925);
nor U6158 (N_6158,N_4608,N_4914);
nor U6159 (N_6159,N_4557,N_4587);
nand U6160 (N_6160,N_4706,N_4756);
nand U6161 (N_6161,N_3805,N_3904);
xor U6162 (N_6162,N_3944,N_4729);
nand U6163 (N_6163,N_4047,N_4913);
nor U6164 (N_6164,N_4858,N_3783);
or U6165 (N_6165,N_4414,N_4728);
nand U6166 (N_6166,N_4107,N_4626);
nor U6167 (N_6167,N_4149,N_4306);
nand U6168 (N_6168,N_4590,N_4589);
nor U6169 (N_6169,N_3783,N_4510);
nand U6170 (N_6170,N_4421,N_4186);
xnor U6171 (N_6171,N_4411,N_4469);
and U6172 (N_6172,N_4430,N_4155);
nand U6173 (N_6173,N_3871,N_4376);
or U6174 (N_6174,N_4868,N_4137);
nor U6175 (N_6175,N_4829,N_4133);
nand U6176 (N_6176,N_3952,N_4713);
xor U6177 (N_6177,N_3832,N_4438);
nor U6178 (N_6178,N_4846,N_4819);
xor U6179 (N_6179,N_3768,N_4627);
nor U6180 (N_6180,N_4205,N_4791);
nand U6181 (N_6181,N_4441,N_4538);
xnor U6182 (N_6182,N_4134,N_4170);
and U6183 (N_6183,N_4742,N_4000);
xor U6184 (N_6184,N_4711,N_4815);
or U6185 (N_6185,N_4997,N_4208);
and U6186 (N_6186,N_4960,N_3861);
xor U6187 (N_6187,N_4954,N_4472);
and U6188 (N_6188,N_4368,N_4003);
nor U6189 (N_6189,N_4756,N_4463);
or U6190 (N_6190,N_4113,N_3920);
and U6191 (N_6191,N_3842,N_4974);
nor U6192 (N_6192,N_4216,N_4870);
nor U6193 (N_6193,N_4470,N_3893);
nand U6194 (N_6194,N_4610,N_4579);
and U6195 (N_6195,N_4260,N_4052);
nand U6196 (N_6196,N_3996,N_4368);
or U6197 (N_6197,N_4924,N_4696);
xor U6198 (N_6198,N_4311,N_3810);
xor U6199 (N_6199,N_3837,N_4101);
and U6200 (N_6200,N_4232,N_4428);
xor U6201 (N_6201,N_4902,N_4910);
nand U6202 (N_6202,N_3914,N_4034);
and U6203 (N_6203,N_3926,N_4941);
or U6204 (N_6204,N_4073,N_4137);
or U6205 (N_6205,N_3775,N_4695);
nand U6206 (N_6206,N_4771,N_4368);
or U6207 (N_6207,N_4239,N_4565);
or U6208 (N_6208,N_4178,N_3770);
or U6209 (N_6209,N_4942,N_3957);
nor U6210 (N_6210,N_4013,N_4101);
nor U6211 (N_6211,N_3871,N_3905);
nand U6212 (N_6212,N_4470,N_4988);
nor U6213 (N_6213,N_4396,N_3779);
or U6214 (N_6214,N_4298,N_4301);
xor U6215 (N_6215,N_4991,N_4175);
and U6216 (N_6216,N_4480,N_4743);
and U6217 (N_6217,N_4451,N_4181);
nand U6218 (N_6218,N_4867,N_4920);
nor U6219 (N_6219,N_3769,N_4486);
nand U6220 (N_6220,N_4570,N_3835);
and U6221 (N_6221,N_4423,N_4546);
nor U6222 (N_6222,N_4190,N_4669);
nand U6223 (N_6223,N_4944,N_4864);
xnor U6224 (N_6224,N_4727,N_3787);
nand U6225 (N_6225,N_4512,N_3845);
xor U6226 (N_6226,N_4235,N_3759);
and U6227 (N_6227,N_4036,N_4842);
nand U6228 (N_6228,N_4202,N_4922);
nand U6229 (N_6229,N_4244,N_3847);
nand U6230 (N_6230,N_4633,N_4990);
nand U6231 (N_6231,N_4141,N_3929);
or U6232 (N_6232,N_4651,N_4320);
xor U6233 (N_6233,N_4797,N_4155);
nand U6234 (N_6234,N_4563,N_4154);
nand U6235 (N_6235,N_4243,N_4297);
nor U6236 (N_6236,N_3858,N_4933);
nand U6237 (N_6237,N_4321,N_4546);
and U6238 (N_6238,N_4933,N_4308);
and U6239 (N_6239,N_3894,N_4301);
xnor U6240 (N_6240,N_4810,N_4150);
nor U6241 (N_6241,N_4599,N_4975);
xnor U6242 (N_6242,N_4099,N_4949);
xnor U6243 (N_6243,N_4512,N_4105);
xnor U6244 (N_6244,N_4810,N_4743);
nand U6245 (N_6245,N_3979,N_4997);
xor U6246 (N_6246,N_3945,N_4298);
and U6247 (N_6247,N_4160,N_4961);
nor U6248 (N_6248,N_3972,N_3894);
and U6249 (N_6249,N_4817,N_3951);
nor U6250 (N_6250,N_5089,N_5273);
and U6251 (N_6251,N_5969,N_5277);
or U6252 (N_6252,N_6143,N_5482);
xnor U6253 (N_6253,N_5788,N_5864);
nor U6254 (N_6254,N_5880,N_6166);
nand U6255 (N_6255,N_5096,N_5526);
nor U6256 (N_6256,N_5087,N_6065);
or U6257 (N_6257,N_5862,N_5955);
nor U6258 (N_6258,N_6035,N_5336);
or U6259 (N_6259,N_5030,N_6148);
nand U6260 (N_6260,N_5530,N_5324);
xor U6261 (N_6261,N_5619,N_5766);
nor U6262 (N_6262,N_5764,N_5114);
nand U6263 (N_6263,N_6144,N_6003);
or U6264 (N_6264,N_5537,N_5347);
and U6265 (N_6265,N_5940,N_5753);
nor U6266 (N_6266,N_5533,N_5255);
nor U6267 (N_6267,N_5228,N_5656);
nand U6268 (N_6268,N_5415,N_5933);
nor U6269 (N_6269,N_6170,N_5921);
nand U6270 (N_6270,N_5980,N_5232);
xor U6271 (N_6271,N_5399,N_5366);
nor U6272 (N_6272,N_5532,N_5683);
and U6273 (N_6273,N_5751,N_5131);
xor U6274 (N_6274,N_5496,N_5443);
and U6275 (N_6275,N_6234,N_6020);
nor U6276 (N_6276,N_5964,N_5538);
and U6277 (N_6277,N_5084,N_5598);
or U6278 (N_6278,N_5982,N_5298);
xnor U6279 (N_6279,N_5004,N_5739);
and U6280 (N_6280,N_5769,N_5717);
or U6281 (N_6281,N_5331,N_5781);
nor U6282 (N_6282,N_6088,N_5300);
nand U6283 (N_6283,N_6004,N_5219);
nor U6284 (N_6284,N_5989,N_5581);
nor U6285 (N_6285,N_5127,N_5514);
and U6286 (N_6286,N_5026,N_5041);
nor U6287 (N_6287,N_5077,N_5264);
and U6288 (N_6288,N_5066,N_5413);
and U6289 (N_6289,N_5835,N_5207);
or U6290 (N_6290,N_6069,N_5469);
xnor U6291 (N_6291,N_5216,N_5322);
or U6292 (N_6292,N_6089,N_6051);
xnor U6293 (N_6293,N_5525,N_5220);
xnor U6294 (N_6294,N_6197,N_6095);
xor U6295 (N_6295,N_5477,N_5950);
nor U6296 (N_6296,N_5328,N_6210);
nand U6297 (N_6297,N_6042,N_5463);
and U6298 (N_6298,N_5778,N_6019);
or U6299 (N_6299,N_5767,N_5777);
xor U6300 (N_6300,N_5897,N_5913);
and U6301 (N_6301,N_5222,N_5179);
nand U6302 (N_6302,N_5020,N_5544);
and U6303 (N_6303,N_5297,N_5224);
or U6304 (N_6304,N_5610,N_5899);
xnor U6305 (N_6305,N_5434,N_5887);
xnor U6306 (N_6306,N_5342,N_5947);
xor U6307 (N_6307,N_5461,N_5645);
nand U6308 (N_6308,N_5616,N_5652);
or U6309 (N_6309,N_6015,N_5249);
nand U6310 (N_6310,N_5548,N_5825);
nor U6311 (N_6311,N_6012,N_5573);
or U6312 (N_6312,N_6079,N_6192);
or U6313 (N_6313,N_5555,N_6081);
nand U6314 (N_6314,N_5569,N_5315);
and U6315 (N_6315,N_5350,N_5499);
or U6316 (N_6316,N_5626,N_6114);
and U6317 (N_6317,N_5786,N_6111);
xor U6318 (N_6318,N_5520,N_5170);
xor U6319 (N_6319,N_5810,N_5735);
or U6320 (N_6320,N_5870,N_5691);
and U6321 (N_6321,N_5775,N_5104);
nor U6322 (N_6322,N_5706,N_5577);
or U6323 (N_6323,N_5960,N_5922);
or U6324 (N_6324,N_5842,N_5100);
nor U6325 (N_6325,N_5423,N_5186);
nand U6326 (N_6326,N_5806,N_5043);
and U6327 (N_6327,N_5001,N_5572);
nand U6328 (N_6328,N_5325,N_6176);
nor U6329 (N_6329,N_5669,N_5408);
nand U6330 (N_6330,N_5741,N_5141);
nand U6331 (N_6331,N_6005,N_5385);
xnor U6332 (N_6332,N_5368,N_6185);
xnor U6333 (N_6333,N_5857,N_5896);
or U6334 (N_6334,N_5106,N_5283);
nand U6335 (N_6335,N_5303,N_5545);
or U6336 (N_6336,N_5090,N_5265);
xnor U6337 (N_6337,N_5789,N_5677);
nand U6338 (N_6338,N_5143,N_5830);
nor U6339 (N_6339,N_5190,N_5063);
nand U6340 (N_6340,N_5308,N_5245);
and U6341 (N_6341,N_5718,N_6094);
xor U6342 (N_6342,N_5177,N_5662);
and U6343 (N_6343,N_5985,N_6105);
or U6344 (N_6344,N_6242,N_5292);
nand U6345 (N_6345,N_5404,N_5396);
nor U6346 (N_6346,N_5348,N_6133);
xnor U6347 (N_6347,N_5681,N_5379);
or U6348 (N_6348,N_5754,N_5456);
nor U6349 (N_6349,N_5098,N_5097);
nor U6350 (N_6350,N_6075,N_5657);
xnor U6351 (N_6351,N_5807,N_6026);
xor U6352 (N_6352,N_5319,N_6092);
xnor U6353 (N_6353,N_5334,N_5129);
nand U6354 (N_6354,N_5266,N_6229);
nor U6355 (N_6355,N_5749,N_5972);
nor U6356 (N_6356,N_5450,N_6188);
or U6357 (N_6357,N_5402,N_5150);
nor U6358 (N_6358,N_5027,N_5258);
nor U6359 (N_6359,N_5172,N_5213);
nand U6360 (N_6360,N_5634,N_5631);
nand U6361 (N_6361,N_5990,N_5958);
xor U6362 (N_6362,N_5783,N_5798);
or U6363 (N_6363,N_5349,N_5279);
xor U6364 (N_6364,N_6097,N_5902);
nand U6365 (N_6365,N_5647,N_5765);
or U6366 (N_6366,N_5688,N_5802);
nor U6367 (N_6367,N_6039,N_5607);
and U6368 (N_6368,N_5863,N_6085);
or U6369 (N_6369,N_5409,N_5109);
and U6370 (N_6370,N_5966,N_5959);
or U6371 (N_6371,N_5113,N_5199);
xnor U6372 (N_6372,N_5497,N_6107);
nor U6373 (N_6373,N_5762,N_6189);
and U6374 (N_6374,N_5791,N_5554);
nand U6375 (N_6375,N_5108,N_6173);
nor U6376 (N_6376,N_5318,N_5794);
nand U6377 (N_6377,N_5163,N_5666);
xnor U6378 (N_6378,N_5246,N_5629);
and U6379 (N_6379,N_5422,N_5599);
nand U6380 (N_6380,N_5618,N_5917);
xnor U6381 (N_6381,N_5390,N_5296);
and U6382 (N_6382,N_5597,N_5595);
xnor U6383 (N_6383,N_5391,N_5589);
xor U6384 (N_6384,N_5214,N_5635);
xnor U6385 (N_6385,N_5949,N_5344);
xnor U6386 (N_6386,N_5551,N_6109);
xnor U6387 (N_6387,N_5035,N_6244);
and U6388 (N_6388,N_5784,N_5210);
and U6389 (N_6389,N_5543,N_5260);
nor U6390 (N_6390,N_5566,N_5375);
xnor U6391 (N_6391,N_5615,N_6016);
and U6392 (N_6392,N_5145,N_5281);
and U6393 (N_6393,N_6228,N_5903);
nand U6394 (N_6394,N_5800,N_5442);
nor U6395 (N_6395,N_5890,N_5871);
nor U6396 (N_6396,N_5481,N_5772);
xor U6397 (N_6397,N_5536,N_5604);
xnor U6398 (N_6398,N_5071,N_5091);
and U6399 (N_6399,N_6046,N_5130);
and U6400 (N_6400,N_5808,N_5371);
nor U6401 (N_6401,N_5837,N_5076);
nor U6402 (N_6402,N_5460,N_5665);
nor U6403 (N_6403,N_6168,N_5680);
and U6404 (N_6404,N_5813,N_5174);
and U6405 (N_6405,N_5011,N_6195);
nand U6406 (N_6406,N_5465,N_5875);
nand U6407 (N_6407,N_5736,N_5447);
or U6408 (N_6408,N_5354,N_5613);
nor U6409 (N_6409,N_5508,N_5419);
or U6410 (N_6410,N_5052,N_5291);
and U6411 (N_6411,N_5158,N_5242);
xnor U6412 (N_6412,N_5171,N_5016);
or U6413 (N_6413,N_5883,N_5998);
xor U6414 (N_6414,N_5564,N_6091);
or U6415 (N_6415,N_5528,N_5462);
or U6416 (N_6416,N_5254,N_5257);
nor U6417 (N_6417,N_5345,N_5702);
xor U6418 (N_6418,N_5911,N_5841);
nand U6419 (N_6419,N_5707,N_5086);
or U6420 (N_6420,N_5079,N_5648);
nand U6421 (N_6421,N_5005,N_5703);
xnor U6422 (N_6422,N_5042,N_5612);
or U6423 (N_6423,N_5023,N_5773);
nand U6424 (N_6424,N_5932,N_5164);
nor U6425 (N_6425,N_5259,N_5803);
and U6426 (N_6426,N_5485,N_6222);
xor U6427 (N_6427,N_5606,N_5776);
xnor U6428 (N_6428,N_5059,N_5270);
nor U6429 (N_6429,N_6231,N_5476);
and U6430 (N_6430,N_6093,N_5128);
and U6431 (N_6431,N_5963,N_6159);
nor U6432 (N_6432,N_6052,N_5760);
nand U6433 (N_6433,N_5819,N_6106);
or U6434 (N_6434,N_5301,N_5697);
or U6435 (N_6435,N_5834,N_5770);
or U6436 (N_6436,N_5268,N_5787);
nand U6437 (N_6437,N_5250,N_5748);
nand U6438 (N_6438,N_6078,N_6090);
or U6439 (N_6439,N_5256,N_5428);
nand U6440 (N_6440,N_6121,N_5455);
or U6441 (N_6441,N_5847,N_5844);
nand U6442 (N_6442,N_5021,N_5865);
or U6443 (N_6443,N_5209,N_5381);
xnor U6444 (N_6444,N_5727,N_5583);
nor U6445 (N_6445,N_5957,N_5248);
nand U6446 (N_6446,N_5335,N_5436);
or U6447 (N_6447,N_5869,N_6216);
nand U6448 (N_6448,N_5991,N_5173);
nor U6449 (N_6449,N_5487,N_6010);
nor U6450 (N_6450,N_6187,N_6021);
and U6451 (N_6451,N_6118,N_5686);
nor U6452 (N_6452,N_5660,N_5853);
or U6453 (N_6453,N_5523,N_5398);
nor U6454 (N_6454,N_5951,N_5439);
nor U6455 (N_6455,N_5643,N_5746);
nand U6456 (N_6456,N_5326,N_5653);
and U6457 (N_6457,N_6177,N_5527);
nor U6458 (N_6458,N_5198,N_6225);
xor U6459 (N_6459,N_6123,N_5912);
or U6460 (N_6460,N_5582,N_5008);
and U6461 (N_6461,N_5710,N_5230);
nand U6462 (N_6462,N_5305,N_6181);
nor U6463 (N_6463,N_5094,N_5571);
and U6464 (N_6464,N_5930,N_5699);
nor U6465 (N_6465,N_5509,N_5506);
and U6466 (N_6466,N_5738,N_5454);
or U6467 (N_6467,N_5970,N_5388);
nor U6468 (N_6468,N_6000,N_5983);
and U6469 (N_6469,N_5904,N_5049);
nand U6470 (N_6470,N_5067,N_5240);
and U6471 (N_6471,N_6041,N_5280);
and U6472 (N_6472,N_5229,N_5851);
nand U6473 (N_6473,N_6080,N_5411);
nor U6474 (N_6474,N_5360,N_6086);
nor U6475 (N_6475,N_5900,N_5977);
xnor U6476 (N_6476,N_5383,N_5441);
nand U6477 (N_6477,N_5032,N_5861);
and U6478 (N_6478,N_5155,N_5828);
or U6479 (N_6479,N_5467,N_6190);
nand U6480 (N_6480,N_5860,N_6066);
nor U6481 (N_6481,N_6014,N_6204);
or U6482 (N_6482,N_5640,N_5147);
xor U6483 (N_6483,N_5517,N_6217);
nor U6484 (N_6484,N_5473,N_5338);
nand U6485 (N_6485,N_6102,N_5797);
and U6486 (N_6486,N_5845,N_5948);
nand U6487 (N_6487,N_5663,N_5560);
nor U6488 (N_6488,N_5636,N_5483);
and U6489 (N_6489,N_5676,N_5457);
nor U6490 (N_6490,N_6165,N_5633);
or U6491 (N_6491,N_5251,N_5208);
xnor U6492 (N_6492,N_5568,N_5227);
nand U6493 (N_6493,N_5596,N_5723);
and U6494 (N_6494,N_5307,N_5472);
xnor U6495 (N_6495,N_5352,N_5805);
nand U6496 (N_6496,N_5642,N_6119);
or U6497 (N_6497,N_5387,N_5888);
and U6498 (N_6498,N_5124,N_5401);
and U6499 (N_6499,N_5015,N_6034);
xor U6500 (N_6500,N_5480,N_5866);
xor U6501 (N_6501,N_5695,N_5756);
nor U6502 (N_6502,N_5962,N_5361);
nor U6503 (N_6503,N_5092,N_5522);
or U6504 (N_6504,N_6202,N_5979);
and U6505 (N_6505,N_5012,N_5547);
xor U6506 (N_6506,N_5540,N_5563);
or U6507 (N_6507,N_5927,N_6226);
nor U6508 (N_6508,N_6221,N_6063);
and U6509 (N_6509,N_6156,N_5142);
xnor U6510 (N_6510,N_6076,N_5730);
and U6511 (N_6511,N_6136,N_5205);
nand U6512 (N_6512,N_6030,N_6215);
xnor U6513 (N_6513,N_5893,N_5272);
or U6514 (N_6514,N_5675,N_5639);
and U6515 (N_6515,N_5311,N_5859);
nor U6516 (N_6516,N_5673,N_5064);
or U6517 (N_6517,N_5057,N_5312);
xor U6518 (N_6518,N_5475,N_5484);
xor U6519 (N_6519,N_5918,N_5936);
or U6520 (N_6520,N_5116,N_6053);
and U6521 (N_6521,N_5693,N_5840);
nand U6522 (N_6522,N_6141,N_5849);
and U6523 (N_6523,N_6132,N_5894);
or U6524 (N_6524,N_5284,N_5341);
xor U6525 (N_6525,N_5356,N_5701);
and U6526 (N_6526,N_5202,N_6047);
xor U6527 (N_6527,N_5306,N_5045);
xnor U6528 (N_6528,N_5630,N_5346);
and U6529 (N_6529,N_5351,N_5855);
nand U6530 (N_6530,N_5121,N_6103);
nor U6531 (N_6531,N_5180,N_6083);
nand U6532 (N_6532,N_6201,N_5774);
or U6533 (N_6533,N_5720,N_5111);
nand U6534 (N_6534,N_6023,N_5987);
and U6535 (N_6535,N_5945,N_5430);
and U6536 (N_6536,N_5226,N_5734);
or U6537 (N_6537,N_5204,N_6087);
or U6538 (N_6538,N_5929,N_5287);
xnor U6539 (N_6539,N_5609,N_5363);
xnor U6540 (N_6540,N_5148,N_5567);
or U6541 (N_6541,N_5200,N_5617);
nand U6542 (N_6542,N_5793,N_5212);
nand U6543 (N_6543,N_5488,N_5188);
nor U6544 (N_6544,N_6218,N_5829);
and U6545 (N_6545,N_5556,N_5288);
nor U6546 (N_6546,N_6127,N_5992);
or U6547 (N_6547,N_5906,N_5167);
nor U6548 (N_6548,N_6011,N_6162);
xnor U6549 (N_6549,N_5275,N_5061);
xor U6550 (N_6550,N_5649,N_5625);
nand U6551 (N_6551,N_5073,N_6149);
xor U6552 (N_6552,N_5452,N_5494);
nand U6553 (N_6553,N_5037,N_5628);
xor U6554 (N_6554,N_5293,N_6050);
nand U6555 (N_6555,N_6163,N_5503);
or U6556 (N_6556,N_5575,N_6104);
and U6557 (N_6557,N_6057,N_5935);
xor U6558 (N_6558,N_6122,N_6008);
nand U6559 (N_6559,N_5974,N_5638);
xor U6560 (N_6560,N_5007,N_5490);
xnor U6561 (N_6561,N_5241,N_5996);
and U6562 (N_6562,N_5299,N_5003);
nor U6563 (N_6563,N_5584,N_5588);
or U6564 (N_6564,N_6224,N_5489);
and U6565 (N_6565,N_5574,N_5758);
nor U6566 (N_6566,N_5136,N_6214);
nor U6567 (N_6567,N_6174,N_5478);
nor U6568 (N_6568,N_6101,N_5211);
nand U6569 (N_6569,N_5608,N_5193);
xnor U6570 (N_6570,N_5981,N_6191);
and U6571 (N_6571,N_5901,N_6061);
xor U6572 (N_6572,N_5592,N_5759);
nand U6573 (N_6573,N_5047,N_5995);
nor U6574 (N_6574,N_5747,N_5197);
nor U6575 (N_6575,N_5337,N_5742);
xor U6576 (N_6576,N_5826,N_5185);
and U6577 (N_6577,N_5729,N_5040);
nor U6578 (N_6578,N_5892,N_5578);
or U6579 (N_6579,N_5750,N_6044);
nand U6580 (N_6580,N_5340,N_6245);
and U6581 (N_6581,N_5846,N_5785);
nand U6582 (N_6582,N_5919,N_5329);
xnor U6583 (N_6583,N_5426,N_5627);
xor U6584 (N_6584,N_5704,N_5101);
nor U6585 (N_6585,N_6045,N_5507);
nand U6586 (N_6586,N_5372,N_5054);
or U6587 (N_6587,N_5838,N_5967);
nand U6588 (N_6588,N_5491,N_6179);
nand U6589 (N_6589,N_5117,N_6152);
or U6590 (N_6590,N_5289,N_5420);
nand U6591 (N_6591,N_6233,N_5692);
and U6592 (N_6592,N_5394,N_5403);
and U6593 (N_6593,N_5370,N_5083);
or U6594 (N_6594,N_6058,N_5817);
nor U6595 (N_6595,N_6184,N_5144);
or U6596 (N_6596,N_5153,N_6055);
and U6597 (N_6597,N_5905,N_5939);
and U6598 (N_6598,N_5790,N_5237);
and U6599 (N_6599,N_5166,N_5058);
nand U6600 (N_6600,N_5429,N_5502);
and U6601 (N_6601,N_6002,N_5424);
and U6602 (N_6602,N_5586,N_6125);
and U6603 (N_6603,N_5558,N_5327);
xnor U6604 (N_6604,N_5668,N_5513);
and U6605 (N_6605,N_6198,N_5261);
nor U6606 (N_6606,N_6072,N_5884);
or U6607 (N_6607,N_5139,N_5024);
nor U6608 (N_6608,N_5392,N_5126);
and U6609 (N_6609,N_5602,N_5768);
nand U6610 (N_6610,N_5529,N_5986);
and U6611 (N_6611,N_5029,N_5238);
xnor U6612 (N_6612,N_6108,N_5938);
xnor U6613 (N_6613,N_5646,N_5889);
and U6614 (N_6614,N_5233,N_5362);
nand U6615 (N_6615,N_6112,N_5405);
nor U6616 (N_6616,N_5072,N_5438);
xnor U6617 (N_6617,N_5122,N_5470);
nand U6618 (N_6618,N_5601,N_5440);
and U6619 (N_6619,N_5715,N_5623);
nand U6620 (N_6620,N_6194,N_5731);
and U6621 (N_6621,N_6032,N_5009);
nor U6622 (N_6622,N_5843,N_6142);
and U6623 (N_6623,N_6017,N_5705);
nor U6624 (N_6624,N_5194,N_5816);
and U6625 (N_6625,N_5504,N_5377);
nor U6626 (N_6626,N_5570,N_5895);
xnor U6627 (N_6627,N_5085,N_5421);
and U6628 (N_6628,N_5169,N_6009);
nand U6629 (N_6629,N_5956,N_5874);
or U6630 (N_6630,N_5332,N_5234);
and U6631 (N_6631,N_5679,N_6200);
xnor U6632 (N_6632,N_6059,N_6182);
nor U6633 (N_6633,N_6161,N_5988);
or U6634 (N_6634,N_5965,N_5670);
nor U6635 (N_6635,N_5152,N_6138);
or U6636 (N_6636,N_5376,N_6237);
nor U6637 (N_6637,N_5358,N_5000);
or U6638 (N_6638,N_5278,N_6248);
or U6639 (N_6639,N_5831,N_6100);
xor U6640 (N_6640,N_6147,N_5565);
and U6641 (N_6641,N_5389,N_5809);
and U6642 (N_6642,N_5304,N_5282);
and U6643 (N_6643,N_5330,N_5053);
nand U6644 (N_6644,N_5678,N_5365);
nand U6645 (N_6645,N_6236,N_5812);
or U6646 (N_6646,N_6208,N_5294);
xor U6647 (N_6647,N_5682,N_6098);
nand U6648 (N_6648,N_5997,N_6212);
or U6649 (N_6649,N_5795,N_5269);
xnor U6650 (N_6650,N_5178,N_6130);
nor U6651 (N_6651,N_5407,N_5267);
nand U6652 (N_6652,N_5123,N_5068);
or U6653 (N_6653,N_5051,N_5740);
or U6654 (N_6654,N_5878,N_5290);
nor U6655 (N_6655,N_5039,N_5953);
and U6656 (N_6656,N_6169,N_5486);
nand U6657 (N_6657,N_5667,N_5822);
xor U6658 (N_6658,N_5309,N_5848);
or U6659 (N_6659,N_5175,N_5432);
and U6660 (N_6660,N_5780,N_5243);
or U6661 (N_6661,N_5712,N_5732);
xor U6662 (N_6662,N_5879,N_5120);
nand U6663 (N_6663,N_5215,N_5044);
or U6664 (N_6664,N_5685,N_5271);
and U6665 (N_6665,N_5135,N_5038);
and U6666 (N_6666,N_5414,N_5374);
and U6667 (N_6667,N_5909,N_5743);
xor U6668 (N_6668,N_5796,N_5709);
or U6669 (N_6669,N_5886,N_6180);
nor U6670 (N_6670,N_6211,N_5534);
or U6671 (N_6671,N_5952,N_6199);
nor U6672 (N_6672,N_5103,N_5553);
xnor U6673 (N_6673,N_5235,N_6232);
or U6674 (N_6674,N_5644,N_5873);
nor U6675 (N_6675,N_5713,N_5737);
xnor U6676 (N_6676,N_5659,N_6031);
or U6677 (N_6677,N_5446,N_5357);
or U6678 (N_6678,N_5632,N_5968);
and U6679 (N_6679,N_6247,N_5099);
and U6680 (N_6680,N_5343,N_5400);
xnor U6681 (N_6681,N_5060,N_5095);
and U6682 (N_6682,N_6064,N_6006);
or U6683 (N_6683,N_5431,N_6230);
and U6684 (N_6684,N_5065,N_6206);
or U6685 (N_6685,N_5002,N_5792);
xnor U6686 (N_6686,N_5195,N_5183);
nand U6687 (N_6687,N_5050,N_6220);
xnor U6688 (N_6688,N_5654,N_5125);
nor U6689 (N_6689,N_6082,N_5019);
xnor U6690 (N_6690,N_5074,N_5276);
and U6691 (N_6691,N_5923,N_6117);
and U6692 (N_6692,N_5105,N_5664);
and U6693 (N_6693,N_5833,N_5934);
nor U6694 (N_6694,N_5885,N_6239);
nand U6695 (N_6695,N_5725,N_5549);
xor U6696 (N_6696,N_5218,N_5317);
or U6697 (N_6697,N_6120,N_5752);
nor U6698 (N_6698,N_6223,N_5641);
xnor U6699 (N_6699,N_6209,N_6013);
nand U6700 (N_6700,N_5839,N_6193);
nand U6701 (N_6701,N_5165,N_5920);
nand U6702 (N_6702,N_5882,N_5433);
or U6703 (N_6703,N_5687,N_5852);
xnor U6704 (N_6704,N_5728,N_5262);
xor U6705 (N_6705,N_5811,N_5159);
nand U6706 (N_6706,N_5637,N_5468);
or U6707 (N_6707,N_6150,N_5316);
and U6708 (N_6708,N_5192,N_5321);
nand U6709 (N_6709,N_5191,N_5771);
or U6710 (N_6710,N_6207,N_5393);
nor U6711 (N_6711,N_5557,N_6060);
nand U6712 (N_6712,N_6196,N_5674);
nand U6713 (N_6713,N_5867,N_5926);
nor U6714 (N_6714,N_5661,N_6246);
and U6715 (N_6715,N_6157,N_6164);
and U6716 (N_6716,N_5263,N_5978);
xor U6717 (N_6717,N_6054,N_5355);
nor U6718 (N_6718,N_5445,N_6007);
nand U6719 (N_6719,N_5055,N_5444);
or U6720 (N_6720,N_6213,N_5132);
nor U6721 (N_6721,N_6022,N_5239);
nand U6722 (N_6722,N_5541,N_5138);
xnor U6723 (N_6723,N_5081,N_5658);
and U6724 (N_6724,N_6077,N_5711);
nand U6725 (N_6725,N_5417,N_5925);
nand U6726 (N_6726,N_5733,N_5196);
nand U6727 (N_6727,N_5600,N_5559);
nor U6728 (N_6728,N_5915,N_5611);
xnor U6729 (N_6729,N_5286,N_5217);
and U6730 (N_6730,N_5036,N_5236);
nand U6731 (N_6731,N_6186,N_5804);
or U6732 (N_6732,N_5156,N_5500);
nand U6733 (N_6733,N_5107,N_5546);
and U6734 (N_6734,N_5539,N_5999);
xnor U6735 (N_6735,N_5745,N_5189);
and U6736 (N_6736,N_5593,N_6096);
nor U6737 (N_6737,N_6145,N_5435);
and U6738 (N_6738,N_5062,N_5779);
xnor U6739 (N_6739,N_5689,N_5716);
xnor U6740 (N_6740,N_5118,N_5359);
and U6741 (N_6741,N_5512,N_5907);
nand U6742 (N_6742,N_6171,N_5157);
and U6743 (N_6743,N_6062,N_5302);
nor U6744 (N_6744,N_5994,N_5872);
nor U6745 (N_6745,N_5033,N_5585);
and U6746 (N_6746,N_5203,N_5594);
and U6747 (N_6747,N_5505,N_5914);
and U6748 (N_6748,N_5941,N_5562);
nor U6749 (N_6749,N_6074,N_5510);
and U6750 (N_6750,N_6018,N_6036);
and U6751 (N_6751,N_5910,N_5542);
nand U6752 (N_6752,N_5018,N_5201);
nor U6753 (N_6753,N_5069,N_5684);
or U6754 (N_6754,N_5724,N_5498);
and U6755 (N_6755,N_6158,N_5459);
nand U6756 (N_6756,N_5168,N_6240);
or U6757 (N_6757,N_6073,N_6033);
or U6758 (N_6758,N_6128,N_5620);
xnor U6759 (N_6759,N_5622,N_5943);
and U6760 (N_6760,N_6048,N_5624);
nand U6761 (N_6761,N_5561,N_5425);
nand U6762 (N_6762,N_5744,N_6160);
nor U6763 (N_6763,N_5088,N_5078);
xnor U6764 (N_6764,N_5453,N_6205);
nor U6765 (N_6765,N_5672,N_5149);
xnor U6766 (N_6766,N_5799,N_5333);
and U6767 (N_6767,N_6001,N_5418);
xnor U6768 (N_6768,N_5184,N_6028);
xor U6769 (N_6769,N_5821,N_5820);
nor U6770 (N_6770,N_6067,N_5782);
xor U6771 (N_6771,N_5877,N_5891);
and U6772 (N_6772,N_5976,N_5763);
xor U6773 (N_6773,N_5310,N_5605);
nand U6774 (N_6774,N_5550,N_5801);
nand U6775 (N_6775,N_5580,N_5836);
nor U6776 (N_6776,N_5493,N_5176);
nor U6777 (N_6777,N_5535,N_5367);
nand U6778 (N_6778,N_5722,N_5815);
xor U6779 (N_6779,N_5946,N_5876);
xor U6780 (N_6780,N_6238,N_5206);
xor U6781 (N_6781,N_5518,N_5590);
nand U6782 (N_6782,N_5295,N_5048);
nor U6783 (N_6783,N_5521,N_5231);
nand U6784 (N_6784,N_5515,N_5154);
nand U6785 (N_6785,N_6183,N_5591);
and U6786 (N_6786,N_5028,N_6124);
and U6787 (N_6787,N_5046,N_6131);
nor U6788 (N_6788,N_6135,N_5285);
or U6789 (N_6789,N_5942,N_5818);
nor U6790 (N_6790,N_5034,N_6155);
or U6791 (N_6791,N_5726,N_5552);
nor U6792 (N_6792,N_5961,N_5313);
or U6793 (N_6793,N_5971,N_5924);
xor U6794 (N_6794,N_6227,N_6025);
and U6795 (N_6795,N_5814,N_5524);
xnor U6796 (N_6796,N_5448,N_5244);
nor U6797 (N_6797,N_5146,N_5650);
nand U6798 (N_6798,N_6129,N_5380);
and U6799 (N_6799,N_5082,N_6137);
or U6800 (N_6800,N_5690,N_5093);
nor U6801 (N_6801,N_5519,N_5973);
xor U6802 (N_6802,N_6110,N_5908);
nor U6803 (N_6803,N_5451,N_5115);
and U6804 (N_6804,N_5579,N_5854);
and U6805 (N_6805,N_6115,N_5671);
nand U6806 (N_6806,N_6027,N_5339);
nor U6807 (N_6807,N_5576,N_6071);
xor U6808 (N_6808,N_5182,N_5110);
and U6809 (N_6809,N_5479,N_5993);
or U6810 (N_6810,N_6167,N_5651);
nor U6811 (N_6811,N_5373,N_5406);
nand U6812 (N_6812,N_5378,N_5931);
nor U6813 (N_6813,N_6024,N_6116);
nand U6814 (N_6814,N_5511,N_5603);
and U6815 (N_6815,N_5253,N_5025);
nor U6816 (N_6816,N_5832,N_6084);
and U6817 (N_6817,N_6235,N_6140);
nand U6818 (N_6818,N_5755,N_6175);
nand U6819 (N_6819,N_6203,N_5070);
or U6820 (N_6820,N_5382,N_5017);
and U6821 (N_6821,N_5464,N_6154);
nand U6822 (N_6822,N_5694,N_5162);
or U6823 (N_6823,N_5881,N_5274);
nor U6824 (N_6824,N_6040,N_5031);
and U6825 (N_6825,N_6029,N_5006);
nor U6826 (N_6826,N_5369,N_5856);
xnor U6827 (N_6827,N_5492,N_6151);
nand U6828 (N_6828,N_5700,N_5137);
and U6829 (N_6829,N_6172,N_5427);
and U6830 (N_6830,N_5187,N_6126);
xor U6831 (N_6831,N_5102,N_5410);
or U6832 (N_6832,N_5696,N_5868);
nor U6833 (N_6833,N_5471,N_5323);
or U6834 (N_6834,N_5621,N_5080);
xnor U6835 (N_6835,N_5698,N_5181);
and U6836 (N_6836,N_5824,N_6068);
or U6837 (N_6837,N_5353,N_5161);
nand U6838 (N_6838,N_5221,N_5655);
xnor U6839 (N_6839,N_6049,N_5140);
nor U6840 (N_6840,N_5761,N_5412);
xor U6841 (N_6841,N_6113,N_5714);
nor U6842 (N_6842,N_5134,N_5397);
xor U6843 (N_6843,N_5010,N_5858);
nor U6844 (N_6844,N_5928,N_5013);
nor U6845 (N_6845,N_6070,N_5151);
xnor U6846 (N_6846,N_6056,N_5364);
and U6847 (N_6847,N_5850,N_5133);
xnor U6848 (N_6848,N_5056,N_5247);
and U6849 (N_6849,N_6038,N_5721);
nor U6850 (N_6850,N_5014,N_5937);
or U6851 (N_6851,N_5898,N_6219);
nor U6852 (N_6852,N_5501,N_5386);
and U6853 (N_6853,N_5719,N_6243);
or U6854 (N_6854,N_5827,N_6043);
nand U6855 (N_6855,N_5416,N_6249);
and U6856 (N_6856,N_6037,N_6139);
nor U6857 (N_6857,N_5516,N_5075);
nand U6858 (N_6858,N_6153,N_5954);
nor U6859 (N_6859,N_5466,N_5223);
nand U6860 (N_6860,N_5395,N_6178);
and U6861 (N_6861,N_5225,N_5252);
or U6862 (N_6862,N_5449,N_5320);
xor U6863 (N_6863,N_5916,N_5384);
nand U6864 (N_6864,N_5474,N_5119);
xor U6865 (N_6865,N_6099,N_5495);
nand U6866 (N_6866,N_5531,N_5823);
and U6867 (N_6867,N_5314,N_5437);
and U6868 (N_6868,N_6241,N_5984);
nor U6869 (N_6869,N_5112,N_6146);
xor U6870 (N_6870,N_5944,N_6134);
nor U6871 (N_6871,N_5587,N_5708);
and U6872 (N_6872,N_5458,N_5022);
nand U6873 (N_6873,N_5975,N_5614);
and U6874 (N_6874,N_5757,N_5160);
and U6875 (N_6875,N_5263,N_5220);
or U6876 (N_6876,N_5133,N_5228);
xor U6877 (N_6877,N_5210,N_6035);
nand U6878 (N_6878,N_5477,N_5926);
and U6879 (N_6879,N_5703,N_5597);
and U6880 (N_6880,N_5654,N_5986);
and U6881 (N_6881,N_6155,N_6068);
nand U6882 (N_6882,N_5883,N_5723);
nand U6883 (N_6883,N_5911,N_5021);
nor U6884 (N_6884,N_5980,N_5890);
nor U6885 (N_6885,N_5287,N_5133);
nor U6886 (N_6886,N_6203,N_5999);
xnor U6887 (N_6887,N_6175,N_5001);
nor U6888 (N_6888,N_5742,N_5621);
or U6889 (N_6889,N_5313,N_5775);
xor U6890 (N_6890,N_6056,N_6095);
and U6891 (N_6891,N_5367,N_5884);
nor U6892 (N_6892,N_6119,N_5052);
or U6893 (N_6893,N_6040,N_5653);
or U6894 (N_6894,N_5427,N_5560);
xor U6895 (N_6895,N_5063,N_5007);
xor U6896 (N_6896,N_5308,N_5613);
or U6897 (N_6897,N_5034,N_5368);
or U6898 (N_6898,N_6231,N_5906);
xor U6899 (N_6899,N_5310,N_5688);
or U6900 (N_6900,N_6078,N_5119);
or U6901 (N_6901,N_6114,N_5444);
nor U6902 (N_6902,N_5992,N_5630);
nor U6903 (N_6903,N_5634,N_5465);
nor U6904 (N_6904,N_5519,N_5816);
and U6905 (N_6905,N_6193,N_5535);
or U6906 (N_6906,N_6013,N_6226);
and U6907 (N_6907,N_5937,N_6187);
nand U6908 (N_6908,N_5452,N_5083);
xor U6909 (N_6909,N_5776,N_6213);
xnor U6910 (N_6910,N_5870,N_5784);
nor U6911 (N_6911,N_6041,N_5303);
or U6912 (N_6912,N_5246,N_6065);
nand U6913 (N_6913,N_5744,N_5331);
and U6914 (N_6914,N_6034,N_5781);
and U6915 (N_6915,N_5443,N_5737);
nor U6916 (N_6916,N_5719,N_5912);
and U6917 (N_6917,N_5920,N_5158);
nand U6918 (N_6918,N_6130,N_5233);
and U6919 (N_6919,N_5997,N_5817);
nand U6920 (N_6920,N_5754,N_5104);
nand U6921 (N_6921,N_5004,N_6176);
and U6922 (N_6922,N_5192,N_5241);
nand U6923 (N_6923,N_6231,N_5795);
xnor U6924 (N_6924,N_6131,N_5943);
nor U6925 (N_6925,N_5630,N_5749);
or U6926 (N_6926,N_5617,N_5368);
and U6927 (N_6927,N_6026,N_5704);
nor U6928 (N_6928,N_6041,N_5663);
xor U6929 (N_6929,N_5795,N_5458);
nor U6930 (N_6930,N_5671,N_5503);
nor U6931 (N_6931,N_5367,N_5292);
nor U6932 (N_6932,N_5501,N_5801);
xnor U6933 (N_6933,N_6020,N_5209);
nand U6934 (N_6934,N_5517,N_5869);
or U6935 (N_6935,N_5476,N_5765);
and U6936 (N_6936,N_5549,N_5319);
and U6937 (N_6937,N_6036,N_5858);
xnor U6938 (N_6938,N_5303,N_5406);
xnor U6939 (N_6939,N_5475,N_5426);
or U6940 (N_6940,N_6058,N_5201);
nand U6941 (N_6941,N_5238,N_5090);
or U6942 (N_6942,N_5329,N_6211);
nor U6943 (N_6943,N_5815,N_5617);
or U6944 (N_6944,N_6132,N_5522);
or U6945 (N_6945,N_5731,N_5462);
and U6946 (N_6946,N_5525,N_5762);
and U6947 (N_6947,N_5266,N_5192);
and U6948 (N_6948,N_5839,N_5314);
nor U6949 (N_6949,N_5321,N_5547);
and U6950 (N_6950,N_5059,N_5374);
xor U6951 (N_6951,N_5104,N_5646);
nor U6952 (N_6952,N_5443,N_5675);
or U6953 (N_6953,N_6099,N_5873);
nor U6954 (N_6954,N_5446,N_5511);
or U6955 (N_6955,N_5986,N_5000);
nand U6956 (N_6956,N_5104,N_5767);
xnor U6957 (N_6957,N_5930,N_5408);
nor U6958 (N_6958,N_5825,N_6127);
nor U6959 (N_6959,N_5962,N_5261);
nand U6960 (N_6960,N_5336,N_5308);
and U6961 (N_6961,N_5083,N_5369);
and U6962 (N_6962,N_5645,N_5332);
nand U6963 (N_6963,N_5080,N_5920);
and U6964 (N_6964,N_5482,N_5962);
or U6965 (N_6965,N_5456,N_5918);
nand U6966 (N_6966,N_5471,N_5880);
nand U6967 (N_6967,N_5046,N_5652);
xnor U6968 (N_6968,N_5956,N_6090);
and U6969 (N_6969,N_5430,N_6019);
nand U6970 (N_6970,N_5020,N_5819);
nand U6971 (N_6971,N_5927,N_6175);
and U6972 (N_6972,N_6028,N_5121);
and U6973 (N_6973,N_5033,N_6191);
and U6974 (N_6974,N_6157,N_6125);
nand U6975 (N_6975,N_5576,N_5714);
nor U6976 (N_6976,N_5660,N_5061);
nor U6977 (N_6977,N_5993,N_5833);
or U6978 (N_6978,N_6168,N_5057);
xnor U6979 (N_6979,N_5024,N_6165);
nor U6980 (N_6980,N_6017,N_5452);
nand U6981 (N_6981,N_5224,N_5552);
nor U6982 (N_6982,N_5953,N_5234);
nand U6983 (N_6983,N_5359,N_5232);
xor U6984 (N_6984,N_5005,N_5277);
or U6985 (N_6985,N_5479,N_6208);
or U6986 (N_6986,N_5753,N_5034);
xnor U6987 (N_6987,N_5180,N_5066);
and U6988 (N_6988,N_5343,N_6050);
or U6989 (N_6989,N_5461,N_5283);
and U6990 (N_6990,N_5876,N_5232);
and U6991 (N_6991,N_5770,N_5267);
nor U6992 (N_6992,N_5386,N_6140);
or U6993 (N_6993,N_5772,N_5192);
nor U6994 (N_6994,N_6039,N_5148);
xor U6995 (N_6995,N_5961,N_5549);
and U6996 (N_6996,N_6193,N_5645);
and U6997 (N_6997,N_5495,N_6220);
xnor U6998 (N_6998,N_5730,N_5865);
nand U6999 (N_6999,N_6151,N_5673);
nand U7000 (N_7000,N_6040,N_6153);
nor U7001 (N_7001,N_5558,N_5078);
or U7002 (N_7002,N_5840,N_6014);
nor U7003 (N_7003,N_5179,N_5022);
xor U7004 (N_7004,N_5711,N_5822);
and U7005 (N_7005,N_5867,N_5825);
and U7006 (N_7006,N_5167,N_5490);
nand U7007 (N_7007,N_5709,N_5043);
and U7008 (N_7008,N_5830,N_5365);
or U7009 (N_7009,N_5287,N_5088);
xor U7010 (N_7010,N_5498,N_5234);
or U7011 (N_7011,N_5046,N_5149);
nor U7012 (N_7012,N_5314,N_6043);
nand U7013 (N_7013,N_5898,N_5975);
xnor U7014 (N_7014,N_5320,N_6241);
or U7015 (N_7015,N_5063,N_5409);
or U7016 (N_7016,N_5585,N_5311);
or U7017 (N_7017,N_5924,N_5262);
xor U7018 (N_7018,N_6161,N_5570);
nand U7019 (N_7019,N_5292,N_5418);
and U7020 (N_7020,N_5457,N_5288);
nor U7021 (N_7021,N_5674,N_5238);
nand U7022 (N_7022,N_6183,N_5708);
nor U7023 (N_7023,N_5691,N_5190);
nor U7024 (N_7024,N_5866,N_5104);
xor U7025 (N_7025,N_6161,N_6114);
nand U7026 (N_7026,N_5279,N_6195);
nand U7027 (N_7027,N_5241,N_5395);
nor U7028 (N_7028,N_6084,N_5845);
nand U7029 (N_7029,N_5719,N_5694);
and U7030 (N_7030,N_5031,N_6036);
xor U7031 (N_7031,N_5808,N_5265);
and U7032 (N_7032,N_5335,N_5452);
nand U7033 (N_7033,N_5754,N_6108);
or U7034 (N_7034,N_5540,N_5119);
and U7035 (N_7035,N_5038,N_5295);
and U7036 (N_7036,N_5304,N_6189);
nand U7037 (N_7037,N_5049,N_6124);
xnor U7038 (N_7038,N_6052,N_5814);
nand U7039 (N_7039,N_5739,N_5094);
and U7040 (N_7040,N_5236,N_5642);
nor U7041 (N_7041,N_5214,N_5436);
xor U7042 (N_7042,N_5337,N_5494);
nand U7043 (N_7043,N_5914,N_5625);
nand U7044 (N_7044,N_5558,N_5344);
or U7045 (N_7045,N_5944,N_5715);
or U7046 (N_7046,N_5273,N_5002);
nand U7047 (N_7047,N_5240,N_5929);
nor U7048 (N_7048,N_5290,N_5924);
xnor U7049 (N_7049,N_5246,N_5938);
nand U7050 (N_7050,N_5645,N_5368);
xor U7051 (N_7051,N_5639,N_6164);
or U7052 (N_7052,N_6120,N_5250);
nor U7053 (N_7053,N_5030,N_5557);
nor U7054 (N_7054,N_5857,N_5024);
nand U7055 (N_7055,N_5718,N_5954);
or U7056 (N_7056,N_5392,N_6161);
xnor U7057 (N_7057,N_5869,N_5748);
xnor U7058 (N_7058,N_5218,N_5292);
and U7059 (N_7059,N_5119,N_6060);
xnor U7060 (N_7060,N_6108,N_5855);
nand U7061 (N_7061,N_5445,N_5899);
nand U7062 (N_7062,N_6240,N_5205);
xor U7063 (N_7063,N_5093,N_5718);
and U7064 (N_7064,N_5278,N_5921);
or U7065 (N_7065,N_5851,N_5883);
and U7066 (N_7066,N_6032,N_5877);
and U7067 (N_7067,N_5374,N_6226);
or U7068 (N_7068,N_5520,N_5200);
nand U7069 (N_7069,N_5241,N_6181);
and U7070 (N_7070,N_5679,N_5072);
and U7071 (N_7071,N_6076,N_5812);
nor U7072 (N_7072,N_5207,N_6083);
and U7073 (N_7073,N_6086,N_6018);
nor U7074 (N_7074,N_5726,N_6190);
or U7075 (N_7075,N_6234,N_6047);
nand U7076 (N_7076,N_5710,N_5930);
xor U7077 (N_7077,N_5832,N_5203);
nor U7078 (N_7078,N_5738,N_5810);
xor U7079 (N_7079,N_5535,N_5464);
xor U7080 (N_7080,N_5889,N_5538);
nand U7081 (N_7081,N_6237,N_6171);
nand U7082 (N_7082,N_5688,N_6028);
and U7083 (N_7083,N_6038,N_5106);
xnor U7084 (N_7084,N_5379,N_6050);
or U7085 (N_7085,N_5158,N_6079);
nor U7086 (N_7086,N_5829,N_5134);
xor U7087 (N_7087,N_5391,N_6071);
nand U7088 (N_7088,N_6109,N_6091);
or U7089 (N_7089,N_5665,N_5245);
and U7090 (N_7090,N_6129,N_5442);
nand U7091 (N_7091,N_5285,N_5012);
xnor U7092 (N_7092,N_5344,N_5042);
xnor U7093 (N_7093,N_5025,N_6136);
or U7094 (N_7094,N_5446,N_5309);
and U7095 (N_7095,N_5397,N_5524);
and U7096 (N_7096,N_5396,N_5403);
or U7097 (N_7097,N_5248,N_6122);
and U7098 (N_7098,N_5354,N_5829);
nand U7099 (N_7099,N_6135,N_5606);
or U7100 (N_7100,N_5142,N_5078);
nor U7101 (N_7101,N_6217,N_6247);
nand U7102 (N_7102,N_5393,N_5379);
or U7103 (N_7103,N_5742,N_6167);
nand U7104 (N_7104,N_5531,N_5600);
or U7105 (N_7105,N_6225,N_5388);
nor U7106 (N_7106,N_5653,N_5575);
nand U7107 (N_7107,N_5613,N_5187);
nor U7108 (N_7108,N_5163,N_5609);
or U7109 (N_7109,N_5344,N_5268);
nand U7110 (N_7110,N_6160,N_5698);
or U7111 (N_7111,N_6155,N_5011);
nand U7112 (N_7112,N_5699,N_6091);
nor U7113 (N_7113,N_6079,N_6107);
nand U7114 (N_7114,N_5876,N_5014);
nor U7115 (N_7115,N_5651,N_5660);
xnor U7116 (N_7116,N_5412,N_5305);
nor U7117 (N_7117,N_5212,N_6094);
or U7118 (N_7118,N_5519,N_5758);
or U7119 (N_7119,N_6206,N_6181);
and U7120 (N_7120,N_5058,N_5576);
and U7121 (N_7121,N_5523,N_6022);
xor U7122 (N_7122,N_5701,N_5287);
nand U7123 (N_7123,N_6109,N_5989);
nor U7124 (N_7124,N_5603,N_5461);
nand U7125 (N_7125,N_5887,N_5214);
or U7126 (N_7126,N_6080,N_6039);
and U7127 (N_7127,N_5904,N_5362);
or U7128 (N_7128,N_5037,N_5020);
or U7129 (N_7129,N_5704,N_5830);
nand U7130 (N_7130,N_5236,N_6171);
or U7131 (N_7131,N_5263,N_5611);
nor U7132 (N_7132,N_6212,N_5110);
xnor U7133 (N_7133,N_5542,N_5493);
nand U7134 (N_7134,N_5272,N_5448);
and U7135 (N_7135,N_6020,N_5760);
and U7136 (N_7136,N_5911,N_5538);
nand U7137 (N_7137,N_6092,N_5053);
or U7138 (N_7138,N_5722,N_6187);
or U7139 (N_7139,N_5261,N_5297);
nand U7140 (N_7140,N_5007,N_5629);
nand U7141 (N_7141,N_5126,N_5681);
nand U7142 (N_7142,N_6017,N_5420);
or U7143 (N_7143,N_5917,N_6045);
xor U7144 (N_7144,N_5051,N_5796);
or U7145 (N_7145,N_6130,N_5830);
xor U7146 (N_7146,N_5312,N_5408);
nor U7147 (N_7147,N_5524,N_5823);
or U7148 (N_7148,N_5226,N_5097);
nand U7149 (N_7149,N_6237,N_6153);
xor U7150 (N_7150,N_5460,N_6005);
nor U7151 (N_7151,N_5109,N_5435);
nor U7152 (N_7152,N_5873,N_5745);
nand U7153 (N_7153,N_6111,N_5190);
or U7154 (N_7154,N_6106,N_5888);
and U7155 (N_7155,N_5107,N_5552);
xnor U7156 (N_7156,N_5031,N_6209);
nand U7157 (N_7157,N_5409,N_5981);
nor U7158 (N_7158,N_5578,N_5842);
xnor U7159 (N_7159,N_5906,N_5424);
nand U7160 (N_7160,N_5549,N_5639);
nor U7161 (N_7161,N_5790,N_6009);
xor U7162 (N_7162,N_5974,N_5036);
xor U7163 (N_7163,N_5454,N_5594);
nand U7164 (N_7164,N_5447,N_5619);
and U7165 (N_7165,N_5406,N_5221);
xnor U7166 (N_7166,N_5901,N_5667);
nor U7167 (N_7167,N_6218,N_5971);
xor U7168 (N_7168,N_5867,N_5740);
nor U7169 (N_7169,N_5827,N_5151);
nand U7170 (N_7170,N_5156,N_5556);
and U7171 (N_7171,N_5775,N_5203);
and U7172 (N_7172,N_5077,N_6145);
or U7173 (N_7173,N_6172,N_5974);
or U7174 (N_7174,N_5399,N_6010);
or U7175 (N_7175,N_5649,N_6175);
and U7176 (N_7176,N_5442,N_5627);
xor U7177 (N_7177,N_5796,N_5625);
or U7178 (N_7178,N_6188,N_5092);
nor U7179 (N_7179,N_5551,N_5320);
xor U7180 (N_7180,N_5728,N_5575);
xor U7181 (N_7181,N_5845,N_5120);
and U7182 (N_7182,N_6188,N_5023);
and U7183 (N_7183,N_6110,N_6243);
or U7184 (N_7184,N_5100,N_5376);
and U7185 (N_7185,N_5238,N_5524);
nor U7186 (N_7186,N_6184,N_5187);
nand U7187 (N_7187,N_5950,N_5249);
and U7188 (N_7188,N_5024,N_5429);
nand U7189 (N_7189,N_5608,N_5819);
or U7190 (N_7190,N_5143,N_6247);
or U7191 (N_7191,N_5313,N_6075);
or U7192 (N_7192,N_6214,N_5133);
nor U7193 (N_7193,N_5059,N_5265);
nand U7194 (N_7194,N_5853,N_5006);
or U7195 (N_7195,N_5199,N_5105);
nand U7196 (N_7196,N_5343,N_5827);
xor U7197 (N_7197,N_5119,N_5020);
xor U7198 (N_7198,N_6093,N_6198);
nand U7199 (N_7199,N_5992,N_5467);
nand U7200 (N_7200,N_5604,N_6129);
xnor U7201 (N_7201,N_5089,N_5263);
and U7202 (N_7202,N_5036,N_5691);
nor U7203 (N_7203,N_5875,N_5870);
nor U7204 (N_7204,N_6002,N_6227);
nand U7205 (N_7205,N_5077,N_5530);
or U7206 (N_7206,N_5153,N_5745);
nor U7207 (N_7207,N_5545,N_6156);
nand U7208 (N_7208,N_5430,N_5136);
or U7209 (N_7209,N_5598,N_5936);
nor U7210 (N_7210,N_5212,N_5121);
nor U7211 (N_7211,N_5350,N_5821);
or U7212 (N_7212,N_6050,N_6185);
and U7213 (N_7213,N_5272,N_5490);
and U7214 (N_7214,N_5252,N_6052);
and U7215 (N_7215,N_5969,N_5350);
or U7216 (N_7216,N_5727,N_5887);
and U7217 (N_7217,N_5835,N_5857);
or U7218 (N_7218,N_6067,N_5956);
and U7219 (N_7219,N_5833,N_5182);
xnor U7220 (N_7220,N_5922,N_6048);
nor U7221 (N_7221,N_6008,N_5123);
or U7222 (N_7222,N_5812,N_5116);
and U7223 (N_7223,N_5036,N_5530);
nand U7224 (N_7224,N_5250,N_5826);
and U7225 (N_7225,N_6084,N_5239);
or U7226 (N_7226,N_5924,N_5784);
or U7227 (N_7227,N_5189,N_5081);
nand U7228 (N_7228,N_5632,N_5709);
nor U7229 (N_7229,N_5598,N_5810);
and U7230 (N_7230,N_5427,N_5021);
xnor U7231 (N_7231,N_5199,N_6100);
or U7232 (N_7232,N_5882,N_5239);
or U7233 (N_7233,N_5294,N_5502);
or U7234 (N_7234,N_5907,N_6101);
nand U7235 (N_7235,N_6245,N_5663);
xnor U7236 (N_7236,N_6199,N_5212);
xnor U7237 (N_7237,N_5388,N_5553);
nand U7238 (N_7238,N_5970,N_5161);
nand U7239 (N_7239,N_5834,N_5753);
and U7240 (N_7240,N_5938,N_5061);
nor U7241 (N_7241,N_6006,N_5672);
nand U7242 (N_7242,N_5918,N_5636);
and U7243 (N_7243,N_5936,N_5422);
and U7244 (N_7244,N_6034,N_5345);
nor U7245 (N_7245,N_5490,N_5997);
or U7246 (N_7246,N_5077,N_5512);
or U7247 (N_7247,N_5222,N_5635);
xnor U7248 (N_7248,N_5773,N_5615);
or U7249 (N_7249,N_5410,N_5840);
xor U7250 (N_7250,N_5834,N_5867);
nand U7251 (N_7251,N_6230,N_5995);
xor U7252 (N_7252,N_5106,N_5907);
nor U7253 (N_7253,N_5032,N_5463);
and U7254 (N_7254,N_5199,N_5364);
nor U7255 (N_7255,N_5908,N_5791);
xnor U7256 (N_7256,N_5289,N_5271);
nor U7257 (N_7257,N_5690,N_5883);
xor U7258 (N_7258,N_6183,N_5875);
nor U7259 (N_7259,N_5596,N_5923);
xor U7260 (N_7260,N_5577,N_5264);
xnor U7261 (N_7261,N_5453,N_6075);
xnor U7262 (N_7262,N_5992,N_5291);
nand U7263 (N_7263,N_5519,N_5769);
xnor U7264 (N_7264,N_6205,N_5983);
nand U7265 (N_7265,N_6130,N_6241);
nor U7266 (N_7266,N_5252,N_6240);
xor U7267 (N_7267,N_5828,N_5975);
nor U7268 (N_7268,N_5524,N_5288);
xnor U7269 (N_7269,N_5798,N_5394);
xnor U7270 (N_7270,N_5664,N_5405);
or U7271 (N_7271,N_5799,N_6143);
nor U7272 (N_7272,N_5542,N_6076);
nor U7273 (N_7273,N_5904,N_5650);
nand U7274 (N_7274,N_5313,N_5205);
and U7275 (N_7275,N_5664,N_5559);
nor U7276 (N_7276,N_5868,N_5007);
nand U7277 (N_7277,N_6187,N_5351);
nor U7278 (N_7278,N_5690,N_5083);
nand U7279 (N_7279,N_6059,N_5203);
nand U7280 (N_7280,N_6087,N_6011);
and U7281 (N_7281,N_5662,N_5335);
nand U7282 (N_7282,N_5863,N_6022);
or U7283 (N_7283,N_5474,N_5764);
xnor U7284 (N_7284,N_5892,N_6011);
and U7285 (N_7285,N_5391,N_5877);
nand U7286 (N_7286,N_6084,N_5541);
or U7287 (N_7287,N_5237,N_5658);
or U7288 (N_7288,N_5757,N_5145);
xor U7289 (N_7289,N_6014,N_5375);
or U7290 (N_7290,N_5126,N_6188);
nand U7291 (N_7291,N_5436,N_5863);
and U7292 (N_7292,N_5799,N_5376);
nor U7293 (N_7293,N_6135,N_5085);
xor U7294 (N_7294,N_5641,N_5108);
xor U7295 (N_7295,N_6240,N_5361);
and U7296 (N_7296,N_5462,N_5466);
nand U7297 (N_7297,N_6055,N_5040);
xnor U7298 (N_7298,N_5038,N_5588);
or U7299 (N_7299,N_5894,N_5612);
nand U7300 (N_7300,N_5134,N_5316);
or U7301 (N_7301,N_5431,N_5800);
nand U7302 (N_7302,N_5046,N_6090);
or U7303 (N_7303,N_5849,N_5587);
xor U7304 (N_7304,N_5164,N_5928);
nand U7305 (N_7305,N_6114,N_6109);
and U7306 (N_7306,N_5514,N_6069);
nor U7307 (N_7307,N_5954,N_5590);
nor U7308 (N_7308,N_5456,N_6038);
nand U7309 (N_7309,N_5579,N_5803);
xor U7310 (N_7310,N_5831,N_5311);
and U7311 (N_7311,N_6233,N_5908);
nor U7312 (N_7312,N_5960,N_5611);
and U7313 (N_7313,N_5451,N_6193);
and U7314 (N_7314,N_5379,N_5501);
nor U7315 (N_7315,N_5396,N_5108);
and U7316 (N_7316,N_5578,N_5633);
xor U7317 (N_7317,N_5744,N_5722);
or U7318 (N_7318,N_5172,N_5776);
xnor U7319 (N_7319,N_5061,N_5575);
and U7320 (N_7320,N_6214,N_5450);
nand U7321 (N_7321,N_5542,N_5154);
nor U7322 (N_7322,N_5873,N_5747);
xor U7323 (N_7323,N_6248,N_5640);
nand U7324 (N_7324,N_5498,N_5079);
nand U7325 (N_7325,N_5270,N_6171);
nand U7326 (N_7326,N_5108,N_5861);
xnor U7327 (N_7327,N_6184,N_6225);
nand U7328 (N_7328,N_5415,N_5262);
xor U7329 (N_7329,N_5191,N_5468);
nor U7330 (N_7330,N_5035,N_5085);
nand U7331 (N_7331,N_5021,N_5371);
nand U7332 (N_7332,N_6135,N_5403);
nand U7333 (N_7333,N_6091,N_5663);
or U7334 (N_7334,N_5824,N_5804);
xnor U7335 (N_7335,N_5122,N_5144);
nor U7336 (N_7336,N_6021,N_5420);
or U7337 (N_7337,N_5991,N_5261);
or U7338 (N_7338,N_5988,N_5264);
or U7339 (N_7339,N_5952,N_5895);
and U7340 (N_7340,N_5811,N_5496);
nor U7341 (N_7341,N_6152,N_5065);
and U7342 (N_7342,N_5248,N_5360);
xnor U7343 (N_7343,N_5988,N_5068);
nor U7344 (N_7344,N_5818,N_6077);
nor U7345 (N_7345,N_5253,N_5221);
nor U7346 (N_7346,N_5332,N_6001);
xnor U7347 (N_7347,N_5607,N_5442);
and U7348 (N_7348,N_5559,N_5037);
nor U7349 (N_7349,N_5712,N_5430);
or U7350 (N_7350,N_5394,N_5559);
nor U7351 (N_7351,N_5470,N_5513);
xnor U7352 (N_7352,N_5120,N_5645);
nor U7353 (N_7353,N_6221,N_5646);
or U7354 (N_7354,N_5911,N_5338);
and U7355 (N_7355,N_5668,N_5720);
or U7356 (N_7356,N_6164,N_5245);
nand U7357 (N_7357,N_5399,N_5735);
nand U7358 (N_7358,N_5977,N_5523);
and U7359 (N_7359,N_5637,N_5526);
and U7360 (N_7360,N_6102,N_5915);
xnor U7361 (N_7361,N_6132,N_5472);
nand U7362 (N_7362,N_6013,N_5786);
or U7363 (N_7363,N_6088,N_6123);
xnor U7364 (N_7364,N_5624,N_5027);
nand U7365 (N_7365,N_5437,N_6222);
nand U7366 (N_7366,N_5955,N_5850);
xnor U7367 (N_7367,N_5166,N_5671);
nor U7368 (N_7368,N_5059,N_6062);
nand U7369 (N_7369,N_5664,N_5686);
or U7370 (N_7370,N_5142,N_6030);
nor U7371 (N_7371,N_5167,N_5697);
nand U7372 (N_7372,N_5208,N_6106);
xor U7373 (N_7373,N_5768,N_5291);
xor U7374 (N_7374,N_6179,N_5022);
nor U7375 (N_7375,N_6124,N_5326);
or U7376 (N_7376,N_5530,N_6207);
xor U7377 (N_7377,N_5902,N_5446);
and U7378 (N_7378,N_5467,N_5600);
or U7379 (N_7379,N_5701,N_6154);
and U7380 (N_7380,N_5184,N_5881);
xor U7381 (N_7381,N_5549,N_5270);
nand U7382 (N_7382,N_6114,N_6218);
and U7383 (N_7383,N_5104,N_6155);
xnor U7384 (N_7384,N_5876,N_5416);
or U7385 (N_7385,N_5189,N_5713);
and U7386 (N_7386,N_5753,N_5416);
xor U7387 (N_7387,N_5814,N_6230);
xnor U7388 (N_7388,N_5238,N_5272);
nand U7389 (N_7389,N_5695,N_5340);
xor U7390 (N_7390,N_5029,N_5970);
and U7391 (N_7391,N_5291,N_5951);
or U7392 (N_7392,N_6010,N_5761);
nand U7393 (N_7393,N_5900,N_5211);
nor U7394 (N_7394,N_5312,N_5097);
xnor U7395 (N_7395,N_5319,N_5256);
and U7396 (N_7396,N_6102,N_5374);
nor U7397 (N_7397,N_5499,N_6187);
or U7398 (N_7398,N_5887,N_5682);
nand U7399 (N_7399,N_5180,N_5283);
or U7400 (N_7400,N_5528,N_5793);
xnor U7401 (N_7401,N_6001,N_6011);
nor U7402 (N_7402,N_5619,N_5072);
or U7403 (N_7403,N_6241,N_5697);
or U7404 (N_7404,N_5955,N_5845);
xor U7405 (N_7405,N_5170,N_5883);
or U7406 (N_7406,N_5772,N_5355);
nand U7407 (N_7407,N_5154,N_5417);
nor U7408 (N_7408,N_5294,N_5339);
nand U7409 (N_7409,N_5678,N_6214);
or U7410 (N_7410,N_5693,N_5761);
nor U7411 (N_7411,N_5259,N_5778);
xnor U7412 (N_7412,N_5748,N_5518);
nand U7413 (N_7413,N_5348,N_6023);
xor U7414 (N_7414,N_5749,N_5396);
or U7415 (N_7415,N_5569,N_5764);
xnor U7416 (N_7416,N_6248,N_5632);
and U7417 (N_7417,N_5215,N_5526);
nor U7418 (N_7418,N_5991,N_6001);
nand U7419 (N_7419,N_5712,N_5026);
nand U7420 (N_7420,N_5546,N_5602);
or U7421 (N_7421,N_5277,N_5507);
or U7422 (N_7422,N_6180,N_5749);
nor U7423 (N_7423,N_6031,N_5884);
xor U7424 (N_7424,N_5695,N_5158);
nor U7425 (N_7425,N_5986,N_5910);
xnor U7426 (N_7426,N_5056,N_6242);
xnor U7427 (N_7427,N_5241,N_5135);
xnor U7428 (N_7428,N_5571,N_5262);
nand U7429 (N_7429,N_5682,N_5668);
xor U7430 (N_7430,N_5195,N_5799);
nand U7431 (N_7431,N_6032,N_5349);
nand U7432 (N_7432,N_6161,N_5869);
or U7433 (N_7433,N_5471,N_5446);
nor U7434 (N_7434,N_5079,N_5205);
and U7435 (N_7435,N_5416,N_5393);
nor U7436 (N_7436,N_5302,N_5715);
nor U7437 (N_7437,N_5040,N_5484);
nand U7438 (N_7438,N_5052,N_5187);
xor U7439 (N_7439,N_5698,N_6001);
nor U7440 (N_7440,N_5724,N_6039);
nand U7441 (N_7441,N_5887,N_5355);
and U7442 (N_7442,N_5407,N_5315);
nor U7443 (N_7443,N_5959,N_6089);
xor U7444 (N_7444,N_5812,N_5437);
xnor U7445 (N_7445,N_6155,N_5177);
and U7446 (N_7446,N_5211,N_5681);
and U7447 (N_7447,N_6052,N_5335);
or U7448 (N_7448,N_5936,N_5410);
xnor U7449 (N_7449,N_5747,N_6084);
nand U7450 (N_7450,N_5873,N_5645);
or U7451 (N_7451,N_6241,N_5397);
nor U7452 (N_7452,N_5038,N_5307);
and U7453 (N_7453,N_5351,N_5219);
or U7454 (N_7454,N_5322,N_6152);
nor U7455 (N_7455,N_5527,N_5432);
and U7456 (N_7456,N_5022,N_5379);
and U7457 (N_7457,N_5546,N_5920);
and U7458 (N_7458,N_6112,N_5739);
xor U7459 (N_7459,N_5722,N_5685);
and U7460 (N_7460,N_5699,N_5409);
or U7461 (N_7461,N_6079,N_5647);
or U7462 (N_7462,N_5403,N_5844);
and U7463 (N_7463,N_5411,N_6149);
xor U7464 (N_7464,N_5445,N_5951);
xor U7465 (N_7465,N_6248,N_5856);
nor U7466 (N_7466,N_5538,N_6133);
or U7467 (N_7467,N_5659,N_6186);
xnor U7468 (N_7468,N_5442,N_5286);
or U7469 (N_7469,N_5919,N_5434);
or U7470 (N_7470,N_6113,N_5850);
and U7471 (N_7471,N_5693,N_5885);
xnor U7472 (N_7472,N_5029,N_5532);
nor U7473 (N_7473,N_5208,N_5598);
nor U7474 (N_7474,N_6079,N_5292);
xnor U7475 (N_7475,N_6173,N_5222);
or U7476 (N_7476,N_5319,N_5375);
and U7477 (N_7477,N_6242,N_6075);
nor U7478 (N_7478,N_5326,N_5640);
or U7479 (N_7479,N_6148,N_5887);
xnor U7480 (N_7480,N_5021,N_5254);
and U7481 (N_7481,N_5229,N_5375);
xor U7482 (N_7482,N_5325,N_5699);
nand U7483 (N_7483,N_5262,N_5529);
xor U7484 (N_7484,N_5651,N_6139);
nand U7485 (N_7485,N_6075,N_5103);
and U7486 (N_7486,N_5683,N_5015);
nand U7487 (N_7487,N_6173,N_6243);
and U7488 (N_7488,N_5428,N_6239);
or U7489 (N_7489,N_5422,N_5349);
xor U7490 (N_7490,N_5411,N_5548);
or U7491 (N_7491,N_5172,N_6153);
or U7492 (N_7492,N_5050,N_5328);
xor U7493 (N_7493,N_5334,N_6215);
or U7494 (N_7494,N_5375,N_5100);
or U7495 (N_7495,N_5805,N_5310);
nand U7496 (N_7496,N_6132,N_6101);
or U7497 (N_7497,N_5100,N_5952);
or U7498 (N_7498,N_5316,N_5288);
nand U7499 (N_7499,N_5410,N_6198);
xnor U7500 (N_7500,N_7437,N_6346);
nand U7501 (N_7501,N_7262,N_6690);
nor U7502 (N_7502,N_6648,N_7343);
nor U7503 (N_7503,N_7201,N_7018);
and U7504 (N_7504,N_6385,N_7153);
nor U7505 (N_7505,N_6500,N_7408);
nor U7506 (N_7506,N_6562,N_6675);
nor U7507 (N_7507,N_6963,N_7365);
nor U7508 (N_7508,N_6968,N_6579);
and U7509 (N_7509,N_7099,N_6732);
and U7510 (N_7510,N_6634,N_7357);
or U7511 (N_7511,N_6373,N_7358);
or U7512 (N_7512,N_6640,N_7474);
or U7513 (N_7513,N_6909,N_6689);
nand U7514 (N_7514,N_6979,N_6281);
xnor U7515 (N_7515,N_6682,N_7156);
and U7516 (N_7516,N_7419,N_6730);
or U7517 (N_7517,N_6734,N_6922);
xnor U7518 (N_7518,N_7088,N_7464);
or U7519 (N_7519,N_7140,N_6704);
xor U7520 (N_7520,N_6866,N_7086);
and U7521 (N_7521,N_6895,N_6923);
and U7522 (N_7522,N_7303,N_7272);
nor U7523 (N_7523,N_6265,N_6506);
xnor U7524 (N_7524,N_7440,N_6822);
nand U7525 (N_7525,N_6448,N_7495);
nor U7526 (N_7526,N_7467,N_6466);
xor U7527 (N_7527,N_7050,N_7042);
and U7528 (N_7528,N_7029,N_6902);
nor U7529 (N_7529,N_6967,N_7055);
xor U7530 (N_7530,N_6830,N_6546);
and U7531 (N_7531,N_6667,N_7380);
nor U7532 (N_7532,N_6992,N_6787);
or U7533 (N_7533,N_7300,N_6994);
nor U7534 (N_7534,N_6557,N_6840);
nand U7535 (N_7535,N_6791,N_6697);
and U7536 (N_7536,N_6336,N_7162);
xor U7537 (N_7537,N_7315,N_6314);
nor U7538 (N_7538,N_7187,N_6808);
nor U7539 (N_7539,N_7136,N_6422);
or U7540 (N_7540,N_6811,N_6999);
nor U7541 (N_7541,N_7445,N_6663);
or U7542 (N_7542,N_6862,N_7487);
or U7543 (N_7543,N_7068,N_7493);
or U7544 (N_7544,N_6632,N_7133);
nor U7545 (N_7545,N_7008,N_6622);
xnor U7546 (N_7546,N_7450,N_6429);
nor U7547 (N_7547,N_6550,N_7031);
nor U7548 (N_7548,N_6720,N_6329);
nand U7549 (N_7549,N_6739,N_6788);
nor U7550 (N_7550,N_6919,N_6617);
and U7551 (N_7551,N_6725,N_6918);
and U7552 (N_7552,N_7383,N_6516);
nor U7553 (N_7553,N_7084,N_6576);
nor U7554 (N_7554,N_6600,N_6790);
nand U7555 (N_7555,N_6616,N_7023);
and U7556 (N_7556,N_6816,N_7320);
nor U7557 (N_7557,N_6916,N_6813);
or U7558 (N_7558,N_6761,N_7482);
nor U7559 (N_7559,N_6392,N_6309);
or U7560 (N_7560,N_7334,N_7232);
nand U7561 (N_7561,N_6888,N_6948);
nor U7562 (N_7562,N_6683,N_7172);
nand U7563 (N_7563,N_6712,N_7298);
nor U7564 (N_7564,N_6936,N_6410);
or U7565 (N_7565,N_6296,N_6766);
xor U7566 (N_7566,N_7499,N_7390);
and U7567 (N_7567,N_6363,N_6850);
nand U7568 (N_7568,N_7335,N_7150);
or U7569 (N_7569,N_6450,N_6267);
xnor U7570 (N_7570,N_6631,N_6501);
xnor U7571 (N_7571,N_6860,N_7190);
nand U7572 (N_7572,N_7052,N_6517);
or U7573 (N_7573,N_6731,N_7095);
xnor U7574 (N_7574,N_6626,N_7484);
nand U7575 (N_7575,N_7064,N_7371);
nor U7576 (N_7576,N_7317,N_6252);
or U7577 (N_7577,N_6623,N_7466);
xnor U7578 (N_7578,N_7227,N_6344);
xnor U7579 (N_7579,N_6807,N_7273);
nand U7580 (N_7580,N_7230,N_6904);
xnor U7581 (N_7581,N_6861,N_7436);
or U7582 (N_7582,N_7032,N_6374);
or U7583 (N_7583,N_6913,N_6603);
xor U7584 (N_7584,N_7087,N_6512);
or U7585 (N_7585,N_7220,N_6912);
nor U7586 (N_7586,N_7145,N_7152);
and U7587 (N_7587,N_6726,N_6433);
nand U7588 (N_7588,N_7169,N_7475);
nor U7589 (N_7589,N_7012,N_7441);
or U7590 (N_7590,N_6742,N_6610);
nand U7591 (N_7591,N_6974,N_7070);
or U7592 (N_7592,N_6377,N_6331);
nor U7593 (N_7593,N_6340,N_7433);
nor U7594 (N_7594,N_7128,N_6881);
nand U7595 (N_7595,N_6621,N_6780);
nor U7596 (N_7596,N_7411,N_6359);
nor U7597 (N_7597,N_7455,N_7129);
nor U7598 (N_7598,N_7400,N_6493);
nor U7599 (N_7599,N_7148,N_7447);
xnor U7600 (N_7600,N_7006,N_6376);
xor U7601 (N_7601,N_7237,N_6727);
nor U7602 (N_7602,N_6815,N_7338);
xor U7603 (N_7603,N_7285,N_7213);
or U7604 (N_7604,N_7120,N_6470);
and U7605 (N_7605,N_6473,N_7065);
and U7606 (N_7606,N_6606,N_6629);
nor U7607 (N_7607,N_7289,N_6875);
xnor U7608 (N_7608,N_7356,N_7339);
nand U7609 (N_7609,N_6812,N_7203);
or U7610 (N_7610,N_7184,N_6491);
nand U7611 (N_7611,N_7132,N_6471);
nor U7612 (N_7612,N_6381,N_6857);
xor U7613 (N_7613,N_6954,N_6927);
xnor U7614 (N_7614,N_7082,N_6308);
xnor U7615 (N_7615,N_6962,N_7001);
or U7616 (N_7616,N_6488,N_7336);
and U7617 (N_7617,N_6400,N_6699);
nor U7618 (N_7618,N_7275,N_7229);
or U7619 (N_7619,N_6800,N_6887);
nand U7620 (N_7620,N_6989,N_6438);
nor U7621 (N_7621,N_7100,N_6736);
nor U7622 (N_7622,N_6669,N_7392);
nand U7623 (N_7623,N_6882,N_6275);
and U7624 (N_7624,N_6903,N_6744);
or U7625 (N_7625,N_7139,N_6520);
xnor U7626 (N_7626,N_7243,N_6393);
nor U7627 (N_7627,N_7496,N_7278);
nor U7628 (N_7628,N_7048,N_6554);
nor U7629 (N_7629,N_7208,N_6404);
xnor U7630 (N_7630,N_6784,N_6848);
xnor U7631 (N_7631,N_6778,N_7395);
nor U7632 (N_7632,N_7186,N_7340);
and U7633 (N_7633,N_7118,N_7264);
and U7634 (N_7634,N_6425,N_6785);
xnor U7635 (N_7635,N_7414,N_6986);
xor U7636 (N_7636,N_6728,N_7083);
or U7637 (N_7637,N_6867,N_6818);
nand U7638 (N_7638,N_6543,N_6596);
nand U7639 (N_7639,N_6297,N_7337);
nor U7640 (N_7640,N_6692,N_6598);
and U7641 (N_7641,N_6581,N_6684);
xor U7642 (N_7642,N_7281,N_6773);
nor U7643 (N_7643,N_6713,N_6553);
or U7644 (N_7644,N_6662,N_7266);
xor U7645 (N_7645,N_6435,N_6388);
or U7646 (N_7646,N_7157,N_6328);
nor U7647 (N_7647,N_6349,N_7171);
or U7648 (N_7648,N_6487,N_7454);
or U7649 (N_7649,N_6321,N_6561);
xnor U7650 (N_7650,N_6523,N_6917);
nand U7651 (N_7651,N_6743,N_7387);
xnor U7652 (N_7652,N_6291,N_6284);
xnor U7653 (N_7653,N_7307,N_7355);
nand U7654 (N_7654,N_7277,N_6462);
or U7655 (N_7655,N_6821,N_6570);
and U7656 (N_7656,N_6796,N_6304);
xor U7657 (N_7657,N_6746,N_7325);
and U7658 (N_7658,N_6318,N_7425);
nand U7659 (N_7659,N_6972,N_6958);
xnor U7660 (N_7660,N_7161,N_7451);
nor U7661 (N_7661,N_6883,N_6300);
nor U7662 (N_7662,N_7022,N_7238);
nand U7663 (N_7663,N_7040,N_6261);
nand U7664 (N_7664,N_6464,N_6337);
xnor U7665 (N_7665,N_6863,N_6611);
nand U7666 (N_7666,N_6484,N_6572);
or U7667 (N_7667,N_7292,N_6467);
and U7668 (N_7668,N_6853,N_7252);
or U7669 (N_7669,N_6371,N_7061);
and U7670 (N_7670,N_6293,N_7056);
or U7671 (N_7671,N_7279,N_7051);
nor U7672 (N_7672,N_7016,N_6456);
nor U7673 (N_7673,N_7134,N_7489);
xor U7674 (N_7674,N_7111,N_7457);
or U7675 (N_7675,N_7348,N_6843);
nand U7676 (N_7676,N_6995,N_7033);
xor U7677 (N_7677,N_6402,N_6431);
nand U7678 (N_7678,N_7304,N_6353);
xnor U7679 (N_7679,N_7116,N_7372);
xor U7680 (N_7680,N_6996,N_6799);
or U7681 (N_7681,N_6672,N_7462);
or U7682 (N_7682,N_7296,N_6702);
or U7683 (N_7683,N_6886,N_6421);
xor U7684 (N_7684,N_7193,N_7361);
or U7685 (N_7685,N_6330,N_6717);
nand U7686 (N_7686,N_6375,N_7045);
nand U7687 (N_7687,N_7453,N_7322);
and U7688 (N_7688,N_6571,N_7043);
nor U7689 (N_7689,N_6608,N_6750);
nor U7690 (N_7690,N_6568,N_6294);
and U7691 (N_7691,N_6414,N_7423);
nor U7692 (N_7692,N_6637,N_6872);
nand U7693 (N_7693,N_7416,N_6652);
nand U7694 (N_7694,N_6348,N_7456);
and U7695 (N_7695,N_6490,N_7074);
and U7696 (N_7696,N_6476,N_6382);
or U7697 (N_7697,N_6580,N_6542);
nor U7698 (N_7698,N_6386,N_6698);
nand U7699 (N_7699,N_6953,N_6826);
xor U7700 (N_7700,N_6599,N_6486);
nand U7701 (N_7701,N_6814,N_7114);
or U7702 (N_7702,N_7398,N_7147);
and U7703 (N_7703,N_6437,N_6443);
or U7704 (N_7704,N_7245,N_6264);
xor U7705 (N_7705,N_7446,N_6459);
nor U7706 (N_7706,N_7288,N_6253);
nor U7707 (N_7707,N_6391,N_7362);
or U7708 (N_7708,N_7364,N_7479);
nand U7709 (N_7709,N_7030,N_7182);
and U7710 (N_7710,N_6420,N_7017);
and U7711 (N_7711,N_7389,N_6356);
and U7712 (N_7712,N_6558,N_7314);
xnor U7713 (N_7713,N_6641,N_6288);
nor U7714 (N_7714,N_6893,N_6380);
xor U7715 (N_7715,N_6878,N_6442);
xor U7716 (N_7716,N_7046,N_7236);
nor U7717 (N_7717,N_7160,N_7477);
nand U7718 (N_7718,N_6372,N_6489);
nor U7719 (N_7719,N_6449,N_7297);
or U7720 (N_7720,N_7490,N_6499);
nor U7721 (N_7721,N_6776,N_6984);
and U7722 (N_7722,N_6505,N_6715);
nand U7723 (N_7723,N_7183,N_7353);
and U7724 (N_7724,N_6492,N_7415);
or U7725 (N_7725,N_6323,N_7219);
or U7726 (N_7726,N_6764,N_6707);
xor U7727 (N_7727,N_7097,N_6914);
or U7728 (N_7728,N_6825,N_6360);
nand U7729 (N_7729,N_6636,N_6564);
xor U7730 (N_7730,N_7407,N_7092);
xnor U7731 (N_7731,N_6469,N_6670);
or U7732 (N_7732,N_6898,N_7439);
nand U7733 (N_7733,N_6426,N_6760);
nor U7734 (N_7734,N_6587,N_6901);
or U7735 (N_7735,N_7347,N_7472);
and U7736 (N_7736,N_6347,N_7077);
and U7737 (N_7737,N_7170,N_6534);
and U7738 (N_7738,N_6703,N_6668);
xnor U7739 (N_7739,N_7234,N_6817);
nand U7740 (N_7740,N_7378,N_7002);
nand U7741 (N_7741,N_6943,N_7422);
and U7742 (N_7742,N_6920,N_7216);
nor U7743 (N_7743,N_6590,N_6678);
xor U7744 (N_7744,N_6977,N_6838);
nand U7745 (N_7745,N_7223,N_7350);
nand U7746 (N_7746,N_6705,N_6477);
nand U7747 (N_7747,N_6524,N_7271);
xnor U7748 (N_7748,N_6889,N_7267);
nand U7749 (N_7749,N_7221,N_6320);
nand U7750 (N_7750,N_7149,N_6475);
or U7751 (N_7751,N_7189,N_7141);
or U7752 (N_7752,N_7379,N_6277);
nor U7753 (N_7753,N_7021,N_7151);
nand U7754 (N_7754,N_6547,N_6642);
nand U7755 (N_7755,N_7282,N_7228);
xnor U7756 (N_7756,N_7205,N_6738);
nand U7757 (N_7757,N_6551,N_6514);
nor U7758 (N_7758,N_6322,N_7177);
nor U7759 (N_7759,N_6649,N_6508);
or U7760 (N_7760,N_6250,N_6269);
or U7761 (N_7761,N_6335,N_6978);
or U7762 (N_7762,N_6498,N_6366);
nand U7763 (N_7763,N_6944,N_7401);
xnor U7764 (N_7764,N_6628,N_6755);
or U7765 (N_7765,N_7473,N_7146);
and U7766 (N_7766,N_6256,N_6327);
or U7767 (N_7767,N_7368,N_7094);
xnor U7768 (N_7768,N_7102,N_6398);
nand U7769 (N_7769,N_6938,N_6947);
and U7770 (N_7770,N_6509,N_7027);
nor U7771 (N_7771,N_6656,N_7175);
and U7772 (N_7772,N_6711,N_7098);
nor U7773 (N_7773,N_7109,N_6960);
xnor U7774 (N_7774,N_6751,N_7209);
nor U7775 (N_7775,N_6820,N_7215);
xnor U7776 (N_7776,N_6258,N_6756);
and U7777 (N_7777,N_6532,N_6529);
nor U7778 (N_7778,N_6729,N_6485);
xor U7779 (N_7779,N_6342,N_7091);
or U7780 (N_7780,N_6941,N_7053);
xor U7781 (N_7781,N_7268,N_7104);
or U7782 (N_7782,N_7342,N_6759);
and U7783 (N_7783,N_7404,N_7393);
nand U7784 (N_7784,N_6719,N_6949);
xor U7785 (N_7785,N_6718,N_6535);
or U7786 (N_7786,N_7117,N_6873);
or U7787 (N_7787,N_7105,N_6769);
or U7788 (N_7788,N_6436,N_7251);
and U7789 (N_7789,N_7212,N_6594);
nor U7790 (N_7790,N_7410,N_7443);
xor U7791 (N_7791,N_6876,N_7274);
and U7792 (N_7792,N_7063,N_6653);
and U7793 (N_7793,N_6326,N_6741);
nor U7794 (N_7794,N_6367,N_6829);
and U7795 (N_7795,N_7305,N_7263);
nor U7796 (N_7796,N_6666,N_7284);
xor U7797 (N_7797,N_7034,N_6583);
nor U7798 (N_7798,N_6604,N_6885);
nand U7799 (N_7799,N_6884,N_7013);
or U7800 (N_7800,N_6567,N_7427);
and U7801 (N_7801,N_6869,N_7176);
nor U7802 (N_7802,N_6383,N_6696);
xnor U7803 (N_7803,N_7463,N_6644);
nor U7804 (N_7804,N_7483,N_6762);
xor U7805 (N_7805,N_7085,N_6521);
xnor U7806 (N_7806,N_6455,N_7486);
nand U7807 (N_7807,N_6671,N_6849);
or U7808 (N_7808,N_7321,N_6721);
or U7809 (N_7809,N_6803,N_7078);
nor U7810 (N_7810,N_6896,N_6651);
and U7811 (N_7811,N_6271,N_7039);
nand U7812 (N_7812,N_6654,N_6428);
nor U7813 (N_7813,N_6618,N_7370);
xor U7814 (N_7814,N_7270,N_7381);
nor U7815 (N_7815,N_6708,N_7351);
nor U7816 (N_7816,N_6679,N_7211);
and U7817 (N_7817,N_6877,N_7256);
or U7818 (N_7818,N_6665,N_7138);
and U7819 (N_7819,N_7424,N_6993);
or U7820 (N_7820,N_6681,N_6797);
and U7821 (N_7821,N_7096,N_6771);
nor U7822 (N_7822,N_6842,N_6806);
or U7823 (N_7823,N_6724,N_7384);
and U7824 (N_7824,N_7326,N_7071);
nor U7825 (N_7825,N_6779,N_7011);
nor U7826 (N_7826,N_6528,N_6864);
and U7827 (N_7827,N_6758,N_6802);
nor U7828 (N_7828,N_6370,N_7310);
or U7829 (N_7829,N_6686,N_6894);
xor U7830 (N_7830,N_6997,N_6573);
nand U7831 (N_7831,N_6339,N_7498);
nor U7832 (N_7832,N_6833,N_6418);
and U7833 (N_7833,N_6351,N_7058);
and U7834 (N_7834,N_6384,N_6539);
and U7835 (N_7835,N_7204,N_7076);
nor U7836 (N_7836,N_6504,N_7276);
xnor U7837 (N_7837,N_7429,N_6819);
xnor U7838 (N_7838,N_6358,N_6441);
or U7839 (N_7839,N_7185,N_6472);
nand U7840 (N_7840,N_7470,N_7460);
nand U7841 (N_7841,N_7382,N_7163);
nor U7842 (N_7842,N_6595,N_6447);
nand U7843 (N_7843,N_6956,N_6440);
or U7844 (N_7844,N_6775,N_7485);
xor U7845 (N_7845,N_6757,N_6891);
nand U7846 (N_7846,N_6983,N_7349);
or U7847 (N_7847,N_6502,N_6763);
and U7848 (N_7848,N_6460,N_6292);
nand U7849 (N_7849,N_7135,N_7412);
or U7850 (N_7850,N_6854,N_6846);
nor U7851 (N_7851,N_6740,N_6439);
xnor U7852 (N_7852,N_7452,N_7009);
xor U7853 (N_7853,N_6343,N_6369);
xnor U7854 (N_7854,N_7036,N_7481);
nor U7855 (N_7855,N_7214,N_6709);
nand U7856 (N_7856,N_6851,N_7000);
and U7857 (N_7857,N_6844,N_6874);
and U7858 (N_7858,N_7198,N_6676);
and U7859 (N_7859,N_6387,N_6933);
or U7860 (N_7860,N_6701,N_6605);
or U7861 (N_7861,N_6494,N_6577);
or U7862 (N_7862,N_6480,N_6985);
or U7863 (N_7863,N_6510,N_7143);
nor U7864 (N_7864,N_6980,N_7283);
xnor U7865 (N_7865,N_7258,N_7253);
nand U7866 (N_7866,N_6687,N_6607);
nor U7867 (N_7867,N_6798,N_6453);
or U7868 (N_7868,N_6908,N_6965);
and U7869 (N_7869,N_7331,N_6262);
or U7870 (N_7870,N_7461,N_6301);
nand U7871 (N_7871,N_6319,N_6620);
or U7872 (N_7872,N_7260,N_6955);
or U7873 (N_7873,N_6781,N_6531);
nand U7874 (N_7874,N_6445,N_6871);
nand U7875 (N_7875,N_6483,N_6299);
or U7876 (N_7876,N_6688,N_7197);
or U7877 (N_7877,N_6973,N_7089);
or U7878 (N_7878,N_6768,N_6563);
or U7879 (N_7879,N_7020,N_6278);
and U7880 (N_7880,N_6839,N_7069);
nand U7881 (N_7881,N_7025,N_6417);
and U7882 (N_7882,N_6513,N_6633);
xor U7883 (N_7883,N_6770,N_7309);
nor U7884 (N_7884,N_6906,N_6952);
nand U7885 (N_7885,N_7377,N_7291);
xnor U7886 (N_7886,N_6619,N_6868);
nor U7887 (N_7887,N_6859,N_6597);
or U7888 (N_7888,N_6530,N_6910);
and U7889 (N_7889,N_7311,N_7014);
and U7890 (N_7890,N_6706,N_7328);
or U7891 (N_7891,N_7257,N_7442);
xor U7892 (N_7892,N_6612,N_6899);
nor U7893 (N_7893,N_7323,N_7494);
or U7894 (N_7894,N_6852,N_6461);
nor U7895 (N_7895,N_7003,N_6627);
nand U7896 (N_7896,N_7476,N_6823);
or U7897 (N_7897,N_7103,N_6541);
and U7898 (N_7898,N_7374,N_6911);
and U7899 (N_7899,N_6354,N_6394);
and U7900 (N_7900,N_6749,N_7155);
or U7901 (N_7901,N_6260,N_6970);
nand U7902 (N_7902,N_6397,N_6457);
nor U7903 (N_7903,N_6987,N_6880);
nand U7904 (N_7904,N_7459,N_6497);
xnor U7905 (N_7905,N_6990,N_7194);
nor U7906 (N_7906,N_6324,N_6411);
or U7907 (N_7907,N_6463,N_6975);
and U7908 (N_7908,N_6522,N_6474);
and U7909 (N_7909,N_6635,N_7038);
xor U7910 (N_7910,N_6793,N_6341);
nor U7911 (N_7911,N_7072,N_6403);
nand U7912 (N_7912,N_7265,N_6276);
and U7913 (N_7913,N_6575,N_6511);
and U7914 (N_7914,N_6971,N_6409);
and U7915 (N_7915,N_6519,N_7075);
xor U7916 (N_7916,N_6602,N_7280);
or U7917 (N_7917,N_7435,N_6824);
or U7918 (N_7918,N_6496,N_6794);
nand U7919 (N_7919,N_6451,N_7241);
xor U7920 (N_7920,N_7402,N_7385);
or U7921 (N_7921,N_7417,N_6415);
xor U7922 (N_7922,N_7324,N_6615);
or U7923 (N_7923,N_7049,N_7035);
and U7924 (N_7924,N_6925,N_6930);
and U7925 (N_7925,N_7196,N_7480);
or U7926 (N_7926,N_6714,N_7130);
xor U7927 (N_7927,N_6931,N_6548);
xnor U7928 (N_7928,N_7388,N_7218);
xor U7929 (N_7929,N_7418,N_6939);
xor U7930 (N_7930,N_7491,N_6801);
or U7931 (N_7931,N_7469,N_7206);
xnor U7932 (N_7932,N_6565,N_7360);
xor U7933 (N_7933,N_7240,N_6638);
and U7934 (N_7934,N_7316,N_6693);
xor U7935 (N_7935,N_6834,N_6915);
xnor U7936 (N_7936,N_7301,N_6691);
nor U7937 (N_7937,N_7354,N_6396);
or U7938 (N_7938,N_6795,N_6325);
and U7939 (N_7939,N_7269,N_7019);
or U7940 (N_7940,N_7405,N_7225);
or U7941 (N_7941,N_7413,N_6536);
and U7942 (N_7942,N_6694,N_6259);
or U7943 (N_7943,N_6828,N_7158);
and U7944 (N_7944,N_6549,N_7290);
or U7945 (N_7945,N_6723,N_7122);
nand U7946 (N_7946,N_6545,N_6745);
nand U7947 (N_7947,N_7492,N_7397);
or U7948 (N_7948,N_6355,N_7449);
and U7949 (N_7949,N_7333,N_6482);
nor U7950 (N_7950,N_6786,N_6934);
or U7951 (N_7951,N_6584,N_6290);
or U7952 (N_7952,N_7233,N_7073);
xnor U7953 (N_7953,N_7359,N_7115);
xor U7954 (N_7954,N_6655,N_6478);
nor U7955 (N_7955,N_6928,N_6589);
xor U7956 (N_7956,N_7468,N_6270);
or U7957 (N_7957,N_6361,N_7312);
and U7958 (N_7958,N_6312,N_7329);
nand U7959 (N_7959,N_6810,N_6660);
nor U7960 (N_7960,N_7458,N_6465);
xnor U7961 (N_7961,N_7173,N_6625);
xnor U7962 (N_7962,N_6303,N_6332);
nor U7963 (N_7963,N_6932,N_7376);
and U7964 (N_7964,N_6272,N_6389);
xnor U7965 (N_7965,N_6350,N_6700);
or U7966 (N_7966,N_6964,N_7131);
nand U7967 (N_7967,N_7344,N_6735);
or U7968 (N_7968,N_6427,N_7255);
and U7969 (N_7969,N_7144,N_6837);
or U7970 (N_7970,N_6544,N_6609);
xnor U7971 (N_7971,N_6338,N_6378);
xor U7972 (N_7972,N_6503,N_6991);
or U7973 (N_7973,N_6365,N_6747);
or U7974 (N_7974,N_7179,N_7247);
nand U7975 (N_7975,N_7409,N_6317);
and U7976 (N_7976,N_6827,N_6674);
nand U7977 (N_7977,N_6279,N_7330);
and U7978 (N_7978,N_7250,N_6832);
nand U7979 (N_7979,N_7199,N_7166);
nor U7980 (N_7980,N_6792,N_6783);
and U7981 (N_7981,N_7394,N_7007);
and U7982 (N_7982,N_6658,N_6283);
xnor U7983 (N_7983,N_6646,N_6804);
nand U7984 (N_7984,N_7192,N_6555);
nor U7985 (N_7985,N_7059,N_6772);
nor U7986 (N_7986,N_6664,N_6677);
or U7987 (N_7987,N_7369,N_7067);
or U7988 (N_7988,N_7341,N_6405);
xor U7989 (N_7989,N_7261,N_6316);
and U7990 (N_7990,N_6255,N_7471);
xor U7991 (N_7991,N_6789,N_7167);
or U7992 (N_7992,N_7231,N_6897);
xnor U7993 (N_7993,N_6643,N_7430);
xnor U7994 (N_7994,N_6419,N_6569);
or U7995 (N_7995,N_6454,N_7079);
and U7996 (N_7996,N_6458,N_6395);
nor U7997 (N_7997,N_6406,N_6659);
nand U7998 (N_7998,N_7178,N_6657);
nand U7999 (N_7999,N_7222,N_6518);
xnor U8000 (N_8000,N_6614,N_7363);
xor U8001 (N_8001,N_7478,N_7137);
nor U8002 (N_8002,N_6313,N_6527);
nor U8003 (N_8003,N_6782,N_6722);
xnor U8004 (N_8004,N_7244,N_7047);
nor U8005 (N_8005,N_6945,N_6890);
xor U8006 (N_8006,N_6847,N_7044);
and U8007 (N_8007,N_6737,N_6716);
xor U8008 (N_8008,N_7028,N_6507);
nor U8009 (N_8009,N_7174,N_7421);
and U8010 (N_8010,N_7420,N_7432);
and U8011 (N_8011,N_6673,N_6900);
nand U8012 (N_8012,N_7286,N_6263);
nand U8013 (N_8013,N_7165,N_7375);
nand U8014 (N_8014,N_6592,N_7180);
and U8015 (N_8015,N_6452,N_6929);
nand U8016 (N_8016,N_7386,N_6298);
nor U8017 (N_8017,N_6752,N_6413);
nand U8018 (N_8018,N_6951,N_6586);
nor U8019 (N_8019,N_7154,N_6407);
nor U8020 (N_8020,N_7367,N_6845);
and U8021 (N_8021,N_6765,N_6302);
xnor U8022 (N_8022,N_6266,N_7207);
nor U8023 (N_8023,N_7426,N_7308);
and U8024 (N_8024,N_7254,N_6585);
nor U8025 (N_8025,N_7090,N_6286);
and U8026 (N_8026,N_7024,N_6865);
xor U8027 (N_8027,N_6998,N_6858);
xor U8028 (N_8028,N_7060,N_6560);
nand U8029 (N_8029,N_6423,N_7306);
and U8030 (N_8030,N_6856,N_6754);
nor U8031 (N_8031,N_7431,N_6926);
xor U8032 (N_8032,N_6578,N_6748);
nand U8033 (N_8033,N_6710,N_7346);
nand U8034 (N_8034,N_6273,N_6556);
and U8035 (N_8035,N_7066,N_6401);
xnor U8036 (N_8036,N_7005,N_6552);
nor U8037 (N_8037,N_7246,N_6613);
or U8038 (N_8038,N_7295,N_7434);
and U8039 (N_8039,N_7101,N_7015);
xnor U8040 (N_8040,N_6988,N_6468);
xor U8041 (N_8041,N_6364,N_6946);
xnor U8042 (N_8042,N_6333,N_6767);
and U8043 (N_8043,N_7054,N_6533);
or U8044 (N_8044,N_7248,N_6582);
or U8045 (N_8045,N_6289,N_6379);
nand U8046 (N_8046,N_6695,N_6434);
xnor U8047 (N_8047,N_6424,N_6495);
nor U8048 (N_8048,N_6280,N_6924);
or U8049 (N_8049,N_7123,N_6591);
nand U8050 (N_8050,N_7302,N_7057);
and U8051 (N_8051,N_7026,N_6310);
xor U8052 (N_8052,N_7366,N_7159);
nand U8053 (N_8053,N_7287,N_7188);
nand U8054 (N_8054,N_6408,N_6835);
or U8055 (N_8055,N_7345,N_6907);
nand U8056 (N_8056,N_6287,N_7226);
or U8057 (N_8057,N_7010,N_6921);
and U8058 (N_8058,N_7106,N_6334);
nor U8059 (N_8059,N_6831,N_7428);
or U8060 (N_8060,N_7107,N_6976);
or U8061 (N_8061,N_6285,N_6661);
nor U8062 (N_8062,N_6753,N_7444);
xnor U8063 (N_8063,N_6959,N_6809);
nor U8064 (N_8064,N_6566,N_6905);
or U8065 (N_8065,N_6981,N_6805);
nand U8066 (N_8066,N_7465,N_6390);
or U8067 (N_8067,N_7202,N_6982);
and U8068 (N_8068,N_7497,N_7119);
xor U8069 (N_8069,N_6345,N_6935);
and U8070 (N_8070,N_6593,N_7293);
nor U8071 (N_8071,N_7112,N_6412);
nand U8072 (N_8072,N_7113,N_6892);
nand U8073 (N_8073,N_7438,N_6515);
or U8074 (N_8074,N_7191,N_6639);
nand U8075 (N_8075,N_6311,N_7373);
or U8076 (N_8076,N_7242,N_7352);
nor U8077 (N_8077,N_6685,N_6841);
and U8078 (N_8078,N_7217,N_7108);
nand U8079 (N_8079,N_6481,N_7294);
or U8080 (N_8080,N_6574,N_7403);
and U8081 (N_8081,N_7391,N_6368);
and U8082 (N_8082,N_6430,N_7126);
xnor U8083 (N_8083,N_6352,N_6733);
nand U8084 (N_8084,N_6950,N_7181);
and U8085 (N_8085,N_6588,N_6957);
xor U8086 (N_8086,N_6416,N_6540);
nor U8087 (N_8087,N_7259,N_7406);
nand U8088 (N_8088,N_6879,N_6966);
or U8089 (N_8089,N_6940,N_7299);
or U8090 (N_8090,N_6836,N_7080);
or U8091 (N_8091,N_6274,N_6526);
nand U8092 (N_8092,N_7318,N_7235);
and U8093 (N_8093,N_6969,N_6624);
xor U8094 (N_8094,N_6444,N_7093);
or U8095 (N_8095,N_7124,N_7164);
xor U8096 (N_8096,N_6295,N_6305);
and U8097 (N_8097,N_7081,N_6282);
nand U8098 (N_8098,N_6254,N_7121);
xor U8099 (N_8099,N_7332,N_6601);
nor U8100 (N_8100,N_6870,N_6647);
and U8101 (N_8101,N_7037,N_6525);
and U8102 (N_8102,N_6251,N_6432);
nand U8103 (N_8103,N_7319,N_7399);
nand U8104 (N_8104,N_6630,N_7488);
and U8105 (N_8105,N_6257,N_6306);
nor U8106 (N_8106,N_6559,N_6362);
xnor U8107 (N_8107,N_6315,N_6357);
or U8108 (N_8108,N_6937,N_7004);
and U8109 (N_8109,N_7249,N_6268);
nor U8110 (N_8110,N_7110,N_7224);
and U8111 (N_8111,N_7127,N_7168);
xor U8112 (N_8112,N_6399,N_6777);
nand U8113 (N_8113,N_6479,N_7041);
xnor U8114 (N_8114,N_6855,N_6537);
or U8115 (N_8115,N_6774,N_7125);
and U8116 (N_8116,N_7062,N_6307);
or U8117 (N_8117,N_7448,N_6538);
nand U8118 (N_8118,N_7200,N_7313);
or U8119 (N_8119,N_6650,N_7210);
nor U8120 (N_8120,N_7327,N_7142);
xnor U8121 (N_8121,N_6680,N_7195);
and U8122 (N_8122,N_6942,N_6645);
or U8123 (N_8123,N_7239,N_7396);
or U8124 (N_8124,N_6446,N_6961);
xnor U8125 (N_8125,N_7063,N_6908);
or U8126 (N_8126,N_6258,N_7384);
nand U8127 (N_8127,N_7042,N_6717);
or U8128 (N_8128,N_7220,N_7014);
nor U8129 (N_8129,N_7186,N_6441);
nor U8130 (N_8130,N_7093,N_7325);
or U8131 (N_8131,N_6258,N_6922);
or U8132 (N_8132,N_6802,N_7241);
and U8133 (N_8133,N_6896,N_7405);
xor U8134 (N_8134,N_6563,N_7294);
nand U8135 (N_8135,N_6349,N_7065);
or U8136 (N_8136,N_6635,N_6416);
xor U8137 (N_8137,N_7485,N_6252);
and U8138 (N_8138,N_7129,N_6299);
or U8139 (N_8139,N_6417,N_6372);
and U8140 (N_8140,N_6472,N_6328);
xor U8141 (N_8141,N_6811,N_7237);
xnor U8142 (N_8142,N_6301,N_6974);
xor U8143 (N_8143,N_6999,N_6398);
and U8144 (N_8144,N_7055,N_6633);
and U8145 (N_8145,N_6364,N_7050);
or U8146 (N_8146,N_6507,N_7426);
or U8147 (N_8147,N_6964,N_6577);
or U8148 (N_8148,N_6896,N_7304);
and U8149 (N_8149,N_7125,N_6456);
xnor U8150 (N_8150,N_6299,N_6316);
xnor U8151 (N_8151,N_6262,N_7241);
and U8152 (N_8152,N_7472,N_6793);
or U8153 (N_8153,N_6403,N_7227);
xnor U8154 (N_8154,N_7335,N_7140);
and U8155 (N_8155,N_7474,N_7473);
nor U8156 (N_8156,N_6312,N_6901);
or U8157 (N_8157,N_7360,N_6441);
and U8158 (N_8158,N_6935,N_6803);
and U8159 (N_8159,N_7075,N_6933);
nor U8160 (N_8160,N_6883,N_7439);
or U8161 (N_8161,N_6642,N_6776);
xor U8162 (N_8162,N_7243,N_7236);
or U8163 (N_8163,N_6957,N_6978);
nor U8164 (N_8164,N_7253,N_6766);
nand U8165 (N_8165,N_7400,N_6760);
or U8166 (N_8166,N_7319,N_6621);
or U8167 (N_8167,N_7089,N_7308);
xnor U8168 (N_8168,N_6594,N_7473);
xnor U8169 (N_8169,N_6328,N_7199);
xor U8170 (N_8170,N_6255,N_7376);
nor U8171 (N_8171,N_6325,N_6683);
xor U8172 (N_8172,N_7396,N_7291);
xor U8173 (N_8173,N_6288,N_7275);
nand U8174 (N_8174,N_6861,N_7347);
or U8175 (N_8175,N_6414,N_6575);
nand U8176 (N_8176,N_7274,N_7133);
and U8177 (N_8177,N_6440,N_7335);
nand U8178 (N_8178,N_7311,N_6423);
nor U8179 (N_8179,N_6967,N_6432);
or U8180 (N_8180,N_6415,N_7076);
or U8181 (N_8181,N_6691,N_6581);
nand U8182 (N_8182,N_6607,N_7027);
or U8183 (N_8183,N_6849,N_7264);
nor U8184 (N_8184,N_7488,N_7486);
and U8185 (N_8185,N_7302,N_6876);
nor U8186 (N_8186,N_6432,N_7371);
or U8187 (N_8187,N_7267,N_6776);
nand U8188 (N_8188,N_6456,N_6417);
or U8189 (N_8189,N_6856,N_6866);
nor U8190 (N_8190,N_6488,N_7224);
nor U8191 (N_8191,N_7133,N_6992);
nand U8192 (N_8192,N_6941,N_7132);
xnor U8193 (N_8193,N_6648,N_6451);
nand U8194 (N_8194,N_6613,N_6828);
nand U8195 (N_8195,N_7274,N_7025);
or U8196 (N_8196,N_6790,N_6586);
xor U8197 (N_8197,N_7076,N_6705);
nand U8198 (N_8198,N_6434,N_7331);
nor U8199 (N_8199,N_6844,N_7294);
xor U8200 (N_8200,N_6681,N_6878);
or U8201 (N_8201,N_6864,N_6800);
and U8202 (N_8202,N_6901,N_6693);
xnor U8203 (N_8203,N_7173,N_7086);
nor U8204 (N_8204,N_7279,N_6688);
nor U8205 (N_8205,N_7248,N_6897);
xnor U8206 (N_8206,N_6492,N_6868);
nand U8207 (N_8207,N_7165,N_7303);
and U8208 (N_8208,N_7347,N_6278);
and U8209 (N_8209,N_7083,N_6847);
and U8210 (N_8210,N_6483,N_6446);
nand U8211 (N_8211,N_6627,N_7410);
and U8212 (N_8212,N_7065,N_6951);
and U8213 (N_8213,N_6327,N_6903);
and U8214 (N_8214,N_6574,N_7017);
and U8215 (N_8215,N_6342,N_6980);
nand U8216 (N_8216,N_7224,N_6454);
or U8217 (N_8217,N_6312,N_6479);
and U8218 (N_8218,N_6698,N_6520);
nor U8219 (N_8219,N_6986,N_7209);
nand U8220 (N_8220,N_7151,N_6679);
xor U8221 (N_8221,N_6624,N_7460);
nor U8222 (N_8222,N_7089,N_6958);
and U8223 (N_8223,N_7039,N_7298);
or U8224 (N_8224,N_7185,N_6695);
nor U8225 (N_8225,N_7490,N_7287);
nand U8226 (N_8226,N_6593,N_6417);
and U8227 (N_8227,N_7294,N_6883);
xnor U8228 (N_8228,N_6812,N_6656);
and U8229 (N_8229,N_7097,N_6298);
nand U8230 (N_8230,N_7221,N_6514);
and U8231 (N_8231,N_7369,N_7211);
nand U8232 (N_8232,N_6403,N_6250);
or U8233 (N_8233,N_6337,N_7359);
or U8234 (N_8234,N_7243,N_6371);
or U8235 (N_8235,N_7461,N_6596);
and U8236 (N_8236,N_6895,N_6753);
or U8237 (N_8237,N_6899,N_6548);
xor U8238 (N_8238,N_7251,N_6635);
xor U8239 (N_8239,N_6729,N_6542);
and U8240 (N_8240,N_6839,N_6818);
nand U8241 (N_8241,N_6595,N_6906);
nor U8242 (N_8242,N_6949,N_6737);
nand U8243 (N_8243,N_6678,N_7275);
and U8244 (N_8244,N_7212,N_6372);
and U8245 (N_8245,N_7346,N_6877);
nand U8246 (N_8246,N_6688,N_7275);
and U8247 (N_8247,N_6691,N_7437);
nor U8248 (N_8248,N_6848,N_7028);
nand U8249 (N_8249,N_6392,N_7479);
or U8250 (N_8250,N_7434,N_7059);
nand U8251 (N_8251,N_6839,N_7384);
and U8252 (N_8252,N_7080,N_6487);
nor U8253 (N_8253,N_6672,N_6776);
nand U8254 (N_8254,N_6360,N_6724);
xnor U8255 (N_8255,N_7285,N_7130);
xnor U8256 (N_8256,N_6743,N_7087);
nor U8257 (N_8257,N_6544,N_7174);
and U8258 (N_8258,N_7495,N_6757);
xor U8259 (N_8259,N_6312,N_6444);
xor U8260 (N_8260,N_7408,N_7172);
nor U8261 (N_8261,N_7210,N_7497);
nor U8262 (N_8262,N_7051,N_7207);
nor U8263 (N_8263,N_6919,N_6671);
or U8264 (N_8264,N_6641,N_6784);
xor U8265 (N_8265,N_6381,N_6800);
or U8266 (N_8266,N_6425,N_6677);
and U8267 (N_8267,N_7475,N_7080);
xnor U8268 (N_8268,N_6734,N_7243);
and U8269 (N_8269,N_6470,N_6262);
or U8270 (N_8270,N_7087,N_6863);
xor U8271 (N_8271,N_6346,N_6648);
or U8272 (N_8272,N_6917,N_6769);
nand U8273 (N_8273,N_6610,N_6919);
or U8274 (N_8274,N_6697,N_7287);
xnor U8275 (N_8275,N_6797,N_7073);
and U8276 (N_8276,N_6906,N_6920);
xnor U8277 (N_8277,N_6751,N_6931);
nand U8278 (N_8278,N_6571,N_7388);
nor U8279 (N_8279,N_6456,N_6298);
or U8280 (N_8280,N_6359,N_6595);
xnor U8281 (N_8281,N_6627,N_7355);
nor U8282 (N_8282,N_7367,N_6379);
nand U8283 (N_8283,N_7380,N_7270);
xor U8284 (N_8284,N_6554,N_6766);
nor U8285 (N_8285,N_7390,N_6280);
nor U8286 (N_8286,N_6699,N_7260);
xnor U8287 (N_8287,N_6604,N_7155);
xor U8288 (N_8288,N_7318,N_6970);
or U8289 (N_8289,N_7290,N_7214);
and U8290 (N_8290,N_6618,N_7216);
or U8291 (N_8291,N_6494,N_6394);
nor U8292 (N_8292,N_7064,N_6583);
and U8293 (N_8293,N_6891,N_6534);
xor U8294 (N_8294,N_7426,N_6332);
or U8295 (N_8295,N_7170,N_7367);
or U8296 (N_8296,N_7255,N_7330);
nor U8297 (N_8297,N_6648,N_6818);
nand U8298 (N_8298,N_6840,N_6529);
and U8299 (N_8299,N_7310,N_6561);
or U8300 (N_8300,N_7316,N_6590);
nor U8301 (N_8301,N_7105,N_6806);
and U8302 (N_8302,N_6542,N_7060);
nand U8303 (N_8303,N_6545,N_6308);
nor U8304 (N_8304,N_7039,N_6620);
or U8305 (N_8305,N_6276,N_6463);
or U8306 (N_8306,N_6976,N_6605);
or U8307 (N_8307,N_7222,N_6657);
xnor U8308 (N_8308,N_7362,N_7258);
xnor U8309 (N_8309,N_6861,N_6564);
and U8310 (N_8310,N_6975,N_7103);
xor U8311 (N_8311,N_7058,N_6878);
xnor U8312 (N_8312,N_6418,N_6972);
nor U8313 (N_8313,N_7396,N_7386);
nand U8314 (N_8314,N_7441,N_7364);
and U8315 (N_8315,N_6765,N_6684);
or U8316 (N_8316,N_7115,N_7488);
xnor U8317 (N_8317,N_6829,N_6637);
xor U8318 (N_8318,N_6678,N_7052);
and U8319 (N_8319,N_6951,N_7233);
xor U8320 (N_8320,N_7392,N_7186);
nor U8321 (N_8321,N_7155,N_6364);
xor U8322 (N_8322,N_6367,N_6948);
xnor U8323 (N_8323,N_6870,N_6651);
xnor U8324 (N_8324,N_7057,N_6431);
and U8325 (N_8325,N_7311,N_6614);
and U8326 (N_8326,N_6317,N_6904);
nand U8327 (N_8327,N_7165,N_7023);
nor U8328 (N_8328,N_6730,N_7094);
xnor U8329 (N_8329,N_7192,N_6405);
and U8330 (N_8330,N_7438,N_7279);
nor U8331 (N_8331,N_6362,N_6845);
or U8332 (N_8332,N_7177,N_7431);
and U8333 (N_8333,N_6914,N_6727);
nand U8334 (N_8334,N_6402,N_7070);
xnor U8335 (N_8335,N_6913,N_7047);
xnor U8336 (N_8336,N_6309,N_6896);
and U8337 (N_8337,N_7165,N_6872);
or U8338 (N_8338,N_7036,N_7090);
and U8339 (N_8339,N_7167,N_7230);
or U8340 (N_8340,N_7405,N_6278);
and U8341 (N_8341,N_6725,N_6805);
nand U8342 (N_8342,N_7035,N_7445);
nand U8343 (N_8343,N_6336,N_6807);
and U8344 (N_8344,N_6475,N_7102);
nor U8345 (N_8345,N_6264,N_6833);
and U8346 (N_8346,N_6346,N_7299);
and U8347 (N_8347,N_7019,N_6815);
and U8348 (N_8348,N_7007,N_6610);
or U8349 (N_8349,N_7430,N_7149);
or U8350 (N_8350,N_6379,N_7312);
xor U8351 (N_8351,N_6341,N_6608);
xor U8352 (N_8352,N_7346,N_6261);
or U8353 (N_8353,N_7391,N_6688);
or U8354 (N_8354,N_6825,N_7022);
or U8355 (N_8355,N_6831,N_6611);
and U8356 (N_8356,N_6759,N_7371);
nand U8357 (N_8357,N_6378,N_6963);
nand U8358 (N_8358,N_7073,N_7342);
nand U8359 (N_8359,N_6552,N_6944);
or U8360 (N_8360,N_6781,N_6961);
or U8361 (N_8361,N_6654,N_6777);
and U8362 (N_8362,N_6795,N_6678);
xnor U8363 (N_8363,N_6690,N_6408);
and U8364 (N_8364,N_7004,N_6736);
or U8365 (N_8365,N_6875,N_7120);
xor U8366 (N_8366,N_6389,N_7490);
and U8367 (N_8367,N_7185,N_6846);
or U8368 (N_8368,N_6972,N_6301);
nor U8369 (N_8369,N_7245,N_6408);
and U8370 (N_8370,N_7205,N_6891);
nand U8371 (N_8371,N_6344,N_7236);
xor U8372 (N_8372,N_6473,N_6746);
xnor U8373 (N_8373,N_7174,N_7347);
and U8374 (N_8374,N_6650,N_6821);
and U8375 (N_8375,N_7081,N_6648);
nor U8376 (N_8376,N_7049,N_6271);
nand U8377 (N_8377,N_7273,N_6965);
nor U8378 (N_8378,N_7332,N_7476);
or U8379 (N_8379,N_7241,N_7058);
xor U8380 (N_8380,N_7183,N_7278);
nand U8381 (N_8381,N_6293,N_6526);
xor U8382 (N_8382,N_6655,N_6951);
nor U8383 (N_8383,N_6656,N_7017);
xor U8384 (N_8384,N_6578,N_6688);
nand U8385 (N_8385,N_6652,N_6731);
or U8386 (N_8386,N_6533,N_7061);
nand U8387 (N_8387,N_6955,N_6352);
nor U8388 (N_8388,N_7262,N_6584);
xnor U8389 (N_8389,N_7489,N_7472);
and U8390 (N_8390,N_7393,N_7139);
xor U8391 (N_8391,N_7239,N_7041);
or U8392 (N_8392,N_6616,N_7320);
nand U8393 (N_8393,N_7292,N_6884);
nor U8394 (N_8394,N_6768,N_6805);
and U8395 (N_8395,N_6642,N_6543);
nor U8396 (N_8396,N_7378,N_7149);
and U8397 (N_8397,N_7342,N_7215);
and U8398 (N_8398,N_7490,N_7308);
nor U8399 (N_8399,N_7069,N_7261);
and U8400 (N_8400,N_7016,N_6572);
nor U8401 (N_8401,N_6885,N_6883);
nor U8402 (N_8402,N_6255,N_7491);
and U8403 (N_8403,N_6690,N_7152);
and U8404 (N_8404,N_6937,N_6632);
nor U8405 (N_8405,N_6255,N_6534);
xor U8406 (N_8406,N_6420,N_7027);
and U8407 (N_8407,N_7307,N_6379);
nand U8408 (N_8408,N_6681,N_6695);
and U8409 (N_8409,N_6406,N_7000);
xor U8410 (N_8410,N_6879,N_6498);
nand U8411 (N_8411,N_6507,N_7203);
xnor U8412 (N_8412,N_7370,N_6692);
or U8413 (N_8413,N_7452,N_7409);
xnor U8414 (N_8414,N_6814,N_7193);
xor U8415 (N_8415,N_7355,N_7251);
xnor U8416 (N_8416,N_7326,N_6604);
nor U8417 (N_8417,N_7350,N_6773);
nor U8418 (N_8418,N_7478,N_6342);
nor U8419 (N_8419,N_6896,N_7147);
or U8420 (N_8420,N_6934,N_6914);
nor U8421 (N_8421,N_7435,N_6718);
and U8422 (N_8422,N_7163,N_6540);
xnor U8423 (N_8423,N_6468,N_7236);
and U8424 (N_8424,N_7155,N_6370);
xor U8425 (N_8425,N_7495,N_6496);
and U8426 (N_8426,N_6565,N_6987);
nand U8427 (N_8427,N_7272,N_7294);
nand U8428 (N_8428,N_7083,N_6492);
or U8429 (N_8429,N_6562,N_6372);
xor U8430 (N_8430,N_6254,N_6731);
nand U8431 (N_8431,N_6989,N_6516);
nand U8432 (N_8432,N_6695,N_6288);
nor U8433 (N_8433,N_7049,N_6375);
nor U8434 (N_8434,N_7065,N_6791);
nor U8435 (N_8435,N_6577,N_6442);
or U8436 (N_8436,N_6549,N_7327);
nor U8437 (N_8437,N_6597,N_6592);
or U8438 (N_8438,N_7291,N_7318);
or U8439 (N_8439,N_6872,N_7181);
xor U8440 (N_8440,N_7419,N_7202);
and U8441 (N_8441,N_6994,N_6536);
nor U8442 (N_8442,N_7118,N_7116);
xor U8443 (N_8443,N_6896,N_7379);
nor U8444 (N_8444,N_6421,N_7108);
or U8445 (N_8445,N_6892,N_7331);
xnor U8446 (N_8446,N_7116,N_7017);
nor U8447 (N_8447,N_6647,N_7311);
and U8448 (N_8448,N_6947,N_6688);
and U8449 (N_8449,N_7402,N_7237);
or U8450 (N_8450,N_7371,N_7401);
or U8451 (N_8451,N_6712,N_7083);
xnor U8452 (N_8452,N_7490,N_6255);
nor U8453 (N_8453,N_6466,N_6864);
xor U8454 (N_8454,N_6566,N_6818);
and U8455 (N_8455,N_6580,N_6426);
xor U8456 (N_8456,N_7382,N_7364);
or U8457 (N_8457,N_7305,N_6420);
nor U8458 (N_8458,N_6396,N_6639);
or U8459 (N_8459,N_7038,N_7151);
or U8460 (N_8460,N_6484,N_6791);
nand U8461 (N_8461,N_7074,N_6564);
nor U8462 (N_8462,N_7221,N_6307);
xnor U8463 (N_8463,N_7486,N_7279);
xnor U8464 (N_8464,N_7162,N_6779);
and U8465 (N_8465,N_7348,N_7402);
and U8466 (N_8466,N_6853,N_6660);
and U8467 (N_8467,N_7376,N_7363);
or U8468 (N_8468,N_7486,N_6616);
and U8469 (N_8469,N_7359,N_6690);
nand U8470 (N_8470,N_6576,N_7023);
nor U8471 (N_8471,N_7497,N_6711);
nor U8472 (N_8472,N_6382,N_7222);
and U8473 (N_8473,N_7462,N_7280);
or U8474 (N_8474,N_7227,N_6252);
nand U8475 (N_8475,N_6858,N_6617);
nand U8476 (N_8476,N_6382,N_7322);
xnor U8477 (N_8477,N_7348,N_7065);
or U8478 (N_8478,N_7482,N_6775);
or U8479 (N_8479,N_6289,N_6303);
nor U8480 (N_8480,N_6760,N_6951);
and U8481 (N_8481,N_6935,N_6261);
nor U8482 (N_8482,N_6886,N_7394);
and U8483 (N_8483,N_6624,N_7287);
nor U8484 (N_8484,N_6948,N_7482);
xor U8485 (N_8485,N_6881,N_6781);
nor U8486 (N_8486,N_6800,N_6756);
and U8487 (N_8487,N_6769,N_7490);
xor U8488 (N_8488,N_7359,N_7479);
and U8489 (N_8489,N_6504,N_7357);
or U8490 (N_8490,N_7233,N_7161);
xor U8491 (N_8491,N_6328,N_6698);
and U8492 (N_8492,N_7399,N_6575);
and U8493 (N_8493,N_7275,N_6855);
and U8494 (N_8494,N_6882,N_7039);
or U8495 (N_8495,N_6607,N_7248);
and U8496 (N_8496,N_6772,N_6387);
and U8497 (N_8497,N_6919,N_7178);
nand U8498 (N_8498,N_7149,N_6384);
xnor U8499 (N_8499,N_6335,N_6838);
nand U8500 (N_8500,N_7010,N_7092);
or U8501 (N_8501,N_6405,N_6915);
nor U8502 (N_8502,N_7053,N_7282);
or U8503 (N_8503,N_7274,N_6270);
nor U8504 (N_8504,N_6562,N_6996);
nor U8505 (N_8505,N_6880,N_6294);
and U8506 (N_8506,N_6799,N_7208);
or U8507 (N_8507,N_7189,N_6269);
xnor U8508 (N_8508,N_6759,N_6293);
xor U8509 (N_8509,N_7372,N_7494);
or U8510 (N_8510,N_7111,N_6888);
or U8511 (N_8511,N_6294,N_6723);
nand U8512 (N_8512,N_6585,N_7299);
nand U8513 (N_8513,N_6555,N_6723);
nor U8514 (N_8514,N_7492,N_7168);
and U8515 (N_8515,N_7059,N_6463);
and U8516 (N_8516,N_7394,N_6482);
and U8517 (N_8517,N_6905,N_6365);
or U8518 (N_8518,N_7289,N_7134);
xor U8519 (N_8519,N_6442,N_6752);
nor U8520 (N_8520,N_6697,N_7425);
nand U8521 (N_8521,N_6708,N_6394);
xor U8522 (N_8522,N_6583,N_6457);
nand U8523 (N_8523,N_6600,N_7352);
nor U8524 (N_8524,N_6934,N_7110);
and U8525 (N_8525,N_6407,N_6360);
nor U8526 (N_8526,N_6448,N_6405);
or U8527 (N_8527,N_6945,N_6922);
and U8528 (N_8528,N_7242,N_6340);
or U8529 (N_8529,N_7406,N_6473);
nand U8530 (N_8530,N_6629,N_7249);
nand U8531 (N_8531,N_6480,N_7246);
and U8532 (N_8532,N_6976,N_6556);
and U8533 (N_8533,N_6259,N_7493);
or U8534 (N_8534,N_6680,N_6355);
and U8535 (N_8535,N_7003,N_6345);
or U8536 (N_8536,N_7394,N_7497);
xnor U8537 (N_8537,N_6870,N_6315);
and U8538 (N_8538,N_7320,N_7152);
nand U8539 (N_8539,N_6371,N_6324);
or U8540 (N_8540,N_6321,N_7489);
or U8541 (N_8541,N_6528,N_7238);
nand U8542 (N_8542,N_6761,N_6762);
nor U8543 (N_8543,N_7330,N_6958);
nand U8544 (N_8544,N_7349,N_6656);
or U8545 (N_8545,N_6972,N_6458);
and U8546 (N_8546,N_6496,N_6659);
nand U8547 (N_8547,N_6300,N_7117);
nand U8548 (N_8548,N_6780,N_6452);
or U8549 (N_8549,N_6831,N_6700);
xor U8550 (N_8550,N_6689,N_6617);
nand U8551 (N_8551,N_6811,N_6353);
nand U8552 (N_8552,N_6313,N_6465);
nand U8553 (N_8553,N_6638,N_7245);
and U8554 (N_8554,N_7400,N_6526);
or U8555 (N_8555,N_6300,N_6434);
xor U8556 (N_8556,N_7487,N_6421);
nand U8557 (N_8557,N_6690,N_6964);
or U8558 (N_8558,N_6708,N_7085);
nand U8559 (N_8559,N_6291,N_7247);
and U8560 (N_8560,N_6495,N_6673);
or U8561 (N_8561,N_6994,N_7135);
and U8562 (N_8562,N_6770,N_6767);
nor U8563 (N_8563,N_6332,N_7139);
nor U8564 (N_8564,N_6716,N_6939);
xnor U8565 (N_8565,N_7218,N_6592);
nand U8566 (N_8566,N_7368,N_6477);
nor U8567 (N_8567,N_7069,N_6643);
nand U8568 (N_8568,N_6541,N_6916);
or U8569 (N_8569,N_6878,N_6752);
nand U8570 (N_8570,N_6795,N_6448);
xor U8571 (N_8571,N_6402,N_7388);
and U8572 (N_8572,N_7346,N_6425);
nor U8573 (N_8573,N_6807,N_7130);
or U8574 (N_8574,N_7150,N_6382);
xnor U8575 (N_8575,N_6506,N_6359);
nand U8576 (N_8576,N_6856,N_7071);
or U8577 (N_8577,N_7279,N_6703);
or U8578 (N_8578,N_7062,N_6935);
and U8579 (N_8579,N_7319,N_7317);
or U8580 (N_8580,N_6898,N_6452);
and U8581 (N_8581,N_6557,N_6502);
nor U8582 (N_8582,N_7017,N_7071);
nand U8583 (N_8583,N_6261,N_7426);
and U8584 (N_8584,N_7277,N_6960);
nor U8585 (N_8585,N_7136,N_7278);
nand U8586 (N_8586,N_6312,N_7086);
or U8587 (N_8587,N_6909,N_7101);
nor U8588 (N_8588,N_7171,N_7220);
or U8589 (N_8589,N_6690,N_6626);
and U8590 (N_8590,N_6668,N_7338);
nor U8591 (N_8591,N_7285,N_6960);
nor U8592 (N_8592,N_6807,N_7151);
xnor U8593 (N_8593,N_7371,N_7443);
or U8594 (N_8594,N_7397,N_6867);
and U8595 (N_8595,N_6617,N_6941);
xor U8596 (N_8596,N_7184,N_6691);
or U8597 (N_8597,N_7424,N_7007);
and U8598 (N_8598,N_7131,N_7326);
or U8599 (N_8599,N_6660,N_6642);
nand U8600 (N_8600,N_7005,N_7073);
and U8601 (N_8601,N_7281,N_7167);
nand U8602 (N_8602,N_6911,N_6553);
xor U8603 (N_8603,N_7483,N_7309);
nor U8604 (N_8604,N_6690,N_6832);
nand U8605 (N_8605,N_6848,N_6861);
or U8606 (N_8606,N_6901,N_6328);
xnor U8607 (N_8607,N_7021,N_6872);
or U8608 (N_8608,N_7033,N_7261);
or U8609 (N_8609,N_6327,N_7048);
nor U8610 (N_8610,N_6348,N_6641);
nand U8611 (N_8611,N_7020,N_6846);
nand U8612 (N_8612,N_6843,N_7442);
or U8613 (N_8613,N_7022,N_7177);
xnor U8614 (N_8614,N_6809,N_6333);
nor U8615 (N_8615,N_7336,N_6743);
nand U8616 (N_8616,N_6951,N_6529);
nor U8617 (N_8617,N_6718,N_7481);
nor U8618 (N_8618,N_6954,N_6388);
and U8619 (N_8619,N_6347,N_7029);
xnor U8620 (N_8620,N_6496,N_6322);
xor U8621 (N_8621,N_7024,N_6735);
and U8622 (N_8622,N_7350,N_6641);
nand U8623 (N_8623,N_6808,N_6538);
nor U8624 (N_8624,N_7146,N_6645);
nand U8625 (N_8625,N_6523,N_6302);
nor U8626 (N_8626,N_6336,N_7152);
nand U8627 (N_8627,N_6596,N_7346);
or U8628 (N_8628,N_6900,N_6908);
xnor U8629 (N_8629,N_6272,N_7041);
nor U8630 (N_8630,N_7201,N_7180);
nand U8631 (N_8631,N_7251,N_6750);
xor U8632 (N_8632,N_6624,N_7044);
nand U8633 (N_8633,N_7194,N_6431);
nor U8634 (N_8634,N_6263,N_7277);
nand U8635 (N_8635,N_7125,N_6906);
nor U8636 (N_8636,N_6415,N_7241);
nand U8637 (N_8637,N_7316,N_6418);
or U8638 (N_8638,N_6533,N_7039);
nand U8639 (N_8639,N_6365,N_6561);
and U8640 (N_8640,N_7344,N_7015);
or U8641 (N_8641,N_6377,N_6449);
xnor U8642 (N_8642,N_6981,N_6898);
nor U8643 (N_8643,N_6372,N_7361);
and U8644 (N_8644,N_7358,N_6543);
and U8645 (N_8645,N_6691,N_6700);
or U8646 (N_8646,N_6339,N_6561);
xnor U8647 (N_8647,N_7096,N_7266);
nor U8648 (N_8648,N_7144,N_6362);
xnor U8649 (N_8649,N_6888,N_6597);
xnor U8650 (N_8650,N_6916,N_6949);
or U8651 (N_8651,N_7121,N_6788);
and U8652 (N_8652,N_6694,N_6664);
and U8653 (N_8653,N_6623,N_7237);
nand U8654 (N_8654,N_6789,N_7314);
and U8655 (N_8655,N_6833,N_6257);
nand U8656 (N_8656,N_6819,N_7018);
nand U8657 (N_8657,N_6737,N_7485);
xor U8658 (N_8658,N_6315,N_7020);
xnor U8659 (N_8659,N_7008,N_7021);
nand U8660 (N_8660,N_7409,N_7352);
nand U8661 (N_8661,N_7188,N_6807);
nor U8662 (N_8662,N_7262,N_6992);
nand U8663 (N_8663,N_7258,N_7107);
and U8664 (N_8664,N_7445,N_7458);
and U8665 (N_8665,N_6831,N_7445);
xnor U8666 (N_8666,N_7189,N_7265);
nand U8667 (N_8667,N_6908,N_6494);
nor U8668 (N_8668,N_7084,N_6713);
nor U8669 (N_8669,N_6780,N_7410);
and U8670 (N_8670,N_6364,N_6905);
nor U8671 (N_8671,N_6264,N_7304);
or U8672 (N_8672,N_6306,N_6970);
and U8673 (N_8673,N_6307,N_7304);
nand U8674 (N_8674,N_7313,N_6708);
nor U8675 (N_8675,N_7201,N_7008);
nand U8676 (N_8676,N_6851,N_6770);
xnor U8677 (N_8677,N_6834,N_7426);
nand U8678 (N_8678,N_7381,N_7211);
or U8679 (N_8679,N_6381,N_6902);
nand U8680 (N_8680,N_7366,N_7400);
nor U8681 (N_8681,N_6592,N_7037);
and U8682 (N_8682,N_6951,N_6868);
nor U8683 (N_8683,N_7104,N_7010);
nor U8684 (N_8684,N_7027,N_7153);
nor U8685 (N_8685,N_6963,N_7442);
xor U8686 (N_8686,N_6390,N_6435);
and U8687 (N_8687,N_7249,N_7453);
xnor U8688 (N_8688,N_6633,N_7274);
xnor U8689 (N_8689,N_7323,N_6932);
xor U8690 (N_8690,N_6324,N_7067);
nand U8691 (N_8691,N_7254,N_6309);
nor U8692 (N_8692,N_7223,N_6365);
xor U8693 (N_8693,N_6643,N_6955);
xor U8694 (N_8694,N_6819,N_7392);
or U8695 (N_8695,N_7306,N_6881);
or U8696 (N_8696,N_6292,N_7319);
and U8697 (N_8697,N_6371,N_7045);
or U8698 (N_8698,N_7227,N_7474);
xor U8699 (N_8699,N_7379,N_6735);
or U8700 (N_8700,N_7462,N_7384);
nor U8701 (N_8701,N_6924,N_7260);
xor U8702 (N_8702,N_7262,N_7160);
and U8703 (N_8703,N_6323,N_6443);
nand U8704 (N_8704,N_7170,N_7324);
and U8705 (N_8705,N_7092,N_7297);
nand U8706 (N_8706,N_6590,N_6653);
and U8707 (N_8707,N_6804,N_6842);
xnor U8708 (N_8708,N_6536,N_7444);
and U8709 (N_8709,N_7387,N_6324);
and U8710 (N_8710,N_7357,N_6853);
or U8711 (N_8711,N_7404,N_6529);
xnor U8712 (N_8712,N_7301,N_7126);
or U8713 (N_8713,N_7442,N_6794);
nand U8714 (N_8714,N_7050,N_7239);
xor U8715 (N_8715,N_6738,N_6443);
or U8716 (N_8716,N_7021,N_6397);
nor U8717 (N_8717,N_7456,N_6436);
xor U8718 (N_8718,N_6514,N_6834);
and U8719 (N_8719,N_6688,N_6565);
xnor U8720 (N_8720,N_6397,N_6906);
and U8721 (N_8721,N_7494,N_6513);
nor U8722 (N_8722,N_6532,N_6592);
or U8723 (N_8723,N_7137,N_6988);
nor U8724 (N_8724,N_7339,N_6290);
xor U8725 (N_8725,N_7182,N_7208);
xor U8726 (N_8726,N_7009,N_7381);
and U8727 (N_8727,N_7023,N_7208);
nand U8728 (N_8728,N_6860,N_6514);
xnor U8729 (N_8729,N_6570,N_6863);
or U8730 (N_8730,N_6576,N_6383);
xnor U8731 (N_8731,N_6424,N_6268);
nor U8732 (N_8732,N_6279,N_6408);
nor U8733 (N_8733,N_6716,N_6448);
xnor U8734 (N_8734,N_6852,N_7098);
nand U8735 (N_8735,N_7185,N_6672);
or U8736 (N_8736,N_7216,N_6506);
xnor U8737 (N_8737,N_6389,N_6804);
nand U8738 (N_8738,N_7417,N_7060);
nor U8739 (N_8739,N_6714,N_6761);
or U8740 (N_8740,N_7116,N_7288);
xnor U8741 (N_8741,N_7114,N_7269);
and U8742 (N_8742,N_6578,N_7436);
xnor U8743 (N_8743,N_7215,N_7331);
nand U8744 (N_8744,N_7126,N_6297);
xnor U8745 (N_8745,N_6368,N_6435);
nand U8746 (N_8746,N_6377,N_7404);
nor U8747 (N_8747,N_6920,N_7377);
nor U8748 (N_8748,N_6876,N_6787);
xor U8749 (N_8749,N_6612,N_6365);
and U8750 (N_8750,N_8597,N_8601);
and U8751 (N_8751,N_8087,N_7910);
xor U8752 (N_8752,N_8438,N_8512);
nor U8753 (N_8753,N_7606,N_8324);
nand U8754 (N_8754,N_7834,N_7529);
and U8755 (N_8755,N_8554,N_8568);
and U8756 (N_8756,N_7814,N_7991);
nor U8757 (N_8757,N_7706,N_7500);
nor U8758 (N_8758,N_8147,N_8581);
and U8759 (N_8759,N_8145,N_7601);
nor U8760 (N_8760,N_7528,N_7597);
nor U8761 (N_8761,N_8136,N_7930);
nor U8762 (N_8762,N_7824,N_7745);
and U8763 (N_8763,N_8281,N_8230);
and U8764 (N_8764,N_7716,N_7977);
xnor U8765 (N_8765,N_8081,N_7852);
and U8766 (N_8766,N_7623,N_8560);
nor U8767 (N_8767,N_8473,N_8090);
nand U8768 (N_8768,N_7857,N_7757);
nand U8769 (N_8769,N_7673,N_7940);
nor U8770 (N_8770,N_8507,N_8284);
and U8771 (N_8771,N_7925,N_8423);
nor U8772 (N_8772,N_7825,N_8579);
xnor U8773 (N_8773,N_8442,N_8315);
xnor U8774 (N_8774,N_8518,N_8550);
and U8775 (N_8775,N_7902,N_8207);
xor U8776 (N_8776,N_7622,N_7633);
nor U8777 (N_8777,N_7683,N_8298);
xor U8778 (N_8778,N_8001,N_7832);
and U8779 (N_8779,N_8437,N_7777);
and U8780 (N_8780,N_7908,N_7647);
and U8781 (N_8781,N_7955,N_7607);
xor U8782 (N_8782,N_8182,N_8338);
and U8783 (N_8783,N_8574,N_7617);
nand U8784 (N_8784,N_7867,N_7754);
or U8785 (N_8785,N_7714,N_7969);
nor U8786 (N_8786,N_8125,N_7533);
nand U8787 (N_8787,N_8365,N_8245);
and U8788 (N_8788,N_8282,N_8428);
xnor U8789 (N_8789,N_7888,N_8570);
nor U8790 (N_8790,N_8166,N_8174);
xor U8791 (N_8791,N_8701,N_8268);
nor U8792 (N_8792,N_7752,N_8356);
xor U8793 (N_8793,N_7621,N_8661);
or U8794 (N_8794,N_7891,N_8368);
nand U8795 (N_8795,N_7804,N_8580);
xor U8796 (N_8796,N_8474,N_8426);
or U8797 (N_8797,N_7643,N_8097);
xnor U8798 (N_8798,N_7799,N_8040);
nor U8799 (N_8799,N_8543,N_7996);
and U8800 (N_8800,N_7952,N_8618);
nand U8801 (N_8801,N_8456,N_8074);
nand U8802 (N_8802,N_8619,N_7510);
and U8803 (N_8803,N_7717,N_8140);
nor U8804 (N_8804,N_8314,N_8589);
and U8805 (N_8805,N_7759,N_8279);
and U8806 (N_8806,N_8533,N_8066);
xnor U8807 (N_8807,N_8340,N_7914);
xnor U8808 (N_8808,N_8471,N_8360);
xnor U8809 (N_8809,N_8736,N_8525);
xnor U8810 (N_8810,N_8121,N_8138);
xnor U8811 (N_8811,N_8400,N_8636);
xnor U8812 (N_8812,N_8034,N_8311);
or U8813 (N_8813,N_7736,N_7593);
xnor U8814 (N_8814,N_7722,N_8515);
or U8815 (N_8815,N_8189,N_7563);
nand U8816 (N_8816,N_7795,N_8466);
and U8817 (N_8817,N_7664,N_7515);
or U8818 (N_8818,N_8077,N_7587);
nand U8819 (N_8819,N_8007,N_8394);
nor U8820 (N_8820,N_7987,N_7794);
or U8821 (N_8821,N_8399,N_7599);
nor U8822 (N_8822,N_7655,N_8639);
nor U8823 (N_8823,N_7895,N_8123);
xnor U8824 (N_8824,N_8729,N_7924);
xor U8825 (N_8825,N_8208,N_7569);
nand U8826 (N_8826,N_7713,N_8130);
nand U8827 (N_8827,N_8067,N_7705);
and U8828 (N_8828,N_8645,N_8584);
xor U8829 (N_8829,N_7922,N_7815);
nor U8830 (N_8830,N_8531,N_8532);
nand U8831 (N_8831,N_7548,N_8609);
nor U8832 (N_8832,N_8627,N_8335);
nor U8833 (N_8833,N_7923,N_8452);
nand U8834 (N_8834,N_8369,N_7567);
nor U8835 (N_8835,N_8488,N_8553);
nor U8836 (N_8836,N_7506,N_8536);
and U8837 (N_8837,N_8716,N_7630);
nand U8838 (N_8838,N_8687,N_7734);
nor U8839 (N_8839,N_7628,N_8603);
xnor U8840 (N_8840,N_8563,N_8173);
nor U8841 (N_8841,N_8339,N_8239);
and U8842 (N_8842,N_8238,N_7792);
nor U8843 (N_8843,N_8705,N_7737);
xor U8844 (N_8844,N_8111,N_8495);
nand U8845 (N_8845,N_8472,N_8300);
nand U8846 (N_8846,N_8254,N_8384);
nand U8847 (N_8847,N_7819,N_7903);
or U8848 (N_8848,N_8707,N_7801);
and U8849 (N_8849,N_7964,N_7917);
and U8850 (N_8850,N_7820,N_8606);
or U8851 (N_8851,N_8629,N_8096);
and U8852 (N_8852,N_7844,N_8725);
nor U8853 (N_8853,N_7501,N_7720);
nand U8854 (N_8854,N_8421,N_8434);
and U8855 (N_8855,N_8212,N_7894);
or U8856 (N_8856,N_8391,N_7892);
nor U8857 (N_8857,N_8195,N_7579);
or U8858 (N_8858,N_8341,N_8075);
or U8859 (N_8859,N_8277,N_8592);
nor U8860 (N_8860,N_8010,N_7562);
nor U8861 (N_8861,N_7702,N_7645);
nor U8862 (N_8862,N_8699,N_8395);
nor U8863 (N_8863,N_8497,N_7707);
nor U8864 (N_8864,N_8477,N_7848);
nor U8865 (N_8865,N_7875,N_8005);
xor U8866 (N_8866,N_7543,N_8351);
and U8867 (N_8867,N_7604,N_7854);
nor U8868 (N_8868,N_7905,N_7840);
nor U8869 (N_8869,N_8662,N_8063);
or U8870 (N_8870,N_8722,N_7658);
nand U8871 (N_8871,N_8444,N_7810);
and U8872 (N_8872,N_8193,N_7670);
and U8873 (N_8873,N_8359,N_8743);
nand U8874 (N_8874,N_8000,N_8236);
or U8875 (N_8875,N_8401,N_7760);
nor U8876 (N_8876,N_8270,N_8711);
or U8877 (N_8877,N_8632,N_8388);
nor U8878 (N_8878,N_8158,N_8229);
nor U8879 (N_8879,N_8186,N_8732);
nor U8880 (N_8880,N_8735,N_7805);
xnor U8881 (N_8881,N_7758,N_8196);
nor U8882 (N_8882,N_7927,N_7790);
xor U8883 (N_8883,N_8069,N_8585);
and U8884 (N_8884,N_7519,N_8119);
nor U8885 (N_8885,N_7853,N_7976);
xnor U8886 (N_8886,N_7863,N_7571);
xnor U8887 (N_8887,N_8008,N_7984);
nand U8888 (N_8888,N_7975,N_7944);
xnor U8889 (N_8889,N_8458,N_8654);
xnor U8890 (N_8890,N_7700,N_8232);
or U8891 (N_8891,N_7635,N_8050);
nand U8892 (N_8892,N_7868,N_7511);
nand U8893 (N_8893,N_7773,N_8604);
and U8894 (N_8894,N_7786,N_8227);
and U8895 (N_8895,N_8266,N_8045);
or U8896 (N_8896,N_7711,N_7576);
xnor U8897 (N_8897,N_7999,N_8179);
xnor U8898 (N_8898,N_7751,N_7907);
or U8899 (N_8899,N_7674,N_8293);
xor U8900 (N_8900,N_8469,N_7833);
xnor U8901 (N_8901,N_8108,N_7989);
nor U8902 (N_8902,N_8332,N_7726);
nand U8903 (N_8903,N_7912,N_8556);
xor U8904 (N_8904,N_8551,N_8464);
xor U8905 (N_8905,N_8591,N_7697);
and U8906 (N_8906,N_7957,N_7514);
nor U8907 (N_8907,N_8415,N_8031);
nand U8908 (N_8908,N_7753,N_7524);
or U8909 (N_8909,N_8126,N_7710);
nor U8910 (N_8910,N_8708,N_7893);
or U8911 (N_8911,N_8514,N_8513);
or U8912 (N_8912,N_7943,N_8484);
xor U8913 (N_8913,N_7941,N_8749);
or U8914 (N_8914,N_8378,N_8188);
nand U8915 (N_8915,N_7849,N_7503);
or U8916 (N_8916,N_8025,N_8738);
and U8917 (N_8917,N_8500,N_7939);
and U8918 (N_8918,N_7998,N_8260);
nand U8919 (N_8919,N_8572,N_8046);
nand U8920 (N_8920,N_7882,N_7559);
or U8921 (N_8921,N_7967,N_8499);
nor U8922 (N_8922,N_7641,N_8567);
and U8923 (N_8923,N_7916,N_8455);
nor U8924 (N_8924,N_7803,N_8262);
or U8925 (N_8925,N_8614,N_8175);
and U8926 (N_8926,N_8163,N_8667);
and U8927 (N_8927,N_7948,N_8176);
or U8928 (N_8928,N_8476,N_7841);
xor U8929 (N_8929,N_8035,N_8521);
nand U8930 (N_8930,N_7701,N_7768);
xor U8931 (N_8931,N_7956,N_7592);
xnor U8932 (N_8932,N_8080,N_8712);
and U8933 (N_8933,N_8151,N_7909);
nor U8934 (N_8934,N_8068,N_7728);
xor U8935 (N_8935,N_8386,N_8573);
nand U8936 (N_8936,N_7818,N_8501);
nand U8937 (N_8937,N_8269,N_7693);
xnor U8938 (N_8938,N_8459,N_8747);
nand U8939 (N_8939,N_8213,N_8013);
nor U8940 (N_8940,N_7933,N_8586);
xnor U8941 (N_8941,N_8343,N_7850);
or U8942 (N_8942,N_8030,N_8660);
and U8943 (N_8943,N_8241,N_7703);
nor U8944 (N_8944,N_8730,N_8047);
nand U8945 (N_8945,N_7959,N_7890);
nor U8946 (N_8946,N_7974,N_8508);
nor U8947 (N_8947,N_8194,N_7618);
nand U8948 (N_8948,N_8146,N_7856);
xor U8949 (N_8949,N_8323,N_7535);
or U8950 (N_8950,N_8100,N_7942);
nand U8951 (N_8951,N_7920,N_7513);
and U8952 (N_8952,N_7546,N_8199);
and U8953 (N_8953,N_7675,N_7509);
nor U8954 (N_8954,N_8510,N_8362);
xor U8955 (N_8955,N_7631,N_8537);
nand U8956 (N_8956,N_8225,N_7522);
or U8957 (N_8957,N_7595,N_8682);
nand U8958 (N_8958,N_7672,N_8628);
xor U8959 (N_8959,N_8498,N_8546);
nor U8960 (N_8960,N_8683,N_7640);
or U8961 (N_8961,N_7541,N_8053);
nor U8962 (N_8962,N_8178,N_8036);
or U8963 (N_8963,N_7808,N_8374);
xor U8964 (N_8964,N_8337,N_7782);
or U8965 (N_8965,N_7538,N_8133);
or U8966 (N_8966,N_8624,N_7869);
or U8967 (N_8967,N_8183,N_8441);
and U8968 (N_8968,N_8114,N_8059);
xor U8969 (N_8969,N_8418,N_7564);
xor U8970 (N_8970,N_8596,N_8052);
and U8971 (N_8971,N_8680,N_8685);
and U8972 (N_8972,N_8168,N_8631);
nand U8973 (N_8973,N_8192,N_7858);
or U8974 (N_8974,N_8169,N_8242);
or U8975 (N_8975,N_7931,N_8427);
and U8976 (N_8976,N_7572,N_7960);
nor U8977 (N_8977,N_7911,N_8303);
nand U8978 (N_8978,N_7507,N_8302);
or U8979 (N_8979,N_7620,N_8430);
or U8980 (N_8980,N_8494,N_8544);
nor U8981 (N_8981,N_8433,N_8608);
or U8982 (N_8982,N_8669,N_8073);
nor U8983 (N_8983,N_8185,N_8659);
nand U8984 (N_8984,N_7687,N_7919);
and U8985 (N_8985,N_7721,N_8079);
nor U8986 (N_8986,N_8569,N_7744);
or U8987 (N_8987,N_7741,N_8061);
xnor U8988 (N_8988,N_7545,N_8594);
nor U8989 (N_8989,N_8617,N_7978);
nor U8990 (N_8990,N_8620,N_8478);
xor U8991 (N_8991,N_7611,N_8291);
and U8992 (N_8992,N_8354,N_8641);
nor U8993 (N_8993,N_7855,N_8390);
or U8994 (N_8994,N_7766,N_7740);
nor U8995 (N_8995,N_7531,N_8558);
xor U8996 (N_8996,N_7906,N_7523);
and U8997 (N_8997,N_8157,N_7921);
or U8998 (N_8998,N_8530,N_7554);
and U8999 (N_8999,N_8634,N_7756);
or U9000 (N_9000,N_7836,N_7870);
nand U9001 (N_9001,N_7504,N_7560);
nor U9002 (N_9002,N_7596,N_8723);
and U9003 (N_9003,N_7685,N_8668);
xor U9004 (N_9004,N_8042,N_8547);
nand U9005 (N_9005,N_8439,N_8425);
nand U9006 (N_9006,N_8342,N_8535);
or U9007 (N_9007,N_8258,N_8054);
nor U9008 (N_9008,N_8719,N_8656);
nor U9009 (N_9009,N_7667,N_8263);
or U9010 (N_9010,N_7694,N_8320);
xnor U9011 (N_9011,N_8529,N_7866);
nand U9012 (N_9012,N_8249,N_7696);
nand U9013 (N_9013,N_8246,N_8327);
nor U9014 (N_9014,N_8445,N_8144);
and U9015 (N_9015,N_8244,N_8648);
or U9016 (N_9016,N_7972,N_7695);
nor U9017 (N_9017,N_7719,N_7918);
xnor U9018 (N_9018,N_8116,N_8317);
nor U9019 (N_9019,N_7612,N_7521);
and U9020 (N_9020,N_8462,N_8237);
xnor U9021 (N_9021,N_8691,N_8152);
nor U9022 (N_9022,N_7778,N_7995);
and U9023 (N_9023,N_7973,N_8220);
or U9024 (N_9024,N_8435,N_7639);
nor U9025 (N_9025,N_7985,N_7838);
xnor U9026 (N_9026,N_7525,N_8102);
nand U9027 (N_9027,N_7632,N_8431);
or U9028 (N_9028,N_7835,N_7518);
and U9029 (N_9029,N_8124,N_8361);
and U9030 (N_9030,N_8409,N_8443);
nand U9031 (N_9031,N_8312,N_7520);
nand U9032 (N_9032,N_7662,N_8009);
nor U9033 (N_9033,N_8318,N_8664);
xnor U9034 (N_9034,N_8387,N_7874);
or U9035 (N_9035,N_8364,N_8223);
and U9036 (N_9036,N_8637,N_8110);
and U9037 (N_9037,N_8727,N_8467);
and U9038 (N_9038,N_8027,N_8329);
nor U9039 (N_9039,N_7516,N_8004);
xor U9040 (N_9040,N_7776,N_8625);
nor U9041 (N_9041,N_8502,N_8105);
nor U9042 (N_9042,N_8170,N_7979);
or U9043 (N_9043,N_8024,N_8275);
nor U9044 (N_9044,N_8306,N_8333);
nor U9045 (N_9045,N_8135,N_7530);
nand U9046 (N_9046,N_7627,N_7885);
and U9047 (N_9047,N_7755,N_8493);
nand U9048 (N_9048,N_8522,N_8653);
and U9049 (N_9049,N_7915,N_8742);
or U9050 (N_9050,N_7608,N_7556);
or U9051 (N_9051,N_7677,N_8267);
and U9052 (N_9052,N_7712,N_7679);
xnor U9053 (N_9053,N_7671,N_8049);
and U9054 (N_9054,N_7963,N_8099);
xnor U9055 (N_9055,N_8256,N_7692);
nor U9056 (N_9056,N_7809,N_7578);
nand U9057 (N_9057,N_7898,N_7536);
xor U9058 (N_9058,N_8156,N_8642);
and U9059 (N_9059,N_8447,N_7534);
xor U9060 (N_9060,N_8575,N_8516);
and U9061 (N_9061,N_8264,N_8429);
nor U9062 (N_9062,N_7889,N_8414);
nand U9063 (N_9063,N_8446,N_8453);
xnor U9064 (N_9064,N_8640,N_8307);
or U9065 (N_9065,N_8381,N_7644);
or U9066 (N_9066,N_8460,N_7602);
nand U9067 (N_9067,N_7651,N_7828);
nand U9068 (N_9068,N_7945,N_8419);
xor U9069 (N_9069,N_7686,N_8345);
and U9070 (N_9070,N_8039,N_7661);
xnor U9071 (N_9071,N_8564,N_8017);
or U9072 (N_9072,N_8688,N_8412);
or U9073 (N_9073,N_8588,N_8093);
xor U9074 (N_9074,N_8086,N_8583);
nand U9075 (N_9075,N_8154,N_8681);
xnor U9076 (N_9076,N_7880,N_7508);
xor U9077 (N_9077,N_7537,N_8150);
xor U9078 (N_9078,N_7738,N_8686);
nand U9079 (N_9079,N_8006,N_7993);
and U9080 (N_9080,N_8299,N_7730);
or U9081 (N_9081,N_8118,N_7680);
nor U9082 (N_9082,N_7724,N_7816);
nor U9083 (N_9083,N_8310,N_8247);
or U9084 (N_9084,N_7802,N_8692);
nand U9085 (N_9085,N_8250,N_8187);
nand U9086 (N_9086,N_8524,N_8094);
xnor U9087 (N_9087,N_8283,N_8630);
or U9088 (N_9088,N_8132,N_8612);
or U9089 (N_9089,N_8702,N_7864);
xnor U9090 (N_9090,N_8635,N_8417);
nand U9091 (N_9091,N_8131,N_8704);
and U9092 (N_9092,N_7542,N_7884);
or U9093 (N_9093,N_8503,N_8259);
xor U9094 (N_9094,N_8280,N_8600);
nor U9095 (N_9095,N_7544,N_8309);
xnor U9096 (N_9096,N_7709,N_7653);
xor U9097 (N_9097,N_8611,N_8257);
and U9098 (N_9098,N_7798,N_7552);
or U9099 (N_9099,N_8571,N_8355);
and U9100 (N_9100,N_8480,N_7772);
nand U9101 (N_9101,N_8101,N_7746);
xor U9102 (N_9102,N_8410,N_7550);
nor U9103 (N_9103,N_8191,N_8328);
xnor U9104 (N_9104,N_7555,N_8454);
and U9105 (N_9105,N_7565,N_8022);
and U9106 (N_9106,N_8545,N_8197);
nor U9107 (N_9107,N_7936,N_7698);
nor U9108 (N_9108,N_8714,N_7899);
or U9109 (N_9109,N_8370,N_8694);
nand U9110 (N_9110,N_8072,N_7600);
or U9111 (N_9111,N_7958,N_7742);
or U9112 (N_9112,N_7865,N_8643);
and U9113 (N_9113,N_8655,N_7512);
xnor U9114 (N_9114,N_7652,N_8398);
xor U9115 (N_9115,N_8511,N_8582);
or U9116 (N_9116,N_8289,N_8406);
nor U9117 (N_9117,N_8023,N_8709);
nor U9118 (N_9118,N_8098,N_7787);
xor U9119 (N_9119,N_7615,N_7904);
and U9120 (N_9120,N_8665,N_8161);
xor U9121 (N_9121,N_8465,N_8697);
and U9122 (N_9122,N_7770,N_8002);
and U9123 (N_9123,N_7876,N_8633);
and U9124 (N_9124,N_7642,N_8344);
nand U9125 (N_9125,N_8720,N_8647);
nand U9126 (N_9126,N_8103,N_8210);
nor U9127 (N_9127,N_7747,N_8095);
nor U9128 (N_9128,N_8235,N_8470);
nor U9129 (N_9129,N_8487,N_8055);
and U9130 (N_9130,N_7823,N_7551);
and U9131 (N_9131,N_8198,N_8448);
nand U9132 (N_9132,N_7937,N_7962);
and U9133 (N_9133,N_7613,N_8078);
nor U9134 (N_9134,N_8089,N_7764);
nor U9135 (N_9135,N_8703,N_7761);
nor U9136 (N_9136,N_7797,N_7605);
or U9137 (N_9137,N_7549,N_8319);
xor U9138 (N_9138,N_8693,N_8593);
and U9139 (N_9139,N_7980,N_8122);
and U9140 (N_9140,N_8221,N_8485);
or U9141 (N_9141,N_7624,N_8613);
nand U9142 (N_9142,N_8292,N_7769);
nand U9143 (N_9143,N_7763,N_7616);
xor U9144 (N_9144,N_8149,N_7900);
nand U9145 (N_9145,N_7791,N_7837);
and U9146 (N_9146,N_8565,N_8217);
nor U9147 (N_9147,N_7935,N_7558);
or U9148 (N_9148,N_8717,N_8367);
and U9149 (N_9149,N_8148,N_8605);
nor U9150 (N_9150,N_8308,N_8255);
nand U9151 (N_9151,N_7657,N_8112);
nor U9152 (N_9152,N_7575,N_8420);
nand U9153 (N_9153,N_8534,N_7946);
and U9154 (N_9154,N_7826,N_8721);
xor U9155 (N_9155,N_8357,N_7750);
or U9156 (N_9156,N_8162,N_8626);
or U9157 (N_9157,N_8422,N_8083);
xnor U9158 (N_9158,N_8517,N_7926);
xor U9159 (N_9159,N_8286,N_8646);
nand U9160 (N_9160,N_7847,N_7663);
and U9161 (N_9161,N_8058,N_7775);
xnor U9162 (N_9162,N_8542,N_8739);
and U9163 (N_9163,N_8128,N_8644);
and U9164 (N_9164,N_8253,N_8224);
nor U9165 (N_9165,N_8167,N_7669);
nand U9166 (N_9166,N_7660,N_8411);
nand U9167 (N_9167,N_8348,N_8143);
nor U9168 (N_9168,N_8372,N_8424);
nor U9169 (N_9169,N_8610,N_8538);
xnor U9170 (N_9170,N_8038,N_8689);
or U9171 (N_9171,N_8084,N_8638);
nor U9172 (N_9172,N_8741,N_8134);
or U9173 (N_9173,N_8177,N_7708);
and U9174 (N_9174,N_8385,N_7934);
and U9175 (N_9175,N_7594,N_8290);
or U9176 (N_9176,N_8621,N_8490);
nor U9177 (N_9177,N_8475,N_8233);
and U9178 (N_9178,N_8171,N_8203);
or U9179 (N_9179,N_8206,N_7928);
and U9180 (N_9180,N_8350,N_8295);
and U9181 (N_9181,N_8461,N_7965);
or U9182 (N_9182,N_8113,N_8276);
and U9183 (N_9183,N_7585,N_8380);
or U9184 (N_9184,N_8407,N_7743);
nor U9185 (N_9185,N_7699,N_7811);
and U9186 (N_9186,N_7582,N_7648);
or U9187 (N_9187,N_7887,N_7527);
xor U9188 (N_9188,N_7843,N_7765);
and U9189 (N_9189,N_8020,N_8032);
or U9190 (N_9190,N_7966,N_8200);
nor U9191 (N_9191,N_8676,N_8451);
and U9192 (N_9192,N_8261,N_8559);
or U9193 (N_9193,N_8043,N_8109);
nand U9194 (N_9194,N_8012,N_8375);
or U9195 (N_9195,N_8598,N_7793);
and U9196 (N_9196,N_8048,N_8623);
xnor U9197 (N_9197,N_8595,N_7951);
and U9198 (N_9198,N_8748,N_8142);
nor U9199 (N_9199,N_8363,N_8321);
or U9200 (N_9200,N_8745,N_8599);
xor U9201 (N_9201,N_8670,N_7739);
nor U9202 (N_9202,N_8003,N_8731);
xor U9203 (N_9203,N_8070,N_7704);
or U9204 (N_9204,N_8226,N_7983);
xor U9205 (N_9205,N_8440,N_8519);
xor U9206 (N_9206,N_8288,N_8706);
nor U9207 (N_9207,N_7584,N_8287);
nand U9208 (N_9208,N_7813,N_8353);
nor U9209 (N_9209,N_8160,N_8204);
xnor U9210 (N_9210,N_8071,N_8377);
nor U9211 (N_9211,N_7668,N_8127);
and U9212 (N_9212,N_8479,N_8540);
and U9213 (N_9213,N_8486,N_7654);
or U9214 (N_9214,N_7532,N_7727);
xor U9215 (N_9215,N_7636,N_7566);
or U9216 (N_9216,N_8155,N_8726);
xnor U9217 (N_9217,N_7970,N_8349);
and U9218 (N_9218,N_8615,N_7817);
xor U9219 (N_9219,N_7505,N_8371);
and U9220 (N_9220,N_8392,N_7517);
nor U9221 (N_9221,N_8404,N_7845);
nand U9222 (N_9222,N_7583,N_8322);
xor U9223 (N_9223,N_8744,N_7732);
nor U9224 (N_9224,N_7547,N_7961);
nor U9225 (N_9225,N_8164,N_8352);
nor U9226 (N_9226,N_7878,N_7689);
nor U9227 (N_9227,N_8265,N_8506);
xnor U9228 (N_9228,N_7950,N_7733);
and U9229 (N_9229,N_8622,N_8405);
nand U9230 (N_9230,N_7789,N_8184);
nor U9231 (N_9231,N_8389,N_7992);
xor U9232 (N_9232,N_8561,N_7881);
nand U9233 (N_9233,N_7540,N_7986);
nor U9234 (N_9234,N_8373,N_7568);
or U9235 (N_9235,N_7862,N_8740);
or U9236 (N_9236,N_8278,N_8679);
nor U9237 (N_9237,N_8033,N_8297);
nand U9238 (N_9238,N_7591,N_7896);
xor U9239 (N_9239,N_8607,N_8092);
xor U9240 (N_9240,N_7767,N_8029);
or U9241 (N_9241,N_8408,N_8234);
or U9242 (N_9242,N_8690,N_7609);
and U9243 (N_9243,N_7598,N_8416);
nor U9244 (N_9244,N_7988,N_8520);
or U9245 (N_9245,N_7812,N_7678);
and U9246 (N_9246,N_8021,N_7577);
or U9247 (N_9247,N_8076,N_7861);
or U9248 (N_9248,N_8737,N_8541);
and U9249 (N_9249,N_8305,N_7897);
xnor U9250 (N_9250,N_7806,N_8139);
xnor U9251 (N_9251,N_8436,N_7859);
and U9252 (N_9252,N_7610,N_8091);
nand U9253 (N_9253,N_8019,N_7589);
nor U9254 (N_9254,N_7827,N_7581);
and U9255 (N_9255,N_7779,N_8733);
xnor U9256 (N_9256,N_8468,N_7553);
or U9257 (N_9257,N_8334,N_8523);
or U9258 (N_9258,N_7748,N_8296);
or U9259 (N_9259,N_8011,N_7557);
or U9260 (N_9260,N_8057,N_8028);
nand U9261 (N_9261,N_7603,N_8016);
and U9262 (N_9262,N_8713,N_8539);
nand U9263 (N_9263,N_8379,N_7997);
nor U9264 (N_9264,N_7586,N_8153);
nand U9265 (N_9265,N_8082,N_7949);
xor U9266 (N_9266,N_7731,N_7851);
and U9267 (N_9267,N_8190,N_7646);
nand U9268 (N_9268,N_8590,N_8273);
xor U9269 (N_9269,N_7929,N_8014);
nand U9270 (N_9270,N_8674,N_8649);
nor U9271 (N_9271,N_8347,N_8172);
nor U9272 (N_9272,N_8678,N_7539);
or U9273 (N_9273,N_8215,N_7691);
or U9274 (N_9274,N_8746,N_7800);
and U9275 (N_9275,N_8313,N_7681);
nand U9276 (N_9276,N_8141,N_7723);
xor U9277 (N_9277,N_8271,N_7666);
xor U9278 (N_9278,N_8718,N_7682);
nand U9279 (N_9279,N_7883,N_8549);
and U9280 (N_9280,N_8576,N_8566);
or U9281 (N_9281,N_8088,N_8165);
xor U9282 (N_9282,N_8650,N_7784);
xor U9283 (N_9283,N_8181,N_8666);
nand U9284 (N_9284,N_8673,N_8684);
and U9285 (N_9285,N_8180,N_7574);
and U9286 (N_9286,N_8728,N_8715);
or U9287 (N_9287,N_7688,N_8677);
and U9288 (N_9288,N_7947,N_8231);
nor U9289 (N_9289,N_7762,N_7879);
or U9290 (N_9290,N_7872,N_7807);
nand U9291 (N_9291,N_7638,N_8129);
xor U9292 (N_9292,N_8432,N_8457);
and U9293 (N_9293,N_8285,N_7982);
and U9294 (N_9294,N_8734,N_8336);
nand U9295 (N_9295,N_7842,N_7877);
nand U9296 (N_9296,N_8304,N_8015);
xor U9297 (N_9297,N_7526,N_7774);
nor U9298 (N_9298,N_8657,N_7676);
nand U9299 (N_9299,N_7871,N_8228);
and U9300 (N_9300,N_8710,N_7649);
nand U9301 (N_9301,N_7829,N_8492);
or U9302 (N_9302,N_8274,N_7725);
nand U9303 (N_9303,N_7788,N_7846);
or U9304 (N_9304,N_7932,N_8366);
and U9305 (N_9305,N_7994,N_8209);
nor U9306 (N_9306,N_7637,N_8060);
xor U9307 (N_9307,N_8402,N_7971);
nand U9308 (N_9308,N_7783,N_8526);
nor U9309 (N_9309,N_8251,N_8555);
xor U9310 (N_9310,N_8672,N_7968);
or U9311 (N_9311,N_8294,N_7735);
nand U9312 (N_9312,N_7570,N_8330);
or U9313 (N_9313,N_7656,N_8698);
nand U9314 (N_9314,N_8700,N_8346);
xnor U9315 (N_9315,N_7831,N_8301);
nand U9316 (N_9316,N_8240,N_8159);
nor U9317 (N_9317,N_8115,N_7981);
and U9318 (N_9318,N_8219,N_7901);
nor U9319 (N_9319,N_8316,N_8107);
or U9320 (N_9320,N_7629,N_8137);
or U9321 (N_9321,N_7822,N_8062);
nand U9322 (N_9322,N_8449,N_7780);
and U9323 (N_9323,N_7873,N_8117);
nand U9324 (N_9324,N_8562,N_7650);
and U9325 (N_9325,N_8397,N_8671);
or U9326 (N_9326,N_8383,N_8587);
nand U9327 (N_9327,N_8382,N_7860);
xor U9328 (N_9328,N_8548,N_8041);
and U9329 (N_9329,N_8044,N_8651);
or U9330 (N_9330,N_8652,N_7913);
and U9331 (N_9331,N_8663,N_8325);
or U9332 (N_9332,N_8326,N_7634);
nor U9333 (N_9333,N_8557,N_8695);
and U9334 (N_9334,N_7590,N_7588);
and U9335 (N_9335,N_8483,N_8202);
nor U9336 (N_9336,N_8243,N_8026);
nand U9337 (N_9337,N_8413,N_8489);
or U9338 (N_9338,N_7715,N_8106);
nand U9339 (N_9339,N_8504,N_8205);
xor U9340 (N_9340,N_8201,N_8216);
or U9341 (N_9341,N_7839,N_7665);
nor U9342 (N_9342,N_7796,N_7573);
nand U9343 (N_9343,N_8577,N_8272);
or U9344 (N_9344,N_8602,N_8065);
xor U9345 (N_9345,N_8481,N_7938);
nand U9346 (N_9346,N_8214,N_8482);
xor U9347 (N_9347,N_8527,N_7729);
or U9348 (N_9348,N_8396,N_7785);
xnor U9349 (N_9349,N_7886,N_8696);
and U9350 (N_9350,N_7781,N_8056);
and U9351 (N_9351,N_8222,N_8463);
nor U9352 (N_9352,N_8252,N_7659);
xor U9353 (N_9353,N_8358,N_8248);
and U9354 (N_9354,N_7625,N_8211);
nand U9355 (N_9355,N_8064,N_8496);
nand U9356 (N_9356,N_8509,N_7718);
and U9357 (N_9357,N_8120,N_8104);
or U9358 (N_9358,N_7614,N_8393);
nand U9359 (N_9359,N_8724,N_8037);
and U9360 (N_9360,N_8528,N_8675);
nor U9361 (N_9361,N_7821,N_8085);
and U9362 (N_9362,N_8376,N_7561);
nand U9363 (N_9363,N_8403,N_8505);
xor U9364 (N_9364,N_7953,N_8331);
and U9365 (N_9365,N_8218,N_8051);
nor U9366 (N_9366,N_8658,N_8018);
xnor U9367 (N_9367,N_7502,N_7684);
and U9368 (N_9368,N_7619,N_8552);
nand U9369 (N_9369,N_7580,N_8578);
or U9370 (N_9370,N_8491,N_8450);
nor U9371 (N_9371,N_7749,N_7771);
and U9372 (N_9372,N_7626,N_7830);
or U9373 (N_9373,N_7690,N_7990);
and U9374 (N_9374,N_8616,N_7954);
or U9375 (N_9375,N_7592,N_8682);
nor U9376 (N_9376,N_8093,N_8728);
nand U9377 (N_9377,N_7700,N_7747);
xnor U9378 (N_9378,N_7816,N_8005);
nor U9379 (N_9379,N_7545,N_8263);
or U9380 (N_9380,N_7581,N_8132);
nand U9381 (N_9381,N_8485,N_7632);
and U9382 (N_9382,N_7952,N_8419);
and U9383 (N_9383,N_8206,N_8584);
nand U9384 (N_9384,N_8545,N_8368);
xnor U9385 (N_9385,N_8723,N_8618);
nand U9386 (N_9386,N_7971,N_8326);
or U9387 (N_9387,N_7933,N_8618);
or U9388 (N_9388,N_7626,N_7709);
or U9389 (N_9389,N_8320,N_8262);
xor U9390 (N_9390,N_8226,N_7882);
and U9391 (N_9391,N_7849,N_7538);
nand U9392 (N_9392,N_8466,N_8736);
or U9393 (N_9393,N_8727,N_8186);
or U9394 (N_9394,N_8411,N_7902);
nor U9395 (N_9395,N_8280,N_7784);
nand U9396 (N_9396,N_8686,N_7993);
and U9397 (N_9397,N_7742,N_8499);
nor U9398 (N_9398,N_7683,N_7891);
nor U9399 (N_9399,N_7952,N_8211);
nor U9400 (N_9400,N_8223,N_8350);
nand U9401 (N_9401,N_7991,N_7528);
and U9402 (N_9402,N_8676,N_8050);
and U9403 (N_9403,N_7707,N_8334);
or U9404 (N_9404,N_8180,N_8022);
nor U9405 (N_9405,N_8181,N_8154);
or U9406 (N_9406,N_8116,N_7908);
xnor U9407 (N_9407,N_8288,N_8293);
nor U9408 (N_9408,N_8196,N_8024);
nand U9409 (N_9409,N_8498,N_7810);
and U9410 (N_9410,N_8058,N_8259);
nor U9411 (N_9411,N_8484,N_8558);
nand U9412 (N_9412,N_7926,N_7809);
nor U9413 (N_9413,N_7940,N_7874);
nor U9414 (N_9414,N_8489,N_8326);
or U9415 (N_9415,N_8222,N_8326);
nor U9416 (N_9416,N_8295,N_8065);
or U9417 (N_9417,N_8459,N_8216);
or U9418 (N_9418,N_7895,N_8606);
nand U9419 (N_9419,N_7599,N_7804);
and U9420 (N_9420,N_8617,N_7513);
nand U9421 (N_9421,N_8748,N_8377);
xor U9422 (N_9422,N_7963,N_7891);
and U9423 (N_9423,N_7781,N_8714);
and U9424 (N_9424,N_8627,N_7939);
nand U9425 (N_9425,N_8232,N_7739);
xnor U9426 (N_9426,N_7936,N_8233);
nor U9427 (N_9427,N_8745,N_8253);
nor U9428 (N_9428,N_7585,N_8447);
or U9429 (N_9429,N_8544,N_8408);
nand U9430 (N_9430,N_7624,N_8339);
nand U9431 (N_9431,N_8017,N_7978);
nand U9432 (N_9432,N_8612,N_8096);
and U9433 (N_9433,N_8603,N_8548);
and U9434 (N_9434,N_7654,N_8624);
nor U9435 (N_9435,N_7879,N_8439);
xor U9436 (N_9436,N_7597,N_7956);
nor U9437 (N_9437,N_8032,N_7723);
or U9438 (N_9438,N_8681,N_7762);
xnor U9439 (N_9439,N_7639,N_7778);
and U9440 (N_9440,N_8586,N_8592);
xor U9441 (N_9441,N_8030,N_8145);
nor U9442 (N_9442,N_7531,N_8650);
nor U9443 (N_9443,N_7687,N_7796);
nand U9444 (N_9444,N_8643,N_7541);
nand U9445 (N_9445,N_8302,N_8388);
and U9446 (N_9446,N_7567,N_7772);
nand U9447 (N_9447,N_8366,N_8729);
nand U9448 (N_9448,N_8331,N_7835);
xor U9449 (N_9449,N_7653,N_7900);
xnor U9450 (N_9450,N_8524,N_7616);
nor U9451 (N_9451,N_8478,N_8568);
nor U9452 (N_9452,N_8026,N_7749);
or U9453 (N_9453,N_8041,N_8573);
and U9454 (N_9454,N_8048,N_8577);
nand U9455 (N_9455,N_7781,N_7715);
xor U9456 (N_9456,N_8568,N_7655);
nor U9457 (N_9457,N_7585,N_7867);
xnor U9458 (N_9458,N_8564,N_7590);
and U9459 (N_9459,N_8235,N_7860);
nor U9460 (N_9460,N_8205,N_7924);
xor U9461 (N_9461,N_7651,N_7720);
nand U9462 (N_9462,N_8390,N_8683);
nor U9463 (N_9463,N_7590,N_8043);
or U9464 (N_9464,N_7863,N_8003);
or U9465 (N_9465,N_7887,N_7745);
and U9466 (N_9466,N_8412,N_7665);
nand U9467 (N_9467,N_7874,N_8118);
and U9468 (N_9468,N_7681,N_7865);
and U9469 (N_9469,N_8646,N_8645);
or U9470 (N_9470,N_7778,N_7597);
xnor U9471 (N_9471,N_7979,N_7807);
and U9472 (N_9472,N_7656,N_8695);
xor U9473 (N_9473,N_7657,N_8283);
nand U9474 (N_9474,N_8674,N_7665);
nor U9475 (N_9475,N_8288,N_8298);
and U9476 (N_9476,N_8420,N_8195);
xnor U9477 (N_9477,N_7732,N_7664);
nor U9478 (N_9478,N_8224,N_8630);
and U9479 (N_9479,N_8041,N_7640);
xor U9480 (N_9480,N_7776,N_8112);
or U9481 (N_9481,N_8296,N_8432);
or U9482 (N_9482,N_8544,N_8438);
nand U9483 (N_9483,N_8034,N_8723);
nor U9484 (N_9484,N_8445,N_8278);
or U9485 (N_9485,N_8298,N_7600);
and U9486 (N_9486,N_8732,N_8303);
xnor U9487 (N_9487,N_8363,N_7853);
and U9488 (N_9488,N_8151,N_7811);
xnor U9489 (N_9489,N_8347,N_8212);
or U9490 (N_9490,N_8301,N_8657);
nor U9491 (N_9491,N_8643,N_8019);
or U9492 (N_9492,N_8747,N_8098);
nor U9493 (N_9493,N_7883,N_7564);
nor U9494 (N_9494,N_8418,N_7922);
nand U9495 (N_9495,N_8299,N_8066);
and U9496 (N_9496,N_7671,N_7828);
nor U9497 (N_9497,N_8224,N_8068);
or U9498 (N_9498,N_8076,N_7552);
and U9499 (N_9499,N_7957,N_7790);
or U9500 (N_9500,N_7997,N_8242);
or U9501 (N_9501,N_8009,N_7584);
and U9502 (N_9502,N_8308,N_8161);
and U9503 (N_9503,N_7991,N_8563);
nand U9504 (N_9504,N_8380,N_8118);
and U9505 (N_9505,N_8659,N_7931);
nand U9506 (N_9506,N_8241,N_8596);
nand U9507 (N_9507,N_7980,N_8675);
or U9508 (N_9508,N_8236,N_8573);
nand U9509 (N_9509,N_8317,N_8198);
or U9510 (N_9510,N_8249,N_8558);
or U9511 (N_9511,N_7865,N_8286);
or U9512 (N_9512,N_7828,N_7512);
nand U9513 (N_9513,N_8322,N_8290);
nor U9514 (N_9514,N_7566,N_8479);
xnor U9515 (N_9515,N_8738,N_7942);
nand U9516 (N_9516,N_7759,N_8435);
or U9517 (N_9517,N_8459,N_7502);
xnor U9518 (N_9518,N_7838,N_7557);
and U9519 (N_9519,N_8529,N_7570);
and U9520 (N_9520,N_8465,N_8029);
and U9521 (N_9521,N_7850,N_8556);
nand U9522 (N_9522,N_7976,N_7670);
nand U9523 (N_9523,N_8315,N_8338);
nand U9524 (N_9524,N_8134,N_7928);
nand U9525 (N_9525,N_7883,N_8273);
nor U9526 (N_9526,N_8486,N_8324);
xor U9527 (N_9527,N_8602,N_8018);
nand U9528 (N_9528,N_8205,N_8362);
or U9529 (N_9529,N_8041,N_8420);
nand U9530 (N_9530,N_7590,N_8643);
or U9531 (N_9531,N_7899,N_8350);
nand U9532 (N_9532,N_7556,N_8053);
nor U9533 (N_9533,N_7879,N_8697);
nand U9534 (N_9534,N_8651,N_7974);
xor U9535 (N_9535,N_8345,N_8362);
or U9536 (N_9536,N_8319,N_8545);
or U9537 (N_9537,N_7733,N_7884);
nor U9538 (N_9538,N_8652,N_7971);
or U9539 (N_9539,N_8656,N_8383);
nand U9540 (N_9540,N_7619,N_8301);
nand U9541 (N_9541,N_7950,N_7509);
nor U9542 (N_9542,N_7630,N_8182);
nand U9543 (N_9543,N_7657,N_8646);
or U9544 (N_9544,N_7660,N_7991);
nand U9545 (N_9545,N_8291,N_8401);
and U9546 (N_9546,N_8634,N_8601);
and U9547 (N_9547,N_8205,N_8744);
xor U9548 (N_9548,N_8683,N_8222);
and U9549 (N_9549,N_7903,N_7660);
xor U9550 (N_9550,N_7771,N_8706);
nand U9551 (N_9551,N_8236,N_8049);
nor U9552 (N_9552,N_8575,N_7694);
nor U9553 (N_9553,N_7768,N_7666);
and U9554 (N_9554,N_7905,N_8252);
and U9555 (N_9555,N_8059,N_8367);
nor U9556 (N_9556,N_7839,N_8049);
or U9557 (N_9557,N_7779,N_8415);
xnor U9558 (N_9558,N_7736,N_7699);
or U9559 (N_9559,N_8436,N_7826);
nor U9560 (N_9560,N_8170,N_8064);
and U9561 (N_9561,N_7792,N_8560);
nand U9562 (N_9562,N_8250,N_8588);
nand U9563 (N_9563,N_8077,N_8038);
or U9564 (N_9564,N_8275,N_7674);
nor U9565 (N_9565,N_8612,N_7676);
xnor U9566 (N_9566,N_8229,N_7509);
or U9567 (N_9567,N_8386,N_7717);
and U9568 (N_9568,N_8474,N_8681);
xnor U9569 (N_9569,N_7603,N_7630);
nand U9570 (N_9570,N_8190,N_8076);
nand U9571 (N_9571,N_8565,N_7617);
nand U9572 (N_9572,N_7620,N_7547);
and U9573 (N_9573,N_8487,N_7519);
nand U9574 (N_9574,N_7988,N_8309);
nor U9575 (N_9575,N_7597,N_8711);
or U9576 (N_9576,N_7547,N_7719);
or U9577 (N_9577,N_8527,N_8275);
or U9578 (N_9578,N_8510,N_8260);
and U9579 (N_9579,N_7625,N_8183);
and U9580 (N_9580,N_8185,N_8351);
nand U9581 (N_9581,N_7596,N_7687);
nand U9582 (N_9582,N_8425,N_8285);
nand U9583 (N_9583,N_8144,N_7548);
xor U9584 (N_9584,N_8534,N_7795);
nand U9585 (N_9585,N_7533,N_8625);
nand U9586 (N_9586,N_8343,N_8053);
nand U9587 (N_9587,N_7639,N_7695);
nor U9588 (N_9588,N_7713,N_7521);
nor U9589 (N_9589,N_7947,N_8521);
nor U9590 (N_9590,N_8723,N_8101);
nand U9591 (N_9591,N_7882,N_8203);
and U9592 (N_9592,N_8476,N_8430);
xnor U9593 (N_9593,N_7543,N_7878);
and U9594 (N_9594,N_7765,N_8726);
nor U9595 (N_9595,N_7949,N_7559);
xor U9596 (N_9596,N_7649,N_8488);
nand U9597 (N_9597,N_8188,N_8439);
nand U9598 (N_9598,N_8507,N_7667);
nor U9599 (N_9599,N_8729,N_8071);
xnor U9600 (N_9600,N_8310,N_7981);
and U9601 (N_9601,N_8266,N_7565);
nor U9602 (N_9602,N_7775,N_7585);
xnor U9603 (N_9603,N_8396,N_7741);
nand U9604 (N_9604,N_8517,N_7690);
and U9605 (N_9605,N_8165,N_8196);
nor U9606 (N_9606,N_8142,N_8400);
or U9607 (N_9607,N_8215,N_8422);
or U9608 (N_9608,N_8424,N_8508);
xor U9609 (N_9609,N_8553,N_8125);
or U9610 (N_9610,N_8275,N_8714);
or U9611 (N_9611,N_8383,N_8101);
nand U9612 (N_9612,N_8604,N_7538);
xor U9613 (N_9613,N_7878,N_8077);
xnor U9614 (N_9614,N_8257,N_8541);
nor U9615 (N_9615,N_8521,N_8253);
nand U9616 (N_9616,N_7719,N_8612);
nor U9617 (N_9617,N_8310,N_8411);
nor U9618 (N_9618,N_7611,N_7541);
nand U9619 (N_9619,N_7501,N_8183);
and U9620 (N_9620,N_8476,N_8089);
or U9621 (N_9621,N_7949,N_8030);
and U9622 (N_9622,N_8604,N_8331);
xnor U9623 (N_9623,N_8044,N_8058);
xnor U9624 (N_9624,N_8419,N_8221);
or U9625 (N_9625,N_8361,N_8366);
nor U9626 (N_9626,N_8014,N_7674);
nor U9627 (N_9627,N_7882,N_7570);
xnor U9628 (N_9628,N_7982,N_8318);
nor U9629 (N_9629,N_7844,N_8703);
xnor U9630 (N_9630,N_8505,N_7989);
nor U9631 (N_9631,N_7677,N_7942);
xnor U9632 (N_9632,N_7807,N_8530);
xor U9633 (N_9633,N_8427,N_8438);
and U9634 (N_9634,N_8209,N_7684);
and U9635 (N_9635,N_8202,N_8520);
and U9636 (N_9636,N_8622,N_8501);
xor U9637 (N_9637,N_8710,N_8725);
nor U9638 (N_9638,N_8537,N_8045);
and U9639 (N_9639,N_7610,N_8273);
or U9640 (N_9640,N_8705,N_8150);
nand U9641 (N_9641,N_8035,N_8426);
and U9642 (N_9642,N_8311,N_7833);
nand U9643 (N_9643,N_8495,N_8600);
xnor U9644 (N_9644,N_7945,N_8615);
and U9645 (N_9645,N_7790,N_7940);
nand U9646 (N_9646,N_7787,N_8010);
and U9647 (N_9647,N_8046,N_8441);
or U9648 (N_9648,N_8175,N_8153);
and U9649 (N_9649,N_7737,N_7717);
and U9650 (N_9650,N_8455,N_7714);
and U9651 (N_9651,N_7634,N_8567);
nand U9652 (N_9652,N_7799,N_8645);
nor U9653 (N_9653,N_8284,N_7705);
and U9654 (N_9654,N_8487,N_8398);
nand U9655 (N_9655,N_7764,N_8220);
nand U9656 (N_9656,N_7535,N_8396);
nor U9657 (N_9657,N_7757,N_8084);
nand U9658 (N_9658,N_8359,N_8607);
nor U9659 (N_9659,N_8382,N_8304);
xor U9660 (N_9660,N_8037,N_8571);
and U9661 (N_9661,N_7505,N_8693);
nand U9662 (N_9662,N_8572,N_7684);
nand U9663 (N_9663,N_7931,N_7512);
xor U9664 (N_9664,N_7891,N_7835);
xor U9665 (N_9665,N_8408,N_7921);
nor U9666 (N_9666,N_8653,N_8680);
and U9667 (N_9667,N_7847,N_8273);
or U9668 (N_9668,N_8456,N_7551);
or U9669 (N_9669,N_8581,N_8555);
xor U9670 (N_9670,N_8187,N_8002);
or U9671 (N_9671,N_8171,N_7641);
or U9672 (N_9672,N_7524,N_8390);
xor U9673 (N_9673,N_8105,N_8715);
and U9674 (N_9674,N_8135,N_8505);
nor U9675 (N_9675,N_7720,N_8391);
or U9676 (N_9676,N_7708,N_7998);
or U9677 (N_9677,N_8334,N_8566);
nand U9678 (N_9678,N_7769,N_7655);
nor U9679 (N_9679,N_7970,N_8545);
or U9680 (N_9680,N_8419,N_7862);
nor U9681 (N_9681,N_7827,N_8122);
xor U9682 (N_9682,N_7853,N_8464);
nand U9683 (N_9683,N_8715,N_8281);
or U9684 (N_9684,N_8247,N_7556);
nand U9685 (N_9685,N_8062,N_8618);
nand U9686 (N_9686,N_8747,N_8283);
nor U9687 (N_9687,N_7544,N_8485);
nand U9688 (N_9688,N_7784,N_8674);
nor U9689 (N_9689,N_8400,N_7961);
nor U9690 (N_9690,N_7626,N_8262);
or U9691 (N_9691,N_8186,N_8674);
nor U9692 (N_9692,N_8163,N_7790);
and U9693 (N_9693,N_7683,N_8364);
xor U9694 (N_9694,N_8443,N_8535);
and U9695 (N_9695,N_7803,N_8729);
and U9696 (N_9696,N_7582,N_8262);
and U9697 (N_9697,N_8689,N_8328);
nor U9698 (N_9698,N_7676,N_7551);
nand U9699 (N_9699,N_8335,N_7935);
or U9700 (N_9700,N_7811,N_8287);
nor U9701 (N_9701,N_7847,N_7579);
xor U9702 (N_9702,N_8204,N_7927);
nor U9703 (N_9703,N_8617,N_8258);
and U9704 (N_9704,N_8538,N_8185);
xor U9705 (N_9705,N_8488,N_8520);
nand U9706 (N_9706,N_7835,N_8489);
and U9707 (N_9707,N_7519,N_8287);
nand U9708 (N_9708,N_8516,N_7983);
and U9709 (N_9709,N_7722,N_7946);
or U9710 (N_9710,N_7823,N_7596);
nor U9711 (N_9711,N_8338,N_8594);
or U9712 (N_9712,N_8589,N_8360);
nand U9713 (N_9713,N_7605,N_8596);
nand U9714 (N_9714,N_8680,N_8342);
nor U9715 (N_9715,N_7667,N_8599);
xnor U9716 (N_9716,N_7646,N_8276);
and U9717 (N_9717,N_7898,N_8459);
or U9718 (N_9718,N_7509,N_7906);
xnor U9719 (N_9719,N_7805,N_8403);
xnor U9720 (N_9720,N_8314,N_8261);
or U9721 (N_9721,N_7517,N_8662);
and U9722 (N_9722,N_7770,N_8652);
nor U9723 (N_9723,N_8109,N_7972);
xor U9724 (N_9724,N_8459,N_8665);
or U9725 (N_9725,N_7886,N_7632);
nor U9726 (N_9726,N_8524,N_8071);
xnor U9727 (N_9727,N_8444,N_7681);
nor U9728 (N_9728,N_8090,N_7815);
xnor U9729 (N_9729,N_8060,N_8591);
or U9730 (N_9730,N_7819,N_7809);
and U9731 (N_9731,N_7863,N_7688);
nand U9732 (N_9732,N_8408,N_8288);
nor U9733 (N_9733,N_8144,N_8471);
xor U9734 (N_9734,N_7959,N_7622);
xnor U9735 (N_9735,N_8081,N_7961);
xnor U9736 (N_9736,N_8513,N_8350);
xnor U9737 (N_9737,N_7921,N_7977);
xnor U9738 (N_9738,N_8679,N_8277);
or U9739 (N_9739,N_7826,N_7876);
and U9740 (N_9740,N_7895,N_8519);
nand U9741 (N_9741,N_8719,N_8288);
and U9742 (N_9742,N_8235,N_7566);
nor U9743 (N_9743,N_8191,N_8459);
xnor U9744 (N_9744,N_7803,N_7758);
xor U9745 (N_9745,N_8392,N_7682);
nor U9746 (N_9746,N_8559,N_8336);
xor U9747 (N_9747,N_7755,N_7691);
and U9748 (N_9748,N_7635,N_8468);
or U9749 (N_9749,N_7777,N_7501);
xor U9750 (N_9750,N_7555,N_7923);
or U9751 (N_9751,N_7886,N_7982);
xnor U9752 (N_9752,N_8106,N_8014);
xnor U9753 (N_9753,N_8735,N_8126);
and U9754 (N_9754,N_8040,N_8473);
or U9755 (N_9755,N_7815,N_8039);
nand U9756 (N_9756,N_7655,N_8495);
nor U9757 (N_9757,N_8124,N_7995);
or U9758 (N_9758,N_8140,N_7544);
or U9759 (N_9759,N_8021,N_7581);
nand U9760 (N_9760,N_8201,N_7682);
nand U9761 (N_9761,N_7890,N_8644);
xnor U9762 (N_9762,N_8415,N_7675);
and U9763 (N_9763,N_7676,N_7771);
xor U9764 (N_9764,N_7596,N_7941);
nor U9765 (N_9765,N_7674,N_8689);
and U9766 (N_9766,N_8605,N_8702);
or U9767 (N_9767,N_8227,N_8442);
nand U9768 (N_9768,N_7696,N_7731);
nor U9769 (N_9769,N_7722,N_8370);
xnor U9770 (N_9770,N_7560,N_8214);
or U9771 (N_9771,N_8708,N_8323);
and U9772 (N_9772,N_8302,N_8407);
and U9773 (N_9773,N_7882,N_7893);
and U9774 (N_9774,N_8073,N_8616);
xnor U9775 (N_9775,N_7872,N_8169);
nor U9776 (N_9776,N_8682,N_8305);
xor U9777 (N_9777,N_8189,N_8058);
nand U9778 (N_9778,N_7603,N_8602);
nor U9779 (N_9779,N_8275,N_8522);
or U9780 (N_9780,N_8188,N_7691);
nand U9781 (N_9781,N_8559,N_8010);
nor U9782 (N_9782,N_7799,N_7670);
or U9783 (N_9783,N_8038,N_8508);
and U9784 (N_9784,N_7652,N_7906);
nand U9785 (N_9785,N_8610,N_8571);
xor U9786 (N_9786,N_7934,N_7542);
or U9787 (N_9787,N_7658,N_7689);
xnor U9788 (N_9788,N_8666,N_8561);
and U9789 (N_9789,N_7903,N_8040);
nand U9790 (N_9790,N_8467,N_7958);
nand U9791 (N_9791,N_7728,N_8303);
nor U9792 (N_9792,N_8328,N_8154);
xnor U9793 (N_9793,N_7546,N_8663);
and U9794 (N_9794,N_7638,N_8343);
and U9795 (N_9795,N_7978,N_8324);
and U9796 (N_9796,N_8400,N_8676);
nor U9797 (N_9797,N_8072,N_8466);
nor U9798 (N_9798,N_7728,N_7931);
or U9799 (N_9799,N_8742,N_8124);
xor U9800 (N_9800,N_7921,N_7788);
nand U9801 (N_9801,N_7558,N_8211);
nor U9802 (N_9802,N_7641,N_7628);
xnor U9803 (N_9803,N_7678,N_7712);
and U9804 (N_9804,N_8077,N_8362);
xnor U9805 (N_9805,N_8224,N_7670);
nand U9806 (N_9806,N_8618,N_8072);
nand U9807 (N_9807,N_8091,N_7763);
nor U9808 (N_9808,N_8567,N_8622);
and U9809 (N_9809,N_8633,N_8412);
xnor U9810 (N_9810,N_8281,N_7516);
and U9811 (N_9811,N_8257,N_8588);
nand U9812 (N_9812,N_8060,N_8394);
nand U9813 (N_9813,N_8149,N_7973);
and U9814 (N_9814,N_8399,N_7796);
or U9815 (N_9815,N_7859,N_7860);
or U9816 (N_9816,N_8175,N_8553);
nand U9817 (N_9817,N_8535,N_8521);
and U9818 (N_9818,N_8059,N_7989);
nor U9819 (N_9819,N_8489,N_8743);
nor U9820 (N_9820,N_8242,N_8669);
xor U9821 (N_9821,N_8700,N_8126);
xnor U9822 (N_9822,N_8743,N_8571);
xor U9823 (N_9823,N_8075,N_7736);
xnor U9824 (N_9824,N_8055,N_7502);
nor U9825 (N_9825,N_8220,N_8577);
nand U9826 (N_9826,N_8144,N_8110);
nor U9827 (N_9827,N_8187,N_8349);
nor U9828 (N_9828,N_8702,N_8047);
nand U9829 (N_9829,N_7661,N_8094);
xnor U9830 (N_9830,N_7897,N_7505);
or U9831 (N_9831,N_8452,N_8130);
nand U9832 (N_9832,N_8498,N_8302);
or U9833 (N_9833,N_7622,N_7844);
or U9834 (N_9834,N_8654,N_8660);
nor U9835 (N_9835,N_8342,N_8106);
xor U9836 (N_9836,N_8301,N_8288);
xor U9837 (N_9837,N_7648,N_8273);
and U9838 (N_9838,N_8731,N_8006);
and U9839 (N_9839,N_8154,N_8011);
and U9840 (N_9840,N_8703,N_8574);
nor U9841 (N_9841,N_7574,N_8531);
or U9842 (N_9842,N_8307,N_8197);
and U9843 (N_9843,N_8159,N_7997);
xnor U9844 (N_9844,N_7726,N_7689);
nand U9845 (N_9845,N_7674,N_8222);
xnor U9846 (N_9846,N_8044,N_7505);
nor U9847 (N_9847,N_8507,N_7719);
nand U9848 (N_9848,N_7983,N_8584);
or U9849 (N_9849,N_7772,N_7502);
xnor U9850 (N_9850,N_8639,N_8014);
or U9851 (N_9851,N_8054,N_8374);
or U9852 (N_9852,N_8315,N_8580);
nand U9853 (N_9853,N_8610,N_7699);
xnor U9854 (N_9854,N_7671,N_7912);
and U9855 (N_9855,N_8333,N_7567);
nand U9856 (N_9856,N_8043,N_8537);
nor U9857 (N_9857,N_8623,N_7861);
or U9858 (N_9858,N_7600,N_7958);
and U9859 (N_9859,N_8420,N_8655);
and U9860 (N_9860,N_8717,N_8702);
and U9861 (N_9861,N_8193,N_8145);
nand U9862 (N_9862,N_8430,N_8606);
nor U9863 (N_9863,N_8054,N_8151);
nor U9864 (N_9864,N_7685,N_8714);
xnor U9865 (N_9865,N_8582,N_7507);
xnor U9866 (N_9866,N_7888,N_7967);
nand U9867 (N_9867,N_8056,N_8371);
or U9868 (N_9868,N_7880,N_8057);
nand U9869 (N_9869,N_7975,N_8706);
nor U9870 (N_9870,N_8404,N_8541);
xnor U9871 (N_9871,N_8070,N_8151);
nand U9872 (N_9872,N_8423,N_7863);
nor U9873 (N_9873,N_8128,N_8351);
and U9874 (N_9874,N_8649,N_8729);
and U9875 (N_9875,N_8533,N_8205);
or U9876 (N_9876,N_7784,N_7802);
nand U9877 (N_9877,N_8638,N_8314);
nand U9878 (N_9878,N_8281,N_7517);
nor U9879 (N_9879,N_7916,N_8449);
or U9880 (N_9880,N_7931,N_7872);
nor U9881 (N_9881,N_8402,N_8191);
and U9882 (N_9882,N_7961,N_8029);
nand U9883 (N_9883,N_7742,N_8508);
and U9884 (N_9884,N_8255,N_8413);
nand U9885 (N_9885,N_7871,N_8493);
or U9886 (N_9886,N_8379,N_8647);
xnor U9887 (N_9887,N_8515,N_7670);
nand U9888 (N_9888,N_7735,N_8500);
nor U9889 (N_9889,N_8075,N_8321);
or U9890 (N_9890,N_8318,N_8720);
or U9891 (N_9891,N_7873,N_8720);
and U9892 (N_9892,N_7823,N_7697);
or U9893 (N_9893,N_8636,N_7692);
nand U9894 (N_9894,N_7791,N_7746);
nand U9895 (N_9895,N_8702,N_8148);
and U9896 (N_9896,N_8285,N_7568);
nor U9897 (N_9897,N_7593,N_8640);
nand U9898 (N_9898,N_7561,N_8639);
nand U9899 (N_9899,N_8477,N_8020);
nand U9900 (N_9900,N_7531,N_7951);
and U9901 (N_9901,N_8169,N_7817);
nand U9902 (N_9902,N_7907,N_8431);
and U9903 (N_9903,N_8037,N_7835);
xor U9904 (N_9904,N_8551,N_7508);
nor U9905 (N_9905,N_7694,N_8189);
or U9906 (N_9906,N_8692,N_7559);
and U9907 (N_9907,N_7700,N_7751);
nor U9908 (N_9908,N_8329,N_7782);
nor U9909 (N_9909,N_7562,N_8200);
nand U9910 (N_9910,N_7889,N_8349);
nand U9911 (N_9911,N_7645,N_8418);
and U9912 (N_9912,N_7754,N_7605);
xnor U9913 (N_9913,N_8326,N_7628);
and U9914 (N_9914,N_8184,N_8581);
xor U9915 (N_9915,N_7873,N_7744);
or U9916 (N_9916,N_8510,N_7762);
xnor U9917 (N_9917,N_7991,N_7977);
or U9918 (N_9918,N_8394,N_8118);
xor U9919 (N_9919,N_8028,N_7873);
nand U9920 (N_9920,N_7673,N_8272);
and U9921 (N_9921,N_8221,N_8514);
xor U9922 (N_9922,N_7866,N_7732);
nor U9923 (N_9923,N_8679,N_8092);
and U9924 (N_9924,N_7986,N_8347);
nor U9925 (N_9925,N_8629,N_8567);
nor U9926 (N_9926,N_8342,N_8201);
and U9927 (N_9927,N_8397,N_8352);
or U9928 (N_9928,N_8422,N_8598);
nor U9929 (N_9929,N_8371,N_8197);
xnor U9930 (N_9930,N_8511,N_8442);
nand U9931 (N_9931,N_8384,N_7933);
nand U9932 (N_9932,N_8257,N_8576);
xnor U9933 (N_9933,N_8424,N_8434);
and U9934 (N_9934,N_8536,N_8349);
nor U9935 (N_9935,N_7636,N_7512);
nor U9936 (N_9936,N_7849,N_7772);
nor U9937 (N_9937,N_8413,N_8306);
and U9938 (N_9938,N_7986,N_8693);
xnor U9939 (N_9939,N_8078,N_8329);
xor U9940 (N_9940,N_8217,N_8282);
nor U9941 (N_9941,N_8053,N_8444);
and U9942 (N_9942,N_8308,N_8339);
and U9943 (N_9943,N_7863,N_8319);
nand U9944 (N_9944,N_8549,N_8351);
nor U9945 (N_9945,N_8054,N_8511);
or U9946 (N_9946,N_8712,N_8394);
and U9947 (N_9947,N_8385,N_7868);
or U9948 (N_9948,N_8366,N_7666);
and U9949 (N_9949,N_8399,N_8285);
and U9950 (N_9950,N_7715,N_8309);
xor U9951 (N_9951,N_8150,N_7891);
and U9952 (N_9952,N_8625,N_8154);
xor U9953 (N_9953,N_8640,N_7937);
and U9954 (N_9954,N_7794,N_8075);
and U9955 (N_9955,N_8264,N_7690);
xnor U9956 (N_9956,N_8135,N_8079);
and U9957 (N_9957,N_8217,N_8505);
nand U9958 (N_9958,N_8155,N_8427);
and U9959 (N_9959,N_8582,N_7924);
and U9960 (N_9960,N_7947,N_7787);
nand U9961 (N_9961,N_8165,N_8331);
nand U9962 (N_9962,N_7566,N_8322);
and U9963 (N_9963,N_8644,N_7565);
and U9964 (N_9964,N_8588,N_8017);
or U9965 (N_9965,N_7917,N_8460);
nor U9966 (N_9966,N_8669,N_7846);
nor U9967 (N_9967,N_7935,N_7588);
or U9968 (N_9968,N_8027,N_8714);
and U9969 (N_9969,N_7604,N_8442);
nor U9970 (N_9970,N_7554,N_7658);
and U9971 (N_9971,N_8583,N_7838);
xor U9972 (N_9972,N_8227,N_8378);
nand U9973 (N_9973,N_8375,N_8448);
nor U9974 (N_9974,N_8554,N_8732);
nor U9975 (N_9975,N_8271,N_8455);
nor U9976 (N_9976,N_7914,N_8285);
xor U9977 (N_9977,N_7972,N_7669);
nand U9978 (N_9978,N_7763,N_8114);
and U9979 (N_9979,N_8251,N_7651);
nor U9980 (N_9980,N_8409,N_7728);
and U9981 (N_9981,N_7692,N_8545);
nor U9982 (N_9982,N_8149,N_7922);
nand U9983 (N_9983,N_7784,N_8061);
nor U9984 (N_9984,N_8556,N_7705);
and U9985 (N_9985,N_8723,N_7932);
and U9986 (N_9986,N_7534,N_8173);
xnor U9987 (N_9987,N_7541,N_7501);
or U9988 (N_9988,N_8436,N_7565);
or U9989 (N_9989,N_8494,N_7753);
xor U9990 (N_9990,N_8011,N_8495);
nor U9991 (N_9991,N_8091,N_8673);
or U9992 (N_9992,N_7556,N_8678);
nor U9993 (N_9993,N_7882,N_7950);
xnor U9994 (N_9994,N_8741,N_8012);
xnor U9995 (N_9995,N_8140,N_7947);
or U9996 (N_9996,N_8144,N_8127);
xnor U9997 (N_9997,N_7501,N_7847);
nor U9998 (N_9998,N_8584,N_7661);
or U9999 (N_9999,N_8664,N_8431);
or U10000 (N_10000,N_9022,N_9782);
nor U10001 (N_10001,N_9273,N_9874);
xor U10002 (N_10002,N_9404,N_9472);
nand U10003 (N_10003,N_8980,N_8789);
and U10004 (N_10004,N_8797,N_9465);
xor U10005 (N_10005,N_9771,N_9192);
or U10006 (N_10006,N_9652,N_9187);
nand U10007 (N_10007,N_9118,N_9966);
or U10008 (N_10008,N_9438,N_8810);
xor U10009 (N_10009,N_9708,N_9279);
nand U10010 (N_10010,N_9325,N_9509);
and U10011 (N_10011,N_8884,N_9016);
or U10012 (N_10012,N_9295,N_9674);
or U10013 (N_10013,N_9568,N_9069);
or U10014 (N_10014,N_9625,N_9834);
and U10015 (N_10015,N_9921,N_9470);
and U10016 (N_10016,N_9504,N_9848);
and U10017 (N_10017,N_9035,N_9501);
or U10018 (N_10018,N_8967,N_9157);
or U10019 (N_10019,N_9887,N_9326);
or U10020 (N_10020,N_9508,N_9707);
or U10021 (N_10021,N_9505,N_9493);
or U10022 (N_10022,N_9705,N_9012);
nand U10023 (N_10023,N_9955,N_9398);
and U10024 (N_10024,N_9116,N_9685);
xor U10025 (N_10025,N_9025,N_9245);
nand U10026 (N_10026,N_9930,N_8928);
and U10027 (N_10027,N_8948,N_9130);
nor U10028 (N_10028,N_8925,N_9695);
nor U10029 (N_10029,N_9626,N_9000);
nor U10030 (N_10030,N_9306,N_9056);
xnor U10031 (N_10031,N_9871,N_9667);
xor U10032 (N_10032,N_8772,N_9064);
or U10033 (N_10033,N_9052,N_9147);
nand U10034 (N_10034,N_8907,N_9765);
nand U10035 (N_10035,N_8920,N_9738);
nor U10036 (N_10036,N_8971,N_9275);
or U10037 (N_10037,N_9133,N_9971);
or U10038 (N_10038,N_8777,N_9589);
or U10039 (N_10039,N_9820,N_9546);
nand U10040 (N_10040,N_9244,N_8996);
xnor U10041 (N_10041,N_9110,N_8995);
or U10042 (N_10042,N_9432,N_9431);
xor U10043 (N_10043,N_9555,N_9489);
and U10044 (N_10044,N_9268,N_9906);
or U10045 (N_10045,N_9922,N_9382);
xnor U10046 (N_10046,N_9554,N_9974);
nand U10047 (N_10047,N_9895,N_9490);
or U10048 (N_10048,N_9635,N_9843);
xor U10049 (N_10049,N_9932,N_9796);
nand U10050 (N_10050,N_9624,N_9338);
or U10051 (N_10051,N_9390,N_9261);
and U10052 (N_10052,N_9727,N_9752);
nor U10053 (N_10053,N_9359,N_9204);
or U10054 (N_10054,N_9480,N_9762);
and U10055 (N_10055,N_9567,N_9371);
or U10056 (N_10056,N_9137,N_9145);
nand U10057 (N_10057,N_8774,N_9754);
xor U10058 (N_10058,N_9597,N_8950);
xor U10059 (N_10059,N_9737,N_8816);
and U10060 (N_10060,N_9867,N_9180);
xor U10061 (N_10061,N_9141,N_9474);
nand U10062 (N_10062,N_9368,N_9911);
or U10063 (N_10063,N_9299,N_9928);
or U10064 (N_10064,N_9592,N_9585);
and U10065 (N_10065,N_9986,N_9476);
or U10066 (N_10066,N_9100,N_9503);
and U10067 (N_10067,N_9030,N_9026);
xnor U10068 (N_10068,N_8973,N_9529);
and U10069 (N_10069,N_9174,N_9783);
nand U10070 (N_10070,N_9557,N_9460);
nor U10071 (N_10071,N_9002,N_9491);
or U10072 (N_10072,N_9082,N_9229);
nor U10073 (N_10073,N_9677,N_9679);
or U10074 (N_10074,N_9896,N_8773);
and U10075 (N_10075,N_9015,N_9029);
and U10076 (N_10076,N_8918,N_9436);
or U10077 (N_10077,N_9463,N_9916);
nand U10078 (N_10078,N_9167,N_9537);
nor U10079 (N_10079,N_8750,N_9191);
xnor U10080 (N_10080,N_9775,N_9709);
xor U10081 (N_10081,N_8921,N_9316);
nor U10082 (N_10082,N_9412,N_9233);
nor U10083 (N_10083,N_9282,N_9722);
xor U10084 (N_10084,N_8759,N_9383);
nand U10085 (N_10085,N_9927,N_9055);
or U10086 (N_10086,N_9880,N_9841);
nor U10087 (N_10087,N_9477,N_9328);
nand U10088 (N_10088,N_8753,N_8901);
nor U10089 (N_10089,N_8868,N_9162);
and U10090 (N_10090,N_9059,N_9214);
nand U10091 (N_10091,N_9993,N_9254);
nand U10092 (N_10092,N_9071,N_9632);
nand U10093 (N_10093,N_9252,N_9348);
xnor U10094 (N_10094,N_9816,N_8775);
nand U10095 (N_10095,N_9031,N_9584);
xnor U10096 (N_10096,N_9269,N_9250);
nand U10097 (N_10097,N_8941,N_9962);
or U10098 (N_10098,N_9826,N_9005);
xnor U10099 (N_10099,N_8904,N_9530);
nor U10100 (N_10100,N_9890,N_9621);
and U10101 (N_10101,N_9561,N_9628);
or U10102 (N_10102,N_9441,N_9303);
nand U10103 (N_10103,N_9660,N_9851);
and U10104 (N_10104,N_9821,N_9779);
nor U10105 (N_10105,N_9217,N_9290);
nor U10106 (N_10106,N_9076,N_9200);
nor U10107 (N_10107,N_9964,N_9284);
nor U10108 (N_10108,N_9414,N_9640);
and U10109 (N_10109,N_9413,N_9336);
nand U10110 (N_10110,N_9040,N_9912);
nor U10111 (N_10111,N_9987,N_9690);
xor U10112 (N_10112,N_8978,N_9602);
nand U10113 (N_10113,N_9433,N_9237);
xnor U10114 (N_10114,N_9149,N_9459);
nor U10115 (N_10115,N_9196,N_8761);
or U10116 (N_10116,N_8998,N_9540);
nor U10117 (N_10117,N_9324,N_8910);
nor U10118 (N_10118,N_9104,N_8785);
nor U10119 (N_10119,N_9623,N_8795);
or U10120 (N_10120,N_9395,N_9999);
and U10121 (N_10121,N_8871,N_9772);
or U10122 (N_10122,N_9142,N_9278);
and U10123 (N_10123,N_9136,N_9760);
or U10124 (N_10124,N_9406,N_9291);
nor U10125 (N_10125,N_8878,N_9298);
xor U10126 (N_10126,N_9017,N_9447);
xor U10127 (N_10127,N_9609,N_9789);
nand U10128 (N_10128,N_8791,N_9270);
and U10129 (N_10129,N_8991,N_9337);
or U10130 (N_10130,N_9037,N_9393);
and U10131 (N_10131,N_9692,N_9044);
or U10132 (N_10132,N_8887,N_9315);
and U10133 (N_10133,N_9575,N_9122);
nor U10134 (N_10134,N_9213,N_9716);
xor U10135 (N_10135,N_9092,N_9862);
or U10136 (N_10136,N_8826,N_9161);
xnor U10137 (N_10137,N_9488,N_9595);
and U10138 (N_10138,N_9688,N_9146);
nor U10139 (N_10139,N_9185,N_9656);
or U10140 (N_10140,N_9812,N_9058);
and U10141 (N_10141,N_9758,N_9662);
nor U10142 (N_10142,N_9645,N_9668);
or U10143 (N_10143,N_9558,N_9687);
and U10144 (N_10144,N_8760,N_9155);
or U10145 (N_10145,N_9255,N_9605);
xnor U10146 (N_10146,N_9564,N_9319);
nand U10147 (N_10147,N_9497,N_9903);
xor U10148 (N_10148,N_9531,N_9225);
nor U10149 (N_10149,N_9067,N_9397);
xor U10150 (N_10150,N_9791,N_9089);
nand U10151 (N_10151,N_9389,N_9551);
nand U10152 (N_10152,N_9202,N_8807);
or U10153 (N_10153,N_9691,N_9926);
and U10154 (N_10154,N_9952,N_9954);
and U10155 (N_10155,N_9020,N_9234);
nand U10156 (N_10156,N_9362,N_9860);
or U10157 (N_10157,N_9096,N_9774);
nand U10158 (N_10158,N_9836,N_8831);
nor U10159 (N_10159,N_9288,N_8969);
nand U10160 (N_10160,N_8906,N_9574);
nor U10161 (N_10161,N_8911,N_9377);
xnor U10162 (N_10162,N_9182,N_8849);
nand U10163 (N_10163,N_9838,N_9419);
and U10164 (N_10164,N_9394,N_9941);
nand U10165 (N_10165,N_9188,N_9294);
nand U10166 (N_10166,N_9201,N_9094);
and U10167 (N_10167,N_8752,N_9620);
nand U10168 (N_10168,N_9405,N_9088);
xor U10169 (N_10169,N_9572,N_8850);
nand U10170 (N_10170,N_9437,N_8877);
and U10171 (N_10171,N_8992,N_9651);
nor U10172 (N_10172,N_9550,N_9773);
and U10173 (N_10173,N_9259,N_9753);
or U10174 (N_10174,N_9346,N_9658);
nor U10175 (N_10175,N_9160,N_9098);
or U10176 (N_10176,N_9251,N_9844);
and U10177 (N_10177,N_9197,N_9481);
or U10178 (N_10178,N_9998,N_8963);
nor U10179 (N_10179,N_9205,N_9942);
and U10180 (N_10180,N_9420,N_9333);
nor U10181 (N_10181,N_8840,N_9190);
xnor U10182 (N_10182,N_9144,N_9973);
and U10183 (N_10183,N_9165,N_9611);
nor U10184 (N_10184,N_8860,N_9776);
or U10185 (N_10185,N_9430,N_8890);
and U10186 (N_10186,N_9947,N_8885);
xor U10187 (N_10187,N_8879,N_9833);
and U10188 (N_10188,N_9724,N_9653);
nor U10189 (N_10189,N_9073,N_9714);
and U10190 (N_10190,N_9126,N_9879);
nor U10191 (N_10191,N_9793,N_9473);
nand U10192 (N_10192,N_8873,N_8851);
nand U10193 (N_10193,N_9853,N_9164);
or U10194 (N_10194,N_9949,N_9455);
nand U10195 (N_10195,N_9766,N_9740);
nor U10196 (N_10196,N_8766,N_9266);
nand U10197 (N_10197,N_9664,N_9899);
or U10198 (N_10198,N_9107,N_9027);
nor U10199 (N_10199,N_9021,N_9230);
nor U10200 (N_10200,N_9258,N_9479);
nor U10201 (N_10201,N_9682,N_9385);
nand U10202 (N_10202,N_9819,N_8899);
or U10203 (N_10203,N_9238,N_9934);
xnor U10204 (N_10204,N_8857,N_9427);
or U10205 (N_10205,N_8839,N_9428);
xnor U10206 (N_10206,N_9041,N_9384);
nand U10207 (N_10207,N_9686,N_9112);
or U10208 (N_10208,N_9070,N_9006);
nand U10209 (N_10209,N_9720,N_9053);
nand U10210 (N_10210,N_9840,N_9829);
and U10211 (N_10211,N_8837,N_9910);
and U10212 (N_10212,N_8786,N_9003);
and U10213 (N_10213,N_8997,N_9777);
or U10214 (N_10214,N_8856,N_8943);
xnor U10215 (N_10215,N_9042,N_9885);
xnor U10216 (N_10216,N_8834,N_9905);
nor U10217 (N_10217,N_9957,N_9097);
xor U10218 (N_10218,N_9093,N_8841);
xor U10219 (N_10219,N_8864,N_9054);
nand U10220 (N_10220,N_9543,N_8821);
and U10221 (N_10221,N_9613,N_8932);
xnor U10222 (N_10222,N_9322,N_9757);
or U10223 (N_10223,N_9102,N_9271);
or U10224 (N_10224,N_9293,N_8970);
xnor U10225 (N_10225,N_8993,N_9712);
nand U10226 (N_10226,N_8889,N_9370);
or U10227 (N_10227,N_9454,N_8802);
nor U10228 (N_10228,N_9131,N_9415);
or U10229 (N_10229,N_9570,N_8838);
xor U10230 (N_10230,N_9235,N_9571);
and U10231 (N_10231,N_9696,N_9748);
nor U10232 (N_10232,N_9719,N_9228);
xnor U10233 (N_10233,N_9732,N_9216);
xnor U10234 (N_10234,N_8828,N_9803);
and U10235 (N_10235,N_9539,N_9123);
xor U10236 (N_10236,N_9081,N_9704);
xor U10237 (N_10237,N_9726,N_8765);
and U10238 (N_10238,N_9068,N_9634);
and U10239 (N_10239,N_8751,N_8869);
or U10240 (N_10240,N_9482,N_9600);
nand U10241 (N_10241,N_9004,N_9372);
nand U10242 (N_10242,N_9787,N_9523);
nand U10243 (N_10243,N_9637,N_9618);
and U10244 (N_10244,N_8900,N_9517);
or U10245 (N_10245,N_8763,N_9979);
and U10246 (N_10246,N_9960,N_9553);
nor U10247 (N_10247,N_9387,N_8846);
and U10248 (N_10248,N_9953,N_8961);
xor U10249 (N_10249,N_9061,N_8917);
or U10250 (N_10250,N_9639,N_9893);
or U10251 (N_10251,N_9670,N_8852);
and U10252 (N_10252,N_9334,N_9591);
nand U10253 (N_10253,N_9521,N_9421);
xor U10254 (N_10254,N_9109,N_9761);
or U10255 (N_10255,N_9730,N_9357);
or U10256 (N_10256,N_8939,N_9689);
and U10257 (N_10257,N_9051,N_9728);
nor U10258 (N_10258,N_8931,N_9864);
and U10259 (N_10259,N_8845,N_9556);
nand U10260 (N_10260,N_8796,N_9702);
xor U10261 (N_10261,N_9701,N_9134);
xnor U10262 (N_10262,N_9125,N_9630);
or U10263 (N_10263,N_9379,N_8934);
nand U10264 (N_10264,N_9260,N_8762);
xor U10265 (N_10265,N_8909,N_9845);
or U10266 (N_10266,N_9717,N_9443);
and U10267 (N_10267,N_9499,N_9650);
and U10268 (N_10268,N_9976,N_8800);
or U10269 (N_10269,N_9296,N_8855);
or U10270 (N_10270,N_9552,N_9856);
nand U10271 (N_10271,N_9579,N_8914);
nand U10272 (N_10272,N_9918,N_9992);
or U10273 (N_10273,N_9559,N_8842);
nand U10274 (N_10274,N_9883,N_9411);
and U10275 (N_10275,N_9839,N_9050);
and U10276 (N_10276,N_9289,N_9920);
or U10277 (N_10277,N_9138,N_9799);
or U10278 (N_10278,N_9512,N_9287);
nand U10279 (N_10279,N_9240,N_9150);
and U10280 (N_10280,N_9086,N_9560);
xor U10281 (N_10281,N_9074,N_9814);
nor U10282 (N_10282,N_9364,N_9001);
and U10283 (N_10283,N_9831,N_8905);
and U10284 (N_10284,N_9329,N_9809);
nor U10285 (N_10285,N_9938,N_8985);
nand U10286 (N_10286,N_9311,N_9566);
xnor U10287 (N_10287,N_8768,N_9510);
and U10288 (N_10288,N_8764,N_8981);
nor U10289 (N_10289,N_9909,N_9478);
or U10290 (N_10290,N_8875,N_9241);
nand U10291 (N_10291,N_9535,N_9946);
and U10292 (N_10292,N_8972,N_9593);
xnor U10293 (N_10293,N_9739,N_9276);
or U10294 (N_10294,N_9795,N_9314);
nor U10295 (N_10295,N_9967,N_8830);
or U10296 (N_10296,N_9528,N_9274);
and U10297 (N_10297,N_8803,N_8798);
or U10298 (N_10298,N_8960,N_9410);
xor U10299 (N_10299,N_9545,N_9914);
nand U10300 (N_10300,N_8872,N_8792);
xor U10301 (N_10301,N_9358,N_9132);
nand U10302 (N_10302,N_8987,N_9292);
nor U10303 (N_10303,N_9475,N_9894);
or U10304 (N_10304,N_9743,N_9469);
or U10305 (N_10305,N_9457,N_9583);
or U10306 (N_10306,N_9057,N_8937);
or U10307 (N_10307,N_8848,N_9193);
nand U10308 (N_10308,N_8903,N_9548);
nand U10309 (N_10309,N_9657,N_9961);
or U10310 (N_10310,N_9194,N_9735);
xnor U10311 (N_10311,N_9373,N_9633);
nor U10312 (N_10312,N_9907,N_9869);
nand U10313 (N_10313,N_9980,N_9090);
nand U10314 (N_10314,N_9283,N_9310);
nor U10315 (N_10315,N_9863,N_9425);
nand U10316 (N_10316,N_9360,N_9562);
nor U10317 (N_10317,N_9643,N_9256);
xnor U10318 (N_10318,N_9231,N_9868);
nor U10319 (N_10319,N_9784,N_9697);
or U10320 (N_10320,N_9576,N_9152);
and U10321 (N_10321,N_9533,N_8865);
or U10322 (N_10322,N_8801,N_9994);
or U10323 (N_10323,N_8926,N_9801);
xnor U10324 (N_10324,N_9019,N_9669);
and U10325 (N_10325,N_9675,N_9904);
nand U10326 (N_10326,N_8893,N_9788);
xnor U10327 (N_10327,N_9308,N_8949);
and U10328 (N_10328,N_8898,N_9997);
nor U10329 (N_10329,N_9400,N_9342);
or U10330 (N_10330,N_9698,N_9492);
nor U10331 (N_10331,N_9642,N_9417);
nor U10332 (N_10332,N_9084,N_9498);
nor U10333 (N_10333,N_9549,N_9984);
nor U10334 (N_10334,N_9159,N_9802);
and U10335 (N_10335,N_9426,N_8862);
or U10336 (N_10336,N_8896,N_9331);
xor U10337 (N_10337,N_9804,N_8858);
nor U10338 (N_10338,N_9350,N_8958);
nand U10339 (N_10339,N_9378,N_9937);
nor U10340 (N_10340,N_9177,N_9915);
xnor U10341 (N_10341,N_9127,N_9063);
or U10342 (N_10342,N_9872,N_8758);
or U10343 (N_10343,N_8923,N_9111);
or U10344 (N_10344,N_8938,N_9148);
nand U10345 (N_10345,N_9341,N_9990);
xor U10346 (N_10346,N_9487,N_8968);
nor U10347 (N_10347,N_8782,N_9518);
or U10348 (N_10348,N_9563,N_9859);
nor U10349 (N_10349,N_9343,N_9154);
nand U10350 (N_10350,N_9532,N_9542);
or U10351 (N_10351,N_9120,N_8986);
and U10352 (N_10352,N_9424,N_9305);
xnor U10353 (N_10353,N_9538,N_9800);
nor U10354 (N_10354,N_9636,N_9627);
nor U10355 (N_10355,N_9654,N_9199);
xor U10356 (N_10356,N_9889,N_8994);
or U10357 (N_10357,N_8902,N_9221);
xor U10358 (N_10358,N_9684,N_9222);
xnor U10359 (N_10359,N_8799,N_8912);
xnor U10360 (N_10360,N_9596,N_9206);
nand U10361 (N_10361,N_9075,N_9815);
nand U10362 (N_10362,N_9694,N_9855);
or U10363 (N_10363,N_9172,N_9590);
and U10364 (N_10364,N_8976,N_9835);
nor U10365 (N_10365,N_9790,N_9113);
nor U10366 (N_10366,N_9536,N_8990);
nand U10367 (N_10367,N_8975,N_8933);
nor U10368 (N_10368,N_9449,N_9736);
nor U10369 (N_10369,N_9923,N_9401);
nor U10370 (N_10370,N_9302,N_9756);
nand U10371 (N_10371,N_9781,N_9085);
or U10372 (N_10372,N_9304,N_9734);
or U10373 (N_10373,N_9117,N_9313);
nand U10374 (N_10374,N_9768,N_9456);
or U10375 (N_10375,N_8947,N_9332);
nor U10376 (N_10376,N_9817,N_9699);
nor U10377 (N_10377,N_9991,N_9806);
and U10378 (N_10378,N_9666,N_9179);
nor U10379 (N_10379,N_8827,N_9087);
nor U10380 (N_10380,N_9265,N_9467);
or U10381 (N_10381,N_8927,N_9671);
or U10382 (N_10382,N_9983,N_8983);
and U10383 (N_10383,N_8836,N_9515);
nor U10384 (N_10384,N_9908,N_9718);
and U10385 (N_10385,N_9227,N_9981);
or U10386 (N_10386,N_9965,N_9236);
xnor U10387 (N_10387,N_9361,N_9151);
and U10388 (N_10388,N_8853,N_9351);
nor U10389 (N_10389,N_9335,N_9386);
or U10390 (N_10390,N_9919,N_9877);
nand U10391 (N_10391,N_9119,N_8892);
and U10392 (N_10392,N_9825,N_9745);
xnor U10393 (N_10393,N_8757,N_9032);
xnor U10394 (N_10394,N_9036,N_8888);
and U10395 (N_10395,N_8809,N_9106);
nor U10396 (N_10396,N_8814,N_9565);
nand U10397 (N_10397,N_9339,N_9211);
nand U10398 (N_10398,N_9519,N_9729);
nor U10399 (N_10399,N_9830,N_9169);
and U10400 (N_10400,N_9970,N_9077);
nand U10401 (N_10401,N_9285,N_8847);
or U10402 (N_10402,N_9023,N_9622);
or U10403 (N_10403,N_8808,N_9770);
and U10404 (N_10404,N_9948,N_8965);
and U10405 (N_10405,N_8787,N_9913);
or U10406 (N_10406,N_9917,N_9985);
nand U10407 (N_10407,N_9170,N_9494);
or U10408 (N_10408,N_8867,N_9253);
or U10409 (N_10409,N_9847,N_9239);
nand U10410 (N_10410,N_8832,N_9811);
and U10411 (N_10411,N_9587,N_8804);
or U10412 (N_10412,N_8916,N_9468);
nand U10413 (N_10413,N_9604,N_8954);
nor U10414 (N_10414,N_9355,N_9140);
xnor U10415 (N_10415,N_9731,N_9822);
or U10416 (N_10416,N_9659,N_9024);
and U10417 (N_10417,N_9603,N_9577);
and U10418 (N_10418,N_9007,N_9321);
nand U10419 (N_10419,N_8824,N_9631);
and U10420 (N_10420,N_9173,N_9312);
nor U10421 (N_10421,N_9391,N_9764);
and U10422 (N_10422,N_9823,N_9451);
and U10423 (N_10423,N_9612,N_9219);
and U10424 (N_10424,N_9725,N_9380);
and U10425 (N_10425,N_9178,N_8881);
xor U10426 (N_10426,N_9902,N_9354);
nor U10427 (N_10427,N_9416,N_9223);
or U10428 (N_10428,N_9062,N_9786);
or U10429 (N_10429,N_9526,N_9248);
nor U10430 (N_10430,N_9242,N_9011);
nand U10431 (N_10431,N_9045,N_8929);
and U10432 (N_10432,N_9402,N_9892);
nor U10433 (N_10433,N_9649,N_9471);
or U10434 (N_10434,N_8935,N_9832);
nor U10435 (N_10435,N_9828,N_8895);
and U10436 (N_10436,N_9139,N_9710);
and U10437 (N_10437,N_9744,N_9409);
nor U10438 (N_10438,N_9163,N_8882);
or U10439 (N_10439,N_8822,N_9115);
nor U10440 (N_10440,N_9440,N_9524);
xor U10441 (N_10441,N_9267,N_9582);
and U10442 (N_10442,N_8770,N_9263);
nand U10443 (N_10443,N_9369,N_9207);
xnor U10444 (N_10444,N_9580,N_9700);
and U10445 (N_10445,N_9616,N_8999);
nor U10446 (N_10446,N_9135,N_9849);
and U10447 (N_10447,N_9511,N_9143);
nand U10448 (N_10448,N_9224,N_9103);
xnor U10449 (N_10449,N_9547,N_9038);
nand U10450 (N_10450,N_9924,N_9759);
nand U10451 (N_10451,N_8982,N_9422);
and U10452 (N_10452,N_8863,N_9852);
and U10453 (N_10453,N_8955,N_9681);
nor U10454 (N_10454,N_8883,N_9573);
nor U10455 (N_10455,N_9995,N_9721);
xor U10456 (N_10456,N_9065,N_8866);
nor U10457 (N_10457,N_9418,N_9769);
and U10458 (N_10458,N_9663,N_9309);
and U10459 (N_10459,N_9824,N_8819);
nor U10460 (N_10460,N_9763,N_9956);
and U10461 (N_10461,N_8959,N_8966);
xor U10462 (N_10462,N_8818,N_9189);
or U10463 (N_10463,N_9901,N_9317);
nand U10464 (N_10464,N_9318,N_9464);
and U10465 (N_10465,N_8780,N_9349);
nor U10466 (N_10466,N_9099,N_9195);
and U10467 (N_10467,N_9606,N_9988);
nand U10468 (N_10468,N_9982,N_9506);
or U10469 (N_10469,N_9661,N_9969);
nand U10470 (N_10470,N_8859,N_9608);
xnor U10471 (N_10471,N_9996,N_8776);
nand U10472 (N_10472,N_9977,N_9807);
nor U10473 (N_10473,N_9866,N_8876);
or U10474 (N_10474,N_9882,N_9376);
or U10475 (N_10475,N_9792,N_9881);
or U10476 (N_10476,N_8771,N_8813);
nor U10477 (N_10477,N_8915,N_9186);
nor U10478 (N_10478,N_9797,N_9014);
or U10479 (N_10479,N_9365,N_8805);
and U10480 (N_10480,N_9876,N_8940);
or U10481 (N_10481,N_9870,N_9644);
nor U10482 (N_10482,N_9678,N_9300);
nand U10483 (N_10483,N_9598,N_9850);
nand U10484 (N_10484,N_9462,N_9778);
nand U10485 (N_10485,N_8894,N_9461);
or U10486 (N_10486,N_9033,N_9435);
or U10487 (N_10487,N_8769,N_9280);
and U10488 (N_10488,N_9891,N_9034);
nand U10489 (N_10489,N_9344,N_9448);
or U10490 (N_10490,N_9407,N_9446);
xnor U10491 (N_10491,N_9028,N_9522);
and U10492 (N_10492,N_9247,N_8794);
and U10493 (N_10493,N_9780,N_9898);
nor U10494 (N_10494,N_8951,N_9935);
and U10495 (N_10495,N_9226,N_9878);
nor U10496 (N_10496,N_9458,N_9875);
nand U10497 (N_10497,N_9706,N_9330);
or U10498 (N_10498,N_9648,N_9733);
xnor U10499 (N_10499,N_9647,N_8781);
and U10500 (N_10500,N_9171,N_9484);
xor U10501 (N_10501,N_9079,N_8988);
nor U10502 (N_10502,N_9156,N_9466);
xnor U10503 (N_10503,N_8945,N_9495);
nand U10504 (N_10504,N_9813,N_9805);
and U10505 (N_10505,N_9713,N_9184);
xnor U10506 (N_10506,N_9375,N_9158);
nand U10507 (N_10507,N_8829,N_9277);
xor U10508 (N_10508,N_9629,N_9741);
xnor U10509 (N_10509,N_9208,N_9673);
and U10510 (N_10510,N_9683,N_9039);
or U10511 (N_10511,N_9210,N_9352);
nor U10512 (N_10512,N_9272,N_9047);
or U10513 (N_10513,N_8835,N_9742);
and U10514 (N_10514,N_8880,N_9886);
xnor U10515 (N_10515,N_9968,N_8874);
nor U10516 (N_10516,N_9818,N_8844);
nor U10517 (N_10517,N_9243,N_9423);
xor U10518 (N_10518,N_9641,N_9665);
nand U10519 (N_10519,N_9212,N_9249);
xnor U10520 (N_10520,N_9452,N_9588);
and U10521 (N_10521,N_9767,N_9978);
xor U10522 (N_10522,N_8922,N_8952);
and U10523 (N_10523,N_9750,N_9327);
nand U10524 (N_10524,N_9933,N_8891);
nand U10525 (N_10525,N_8754,N_9049);
nor U10526 (N_10526,N_9601,N_9008);
nand U10527 (N_10527,N_8870,N_8979);
xnor U10528 (N_10528,N_9514,N_9453);
nand U10529 (N_10529,N_9963,N_9166);
xor U10530 (N_10530,N_9072,N_9345);
nor U10531 (N_10531,N_8811,N_9366);
or U10532 (N_10532,N_9785,N_9951);
or U10533 (N_10533,N_9183,N_9569);
nor U10534 (N_10534,N_9010,N_9181);
xor U10535 (N_10535,N_9198,N_9507);
and U10536 (N_10536,N_9842,N_9972);
nand U10537 (N_10537,N_9958,N_8962);
nand U10538 (N_10538,N_9450,N_9746);
or U10539 (N_10539,N_9403,N_9486);
xnor U10540 (N_10540,N_9396,N_9578);
or U10541 (N_10541,N_9046,N_9399);
nand U10542 (N_10542,N_9286,N_9827);
nor U10543 (N_10543,N_9900,N_9617);
nor U10544 (N_10544,N_9794,N_8793);
nor U10545 (N_10545,N_9747,N_8755);
nor U10546 (N_10546,N_9363,N_9374);
nand U10547 (N_10547,N_8820,N_9693);
nand U10548 (N_10548,N_9444,N_9124);
nor U10549 (N_10549,N_9091,N_9615);
and U10550 (N_10550,N_9168,N_9516);
xnor U10551 (N_10551,N_9320,N_9755);
or U10552 (N_10552,N_9392,N_9083);
xor U10553 (N_10553,N_9340,N_9837);
or U10554 (N_10554,N_9607,N_9175);
and U10555 (N_10555,N_9865,N_9959);
nand U10556 (N_10556,N_9940,N_9153);
xnor U10557 (N_10557,N_9599,N_9232);
and U10558 (N_10558,N_9215,N_9209);
nand U10559 (N_10559,N_8815,N_9262);
xnor U10560 (N_10560,N_8977,N_9534);
or U10561 (N_10561,N_9105,N_9619);
nand U10562 (N_10562,N_9281,N_9513);
xnor U10563 (N_10563,N_8936,N_9078);
or U10564 (N_10564,N_9703,N_9925);
and U10565 (N_10565,N_8812,N_9945);
nand U10566 (N_10566,N_9060,N_9176);
xnor U10567 (N_10567,N_9808,N_9989);
xnor U10568 (N_10568,N_8817,N_9323);
nor U10569 (N_10569,N_9544,N_9114);
nor U10570 (N_10570,N_9723,N_8778);
or U10571 (N_10571,N_9749,N_9121);
nor U10572 (N_10572,N_9715,N_8784);
xnor U10573 (N_10573,N_9810,N_9586);
or U10574 (N_10574,N_8984,N_8908);
nor U10575 (N_10575,N_8783,N_8779);
xnor U10576 (N_10576,N_8957,N_9939);
nand U10577 (N_10577,N_9931,N_9367);
and U10578 (N_10578,N_9610,N_9520);
nor U10579 (N_10579,N_9246,N_9408);
nor U10580 (N_10580,N_9496,N_8974);
nor U10581 (N_10581,N_8861,N_9798);
or U10582 (N_10582,N_8790,N_8946);
nor U10583 (N_10583,N_9646,N_9858);
xnor U10584 (N_10584,N_9066,N_9381);
nor U10585 (N_10585,N_9936,N_8854);
nor U10586 (N_10586,N_9672,N_8930);
or U10587 (N_10587,N_9264,N_8919);
nand U10588 (N_10588,N_9043,N_9009);
xnor U10589 (N_10589,N_9018,N_9638);
nand U10590 (N_10590,N_9594,N_9080);
or U10591 (N_10591,N_9307,N_8964);
or U10592 (N_10592,N_8756,N_9676);
xor U10593 (N_10593,N_9711,N_9101);
nor U10594 (N_10594,N_8833,N_9485);
nor U10595 (N_10595,N_9944,N_9128);
nor U10596 (N_10596,N_9257,N_8956);
xor U10597 (N_10597,N_9861,N_9439);
and U10598 (N_10598,N_9013,N_9854);
nor U10599 (N_10599,N_8825,N_9525);
nand U10600 (N_10600,N_9888,N_8944);
and U10601 (N_10601,N_9353,N_9751);
and U10602 (N_10602,N_9614,N_9655);
xnor U10603 (N_10603,N_8924,N_9502);
nor U10604 (N_10604,N_9347,N_9943);
or U10605 (N_10605,N_9129,N_9429);
nand U10606 (N_10606,N_8843,N_9884);
xor U10607 (N_10607,N_8953,N_8989);
and U10608 (N_10608,N_9846,N_8942);
nor U10609 (N_10609,N_9108,N_9434);
or U10610 (N_10610,N_9527,N_9929);
and U10611 (N_10611,N_8897,N_8788);
xor U10612 (N_10612,N_8886,N_9388);
or U10613 (N_10613,N_9680,N_9873);
and U10614 (N_10614,N_9095,N_9218);
xnor U10615 (N_10615,N_9445,N_9483);
nor U10616 (N_10616,N_9442,N_9950);
nand U10617 (N_10617,N_9581,N_8767);
or U10618 (N_10618,N_9220,N_9297);
nand U10619 (N_10619,N_8913,N_9897);
nor U10620 (N_10620,N_9857,N_8806);
nor U10621 (N_10621,N_9500,N_9203);
xor U10622 (N_10622,N_8823,N_9301);
and U10623 (N_10623,N_9975,N_9048);
or U10624 (N_10624,N_9356,N_9541);
nor U10625 (N_10625,N_9858,N_8833);
xor U10626 (N_10626,N_8795,N_9686);
xor U10627 (N_10627,N_9234,N_9146);
nor U10628 (N_10628,N_9296,N_9040);
xor U10629 (N_10629,N_9573,N_8839);
nand U10630 (N_10630,N_9485,N_9551);
xnor U10631 (N_10631,N_9475,N_9406);
nor U10632 (N_10632,N_8958,N_9214);
or U10633 (N_10633,N_9326,N_9554);
xnor U10634 (N_10634,N_9584,N_9371);
nand U10635 (N_10635,N_8886,N_9883);
nand U10636 (N_10636,N_9587,N_9040);
xnor U10637 (N_10637,N_9997,N_9677);
nand U10638 (N_10638,N_9892,N_9241);
xnor U10639 (N_10639,N_9306,N_9528);
nand U10640 (N_10640,N_9611,N_9320);
nand U10641 (N_10641,N_8769,N_8794);
xor U10642 (N_10642,N_9827,N_9120);
xnor U10643 (N_10643,N_9670,N_9323);
nor U10644 (N_10644,N_9261,N_9606);
nor U10645 (N_10645,N_9418,N_9523);
or U10646 (N_10646,N_8875,N_9265);
nor U10647 (N_10647,N_9296,N_9906);
nand U10648 (N_10648,N_9656,N_9334);
nand U10649 (N_10649,N_9906,N_9114);
nand U10650 (N_10650,N_8951,N_9580);
nand U10651 (N_10651,N_9012,N_9476);
nor U10652 (N_10652,N_9061,N_9651);
and U10653 (N_10653,N_9614,N_8807);
nand U10654 (N_10654,N_9907,N_9079);
and U10655 (N_10655,N_9317,N_9134);
or U10656 (N_10656,N_9393,N_8907);
nand U10657 (N_10657,N_9277,N_8980);
or U10658 (N_10658,N_9308,N_9632);
nand U10659 (N_10659,N_9886,N_9744);
nand U10660 (N_10660,N_9570,N_8866);
nand U10661 (N_10661,N_9903,N_9588);
nand U10662 (N_10662,N_9066,N_9767);
and U10663 (N_10663,N_9662,N_9005);
or U10664 (N_10664,N_8854,N_9586);
or U10665 (N_10665,N_9437,N_9953);
nor U10666 (N_10666,N_9062,N_9215);
xor U10667 (N_10667,N_9745,N_8995);
nand U10668 (N_10668,N_9897,N_9858);
and U10669 (N_10669,N_9128,N_9504);
xor U10670 (N_10670,N_9414,N_8979);
nand U10671 (N_10671,N_9486,N_9207);
nand U10672 (N_10672,N_9197,N_9203);
or U10673 (N_10673,N_9872,N_9923);
nor U10674 (N_10674,N_9613,N_9993);
xor U10675 (N_10675,N_9720,N_9650);
nand U10676 (N_10676,N_9757,N_8833);
nand U10677 (N_10677,N_9722,N_9122);
nand U10678 (N_10678,N_8777,N_9032);
xor U10679 (N_10679,N_8901,N_9202);
xnor U10680 (N_10680,N_9357,N_9042);
nor U10681 (N_10681,N_9993,N_8922);
xnor U10682 (N_10682,N_9546,N_9922);
nand U10683 (N_10683,N_9178,N_9643);
or U10684 (N_10684,N_8802,N_8899);
xor U10685 (N_10685,N_9082,N_9057);
xor U10686 (N_10686,N_8912,N_9114);
xnor U10687 (N_10687,N_9047,N_9270);
nor U10688 (N_10688,N_9754,N_8928);
nor U10689 (N_10689,N_9186,N_9873);
xor U10690 (N_10690,N_9578,N_9703);
nand U10691 (N_10691,N_9919,N_9633);
nand U10692 (N_10692,N_9751,N_9811);
nor U10693 (N_10693,N_9593,N_9379);
xor U10694 (N_10694,N_8892,N_8852);
and U10695 (N_10695,N_9139,N_9542);
nor U10696 (N_10696,N_8836,N_9079);
or U10697 (N_10697,N_8843,N_9408);
or U10698 (N_10698,N_8753,N_9860);
nand U10699 (N_10699,N_9137,N_9024);
and U10700 (N_10700,N_9691,N_9548);
and U10701 (N_10701,N_9265,N_9964);
and U10702 (N_10702,N_9217,N_9401);
nand U10703 (N_10703,N_9134,N_8810);
and U10704 (N_10704,N_9147,N_9059);
and U10705 (N_10705,N_9884,N_8927);
xor U10706 (N_10706,N_9202,N_9715);
nand U10707 (N_10707,N_8941,N_9170);
xor U10708 (N_10708,N_9607,N_9652);
xnor U10709 (N_10709,N_9971,N_9606);
and U10710 (N_10710,N_8949,N_9872);
nor U10711 (N_10711,N_8763,N_8901);
nand U10712 (N_10712,N_9574,N_9576);
nor U10713 (N_10713,N_9513,N_8827);
nor U10714 (N_10714,N_9944,N_9264);
and U10715 (N_10715,N_9371,N_8949);
or U10716 (N_10716,N_9228,N_8806);
nor U10717 (N_10717,N_9184,N_9182);
nor U10718 (N_10718,N_9032,N_9375);
or U10719 (N_10719,N_9204,N_9449);
nand U10720 (N_10720,N_9087,N_9432);
nor U10721 (N_10721,N_9167,N_9000);
and U10722 (N_10722,N_8822,N_9501);
and U10723 (N_10723,N_9174,N_8859);
xor U10724 (N_10724,N_9852,N_8770);
xor U10725 (N_10725,N_9043,N_9732);
or U10726 (N_10726,N_9102,N_8764);
or U10727 (N_10727,N_9054,N_8812);
or U10728 (N_10728,N_8863,N_8949);
nor U10729 (N_10729,N_9043,N_8799);
and U10730 (N_10730,N_9684,N_9045);
or U10731 (N_10731,N_9716,N_9802);
or U10732 (N_10732,N_9455,N_9622);
nor U10733 (N_10733,N_9776,N_9264);
nor U10734 (N_10734,N_8791,N_9874);
nor U10735 (N_10735,N_9149,N_9833);
nor U10736 (N_10736,N_9840,N_8801);
and U10737 (N_10737,N_9740,N_9419);
nor U10738 (N_10738,N_9788,N_9389);
and U10739 (N_10739,N_8815,N_8987);
and U10740 (N_10740,N_9990,N_9545);
or U10741 (N_10741,N_8925,N_9258);
xnor U10742 (N_10742,N_8903,N_9121);
nor U10743 (N_10743,N_9806,N_9689);
nor U10744 (N_10744,N_8833,N_9709);
xor U10745 (N_10745,N_9711,N_9182);
and U10746 (N_10746,N_9198,N_9121);
and U10747 (N_10747,N_8860,N_9633);
or U10748 (N_10748,N_9308,N_9577);
nor U10749 (N_10749,N_9096,N_9898);
and U10750 (N_10750,N_9355,N_9481);
xnor U10751 (N_10751,N_9095,N_9625);
xor U10752 (N_10752,N_9496,N_9317);
or U10753 (N_10753,N_9141,N_9274);
or U10754 (N_10754,N_9558,N_9622);
xnor U10755 (N_10755,N_8805,N_9179);
and U10756 (N_10756,N_9583,N_9953);
nand U10757 (N_10757,N_9098,N_9520);
nand U10758 (N_10758,N_8843,N_9534);
xnor U10759 (N_10759,N_9251,N_8815);
or U10760 (N_10760,N_8907,N_9873);
nor U10761 (N_10761,N_9321,N_9479);
nor U10762 (N_10762,N_9349,N_9541);
nor U10763 (N_10763,N_8916,N_9697);
xnor U10764 (N_10764,N_9849,N_9994);
or U10765 (N_10765,N_8975,N_9228);
or U10766 (N_10766,N_9383,N_9581);
and U10767 (N_10767,N_9615,N_9587);
xnor U10768 (N_10768,N_9810,N_8838);
nand U10769 (N_10769,N_9613,N_9932);
and U10770 (N_10770,N_9361,N_9772);
and U10771 (N_10771,N_9296,N_8841);
xor U10772 (N_10772,N_8938,N_9303);
and U10773 (N_10773,N_8764,N_9809);
nor U10774 (N_10774,N_9738,N_8809);
nand U10775 (N_10775,N_9227,N_8920);
nand U10776 (N_10776,N_9206,N_9387);
nand U10777 (N_10777,N_9527,N_9127);
nand U10778 (N_10778,N_9459,N_8837);
nand U10779 (N_10779,N_9607,N_8766);
nand U10780 (N_10780,N_9923,N_9595);
nor U10781 (N_10781,N_9245,N_9428);
nor U10782 (N_10782,N_9977,N_9623);
nand U10783 (N_10783,N_9184,N_8868);
nand U10784 (N_10784,N_9052,N_9458);
nor U10785 (N_10785,N_9740,N_9729);
nor U10786 (N_10786,N_9649,N_9129);
xor U10787 (N_10787,N_8995,N_8897);
nor U10788 (N_10788,N_9146,N_9509);
and U10789 (N_10789,N_8997,N_9574);
nor U10790 (N_10790,N_9587,N_9196);
and U10791 (N_10791,N_9438,N_9488);
or U10792 (N_10792,N_9536,N_9097);
nand U10793 (N_10793,N_9778,N_9544);
nor U10794 (N_10794,N_9699,N_9499);
xor U10795 (N_10795,N_9758,N_9208);
or U10796 (N_10796,N_9960,N_9285);
xor U10797 (N_10797,N_8809,N_9287);
and U10798 (N_10798,N_8974,N_8755);
nor U10799 (N_10799,N_9425,N_9381);
and U10800 (N_10800,N_9552,N_9782);
and U10801 (N_10801,N_9397,N_9707);
and U10802 (N_10802,N_9688,N_9826);
xnor U10803 (N_10803,N_9393,N_9771);
xor U10804 (N_10804,N_9447,N_8988);
nand U10805 (N_10805,N_9105,N_9807);
xnor U10806 (N_10806,N_9399,N_9127);
nand U10807 (N_10807,N_8864,N_9324);
or U10808 (N_10808,N_9054,N_9277);
and U10809 (N_10809,N_9819,N_9569);
nand U10810 (N_10810,N_8752,N_9334);
nor U10811 (N_10811,N_9142,N_8862);
nor U10812 (N_10812,N_9765,N_8928);
nor U10813 (N_10813,N_9365,N_8775);
nor U10814 (N_10814,N_9350,N_9938);
xnor U10815 (N_10815,N_8915,N_9869);
or U10816 (N_10816,N_9445,N_9008);
nor U10817 (N_10817,N_9772,N_8947);
nor U10818 (N_10818,N_9990,N_9221);
nand U10819 (N_10819,N_9743,N_9070);
and U10820 (N_10820,N_9319,N_9475);
nor U10821 (N_10821,N_8904,N_8873);
or U10822 (N_10822,N_9608,N_9588);
or U10823 (N_10823,N_9128,N_9998);
and U10824 (N_10824,N_8843,N_9906);
nor U10825 (N_10825,N_9629,N_9140);
xnor U10826 (N_10826,N_9069,N_9864);
or U10827 (N_10827,N_9823,N_8860);
or U10828 (N_10828,N_9689,N_9767);
nand U10829 (N_10829,N_9966,N_9804);
xor U10830 (N_10830,N_8871,N_9626);
nand U10831 (N_10831,N_9665,N_9860);
and U10832 (N_10832,N_9226,N_9575);
and U10833 (N_10833,N_9240,N_9861);
or U10834 (N_10834,N_8909,N_8755);
and U10835 (N_10835,N_9141,N_9723);
and U10836 (N_10836,N_9201,N_9818);
nand U10837 (N_10837,N_8969,N_9446);
and U10838 (N_10838,N_9919,N_9842);
nand U10839 (N_10839,N_9009,N_9456);
nand U10840 (N_10840,N_9560,N_9966);
nand U10841 (N_10841,N_9048,N_9317);
and U10842 (N_10842,N_8988,N_9220);
xnor U10843 (N_10843,N_9793,N_9567);
xor U10844 (N_10844,N_9933,N_9920);
nand U10845 (N_10845,N_9654,N_9364);
xor U10846 (N_10846,N_9186,N_9620);
nand U10847 (N_10847,N_8887,N_9566);
nor U10848 (N_10848,N_9263,N_9724);
and U10849 (N_10849,N_9253,N_8835);
nand U10850 (N_10850,N_9618,N_9458);
and U10851 (N_10851,N_9691,N_9851);
and U10852 (N_10852,N_9225,N_9128);
and U10853 (N_10853,N_9935,N_8905);
and U10854 (N_10854,N_9779,N_8751);
or U10855 (N_10855,N_9138,N_9362);
or U10856 (N_10856,N_9168,N_9145);
xor U10857 (N_10857,N_9414,N_8953);
and U10858 (N_10858,N_9721,N_9179);
xor U10859 (N_10859,N_8803,N_8818);
nand U10860 (N_10860,N_8893,N_9110);
or U10861 (N_10861,N_9302,N_9202);
and U10862 (N_10862,N_9834,N_9438);
xor U10863 (N_10863,N_9304,N_8843);
xor U10864 (N_10864,N_9551,N_9623);
nand U10865 (N_10865,N_8881,N_8914);
and U10866 (N_10866,N_9000,N_9772);
nor U10867 (N_10867,N_8763,N_9895);
nand U10868 (N_10868,N_9367,N_9504);
nor U10869 (N_10869,N_9114,N_9158);
xor U10870 (N_10870,N_9052,N_9840);
nand U10871 (N_10871,N_9306,N_9059);
and U10872 (N_10872,N_9348,N_8865);
nand U10873 (N_10873,N_9059,N_9846);
nor U10874 (N_10874,N_9761,N_9736);
nor U10875 (N_10875,N_9724,N_9166);
nand U10876 (N_10876,N_8918,N_9663);
nor U10877 (N_10877,N_9683,N_9249);
nand U10878 (N_10878,N_8906,N_9805);
and U10879 (N_10879,N_9060,N_8939);
nand U10880 (N_10880,N_9040,N_8822);
nor U10881 (N_10881,N_8920,N_8949);
nand U10882 (N_10882,N_9735,N_8964);
or U10883 (N_10883,N_9639,N_8837);
nor U10884 (N_10884,N_9181,N_9449);
nor U10885 (N_10885,N_9114,N_9852);
nand U10886 (N_10886,N_8894,N_9675);
xnor U10887 (N_10887,N_9085,N_9091);
nand U10888 (N_10888,N_9221,N_8783);
nand U10889 (N_10889,N_9531,N_9448);
or U10890 (N_10890,N_9167,N_8963);
nor U10891 (N_10891,N_9598,N_9487);
or U10892 (N_10892,N_9824,N_9464);
nand U10893 (N_10893,N_9770,N_9104);
or U10894 (N_10894,N_8894,N_9280);
and U10895 (N_10895,N_9038,N_9264);
and U10896 (N_10896,N_9591,N_9947);
xnor U10897 (N_10897,N_9267,N_9594);
nand U10898 (N_10898,N_9079,N_9529);
or U10899 (N_10899,N_9179,N_9048);
and U10900 (N_10900,N_8806,N_9486);
and U10901 (N_10901,N_9342,N_9349);
xnor U10902 (N_10902,N_9454,N_9967);
nor U10903 (N_10903,N_9063,N_9515);
xnor U10904 (N_10904,N_9464,N_9602);
and U10905 (N_10905,N_9573,N_8770);
xor U10906 (N_10906,N_9523,N_9261);
or U10907 (N_10907,N_9716,N_9689);
xor U10908 (N_10908,N_9037,N_9117);
xnor U10909 (N_10909,N_8845,N_9592);
or U10910 (N_10910,N_9264,N_9978);
nor U10911 (N_10911,N_8964,N_9019);
xnor U10912 (N_10912,N_8808,N_9741);
nor U10913 (N_10913,N_9376,N_9886);
nand U10914 (N_10914,N_9494,N_8842);
or U10915 (N_10915,N_9688,N_9194);
nand U10916 (N_10916,N_9661,N_9641);
xnor U10917 (N_10917,N_9616,N_8894);
or U10918 (N_10918,N_9809,N_9686);
and U10919 (N_10919,N_9174,N_8790);
and U10920 (N_10920,N_9214,N_9249);
or U10921 (N_10921,N_9070,N_9039);
nor U10922 (N_10922,N_9000,N_9891);
and U10923 (N_10923,N_9046,N_9651);
and U10924 (N_10924,N_9249,N_8912);
xnor U10925 (N_10925,N_9881,N_9594);
xor U10926 (N_10926,N_9979,N_9215);
xnor U10927 (N_10927,N_9915,N_9324);
and U10928 (N_10928,N_9542,N_9739);
or U10929 (N_10929,N_9270,N_9300);
nor U10930 (N_10930,N_9051,N_9011);
and U10931 (N_10931,N_9436,N_9811);
xnor U10932 (N_10932,N_9233,N_9025);
nor U10933 (N_10933,N_9098,N_8953);
nor U10934 (N_10934,N_9895,N_9383);
and U10935 (N_10935,N_8915,N_9013);
or U10936 (N_10936,N_8941,N_9580);
or U10937 (N_10937,N_9446,N_9319);
and U10938 (N_10938,N_9177,N_9004);
xor U10939 (N_10939,N_8940,N_9382);
or U10940 (N_10940,N_8908,N_8944);
nand U10941 (N_10941,N_9777,N_9868);
or U10942 (N_10942,N_9377,N_8787);
or U10943 (N_10943,N_9390,N_9592);
nand U10944 (N_10944,N_9000,N_9076);
xnor U10945 (N_10945,N_9529,N_9542);
and U10946 (N_10946,N_9245,N_8972);
and U10947 (N_10947,N_9270,N_9993);
xnor U10948 (N_10948,N_9516,N_9355);
or U10949 (N_10949,N_8771,N_9750);
and U10950 (N_10950,N_9884,N_9221);
xnor U10951 (N_10951,N_8868,N_9705);
nand U10952 (N_10952,N_8886,N_9836);
nand U10953 (N_10953,N_8920,N_8922);
nor U10954 (N_10954,N_8771,N_8973);
or U10955 (N_10955,N_9409,N_9526);
or U10956 (N_10956,N_9254,N_9870);
xor U10957 (N_10957,N_8900,N_9390);
and U10958 (N_10958,N_9969,N_9642);
or U10959 (N_10959,N_9218,N_9601);
nor U10960 (N_10960,N_9842,N_9454);
and U10961 (N_10961,N_9837,N_9117);
nand U10962 (N_10962,N_9120,N_9740);
xor U10963 (N_10963,N_9085,N_8940);
nor U10964 (N_10964,N_9307,N_9589);
or U10965 (N_10965,N_8989,N_8837);
nor U10966 (N_10966,N_9579,N_9276);
or U10967 (N_10967,N_9026,N_9920);
nand U10968 (N_10968,N_9949,N_9656);
nor U10969 (N_10969,N_9941,N_9259);
and U10970 (N_10970,N_9257,N_9029);
nand U10971 (N_10971,N_9797,N_9850);
and U10972 (N_10972,N_9351,N_9262);
nand U10973 (N_10973,N_9433,N_9519);
nor U10974 (N_10974,N_9531,N_8949);
and U10975 (N_10975,N_9743,N_9625);
and U10976 (N_10976,N_9156,N_9030);
xnor U10977 (N_10977,N_8876,N_9824);
nand U10978 (N_10978,N_9727,N_9192);
or U10979 (N_10979,N_9600,N_8771);
nand U10980 (N_10980,N_8797,N_9990);
nor U10981 (N_10981,N_8754,N_9395);
nand U10982 (N_10982,N_9500,N_9363);
or U10983 (N_10983,N_9273,N_9015);
nor U10984 (N_10984,N_9305,N_9480);
nor U10985 (N_10985,N_9014,N_8948);
and U10986 (N_10986,N_9331,N_9153);
xnor U10987 (N_10987,N_9224,N_9213);
and U10988 (N_10988,N_9374,N_9708);
nor U10989 (N_10989,N_9683,N_9278);
and U10990 (N_10990,N_8958,N_9857);
nor U10991 (N_10991,N_9509,N_8805);
xor U10992 (N_10992,N_8992,N_8768);
or U10993 (N_10993,N_9277,N_8864);
and U10994 (N_10994,N_9047,N_9498);
or U10995 (N_10995,N_9071,N_9037);
or U10996 (N_10996,N_9441,N_8872);
xnor U10997 (N_10997,N_9533,N_9187);
and U10998 (N_10998,N_9195,N_8795);
nor U10999 (N_10999,N_9111,N_9673);
nand U11000 (N_11000,N_9106,N_9830);
xnor U11001 (N_11001,N_9803,N_9730);
nor U11002 (N_11002,N_9911,N_9942);
or U11003 (N_11003,N_9162,N_9649);
xor U11004 (N_11004,N_9453,N_9380);
nor U11005 (N_11005,N_8836,N_9801);
and U11006 (N_11006,N_9597,N_9806);
or U11007 (N_11007,N_9331,N_9511);
nand U11008 (N_11008,N_9921,N_9902);
nor U11009 (N_11009,N_9997,N_8815);
xnor U11010 (N_11010,N_8829,N_8822);
or U11011 (N_11011,N_9258,N_9389);
nor U11012 (N_11012,N_9806,N_9621);
xor U11013 (N_11013,N_9195,N_9249);
nor U11014 (N_11014,N_9080,N_9187);
nor U11015 (N_11015,N_9212,N_9985);
nand U11016 (N_11016,N_9470,N_8818);
and U11017 (N_11017,N_9683,N_9791);
nor U11018 (N_11018,N_9273,N_9771);
nor U11019 (N_11019,N_8982,N_9146);
or U11020 (N_11020,N_9735,N_9785);
nand U11021 (N_11021,N_9437,N_9174);
xor U11022 (N_11022,N_9589,N_9248);
xor U11023 (N_11023,N_9741,N_9404);
or U11024 (N_11024,N_9209,N_8982);
or U11025 (N_11025,N_9300,N_9423);
and U11026 (N_11026,N_9665,N_9121);
nand U11027 (N_11027,N_9846,N_9095);
and U11028 (N_11028,N_9873,N_9950);
and U11029 (N_11029,N_9252,N_9497);
nand U11030 (N_11030,N_9216,N_9587);
nand U11031 (N_11031,N_9563,N_8838);
nand U11032 (N_11032,N_9079,N_9839);
nor U11033 (N_11033,N_9253,N_9738);
xnor U11034 (N_11034,N_8920,N_9063);
and U11035 (N_11035,N_9629,N_9671);
xnor U11036 (N_11036,N_9607,N_9921);
nor U11037 (N_11037,N_9679,N_8961);
nor U11038 (N_11038,N_9692,N_9033);
nand U11039 (N_11039,N_9920,N_9350);
or U11040 (N_11040,N_9480,N_9053);
or U11041 (N_11041,N_8841,N_9285);
and U11042 (N_11042,N_9946,N_9776);
nor U11043 (N_11043,N_8776,N_9597);
and U11044 (N_11044,N_9693,N_9339);
nor U11045 (N_11045,N_9219,N_8785);
xor U11046 (N_11046,N_9112,N_8889);
nor U11047 (N_11047,N_9778,N_9236);
and U11048 (N_11048,N_9990,N_9030);
nor U11049 (N_11049,N_9418,N_9582);
xnor U11050 (N_11050,N_8922,N_8961);
or U11051 (N_11051,N_9628,N_9050);
or U11052 (N_11052,N_8968,N_9460);
nor U11053 (N_11053,N_9824,N_9705);
or U11054 (N_11054,N_9149,N_8905);
nor U11055 (N_11055,N_8854,N_8814);
and U11056 (N_11056,N_9848,N_8768);
or U11057 (N_11057,N_9065,N_9250);
and U11058 (N_11058,N_9939,N_9736);
or U11059 (N_11059,N_9775,N_9879);
and U11060 (N_11060,N_9253,N_9859);
or U11061 (N_11061,N_8824,N_9585);
and U11062 (N_11062,N_9748,N_9828);
nor U11063 (N_11063,N_8957,N_9580);
nor U11064 (N_11064,N_9469,N_9082);
and U11065 (N_11065,N_9449,N_9858);
nor U11066 (N_11066,N_9993,N_8768);
and U11067 (N_11067,N_9093,N_9976);
and U11068 (N_11068,N_9472,N_8820);
nor U11069 (N_11069,N_9815,N_9132);
nor U11070 (N_11070,N_9126,N_8769);
nand U11071 (N_11071,N_9040,N_9703);
and U11072 (N_11072,N_8842,N_8830);
nor U11073 (N_11073,N_9180,N_9153);
nand U11074 (N_11074,N_9570,N_9312);
nor U11075 (N_11075,N_9670,N_9202);
xor U11076 (N_11076,N_9645,N_9993);
and U11077 (N_11077,N_9597,N_9711);
and U11078 (N_11078,N_9854,N_9622);
nand U11079 (N_11079,N_9338,N_9786);
nand U11080 (N_11080,N_9123,N_9241);
and U11081 (N_11081,N_9511,N_9120);
xnor U11082 (N_11082,N_9887,N_9129);
nand U11083 (N_11083,N_9651,N_9227);
nand U11084 (N_11084,N_9992,N_9454);
nor U11085 (N_11085,N_9554,N_9281);
nor U11086 (N_11086,N_9617,N_8964);
xnor U11087 (N_11087,N_9551,N_9875);
xnor U11088 (N_11088,N_9663,N_9853);
nor U11089 (N_11089,N_9728,N_9152);
or U11090 (N_11090,N_9643,N_9864);
or U11091 (N_11091,N_9377,N_9750);
or U11092 (N_11092,N_8920,N_9941);
or U11093 (N_11093,N_8952,N_9549);
and U11094 (N_11094,N_9471,N_8861);
nor U11095 (N_11095,N_8963,N_9613);
nand U11096 (N_11096,N_9631,N_9005);
nand U11097 (N_11097,N_9928,N_8794);
xor U11098 (N_11098,N_8871,N_9693);
and U11099 (N_11099,N_9553,N_9557);
nand U11100 (N_11100,N_9892,N_9042);
nand U11101 (N_11101,N_9125,N_9896);
or U11102 (N_11102,N_9248,N_8759);
xor U11103 (N_11103,N_9993,N_9640);
xnor U11104 (N_11104,N_9640,N_9650);
or U11105 (N_11105,N_9843,N_9359);
nor U11106 (N_11106,N_9444,N_9972);
nand U11107 (N_11107,N_9260,N_9727);
or U11108 (N_11108,N_9991,N_9218);
and U11109 (N_11109,N_9147,N_9524);
nor U11110 (N_11110,N_9892,N_9011);
xnor U11111 (N_11111,N_8892,N_9816);
nor U11112 (N_11112,N_9526,N_9797);
nand U11113 (N_11113,N_9767,N_9077);
xnor U11114 (N_11114,N_9367,N_8778);
or U11115 (N_11115,N_9268,N_9446);
nand U11116 (N_11116,N_9360,N_9880);
nand U11117 (N_11117,N_9487,N_8950);
nand U11118 (N_11118,N_9262,N_9381);
xor U11119 (N_11119,N_9456,N_9052);
or U11120 (N_11120,N_9844,N_9384);
nand U11121 (N_11121,N_9209,N_9963);
nand U11122 (N_11122,N_8852,N_9393);
xor U11123 (N_11123,N_9628,N_9568);
or U11124 (N_11124,N_9320,N_8833);
and U11125 (N_11125,N_9329,N_9254);
and U11126 (N_11126,N_9992,N_8989);
nor U11127 (N_11127,N_8819,N_9437);
or U11128 (N_11128,N_9585,N_8851);
and U11129 (N_11129,N_9194,N_9710);
xor U11130 (N_11130,N_9004,N_9871);
nand U11131 (N_11131,N_9437,N_8801);
or U11132 (N_11132,N_9046,N_9944);
xor U11133 (N_11133,N_9017,N_9306);
xor U11134 (N_11134,N_9555,N_9076);
and U11135 (N_11135,N_9296,N_9646);
or U11136 (N_11136,N_9712,N_9449);
and U11137 (N_11137,N_9715,N_8941);
xnor U11138 (N_11138,N_8995,N_9101);
or U11139 (N_11139,N_9700,N_9656);
or U11140 (N_11140,N_9823,N_9708);
nor U11141 (N_11141,N_9810,N_9254);
or U11142 (N_11142,N_9932,N_9921);
and U11143 (N_11143,N_9683,N_9126);
nor U11144 (N_11144,N_9065,N_9301);
and U11145 (N_11145,N_9737,N_9479);
or U11146 (N_11146,N_9939,N_9948);
and U11147 (N_11147,N_8976,N_9404);
and U11148 (N_11148,N_9263,N_8782);
nand U11149 (N_11149,N_9695,N_8838);
nor U11150 (N_11150,N_9410,N_9944);
xnor U11151 (N_11151,N_8811,N_9102);
nor U11152 (N_11152,N_8797,N_9405);
nand U11153 (N_11153,N_8765,N_9157);
nor U11154 (N_11154,N_9765,N_8781);
nand U11155 (N_11155,N_8767,N_9023);
or U11156 (N_11156,N_9907,N_9619);
xnor U11157 (N_11157,N_8967,N_8943);
nand U11158 (N_11158,N_9690,N_9591);
xnor U11159 (N_11159,N_9073,N_9503);
nor U11160 (N_11160,N_9125,N_9853);
nor U11161 (N_11161,N_9048,N_8779);
nor U11162 (N_11162,N_9836,N_9321);
or U11163 (N_11163,N_9107,N_9826);
or U11164 (N_11164,N_8765,N_9622);
xnor U11165 (N_11165,N_9354,N_9837);
or U11166 (N_11166,N_8936,N_9392);
nand U11167 (N_11167,N_9565,N_9031);
xnor U11168 (N_11168,N_9815,N_9610);
or U11169 (N_11169,N_9938,N_8840);
nand U11170 (N_11170,N_9183,N_8981);
nor U11171 (N_11171,N_9279,N_9044);
xor U11172 (N_11172,N_9703,N_9761);
or U11173 (N_11173,N_8875,N_9403);
nor U11174 (N_11174,N_9011,N_9482);
or U11175 (N_11175,N_9533,N_9303);
or U11176 (N_11176,N_8785,N_9391);
and U11177 (N_11177,N_8861,N_9949);
nor U11178 (N_11178,N_9272,N_9441);
and U11179 (N_11179,N_8877,N_9764);
nand U11180 (N_11180,N_9411,N_9735);
or U11181 (N_11181,N_8998,N_9399);
nand U11182 (N_11182,N_9668,N_9175);
nor U11183 (N_11183,N_8974,N_9743);
nor U11184 (N_11184,N_9551,N_9953);
and U11185 (N_11185,N_8841,N_9029);
xor U11186 (N_11186,N_8886,N_9072);
nor U11187 (N_11187,N_9647,N_8854);
nand U11188 (N_11188,N_9104,N_9026);
or U11189 (N_11189,N_9625,N_9631);
and U11190 (N_11190,N_9267,N_9225);
or U11191 (N_11191,N_9602,N_9105);
nand U11192 (N_11192,N_9948,N_9380);
xor U11193 (N_11193,N_9323,N_9712);
or U11194 (N_11194,N_8851,N_8861);
xor U11195 (N_11195,N_9631,N_9781);
nand U11196 (N_11196,N_9991,N_9759);
and U11197 (N_11197,N_9389,N_9631);
or U11198 (N_11198,N_8982,N_9877);
and U11199 (N_11199,N_9140,N_9276);
or U11200 (N_11200,N_8810,N_9318);
nand U11201 (N_11201,N_8767,N_9766);
and U11202 (N_11202,N_9618,N_8964);
nand U11203 (N_11203,N_9549,N_9244);
or U11204 (N_11204,N_9431,N_9645);
or U11205 (N_11205,N_8976,N_8966);
and U11206 (N_11206,N_9459,N_9649);
and U11207 (N_11207,N_8953,N_8750);
or U11208 (N_11208,N_9810,N_9725);
nor U11209 (N_11209,N_9626,N_9555);
and U11210 (N_11210,N_9737,N_9090);
nand U11211 (N_11211,N_9071,N_9851);
nand U11212 (N_11212,N_9598,N_8793);
xor U11213 (N_11213,N_9507,N_9335);
or U11214 (N_11214,N_8920,N_9269);
or U11215 (N_11215,N_8944,N_9913);
nor U11216 (N_11216,N_9825,N_8962);
nor U11217 (N_11217,N_9404,N_9650);
and U11218 (N_11218,N_9338,N_9978);
xor U11219 (N_11219,N_9441,N_9012);
or U11220 (N_11220,N_9977,N_9736);
xnor U11221 (N_11221,N_8993,N_9722);
or U11222 (N_11222,N_8969,N_9883);
or U11223 (N_11223,N_9060,N_9454);
xor U11224 (N_11224,N_9895,N_9843);
nand U11225 (N_11225,N_9164,N_9474);
nand U11226 (N_11226,N_9526,N_9654);
and U11227 (N_11227,N_9943,N_9807);
xor U11228 (N_11228,N_9079,N_9344);
or U11229 (N_11229,N_9298,N_8883);
nand U11230 (N_11230,N_9650,N_9822);
nor U11231 (N_11231,N_9499,N_9680);
nor U11232 (N_11232,N_9809,N_9018);
and U11233 (N_11233,N_9377,N_9413);
and U11234 (N_11234,N_9813,N_9488);
nor U11235 (N_11235,N_9554,N_8798);
and U11236 (N_11236,N_8996,N_9599);
xnor U11237 (N_11237,N_9796,N_9566);
nand U11238 (N_11238,N_9922,N_9784);
xnor U11239 (N_11239,N_9651,N_9535);
nor U11240 (N_11240,N_9657,N_9856);
nor U11241 (N_11241,N_9997,N_9757);
nor U11242 (N_11242,N_9888,N_9767);
or U11243 (N_11243,N_9898,N_8949);
nor U11244 (N_11244,N_9594,N_9898);
or U11245 (N_11245,N_9326,N_9711);
nand U11246 (N_11246,N_9506,N_9794);
nand U11247 (N_11247,N_8817,N_8977);
nand U11248 (N_11248,N_9125,N_8864);
and U11249 (N_11249,N_9858,N_9980);
nor U11250 (N_11250,N_10300,N_10683);
nand U11251 (N_11251,N_11030,N_11134);
nand U11252 (N_11252,N_10768,N_10024);
xnor U11253 (N_11253,N_10250,N_11231);
or U11254 (N_11254,N_11229,N_10177);
xnor U11255 (N_11255,N_10821,N_10132);
xnor U11256 (N_11256,N_10858,N_11100);
nand U11257 (N_11257,N_10744,N_10442);
and U11258 (N_11258,N_10457,N_10546);
or U11259 (N_11259,N_11212,N_11141);
xnor U11260 (N_11260,N_10819,N_11065);
and U11261 (N_11261,N_11014,N_11117);
nor U11262 (N_11262,N_10303,N_11160);
xnor U11263 (N_11263,N_11159,N_11122);
nor U11264 (N_11264,N_11018,N_10071);
nor U11265 (N_11265,N_10023,N_10021);
xnor U11266 (N_11266,N_10319,N_10929);
xnor U11267 (N_11267,N_10262,N_11079);
nand U11268 (N_11268,N_10931,N_10043);
or U11269 (N_11269,N_11230,N_11237);
or U11270 (N_11270,N_10728,N_10597);
nand U11271 (N_11271,N_10778,N_11185);
nand U11272 (N_11272,N_10879,N_10786);
and U11273 (N_11273,N_11011,N_10473);
xor U11274 (N_11274,N_10474,N_10305);
nor U11275 (N_11275,N_10409,N_11202);
xnor U11276 (N_11276,N_10137,N_10689);
and U11277 (N_11277,N_11218,N_10314);
xnor U11278 (N_11278,N_11045,N_10574);
and U11279 (N_11279,N_10708,N_10167);
nor U11280 (N_11280,N_10184,N_10309);
nand U11281 (N_11281,N_10391,N_11094);
xor U11282 (N_11282,N_10567,N_10377);
xor U11283 (N_11283,N_10073,N_10989);
nand U11284 (N_11284,N_10553,N_10990);
xor U11285 (N_11285,N_10948,N_10548);
and U11286 (N_11286,N_10238,N_10783);
nand U11287 (N_11287,N_10290,N_10699);
and U11288 (N_11288,N_11223,N_10555);
xnor U11289 (N_11289,N_10974,N_11188);
xnor U11290 (N_11290,N_10413,N_10185);
or U11291 (N_11291,N_10444,N_10613);
and U11292 (N_11292,N_11196,N_10633);
nand U11293 (N_11293,N_10750,N_10253);
nor U11294 (N_11294,N_10845,N_10440);
xnor U11295 (N_11295,N_10392,N_10153);
and U11296 (N_11296,N_10826,N_11103);
or U11297 (N_11297,N_10266,N_10147);
and U11298 (N_11298,N_10551,N_11001);
nand U11299 (N_11299,N_11056,N_10718);
and U11300 (N_11300,N_10732,N_10631);
nand U11301 (N_11301,N_11204,N_10541);
and U11302 (N_11302,N_10347,N_10471);
xor U11303 (N_11303,N_11038,N_10454);
or U11304 (N_11304,N_10249,N_10124);
or U11305 (N_11305,N_10372,N_10706);
or U11306 (N_11306,N_11126,N_11035);
xor U11307 (N_11307,N_10832,N_10557);
and U11308 (N_11308,N_10014,N_10745);
xnor U11309 (N_11309,N_10885,N_10644);
nand U11310 (N_11310,N_10374,N_11092);
nor U11311 (N_11311,N_11049,N_10010);
xor U11312 (N_11312,N_10403,N_10719);
nor U11313 (N_11313,N_10388,N_10018);
nor U11314 (N_11314,N_10123,N_11099);
xor U11315 (N_11315,N_10316,N_11044);
or U11316 (N_11316,N_10339,N_10582);
nand U11317 (N_11317,N_10459,N_10386);
nand U11318 (N_11318,N_10795,N_11005);
or U11319 (N_11319,N_10060,N_10500);
xnor U11320 (N_11320,N_10489,N_10129);
nor U11321 (N_11321,N_10009,N_10810);
nand U11322 (N_11322,N_10517,N_11215);
and U11323 (N_11323,N_10222,N_10804);
nand U11324 (N_11324,N_10690,N_10201);
and U11325 (N_11325,N_10282,N_11072);
or U11326 (N_11326,N_11187,N_11211);
or U11327 (N_11327,N_10126,N_10875);
and U11328 (N_11328,N_10350,N_10040);
or U11329 (N_11329,N_11095,N_11082);
nand U11330 (N_11330,N_10855,N_10150);
or U11331 (N_11331,N_11124,N_11101);
xor U11332 (N_11332,N_10481,N_10534);
nand U11333 (N_11333,N_11058,N_10439);
or U11334 (N_11334,N_11174,N_10711);
and U11335 (N_11335,N_10315,N_10881);
nor U11336 (N_11336,N_10743,N_10484);
and U11337 (N_11337,N_11000,N_10285);
nor U11338 (N_11338,N_10993,N_10346);
and U11339 (N_11339,N_10790,N_10479);
xor U11340 (N_11340,N_10635,N_10287);
nand U11341 (N_11341,N_10569,N_10994);
nand U11342 (N_11342,N_10427,N_10660);
nand U11343 (N_11343,N_10416,N_10006);
nor U11344 (N_11344,N_10629,N_10306);
and U11345 (N_11345,N_10531,N_11021);
xor U11346 (N_11346,N_10170,N_10692);
xor U11347 (N_11347,N_10142,N_11017);
and U11348 (N_11348,N_10755,N_10550);
or U11349 (N_11349,N_10203,N_10599);
xor U11350 (N_11350,N_11031,N_10687);
nor U11351 (N_11351,N_10779,N_10351);
xor U11352 (N_11352,N_10611,N_11074);
or U11353 (N_11353,N_10322,N_10115);
nand U11354 (N_11354,N_10589,N_10381);
xor U11355 (N_11355,N_10638,N_10894);
xnor U11356 (N_11356,N_10402,N_11020);
nor U11357 (N_11357,N_10095,N_11104);
or U11358 (N_11358,N_10963,N_10691);
xnor U11359 (N_11359,N_10468,N_11144);
xor U11360 (N_11360,N_10776,N_10672);
and U11361 (N_11361,N_10079,N_11243);
xnor U11362 (N_11362,N_10872,N_10664);
xnor U11363 (N_11363,N_10195,N_10164);
xnor U11364 (N_11364,N_11200,N_11029);
and U11365 (N_11365,N_10148,N_10501);
and U11366 (N_11366,N_10463,N_10362);
xnor U11367 (N_11367,N_11197,N_11227);
nor U11368 (N_11368,N_10312,N_10647);
xor U11369 (N_11369,N_11016,N_10280);
and U11370 (N_11370,N_10231,N_10470);
or U11371 (N_11371,N_10458,N_10882);
or U11372 (N_11372,N_10091,N_10332);
nand U11373 (N_11373,N_10625,N_10752);
xor U11374 (N_11374,N_10536,N_11033);
xor U11375 (N_11375,N_10900,N_11151);
and U11376 (N_11376,N_10673,N_10295);
or U11377 (N_11377,N_10601,N_11075);
or U11378 (N_11378,N_10183,N_10450);
nand U11379 (N_11379,N_10982,N_10037);
nand U11380 (N_11380,N_10273,N_10921);
nor U11381 (N_11381,N_10874,N_10966);
nand U11382 (N_11382,N_11039,N_10704);
and U11383 (N_11383,N_10802,N_11125);
and U11384 (N_11384,N_11127,N_10740);
and U11385 (N_11385,N_10587,N_11164);
or U11386 (N_11386,N_11111,N_10051);
and U11387 (N_11387,N_10630,N_10585);
or U11388 (N_11388,N_10063,N_10181);
xnor U11389 (N_11389,N_10724,N_10584);
and U11390 (N_11390,N_11010,N_10674);
nor U11391 (N_11391,N_10429,N_10800);
xnor U11392 (N_11392,N_10256,N_10090);
and U11393 (N_11393,N_10624,N_10056);
nand U11394 (N_11394,N_11064,N_10682);
or U11395 (N_11395,N_10452,N_10632);
nand U11396 (N_11396,N_10572,N_10186);
or U11397 (N_11397,N_10737,N_10277);
or U11398 (N_11398,N_10808,N_10566);
and U11399 (N_11399,N_10760,N_10415);
or U11400 (N_11400,N_11050,N_10862);
and U11401 (N_11401,N_10902,N_10970);
nand U11402 (N_11402,N_10108,N_10722);
xor U11403 (N_11403,N_10431,N_10803);
and U11404 (N_11404,N_10612,N_10816);
or U11405 (N_11405,N_10053,N_10324);
nor U11406 (N_11406,N_10843,N_10485);
and U11407 (N_11407,N_10304,N_10270);
nor U11408 (N_11408,N_10671,N_10155);
xnor U11409 (N_11409,N_11096,N_11036);
xor U11410 (N_11410,N_10087,N_10964);
nor U11411 (N_11411,N_10257,N_10396);
and U11412 (N_11412,N_10478,N_10128);
nor U11413 (N_11413,N_10364,N_10775);
nor U11414 (N_11414,N_11119,N_10999);
nand U11415 (N_11415,N_10941,N_10070);
nor U11416 (N_11416,N_10318,N_10488);
or U11417 (N_11417,N_10038,N_10446);
xor U11418 (N_11418,N_10193,N_10356);
nand U11419 (N_11419,N_10714,N_10017);
nand U11420 (N_11420,N_11097,N_10705);
or U11421 (N_11421,N_10527,N_10157);
or U11422 (N_11422,N_10015,N_10477);
xnor U11423 (N_11423,N_10449,N_10092);
and U11424 (N_11424,N_10552,N_10269);
or U11425 (N_11425,N_10873,N_10221);
xnor U11426 (N_11426,N_10279,N_10437);
and U11427 (N_11427,N_10716,N_10109);
xor U11428 (N_11428,N_10297,N_11047);
nor U11429 (N_11429,N_10748,N_10529);
and U11430 (N_11430,N_10456,N_10972);
and U11431 (N_11431,N_10214,N_10365);
and U11432 (N_11432,N_11172,N_10395);
nand U11433 (N_11433,N_10796,N_10264);
or U11434 (N_11434,N_11087,N_10292);
nand U11435 (N_11435,N_10759,N_10807);
xor U11436 (N_11436,N_11228,N_10676);
xor U11437 (N_11437,N_10204,N_11048);
or U11438 (N_11438,N_10844,N_10588);
or U11439 (N_11439,N_10856,N_10301);
nor U11440 (N_11440,N_10554,N_10665);
xor U11441 (N_11441,N_11246,N_10865);
nand U11442 (N_11442,N_11224,N_10224);
nand U11443 (N_11443,N_10240,N_10048);
xnor U11444 (N_11444,N_11066,N_10219);
and U11445 (N_11445,N_11120,N_10399);
nand U11446 (N_11446,N_11140,N_10663);
nor U11447 (N_11447,N_10729,N_10475);
or U11448 (N_11448,N_10205,N_10887);
nand U11449 (N_11449,N_10892,N_11203);
or U11450 (N_11450,N_10677,N_10945);
xnor U11451 (N_11451,N_10258,N_10739);
nor U11452 (N_11452,N_10507,N_11245);
nor U11453 (N_11453,N_10410,N_10251);
or U11454 (N_11454,N_10940,N_10216);
nand U11455 (N_11455,N_10451,N_10522);
or U11456 (N_11456,N_10684,N_10904);
and U11457 (N_11457,N_10230,N_11062);
or U11458 (N_11458,N_10571,N_10293);
nand U11459 (N_11459,N_10641,N_10189);
xnor U11460 (N_11460,N_10976,N_10893);
nand U11461 (N_11461,N_11162,N_11234);
and U11462 (N_11462,N_10511,N_10762);
xor U11463 (N_11463,N_11091,N_10307);
and U11464 (N_11464,N_10502,N_10514);
nor U11465 (N_11465,N_11163,N_11138);
xnor U11466 (N_11466,N_11239,N_10105);
xor U11467 (N_11467,N_10889,N_10294);
nor U11468 (N_11468,N_10734,N_10031);
and U11469 (N_11469,N_10328,N_10828);
or U11470 (N_11470,N_11154,N_10371);
and U11471 (N_11471,N_10116,N_10149);
xor U11472 (N_11472,N_10104,N_10077);
and U11473 (N_11473,N_10117,N_11106);
and U11474 (N_11474,N_10029,N_10486);
or U11475 (N_11475,N_10561,N_10254);
xor U11476 (N_11476,N_11032,N_10125);
or U11477 (N_11477,N_11123,N_10175);
and U11478 (N_11478,N_10498,N_10311);
and U11479 (N_11479,N_11165,N_10590);
and U11480 (N_11480,N_10370,N_10136);
xnor U11481 (N_11481,N_10131,N_10770);
or U11482 (N_11482,N_10575,N_11051);
xor U11483 (N_11483,N_11040,N_10179);
and U11484 (N_11484,N_10846,N_10138);
nor U11485 (N_11485,N_10841,N_10628);
and U11486 (N_11486,N_11135,N_10606);
xor U11487 (N_11487,N_11086,N_10535);
and U11488 (N_11488,N_10325,N_11057);
and U11489 (N_11489,N_11191,N_10243);
nor U11490 (N_11490,N_10418,N_10905);
or U11491 (N_11491,N_10639,N_10331);
nor U11492 (N_11492,N_10655,N_10906);
nor U11493 (N_11493,N_10504,N_10085);
nand U11494 (N_11494,N_11219,N_10423);
or U11495 (N_11495,N_10642,N_10036);
or U11496 (N_11496,N_10093,N_10291);
xor U11497 (N_11497,N_10560,N_10330);
xnor U11498 (N_11498,N_10637,N_10151);
nand U11499 (N_11499,N_10910,N_10576);
xor U11500 (N_11500,N_10895,N_10919);
nor U11501 (N_11501,N_10525,N_10499);
nor U11502 (N_11502,N_10286,N_10492);
xor U11503 (N_11503,N_10952,N_10605);
or U11504 (N_11504,N_11167,N_10688);
nor U11505 (N_11505,N_10389,N_10035);
xnor U11506 (N_11506,N_10465,N_10333);
and U11507 (N_11507,N_10384,N_10533);
nand U11508 (N_11508,N_10650,N_10933);
nand U11509 (N_11509,N_10842,N_10069);
or U11510 (N_11510,N_11153,N_11176);
nor U11511 (N_11511,N_10352,N_11034);
nand U11512 (N_11512,N_10764,N_10949);
nand U11513 (N_11513,N_10831,N_10382);
xnor U11514 (N_11514,N_10455,N_10114);
and U11515 (N_11515,N_11149,N_10013);
nand U11516 (N_11516,N_10610,N_10788);
or U11517 (N_11517,N_10765,N_10614);
or U11518 (N_11518,N_10738,N_10154);
nor U11519 (N_11519,N_10793,N_10327);
or U11520 (N_11520,N_10275,N_10991);
nor U11521 (N_11521,N_10710,N_11244);
and U11522 (N_11522,N_10074,N_10353);
nor U11523 (N_11523,N_10233,N_11142);
or U11524 (N_11524,N_10202,N_10076);
nand U11525 (N_11525,N_11166,N_10573);
xor U11526 (N_11526,N_11190,N_10022);
nand U11527 (N_11527,N_10354,N_10908);
nor U11528 (N_11528,N_10016,N_10265);
or U11529 (N_11529,N_11027,N_11012);
nor U11530 (N_11530,N_10884,N_10012);
nand U11531 (N_11531,N_10461,N_10857);
nor U11532 (N_11532,N_10834,N_10996);
and U11533 (N_11533,N_10656,N_11109);
and U11534 (N_11534,N_10135,N_10443);
nand U11535 (N_11535,N_10696,N_11004);
nor U11536 (N_11536,N_10196,N_10246);
or U11537 (N_11537,N_10133,N_10868);
nand U11538 (N_11538,N_10827,N_10646);
nor U11539 (N_11539,N_10595,N_10695);
and U11540 (N_11540,N_10958,N_10234);
nand U11541 (N_11541,N_10206,N_10886);
and U11542 (N_11542,N_10955,N_11222);
nor U11543 (N_11543,N_10782,N_11114);
and U11544 (N_11544,N_10944,N_10797);
xnor U11545 (N_11545,N_10068,N_10420);
or U11546 (N_11546,N_10447,N_10947);
xor U11547 (N_11547,N_10707,N_10220);
nand U11548 (N_11548,N_11139,N_10348);
and U11549 (N_11549,N_11242,N_11150);
nand U11550 (N_11550,N_10918,N_10727);
xnor U11551 (N_11551,N_10122,N_11078);
nor U11552 (N_11552,N_10592,N_10667);
nor U11553 (N_11553,N_10191,N_10995);
or U11554 (N_11554,N_10713,N_10515);
and U11555 (N_11555,N_10008,N_10101);
and U11556 (N_11556,N_10494,N_10658);
nor U11557 (N_11557,N_11080,N_10594);
or U11558 (N_11558,N_10143,N_10603);
xnor U11559 (N_11559,N_10987,N_10602);
or U11560 (N_11560,N_10049,N_10657);
nor U11561 (N_11561,N_10368,N_10888);
or U11562 (N_11562,N_10239,N_10397);
nand U11563 (N_11563,N_10961,N_10953);
nor U11564 (N_11564,N_10361,N_11248);
and U11565 (N_11565,N_10213,N_10914);
xnor U11566 (N_11566,N_10299,N_10758);
xor U11567 (N_11567,N_10199,N_10390);
and U11568 (N_11568,N_10472,N_10980);
xnor U11569 (N_11569,N_10067,N_11148);
nor U11570 (N_11570,N_11077,N_10245);
nand U11571 (N_11571,N_10767,N_10957);
nand U11572 (N_11572,N_10120,N_10913);
and U11573 (N_11573,N_10530,N_11023);
nor U11574 (N_11574,N_10441,N_10815);
and U11575 (N_11575,N_10398,N_10385);
xnor U11576 (N_11576,N_10380,N_10032);
or U11577 (N_11577,N_10626,N_10259);
and U11578 (N_11578,N_10055,N_10824);
nand U11579 (N_11579,N_10877,N_10697);
or U11580 (N_11580,N_10047,N_10805);
nor U11581 (N_11581,N_11178,N_10172);
nand U11582 (N_11582,N_10469,N_10025);
or U11583 (N_11583,N_10518,N_11085);
nor U11584 (N_11584,N_11037,N_10591);
and U11585 (N_11585,N_10538,N_10360);
nand U11586 (N_11586,N_10645,N_11076);
and U11587 (N_11587,N_10891,N_10345);
nor U11588 (N_11588,N_10806,N_10519);
xnor U11589 (N_11589,N_10822,N_11024);
and U11590 (N_11590,N_10973,N_10383);
nand U11591 (N_11591,N_10627,N_10621);
nand U11592 (N_11592,N_11088,N_11067);
xnor U11593 (N_11593,N_10263,N_10281);
nor U11594 (N_11594,N_11093,N_10198);
xor U11595 (N_11595,N_11006,N_10011);
or U11596 (N_11596,N_10897,N_10366);
xor U11597 (N_11597,N_10864,N_10769);
or U11598 (N_11598,N_11208,N_10742);
nor U11599 (N_11599,N_10419,N_10041);
xor U11600 (N_11600,N_11136,N_10811);
nand U11601 (N_11601,N_10814,N_10866);
nand U11602 (N_11602,N_11207,N_10753);
or U11603 (N_11603,N_10227,N_10180);
or U11604 (N_11604,N_10833,N_10083);
nand U11605 (N_11605,N_10118,N_10661);
nor U11606 (N_11606,N_10237,N_10241);
and U11607 (N_11607,N_10559,N_10171);
nor U11608 (N_11608,N_11184,N_10867);
nand U11609 (N_11609,N_10190,N_10242);
xnor U11610 (N_11610,N_11108,N_10939);
or U11611 (N_11611,N_11173,N_10825);
and U11612 (N_11612,N_10720,N_10809);
xor U11613 (N_11613,N_10448,N_11081);
xnor U11614 (N_11614,N_10408,N_11061);
nor U11615 (N_11615,N_11009,N_10176);
nor U11616 (N_11616,N_10852,N_11249);
and U11617 (N_11617,N_11131,N_10166);
xor U11618 (N_11618,N_10917,N_11180);
nor U11619 (N_11619,N_10777,N_10730);
nor U11620 (N_11620,N_10899,N_10404);
xnor U11621 (N_11621,N_11143,N_10033);
nand U11622 (N_11622,N_10977,N_10901);
or U11623 (N_11623,N_10562,N_10100);
and U11624 (N_11624,N_10424,N_10218);
and U11625 (N_11625,N_11169,N_11003);
nand U11626 (N_11626,N_10757,N_10912);
and U11627 (N_11627,N_10247,N_10969);
and U11628 (N_11628,N_10523,N_10476);
nor U11629 (N_11629,N_10653,N_10934);
or U11630 (N_11630,N_10820,N_11046);
nand U11631 (N_11631,N_10462,N_10144);
nor U11632 (N_11632,N_10088,N_10721);
nand U11633 (N_11633,N_10784,N_10935);
and U11634 (N_11634,N_10062,N_10871);
nand U11635 (N_11635,N_10435,N_10042);
nand U11636 (N_11636,N_11022,N_10583);
nor U11637 (N_11637,N_10159,N_10978);
or U11638 (N_11638,N_10986,N_11225);
nand U11639 (N_11639,N_10057,N_10414);
nor U11640 (N_11640,N_10607,N_10799);
and U11641 (N_11641,N_10173,N_10979);
nand U11642 (N_11642,N_10421,N_10680);
or U11643 (N_11643,N_10344,N_10103);
nor U11644 (N_11644,N_10428,N_10493);
nand U11645 (N_11645,N_10323,N_10197);
or U11646 (N_11646,N_10508,N_10640);
nand U11647 (N_11647,N_10460,N_10836);
xnor U11648 (N_11648,N_10054,N_10618);
xnor U11649 (N_11649,N_10355,N_10211);
nand U11650 (N_11650,N_10787,N_10001);
xnor U11651 (N_11651,N_10066,N_10229);
xnor U11652 (N_11652,N_10102,N_10712);
or U11653 (N_11653,N_10997,N_10308);
xnor U11654 (N_11654,N_10425,N_10225);
and U11655 (N_11655,N_10542,N_11026);
or U11656 (N_11656,N_10608,N_10127);
xnor U11657 (N_11657,N_10169,N_10310);
nand U11658 (N_11658,N_10400,N_10453);
xor U11659 (N_11659,N_10537,N_10524);
and U11660 (N_11660,N_11220,N_10878);
nand U11661 (N_11661,N_10698,N_10194);
nand U11662 (N_11662,N_10920,N_10505);
nand U11663 (N_11663,N_11083,N_10210);
nand U11664 (N_11664,N_10916,N_10593);
xor U11665 (N_11665,N_11028,N_10766);
and U11666 (N_11666,N_10731,N_10369);
nand U11667 (N_11667,N_10089,N_10061);
nand U11668 (N_11668,N_10097,N_10984);
xor U11669 (N_11669,N_11069,N_10110);
or U11670 (N_11670,N_11137,N_10526);
and U11671 (N_11671,N_10178,N_10785);
nand U11672 (N_11672,N_10998,N_10174);
nand U11673 (N_11673,N_11121,N_10558);
and U11674 (N_11674,N_10643,N_10046);
xnor U11675 (N_11675,N_11226,N_10791);
and U11676 (N_11676,N_10848,N_10387);
nor U11677 (N_11677,N_10094,N_10340);
nor U11678 (N_11678,N_10938,N_10539);
nor U11679 (N_11679,N_10975,N_10107);
xnor U11680 (N_11680,N_11233,N_11055);
or U11681 (N_11681,N_10649,N_10072);
nand U11682 (N_11682,N_10432,N_10545);
and U11683 (N_11683,N_10436,N_11145);
and U11684 (N_11684,N_10715,N_10495);
nand U11685 (N_11685,N_10121,N_11155);
nand U11686 (N_11686,N_10326,N_11177);
xor U11687 (N_11687,N_10491,N_11007);
xor U11688 (N_11688,N_11199,N_10276);
or U11689 (N_11689,N_11210,N_10774);
nand U11690 (N_11690,N_10223,N_11008);
or U11691 (N_11691,N_10965,N_10598);
nand U11692 (N_11692,N_11201,N_10907);
and U11693 (N_11693,N_10433,N_10763);
nand U11694 (N_11694,N_10394,N_10510);
xor U11695 (N_11695,N_10749,N_10754);
and U11696 (N_11696,N_11182,N_10577);
nand U11697 (N_11697,N_11175,N_10792);
and U11698 (N_11698,N_11052,N_10565);
xnor U11699 (N_11699,N_10373,N_10761);
or U11700 (N_11700,N_10840,N_11132);
nor U11701 (N_11701,N_10623,N_10968);
or U11702 (N_11702,N_10798,N_11171);
nor U11703 (N_11703,N_10532,N_10430);
or U11704 (N_11704,N_10570,N_10823);
xor U11705 (N_11705,N_11043,N_11054);
nor U11706 (N_11706,N_10951,N_10839);
xnor U11707 (N_11707,N_10052,N_10751);
nor U11708 (N_11708,N_10943,N_11157);
xnor U11709 (N_11709,N_10932,N_10268);
nor U11710 (N_11710,N_10870,N_10516);
or U11711 (N_11711,N_10379,N_10813);
and U11712 (N_11712,N_10735,N_10564);
and U11713 (N_11713,N_10119,N_10039);
or U11714 (N_11714,N_10685,N_10981);
and U11715 (N_11715,N_10165,N_10417);
nand U11716 (N_11716,N_10506,N_10771);
or U11717 (N_11717,N_10876,N_10668);
or U11718 (N_11718,N_10869,N_10426);
xor U11719 (N_11719,N_10342,N_10686);
or U11720 (N_11720,N_10000,N_10817);
and U11721 (N_11721,N_10600,N_10634);
xor U11722 (N_11722,N_10781,N_11113);
or U11723 (N_11723,N_10863,N_10080);
nand U11724 (N_11724,N_10956,N_10509);
nor U11725 (N_11725,N_10134,N_10925);
xor U11726 (N_11726,N_10544,N_10217);
or U11727 (N_11727,N_11098,N_11156);
or U11728 (N_11728,N_10146,N_10075);
xnor U11729 (N_11729,N_10106,N_10329);
xor U11730 (N_11730,N_11060,N_11129);
or U11731 (N_11731,N_10700,N_10670);
nor U11732 (N_11732,N_11183,N_10694);
nor U11733 (N_11733,N_10983,N_11089);
nand U11734 (N_11734,N_10801,N_10675);
xor U11735 (N_11735,N_10849,N_11002);
and U11736 (N_11736,N_10349,N_10082);
nand U11737 (N_11737,N_10378,N_11105);
nor U11738 (N_11738,N_10909,N_10065);
or U11739 (N_11739,N_10512,N_10651);
xnor U11740 (N_11740,N_10928,N_10438);
nand U11741 (N_11741,N_10226,N_10654);
nand U11742 (N_11742,N_11102,N_10992);
nand U11743 (N_11743,N_11189,N_10622);
nor U11744 (N_11744,N_10411,N_10313);
and U11745 (N_11745,N_10890,N_10335);
nand U11746 (N_11746,N_10099,N_10019);
and U11747 (N_11747,N_10261,N_11192);
nand U11748 (N_11748,N_10289,N_10703);
nor U11749 (N_11749,N_10837,N_10407);
and U11750 (N_11750,N_10139,N_10596);
nor U11751 (N_11751,N_10003,N_10026);
nand U11752 (N_11752,N_10212,N_10232);
nor U11753 (N_11753,N_10283,N_10861);
and U11754 (N_11754,N_10208,N_10467);
or U11755 (N_11755,N_10922,N_11130);
nor U11756 (N_11756,N_10883,N_10278);
xor U11757 (N_11757,N_10942,N_10528);
nor U11758 (N_11758,N_11025,N_11205);
xor U11759 (N_11759,N_11247,N_10375);
nor U11760 (N_11760,N_11198,N_10847);
xnor U11761 (N_11761,N_10678,N_10434);
and U11762 (N_11762,N_10096,N_10860);
and U11763 (N_11763,N_11070,N_10568);
xor U11764 (N_11764,N_10367,N_11170);
or U11765 (N_11765,N_11073,N_10636);
xnor U11766 (N_11766,N_11193,N_10343);
nand U11767 (N_11767,N_11158,N_10236);
nand U11768 (N_11768,N_10005,N_10985);
or U11769 (N_11769,N_10248,N_11084);
and U11770 (N_11770,N_10556,N_10609);
nand U11771 (N_11771,N_10662,N_10255);
and U11772 (N_11772,N_10746,N_10896);
or U11773 (N_11773,N_10112,N_10818);
xor U11774 (N_11774,N_10002,N_10543);
and U11775 (N_11775,N_10487,N_10152);
or U11776 (N_11776,N_11214,N_10702);
nand U11777 (N_11777,N_11118,N_10274);
and U11778 (N_11778,N_10926,N_11186);
nand U11779 (N_11779,N_10617,N_11241);
nor U11780 (N_11780,N_10619,N_10004);
and U11781 (N_11781,N_10464,N_10679);
and U11782 (N_11782,N_10923,N_10959);
and U11783 (N_11783,N_10086,N_10401);
nand U11784 (N_11784,N_10579,N_10334);
and U11785 (N_11785,N_10497,N_10717);
or U11786 (N_11786,N_10406,N_10158);
nand U11787 (N_11787,N_11221,N_10563);
nor U11788 (N_11788,N_10228,N_11181);
nor U11789 (N_11789,N_10780,N_10341);
and U11790 (N_11790,N_10967,N_10701);
nor U11791 (N_11791,N_10520,N_10028);
nand U11792 (N_11792,N_10483,N_10988);
and U11793 (N_11793,N_10578,N_10272);
xnor U11794 (N_11794,N_11107,N_10681);
nand U11795 (N_11795,N_11146,N_10163);
xnor U11796 (N_11796,N_10773,N_11179);
or U11797 (N_11797,N_10405,N_10244);
and U11798 (N_11798,N_10496,N_10581);
xnor U11799 (N_11799,N_10880,N_10726);
or U11800 (N_11800,N_10412,N_11168);
xor U11801 (N_11801,N_10209,N_10971);
or U11802 (N_11802,N_10937,N_10480);
nor U11803 (N_11803,N_11112,N_10020);
or U11804 (N_11804,N_11071,N_10915);
xor U11805 (N_11805,N_10260,N_10376);
nand U11806 (N_11806,N_10188,N_10747);
or U11807 (N_11807,N_10187,N_10288);
nor U11808 (N_11808,N_10050,N_10741);
or U11809 (N_11809,N_10320,N_11235);
xnor U11810 (N_11810,N_11013,N_10669);
xor U11811 (N_11811,N_11133,N_10267);
or U11812 (N_11812,N_10693,N_10911);
xnor U11813 (N_11813,N_10338,N_11206);
or U11814 (N_11814,N_10363,N_11147);
nor U11815 (N_11815,N_10161,N_10359);
nor U11816 (N_11816,N_10789,N_10829);
or U11817 (N_11817,N_10547,N_10903);
or U11818 (N_11818,N_10207,N_10298);
and U11819 (N_11819,N_10358,N_10513);
and U11820 (N_11820,N_10736,N_10111);
or U11821 (N_11821,N_10044,N_10098);
nand U11822 (N_11822,N_11019,N_10081);
nand U11823 (N_11823,N_10182,N_10393);
nand U11824 (N_11824,N_10859,N_11042);
xnor U11825 (N_11825,N_10058,N_10296);
nor U11826 (N_11826,N_10215,N_10130);
or U11827 (N_11827,N_11194,N_10252);
or U11828 (N_11828,N_11238,N_10027);
xor U11829 (N_11829,N_11116,N_11216);
xor U11830 (N_11830,N_10007,N_10930);
and U11831 (N_11831,N_10954,N_11059);
nand U11832 (N_11832,N_10666,N_10615);
nor U11833 (N_11833,N_10604,N_11068);
and U11834 (N_11834,N_10140,N_10851);
and U11835 (N_11835,N_11015,N_10337);
nand U11836 (N_11836,N_10652,N_10659);
nand U11837 (N_11837,N_10924,N_11213);
xor U11838 (N_11838,N_10302,N_10113);
xor U11839 (N_11839,N_10616,N_10145);
and U11840 (N_11840,N_11240,N_10962);
or U11841 (N_11841,N_10549,N_10192);
nor U11842 (N_11842,N_10064,N_10540);
and U11843 (N_11843,N_11195,N_10357);
xor U11844 (N_11844,N_10835,N_10830);
xnor U11845 (N_11845,N_10284,N_10723);
and U11846 (N_11846,N_10725,N_10162);
and U11847 (N_11847,N_10927,N_10466);
xnor U11848 (N_11848,N_10482,N_10045);
or U11849 (N_11849,N_10490,N_10838);
and U11850 (N_11850,N_10271,N_11236);
and U11851 (N_11851,N_10034,N_11110);
nor U11852 (N_11852,N_10709,N_10812);
or U11853 (N_11853,N_11115,N_11041);
xnor U11854 (N_11854,N_11161,N_10521);
or U11855 (N_11855,N_10946,N_10580);
nor U11856 (N_11856,N_11209,N_10936);
nand U11857 (N_11857,N_10772,N_10898);
and U11858 (N_11858,N_10620,N_10960);
xor U11859 (N_11859,N_10235,N_11090);
nor U11860 (N_11860,N_10648,N_11217);
and U11861 (N_11861,N_10794,N_10850);
or U11862 (N_11862,N_10853,N_10321);
or U11863 (N_11863,N_10854,N_11128);
nor U11864 (N_11864,N_10200,N_11063);
nor U11865 (N_11865,N_10030,N_11232);
and U11866 (N_11866,N_10733,N_10141);
xnor U11867 (N_11867,N_10586,N_11053);
nor U11868 (N_11868,N_10950,N_10168);
nand U11869 (N_11869,N_10445,N_10317);
nand U11870 (N_11870,N_10422,N_10503);
nor U11871 (N_11871,N_10078,N_10756);
and U11872 (N_11872,N_10059,N_10084);
and U11873 (N_11873,N_10160,N_10156);
nand U11874 (N_11874,N_11152,N_10336);
xor U11875 (N_11875,N_10266,N_10784);
nand U11876 (N_11876,N_10178,N_10564);
xor U11877 (N_11877,N_10203,N_10393);
xor U11878 (N_11878,N_10672,N_10845);
nor U11879 (N_11879,N_11100,N_11002);
nand U11880 (N_11880,N_11130,N_10022);
xnor U11881 (N_11881,N_10530,N_10568);
xor U11882 (N_11882,N_10980,N_10067);
nand U11883 (N_11883,N_10972,N_10092);
or U11884 (N_11884,N_11107,N_11003);
nor U11885 (N_11885,N_10035,N_10363);
xor U11886 (N_11886,N_10427,N_10689);
and U11887 (N_11887,N_10279,N_10108);
nor U11888 (N_11888,N_11150,N_10681);
nand U11889 (N_11889,N_10116,N_10481);
nand U11890 (N_11890,N_10197,N_10209);
nand U11891 (N_11891,N_10716,N_10028);
or U11892 (N_11892,N_10968,N_10367);
and U11893 (N_11893,N_10312,N_11139);
xnor U11894 (N_11894,N_10184,N_10281);
or U11895 (N_11895,N_10187,N_11138);
xnor U11896 (N_11896,N_11039,N_10798);
nand U11897 (N_11897,N_11123,N_10288);
and U11898 (N_11898,N_10613,N_10099);
nor U11899 (N_11899,N_10865,N_10350);
or U11900 (N_11900,N_10804,N_10580);
nand U11901 (N_11901,N_10112,N_11157);
nor U11902 (N_11902,N_10704,N_11172);
and U11903 (N_11903,N_11193,N_10810);
or U11904 (N_11904,N_10999,N_10001);
xor U11905 (N_11905,N_10548,N_10898);
and U11906 (N_11906,N_10007,N_10211);
nor U11907 (N_11907,N_10386,N_10594);
xnor U11908 (N_11908,N_10640,N_10513);
nand U11909 (N_11909,N_10317,N_10585);
xor U11910 (N_11910,N_10901,N_10243);
or U11911 (N_11911,N_10155,N_10420);
or U11912 (N_11912,N_10711,N_10079);
nor U11913 (N_11913,N_10305,N_10216);
xnor U11914 (N_11914,N_11150,N_11240);
or U11915 (N_11915,N_10829,N_10395);
nand U11916 (N_11916,N_10497,N_10219);
and U11917 (N_11917,N_10078,N_10375);
and U11918 (N_11918,N_10292,N_10201);
or U11919 (N_11919,N_10439,N_10283);
nand U11920 (N_11920,N_10185,N_10348);
or U11921 (N_11921,N_10285,N_10989);
xor U11922 (N_11922,N_10838,N_10593);
and U11923 (N_11923,N_10178,N_11103);
xnor U11924 (N_11924,N_10953,N_10907);
nor U11925 (N_11925,N_10597,N_10330);
and U11926 (N_11926,N_10436,N_10587);
and U11927 (N_11927,N_11200,N_11130);
or U11928 (N_11928,N_10165,N_10109);
nor U11929 (N_11929,N_10503,N_10797);
nor U11930 (N_11930,N_11031,N_10783);
xnor U11931 (N_11931,N_10721,N_10504);
xor U11932 (N_11932,N_10325,N_10463);
xor U11933 (N_11933,N_10264,N_10452);
nor U11934 (N_11934,N_11047,N_10164);
and U11935 (N_11935,N_10215,N_10018);
or U11936 (N_11936,N_10329,N_10097);
xor U11937 (N_11937,N_11188,N_10828);
nand U11938 (N_11938,N_10434,N_10599);
or U11939 (N_11939,N_10667,N_10814);
xnor U11940 (N_11940,N_11146,N_10662);
xor U11941 (N_11941,N_10562,N_10518);
nand U11942 (N_11942,N_11040,N_11016);
nor U11943 (N_11943,N_10019,N_10540);
or U11944 (N_11944,N_10311,N_10844);
xnor U11945 (N_11945,N_10969,N_10885);
nand U11946 (N_11946,N_10922,N_11065);
or U11947 (N_11947,N_10950,N_10081);
xnor U11948 (N_11948,N_10977,N_10675);
and U11949 (N_11949,N_10247,N_10185);
nor U11950 (N_11950,N_10948,N_10392);
and U11951 (N_11951,N_11121,N_10465);
or U11952 (N_11952,N_11067,N_10814);
or U11953 (N_11953,N_11110,N_11045);
nand U11954 (N_11954,N_10573,N_11050);
and U11955 (N_11955,N_10893,N_10189);
or U11956 (N_11956,N_10343,N_11101);
nor U11957 (N_11957,N_10185,N_10575);
xnor U11958 (N_11958,N_10795,N_10038);
or U11959 (N_11959,N_10635,N_10690);
or U11960 (N_11960,N_10661,N_10382);
nor U11961 (N_11961,N_10001,N_11203);
or U11962 (N_11962,N_10623,N_10074);
xor U11963 (N_11963,N_10508,N_10602);
xnor U11964 (N_11964,N_10286,N_10094);
xor U11965 (N_11965,N_10228,N_10857);
or U11966 (N_11966,N_10557,N_10391);
or U11967 (N_11967,N_10092,N_10581);
and U11968 (N_11968,N_11158,N_10354);
and U11969 (N_11969,N_11139,N_11176);
and U11970 (N_11970,N_10518,N_10085);
xnor U11971 (N_11971,N_10176,N_11176);
and U11972 (N_11972,N_10100,N_11201);
or U11973 (N_11973,N_10612,N_10279);
nand U11974 (N_11974,N_10299,N_10889);
xor U11975 (N_11975,N_10125,N_10729);
or U11976 (N_11976,N_10352,N_10328);
or U11977 (N_11977,N_10695,N_10884);
nand U11978 (N_11978,N_10674,N_10634);
nor U11979 (N_11979,N_10060,N_10390);
and U11980 (N_11980,N_10050,N_10063);
nand U11981 (N_11981,N_10991,N_10326);
and U11982 (N_11982,N_10963,N_10259);
and U11983 (N_11983,N_11177,N_10862);
and U11984 (N_11984,N_10018,N_10325);
nand U11985 (N_11985,N_10530,N_10760);
or U11986 (N_11986,N_10574,N_10840);
nor U11987 (N_11987,N_10970,N_10589);
nor U11988 (N_11988,N_10476,N_10820);
xor U11989 (N_11989,N_10053,N_11111);
nand U11990 (N_11990,N_10737,N_10831);
nor U11991 (N_11991,N_10264,N_10780);
nand U11992 (N_11992,N_11053,N_10792);
or U11993 (N_11993,N_10631,N_11025);
xnor U11994 (N_11994,N_10437,N_10808);
or U11995 (N_11995,N_10366,N_10405);
and U11996 (N_11996,N_11230,N_10444);
and U11997 (N_11997,N_10364,N_10799);
and U11998 (N_11998,N_11136,N_11100);
and U11999 (N_11999,N_11212,N_10249);
nand U12000 (N_12000,N_10590,N_10365);
or U12001 (N_12001,N_10758,N_10349);
xnor U12002 (N_12002,N_10887,N_10984);
nand U12003 (N_12003,N_10476,N_10235);
nand U12004 (N_12004,N_11014,N_10290);
nand U12005 (N_12005,N_10742,N_10795);
xor U12006 (N_12006,N_10404,N_11240);
or U12007 (N_12007,N_11065,N_10228);
or U12008 (N_12008,N_11061,N_10168);
nand U12009 (N_12009,N_11181,N_10869);
nand U12010 (N_12010,N_10398,N_10735);
or U12011 (N_12011,N_10166,N_10242);
nor U12012 (N_12012,N_10095,N_10496);
nand U12013 (N_12013,N_10647,N_10836);
nand U12014 (N_12014,N_11162,N_10671);
nor U12015 (N_12015,N_10197,N_10096);
or U12016 (N_12016,N_10043,N_10378);
xnor U12017 (N_12017,N_10644,N_11117);
xor U12018 (N_12018,N_10893,N_10884);
and U12019 (N_12019,N_11028,N_10748);
nand U12020 (N_12020,N_11133,N_10562);
nand U12021 (N_12021,N_10416,N_10524);
or U12022 (N_12022,N_10692,N_11042);
nor U12023 (N_12023,N_10530,N_10208);
or U12024 (N_12024,N_10067,N_11012);
nand U12025 (N_12025,N_10046,N_11057);
and U12026 (N_12026,N_10744,N_10175);
and U12027 (N_12027,N_10172,N_10126);
nand U12028 (N_12028,N_10123,N_10913);
nor U12029 (N_12029,N_10862,N_10585);
nand U12030 (N_12030,N_10625,N_10145);
or U12031 (N_12031,N_10948,N_10328);
nand U12032 (N_12032,N_10364,N_11121);
nor U12033 (N_12033,N_10880,N_10606);
nor U12034 (N_12034,N_10643,N_10192);
or U12035 (N_12035,N_10642,N_11191);
xnor U12036 (N_12036,N_11082,N_10992);
xor U12037 (N_12037,N_10779,N_10851);
xor U12038 (N_12038,N_10791,N_10175);
and U12039 (N_12039,N_11219,N_10993);
and U12040 (N_12040,N_10934,N_10986);
nor U12041 (N_12041,N_10218,N_11015);
nor U12042 (N_12042,N_10723,N_10971);
or U12043 (N_12043,N_10647,N_10889);
nor U12044 (N_12044,N_10169,N_10864);
or U12045 (N_12045,N_10209,N_10127);
or U12046 (N_12046,N_10559,N_10599);
nand U12047 (N_12047,N_10663,N_10544);
xnor U12048 (N_12048,N_10101,N_10537);
or U12049 (N_12049,N_10878,N_10459);
nor U12050 (N_12050,N_10748,N_11234);
and U12051 (N_12051,N_10336,N_10503);
xnor U12052 (N_12052,N_10652,N_11174);
xnor U12053 (N_12053,N_10539,N_10313);
nor U12054 (N_12054,N_10172,N_10045);
and U12055 (N_12055,N_10269,N_10323);
nand U12056 (N_12056,N_10615,N_10621);
and U12057 (N_12057,N_10866,N_10224);
nand U12058 (N_12058,N_11132,N_10465);
xor U12059 (N_12059,N_11143,N_11103);
and U12060 (N_12060,N_10699,N_10193);
and U12061 (N_12061,N_10254,N_11214);
or U12062 (N_12062,N_11043,N_11215);
xor U12063 (N_12063,N_11028,N_11213);
and U12064 (N_12064,N_10864,N_10609);
nand U12065 (N_12065,N_10618,N_10446);
and U12066 (N_12066,N_10124,N_10691);
xor U12067 (N_12067,N_10468,N_11085);
nand U12068 (N_12068,N_10576,N_10722);
and U12069 (N_12069,N_11111,N_10751);
nand U12070 (N_12070,N_10337,N_10177);
nor U12071 (N_12071,N_10555,N_10864);
nor U12072 (N_12072,N_10887,N_10592);
or U12073 (N_12073,N_10520,N_10491);
nand U12074 (N_12074,N_10441,N_10709);
or U12075 (N_12075,N_10501,N_10571);
nand U12076 (N_12076,N_10626,N_10954);
nand U12077 (N_12077,N_10535,N_10497);
and U12078 (N_12078,N_11078,N_10510);
or U12079 (N_12079,N_10822,N_11021);
and U12080 (N_12080,N_10352,N_10946);
nor U12081 (N_12081,N_11021,N_10701);
or U12082 (N_12082,N_10845,N_10076);
or U12083 (N_12083,N_10109,N_10861);
xnor U12084 (N_12084,N_10018,N_10790);
or U12085 (N_12085,N_10788,N_10455);
or U12086 (N_12086,N_10753,N_11074);
nand U12087 (N_12087,N_10923,N_10135);
xnor U12088 (N_12088,N_10625,N_11118);
or U12089 (N_12089,N_10488,N_11207);
nor U12090 (N_12090,N_10115,N_10645);
and U12091 (N_12091,N_11125,N_11036);
nor U12092 (N_12092,N_10703,N_10898);
and U12093 (N_12093,N_10378,N_10534);
and U12094 (N_12094,N_11073,N_10388);
nand U12095 (N_12095,N_10934,N_10120);
nor U12096 (N_12096,N_10823,N_10216);
xor U12097 (N_12097,N_10778,N_10940);
nand U12098 (N_12098,N_10085,N_11039);
and U12099 (N_12099,N_10815,N_10725);
nor U12100 (N_12100,N_10265,N_10731);
xor U12101 (N_12101,N_10553,N_10318);
nor U12102 (N_12102,N_10534,N_10612);
xor U12103 (N_12103,N_10758,N_10251);
nand U12104 (N_12104,N_10425,N_10227);
and U12105 (N_12105,N_10348,N_10355);
and U12106 (N_12106,N_10055,N_10778);
nand U12107 (N_12107,N_10137,N_10903);
nand U12108 (N_12108,N_10690,N_11002);
and U12109 (N_12109,N_10170,N_11096);
xnor U12110 (N_12110,N_10522,N_10834);
and U12111 (N_12111,N_10389,N_10891);
nand U12112 (N_12112,N_11146,N_10125);
and U12113 (N_12113,N_10430,N_10527);
xnor U12114 (N_12114,N_11152,N_10041);
nand U12115 (N_12115,N_10755,N_11152);
and U12116 (N_12116,N_11135,N_11025);
xnor U12117 (N_12117,N_10949,N_10158);
nand U12118 (N_12118,N_10879,N_10980);
xor U12119 (N_12119,N_11105,N_10401);
or U12120 (N_12120,N_10871,N_10457);
or U12121 (N_12121,N_11234,N_10454);
nor U12122 (N_12122,N_10414,N_11166);
and U12123 (N_12123,N_10665,N_10234);
or U12124 (N_12124,N_11210,N_10529);
or U12125 (N_12125,N_10659,N_10014);
and U12126 (N_12126,N_10106,N_10420);
nor U12127 (N_12127,N_11161,N_10272);
xnor U12128 (N_12128,N_10068,N_10433);
or U12129 (N_12129,N_10278,N_10132);
nand U12130 (N_12130,N_10093,N_10477);
or U12131 (N_12131,N_10423,N_11093);
nand U12132 (N_12132,N_10464,N_10448);
or U12133 (N_12133,N_10956,N_10136);
xor U12134 (N_12134,N_10369,N_10400);
nand U12135 (N_12135,N_10240,N_10543);
xor U12136 (N_12136,N_10328,N_10788);
and U12137 (N_12137,N_11185,N_11124);
nor U12138 (N_12138,N_10098,N_10778);
xnor U12139 (N_12139,N_10552,N_11005);
xor U12140 (N_12140,N_10110,N_10516);
or U12141 (N_12141,N_10015,N_10088);
xnor U12142 (N_12142,N_11096,N_10146);
nand U12143 (N_12143,N_10377,N_10577);
nor U12144 (N_12144,N_10513,N_10447);
and U12145 (N_12145,N_10549,N_10825);
or U12146 (N_12146,N_10680,N_11086);
xnor U12147 (N_12147,N_10207,N_11126);
nand U12148 (N_12148,N_10384,N_11230);
nand U12149 (N_12149,N_10525,N_10232);
nor U12150 (N_12150,N_10707,N_10064);
or U12151 (N_12151,N_10361,N_10103);
nand U12152 (N_12152,N_10421,N_10711);
xor U12153 (N_12153,N_10936,N_11196);
nand U12154 (N_12154,N_10676,N_10677);
and U12155 (N_12155,N_10022,N_10118);
nand U12156 (N_12156,N_11239,N_10632);
and U12157 (N_12157,N_11038,N_11098);
or U12158 (N_12158,N_10736,N_10182);
xnor U12159 (N_12159,N_10431,N_11161);
nor U12160 (N_12160,N_10043,N_10643);
and U12161 (N_12161,N_11091,N_10251);
nor U12162 (N_12162,N_10234,N_10687);
and U12163 (N_12163,N_10724,N_10174);
nor U12164 (N_12164,N_10941,N_11219);
and U12165 (N_12165,N_11171,N_10026);
nor U12166 (N_12166,N_10498,N_11197);
nor U12167 (N_12167,N_10506,N_10828);
nor U12168 (N_12168,N_10662,N_11199);
xnor U12169 (N_12169,N_11206,N_10916);
xor U12170 (N_12170,N_10110,N_10540);
and U12171 (N_12171,N_10332,N_10287);
and U12172 (N_12172,N_11130,N_10976);
nand U12173 (N_12173,N_10393,N_10119);
and U12174 (N_12174,N_10218,N_11033);
nand U12175 (N_12175,N_10882,N_10234);
or U12176 (N_12176,N_11052,N_11193);
or U12177 (N_12177,N_10386,N_10661);
nor U12178 (N_12178,N_10576,N_10004);
or U12179 (N_12179,N_10605,N_10700);
nand U12180 (N_12180,N_10722,N_10781);
or U12181 (N_12181,N_10653,N_10956);
or U12182 (N_12182,N_11145,N_11159);
nor U12183 (N_12183,N_10616,N_10072);
or U12184 (N_12184,N_10528,N_10210);
xor U12185 (N_12185,N_10153,N_10989);
nor U12186 (N_12186,N_10108,N_10395);
nor U12187 (N_12187,N_10401,N_10026);
nand U12188 (N_12188,N_10913,N_10442);
nand U12189 (N_12189,N_10690,N_10100);
nand U12190 (N_12190,N_11122,N_10317);
and U12191 (N_12191,N_10070,N_10991);
nand U12192 (N_12192,N_10189,N_10880);
and U12193 (N_12193,N_10012,N_10326);
xnor U12194 (N_12194,N_11226,N_10905);
nand U12195 (N_12195,N_10142,N_10963);
xnor U12196 (N_12196,N_11117,N_10678);
xnor U12197 (N_12197,N_10482,N_10934);
or U12198 (N_12198,N_10652,N_10055);
or U12199 (N_12199,N_10655,N_10588);
nor U12200 (N_12200,N_11002,N_10127);
xor U12201 (N_12201,N_10689,N_10176);
and U12202 (N_12202,N_10030,N_11186);
and U12203 (N_12203,N_10994,N_10894);
nor U12204 (N_12204,N_10697,N_10420);
xor U12205 (N_12205,N_11206,N_11044);
nor U12206 (N_12206,N_10477,N_10232);
xnor U12207 (N_12207,N_10281,N_10191);
nor U12208 (N_12208,N_10904,N_11033);
and U12209 (N_12209,N_10234,N_10859);
nor U12210 (N_12210,N_11155,N_11233);
and U12211 (N_12211,N_10628,N_10852);
nor U12212 (N_12212,N_10505,N_10525);
or U12213 (N_12213,N_10575,N_10641);
and U12214 (N_12214,N_10027,N_10916);
and U12215 (N_12215,N_10379,N_10285);
and U12216 (N_12216,N_10216,N_10493);
xnor U12217 (N_12217,N_10389,N_10934);
or U12218 (N_12218,N_10411,N_10951);
xnor U12219 (N_12219,N_10831,N_10206);
nor U12220 (N_12220,N_10227,N_10413);
nor U12221 (N_12221,N_10849,N_10178);
and U12222 (N_12222,N_10828,N_10721);
and U12223 (N_12223,N_10768,N_10078);
and U12224 (N_12224,N_10818,N_10980);
nor U12225 (N_12225,N_10808,N_10850);
nand U12226 (N_12226,N_10611,N_10258);
or U12227 (N_12227,N_10346,N_11192);
or U12228 (N_12228,N_11050,N_10012);
nor U12229 (N_12229,N_10936,N_10489);
and U12230 (N_12230,N_11206,N_10924);
xnor U12231 (N_12231,N_10381,N_10742);
and U12232 (N_12232,N_10309,N_10369);
xnor U12233 (N_12233,N_11076,N_10844);
or U12234 (N_12234,N_11027,N_10372);
and U12235 (N_12235,N_10423,N_10583);
xnor U12236 (N_12236,N_10943,N_11037);
nor U12237 (N_12237,N_10483,N_10816);
nand U12238 (N_12238,N_10229,N_10141);
nor U12239 (N_12239,N_10754,N_10478);
nand U12240 (N_12240,N_10206,N_10799);
nor U12241 (N_12241,N_11212,N_10669);
nand U12242 (N_12242,N_10202,N_11112);
and U12243 (N_12243,N_10831,N_11135);
and U12244 (N_12244,N_10246,N_10438);
and U12245 (N_12245,N_10817,N_10246);
nand U12246 (N_12246,N_10536,N_10682);
or U12247 (N_12247,N_11134,N_10306);
nor U12248 (N_12248,N_10410,N_10548);
or U12249 (N_12249,N_10205,N_10511);
or U12250 (N_12250,N_10307,N_11058);
or U12251 (N_12251,N_11132,N_10216);
or U12252 (N_12252,N_10638,N_10150);
or U12253 (N_12253,N_10150,N_11065);
nor U12254 (N_12254,N_10970,N_10850);
nor U12255 (N_12255,N_10213,N_10901);
or U12256 (N_12256,N_10587,N_10179);
xnor U12257 (N_12257,N_10980,N_10892);
or U12258 (N_12258,N_10692,N_11052);
xor U12259 (N_12259,N_11004,N_10739);
or U12260 (N_12260,N_10592,N_10490);
nor U12261 (N_12261,N_10531,N_10740);
and U12262 (N_12262,N_10881,N_10131);
nand U12263 (N_12263,N_10726,N_10683);
nand U12264 (N_12264,N_10631,N_11088);
xor U12265 (N_12265,N_10172,N_10408);
or U12266 (N_12266,N_10561,N_10178);
nand U12267 (N_12267,N_10808,N_10669);
nor U12268 (N_12268,N_10304,N_10496);
or U12269 (N_12269,N_10158,N_11016);
and U12270 (N_12270,N_10547,N_10461);
and U12271 (N_12271,N_10375,N_10700);
nor U12272 (N_12272,N_10423,N_10210);
or U12273 (N_12273,N_10571,N_10854);
nand U12274 (N_12274,N_11209,N_10070);
nand U12275 (N_12275,N_10266,N_10598);
xnor U12276 (N_12276,N_10438,N_10079);
xor U12277 (N_12277,N_11094,N_11159);
xnor U12278 (N_12278,N_10219,N_10268);
xnor U12279 (N_12279,N_10378,N_10870);
and U12280 (N_12280,N_10658,N_11036);
xnor U12281 (N_12281,N_10665,N_10286);
and U12282 (N_12282,N_11101,N_11027);
xnor U12283 (N_12283,N_10701,N_10406);
xnor U12284 (N_12284,N_10624,N_10685);
and U12285 (N_12285,N_10301,N_10669);
and U12286 (N_12286,N_10883,N_10466);
xor U12287 (N_12287,N_10509,N_10720);
xnor U12288 (N_12288,N_10288,N_10816);
and U12289 (N_12289,N_11168,N_11056);
or U12290 (N_12290,N_10464,N_10748);
nand U12291 (N_12291,N_10493,N_10336);
nor U12292 (N_12292,N_10628,N_10851);
and U12293 (N_12293,N_10489,N_10487);
xor U12294 (N_12294,N_11128,N_10366);
nor U12295 (N_12295,N_10486,N_10128);
or U12296 (N_12296,N_10638,N_10377);
and U12297 (N_12297,N_10786,N_10671);
nor U12298 (N_12298,N_10407,N_10757);
nand U12299 (N_12299,N_10099,N_11137);
and U12300 (N_12300,N_10047,N_11097);
nor U12301 (N_12301,N_10405,N_10575);
nor U12302 (N_12302,N_11056,N_10225);
nand U12303 (N_12303,N_10952,N_11235);
nor U12304 (N_12304,N_10884,N_10315);
and U12305 (N_12305,N_11118,N_10600);
nand U12306 (N_12306,N_10171,N_10115);
nor U12307 (N_12307,N_11090,N_11132);
and U12308 (N_12308,N_10066,N_10872);
and U12309 (N_12309,N_10289,N_11019);
or U12310 (N_12310,N_11194,N_10013);
or U12311 (N_12311,N_10920,N_10131);
or U12312 (N_12312,N_10175,N_11157);
nor U12313 (N_12313,N_11234,N_10479);
and U12314 (N_12314,N_10006,N_10921);
or U12315 (N_12315,N_10545,N_11243);
and U12316 (N_12316,N_10332,N_11208);
or U12317 (N_12317,N_10489,N_10070);
nand U12318 (N_12318,N_11169,N_10790);
or U12319 (N_12319,N_10661,N_10625);
nand U12320 (N_12320,N_10293,N_10579);
and U12321 (N_12321,N_11038,N_10768);
nand U12322 (N_12322,N_10282,N_10867);
or U12323 (N_12323,N_11071,N_10958);
nand U12324 (N_12324,N_10805,N_10396);
nor U12325 (N_12325,N_10575,N_10452);
nor U12326 (N_12326,N_10340,N_10230);
nor U12327 (N_12327,N_10139,N_10295);
nor U12328 (N_12328,N_10102,N_10184);
nor U12329 (N_12329,N_10514,N_10803);
nand U12330 (N_12330,N_11104,N_11199);
xor U12331 (N_12331,N_10101,N_10979);
and U12332 (N_12332,N_10044,N_10553);
or U12333 (N_12333,N_10389,N_10924);
xnor U12334 (N_12334,N_10502,N_11010);
or U12335 (N_12335,N_10708,N_10280);
and U12336 (N_12336,N_10438,N_10915);
xor U12337 (N_12337,N_11196,N_10779);
nand U12338 (N_12338,N_10002,N_11043);
xor U12339 (N_12339,N_10571,N_10799);
nor U12340 (N_12340,N_10870,N_10939);
or U12341 (N_12341,N_10958,N_10635);
xor U12342 (N_12342,N_10604,N_10775);
or U12343 (N_12343,N_10919,N_10088);
or U12344 (N_12344,N_10709,N_10938);
nand U12345 (N_12345,N_10198,N_10747);
or U12346 (N_12346,N_11078,N_10331);
nand U12347 (N_12347,N_11094,N_10415);
xor U12348 (N_12348,N_10586,N_10309);
or U12349 (N_12349,N_10231,N_10263);
xnor U12350 (N_12350,N_11240,N_11044);
nor U12351 (N_12351,N_10930,N_10807);
or U12352 (N_12352,N_10660,N_10875);
nand U12353 (N_12353,N_10697,N_10309);
nand U12354 (N_12354,N_10166,N_10027);
nand U12355 (N_12355,N_10925,N_10279);
xor U12356 (N_12356,N_10458,N_10930);
nor U12357 (N_12357,N_10904,N_10315);
nand U12358 (N_12358,N_10071,N_10637);
and U12359 (N_12359,N_10472,N_10979);
xor U12360 (N_12360,N_10309,N_11249);
or U12361 (N_12361,N_11009,N_11134);
xor U12362 (N_12362,N_10085,N_10068);
or U12363 (N_12363,N_10986,N_10265);
or U12364 (N_12364,N_10004,N_11049);
nor U12365 (N_12365,N_10564,N_10422);
and U12366 (N_12366,N_10469,N_10154);
nor U12367 (N_12367,N_11200,N_10287);
nor U12368 (N_12368,N_11217,N_10231);
or U12369 (N_12369,N_10348,N_10128);
and U12370 (N_12370,N_10301,N_10765);
xnor U12371 (N_12371,N_10641,N_10588);
nor U12372 (N_12372,N_10433,N_10472);
nor U12373 (N_12373,N_10459,N_10513);
or U12374 (N_12374,N_10184,N_10551);
nand U12375 (N_12375,N_10856,N_10364);
nand U12376 (N_12376,N_10912,N_11223);
nor U12377 (N_12377,N_10872,N_10272);
nand U12378 (N_12378,N_10402,N_10293);
nand U12379 (N_12379,N_10467,N_10313);
nand U12380 (N_12380,N_10824,N_11140);
xnor U12381 (N_12381,N_11175,N_10422);
nor U12382 (N_12382,N_11158,N_10559);
or U12383 (N_12383,N_10696,N_11031);
or U12384 (N_12384,N_10173,N_10560);
xor U12385 (N_12385,N_11160,N_11043);
or U12386 (N_12386,N_11063,N_10861);
and U12387 (N_12387,N_10396,N_10451);
nor U12388 (N_12388,N_10235,N_10722);
and U12389 (N_12389,N_10059,N_11171);
nand U12390 (N_12390,N_10680,N_10284);
nor U12391 (N_12391,N_10219,N_10848);
nor U12392 (N_12392,N_11026,N_10913);
nand U12393 (N_12393,N_10633,N_10489);
and U12394 (N_12394,N_11137,N_11136);
nor U12395 (N_12395,N_10549,N_10514);
nor U12396 (N_12396,N_10623,N_10435);
xnor U12397 (N_12397,N_10414,N_10509);
and U12398 (N_12398,N_10782,N_10144);
or U12399 (N_12399,N_11134,N_11203);
and U12400 (N_12400,N_10541,N_10728);
and U12401 (N_12401,N_10898,N_10327);
nor U12402 (N_12402,N_10105,N_10190);
nor U12403 (N_12403,N_10152,N_11000);
nand U12404 (N_12404,N_10690,N_10014);
nand U12405 (N_12405,N_10211,N_10419);
and U12406 (N_12406,N_10114,N_11014);
and U12407 (N_12407,N_10551,N_10732);
nor U12408 (N_12408,N_10257,N_11157);
and U12409 (N_12409,N_10403,N_10615);
nor U12410 (N_12410,N_10703,N_11026);
nand U12411 (N_12411,N_11146,N_11048);
and U12412 (N_12412,N_10435,N_10540);
nand U12413 (N_12413,N_10997,N_11180);
nand U12414 (N_12414,N_11162,N_10600);
nand U12415 (N_12415,N_11152,N_10196);
and U12416 (N_12416,N_10272,N_11129);
nand U12417 (N_12417,N_11080,N_10728);
nand U12418 (N_12418,N_10961,N_11093);
nand U12419 (N_12419,N_10064,N_10024);
and U12420 (N_12420,N_10536,N_10230);
and U12421 (N_12421,N_10029,N_11107);
xor U12422 (N_12422,N_10496,N_11035);
xnor U12423 (N_12423,N_10762,N_10207);
or U12424 (N_12424,N_10672,N_10007);
nor U12425 (N_12425,N_10733,N_11153);
or U12426 (N_12426,N_11034,N_11158);
or U12427 (N_12427,N_11038,N_10982);
xnor U12428 (N_12428,N_10088,N_10920);
nor U12429 (N_12429,N_10232,N_10451);
nor U12430 (N_12430,N_10636,N_10419);
xnor U12431 (N_12431,N_10377,N_10680);
and U12432 (N_12432,N_10369,N_10923);
nand U12433 (N_12433,N_10390,N_10871);
or U12434 (N_12434,N_10275,N_11170);
xor U12435 (N_12435,N_10294,N_10614);
nand U12436 (N_12436,N_10960,N_10236);
nand U12437 (N_12437,N_10293,N_10022);
xor U12438 (N_12438,N_10037,N_10555);
and U12439 (N_12439,N_10729,N_10423);
nor U12440 (N_12440,N_11045,N_10565);
or U12441 (N_12441,N_11188,N_10694);
or U12442 (N_12442,N_11224,N_10820);
nand U12443 (N_12443,N_10558,N_10578);
nand U12444 (N_12444,N_10888,N_10097);
nor U12445 (N_12445,N_10731,N_10935);
xnor U12446 (N_12446,N_11219,N_10341);
or U12447 (N_12447,N_10248,N_10847);
nor U12448 (N_12448,N_10316,N_10234);
nor U12449 (N_12449,N_11080,N_10269);
nor U12450 (N_12450,N_10149,N_11081);
nand U12451 (N_12451,N_10572,N_10710);
nand U12452 (N_12452,N_10190,N_10083);
nand U12453 (N_12453,N_10438,N_11080);
or U12454 (N_12454,N_10401,N_10950);
and U12455 (N_12455,N_10557,N_10616);
and U12456 (N_12456,N_10594,N_10058);
or U12457 (N_12457,N_10691,N_10036);
or U12458 (N_12458,N_10780,N_10472);
nand U12459 (N_12459,N_10727,N_10344);
xnor U12460 (N_12460,N_10597,N_10579);
xor U12461 (N_12461,N_11062,N_11132);
nor U12462 (N_12462,N_10456,N_10094);
xor U12463 (N_12463,N_10641,N_11194);
nor U12464 (N_12464,N_10990,N_10733);
nand U12465 (N_12465,N_10110,N_10752);
xor U12466 (N_12466,N_10662,N_11215);
nand U12467 (N_12467,N_11059,N_10190);
or U12468 (N_12468,N_11142,N_10721);
or U12469 (N_12469,N_10926,N_10359);
nor U12470 (N_12470,N_10560,N_11234);
nor U12471 (N_12471,N_10629,N_10628);
and U12472 (N_12472,N_10879,N_10888);
xor U12473 (N_12473,N_10340,N_10821);
or U12474 (N_12474,N_10158,N_10407);
nand U12475 (N_12475,N_10086,N_10680);
nor U12476 (N_12476,N_10814,N_10213);
or U12477 (N_12477,N_11052,N_10887);
nand U12478 (N_12478,N_10818,N_10333);
and U12479 (N_12479,N_10378,N_11232);
nor U12480 (N_12480,N_10151,N_10128);
xor U12481 (N_12481,N_10437,N_10533);
nor U12482 (N_12482,N_10951,N_10130);
nand U12483 (N_12483,N_10588,N_10704);
xnor U12484 (N_12484,N_10606,N_10847);
nor U12485 (N_12485,N_11084,N_10487);
and U12486 (N_12486,N_10235,N_10294);
or U12487 (N_12487,N_10869,N_10366);
xnor U12488 (N_12488,N_10706,N_10750);
and U12489 (N_12489,N_10563,N_10275);
and U12490 (N_12490,N_10635,N_10722);
xnor U12491 (N_12491,N_10369,N_11119);
nor U12492 (N_12492,N_10339,N_10226);
nand U12493 (N_12493,N_10187,N_10891);
nand U12494 (N_12494,N_10993,N_10246);
nor U12495 (N_12495,N_10162,N_11176);
xnor U12496 (N_12496,N_10472,N_10579);
xor U12497 (N_12497,N_11068,N_11212);
or U12498 (N_12498,N_10213,N_11007);
xor U12499 (N_12499,N_10585,N_10622);
xnor U12500 (N_12500,N_12457,N_11264);
or U12501 (N_12501,N_12013,N_12453);
nor U12502 (N_12502,N_11369,N_11373);
nand U12503 (N_12503,N_12159,N_11402);
or U12504 (N_12504,N_12354,N_12221);
nand U12505 (N_12505,N_11468,N_12071);
and U12506 (N_12506,N_11571,N_12399);
nand U12507 (N_12507,N_12017,N_12476);
or U12508 (N_12508,N_11882,N_11986);
nand U12509 (N_12509,N_11613,N_12056);
xor U12510 (N_12510,N_11660,N_12258);
nand U12511 (N_12511,N_11721,N_11367);
nor U12512 (N_12512,N_12194,N_12295);
nand U12513 (N_12513,N_11553,N_12424);
nand U12514 (N_12514,N_12038,N_12143);
xnor U12515 (N_12515,N_11623,N_11636);
or U12516 (N_12516,N_12296,N_12185);
nor U12517 (N_12517,N_12487,N_12462);
xnor U12518 (N_12518,N_11634,N_11513);
and U12519 (N_12519,N_11730,N_11763);
nor U12520 (N_12520,N_12379,N_12235);
nand U12521 (N_12521,N_11315,N_12483);
nand U12522 (N_12522,N_11698,N_12035);
nor U12523 (N_12523,N_12302,N_11655);
nor U12524 (N_12524,N_11479,N_11328);
nand U12525 (N_12525,N_11612,N_11699);
or U12526 (N_12526,N_11538,N_11288);
nor U12527 (N_12527,N_11833,N_11378);
nor U12528 (N_12528,N_12468,N_12313);
nand U12529 (N_12529,N_12232,N_11706);
nand U12530 (N_12530,N_11371,N_12492);
xnor U12531 (N_12531,N_12073,N_12496);
nor U12532 (N_12532,N_12198,N_12342);
xor U12533 (N_12533,N_11311,N_11361);
nand U12534 (N_12534,N_11967,N_12175);
xor U12535 (N_12535,N_12050,N_11608);
nor U12536 (N_12536,N_12270,N_11422);
and U12537 (N_12537,N_11950,N_11823);
or U12538 (N_12538,N_11801,N_11624);
nand U12539 (N_12539,N_11802,N_11459);
and U12540 (N_12540,N_11509,N_12361);
or U12541 (N_12541,N_11320,N_11670);
xor U12542 (N_12542,N_11971,N_11872);
nand U12543 (N_12543,N_11521,N_11598);
nand U12544 (N_12544,N_12455,N_12331);
nor U12545 (N_12545,N_12176,N_11300);
and U12546 (N_12546,N_11905,N_11672);
xor U12547 (N_12547,N_11541,N_11516);
nand U12548 (N_12548,N_11886,N_11847);
nand U12549 (N_12549,N_11430,N_12420);
xor U12550 (N_12550,N_12266,N_11867);
or U12551 (N_12551,N_12172,N_11734);
and U12552 (N_12552,N_11291,N_11930);
nor U12553 (N_12553,N_11473,N_11250);
nor U12554 (N_12554,N_11309,N_11918);
nor U12555 (N_12555,N_11267,N_11354);
xnor U12556 (N_12556,N_12392,N_11476);
or U12557 (N_12557,N_11704,N_12099);
nor U12558 (N_12558,N_11737,N_11607);
or U12559 (N_12559,N_11832,N_12314);
nor U12560 (N_12560,N_12243,N_11983);
or U12561 (N_12561,N_11390,N_11920);
xor U12562 (N_12562,N_12464,N_11335);
xor U12563 (N_12563,N_11331,N_12223);
and U12564 (N_12564,N_11396,N_12166);
xor U12565 (N_12565,N_12054,N_11449);
nor U12566 (N_12566,N_11962,N_12103);
nor U12567 (N_12567,N_11979,N_11363);
xor U12568 (N_12568,N_11880,N_11626);
xor U12569 (N_12569,N_12061,N_11691);
or U12570 (N_12570,N_11951,N_11263);
nand U12571 (N_12571,N_11419,N_12162);
and U12572 (N_12572,N_11888,N_11965);
nor U12573 (N_12573,N_12454,N_12240);
and U12574 (N_12574,N_12131,N_12092);
nor U12575 (N_12575,N_12350,N_12432);
nand U12576 (N_12576,N_11646,N_12231);
or U12577 (N_12577,N_12308,N_11532);
nand U12578 (N_12578,N_12470,N_11540);
nand U12579 (N_12579,N_12316,N_12422);
or U12580 (N_12580,N_11506,N_11450);
xnor U12581 (N_12581,N_11330,N_11701);
or U12582 (N_12582,N_12477,N_12493);
nand U12583 (N_12583,N_11425,N_11527);
and U12584 (N_12584,N_12499,N_12444);
xnor U12585 (N_12585,N_11935,N_12052);
or U12586 (N_12586,N_11818,N_12337);
nor U12587 (N_12587,N_11929,N_12100);
xnor U12588 (N_12588,N_12059,N_11819);
and U12589 (N_12589,N_11340,N_12309);
xnor U12590 (N_12590,N_12006,N_12480);
xor U12591 (N_12591,N_12352,N_11878);
and U12592 (N_12592,N_12484,N_12135);
or U12593 (N_12593,N_12441,N_11671);
nand U12594 (N_12594,N_11939,N_12149);
xor U12595 (N_12595,N_11972,N_11658);
nor U12596 (N_12596,N_11941,N_12426);
nand U12597 (N_12597,N_12490,N_11418);
or U12598 (N_12598,N_11739,N_11545);
xnor U12599 (N_12599,N_11649,N_11280);
xor U12600 (N_12600,N_12207,N_11585);
and U12601 (N_12601,N_12163,N_11502);
xor U12602 (N_12602,N_11394,N_11455);
nand U12603 (N_12603,N_11831,N_12395);
xnor U12604 (N_12604,N_11495,N_11314);
and U12605 (N_12605,N_11544,N_11357);
nor U12606 (N_12606,N_11915,N_12319);
or U12607 (N_12607,N_11557,N_11548);
xnor U12608 (N_12608,N_12069,N_11728);
nand U12609 (N_12609,N_11835,N_11994);
and U12610 (N_12610,N_12153,N_11355);
and U12611 (N_12611,N_12126,N_12091);
or U12612 (N_12612,N_11253,N_11407);
xor U12613 (N_12613,N_12030,N_11324);
nor U12614 (N_12614,N_11955,N_11411);
and U12615 (N_12615,N_12081,N_11834);
nand U12616 (N_12616,N_11817,N_11445);
xnor U12617 (N_12617,N_12344,N_11283);
or U12618 (N_12618,N_11559,N_12357);
or U12619 (N_12619,N_11707,N_11630);
and U12620 (N_12620,N_12307,N_11305);
and U12621 (N_12621,N_11567,N_12396);
nor U12622 (N_12622,N_11849,N_11260);
xnor U12623 (N_12623,N_11491,N_11720);
xnor U12624 (N_12624,N_12388,N_12239);
and U12625 (N_12625,N_12467,N_12274);
nor U12626 (N_12626,N_12459,N_11617);
xor U12627 (N_12627,N_11751,N_12475);
nand U12628 (N_12628,N_11265,N_12315);
or U12629 (N_12629,N_12471,N_11599);
or U12630 (N_12630,N_11957,N_12401);
or U12631 (N_12631,N_11470,N_12353);
and U12632 (N_12632,N_11710,N_12409);
or U12633 (N_12633,N_12443,N_11807);
and U12634 (N_12634,N_11583,N_12024);
nand U12635 (N_12635,N_11257,N_12021);
nand U12636 (N_12636,N_11622,N_11657);
nor U12637 (N_12637,N_12387,N_12124);
and U12638 (N_12638,N_11687,N_12288);
or U12639 (N_12639,N_12064,N_12275);
or U12640 (N_12640,N_11290,N_11385);
xor U12641 (N_12641,N_11594,N_11959);
and U12642 (N_12642,N_12322,N_11753);
nor U12643 (N_12643,N_12215,N_12283);
nor U12644 (N_12644,N_12226,N_12062);
nand U12645 (N_12645,N_11754,N_11944);
nand U12646 (N_12646,N_11727,N_11619);
xor U12647 (N_12647,N_12220,N_11947);
and U12648 (N_12648,N_12106,N_11813);
nor U12649 (N_12649,N_12097,N_11282);
nor U12650 (N_12650,N_11362,N_12276);
xor U12651 (N_12651,N_11399,N_12389);
xor U12652 (N_12652,N_12386,N_11916);
and U12653 (N_12653,N_12053,N_11684);
or U12654 (N_12654,N_11996,N_12028);
xor U12655 (N_12655,N_12112,N_11816);
or U12656 (N_12656,N_11934,N_11978);
and U12657 (N_12657,N_12261,N_12347);
and U12658 (N_12658,N_11474,N_11436);
or U12659 (N_12659,N_12320,N_12324);
nand U12660 (N_12660,N_11365,N_11884);
nor U12661 (N_12661,N_11252,N_12268);
nand U12662 (N_12662,N_11457,N_11960);
xor U12663 (N_12663,N_11803,N_11744);
nor U12664 (N_12664,N_12078,N_11862);
xnor U12665 (N_12665,N_12383,N_11787);
nand U12666 (N_12666,N_11377,N_11524);
nand U12667 (N_12667,N_11987,N_11830);
nor U12668 (N_12668,N_11379,N_11633);
nand U12669 (N_12669,N_12249,N_11881);
xnor U12670 (N_12670,N_12070,N_12299);
nand U12671 (N_12671,N_12425,N_12148);
nand U12672 (N_12672,N_11278,N_12391);
and U12673 (N_12673,N_12278,N_12244);
nand U12674 (N_12674,N_11759,N_11773);
or U12675 (N_12675,N_11562,N_12290);
nand U12676 (N_12676,N_11820,N_11907);
and U12677 (N_12677,N_12257,N_12216);
or U12678 (N_12678,N_12005,N_11580);
nor U12679 (N_12679,N_12193,N_12170);
xnor U12680 (N_12680,N_12087,N_12248);
and U12681 (N_12681,N_12079,N_11417);
xor U12682 (N_12682,N_11554,N_12406);
and U12683 (N_12683,N_11376,N_12136);
and U12684 (N_12684,N_11799,N_12115);
or U12685 (N_12685,N_11480,N_11713);
or U12686 (N_12686,N_11866,N_11871);
nand U12687 (N_12687,N_12356,N_12177);
xnor U12688 (N_12688,N_11964,N_11453);
xnor U12689 (N_12689,N_12210,N_12074);
or U12690 (N_12690,N_11403,N_12104);
nand U12691 (N_12691,N_12109,N_11952);
nand U12692 (N_12692,N_11785,N_11946);
and U12693 (N_12693,N_12430,N_11368);
xor U12694 (N_12694,N_11500,N_11327);
or U12695 (N_12695,N_11464,N_11772);
or U12696 (N_12696,N_12362,N_11752);
and U12697 (N_12697,N_11384,N_11621);
or U12698 (N_12698,N_11561,N_11606);
nand U12699 (N_12699,N_11990,N_12417);
xnor U12700 (N_12700,N_11398,N_11645);
or U12701 (N_12701,N_11579,N_12334);
nor U12702 (N_12702,N_12125,N_11931);
or U12703 (N_12703,N_11597,N_11928);
xnor U12704 (N_12704,N_11281,N_11405);
nor U12705 (N_12705,N_11779,N_11269);
and U12706 (N_12706,N_11894,N_11841);
and U12707 (N_12707,N_12128,N_11413);
or U12708 (N_12708,N_11589,N_12330);
nand U12709 (N_12709,N_12310,N_11575);
xnor U12710 (N_12710,N_12394,N_12118);
nand U12711 (N_12711,N_11942,N_11356);
and U12712 (N_12712,N_11504,N_12123);
nor U12713 (N_12713,N_11348,N_11522);
nand U12714 (N_12714,N_12042,N_11338);
and U12715 (N_12715,N_12019,N_11614);
xnor U12716 (N_12716,N_11973,N_12335);
or U12717 (N_12717,N_11656,N_11953);
xor U12718 (N_12718,N_11761,N_11879);
xor U12719 (N_12719,N_11900,N_11556);
xnor U12720 (N_12720,N_12068,N_11899);
nand U12721 (N_12721,N_11302,N_12084);
or U12722 (N_12722,N_12340,N_12398);
or U12723 (N_12723,N_11981,N_12433);
and U12724 (N_12724,N_11381,N_12152);
xnor U12725 (N_12725,N_11673,N_12156);
nor U12726 (N_12726,N_11452,N_11668);
or U12727 (N_12727,N_11366,N_11471);
and U12728 (N_12728,N_11873,N_11956);
and U12729 (N_12729,N_12348,N_11789);
and U12730 (N_12730,N_11653,N_12375);
and U12731 (N_12731,N_11401,N_12206);
and U12732 (N_12732,N_12098,N_12138);
or U12733 (N_12733,N_11272,N_12498);
and U12734 (N_12734,N_12345,N_11296);
or U12735 (N_12735,N_11814,N_12481);
nand U12736 (N_12736,N_11889,N_11898);
and U12737 (N_12737,N_11826,N_11937);
nand U12738 (N_12738,N_12113,N_12486);
or U12739 (N_12739,N_12045,N_11908);
xnor U12740 (N_12740,N_12048,N_12102);
nor U12741 (N_12741,N_11836,N_11319);
nor U12742 (N_12742,N_11654,N_11462);
nand U12743 (N_12743,N_11484,N_12402);
or U12744 (N_12744,N_11891,N_11736);
nor U12745 (N_12745,N_11518,N_12479);
nor U12746 (N_12746,N_12051,N_11729);
xor U12747 (N_12747,N_12305,N_11805);
or U12748 (N_12748,N_12328,N_11812);
nand U12749 (N_12749,N_11708,N_11749);
xor U12750 (N_12750,N_12411,N_12437);
xnor U12751 (N_12751,N_12197,N_12405);
nand U12752 (N_12752,N_11321,N_11463);
xor U12753 (N_12753,N_11828,N_11664);
nand U12754 (N_12754,N_11925,N_11611);
and U12755 (N_12755,N_11375,N_11844);
xnor U12756 (N_12756,N_11578,N_11932);
nand U12757 (N_12757,N_12196,N_12026);
and U12758 (N_12758,N_11352,N_11897);
or U12759 (N_12759,N_12174,N_11682);
or U12760 (N_12760,N_11917,N_12036);
xnor U12761 (N_12761,N_11991,N_11725);
or U12762 (N_12762,N_11688,N_12183);
xnor U12763 (N_12763,N_11793,N_12082);
and U12764 (N_12764,N_12397,N_11782);
and U12765 (N_12765,N_12473,N_11927);
or U12766 (N_12766,N_11912,N_11475);
xnor U12767 (N_12767,N_11251,N_12141);
nor U12768 (N_12768,N_11359,N_11890);
nand U12769 (N_12769,N_12456,N_11409);
or U12770 (N_12770,N_11806,N_12241);
xor U12771 (N_12771,N_12321,N_11317);
xnor U12772 (N_12772,N_11685,N_12349);
nor U12773 (N_12773,N_11514,N_11313);
xor U12774 (N_12774,N_11859,N_11926);
nand U12775 (N_12775,N_12063,N_11530);
or U12776 (N_12776,N_12450,N_11854);
and U12777 (N_12777,N_11883,N_11428);
and U12778 (N_12778,N_12090,N_11326);
or U12779 (N_12779,N_11631,N_11998);
nand U12780 (N_12780,N_12372,N_11546);
or U12781 (N_12781,N_11702,N_12360);
nor U12782 (N_12782,N_12368,N_12238);
and U12783 (N_12783,N_11298,N_11542);
or U12784 (N_12784,N_11286,N_12023);
and U12785 (N_12785,N_11681,N_12117);
or U12786 (N_12786,N_11601,N_12014);
and U12787 (N_12787,N_11712,N_11602);
xor U12788 (N_12788,N_11954,N_12482);
nand U12789 (N_12789,N_11757,N_12000);
or U12790 (N_12790,N_11770,N_11731);
and U12791 (N_12791,N_11345,N_11896);
and U12792 (N_12792,N_12363,N_11639);
nand U12793 (N_12793,N_11781,N_11489);
or U12794 (N_12794,N_11266,N_11439);
nand U12795 (N_12795,N_11458,N_12008);
xnor U12796 (N_12796,N_11690,N_12385);
xor U12797 (N_12797,N_11662,N_11674);
or U12798 (N_12798,N_11337,N_12204);
or U12799 (N_12799,N_12250,N_11570);
nor U12800 (N_12800,N_11349,N_11582);
or U12801 (N_12801,N_11414,N_11400);
or U12802 (N_12802,N_12466,N_12093);
nor U12803 (N_12803,N_11270,N_11910);
and U12804 (N_12804,N_12116,N_12129);
nand U12805 (N_12805,N_11625,N_11408);
or U12806 (N_12806,N_11842,N_11755);
and U12807 (N_12807,N_11395,N_11472);
nor U12808 (N_12808,N_11564,N_12242);
nand U12809 (N_12809,N_11988,N_11767);
nand U12810 (N_12810,N_12246,N_11496);
nor U12811 (N_12811,N_12155,N_12080);
xnor U12812 (N_12812,N_12173,N_12209);
or U12813 (N_12813,N_11709,N_12157);
or U12814 (N_12814,N_12323,N_11507);
and U12815 (N_12815,N_11304,N_11444);
and U12816 (N_12816,N_12291,N_12474);
and U12817 (N_12817,N_12111,N_12140);
and U12818 (N_12818,N_11794,N_12269);
nand U12819 (N_12819,N_11256,N_12076);
and U12820 (N_12820,N_11745,N_11482);
nor U12821 (N_12821,N_12094,N_11437);
and U12822 (N_12822,N_11632,N_11969);
or U12823 (N_12823,N_11650,N_11858);
and U12824 (N_12824,N_11483,N_11719);
and U12825 (N_12825,N_12077,N_12224);
nor U12826 (N_12826,N_12469,N_12317);
nand U12827 (N_12827,N_11467,N_11914);
or U12828 (N_12828,N_12001,N_11603);
nor U12829 (N_12829,N_11863,N_11995);
or U12830 (N_12830,N_11762,N_11647);
and U12831 (N_12831,N_11528,N_11857);
xor U12832 (N_12832,N_12066,N_11764);
xor U12833 (N_12833,N_11543,N_11689);
or U12834 (N_12834,N_11526,N_12214);
xor U12835 (N_12835,N_11776,N_11353);
nor U12836 (N_12836,N_11984,N_11628);
nor U12837 (N_12837,N_11895,N_12010);
nand U12838 (N_12838,N_12095,N_12413);
xnor U12839 (N_12839,N_12228,N_12438);
xnor U12840 (N_12840,N_11887,N_11663);
and U12841 (N_12841,N_11271,N_11275);
nand U12842 (N_12842,N_11620,N_12089);
or U12843 (N_12843,N_11609,N_12286);
xnor U12844 (N_12844,N_12312,N_11748);
xor U12845 (N_12845,N_12018,N_11434);
or U12846 (N_12846,N_11446,N_12370);
nor U12847 (N_12847,N_11694,N_11966);
or U12848 (N_12848,N_12447,N_12083);
and U12849 (N_12849,N_11312,N_12255);
and U12850 (N_12850,N_11547,N_11629);
xnor U12851 (N_12851,N_11566,N_12127);
nor U12852 (N_12852,N_11961,N_11261);
nand U12853 (N_12853,N_11572,N_12096);
and U12854 (N_12854,N_11768,N_12440);
nand U12855 (N_12855,N_11989,N_11693);
nand U12856 (N_12856,N_11431,N_12415);
or U12857 (N_12857,N_11716,N_11865);
nand U12858 (N_12858,N_12364,N_12343);
or U12859 (N_12859,N_12376,N_11374);
xnor U12860 (N_12860,N_11740,N_12303);
nor U12861 (N_12861,N_12145,N_12192);
nor U12862 (N_12862,N_12213,N_11534);
or U12863 (N_12863,N_12142,N_11397);
nor U12864 (N_12864,N_11676,N_11922);
xnor U12865 (N_12865,N_11974,N_12040);
nand U12866 (N_12866,N_12154,N_12212);
and U12867 (N_12867,N_12289,N_12245);
xnor U12868 (N_12868,N_12107,N_11977);
and U12869 (N_12869,N_11587,N_11892);
and U12870 (N_12870,N_11638,N_11700);
xor U12871 (N_12871,N_12043,N_12182);
nand U12872 (N_12872,N_11339,N_11536);
or U12873 (N_12873,N_11387,N_11301);
xor U12874 (N_12874,N_12461,N_11565);
xor U12875 (N_12875,N_11466,N_12373);
or U12876 (N_12876,N_12122,N_11771);
or U12877 (N_12877,N_11370,N_12448);
nor U12878 (N_12878,N_11860,N_11796);
xor U12879 (N_12879,N_11618,N_11490);
or U12880 (N_12880,N_11287,N_12439);
nand U12881 (N_12881,N_11276,N_11515);
xor U12882 (N_12882,N_11864,N_12004);
nand U12883 (N_12883,N_11268,N_12429);
xor U12884 (N_12884,N_11550,N_12199);
nand U12885 (N_12885,N_12287,N_11393);
or U12886 (N_12886,N_12404,N_11277);
nand U12887 (N_12887,N_11577,N_12032);
nor U12888 (N_12888,N_11552,N_11294);
xor U12889 (N_12889,N_11284,N_12445);
nand U12890 (N_12890,N_11877,N_12072);
and U12891 (N_12891,N_11350,N_12171);
and U12892 (N_12892,N_11869,N_11677);
nor U12893 (N_12893,N_11307,N_12012);
xor U12894 (N_12894,N_12279,N_11809);
or U12895 (N_12895,N_11870,N_11695);
or U12896 (N_12896,N_11938,N_11503);
or U12897 (N_12897,N_11798,N_11850);
nand U12898 (N_12898,N_11590,N_11593);
or U12899 (N_12899,N_11837,N_12367);
and U12900 (N_12900,N_12284,N_12222);
or U12901 (N_12901,N_11643,N_11913);
nor U12902 (N_12902,N_12263,N_11641);
xor U12903 (N_12903,N_11853,N_11600);
nand U12904 (N_12904,N_12460,N_12400);
nor U12905 (N_12905,N_11711,N_12449);
or U12906 (N_12906,N_12346,N_11999);
xor U12907 (N_12907,N_11610,N_12421);
xnor U12908 (N_12908,N_11845,N_11410);
xnor U12909 (N_12909,N_11923,N_11644);
xor U12910 (N_12910,N_11911,N_11318);
xnor U12911 (N_12911,N_12229,N_11992);
xnor U12912 (N_12912,N_12325,N_11874);
or U12913 (N_12913,N_12416,N_12234);
nor U12914 (N_12914,N_11786,N_12306);
nor U12915 (N_12915,N_12427,N_11465);
nand U12916 (N_12916,N_12336,N_12139);
nand U12917 (N_12917,N_12495,N_11921);
nand U12918 (N_12918,N_12189,N_11511);
or U12919 (N_12919,N_11380,N_11940);
or U12920 (N_12920,N_12446,N_11438);
nand U12921 (N_12921,N_11783,N_11642);
or U12922 (N_12922,N_11306,N_11460);
nand U12923 (N_12923,N_12119,N_12463);
and U12924 (N_12924,N_11274,N_11824);
xnor U12925 (N_12925,N_12442,N_11519);
nor U12926 (N_12926,N_12219,N_11469);
nor U12927 (N_12927,N_11325,N_12164);
xor U12928 (N_12928,N_12179,N_12132);
xor U12929 (N_12929,N_11415,N_12205);
xnor U12930 (N_12930,N_12202,N_11584);
nand U12931 (N_12931,N_11510,N_12034);
nor U12932 (N_12932,N_11456,N_11481);
nor U12933 (N_12933,N_12300,N_11343);
nand U12934 (N_12934,N_11963,N_11715);
xor U12935 (N_12935,N_12494,N_12451);
nor U12936 (N_12936,N_11581,N_12489);
xnor U12937 (N_12937,N_12434,N_11316);
xnor U12938 (N_12938,N_11383,N_11722);
nand U12939 (N_12939,N_11520,N_12031);
xnor U12940 (N_12940,N_12150,N_11665);
nor U12941 (N_12941,N_12169,N_11427);
and U12942 (N_12942,N_11323,N_11958);
nand U12943 (N_12943,N_11821,N_11651);
nand U12944 (N_12944,N_12025,N_12203);
nand U12945 (N_12945,N_11846,N_12264);
or U12946 (N_12946,N_11588,N_12191);
nand U12947 (N_12947,N_12338,N_11735);
nand U12948 (N_12948,N_11738,N_11448);
or U12949 (N_12949,N_12247,N_11637);
and U12950 (N_12950,N_12058,N_11478);
nand U12951 (N_12951,N_12297,N_11827);
nand U12952 (N_12952,N_11903,N_11346);
or U12953 (N_12953,N_12165,N_12130);
nor U12954 (N_12954,N_11443,N_12168);
nand U12955 (N_12955,N_11856,N_12254);
nor U12956 (N_12956,N_11441,N_11531);
nor U12957 (N_12957,N_11750,N_12160);
nand U12958 (N_12958,N_11297,N_12146);
nand U12959 (N_12959,N_11901,N_11303);
or U12960 (N_12960,N_11774,N_12151);
nor U12961 (N_12961,N_11948,N_11822);
or U12962 (N_12962,N_11993,N_11741);
xor U12963 (N_12963,N_11810,N_12272);
nor U12964 (N_12964,N_11539,N_12178);
and U12965 (N_12965,N_12252,N_12039);
xnor U12966 (N_12966,N_12412,N_12282);
or U12967 (N_12967,N_11497,N_12259);
nand U12968 (N_12968,N_12253,N_11537);
nor U12969 (N_12969,N_11906,N_11364);
and U12970 (N_12970,N_12158,N_11840);
or U12971 (N_12971,N_12225,N_12002);
xor U12972 (N_12972,N_12384,N_11360);
xor U12973 (N_12973,N_12351,N_11555);
nand U12974 (N_12974,N_12418,N_11997);
nand U12975 (N_12975,N_11604,N_12120);
nor U12976 (N_12976,N_11791,N_12237);
and U12977 (N_12977,N_12359,N_11299);
nor U12978 (N_12978,N_12293,N_11429);
or U12979 (N_12979,N_12301,N_12472);
xor U12980 (N_12980,N_11747,N_11800);
and U12981 (N_12981,N_11766,N_12497);
and U12982 (N_12982,N_11902,N_11667);
xor U12983 (N_12983,N_12047,N_11838);
nor U12984 (N_12984,N_12333,N_11332);
or U12985 (N_12985,N_11568,N_11498);
xor U12986 (N_12986,N_12267,N_11295);
nor U12987 (N_12987,N_11372,N_12167);
nand U12988 (N_12988,N_12108,N_12251);
or U12989 (N_12989,N_11758,N_11705);
xor U12990 (N_12990,N_11388,N_11815);
and U12991 (N_12991,N_11652,N_11924);
nand U12992 (N_12992,N_11875,N_12184);
and U12993 (N_12993,N_11732,N_11627);
nor U12994 (N_12994,N_11679,N_11392);
and U12995 (N_12995,N_11985,N_11683);
nand U12996 (N_12996,N_12410,N_11616);
or U12997 (N_12997,N_11461,N_11592);
or U12998 (N_12998,N_11477,N_11718);
or U12999 (N_12999,N_11742,N_11943);
xnor U13000 (N_13000,N_11851,N_11426);
nand U13001 (N_13001,N_11535,N_12371);
xnor U13002 (N_13002,N_12067,N_12060);
or U13003 (N_13003,N_11386,N_12265);
xnor U13004 (N_13004,N_12478,N_11666);
xor U13005 (N_13005,N_11760,N_11726);
nor U13006 (N_13006,N_12009,N_11795);
or U13007 (N_13007,N_11308,N_12408);
and U13008 (N_13008,N_11868,N_11790);
or U13009 (N_13009,N_11336,N_11696);
nor U13010 (N_13010,N_12435,N_12431);
nand U13011 (N_13011,N_11255,N_11358);
xor U13012 (N_13012,N_11788,N_12181);
or U13013 (N_13013,N_11640,N_12022);
xnor U13014 (N_13014,N_11433,N_11591);
nor U13015 (N_13015,N_11848,N_12374);
nand U13016 (N_13016,N_12318,N_11382);
or U13017 (N_13017,N_11292,N_11804);
nor U13018 (N_13018,N_12236,N_11784);
nor U13019 (N_13019,N_12285,N_11505);
or U13020 (N_13020,N_12369,N_11733);
xor U13021 (N_13021,N_11508,N_12211);
nand U13022 (N_13022,N_11855,N_12085);
and U13023 (N_13023,N_11797,N_12365);
or U13024 (N_13024,N_12044,N_11949);
or U13025 (N_13025,N_11416,N_11825);
or U13026 (N_13026,N_12137,N_12329);
xor U13027 (N_13027,N_12208,N_12262);
xor U13028 (N_13028,N_11697,N_11447);
and U13029 (N_13029,N_12485,N_11549);
xnor U13030 (N_13030,N_11533,N_11852);
or U13031 (N_13031,N_11723,N_12147);
or U13032 (N_13032,N_11945,N_12055);
xor U13033 (N_13033,N_12110,N_12121);
and U13034 (N_13034,N_12088,N_11391);
or U13035 (N_13035,N_12218,N_11829);
xnor U13036 (N_13036,N_12188,N_12003);
xnor U13037 (N_13037,N_12027,N_11499);
or U13038 (N_13038,N_11342,N_11765);
nand U13039 (N_13039,N_12015,N_11780);
nand U13040 (N_13040,N_11605,N_12230);
xor U13041 (N_13041,N_12260,N_11976);
and U13042 (N_13042,N_11904,N_12407);
or U13043 (N_13043,N_12271,N_11493);
or U13044 (N_13044,N_12114,N_11279);
xor U13045 (N_13045,N_12101,N_11254);
or U13046 (N_13046,N_11258,N_12458);
nor U13047 (N_13047,N_11485,N_11440);
or U13048 (N_13048,N_11406,N_11285);
xor U13049 (N_13049,N_11980,N_11322);
or U13050 (N_13050,N_12280,N_11273);
nand U13051 (N_13051,N_11347,N_11344);
nor U13052 (N_13052,N_11678,N_11451);
nand U13053 (N_13053,N_12011,N_12033);
or U13054 (N_13054,N_11919,N_11576);
or U13055 (N_13055,N_11686,N_12326);
nor U13056 (N_13056,N_12393,N_12133);
or U13057 (N_13057,N_12273,N_12381);
nand U13058 (N_13058,N_12355,N_11421);
and U13059 (N_13059,N_11777,N_12403);
xor U13060 (N_13060,N_11778,N_12341);
and U13061 (N_13061,N_11586,N_12377);
nor U13062 (N_13062,N_11635,N_11669);
xnor U13063 (N_13063,N_12488,N_11724);
nor U13064 (N_13064,N_11423,N_11714);
or U13065 (N_13065,N_11341,N_11792);
and U13066 (N_13066,N_11389,N_11661);
nand U13067 (N_13067,N_11412,N_11648);
or U13068 (N_13068,N_12201,N_12390);
or U13069 (N_13069,N_12075,N_11775);
or U13070 (N_13070,N_11743,N_11432);
nor U13071 (N_13071,N_11936,N_11909);
nor U13072 (N_13072,N_11529,N_11970);
nor U13073 (N_13073,N_12436,N_11501);
and U13074 (N_13074,N_12298,N_11861);
xor U13075 (N_13075,N_11487,N_12292);
nand U13076 (N_13076,N_12195,N_12180);
or U13077 (N_13077,N_11523,N_12378);
and U13078 (N_13078,N_12049,N_12144);
or U13079 (N_13079,N_11486,N_12465);
or U13080 (N_13080,N_11675,N_11659);
and U13081 (N_13081,N_12065,N_11596);
xnor U13082 (N_13082,N_12294,N_11262);
xnor U13083 (N_13083,N_12161,N_11769);
xor U13084 (N_13084,N_12233,N_11494);
nor U13085 (N_13085,N_11843,N_12332);
nand U13086 (N_13086,N_11488,N_11259);
and U13087 (N_13087,N_11558,N_11680);
or U13088 (N_13088,N_11756,N_11424);
xor U13089 (N_13089,N_11492,N_11975);
nor U13090 (N_13090,N_12414,N_11717);
xor U13091 (N_13091,N_12227,N_11310);
or U13092 (N_13092,N_11435,N_11351);
or U13093 (N_13093,N_11329,N_11808);
nor U13094 (N_13094,N_11293,N_11811);
and U13095 (N_13095,N_12311,N_12366);
xnor U13096 (N_13096,N_12491,N_12304);
or U13097 (N_13097,N_12256,N_12380);
nand U13098 (N_13098,N_12217,N_12186);
xnor U13099 (N_13099,N_11334,N_12277);
or U13100 (N_13100,N_11876,N_12041);
nor U13101 (N_13101,N_11333,N_12428);
nor U13102 (N_13102,N_12007,N_11289);
nand U13103 (N_13103,N_12281,N_12105);
xor U13104 (N_13104,N_12046,N_12327);
xor U13105 (N_13105,N_11703,N_11982);
or U13106 (N_13106,N_12358,N_11893);
nor U13107 (N_13107,N_12187,N_12339);
nor U13108 (N_13108,N_12134,N_12452);
xor U13109 (N_13109,N_12419,N_11563);
and U13110 (N_13110,N_11595,N_12382);
nor U13111 (N_13111,N_12200,N_11512);
nor U13112 (N_13112,N_11615,N_11517);
xor U13113 (N_13113,N_11454,N_11885);
and U13114 (N_13114,N_12020,N_11420);
nand U13115 (N_13115,N_11442,N_11746);
nand U13116 (N_13116,N_11569,N_11692);
nor U13117 (N_13117,N_11551,N_11404);
or U13118 (N_13118,N_11574,N_12423);
nor U13119 (N_13119,N_12190,N_12016);
nand U13120 (N_13120,N_11968,N_12029);
nor U13121 (N_13121,N_12057,N_11839);
or U13122 (N_13122,N_11933,N_12086);
or U13123 (N_13123,N_12037,N_11560);
or U13124 (N_13124,N_11525,N_11573);
or U13125 (N_13125,N_11681,N_12444);
or U13126 (N_13126,N_11779,N_11306);
or U13127 (N_13127,N_11910,N_11863);
nor U13128 (N_13128,N_11650,N_11779);
nand U13129 (N_13129,N_12070,N_11945);
xor U13130 (N_13130,N_11376,N_11965);
and U13131 (N_13131,N_11309,N_12185);
nand U13132 (N_13132,N_12162,N_11913);
nor U13133 (N_13133,N_11778,N_11537);
or U13134 (N_13134,N_12479,N_11876);
nor U13135 (N_13135,N_12083,N_11777);
and U13136 (N_13136,N_12356,N_11300);
nor U13137 (N_13137,N_12157,N_11728);
or U13138 (N_13138,N_12458,N_12305);
xnor U13139 (N_13139,N_12116,N_11573);
and U13140 (N_13140,N_12067,N_11686);
or U13141 (N_13141,N_11941,N_11660);
xor U13142 (N_13142,N_12297,N_11653);
nand U13143 (N_13143,N_11635,N_11975);
or U13144 (N_13144,N_12320,N_12059);
xor U13145 (N_13145,N_12241,N_11383);
nor U13146 (N_13146,N_12382,N_11842);
and U13147 (N_13147,N_11381,N_12258);
nand U13148 (N_13148,N_11410,N_12397);
xor U13149 (N_13149,N_11835,N_11285);
xor U13150 (N_13150,N_11433,N_12269);
and U13151 (N_13151,N_11389,N_11412);
and U13152 (N_13152,N_11756,N_12063);
nand U13153 (N_13153,N_12250,N_12376);
xor U13154 (N_13154,N_12183,N_11763);
and U13155 (N_13155,N_11813,N_11521);
and U13156 (N_13156,N_11653,N_11520);
and U13157 (N_13157,N_11502,N_12250);
nand U13158 (N_13158,N_12097,N_12256);
nor U13159 (N_13159,N_11927,N_12428);
xnor U13160 (N_13160,N_11565,N_11302);
nand U13161 (N_13161,N_11359,N_11729);
or U13162 (N_13162,N_12223,N_11684);
nor U13163 (N_13163,N_12486,N_11838);
xnor U13164 (N_13164,N_11306,N_11859);
or U13165 (N_13165,N_12267,N_11280);
nor U13166 (N_13166,N_12245,N_11671);
nand U13167 (N_13167,N_12238,N_11311);
or U13168 (N_13168,N_11796,N_11347);
nor U13169 (N_13169,N_11635,N_11767);
and U13170 (N_13170,N_12221,N_11698);
or U13171 (N_13171,N_11756,N_12089);
or U13172 (N_13172,N_11444,N_11863);
nor U13173 (N_13173,N_12196,N_12405);
or U13174 (N_13174,N_11250,N_12080);
and U13175 (N_13175,N_11680,N_11388);
xor U13176 (N_13176,N_11413,N_12037);
and U13177 (N_13177,N_11309,N_11447);
nand U13178 (N_13178,N_12153,N_11811);
and U13179 (N_13179,N_12498,N_11274);
and U13180 (N_13180,N_12363,N_12272);
nor U13181 (N_13181,N_11802,N_11950);
xnor U13182 (N_13182,N_11661,N_11567);
or U13183 (N_13183,N_11320,N_11556);
nand U13184 (N_13184,N_11909,N_12394);
nor U13185 (N_13185,N_11965,N_12449);
nor U13186 (N_13186,N_11565,N_12371);
or U13187 (N_13187,N_12277,N_12348);
and U13188 (N_13188,N_11534,N_12117);
and U13189 (N_13189,N_11815,N_11794);
or U13190 (N_13190,N_11597,N_11873);
nand U13191 (N_13191,N_12029,N_11489);
nor U13192 (N_13192,N_11379,N_12058);
nor U13193 (N_13193,N_11432,N_12168);
nand U13194 (N_13194,N_11980,N_11613);
nor U13195 (N_13195,N_12007,N_11371);
and U13196 (N_13196,N_11638,N_11450);
or U13197 (N_13197,N_12092,N_12176);
nand U13198 (N_13198,N_11853,N_12103);
and U13199 (N_13199,N_11592,N_12111);
xnor U13200 (N_13200,N_12049,N_12150);
nor U13201 (N_13201,N_11597,N_11700);
or U13202 (N_13202,N_11736,N_12109);
nor U13203 (N_13203,N_12149,N_12371);
or U13204 (N_13204,N_11788,N_12231);
and U13205 (N_13205,N_11505,N_12245);
nor U13206 (N_13206,N_12407,N_12172);
or U13207 (N_13207,N_12072,N_11632);
nor U13208 (N_13208,N_11948,N_12004);
nor U13209 (N_13209,N_11505,N_11797);
nor U13210 (N_13210,N_11587,N_11948);
or U13211 (N_13211,N_11313,N_11271);
and U13212 (N_13212,N_11758,N_11782);
nor U13213 (N_13213,N_11618,N_11638);
and U13214 (N_13214,N_11319,N_11253);
and U13215 (N_13215,N_12150,N_12134);
or U13216 (N_13216,N_11799,N_11608);
or U13217 (N_13217,N_11506,N_11933);
and U13218 (N_13218,N_11328,N_11610);
xor U13219 (N_13219,N_11987,N_11780);
nor U13220 (N_13220,N_12218,N_12396);
or U13221 (N_13221,N_12039,N_12176);
or U13222 (N_13222,N_12225,N_11745);
and U13223 (N_13223,N_12063,N_11731);
nor U13224 (N_13224,N_12205,N_12112);
nor U13225 (N_13225,N_11851,N_12431);
nor U13226 (N_13226,N_11438,N_12443);
nor U13227 (N_13227,N_11274,N_11448);
xnor U13228 (N_13228,N_11822,N_12432);
nor U13229 (N_13229,N_12384,N_12020);
xor U13230 (N_13230,N_12028,N_12296);
xnor U13231 (N_13231,N_11282,N_12133);
and U13232 (N_13232,N_11257,N_11399);
nor U13233 (N_13233,N_12059,N_11332);
nor U13234 (N_13234,N_11629,N_11726);
nand U13235 (N_13235,N_11267,N_12278);
nor U13236 (N_13236,N_12100,N_11598);
or U13237 (N_13237,N_11415,N_11537);
nor U13238 (N_13238,N_11369,N_12250);
or U13239 (N_13239,N_11685,N_12023);
and U13240 (N_13240,N_11566,N_11822);
nand U13241 (N_13241,N_11493,N_12490);
nand U13242 (N_13242,N_11978,N_12492);
nand U13243 (N_13243,N_11277,N_11553);
xor U13244 (N_13244,N_11821,N_12381);
nor U13245 (N_13245,N_11588,N_11745);
nor U13246 (N_13246,N_12202,N_12002);
nand U13247 (N_13247,N_12218,N_12175);
and U13248 (N_13248,N_12283,N_12095);
and U13249 (N_13249,N_11760,N_12212);
or U13250 (N_13250,N_11860,N_12310);
nand U13251 (N_13251,N_11565,N_12079);
and U13252 (N_13252,N_11261,N_12122);
nor U13253 (N_13253,N_11415,N_11952);
nand U13254 (N_13254,N_11407,N_11308);
and U13255 (N_13255,N_11788,N_11267);
xnor U13256 (N_13256,N_11320,N_12468);
nand U13257 (N_13257,N_11683,N_11747);
and U13258 (N_13258,N_12390,N_11323);
and U13259 (N_13259,N_11427,N_11423);
or U13260 (N_13260,N_12384,N_11768);
nand U13261 (N_13261,N_12365,N_11434);
nor U13262 (N_13262,N_12110,N_11855);
xnor U13263 (N_13263,N_12344,N_12415);
nor U13264 (N_13264,N_11803,N_12051);
nor U13265 (N_13265,N_11693,N_12483);
or U13266 (N_13266,N_11866,N_11843);
nand U13267 (N_13267,N_11745,N_12464);
or U13268 (N_13268,N_11630,N_12370);
nor U13269 (N_13269,N_12425,N_11885);
xnor U13270 (N_13270,N_11624,N_11411);
xor U13271 (N_13271,N_11578,N_12124);
or U13272 (N_13272,N_11288,N_12133);
xnor U13273 (N_13273,N_12300,N_12011);
nor U13274 (N_13274,N_12033,N_11909);
xor U13275 (N_13275,N_12145,N_11943);
and U13276 (N_13276,N_12132,N_12196);
nand U13277 (N_13277,N_11543,N_12117);
or U13278 (N_13278,N_12284,N_12498);
and U13279 (N_13279,N_11507,N_12342);
and U13280 (N_13280,N_11893,N_11543);
and U13281 (N_13281,N_12113,N_12202);
or U13282 (N_13282,N_11555,N_11737);
or U13283 (N_13283,N_12367,N_11500);
and U13284 (N_13284,N_11373,N_12242);
or U13285 (N_13285,N_11327,N_11835);
or U13286 (N_13286,N_11564,N_11444);
or U13287 (N_13287,N_11485,N_12373);
xor U13288 (N_13288,N_12179,N_11408);
xnor U13289 (N_13289,N_11550,N_12078);
nand U13290 (N_13290,N_12218,N_12243);
nor U13291 (N_13291,N_12312,N_11291);
xnor U13292 (N_13292,N_12130,N_12062);
or U13293 (N_13293,N_11463,N_11926);
and U13294 (N_13294,N_11696,N_11718);
nor U13295 (N_13295,N_11755,N_11469);
nand U13296 (N_13296,N_11914,N_11482);
nand U13297 (N_13297,N_12395,N_12140);
or U13298 (N_13298,N_11944,N_11491);
or U13299 (N_13299,N_11580,N_11358);
or U13300 (N_13300,N_11345,N_12355);
nand U13301 (N_13301,N_12136,N_11448);
and U13302 (N_13302,N_11363,N_11514);
nand U13303 (N_13303,N_11930,N_11597);
nand U13304 (N_13304,N_11532,N_11832);
nor U13305 (N_13305,N_11656,N_11474);
xnor U13306 (N_13306,N_11517,N_12054);
and U13307 (N_13307,N_11953,N_11789);
nor U13308 (N_13308,N_12030,N_11522);
nand U13309 (N_13309,N_11961,N_12034);
nor U13310 (N_13310,N_11820,N_11768);
nand U13311 (N_13311,N_11790,N_11337);
or U13312 (N_13312,N_11798,N_12342);
or U13313 (N_13313,N_11312,N_12397);
nor U13314 (N_13314,N_12188,N_11265);
and U13315 (N_13315,N_12021,N_11355);
nor U13316 (N_13316,N_12347,N_11669);
nand U13317 (N_13317,N_11533,N_11960);
and U13318 (N_13318,N_12374,N_12349);
nor U13319 (N_13319,N_11446,N_12402);
or U13320 (N_13320,N_12196,N_11443);
nor U13321 (N_13321,N_11946,N_12347);
xor U13322 (N_13322,N_11634,N_11959);
and U13323 (N_13323,N_12219,N_12416);
nand U13324 (N_13324,N_12186,N_11676);
nor U13325 (N_13325,N_11481,N_12316);
or U13326 (N_13326,N_11717,N_11537);
xor U13327 (N_13327,N_12465,N_11645);
xor U13328 (N_13328,N_12082,N_12077);
and U13329 (N_13329,N_11584,N_12445);
and U13330 (N_13330,N_12106,N_12086);
or U13331 (N_13331,N_11720,N_12292);
and U13332 (N_13332,N_12158,N_12049);
nor U13333 (N_13333,N_11903,N_12380);
nor U13334 (N_13334,N_12182,N_11502);
nand U13335 (N_13335,N_11527,N_11468);
nand U13336 (N_13336,N_12397,N_11874);
nand U13337 (N_13337,N_12427,N_11409);
or U13338 (N_13338,N_11562,N_11631);
xnor U13339 (N_13339,N_12152,N_11366);
and U13340 (N_13340,N_11501,N_12256);
nor U13341 (N_13341,N_12312,N_11749);
and U13342 (N_13342,N_11636,N_12430);
nor U13343 (N_13343,N_12391,N_11838);
and U13344 (N_13344,N_11750,N_11401);
nor U13345 (N_13345,N_12236,N_12122);
nor U13346 (N_13346,N_11651,N_11776);
nand U13347 (N_13347,N_11507,N_11373);
nand U13348 (N_13348,N_12036,N_11585);
xnor U13349 (N_13349,N_12047,N_12333);
xnor U13350 (N_13350,N_12328,N_11430);
and U13351 (N_13351,N_12088,N_11505);
nand U13352 (N_13352,N_11736,N_11734);
nand U13353 (N_13353,N_11917,N_12179);
or U13354 (N_13354,N_12036,N_12277);
xnor U13355 (N_13355,N_12460,N_11668);
nand U13356 (N_13356,N_11533,N_11946);
nor U13357 (N_13357,N_12404,N_12262);
nor U13358 (N_13358,N_11252,N_11665);
xnor U13359 (N_13359,N_11477,N_11975);
or U13360 (N_13360,N_11455,N_11390);
nand U13361 (N_13361,N_12088,N_11339);
or U13362 (N_13362,N_11814,N_12301);
nor U13363 (N_13363,N_11622,N_12094);
nand U13364 (N_13364,N_11331,N_12376);
nor U13365 (N_13365,N_12267,N_11937);
xnor U13366 (N_13366,N_11772,N_12243);
or U13367 (N_13367,N_12315,N_11666);
nand U13368 (N_13368,N_12033,N_11738);
xnor U13369 (N_13369,N_11872,N_11330);
or U13370 (N_13370,N_12366,N_11686);
xor U13371 (N_13371,N_11298,N_12141);
nand U13372 (N_13372,N_12038,N_12430);
or U13373 (N_13373,N_11939,N_11937);
nand U13374 (N_13374,N_12395,N_12033);
or U13375 (N_13375,N_11351,N_11534);
nand U13376 (N_13376,N_11694,N_11491);
nor U13377 (N_13377,N_11487,N_11910);
xor U13378 (N_13378,N_11736,N_11300);
nor U13379 (N_13379,N_12125,N_12351);
and U13380 (N_13380,N_12033,N_11768);
nand U13381 (N_13381,N_11841,N_11363);
nor U13382 (N_13382,N_12478,N_11851);
nor U13383 (N_13383,N_12089,N_12245);
nand U13384 (N_13384,N_11933,N_11352);
nand U13385 (N_13385,N_11792,N_11310);
or U13386 (N_13386,N_11560,N_11925);
nor U13387 (N_13387,N_11614,N_11692);
nor U13388 (N_13388,N_11423,N_11747);
and U13389 (N_13389,N_11962,N_12170);
nand U13390 (N_13390,N_11996,N_11275);
nand U13391 (N_13391,N_11589,N_12499);
nor U13392 (N_13392,N_11781,N_11925);
nor U13393 (N_13393,N_11838,N_12175);
xnor U13394 (N_13394,N_11493,N_11446);
and U13395 (N_13395,N_11840,N_12096);
or U13396 (N_13396,N_11286,N_11324);
and U13397 (N_13397,N_11479,N_11278);
nor U13398 (N_13398,N_11870,N_12008);
nor U13399 (N_13399,N_12208,N_11255);
and U13400 (N_13400,N_11544,N_11491);
xor U13401 (N_13401,N_12271,N_11872);
nor U13402 (N_13402,N_12021,N_12153);
nor U13403 (N_13403,N_11945,N_12330);
or U13404 (N_13404,N_11606,N_12126);
nor U13405 (N_13405,N_12109,N_11604);
nand U13406 (N_13406,N_11493,N_12055);
nand U13407 (N_13407,N_11608,N_11853);
or U13408 (N_13408,N_11965,N_11589);
nand U13409 (N_13409,N_11509,N_11298);
or U13410 (N_13410,N_11491,N_11410);
and U13411 (N_13411,N_11826,N_11827);
or U13412 (N_13412,N_12089,N_11325);
or U13413 (N_13413,N_12029,N_11452);
nand U13414 (N_13414,N_12235,N_11855);
and U13415 (N_13415,N_11411,N_12070);
and U13416 (N_13416,N_11432,N_11317);
xnor U13417 (N_13417,N_11386,N_11644);
or U13418 (N_13418,N_11291,N_11588);
xor U13419 (N_13419,N_12354,N_12462);
nor U13420 (N_13420,N_12495,N_12251);
or U13421 (N_13421,N_12432,N_11547);
nor U13422 (N_13422,N_12375,N_11879);
xnor U13423 (N_13423,N_11628,N_12480);
xnor U13424 (N_13424,N_11498,N_11272);
nor U13425 (N_13425,N_12234,N_12268);
nand U13426 (N_13426,N_12374,N_11357);
or U13427 (N_13427,N_12051,N_11693);
nand U13428 (N_13428,N_12476,N_11775);
xnor U13429 (N_13429,N_11363,N_11671);
xor U13430 (N_13430,N_11923,N_11332);
xnor U13431 (N_13431,N_12110,N_12201);
nor U13432 (N_13432,N_11281,N_12241);
nor U13433 (N_13433,N_11427,N_11990);
nand U13434 (N_13434,N_11394,N_11827);
xor U13435 (N_13435,N_12219,N_12243);
or U13436 (N_13436,N_12264,N_11794);
and U13437 (N_13437,N_12436,N_11881);
and U13438 (N_13438,N_11573,N_11982);
or U13439 (N_13439,N_11483,N_12282);
xor U13440 (N_13440,N_11987,N_11899);
nand U13441 (N_13441,N_12472,N_12082);
or U13442 (N_13442,N_12187,N_11303);
nor U13443 (N_13443,N_12198,N_11977);
nor U13444 (N_13444,N_12317,N_11809);
and U13445 (N_13445,N_12416,N_11692);
nor U13446 (N_13446,N_11563,N_11806);
and U13447 (N_13447,N_12338,N_12059);
nand U13448 (N_13448,N_11709,N_12241);
nand U13449 (N_13449,N_12270,N_11491);
nand U13450 (N_13450,N_11848,N_12322);
and U13451 (N_13451,N_11826,N_12415);
nand U13452 (N_13452,N_11505,N_12379);
nand U13453 (N_13453,N_11476,N_11939);
nand U13454 (N_13454,N_11883,N_12004);
and U13455 (N_13455,N_11347,N_11676);
nor U13456 (N_13456,N_12124,N_11469);
xor U13457 (N_13457,N_12423,N_12190);
or U13458 (N_13458,N_12350,N_12072);
nor U13459 (N_13459,N_11334,N_12000);
nand U13460 (N_13460,N_11814,N_12272);
nor U13461 (N_13461,N_11441,N_11968);
or U13462 (N_13462,N_11648,N_12129);
or U13463 (N_13463,N_12267,N_12359);
and U13464 (N_13464,N_12463,N_11755);
and U13465 (N_13465,N_11935,N_11626);
or U13466 (N_13466,N_11878,N_11490);
nor U13467 (N_13467,N_11951,N_12023);
nand U13468 (N_13468,N_11320,N_12035);
xnor U13469 (N_13469,N_11443,N_11380);
or U13470 (N_13470,N_12099,N_11612);
and U13471 (N_13471,N_11674,N_11517);
xor U13472 (N_13472,N_12457,N_12086);
nand U13473 (N_13473,N_11947,N_11331);
and U13474 (N_13474,N_12058,N_11705);
xor U13475 (N_13475,N_11716,N_11486);
and U13476 (N_13476,N_11746,N_11516);
nand U13477 (N_13477,N_12373,N_11499);
xor U13478 (N_13478,N_12216,N_12239);
nand U13479 (N_13479,N_12334,N_11962);
nor U13480 (N_13480,N_12313,N_11667);
or U13481 (N_13481,N_12477,N_12190);
xnor U13482 (N_13482,N_12161,N_11530);
nor U13483 (N_13483,N_11629,N_11723);
or U13484 (N_13484,N_11700,N_11983);
or U13485 (N_13485,N_11817,N_11582);
nand U13486 (N_13486,N_11362,N_11287);
and U13487 (N_13487,N_11490,N_11786);
nand U13488 (N_13488,N_12003,N_11365);
and U13489 (N_13489,N_12430,N_12319);
xnor U13490 (N_13490,N_11785,N_11743);
and U13491 (N_13491,N_12019,N_11605);
nand U13492 (N_13492,N_12433,N_12426);
or U13493 (N_13493,N_12374,N_11298);
xor U13494 (N_13494,N_11973,N_11951);
and U13495 (N_13495,N_12164,N_11941);
or U13496 (N_13496,N_11743,N_11631);
xor U13497 (N_13497,N_12160,N_11326);
nand U13498 (N_13498,N_12022,N_11996);
and U13499 (N_13499,N_12194,N_12141);
nand U13500 (N_13500,N_11613,N_12405);
nand U13501 (N_13501,N_11882,N_12104);
and U13502 (N_13502,N_11510,N_11840);
xnor U13503 (N_13503,N_11321,N_12354);
nor U13504 (N_13504,N_12332,N_11463);
xnor U13505 (N_13505,N_11360,N_12242);
xnor U13506 (N_13506,N_11701,N_11538);
or U13507 (N_13507,N_12153,N_12081);
or U13508 (N_13508,N_12432,N_11978);
nand U13509 (N_13509,N_11834,N_11486);
and U13510 (N_13510,N_11753,N_12239);
or U13511 (N_13511,N_12334,N_11667);
nand U13512 (N_13512,N_11577,N_11640);
or U13513 (N_13513,N_11980,N_12068);
or U13514 (N_13514,N_11933,N_11781);
and U13515 (N_13515,N_11331,N_11721);
xnor U13516 (N_13516,N_11845,N_11912);
and U13517 (N_13517,N_11865,N_11533);
nor U13518 (N_13518,N_11703,N_12079);
nor U13519 (N_13519,N_11681,N_12036);
nand U13520 (N_13520,N_11263,N_12076);
xor U13521 (N_13521,N_12292,N_12282);
xnor U13522 (N_13522,N_12317,N_11784);
xor U13523 (N_13523,N_12012,N_11808);
nand U13524 (N_13524,N_12365,N_12055);
xnor U13525 (N_13525,N_12354,N_12280);
nand U13526 (N_13526,N_11650,N_12446);
and U13527 (N_13527,N_12224,N_12061);
nor U13528 (N_13528,N_11729,N_11845);
or U13529 (N_13529,N_11301,N_11286);
xor U13530 (N_13530,N_12343,N_11476);
nor U13531 (N_13531,N_11327,N_11382);
xnor U13532 (N_13532,N_11251,N_12364);
nor U13533 (N_13533,N_11628,N_11849);
xor U13534 (N_13534,N_12283,N_12453);
nand U13535 (N_13535,N_11520,N_11956);
and U13536 (N_13536,N_11687,N_11542);
nand U13537 (N_13537,N_12313,N_11776);
xnor U13538 (N_13538,N_11492,N_11346);
and U13539 (N_13539,N_11679,N_11702);
nor U13540 (N_13540,N_11792,N_11739);
xor U13541 (N_13541,N_12354,N_11968);
nor U13542 (N_13542,N_11625,N_12396);
nand U13543 (N_13543,N_11919,N_12182);
xnor U13544 (N_13544,N_11590,N_11694);
nor U13545 (N_13545,N_11426,N_12467);
or U13546 (N_13546,N_11993,N_11472);
and U13547 (N_13547,N_11638,N_12451);
xnor U13548 (N_13548,N_11973,N_11878);
or U13549 (N_13549,N_11856,N_11561);
or U13550 (N_13550,N_11617,N_12228);
or U13551 (N_13551,N_11646,N_12398);
nand U13552 (N_13552,N_11700,N_12291);
xnor U13553 (N_13553,N_12339,N_12014);
or U13554 (N_13554,N_12107,N_12254);
xnor U13555 (N_13555,N_11718,N_11984);
nor U13556 (N_13556,N_11530,N_11917);
xnor U13557 (N_13557,N_12273,N_11714);
nor U13558 (N_13558,N_12142,N_12437);
nand U13559 (N_13559,N_12347,N_12331);
nand U13560 (N_13560,N_12135,N_12273);
xor U13561 (N_13561,N_11368,N_12457);
and U13562 (N_13562,N_12259,N_11521);
nor U13563 (N_13563,N_11498,N_12472);
or U13564 (N_13564,N_11855,N_12244);
and U13565 (N_13565,N_12355,N_12104);
nand U13566 (N_13566,N_11321,N_11686);
nand U13567 (N_13567,N_12157,N_12226);
nand U13568 (N_13568,N_12285,N_11530);
or U13569 (N_13569,N_11883,N_11681);
xnor U13570 (N_13570,N_11700,N_11435);
xnor U13571 (N_13571,N_11398,N_11680);
nor U13572 (N_13572,N_12232,N_12353);
nand U13573 (N_13573,N_11655,N_12355);
xor U13574 (N_13574,N_12368,N_11915);
nand U13575 (N_13575,N_11574,N_12152);
nor U13576 (N_13576,N_11699,N_12436);
xnor U13577 (N_13577,N_11365,N_12425);
nor U13578 (N_13578,N_12318,N_12476);
and U13579 (N_13579,N_11313,N_12275);
or U13580 (N_13580,N_11709,N_12335);
xnor U13581 (N_13581,N_11286,N_11833);
nand U13582 (N_13582,N_11808,N_11876);
nand U13583 (N_13583,N_12354,N_12038);
nand U13584 (N_13584,N_12477,N_12383);
nand U13585 (N_13585,N_11926,N_11413);
nor U13586 (N_13586,N_11866,N_12351);
nor U13587 (N_13587,N_11886,N_11396);
nor U13588 (N_13588,N_11741,N_11682);
xor U13589 (N_13589,N_11447,N_11991);
xnor U13590 (N_13590,N_11816,N_12259);
or U13591 (N_13591,N_11378,N_12186);
and U13592 (N_13592,N_12129,N_12328);
xnor U13593 (N_13593,N_11508,N_11756);
nand U13594 (N_13594,N_11666,N_12244);
nand U13595 (N_13595,N_11642,N_12246);
and U13596 (N_13596,N_11305,N_11551);
xnor U13597 (N_13597,N_11942,N_11354);
nor U13598 (N_13598,N_11613,N_12341);
and U13599 (N_13599,N_11449,N_12143);
nand U13600 (N_13600,N_11876,N_11724);
nor U13601 (N_13601,N_11877,N_12109);
xor U13602 (N_13602,N_12217,N_12026);
and U13603 (N_13603,N_12312,N_11340);
or U13604 (N_13604,N_11666,N_12168);
xor U13605 (N_13605,N_11253,N_12279);
and U13606 (N_13606,N_12448,N_12115);
nand U13607 (N_13607,N_11805,N_11265);
nor U13608 (N_13608,N_11747,N_12090);
xnor U13609 (N_13609,N_12490,N_11459);
nor U13610 (N_13610,N_11473,N_12041);
nor U13611 (N_13611,N_12008,N_12292);
nor U13612 (N_13612,N_12019,N_12387);
nor U13613 (N_13613,N_12135,N_11736);
xnor U13614 (N_13614,N_11661,N_11734);
or U13615 (N_13615,N_11422,N_11995);
xnor U13616 (N_13616,N_11875,N_12072);
nor U13617 (N_13617,N_11724,N_12182);
nand U13618 (N_13618,N_11601,N_12446);
nor U13619 (N_13619,N_11437,N_11380);
or U13620 (N_13620,N_12045,N_11751);
and U13621 (N_13621,N_11488,N_12433);
and U13622 (N_13622,N_12293,N_12394);
and U13623 (N_13623,N_11548,N_11984);
and U13624 (N_13624,N_12452,N_12496);
xnor U13625 (N_13625,N_11321,N_11287);
and U13626 (N_13626,N_11566,N_11679);
and U13627 (N_13627,N_11978,N_11540);
or U13628 (N_13628,N_11638,N_11878);
xor U13629 (N_13629,N_11838,N_12371);
nand U13630 (N_13630,N_11392,N_11451);
nand U13631 (N_13631,N_11484,N_11738);
xor U13632 (N_13632,N_12157,N_12347);
xnor U13633 (N_13633,N_11492,N_12054);
or U13634 (N_13634,N_12401,N_12480);
or U13635 (N_13635,N_12200,N_11385);
xnor U13636 (N_13636,N_12128,N_12432);
xor U13637 (N_13637,N_11927,N_11695);
and U13638 (N_13638,N_12236,N_12462);
nor U13639 (N_13639,N_11716,N_11710);
xnor U13640 (N_13640,N_12215,N_12397);
or U13641 (N_13641,N_12165,N_11584);
or U13642 (N_13642,N_12390,N_12153);
or U13643 (N_13643,N_11449,N_12030);
xnor U13644 (N_13644,N_11299,N_11339);
or U13645 (N_13645,N_12058,N_12210);
or U13646 (N_13646,N_12093,N_11324);
nand U13647 (N_13647,N_11278,N_11564);
nand U13648 (N_13648,N_11754,N_11744);
and U13649 (N_13649,N_12271,N_12086);
nand U13650 (N_13650,N_11696,N_12236);
xor U13651 (N_13651,N_11825,N_12248);
and U13652 (N_13652,N_12001,N_11542);
nor U13653 (N_13653,N_12099,N_11528);
xor U13654 (N_13654,N_11905,N_11670);
and U13655 (N_13655,N_12085,N_11684);
nand U13656 (N_13656,N_11943,N_11531);
or U13657 (N_13657,N_12015,N_12046);
or U13658 (N_13658,N_11582,N_11309);
nor U13659 (N_13659,N_12220,N_11555);
nor U13660 (N_13660,N_11611,N_11536);
and U13661 (N_13661,N_12404,N_11593);
nand U13662 (N_13662,N_12254,N_11628);
or U13663 (N_13663,N_11482,N_11899);
or U13664 (N_13664,N_11619,N_11811);
or U13665 (N_13665,N_11535,N_11526);
and U13666 (N_13666,N_11534,N_11710);
or U13667 (N_13667,N_11989,N_12060);
and U13668 (N_13668,N_11458,N_11673);
nand U13669 (N_13669,N_12283,N_11769);
xor U13670 (N_13670,N_11507,N_11938);
and U13671 (N_13671,N_11599,N_12388);
xor U13672 (N_13672,N_12403,N_11662);
xor U13673 (N_13673,N_11475,N_11560);
and U13674 (N_13674,N_11800,N_11384);
xor U13675 (N_13675,N_11955,N_12326);
or U13676 (N_13676,N_11891,N_11950);
nor U13677 (N_13677,N_11628,N_11682);
and U13678 (N_13678,N_12165,N_11655);
nor U13679 (N_13679,N_11493,N_11801);
nor U13680 (N_13680,N_11620,N_12184);
xor U13681 (N_13681,N_12276,N_11941);
nand U13682 (N_13682,N_11880,N_11355);
nand U13683 (N_13683,N_12251,N_11384);
nor U13684 (N_13684,N_12004,N_12319);
xnor U13685 (N_13685,N_11481,N_12087);
nand U13686 (N_13686,N_12216,N_12169);
nor U13687 (N_13687,N_11277,N_12090);
xnor U13688 (N_13688,N_11645,N_12434);
or U13689 (N_13689,N_11972,N_11525);
nor U13690 (N_13690,N_11957,N_11825);
or U13691 (N_13691,N_11463,N_12438);
xnor U13692 (N_13692,N_11374,N_11697);
xor U13693 (N_13693,N_12277,N_12245);
or U13694 (N_13694,N_11858,N_11580);
and U13695 (N_13695,N_11822,N_11706);
or U13696 (N_13696,N_11816,N_11715);
nand U13697 (N_13697,N_12266,N_11586);
xnor U13698 (N_13698,N_12091,N_11984);
and U13699 (N_13699,N_11371,N_11703);
nand U13700 (N_13700,N_11365,N_11906);
and U13701 (N_13701,N_11312,N_11561);
nor U13702 (N_13702,N_12043,N_12036);
xnor U13703 (N_13703,N_11487,N_11477);
and U13704 (N_13704,N_11462,N_12174);
or U13705 (N_13705,N_12325,N_11545);
nor U13706 (N_13706,N_11597,N_12275);
and U13707 (N_13707,N_11319,N_12142);
nand U13708 (N_13708,N_11618,N_11607);
nand U13709 (N_13709,N_11699,N_11300);
or U13710 (N_13710,N_11577,N_11479);
and U13711 (N_13711,N_12342,N_11309);
xnor U13712 (N_13712,N_12039,N_11894);
nor U13713 (N_13713,N_11852,N_11353);
xor U13714 (N_13714,N_11453,N_11733);
and U13715 (N_13715,N_11694,N_11362);
or U13716 (N_13716,N_11459,N_12206);
nand U13717 (N_13717,N_11891,N_12255);
xor U13718 (N_13718,N_11755,N_11376);
nor U13719 (N_13719,N_11965,N_11447);
xnor U13720 (N_13720,N_11717,N_12449);
or U13721 (N_13721,N_11833,N_12313);
and U13722 (N_13722,N_11400,N_12002);
nand U13723 (N_13723,N_12344,N_12346);
and U13724 (N_13724,N_12413,N_11750);
nand U13725 (N_13725,N_12302,N_12063);
nand U13726 (N_13726,N_11904,N_11265);
nand U13727 (N_13727,N_11510,N_12227);
xor U13728 (N_13728,N_11985,N_11739);
nor U13729 (N_13729,N_11328,N_11398);
and U13730 (N_13730,N_12112,N_11699);
nor U13731 (N_13731,N_11953,N_12223);
or U13732 (N_13732,N_12300,N_11318);
nand U13733 (N_13733,N_12334,N_12107);
or U13734 (N_13734,N_11279,N_12457);
nand U13735 (N_13735,N_12456,N_12469);
and U13736 (N_13736,N_11883,N_11403);
and U13737 (N_13737,N_12241,N_11719);
xnor U13738 (N_13738,N_12493,N_12355);
xnor U13739 (N_13739,N_11422,N_12257);
or U13740 (N_13740,N_12278,N_11962);
nor U13741 (N_13741,N_11390,N_12122);
xor U13742 (N_13742,N_11410,N_11768);
and U13743 (N_13743,N_11304,N_11390);
nor U13744 (N_13744,N_11687,N_11430);
nand U13745 (N_13745,N_11535,N_11769);
xor U13746 (N_13746,N_12149,N_11530);
and U13747 (N_13747,N_11378,N_11950);
xnor U13748 (N_13748,N_12356,N_12453);
and U13749 (N_13749,N_12384,N_11467);
xnor U13750 (N_13750,N_13572,N_12831);
or U13751 (N_13751,N_13634,N_12754);
nor U13752 (N_13752,N_13594,N_13614);
nor U13753 (N_13753,N_12809,N_13600);
nand U13754 (N_13754,N_12784,N_12583);
nor U13755 (N_13755,N_13025,N_13390);
nor U13756 (N_13756,N_12752,N_13183);
and U13757 (N_13757,N_13420,N_13586);
nor U13758 (N_13758,N_13457,N_13418);
and U13759 (N_13759,N_13492,N_12565);
xor U13760 (N_13760,N_12953,N_13355);
nor U13761 (N_13761,N_13404,N_13141);
and U13762 (N_13762,N_13437,N_13607);
xnor U13763 (N_13763,N_12526,N_13350);
and U13764 (N_13764,N_13721,N_13646);
or U13765 (N_13765,N_13740,N_13555);
nor U13766 (N_13766,N_13160,N_12760);
and U13767 (N_13767,N_13014,N_12668);
or U13768 (N_13768,N_13063,N_12511);
or U13769 (N_13769,N_13387,N_12876);
nor U13770 (N_13770,N_13030,N_13367);
xnor U13771 (N_13771,N_12518,N_13294);
and U13772 (N_13772,N_13015,N_13299);
xnor U13773 (N_13773,N_13202,N_12884);
nor U13774 (N_13774,N_13523,N_12543);
nor U13775 (N_13775,N_12827,N_12755);
or U13776 (N_13776,N_13322,N_12599);
xnor U13777 (N_13777,N_12531,N_13538);
nand U13778 (N_13778,N_13564,N_13301);
nand U13779 (N_13779,N_13349,N_13049);
nor U13780 (N_13780,N_12747,N_12657);
nand U13781 (N_13781,N_13217,N_13267);
and U13782 (N_13782,N_13507,N_12708);
nor U13783 (N_13783,N_13700,N_12846);
xor U13784 (N_13784,N_12776,N_13051);
nor U13785 (N_13785,N_12765,N_12503);
or U13786 (N_13786,N_13497,N_12701);
nand U13787 (N_13787,N_12553,N_12537);
nand U13788 (N_13788,N_12541,N_12905);
nor U13789 (N_13789,N_13375,N_12629);
and U13790 (N_13790,N_13466,N_13569);
nand U13791 (N_13791,N_13529,N_12542);
nand U13792 (N_13792,N_13442,N_12788);
xnor U13793 (N_13793,N_13577,N_13395);
nor U13794 (N_13794,N_13251,N_13303);
xor U13795 (N_13795,N_12912,N_13312);
nand U13796 (N_13796,N_13280,N_13494);
nor U13797 (N_13797,N_13239,N_13173);
xnor U13798 (N_13798,N_13552,N_13091);
or U13799 (N_13799,N_12660,N_13238);
nor U13800 (N_13800,N_12648,N_12800);
nand U13801 (N_13801,N_12898,N_12900);
and U13802 (N_13802,N_13372,N_13508);
nand U13803 (N_13803,N_13535,N_12761);
and U13804 (N_13804,N_13416,N_12603);
xnor U13805 (N_13805,N_13448,N_12814);
and U13806 (N_13806,N_13174,N_13369);
or U13807 (N_13807,N_13140,N_12819);
or U13808 (N_13808,N_13326,N_12966);
nand U13809 (N_13809,N_13116,N_12714);
and U13810 (N_13810,N_13084,N_13444);
and U13811 (N_13811,N_12895,N_13727);
nand U13812 (N_13812,N_13694,N_12624);
xnor U13813 (N_13813,N_12763,N_12973);
and U13814 (N_13814,N_13113,N_12727);
nand U13815 (N_13815,N_13467,N_12709);
and U13816 (N_13816,N_12866,N_12934);
nand U13817 (N_13817,N_13119,N_13676);
xnor U13818 (N_13818,N_12721,N_12829);
nand U13819 (N_13819,N_13479,N_13641);
and U13820 (N_13820,N_12688,N_12567);
and U13821 (N_13821,N_12970,N_13002);
nor U13822 (N_13822,N_13132,N_13595);
nand U13823 (N_13823,N_13547,N_13008);
or U13824 (N_13824,N_13582,N_12611);
or U13825 (N_13825,N_13500,N_13710);
or U13826 (N_13826,N_12595,N_13283);
nand U13827 (N_13827,N_13075,N_12997);
xor U13828 (N_13828,N_13415,N_13168);
nand U13829 (N_13829,N_13624,N_13636);
nor U13830 (N_13830,N_12949,N_12628);
xnor U13831 (N_13831,N_13685,N_13601);
nor U13832 (N_13832,N_13164,N_13240);
nand U13833 (N_13833,N_12910,N_13150);
nor U13834 (N_13834,N_12520,N_13609);
nand U13835 (N_13835,N_13034,N_13452);
nand U13836 (N_13836,N_12886,N_12664);
nor U13837 (N_13837,N_13276,N_13617);
nor U13838 (N_13838,N_13257,N_13412);
nand U13839 (N_13839,N_12878,N_12820);
nand U13840 (N_13840,N_13458,N_13491);
and U13841 (N_13841,N_12710,N_12773);
nand U13842 (N_13842,N_13275,N_12625);
nand U13843 (N_13843,N_13287,N_13481);
nand U13844 (N_13844,N_13521,N_13201);
nor U13845 (N_13845,N_13365,N_13259);
or U13846 (N_13846,N_12667,N_13623);
and U13847 (N_13847,N_12848,N_13510);
or U13848 (N_13848,N_13172,N_13498);
nor U13849 (N_13849,N_13593,N_12570);
and U13850 (N_13850,N_13425,N_12580);
or U13851 (N_13851,N_13035,N_13602);
nand U13852 (N_13852,N_12892,N_13081);
nor U13853 (N_13853,N_13319,N_13263);
or U13854 (N_13854,N_13225,N_13208);
nand U13855 (N_13855,N_13477,N_12587);
or U13856 (N_13856,N_13731,N_12746);
and U13857 (N_13857,N_13255,N_12988);
or U13858 (N_13858,N_12575,N_12823);
xnor U13859 (N_13859,N_13126,N_13249);
and U13860 (N_13860,N_13707,N_13683);
nand U13861 (N_13861,N_13668,N_13188);
xor U13862 (N_13862,N_13468,N_13534);
nand U13863 (N_13863,N_12920,N_12529);
xor U13864 (N_13864,N_12641,N_13677);
xor U13865 (N_13865,N_12929,N_13264);
nor U13866 (N_13866,N_13664,N_12650);
and U13867 (N_13867,N_13662,N_13094);
and U13868 (N_13868,N_12644,N_12513);
nor U13869 (N_13869,N_13336,N_13268);
or U13870 (N_13870,N_13407,N_13509);
nand U13871 (N_13871,N_13151,N_12725);
and U13872 (N_13872,N_13243,N_12914);
nand U13873 (N_13873,N_13392,N_13179);
nand U13874 (N_13874,N_12992,N_13525);
nand U13875 (N_13875,N_13745,N_13124);
xor U13876 (N_13876,N_13675,N_13310);
nand U13877 (N_13877,N_12706,N_12535);
nand U13878 (N_13878,N_13161,N_13660);
or U13879 (N_13879,N_12781,N_12649);
or U13880 (N_13880,N_13199,N_13135);
nor U13881 (N_13881,N_12850,N_12861);
or U13882 (N_13882,N_13578,N_12692);
nand U13883 (N_13883,N_12837,N_13215);
nor U13884 (N_13884,N_12843,N_12798);
nor U13885 (N_13885,N_13060,N_13421);
and U13886 (N_13886,N_12830,N_12631);
nor U13887 (N_13887,N_13433,N_13456);
nand U13888 (N_13888,N_13020,N_13105);
nand U13889 (N_13889,N_12960,N_13180);
xnor U13890 (N_13890,N_13347,N_13483);
xnor U13891 (N_13891,N_12715,N_12944);
and U13892 (N_13892,N_12569,N_12534);
nor U13893 (N_13893,N_13170,N_12919);
or U13894 (N_13894,N_12998,N_13505);
and U13895 (N_13895,N_13134,N_13110);
nor U13896 (N_13896,N_13650,N_13695);
and U13897 (N_13897,N_13331,N_12612);
xnor U13898 (N_13898,N_13464,N_12557);
nor U13899 (N_13899,N_13562,N_13001);
xnor U13900 (N_13900,N_13496,N_12869);
nor U13901 (N_13901,N_13654,N_13591);
xor U13902 (N_13902,N_12604,N_13717);
nand U13903 (N_13903,N_13450,N_12937);
nand U13904 (N_13904,N_12958,N_13621);
nand U13905 (N_13905,N_13175,N_13226);
xor U13906 (N_13906,N_12844,N_13645);
xor U13907 (N_13907,N_12608,N_13305);
nand U13908 (N_13908,N_13428,N_12681);
xnor U13909 (N_13909,N_13596,N_13203);
or U13910 (N_13910,N_13682,N_13096);
nor U13911 (N_13911,N_12510,N_13478);
nand U13912 (N_13912,N_13061,N_12505);
xor U13913 (N_13913,N_13743,N_13561);
and U13914 (N_13914,N_12787,N_13320);
nor U13915 (N_13915,N_13380,N_13085);
nor U13916 (N_13916,N_13028,N_13269);
nor U13917 (N_13917,N_13482,N_12780);
nand U13918 (N_13918,N_13068,N_13518);
nor U13919 (N_13919,N_13459,N_13426);
and U13920 (N_13920,N_12556,N_13233);
nor U13921 (N_13921,N_13473,N_12945);
nor U13922 (N_13922,N_13619,N_12699);
nor U13923 (N_13923,N_12769,N_13551);
nand U13924 (N_13924,N_13246,N_13629);
and U13925 (N_13925,N_12799,N_13036);
and U13926 (N_13926,N_12620,N_12768);
nand U13927 (N_13927,N_12842,N_12855);
or U13928 (N_13928,N_13353,N_13351);
or U13929 (N_13929,N_12658,N_13689);
and U13930 (N_13930,N_13746,N_13204);
or U13931 (N_13931,N_12555,N_13651);
nand U13932 (N_13932,N_12874,N_13079);
nor U13933 (N_13933,N_12563,N_12736);
nor U13934 (N_13934,N_12528,N_13245);
xor U13935 (N_13935,N_13133,N_13697);
nor U13936 (N_13936,N_13566,N_13658);
xnor U13937 (N_13937,N_13388,N_12775);
nand U13938 (N_13938,N_13328,N_13129);
xnor U13939 (N_13939,N_13401,N_13222);
xnor U13940 (N_13940,N_12821,N_12858);
xor U13941 (N_13941,N_13516,N_12803);
nand U13942 (N_13942,N_12750,N_12719);
or U13943 (N_13943,N_12815,N_13678);
nor U13944 (N_13944,N_12981,N_13059);
nor U13945 (N_13945,N_13252,N_13206);
and U13946 (N_13946,N_13608,N_13329);
nor U13947 (N_13947,N_13258,N_12693);
nor U13948 (N_13948,N_13106,N_13053);
and U13949 (N_13949,N_12753,N_12955);
nand U13950 (N_13950,N_12965,N_13220);
xnor U13951 (N_13951,N_12550,N_13099);
nor U13952 (N_13952,N_13356,N_12656);
nor U13953 (N_13953,N_13453,N_13413);
and U13954 (N_13954,N_12882,N_12610);
nand U13955 (N_13955,N_13432,N_12530);
nor U13956 (N_13956,N_13234,N_12839);
or U13957 (N_13957,N_12952,N_13363);
nand U13958 (N_13958,N_13130,N_13352);
nor U13959 (N_13959,N_13325,N_13589);
nor U13960 (N_13960,N_13019,N_13396);
nand U13961 (N_13961,N_13089,N_13346);
nor U13962 (N_13962,N_12947,N_12507);
xnor U13963 (N_13963,N_13343,N_12717);
xnor U13964 (N_13964,N_13655,N_12740);
nor U13965 (N_13965,N_13573,N_12732);
nand U13966 (N_13966,N_12979,N_12852);
xor U13967 (N_13967,N_12700,N_12812);
or U13968 (N_13968,N_13469,N_12805);
xor U13969 (N_13969,N_13144,N_12909);
nand U13970 (N_13970,N_12825,N_13604);
or U13971 (N_13971,N_13190,N_12993);
nor U13972 (N_13972,N_13315,N_13272);
and U13973 (N_13973,N_12857,N_13550);
nand U13974 (N_13974,N_12893,N_13253);
nand U13975 (N_13975,N_13524,N_12508);
nand U13976 (N_13976,N_12590,N_13649);
nand U13977 (N_13977,N_12875,N_12916);
xor U13978 (N_13978,N_12524,N_12921);
nor U13979 (N_13979,N_13409,N_13295);
nand U13980 (N_13980,N_12698,N_13581);
or U13981 (N_13981,N_13149,N_12730);
and U13982 (N_13982,N_12606,N_13712);
xor U13983 (N_13983,N_13157,N_13182);
xor U13984 (N_13984,N_13537,N_13670);
or U13985 (N_13985,N_12728,N_12943);
or U13986 (N_13986,N_12990,N_12972);
nand U13987 (N_13987,N_12817,N_12642);
xor U13988 (N_13988,N_12593,N_13335);
nand U13989 (N_13989,N_13513,N_12907);
and U13990 (N_13990,N_13570,N_13207);
nand U13991 (N_13991,N_13377,N_13383);
and U13992 (N_13992,N_13115,N_13041);
and U13993 (N_13993,N_12976,N_13309);
and U13994 (N_13994,N_13023,N_13490);
and U13995 (N_13995,N_13114,N_13127);
nor U13996 (N_13996,N_13200,N_13337);
nand U13997 (N_13997,N_12836,N_12963);
or U13998 (N_13998,N_13038,N_12742);
xnor U13999 (N_13999,N_12926,N_12885);
xnor U14000 (N_14000,N_13656,N_13638);
nand U14001 (N_14001,N_13422,N_12635);
or U14002 (N_14002,N_13394,N_13307);
nor U14003 (N_14003,N_12654,N_12984);
or U14004 (N_14004,N_13567,N_12774);
xnor U14005 (N_14005,N_13027,N_12991);
and U14006 (N_14006,N_12581,N_12527);
xor U14007 (N_14007,N_12764,N_13576);
xnor U14008 (N_14008,N_13410,N_13613);
nor U14009 (N_14009,N_12501,N_13587);
nor U14010 (N_14010,N_13158,N_12822);
nor U14011 (N_14011,N_13332,N_12643);
nor U14012 (N_14012,N_12655,N_12633);
or U14013 (N_14013,N_13112,N_12927);
xnor U14014 (N_14014,N_13288,N_13087);
and U14015 (N_14015,N_13622,N_12665);
xnor U14016 (N_14016,N_13663,N_12637);
nor U14017 (N_14017,N_12645,N_13317);
nor U14018 (N_14018,N_13431,N_13612);
and U14019 (N_14019,N_13000,N_13393);
and U14020 (N_14020,N_12801,N_13072);
or U14021 (N_14021,N_12577,N_13511);
nand U14022 (N_14022,N_12999,N_13358);
xnor U14023 (N_14023,N_13659,N_13493);
nor U14024 (N_14024,N_13644,N_13533);
and U14025 (N_14025,N_13443,N_13739);
or U14026 (N_14026,N_13308,N_13704);
xor U14027 (N_14027,N_12516,N_12720);
and U14028 (N_14028,N_13440,N_13147);
and U14029 (N_14029,N_13403,N_13434);
nand U14030 (N_14030,N_12521,N_12666);
nor U14031 (N_14031,N_13417,N_13300);
or U14032 (N_14032,N_13118,N_13445);
xor U14033 (N_14033,N_12770,N_12639);
or U14034 (N_14034,N_13748,N_12942);
and U14035 (N_14035,N_13583,N_13101);
and U14036 (N_14036,N_13361,N_13429);
xor U14037 (N_14037,N_13250,N_13736);
nor U14038 (N_14038,N_13009,N_12930);
xnor U14039 (N_14039,N_13495,N_13720);
nand U14040 (N_14040,N_13040,N_13185);
nor U14041 (N_14041,N_13423,N_13184);
nand U14042 (N_14042,N_13177,N_13642);
nor U14043 (N_14043,N_12703,N_12523);
nand U14044 (N_14044,N_12881,N_13078);
or U14045 (N_14045,N_13050,N_13620);
xor U14046 (N_14046,N_13667,N_13397);
nand U14047 (N_14047,N_12807,N_13155);
nand U14048 (N_14048,N_13323,N_12562);
xor U14049 (N_14049,N_13166,N_12946);
nor U14050 (N_14050,N_12757,N_12586);
or U14051 (N_14051,N_12538,N_12684);
nand U14052 (N_14052,N_12982,N_12661);
xnor U14053 (N_14053,N_13626,N_13539);
nor U14054 (N_14054,N_13064,N_13398);
nor U14055 (N_14055,N_12804,N_13556);
or U14056 (N_14056,N_12585,N_12879);
and U14057 (N_14057,N_13705,N_12908);
nor U14058 (N_14058,N_13043,N_12794);
xnor U14059 (N_14059,N_13120,N_12578);
and U14060 (N_14060,N_13230,N_12544);
and U14061 (N_14061,N_13430,N_13474);
and U14062 (N_14062,N_12572,N_12672);
nand U14063 (N_14063,N_12536,N_12670);
and U14064 (N_14064,N_13324,N_12500);
or U14065 (N_14065,N_13679,N_12864);
nor U14066 (N_14066,N_13055,N_12880);
xnor U14067 (N_14067,N_13005,N_13631);
and U14068 (N_14068,N_12647,N_13730);
nor U14069 (N_14069,N_12828,N_13266);
xor U14070 (N_14070,N_13057,N_12561);
xor U14071 (N_14071,N_12579,N_12724);
or U14072 (N_14072,N_13598,N_12677);
xor U14073 (N_14073,N_13546,N_13709);
nand U14074 (N_14074,N_13687,N_13599);
and U14075 (N_14075,N_13108,N_13384);
xnor U14076 (N_14076,N_13153,N_13368);
nand U14077 (N_14077,N_12696,N_13665);
xor U14078 (N_14078,N_12834,N_12896);
xor U14079 (N_14079,N_13545,N_12786);
nand U14080 (N_14080,N_13643,N_12867);
xnor U14081 (N_14081,N_13512,N_12903);
nor U14082 (N_14082,N_13066,N_13506);
xor U14083 (N_14083,N_13530,N_13327);
xor U14084 (N_14084,N_13714,N_12634);
xnor U14085 (N_14085,N_13152,N_13159);
xnor U14086 (N_14086,N_12969,N_13022);
and U14087 (N_14087,N_12616,N_12597);
or U14088 (N_14088,N_13360,N_13724);
nor U14089 (N_14089,N_13042,N_12676);
or U14090 (N_14090,N_13104,N_12589);
and U14091 (N_14091,N_12795,N_12968);
or U14092 (N_14092,N_12948,N_13411);
xor U14093 (N_14093,N_12872,N_12689);
xnor U14094 (N_14094,N_12959,N_12932);
xnor U14095 (N_14095,N_13376,N_12554);
nand U14096 (N_14096,N_12694,N_12957);
xnor U14097 (N_14097,N_13070,N_12704);
or U14098 (N_14098,N_13029,N_12762);
and U14099 (N_14099,N_13242,N_12552);
nor U14100 (N_14100,N_13205,N_12918);
and U14101 (N_14101,N_12729,N_12766);
and U14102 (N_14102,N_13558,N_13293);
and U14103 (N_14103,N_13405,N_12756);
xnor U14104 (N_14104,N_13447,N_12854);
or U14105 (N_14105,N_13639,N_12749);
and U14106 (N_14106,N_13306,N_12797);
nor U14107 (N_14107,N_12978,N_13499);
or U14108 (N_14108,N_12767,N_13548);
nand U14109 (N_14109,N_12539,N_13735);
nor U14110 (N_14110,N_12935,N_13742);
and U14111 (N_14111,N_13344,N_13193);
and U14112 (N_14112,N_12682,N_13406);
nor U14113 (N_14113,N_12790,N_12811);
nor U14114 (N_14114,N_13359,N_13633);
nor U14115 (N_14115,N_13391,N_13145);
xnor U14116 (N_14116,N_13291,N_12726);
or U14117 (N_14117,N_13378,N_13673);
or U14118 (N_14118,N_12782,N_13542);
nand U14119 (N_14119,N_13637,N_13711);
xnor U14120 (N_14120,N_13543,N_13235);
nand U14121 (N_14121,N_12925,N_13733);
xnor U14122 (N_14122,N_13674,N_13610);
nand U14123 (N_14123,N_12983,N_13402);
and U14124 (N_14124,N_13071,N_13098);
nand U14125 (N_14125,N_13374,N_13178);
nand U14126 (N_14126,N_12877,N_12713);
xor U14127 (N_14127,N_12652,N_12928);
or U14128 (N_14128,N_12659,N_12564);
nand U14129 (N_14129,N_12824,N_13590);
or U14130 (N_14130,N_12517,N_13515);
nand U14131 (N_14131,N_12890,N_12987);
and U14132 (N_14132,N_13054,N_12705);
xnor U14133 (N_14133,N_12940,N_12626);
nand U14134 (N_14134,N_12964,N_12941);
xnor U14135 (N_14135,N_13379,N_12924);
xnor U14136 (N_14136,N_13554,N_12617);
nor U14137 (N_14137,N_13248,N_13128);
or U14138 (N_14138,N_13143,N_12791);
and U14139 (N_14139,N_12818,N_13648);
nor U14140 (N_14140,N_13097,N_13348);
or U14141 (N_14141,N_13640,N_13018);
nor U14142 (N_14142,N_12678,N_13262);
nand U14143 (N_14143,N_13165,N_12954);
xnor U14144 (N_14144,N_13285,N_13345);
xnor U14145 (N_14145,N_13436,N_13065);
nand U14146 (N_14146,N_13304,N_13321);
and U14147 (N_14147,N_12640,N_13615);
and U14148 (N_14148,N_12618,N_12588);
nor U14149 (N_14149,N_13585,N_13354);
nor U14150 (N_14150,N_13502,N_13460);
or U14151 (N_14151,N_12697,N_12549);
nand U14152 (N_14152,N_13454,N_13504);
nor U14153 (N_14153,N_13635,N_12931);
and U14154 (N_14154,N_12810,N_13194);
nand U14155 (N_14155,N_12826,N_12522);
or U14156 (N_14156,N_13139,N_13451);
xnor U14157 (N_14157,N_12514,N_13031);
nand U14158 (N_14158,N_12950,N_13462);
or U14159 (N_14159,N_13625,N_13540);
nand U14160 (N_14160,N_13273,N_13181);
xor U14161 (N_14161,N_13501,N_13284);
nor U14162 (N_14162,N_13652,N_13290);
nor U14163 (N_14163,N_12887,N_12568);
xor U14164 (N_14164,N_12591,N_13080);
nor U14165 (N_14165,N_12547,N_12690);
nand U14166 (N_14166,N_13461,N_12687);
nor U14167 (N_14167,N_13270,N_13111);
nand U14168 (N_14168,N_13292,N_12751);
and U14169 (N_14169,N_13296,N_13439);
nand U14170 (N_14170,N_13485,N_12638);
nand U14171 (N_14171,N_13247,N_13381);
xnor U14172 (N_14172,N_13568,N_12707);
and U14173 (N_14173,N_13039,N_12838);
nor U14174 (N_14174,N_12546,N_13357);
or U14175 (N_14175,N_13122,N_13399);
nor U14176 (N_14176,N_13047,N_13256);
xnor U14177 (N_14177,N_13187,N_12601);
nor U14178 (N_14178,N_13012,N_12632);
or U14179 (N_14179,N_12985,N_12833);
or U14180 (N_14180,N_12739,N_13544);
xor U14181 (N_14181,N_12783,N_12662);
nand U14182 (N_14182,N_13298,N_13486);
and U14183 (N_14183,N_12911,N_13647);
nand U14184 (N_14184,N_13435,N_12995);
or U14185 (N_14185,N_12777,N_12598);
and U14186 (N_14186,N_13463,N_13691);
xnor U14187 (N_14187,N_12913,N_13520);
or U14188 (N_14188,N_13074,N_13703);
and U14189 (N_14189,N_12738,N_12971);
nor U14190 (N_14190,N_13167,N_13661);
nand U14191 (N_14191,N_13227,N_13191);
nand U14192 (N_14192,N_12744,N_12986);
or U14193 (N_14193,N_13236,N_12594);
xnor U14194 (N_14194,N_12735,N_12596);
or U14195 (N_14195,N_12683,N_12863);
or U14196 (N_14196,N_12551,N_13209);
xor U14197 (N_14197,N_13519,N_13282);
xor U14198 (N_14198,N_13475,N_13016);
nand U14199 (N_14199,N_13732,N_13389);
and U14200 (N_14200,N_13557,N_13488);
nand U14201 (N_14201,N_13062,N_13719);
nor U14202 (N_14202,N_13069,N_13716);
xor U14203 (N_14203,N_12771,N_13261);
xnor U14204 (N_14204,N_12994,N_12915);
nand U14205 (N_14205,N_12675,N_12785);
nand U14206 (N_14206,N_13092,N_13414);
or U14207 (N_14207,N_13192,N_13142);
nor U14208 (N_14208,N_13588,N_13076);
nor U14209 (N_14209,N_13163,N_12851);
or U14210 (N_14210,N_12980,N_12845);
or U14211 (N_14211,N_13297,N_12956);
nand U14212 (N_14212,N_13722,N_13702);
and U14213 (N_14213,N_13314,N_13522);
xor U14214 (N_14214,N_13370,N_13455);
or U14215 (N_14215,N_12792,N_13690);
nand U14216 (N_14216,N_12899,N_12623);
xor U14217 (N_14217,N_12977,N_13154);
xor U14218 (N_14218,N_13339,N_12619);
and U14219 (N_14219,N_12891,N_12685);
nand U14220 (N_14220,N_13340,N_12600);
xor U14221 (N_14221,N_13169,N_12651);
and U14222 (N_14222,N_12967,N_12663);
and U14223 (N_14223,N_13013,N_13366);
xnor U14224 (N_14224,N_13470,N_12559);
or U14225 (N_14225,N_12607,N_13669);
nor U14226 (N_14226,N_13077,N_13630);
nor U14227 (N_14227,N_12975,N_13052);
or U14228 (N_14228,N_12802,N_12576);
or U14229 (N_14229,N_12722,N_13254);
or U14230 (N_14230,N_12759,N_12856);
or U14231 (N_14231,N_12630,N_12716);
nand U14232 (N_14232,N_13575,N_13371);
nand U14233 (N_14233,N_13471,N_13232);
xnor U14234 (N_14234,N_12574,N_13563);
xor U14235 (N_14235,N_13228,N_12758);
xor U14236 (N_14236,N_13083,N_13713);
nor U14237 (N_14237,N_13277,N_13006);
nor U14238 (N_14238,N_13046,N_13058);
and U14239 (N_14239,N_12859,N_13044);
and U14240 (N_14240,N_12894,N_12515);
or U14241 (N_14241,N_12686,N_12584);
nand U14242 (N_14242,N_12862,N_13737);
or U14243 (N_14243,N_13017,N_12674);
nand U14244 (N_14244,N_13362,N_12653);
nand U14245 (N_14245,N_13316,N_12873);
or U14246 (N_14246,N_12545,N_13278);
nand U14247 (N_14247,N_12695,N_13465);
or U14248 (N_14248,N_12939,N_12868);
nand U14249 (N_14249,N_12849,N_12860);
and U14250 (N_14250,N_13197,N_13244);
xnor U14251 (N_14251,N_13584,N_12540);
or U14252 (N_14252,N_13313,N_13734);
and U14253 (N_14253,N_12870,N_13441);
and U14254 (N_14254,N_12847,N_12883);
nor U14255 (N_14255,N_13382,N_13010);
nand U14256 (N_14256,N_13487,N_12906);
nor U14257 (N_14257,N_12602,N_13427);
and U14258 (N_14258,N_12718,N_13032);
nand U14259 (N_14259,N_13528,N_12793);
and U14260 (N_14260,N_12504,N_12571);
nor U14261 (N_14261,N_12614,N_12669);
and U14262 (N_14262,N_13517,N_12573);
and U14263 (N_14263,N_13503,N_13541);
xnor U14264 (N_14264,N_13281,N_13592);
and U14265 (N_14265,N_12840,N_12532);
nor U14266 (N_14266,N_13224,N_13706);
or U14267 (N_14267,N_12901,N_13196);
nor U14268 (N_14268,N_13680,N_13274);
or U14269 (N_14269,N_12533,N_12936);
and U14270 (N_14270,N_12779,N_13214);
xnor U14271 (N_14271,N_12933,N_13472);
and U14272 (N_14272,N_12923,N_13218);
nor U14273 (N_14273,N_12974,N_13693);
nor U14274 (N_14274,N_13333,N_12961);
or U14275 (N_14275,N_12646,N_12566);
or U14276 (N_14276,N_13189,N_13666);
nor U14277 (N_14277,N_13090,N_13726);
and U14278 (N_14278,N_13657,N_13219);
xor U14279 (N_14279,N_13056,N_12621);
nor U14280 (N_14280,N_13653,N_13729);
nand U14281 (N_14281,N_13408,N_13446);
nand U14282 (N_14282,N_13216,N_13073);
or U14283 (N_14283,N_13565,N_12711);
nand U14284 (N_14284,N_12743,N_13171);
nor U14285 (N_14285,N_12712,N_13627);
nand U14286 (N_14286,N_13033,N_13210);
nand U14287 (N_14287,N_13229,N_13103);
and U14288 (N_14288,N_13198,N_13004);
xnor U14289 (N_14289,N_12865,N_13364);
or U14290 (N_14290,N_13086,N_13438);
nor U14291 (N_14291,N_12592,N_13606);
nor U14292 (N_14292,N_13195,N_13549);
xor U14293 (N_14293,N_13211,N_13102);
nand U14294 (N_14294,N_13749,N_13489);
nand U14295 (N_14295,N_12731,N_13480);
nor U14296 (N_14296,N_12741,N_13003);
and U14297 (N_14297,N_13671,N_13279);
or U14298 (N_14298,N_13176,N_13237);
and U14299 (N_14299,N_13632,N_13688);
or U14300 (N_14300,N_12745,N_13011);
and U14301 (N_14301,N_13628,N_13424);
and U14302 (N_14302,N_12917,N_12808);
xnor U14303 (N_14303,N_12502,N_12558);
and U14304 (N_14304,N_13728,N_13107);
xor U14305 (N_14305,N_12560,N_12506);
nand U14306 (N_14306,N_13223,N_12989);
nand U14307 (N_14307,N_13338,N_13146);
or U14308 (N_14308,N_12922,N_12615);
nor U14309 (N_14309,N_13579,N_13123);
or U14310 (N_14310,N_12691,N_13718);
nand U14311 (N_14311,N_13715,N_13026);
and U14312 (N_14312,N_13067,N_13526);
nand U14313 (N_14313,N_12734,N_12796);
nand U14314 (N_14314,N_12938,N_12519);
xor U14315 (N_14315,N_13616,N_13527);
nor U14316 (N_14316,N_12509,N_12778);
nor U14317 (N_14317,N_13574,N_12806);
nor U14318 (N_14318,N_13088,N_13289);
nor U14319 (N_14319,N_13117,N_12627);
or U14320 (N_14320,N_12636,N_12889);
or U14321 (N_14321,N_12679,N_13137);
and U14322 (N_14322,N_13385,N_13231);
nand U14323 (N_14323,N_13121,N_12582);
nand U14324 (N_14324,N_12832,N_13559);
nand U14325 (N_14325,N_13136,N_13611);
nor U14326 (N_14326,N_12512,N_13449);
and U14327 (N_14327,N_13048,N_12816);
nand U14328 (N_14328,N_13476,N_12951);
xnor U14329 (N_14329,N_12548,N_12813);
xnor U14330 (N_14330,N_13212,N_13699);
or U14331 (N_14331,N_13708,N_13419);
or U14332 (N_14332,N_13138,N_13386);
and U14333 (N_14333,N_12748,N_13672);
xor U14334 (N_14334,N_12841,N_13684);
and U14335 (N_14335,N_12723,N_13618);
or U14336 (N_14336,N_12888,N_12789);
nand U14337 (N_14337,N_13221,N_13514);
nor U14338 (N_14338,N_13698,N_13330);
and U14339 (N_14339,N_12962,N_13692);
nor U14340 (N_14340,N_13271,N_12902);
or U14341 (N_14341,N_13045,N_13571);
or U14342 (N_14342,N_13580,N_12605);
nor U14343 (N_14343,N_13701,N_13723);
nor U14344 (N_14344,N_12702,N_12835);
nor U14345 (N_14345,N_13605,N_13318);
and U14346 (N_14346,N_13095,N_13125);
and U14347 (N_14347,N_13109,N_13696);
nor U14348 (N_14348,N_13400,N_13131);
and U14349 (N_14349,N_12772,N_12733);
or U14350 (N_14350,N_13603,N_13373);
and U14351 (N_14351,N_13100,N_13686);
nand U14352 (N_14352,N_13725,N_13265);
nand U14353 (N_14353,N_13341,N_13037);
and U14354 (N_14354,N_13560,N_13148);
nor U14355 (N_14355,N_13597,N_13021);
nand U14356 (N_14356,N_13186,N_13082);
or U14357 (N_14357,N_13536,N_12897);
nor U14358 (N_14358,N_12673,N_13260);
nor U14359 (N_14359,N_13007,N_12609);
nor U14360 (N_14360,N_13532,N_12622);
nand U14361 (N_14361,N_13241,N_12871);
or U14362 (N_14362,N_12996,N_13681);
or U14363 (N_14363,N_13553,N_13213);
nand U14364 (N_14364,N_12613,N_13334);
and U14365 (N_14365,N_13093,N_13286);
and U14366 (N_14366,N_13747,N_12853);
nand U14367 (N_14367,N_13342,N_13162);
xor U14368 (N_14368,N_13311,N_12525);
nor U14369 (N_14369,N_13738,N_13302);
nor U14370 (N_14370,N_12680,N_13484);
or U14371 (N_14371,N_12737,N_13531);
and U14372 (N_14372,N_13156,N_13024);
nand U14373 (N_14373,N_13741,N_12904);
nor U14374 (N_14374,N_13744,N_12671);
or U14375 (N_14375,N_13333,N_13497);
nor U14376 (N_14376,N_13711,N_12924);
nand U14377 (N_14377,N_13093,N_13699);
or U14378 (N_14378,N_13045,N_12874);
nor U14379 (N_14379,N_12964,N_13272);
xnor U14380 (N_14380,N_13063,N_13094);
nor U14381 (N_14381,N_12690,N_12898);
nand U14382 (N_14382,N_13476,N_12582);
nand U14383 (N_14383,N_13700,N_13368);
xnor U14384 (N_14384,N_12692,N_13155);
and U14385 (N_14385,N_13679,N_13505);
nand U14386 (N_14386,N_13411,N_13434);
xnor U14387 (N_14387,N_13332,N_13354);
nor U14388 (N_14388,N_12718,N_12912);
or U14389 (N_14389,N_13445,N_13335);
or U14390 (N_14390,N_13096,N_13399);
xor U14391 (N_14391,N_12634,N_13582);
xor U14392 (N_14392,N_13296,N_13088);
nand U14393 (N_14393,N_12975,N_12929);
or U14394 (N_14394,N_13292,N_12699);
and U14395 (N_14395,N_13012,N_12773);
or U14396 (N_14396,N_12610,N_13355);
nor U14397 (N_14397,N_13251,N_12573);
xnor U14398 (N_14398,N_13450,N_12794);
or U14399 (N_14399,N_12675,N_13318);
nand U14400 (N_14400,N_13028,N_12818);
nand U14401 (N_14401,N_13735,N_13030);
and U14402 (N_14402,N_13585,N_13028);
or U14403 (N_14403,N_13090,N_13002);
xnor U14404 (N_14404,N_13601,N_12735);
and U14405 (N_14405,N_13181,N_13051);
nand U14406 (N_14406,N_12510,N_12955);
nor U14407 (N_14407,N_13360,N_12573);
xor U14408 (N_14408,N_12832,N_13451);
or U14409 (N_14409,N_12844,N_12603);
nor U14410 (N_14410,N_13540,N_13741);
nand U14411 (N_14411,N_13525,N_13041);
and U14412 (N_14412,N_12578,N_13091);
or U14413 (N_14413,N_13015,N_12903);
or U14414 (N_14414,N_12819,N_12567);
or U14415 (N_14415,N_13707,N_12840);
nor U14416 (N_14416,N_13146,N_12748);
nor U14417 (N_14417,N_12844,N_12738);
nand U14418 (N_14418,N_13328,N_13118);
and U14419 (N_14419,N_13094,N_13202);
or U14420 (N_14420,N_13738,N_13160);
nor U14421 (N_14421,N_13391,N_12803);
xnor U14422 (N_14422,N_13326,N_13140);
or U14423 (N_14423,N_12559,N_13205);
xor U14424 (N_14424,N_13078,N_13456);
and U14425 (N_14425,N_12788,N_13525);
and U14426 (N_14426,N_13061,N_13065);
xor U14427 (N_14427,N_13708,N_12555);
xor U14428 (N_14428,N_13221,N_13206);
and U14429 (N_14429,N_13255,N_13421);
nor U14430 (N_14430,N_12739,N_13729);
and U14431 (N_14431,N_12928,N_13232);
or U14432 (N_14432,N_13501,N_13265);
or U14433 (N_14433,N_12566,N_13667);
nor U14434 (N_14434,N_12595,N_13253);
xor U14435 (N_14435,N_13104,N_12600);
and U14436 (N_14436,N_13055,N_13458);
xor U14437 (N_14437,N_13641,N_13387);
or U14438 (N_14438,N_13118,N_13145);
xnor U14439 (N_14439,N_13607,N_13693);
and U14440 (N_14440,N_12988,N_12956);
nor U14441 (N_14441,N_12708,N_13740);
or U14442 (N_14442,N_12809,N_13562);
xnor U14443 (N_14443,N_13733,N_13049);
and U14444 (N_14444,N_13149,N_13164);
xor U14445 (N_14445,N_13747,N_12969);
xnor U14446 (N_14446,N_12869,N_13738);
nand U14447 (N_14447,N_12998,N_13118);
or U14448 (N_14448,N_13027,N_13357);
nand U14449 (N_14449,N_13539,N_12942);
nor U14450 (N_14450,N_13658,N_13233);
or U14451 (N_14451,N_13672,N_12572);
xor U14452 (N_14452,N_13667,N_13175);
nand U14453 (N_14453,N_13721,N_12959);
and U14454 (N_14454,N_12634,N_13739);
nand U14455 (N_14455,N_12700,N_13275);
and U14456 (N_14456,N_13662,N_13691);
xor U14457 (N_14457,N_13339,N_12548);
nor U14458 (N_14458,N_13701,N_12529);
and U14459 (N_14459,N_12771,N_12677);
and U14460 (N_14460,N_13117,N_13434);
nor U14461 (N_14461,N_12808,N_12955);
xor U14462 (N_14462,N_12842,N_12663);
nand U14463 (N_14463,N_13556,N_12798);
nand U14464 (N_14464,N_13718,N_12579);
nand U14465 (N_14465,N_13711,N_12983);
nand U14466 (N_14466,N_13374,N_13478);
xnor U14467 (N_14467,N_12907,N_13596);
nand U14468 (N_14468,N_12743,N_13436);
nor U14469 (N_14469,N_13384,N_13557);
nor U14470 (N_14470,N_12792,N_13188);
and U14471 (N_14471,N_12924,N_12911);
xnor U14472 (N_14472,N_13122,N_13081);
or U14473 (N_14473,N_12742,N_12521);
and U14474 (N_14474,N_12835,N_12940);
nor U14475 (N_14475,N_12833,N_13366);
xor U14476 (N_14476,N_12657,N_13329);
or U14477 (N_14477,N_12855,N_13592);
nand U14478 (N_14478,N_13158,N_13493);
or U14479 (N_14479,N_13663,N_12745);
nor U14480 (N_14480,N_12720,N_12562);
and U14481 (N_14481,N_13636,N_12945);
or U14482 (N_14482,N_13387,N_13252);
nand U14483 (N_14483,N_13198,N_12914);
xnor U14484 (N_14484,N_13254,N_13628);
nor U14485 (N_14485,N_13176,N_12777);
nand U14486 (N_14486,N_12826,N_12806);
nand U14487 (N_14487,N_13148,N_12973);
nor U14488 (N_14488,N_12768,N_12754);
and U14489 (N_14489,N_13140,N_12573);
nand U14490 (N_14490,N_13104,N_13614);
xor U14491 (N_14491,N_12662,N_12734);
and U14492 (N_14492,N_12908,N_12503);
nor U14493 (N_14493,N_13700,N_13433);
or U14494 (N_14494,N_12554,N_12807);
and U14495 (N_14495,N_12897,N_13349);
xnor U14496 (N_14496,N_12571,N_12558);
nand U14497 (N_14497,N_12900,N_13251);
nand U14498 (N_14498,N_12693,N_13072);
nand U14499 (N_14499,N_13183,N_13046);
and U14500 (N_14500,N_13379,N_12598);
nand U14501 (N_14501,N_13357,N_12659);
or U14502 (N_14502,N_13643,N_13145);
xor U14503 (N_14503,N_13738,N_12621);
xor U14504 (N_14504,N_13306,N_12721);
nand U14505 (N_14505,N_13462,N_12936);
nor U14506 (N_14506,N_12522,N_12925);
or U14507 (N_14507,N_13569,N_13317);
xor U14508 (N_14508,N_12552,N_13014);
nor U14509 (N_14509,N_12932,N_13266);
nor U14510 (N_14510,N_13082,N_12571);
nor U14511 (N_14511,N_12549,N_12751);
nor U14512 (N_14512,N_13700,N_12896);
nor U14513 (N_14513,N_12727,N_13205);
or U14514 (N_14514,N_12918,N_13660);
xnor U14515 (N_14515,N_13611,N_12845);
nor U14516 (N_14516,N_13228,N_12896);
nand U14517 (N_14517,N_13551,N_13524);
and U14518 (N_14518,N_12762,N_13269);
and U14519 (N_14519,N_12731,N_13472);
or U14520 (N_14520,N_12935,N_13259);
or U14521 (N_14521,N_13057,N_13455);
and U14522 (N_14522,N_12818,N_13443);
and U14523 (N_14523,N_13618,N_13511);
nand U14524 (N_14524,N_12697,N_13203);
and U14525 (N_14525,N_13227,N_13186);
nor U14526 (N_14526,N_13288,N_13066);
xor U14527 (N_14527,N_13721,N_12778);
or U14528 (N_14528,N_12885,N_13474);
nor U14529 (N_14529,N_12880,N_13617);
nor U14530 (N_14530,N_13310,N_13048);
nand U14531 (N_14531,N_12966,N_13743);
nor U14532 (N_14532,N_12571,N_13573);
or U14533 (N_14533,N_13032,N_13134);
or U14534 (N_14534,N_13420,N_12902);
and U14535 (N_14535,N_13160,N_12722);
and U14536 (N_14536,N_12850,N_12979);
or U14537 (N_14537,N_13553,N_13570);
nand U14538 (N_14538,N_12947,N_12544);
and U14539 (N_14539,N_12762,N_13452);
xor U14540 (N_14540,N_12922,N_12770);
or U14541 (N_14541,N_13582,N_13649);
or U14542 (N_14542,N_12955,N_13325);
xor U14543 (N_14543,N_13478,N_13260);
xor U14544 (N_14544,N_13269,N_13161);
or U14545 (N_14545,N_12617,N_13216);
xnor U14546 (N_14546,N_13044,N_12866);
nand U14547 (N_14547,N_13444,N_13636);
or U14548 (N_14548,N_12614,N_12794);
and U14549 (N_14549,N_12811,N_12624);
or U14550 (N_14550,N_12914,N_13410);
nor U14551 (N_14551,N_12877,N_12647);
nor U14552 (N_14552,N_13405,N_13184);
nor U14553 (N_14553,N_13490,N_13328);
xnor U14554 (N_14554,N_13349,N_12641);
and U14555 (N_14555,N_13173,N_12847);
nand U14556 (N_14556,N_12854,N_12712);
or U14557 (N_14557,N_13041,N_12619);
nor U14558 (N_14558,N_13349,N_13619);
xor U14559 (N_14559,N_12813,N_12895);
nor U14560 (N_14560,N_13232,N_13002);
xor U14561 (N_14561,N_12981,N_12813);
xor U14562 (N_14562,N_13221,N_12903);
xor U14563 (N_14563,N_13610,N_12930);
and U14564 (N_14564,N_13467,N_12526);
nand U14565 (N_14565,N_13378,N_13640);
and U14566 (N_14566,N_12555,N_12886);
and U14567 (N_14567,N_12829,N_13210);
xnor U14568 (N_14568,N_13183,N_13085);
and U14569 (N_14569,N_12953,N_13127);
xor U14570 (N_14570,N_13453,N_12804);
xor U14571 (N_14571,N_13624,N_13052);
xnor U14572 (N_14572,N_12893,N_13098);
xor U14573 (N_14573,N_12917,N_13180);
or U14574 (N_14574,N_13451,N_13102);
nand U14575 (N_14575,N_13413,N_12957);
or U14576 (N_14576,N_13586,N_12765);
xnor U14577 (N_14577,N_12773,N_13320);
xor U14578 (N_14578,N_12917,N_12554);
nand U14579 (N_14579,N_12639,N_13462);
or U14580 (N_14580,N_13275,N_13307);
or U14581 (N_14581,N_13180,N_12884);
and U14582 (N_14582,N_12818,N_13174);
and U14583 (N_14583,N_13696,N_13532);
xor U14584 (N_14584,N_12741,N_12678);
nand U14585 (N_14585,N_12542,N_12715);
xnor U14586 (N_14586,N_13488,N_13160);
nand U14587 (N_14587,N_13488,N_12870);
nand U14588 (N_14588,N_13390,N_13315);
and U14589 (N_14589,N_12704,N_12895);
xor U14590 (N_14590,N_13076,N_13747);
or U14591 (N_14591,N_13487,N_12823);
nor U14592 (N_14592,N_12787,N_13661);
or U14593 (N_14593,N_13420,N_13724);
and U14594 (N_14594,N_12639,N_13132);
nand U14595 (N_14595,N_12957,N_12861);
nand U14596 (N_14596,N_13725,N_13544);
or U14597 (N_14597,N_13062,N_13588);
nand U14598 (N_14598,N_12647,N_13018);
and U14599 (N_14599,N_12631,N_12523);
nor U14600 (N_14600,N_12579,N_12803);
nor U14601 (N_14601,N_13656,N_12810);
or U14602 (N_14602,N_12606,N_13524);
nand U14603 (N_14603,N_12524,N_13462);
nand U14604 (N_14604,N_12863,N_13459);
and U14605 (N_14605,N_12882,N_12514);
and U14606 (N_14606,N_13334,N_13689);
and U14607 (N_14607,N_12939,N_13555);
nor U14608 (N_14608,N_13059,N_13519);
or U14609 (N_14609,N_12702,N_12991);
nor U14610 (N_14610,N_13459,N_13566);
or U14611 (N_14611,N_12574,N_12649);
nand U14612 (N_14612,N_13467,N_13569);
nand U14613 (N_14613,N_13473,N_13422);
xnor U14614 (N_14614,N_12810,N_13001);
nand U14615 (N_14615,N_13015,N_13647);
nand U14616 (N_14616,N_12998,N_12711);
nor U14617 (N_14617,N_12903,N_12518);
xor U14618 (N_14618,N_12621,N_12866);
xnor U14619 (N_14619,N_13442,N_12813);
or U14620 (N_14620,N_13532,N_13638);
nand U14621 (N_14621,N_13179,N_13429);
nor U14622 (N_14622,N_12778,N_13002);
and U14623 (N_14623,N_12886,N_12595);
nor U14624 (N_14624,N_13164,N_13443);
nand U14625 (N_14625,N_13693,N_12571);
nor U14626 (N_14626,N_13439,N_12857);
xor U14627 (N_14627,N_13574,N_12718);
or U14628 (N_14628,N_12788,N_13512);
and U14629 (N_14629,N_13295,N_12525);
or U14630 (N_14630,N_12822,N_13665);
and U14631 (N_14631,N_13716,N_13038);
nand U14632 (N_14632,N_12670,N_12504);
or U14633 (N_14633,N_13008,N_12705);
and U14634 (N_14634,N_13651,N_12953);
nor U14635 (N_14635,N_12546,N_13661);
nand U14636 (N_14636,N_12655,N_13330);
and U14637 (N_14637,N_13127,N_12729);
nand U14638 (N_14638,N_13425,N_13126);
nand U14639 (N_14639,N_13269,N_13699);
nand U14640 (N_14640,N_13025,N_12622);
nor U14641 (N_14641,N_12912,N_12709);
xor U14642 (N_14642,N_12606,N_13348);
nand U14643 (N_14643,N_13612,N_13394);
and U14644 (N_14644,N_12639,N_12985);
or U14645 (N_14645,N_13723,N_12790);
or U14646 (N_14646,N_13468,N_13277);
nor U14647 (N_14647,N_13435,N_13456);
xnor U14648 (N_14648,N_12696,N_13349);
xor U14649 (N_14649,N_13219,N_13590);
or U14650 (N_14650,N_12812,N_13124);
nor U14651 (N_14651,N_12952,N_13530);
or U14652 (N_14652,N_13417,N_13164);
nand U14653 (N_14653,N_12864,N_13258);
xnor U14654 (N_14654,N_12548,N_12883);
xnor U14655 (N_14655,N_13429,N_12539);
nand U14656 (N_14656,N_12519,N_13360);
xnor U14657 (N_14657,N_13042,N_12954);
and U14658 (N_14658,N_13416,N_12729);
xnor U14659 (N_14659,N_12513,N_13649);
nor U14660 (N_14660,N_12808,N_13007);
nand U14661 (N_14661,N_13049,N_13487);
and U14662 (N_14662,N_13737,N_13067);
nor U14663 (N_14663,N_12907,N_13328);
and U14664 (N_14664,N_13399,N_13161);
and U14665 (N_14665,N_13031,N_13044);
or U14666 (N_14666,N_13037,N_13301);
or U14667 (N_14667,N_12895,N_13533);
nand U14668 (N_14668,N_12842,N_13257);
nand U14669 (N_14669,N_13525,N_13690);
nand U14670 (N_14670,N_12633,N_12803);
and U14671 (N_14671,N_13527,N_12737);
nor U14672 (N_14672,N_13576,N_13544);
xnor U14673 (N_14673,N_12704,N_12799);
nor U14674 (N_14674,N_13574,N_12905);
nand U14675 (N_14675,N_12877,N_13107);
or U14676 (N_14676,N_13605,N_13216);
nor U14677 (N_14677,N_13500,N_13022);
xor U14678 (N_14678,N_12978,N_13661);
or U14679 (N_14679,N_12610,N_12705);
or U14680 (N_14680,N_12608,N_13178);
nor U14681 (N_14681,N_13130,N_12656);
nor U14682 (N_14682,N_12949,N_13528);
nor U14683 (N_14683,N_13332,N_13365);
or U14684 (N_14684,N_12962,N_13114);
nand U14685 (N_14685,N_13739,N_13555);
xor U14686 (N_14686,N_13199,N_12655);
nor U14687 (N_14687,N_12836,N_13410);
nor U14688 (N_14688,N_13481,N_13525);
or U14689 (N_14689,N_13018,N_13432);
and U14690 (N_14690,N_13698,N_12534);
or U14691 (N_14691,N_12871,N_13665);
nand U14692 (N_14692,N_12624,N_12982);
nand U14693 (N_14693,N_13447,N_13087);
nor U14694 (N_14694,N_13331,N_12787);
or U14695 (N_14695,N_13175,N_13357);
xor U14696 (N_14696,N_13670,N_12667);
xor U14697 (N_14697,N_13429,N_13530);
nor U14698 (N_14698,N_13231,N_13255);
nor U14699 (N_14699,N_13468,N_13401);
nor U14700 (N_14700,N_13339,N_13527);
and U14701 (N_14701,N_12516,N_12812);
or U14702 (N_14702,N_12788,N_12547);
and U14703 (N_14703,N_12604,N_13244);
or U14704 (N_14704,N_12665,N_13568);
nor U14705 (N_14705,N_13246,N_12662);
or U14706 (N_14706,N_13170,N_12677);
or U14707 (N_14707,N_13728,N_13018);
nand U14708 (N_14708,N_12894,N_13723);
and U14709 (N_14709,N_12861,N_13240);
nor U14710 (N_14710,N_12704,N_13608);
xor U14711 (N_14711,N_13036,N_12998);
or U14712 (N_14712,N_12738,N_12923);
xor U14713 (N_14713,N_12869,N_13260);
nand U14714 (N_14714,N_13048,N_12810);
xnor U14715 (N_14715,N_12800,N_13394);
or U14716 (N_14716,N_13135,N_13377);
xnor U14717 (N_14717,N_12856,N_13639);
or U14718 (N_14718,N_13533,N_13483);
and U14719 (N_14719,N_12777,N_13108);
and U14720 (N_14720,N_13134,N_13193);
xor U14721 (N_14721,N_13292,N_12638);
and U14722 (N_14722,N_13470,N_13685);
nand U14723 (N_14723,N_12519,N_12859);
nor U14724 (N_14724,N_13067,N_13301);
nor U14725 (N_14725,N_13052,N_13347);
and U14726 (N_14726,N_12675,N_13124);
xnor U14727 (N_14727,N_12893,N_12979);
or U14728 (N_14728,N_12613,N_13510);
nand U14729 (N_14729,N_13274,N_13223);
nor U14730 (N_14730,N_13059,N_12826);
or U14731 (N_14731,N_12761,N_13737);
xor U14732 (N_14732,N_12676,N_13444);
and U14733 (N_14733,N_13163,N_12752);
nor U14734 (N_14734,N_12738,N_13196);
nand U14735 (N_14735,N_13251,N_13525);
and U14736 (N_14736,N_13580,N_13239);
or U14737 (N_14737,N_12913,N_13022);
and U14738 (N_14738,N_12513,N_12658);
and U14739 (N_14739,N_13356,N_13387);
and U14740 (N_14740,N_13550,N_13206);
nor U14741 (N_14741,N_13639,N_13264);
nand U14742 (N_14742,N_13583,N_12663);
nand U14743 (N_14743,N_12878,N_12617);
nand U14744 (N_14744,N_13133,N_13458);
nor U14745 (N_14745,N_13211,N_12528);
nor U14746 (N_14746,N_12536,N_12602);
or U14747 (N_14747,N_13338,N_13620);
xor U14748 (N_14748,N_12580,N_13255);
nor U14749 (N_14749,N_12714,N_12876);
nand U14750 (N_14750,N_12867,N_12993);
or U14751 (N_14751,N_12834,N_12625);
nor U14752 (N_14752,N_13320,N_13381);
nand U14753 (N_14753,N_12708,N_13295);
nor U14754 (N_14754,N_13466,N_13322);
xor U14755 (N_14755,N_13045,N_13065);
nand U14756 (N_14756,N_12632,N_13239);
nor U14757 (N_14757,N_13165,N_13430);
xor U14758 (N_14758,N_13223,N_13245);
nor U14759 (N_14759,N_12520,N_12639);
nor U14760 (N_14760,N_13661,N_13360);
xnor U14761 (N_14761,N_13094,N_12723);
and U14762 (N_14762,N_13193,N_13518);
nor U14763 (N_14763,N_13035,N_12940);
xor U14764 (N_14764,N_13631,N_12986);
nor U14765 (N_14765,N_13121,N_12848);
or U14766 (N_14766,N_13179,N_13101);
or U14767 (N_14767,N_13616,N_13585);
nor U14768 (N_14768,N_13483,N_12920);
nor U14769 (N_14769,N_13257,N_12789);
nand U14770 (N_14770,N_13112,N_12513);
and U14771 (N_14771,N_12682,N_13470);
or U14772 (N_14772,N_12536,N_13471);
nand U14773 (N_14773,N_12886,N_13355);
and U14774 (N_14774,N_13717,N_13636);
nor U14775 (N_14775,N_13156,N_12779);
nand U14776 (N_14776,N_12963,N_12843);
or U14777 (N_14777,N_13095,N_13433);
nor U14778 (N_14778,N_13304,N_13588);
nand U14779 (N_14779,N_13659,N_13215);
nor U14780 (N_14780,N_13349,N_13524);
or U14781 (N_14781,N_13014,N_13507);
xor U14782 (N_14782,N_13507,N_12838);
nor U14783 (N_14783,N_12566,N_13320);
nor U14784 (N_14784,N_12618,N_13191);
nor U14785 (N_14785,N_13180,N_13304);
nand U14786 (N_14786,N_13379,N_13672);
or U14787 (N_14787,N_13692,N_13391);
xnor U14788 (N_14788,N_12883,N_12871);
xnor U14789 (N_14789,N_13595,N_13003);
nor U14790 (N_14790,N_13595,N_13550);
or U14791 (N_14791,N_13685,N_13594);
xnor U14792 (N_14792,N_12737,N_12985);
nor U14793 (N_14793,N_13562,N_13588);
or U14794 (N_14794,N_13746,N_13139);
or U14795 (N_14795,N_12931,N_13337);
xnor U14796 (N_14796,N_13365,N_12827);
or U14797 (N_14797,N_13613,N_13712);
nor U14798 (N_14798,N_12718,N_13475);
nand U14799 (N_14799,N_12916,N_13377);
nor U14800 (N_14800,N_13373,N_12911);
xnor U14801 (N_14801,N_13508,N_12922);
nor U14802 (N_14802,N_12802,N_13204);
and U14803 (N_14803,N_12906,N_13444);
nand U14804 (N_14804,N_13743,N_13618);
and U14805 (N_14805,N_12952,N_13178);
and U14806 (N_14806,N_12642,N_13117);
or U14807 (N_14807,N_13236,N_12817);
or U14808 (N_14808,N_12790,N_12733);
xnor U14809 (N_14809,N_12654,N_12877);
xor U14810 (N_14810,N_12983,N_13719);
and U14811 (N_14811,N_13360,N_12678);
xor U14812 (N_14812,N_12864,N_13264);
or U14813 (N_14813,N_13212,N_12570);
and U14814 (N_14814,N_12913,N_12583);
nand U14815 (N_14815,N_13271,N_12764);
nand U14816 (N_14816,N_13180,N_13040);
nor U14817 (N_14817,N_12823,N_13734);
nand U14818 (N_14818,N_13609,N_12676);
nand U14819 (N_14819,N_13679,N_13130);
and U14820 (N_14820,N_12900,N_12586);
xor U14821 (N_14821,N_12737,N_13393);
and U14822 (N_14822,N_13706,N_12893);
nand U14823 (N_14823,N_13104,N_12724);
and U14824 (N_14824,N_12892,N_12848);
nand U14825 (N_14825,N_13125,N_12693);
and U14826 (N_14826,N_13121,N_13042);
or U14827 (N_14827,N_13097,N_12926);
nor U14828 (N_14828,N_13679,N_13017);
nor U14829 (N_14829,N_12650,N_12608);
nand U14830 (N_14830,N_12702,N_13394);
and U14831 (N_14831,N_13163,N_12614);
or U14832 (N_14832,N_13205,N_12549);
nor U14833 (N_14833,N_13175,N_12651);
nor U14834 (N_14834,N_13526,N_12728);
and U14835 (N_14835,N_13191,N_12820);
and U14836 (N_14836,N_13149,N_12803);
nor U14837 (N_14837,N_13431,N_13149);
xnor U14838 (N_14838,N_13703,N_13396);
or U14839 (N_14839,N_12866,N_13420);
nand U14840 (N_14840,N_13284,N_13681);
nor U14841 (N_14841,N_13378,N_13337);
and U14842 (N_14842,N_13416,N_13685);
nor U14843 (N_14843,N_13213,N_12766);
xnor U14844 (N_14844,N_13626,N_12930);
and U14845 (N_14845,N_13115,N_12606);
nor U14846 (N_14846,N_12633,N_12814);
or U14847 (N_14847,N_13155,N_12795);
nand U14848 (N_14848,N_12675,N_13074);
and U14849 (N_14849,N_13527,N_12866);
nand U14850 (N_14850,N_13703,N_13685);
nor U14851 (N_14851,N_12955,N_12999);
and U14852 (N_14852,N_13165,N_12914);
nand U14853 (N_14853,N_13687,N_13458);
and U14854 (N_14854,N_13096,N_12588);
nor U14855 (N_14855,N_12986,N_12900);
nand U14856 (N_14856,N_12558,N_12643);
or U14857 (N_14857,N_13339,N_12906);
and U14858 (N_14858,N_13589,N_12629);
nor U14859 (N_14859,N_12512,N_13505);
and U14860 (N_14860,N_13695,N_13316);
xor U14861 (N_14861,N_12947,N_13181);
xor U14862 (N_14862,N_12836,N_13742);
xor U14863 (N_14863,N_12567,N_12517);
or U14864 (N_14864,N_13567,N_13400);
or U14865 (N_14865,N_12837,N_13099);
or U14866 (N_14866,N_13393,N_13650);
nand U14867 (N_14867,N_13715,N_13179);
xor U14868 (N_14868,N_13351,N_13388);
and U14869 (N_14869,N_13255,N_13415);
nand U14870 (N_14870,N_13256,N_12788);
nor U14871 (N_14871,N_13706,N_12988);
nand U14872 (N_14872,N_13742,N_12671);
nor U14873 (N_14873,N_13717,N_13625);
nand U14874 (N_14874,N_12894,N_12798);
nand U14875 (N_14875,N_13713,N_12617);
nand U14876 (N_14876,N_13609,N_13302);
or U14877 (N_14877,N_13090,N_12830);
nor U14878 (N_14878,N_13726,N_12672);
nand U14879 (N_14879,N_12760,N_13237);
nor U14880 (N_14880,N_12897,N_12920);
or U14881 (N_14881,N_13391,N_13244);
nor U14882 (N_14882,N_13329,N_13510);
nand U14883 (N_14883,N_13617,N_12521);
nand U14884 (N_14884,N_12957,N_13500);
or U14885 (N_14885,N_12738,N_12832);
xor U14886 (N_14886,N_12811,N_12736);
or U14887 (N_14887,N_13207,N_13498);
and U14888 (N_14888,N_12942,N_13304);
xor U14889 (N_14889,N_12522,N_13335);
xnor U14890 (N_14890,N_12880,N_13002);
xnor U14891 (N_14891,N_13596,N_12855);
and U14892 (N_14892,N_12730,N_13387);
xor U14893 (N_14893,N_12862,N_12828);
nor U14894 (N_14894,N_12601,N_13180);
or U14895 (N_14895,N_12927,N_12796);
nor U14896 (N_14896,N_13304,N_13607);
xor U14897 (N_14897,N_13468,N_12553);
xor U14898 (N_14898,N_13705,N_13463);
nor U14899 (N_14899,N_13480,N_12505);
xnor U14900 (N_14900,N_12574,N_12875);
and U14901 (N_14901,N_12771,N_13331);
nand U14902 (N_14902,N_12904,N_12501);
nor U14903 (N_14903,N_13493,N_12970);
xor U14904 (N_14904,N_13680,N_13157);
nor U14905 (N_14905,N_13533,N_13622);
nand U14906 (N_14906,N_12619,N_13579);
and U14907 (N_14907,N_12798,N_13335);
xnor U14908 (N_14908,N_13554,N_13699);
or U14909 (N_14909,N_12779,N_13600);
xor U14910 (N_14910,N_13252,N_13433);
or U14911 (N_14911,N_13145,N_13383);
and U14912 (N_14912,N_12817,N_12753);
and U14913 (N_14913,N_12626,N_13606);
nand U14914 (N_14914,N_13006,N_12902);
or U14915 (N_14915,N_13115,N_13468);
xnor U14916 (N_14916,N_12828,N_13582);
and U14917 (N_14917,N_13684,N_13147);
nand U14918 (N_14918,N_12840,N_13646);
xor U14919 (N_14919,N_13495,N_12694);
or U14920 (N_14920,N_13219,N_13163);
nand U14921 (N_14921,N_13038,N_12722);
nor U14922 (N_14922,N_12509,N_13097);
xor U14923 (N_14923,N_12998,N_13346);
and U14924 (N_14924,N_13065,N_12572);
or U14925 (N_14925,N_13536,N_12514);
nand U14926 (N_14926,N_13278,N_12709);
or U14927 (N_14927,N_13430,N_13692);
xnor U14928 (N_14928,N_13158,N_13002);
xor U14929 (N_14929,N_13692,N_13612);
nor U14930 (N_14930,N_12987,N_13629);
xor U14931 (N_14931,N_13324,N_13738);
nand U14932 (N_14932,N_12958,N_12620);
nor U14933 (N_14933,N_13640,N_12779);
or U14934 (N_14934,N_13651,N_13229);
xnor U14935 (N_14935,N_12866,N_13191);
and U14936 (N_14936,N_12783,N_12599);
nand U14937 (N_14937,N_13445,N_13073);
nand U14938 (N_14938,N_13336,N_13485);
nand U14939 (N_14939,N_12790,N_13558);
nand U14940 (N_14940,N_12606,N_12689);
nor U14941 (N_14941,N_12855,N_13394);
nor U14942 (N_14942,N_12886,N_12924);
nand U14943 (N_14943,N_13444,N_12808);
nand U14944 (N_14944,N_13660,N_13189);
xor U14945 (N_14945,N_12673,N_13473);
nor U14946 (N_14946,N_13356,N_13110);
and U14947 (N_14947,N_13425,N_12776);
nand U14948 (N_14948,N_13458,N_13214);
and U14949 (N_14949,N_12794,N_13038);
and U14950 (N_14950,N_12904,N_13365);
xnor U14951 (N_14951,N_12601,N_13376);
xnor U14952 (N_14952,N_13306,N_13210);
nor U14953 (N_14953,N_13520,N_13459);
and U14954 (N_14954,N_13363,N_13161);
or U14955 (N_14955,N_13026,N_13305);
nand U14956 (N_14956,N_13524,N_12533);
or U14957 (N_14957,N_12783,N_13738);
nor U14958 (N_14958,N_13026,N_12709);
nor U14959 (N_14959,N_13612,N_12637);
or U14960 (N_14960,N_13530,N_12549);
or U14961 (N_14961,N_13254,N_13531);
nor U14962 (N_14962,N_13493,N_13556);
nor U14963 (N_14963,N_13218,N_12848);
xor U14964 (N_14964,N_12667,N_13533);
and U14965 (N_14965,N_12761,N_13491);
and U14966 (N_14966,N_13725,N_12847);
or U14967 (N_14967,N_13707,N_12707);
or U14968 (N_14968,N_13677,N_13099);
and U14969 (N_14969,N_12756,N_13558);
and U14970 (N_14970,N_13047,N_13455);
nand U14971 (N_14971,N_12618,N_13337);
nor U14972 (N_14972,N_13543,N_12547);
nand U14973 (N_14973,N_12941,N_12549);
and U14974 (N_14974,N_12871,N_13313);
xnor U14975 (N_14975,N_12505,N_13692);
and U14976 (N_14976,N_12943,N_12709);
nor U14977 (N_14977,N_13435,N_13749);
nand U14978 (N_14978,N_13548,N_12846);
and U14979 (N_14979,N_12983,N_13740);
nand U14980 (N_14980,N_13365,N_13677);
or U14981 (N_14981,N_13043,N_12747);
or U14982 (N_14982,N_13706,N_13415);
nand U14983 (N_14983,N_13533,N_12793);
or U14984 (N_14984,N_13525,N_13153);
or U14985 (N_14985,N_12949,N_13443);
and U14986 (N_14986,N_13167,N_13620);
and U14987 (N_14987,N_13640,N_12921);
and U14988 (N_14988,N_13440,N_12932);
nand U14989 (N_14989,N_12561,N_13394);
nor U14990 (N_14990,N_12683,N_12655);
nand U14991 (N_14991,N_12858,N_12911);
xnor U14992 (N_14992,N_13635,N_12634);
xor U14993 (N_14993,N_13722,N_13550);
nor U14994 (N_14994,N_13121,N_13487);
xor U14995 (N_14995,N_12843,N_12686);
nand U14996 (N_14996,N_13451,N_13448);
and U14997 (N_14997,N_13284,N_13027);
nor U14998 (N_14998,N_12695,N_13199);
nand U14999 (N_14999,N_13581,N_13110);
nand U15000 (N_15000,N_14304,N_14802);
xor U15001 (N_15001,N_14529,N_14643);
nor U15002 (N_15002,N_13820,N_14476);
nand U15003 (N_15003,N_14932,N_14846);
nor U15004 (N_15004,N_14160,N_14603);
xor U15005 (N_15005,N_14791,N_14209);
and U15006 (N_15006,N_14179,N_14089);
xor U15007 (N_15007,N_14213,N_13999);
xor U15008 (N_15008,N_13787,N_14579);
or U15009 (N_15009,N_14972,N_14036);
and U15010 (N_15010,N_14428,N_14748);
nor U15011 (N_15011,N_14020,N_14436);
and U15012 (N_15012,N_13961,N_14946);
xnor U15013 (N_15013,N_14597,N_14426);
nand U15014 (N_15014,N_14726,N_14374);
or U15015 (N_15015,N_14134,N_14687);
nor U15016 (N_15016,N_14698,N_14188);
nand U15017 (N_15017,N_14879,N_13895);
and U15018 (N_15018,N_14614,N_13764);
nand U15019 (N_15019,N_14083,N_14752);
xor U15020 (N_15020,N_14014,N_14002);
nor U15021 (N_15021,N_13831,N_14445);
nor U15022 (N_15022,N_14300,N_13914);
and U15023 (N_15023,N_14427,N_14666);
nand U15024 (N_15024,N_14238,N_14406);
nand U15025 (N_15025,N_14017,N_14654);
and U15026 (N_15026,N_14249,N_13942);
or U15027 (N_15027,N_14039,N_14977);
xnor U15028 (N_15028,N_14743,N_13751);
and U15029 (N_15029,N_14463,N_14389);
xnor U15030 (N_15030,N_13958,N_14670);
nor U15031 (N_15031,N_14561,N_14208);
or U15032 (N_15032,N_14587,N_14874);
xor U15033 (N_15033,N_14660,N_14093);
nand U15034 (N_15034,N_14585,N_14868);
nand U15035 (N_15035,N_14661,N_13985);
nand U15036 (N_15036,N_13841,N_13889);
nand U15037 (N_15037,N_14756,N_14404);
or U15038 (N_15038,N_13983,N_14328);
nor U15039 (N_15039,N_14184,N_14609);
or U15040 (N_15040,N_14566,N_14187);
nand U15041 (N_15041,N_14851,N_14363);
or U15042 (N_15042,N_14196,N_14120);
nor U15043 (N_15043,N_14469,N_14254);
xor U15044 (N_15044,N_14084,N_14466);
nor U15045 (N_15045,N_14430,N_14984);
xnor U15046 (N_15046,N_14700,N_14556);
nor U15047 (N_15047,N_14057,N_14728);
or U15048 (N_15048,N_14681,N_14736);
nand U15049 (N_15049,N_14560,N_13995);
nor U15050 (N_15050,N_13778,N_14907);
xor U15051 (N_15051,N_14147,N_13872);
nand U15052 (N_15052,N_13753,N_14702);
nand U15053 (N_15053,N_13941,N_14313);
and U15054 (N_15054,N_13801,N_14200);
nand U15055 (N_15055,N_14862,N_13869);
xor U15056 (N_15056,N_14491,N_14803);
or U15057 (N_15057,N_14858,N_14572);
and U15058 (N_15058,N_14709,N_14864);
or U15059 (N_15059,N_13975,N_14853);
xnor U15060 (N_15060,N_14598,N_14279);
nor U15061 (N_15061,N_13808,N_14462);
xor U15062 (N_15062,N_14171,N_13885);
nor U15063 (N_15063,N_14873,N_14575);
xor U15064 (N_15064,N_14206,N_14344);
or U15065 (N_15065,N_13913,N_14633);
nor U15066 (N_15066,N_14338,N_13892);
xor U15067 (N_15067,N_13937,N_13911);
nand U15068 (N_15068,N_13828,N_14302);
and U15069 (N_15069,N_14408,N_14896);
and U15070 (N_15070,N_14886,N_14353);
or U15071 (N_15071,N_14980,N_14753);
nand U15072 (N_15072,N_13873,N_14016);
nand U15073 (N_15073,N_14034,N_14659);
or U15074 (N_15074,N_14905,N_14174);
nand U15075 (N_15075,N_14773,N_14554);
and U15076 (N_15076,N_14190,N_14033);
or U15077 (N_15077,N_13994,N_14453);
and U15078 (N_15078,N_14382,N_14695);
xnor U15079 (N_15079,N_14314,N_14674);
or U15080 (N_15080,N_14251,N_14100);
and U15081 (N_15081,N_14724,N_14964);
xnor U15082 (N_15082,N_14267,N_14876);
or U15083 (N_15083,N_14336,N_14895);
and U15084 (N_15084,N_14844,N_14899);
nor U15085 (N_15085,N_14542,N_14216);
or U15086 (N_15086,N_14000,N_13771);
nand U15087 (N_15087,N_14103,N_13943);
nor U15088 (N_15088,N_14278,N_14757);
nor U15089 (N_15089,N_14318,N_14523);
xnor U15090 (N_15090,N_14717,N_14348);
or U15091 (N_15091,N_14001,N_14524);
or U15092 (N_15092,N_14506,N_14589);
or U15093 (N_15093,N_14533,N_13815);
or U15094 (N_15094,N_13905,N_14013);
xnor U15095 (N_15095,N_14857,N_14845);
nand U15096 (N_15096,N_14418,N_13978);
nand U15097 (N_15097,N_14644,N_14971);
nor U15098 (N_15098,N_14714,N_14610);
nor U15099 (N_15099,N_14085,N_14168);
and U15100 (N_15100,N_14619,N_14559);
and U15101 (N_15101,N_13916,N_13891);
nand U15102 (N_15102,N_14118,N_14394);
or U15103 (N_15103,N_14230,N_14163);
and U15104 (N_15104,N_14543,N_14782);
or U15105 (N_15105,N_14326,N_14343);
xor U15106 (N_15106,N_14499,N_14412);
xnor U15107 (N_15107,N_13923,N_13982);
nor U15108 (N_15108,N_14961,N_14958);
nand U15109 (N_15109,N_14805,N_13996);
or U15110 (N_15110,N_14825,N_14970);
nor U15111 (N_15111,N_14903,N_14357);
nor U15112 (N_15112,N_14552,N_14890);
nor U15113 (N_15113,N_14226,N_14535);
nand U15114 (N_15114,N_14119,N_14071);
or U15115 (N_15115,N_14191,N_14095);
and U15116 (N_15116,N_14983,N_13966);
or U15117 (N_15117,N_13962,N_14305);
and U15118 (N_15118,N_14117,N_13919);
or U15119 (N_15119,N_14411,N_14078);
and U15120 (N_15120,N_14833,N_13785);
and U15121 (N_15121,N_14451,N_13921);
nor U15122 (N_15122,N_14658,N_14058);
nor U15123 (N_15123,N_14799,N_14031);
nand U15124 (N_15124,N_14221,N_14628);
xnor U15125 (N_15125,N_14632,N_14713);
nand U15126 (N_15126,N_13781,N_14052);
xnor U15127 (N_15127,N_14586,N_14708);
nand U15128 (N_15128,N_14433,N_14848);
nor U15129 (N_15129,N_13890,N_14291);
and U15130 (N_15130,N_14235,N_14861);
or U15131 (N_15131,N_14838,N_14537);
or U15132 (N_15132,N_14153,N_14106);
nand U15133 (N_15133,N_13964,N_14594);
nor U15134 (N_15134,N_13901,N_14250);
nand U15135 (N_15135,N_13777,N_14446);
and U15136 (N_15136,N_14288,N_14136);
and U15137 (N_15137,N_14038,N_14028);
nor U15138 (N_15138,N_13990,N_14203);
nand U15139 (N_15139,N_14274,N_14934);
nand U15140 (N_15140,N_13939,N_14869);
and U15141 (N_15141,N_13802,N_14144);
xor U15142 (N_15142,N_14360,N_14494);
xnor U15143 (N_15143,N_14477,N_14593);
and U15144 (N_15144,N_14841,N_14173);
nand U15145 (N_15145,N_14459,N_14742);
nor U15146 (N_15146,N_13915,N_14116);
xor U15147 (N_15147,N_14590,N_14637);
nand U15148 (N_15148,N_13897,N_14636);
and U15149 (N_15149,N_13856,N_14781);
or U15150 (N_15150,N_14259,N_14063);
and U15151 (N_15151,N_14933,N_14067);
nor U15152 (N_15152,N_14218,N_14830);
and U15153 (N_15153,N_14673,N_14088);
and U15154 (N_15154,N_14827,N_14169);
xor U15155 (N_15155,N_14545,N_14293);
xnor U15156 (N_15156,N_14828,N_14652);
or U15157 (N_15157,N_14925,N_14049);
nand U15158 (N_15158,N_14010,N_14831);
and U15159 (N_15159,N_14887,N_14935);
or U15160 (N_15160,N_14098,N_14776);
nand U15161 (N_15161,N_14908,N_14025);
and U15162 (N_15162,N_14046,N_14091);
xnor U15163 (N_15163,N_13989,N_14722);
or U15164 (N_15164,N_14316,N_14750);
nand U15165 (N_15165,N_14821,N_14795);
xnor U15166 (N_15166,N_14454,N_14581);
or U15167 (N_15167,N_14792,N_14176);
nor U15168 (N_15168,N_14749,N_14420);
or U15169 (N_15169,N_13974,N_14145);
xor U15170 (N_15170,N_14580,N_14435);
nand U15171 (N_15171,N_14810,N_14417);
nor U15172 (N_15172,N_13804,N_13973);
nor U15173 (N_15173,N_13826,N_14503);
xnor U15174 (N_15174,N_14967,N_14528);
or U15175 (N_15175,N_13797,N_14149);
nand U15176 (N_15176,N_14051,N_13799);
nand U15177 (N_15177,N_14788,N_14504);
xnor U15178 (N_15178,N_14982,N_14269);
xor U15179 (N_15179,N_14281,N_14225);
and U15180 (N_15180,N_13948,N_14415);
nor U15181 (N_15181,N_14732,N_14180);
xnor U15182 (N_15182,N_14512,N_13870);
nor U15183 (N_15183,N_14947,N_14604);
and U15184 (N_15184,N_14555,N_13900);
nand U15185 (N_15185,N_14495,N_14073);
and U15186 (N_15186,N_13861,N_14806);
or U15187 (N_15187,N_14201,N_14521);
xnor U15188 (N_15188,N_14836,N_13822);
xor U15189 (N_15189,N_14975,N_14087);
xor U15190 (N_15190,N_14276,N_14655);
nor U15191 (N_15191,N_14904,N_14335);
nand U15192 (N_15192,N_14738,N_14892);
xor U15193 (N_15193,N_14944,N_14968);
nor U15194 (N_15194,N_13762,N_14847);
xnor U15195 (N_15195,N_13920,N_14544);
xor U15196 (N_15196,N_14735,N_14854);
nand U15197 (N_15197,N_14684,N_13761);
nand U15198 (N_15198,N_14998,N_14143);
and U15199 (N_15199,N_14930,N_14591);
nor U15200 (N_15200,N_14157,N_14626);
xnor U15201 (N_15201,N_14719,N_13795);
and U15202 (N_15202,N_14730,N_14835);
or U15203 (N_15203,N_13863,N_14917);
nor U15204 (N_15204,N_14397,N_14541);
xnor U15205 (N_15205,N_14648,N_14677);
and U15206 (N_15206,N_13894,N_14532);
and U15207 (N_15207,N_14790,N_14161);
xnor U15208 (N_15208,N_14508,N_14260);
or U15209 (N_15209,N_14771,N_13832);
nor U15210 (N_15210,N_14355,N_13926);
nor U15211 (N_15211,N_13965,N_13903);
and U15212 (N_15212,N_14320,N_13859);
and U15213 (N_15213,N_14650,N_14496);
and U15214 (N_15214,N_14871,N_14723);
or U15215 (N_15215,N_14897,N_13852);
or U15216 (N_15216,N_14929,N_14400);
nand U15217 (N_15217,N_14819,N_13925);
nor U15218 (N_15218,N_14207,N_13775);
xnor U15219 (N_15219,N_14181,N_14409);
xor U15220 (N_15220,N_14922,N_14152);
nand U15221 (N_15221,N_14019,N_13940);
xnor U15222 (N_15222,N_14672,N_14105);
nor U15223 (N_15223,N_13956,N_14332);
nor U15224 (N_15224,N_14721,N_14139);
or U15225 (N_15225,N_14731,N_14502);
xnor U15226 (N_15226,N_14364,N_14622);
xor U15227 (N_15227,N_14410,N_14202);
or U15228 (N_15228,N_13806,N_14829);
nor U15229 (N_15229,N_13848,N_14156);
and U15230 (N_15230,N_14960,N_14900);
nand U15231 (N_15231,N_14909,N_14621);
or U15232 (N_15232,N_13879,N_14642);
xor U15233 (N_15233,N_14867,N_14839);
nand U15234 (N_15234,N_14330,N_14951);
nor U15235 (N_15235,N_13931,N_13928);
nand U15236 (N_15236,N_13997,N_14573);
or U15237 (N_15237,N_14124,N_14490);
nor U15238 (N_15238,N_14710,N_14458);
or U15239 (N_15239,N_14030,N_14077);
and U15240 (N_15240,N_14814,N_14205);
xor U15241 (N_15241,N_14809,N_14263);
or U15242 (N_15242,N_14372,N_14950);
or U15243 (N_15243,N_13823,N_14759);
and U15244 (N_15244,N_13838,N_14475);
nor U15245 (N_15245,N_14519,N_14423);
nor U15246 (N_15246,N_14737,N_13846);
xor U15247 (N_15247,N_14793,N_14901);
xor U15248 (N_15248,N_14640,N_14099);
and U15249 (N_15249,N_14718,N_14405);
nor U15250 (N_15250,N_14081,N_14921);
and U15251 (N_15251,N_14277,N_14135);
or U15252 (N_15252,N_14647,N_14527);
nor U15253 (N_15253,N_13936,N_13779);
and U15254 (N_15254,N_14125,N_13782);
nand U15255 (N_15255,N_14347,N_14388);
nor U15256 (N_15256,N_14399,N_14510);
nor U15257 (N_15257,N_14162,N_14992);
or U15258 (N_15258,N_13998,N_14365);
nor U15259 (N_15259,N_14965,N_14480);
or U15260 (N_15260,N_14891,N_14244);
nor U15261 (N_15261,N_14973,N_14910);
or U15262 (N_15262,N_13763,N_14309);
or U15263 (N_15263,N_14325,N_14689);
nand U15264 (N_15264,N_13881,N_14815);
and U15265 (N_15265,N_13840,N_13865);
nor U15266 (N_15266,N_14231,N_14055);
nor U15267 (N_15267,N_14070,N_14978);
and U15268 (N_15268,N_14807,N_14222);
nor U15269 (N_15269,N_14682,N_14761);
or U15270 (N_15270,N_14403,N_14322);
xnor U15271 (N_15271,N_13899,N_14424);
nand U15272 (N_15272,N_14849,N_14056);
nand U15273 (N_15273,N_13794,N_14999);
xnor U15274 (N_15274,N_14988,N_14624);
xor U15275 (N_15275,N_14247,N_14333);
xor U15276 (N_15276,N_14941,N_14669);
nand U15277 (N_15277,N_14366,N_14349);
nand U15278 (N_15278,N_14959,N_14818);
nand U15279 (N_15279,N_13875,N_14870);
or U15280 (N_15280,N_14264,N_14004);
nor U15281 (N_15281,N_13824,N_14346);
xnor U15282 (N_15282,N_14352,N_14101);
nand U15283 (N_15283,N_14482,N_13877);
nor U15284 (N_15284,N_13774,N_13986);
nor U15285 (N_15285,N_14568,N_14197);
nor U15286 (N_15286,N_14878,N_14635);
xor U15287 (N_15287,N_13908,N_14765);
xnor U15288 (N_15288,N_13977,N_13788);
nor U15289 (N_15289,N_14913,N_14567);
nand U15290 (N_15290,N_14690,N_14166);
or U15291 (N_15291,N_14448,N_14111);
xor U15292 (N_15292,N_14455,N_14741);
or U15293 (N_15293,N_14214,N_14246);
and U15294 (N_15294,N_14268,N_14398);
nand U15295 (N_15295,N_14142,N_14323);
or U15296 (N_15296,N_14104,N_14704);
nand U15297 (N_15297,N_14299,N_13759);
and U15298 (N_15298,N_13796,N_14003);
nand U15299 (N_15299,N_14434,N_14024);
or U15300 (N_15300,N_13791,N_14054);
xnor U15301 (N_15301,N_14767,N_13857);
nor U15302 (N_15302,N_13946,N_14356);
xor U15303 (N_15303,N_14351,N_14359);
xor U15304 (N_15304,N_13752,N_14608);
nand U15305 (N_15305,N_14075,N_14072);
nand U15306 (N_15306,N_14138,N_14262);
and U15307 (N_15307,N_14651,N_14813);
or U15308 (N_15308,N_13810,N_14855);
and U15309 (N_15309,N_14997,N_14109);
nand U15310 (N_15310,N_14062,N_14431);
xor U15311 (N_15311,N_13845,N_13790);
xnor U15312 (N_15312,N_13807,N_13984);
or U15313 (N_15313,N_14966,N_14286);
nand U15314 (N_15314,N_14367,N_14170);
nand U15315 (N_15315,N_14600,N_14165);
xnor U15316 (N_15316,N_14429,N_14680);
xor U15317 (N_15317,N_14114,N_14937);
nand U15318 (N_15318,N_14008,N_14625);
and U15319 (N_15319,N_13910,N_13853);
nor U15320 (N_15320,N_14112,N_14327);
nand U15321 (N_15321,N_14043,N_14665);
nand U15322 (N_15322,N_13839,N_14564);
nor U15323 (N_15323,N_14257,N_14154);
and U15324 (N_15324,N_14059,N_14612);
or U15325 (N_15325,N_13909,N_13854);
or U15326 (N_15326,N_14740,N_13862);
or U15327 (N_15327,N_14065,N_14863);
or U15328 (N_15328,N_14956,N_13967);
nor U15329 (N_15329,N_14602,N_14082);
xnor U15330 (N_15330,N_13819,N_13934);
or U15331 (N_15331,N_13829,N_13992);
nand U15332 (N_15332,N_14536,N_14126);
nor U15333 (N_15333,N_14725,N_14498);
xnor U15334 (N_15334,N_14437,N_14339);
xnor U15335 (N_15335,N_14954,N_13772);
nor U15336 (N_15336,N_14468,N_14701);
nor U15337 (N_15337,N_13987,N_14151);
nand U15338 (N_15338,N_13972,N_14786);
xor U15339 (N_15339,N_14957,N_14796);
xor U15340 (N_15340,N_14639,N_13803);
xnor U15341 (N_15341,N_14076,N_13850);
nor U15342 (N_15342,N_14927,N_14478);
nor U15343 (N_15343,N_14306,N_14938);
and U15344 (N_15344,N_14223,N_14245);
or U15345 (N_15345,N_14520,N_14185);
or U15346 (N_15346,N_14271,N_14471);
nor U15347 (N_15347,N_14228,N_13830);
nand U15348 (N_15348,N_14270,N_14832);
or U15349 (N_15349,N_14668,N_14345);
and U15350 (N_15350,N_14615,N_14122);
and U15351 (N_15351,N_13750,N_14511);
and U15352 (N_15352,N_14432,N_14241);
and U15353 (N_15353,N_14007,N_14993);
and U15354 (N_15354,N_14285,N_14422);
and U15355 (N_15355,N_14461,N_14906);
or U15356 (N_15356,N_14745,N_13980);
xor U15357 (N_15357,N_14069,N_13949);
xor U15358 (N_15358,N_14565,N_14307);
nor U15359 (N_15359,N_14920,N_14376);
or U15360 (N_15360,N_14885,N_14777);
xor U15361 (N_15361,N_13784,N_14611);
and U15362 (N_15362,N_14159,N_14419);
and U15363 (N_15363,N_14295,N_14616);
or U15364 (N_15364,N_14509,N_14762);
and U15365 (N_15365,N_14204,N_14686);
and U15366 (N_15366,N_13906,N_14557);
and U15367 (N_15367,N_14391,N_14607);
and U15368 (N_15368,N_14606,N_14823);
xor U15369 (N_15369,N_14447,N_13864);
nand U15370 (N_15370,N_14787,N_14487);
and U15371 (N_15371,N_14370,N_14808);
or U15372 (N_15372,N_14047,N_13770);
or U15373 (N_15373,N_14766,N_13768);
or U15374 (N_15374,N_14942,N_14485);
nor U15375 (N_15375,N_13760,N_14694);
nor U15376 (N_15376,N_14953,N_14439);
nor U15377 (N_15377,N_14387,N_14840);
xor U15378 (N_15378,N_14729,N_14340);
xnor U15379 (N_15379,N_14746,N_14884);
nor U15380 (N_15380,N_13814,N_13950);
nor U15381 (N_15381,N_14720,N_14852);
xor U15382 (N_15382,N_14210,N_13798);
xnor U15383 (N_15383,N_14483,N_14866);
nor U15384 (N_15384,N_14902,N_14785);
or U15385 (N_15385,N_14744,N_14195);
xnor U15386 (N_15386,N_14383,N_14018);
or U15387 (N_15387,N_14627,N_14385);
and U15388 (N_15388,N_14182,N_14456);
xnor U15389 (N_15389,N_14712,N_14479);
nand U15390 (N_15390,N_14378,N_14464);
or U15391 (N_15391,N_14553,N_14688);
or U15392 (N_15392,N_14193,N_14525);
nand U15393 (N_15393,N_13904,N_13874);
xor U15394 (N_15394,N_14898,N_14473);
or U15395 (N_15395,N_13755,N_14540);
xor U15396 (N_15396,N_14060,N_14631);
xnor U15397 (N_15397,N_14401,N_14646);
nor U15398 (N_15398,N_13860,N_14969);
nor U15399 (N_15399,N_14023,N_14407);
and U15400 (N_15400,N_14183,N_13855);
or U15401 (N_15401,N_14396,N_14706);
and U15402 (N_15402,N_13851,N_14577);
and U15403 (N_15403,N_14470,N_14272);
nand U15404 (N_15404,N_13836,N_14113);
nor U15405 (N_15405,N_14826,N_14402);
nand U15406 (N_15406,N_14817,N_14450);
nand U15407 (N_15407,N_14948,N_13793);
nor U15408 (N_15408,N_13783,N_13789);
nand U15409 (N_15409,N_14517,N_14530);
or U15410 (N_15410,N_14442,N_13968);
nor U15411 (N_15411,N_14576,N_14514);
or U15412 (N_15412,N_14444,N_14044);
nand U15413 (N_15413,N_14368,N_14547);
nand U15414 (N_15414,N_14265,N_14843);
or U15415 (N_15415,N_14497,N_14918);
or U15416 (N_15416,N_14150,N_14675);
and U15417 (N_15417,N_14513,N_14697);
or U15418 (N_15418,N_13773,N_14613);
and U15419 (N_15419,N_14312,N_13827);
and U15420 (N_15420,N_13960,N_14774);
nand U15421 (N_15421,N_14707,N_14623);
xor U15422 (N_15422,N_14751,N_14115);
nor U15423 (N_15423,N_14009,N_14501);
and U15424 (N_15424,N_13927,N_14859);
nor U15425 (N_15425,N_14949,N_14772);
nand U15426 (N_15426,N_14940,N_13912);
or U15427 (N_15427,N_14198,N_13991);
and U15428 (N_15428,N_13922,N_14341);
and U15429 (N_15429,N_14856,N_14562);
and U15430 (N_15430,N_14518,N_13918);
nand U15431 (N_15431,N_13929,N_14488);
xor U15432 (N_15432,N_13938,N_13871);
nor U15433 (N_15433,N_14693,N_14239);
or U15434 (N_15434,N_14261,N_14783);
nor U15435 (N_15435,N_14943,N_14911);
xnor U15436 (N_15436,N_14303,N_14522);
nand U15437 (N_15437,N_13887,N_13883);
nor U15438 (N_15438,N_14440,N_14097);
and U15439 (N_15439,N_14102,N_14337);
or U15440 (N_15440,N_14045,N_14061);
or U15441 (N_15441,N_14493,N_14457);
or U15442 (N_15442,N_14186,N_13886);
nand U15443 (N_15443,N_14538,N_14240);
and U15444 (N_15444,N_14130,N_13805);
nor U15445 (N_15445,N_14253,N_14164);
xor U15446 (N_15446,N_14236,N_14711);
nand U15447 (N_15447,N_14292,N_14199);
nand U15448 (N_15448,N_14224,N_13835);
xor U15449 (N_15449,N_13780,N_14110);
and U15450 (N_15450,N_14287,N_14486);
nand U15451 (N_15451,N_14392,N_14243);
nand U15452 (N_15452,N_14692,N_14916);
xor U15453 (N_15453,N_14283,N_14974);
nor U15454 (N_15454,N_14311,N_13868);
nand U15455 (N_15455,N_14797,N_14395);
and U15456 (N_15456,N_14148,N_14979);
nor U15457 (N_15457,N_14880,N_13970);
xor U15458 (N_15458,N_13834,N_13811);
or U15459 (N_15459,N_14258,N_13765);
nor U15460 (N_15460,N_14595,N_14317);
or U15461 (N_15461,N_14123,N_14233);
nor U15462 (N_15462,N_14484,N_14936);
or U15463 (N_15463,N_14298,N_14137);
or U15464 (N_15464,N_14784,N_14308);
nor U15465 (N_15465,N_14474,N_14079);
and U15466 (N_15466,N_14893,N_14516);
or U15467 (N_15467,N_14481,N_14361);
or U15468 (N_15468,N_14386,N_13756);
xnor U15469 (N_15469,N_14329,N_14127);
nor U15470 (N_15470,N_13866,N_14769);
nor U15471 (N_15471,N_13844,N_14390);
xnor U15472 (N_15472,N_14842,N_14342);
nor U15473 (N_15473,N_14131,N_14449);
and U15474 (N_15474,N_13935,N_14733);
xor U15475 (N_15475,N_14212,N_13766);
nor U15476 (N_15476,N_13818,N_14894);
and U15477 (N_15477,N_13884,N_13953);
xor U15478 (N_15478,N_14715,N_14438);
nor U15479 (N_15479,N_13813,N_14377);
nor U15480 (N_15480,N_14066,N_14605);
or U15481 (N_15481,N_14443,N_14549);
nand U15482 (N_15482,N_14027,N_13817);
or U15483 (N_15483,N_14011,N_14234);
xnor U15484 (N_15484,N_14500,N_14121);
xnor U15485 (N_15485,N_14986,N_14985);
or U15486 (N_15486,N_14297,N_13842);
or U15487 (N_15487,N_14641,N_14369);
nor U15488 (N_15488,N_13959,N_14108);
nor U15489 (N_15489,N_14574,N_14050);
or U15490 (N_15490,N_14515,N_14215);
and U15491 (N_15491,N_14256,N_13876);
and U15492 (N_15492,N_14505,N_14252);
or U15493 (N_15493,N_13880,N_14939);
or U15494 (N_15494,N_13792,N_14158);
nand U15495 (N_15495,N_14232,N_14194);
or U15496 (N_15496,N_14354,N_14931);
nor U15497 (N_15497,N_14667,N_14758);
nand U15498 (N_15498,N_14889,N_14996);
and U15499 (N_15499,N_14834,N_14571);
xnor U15500 (N_15500,N_14596,N_14923);
nand U15501 (N_15501,N_14092,N_14452);
xnor U15502 (N_15502,N_14928,N_14192);
xor U15503 (N_15503,N_14888,N_14629);
and U15504 (N_15504,N_14952,N_14375);
or U15505 (N_15505,N_14578,N_13878);
or U15506 (N_15506,N_14801,N_13821);
and U15507 (N_15507,N_14915,N_14217);
xnor U15508 (N_15508,N_13833,N_14381);
nand U15509 (N_15509,N_14551,N_14032);
and U15510 (N_15510,N_14371,N_14789);
and U15511 (N_15511,N_14800,N_14877);
nand U15512 (N_15512,N_14315,N_14211);
xnor U15513 (N_15513,N_13981,N_14981);
nand U15514 (N_15514,N_13812,N_14739);
nand U15515 (N_15515,N_14042,N_14919);
nand U15516 (N_15516,N_14837,N_14912);
and U15517 (N_15517,N_14558,N_14350);
or U15518 (N_15518,N_14583,N_13902);
xnor U15519 (N_15519,N_14653,N_13896);
and U15520 (N_15520,N_14133,N_14685);
and U15521 (N_15521,N_14086,N_14747);
or U15522 (N_15522,N_14882,N_14296);
nand U15523 (N_15523,N_13825,N_14976);
xnor U15524 (N_15524,N_14656,N_14413);
and U15525 (N_15525,N_14248,N_13976);
xor U15526 (N_15526,N_14768,N_14645);
and U15527 (N_15527,N_14764,N_13930);
or U15528 (N_15528,N_14358,N_14319);
nand U15529 (N_15529,N_14273,N_13776);
xnor U15530 (N_15530,N_14472,N_13917);
nand U15531 (N_15531,N_14294,N_14763);
nor U15532 (N_15532,N_14822,N_14175);
xor U15533 (N_15533,N_14816,N_14229);
nand U15534 (N_15534,N_14321,N_14546);
nand U15535 (N_15535,N_14570,N_14875);
nand U15536 (N_15536,N_14727,N_14563);
nand U15537 (N_15537,N_14290,N_14955);
and U15538 (N_15538,N_14373,N_14865);
or U15539 (N_15539,N_14022,N_14107);
nand U15540 (N_15540,N_14021,N_14582);
and U15541 (N_15541,N_14146,N_14178);
nand U15542 (N_15542,N_14649,N_14584);
nor U15543 (N_15543,N_14678,N_14991);
or U15544 (N_15544,N_14760,N_14699);
xor U15545 (N_15545,N_14189,N_14096);
or U15546 (N_15546,N_14414,N_13963);
nand U15547 (N_15547,N_14638,N_14266);
xor U15548 (N_15548,N_14548,N_14467);
or U15549 (N_15549,N_14132,N_14618);
nand U15550 (N_15550,N_14037,N_14053);
and U15551 (N_15551,N_14465,N_14824);
or U15552 (N_15552,N_14155,N_13888);
or U15553 (N_15553,N_14227,N_14945);
nand U15554 (N_15554,N_14064,N_14812);
or U15555 (N_15555,N_14811,N_14990);
or U15556 (N_15556,N_14794,N_14592);
xnor U15557 (N_15557,N_13947,N_14040);
nand U15558 (N_15558,N_13979,N_13971);
nor U15559 (N_15559,N_13954,N_14128);
nand U15560 (N_15560,N_14601,N_14754);
or U15561 (N_15561,N_13816,N_14630);
nor U15562 (N_15562,N_14140,N_14798);
xnor U15563 (N_15563,N_14989,N_14778);
or U15564 (N_15564,N_13758,N_14275);
and U15565 (N_15565,N_14167,N_14015);
nor U15566 (N_15566,N_13843,N_14393);
or U15567 (N_15567,N_14872,N_14634);
and U15568 (N_15568,N_14362,N_14663);
or U15569 (N_15569,N_14679,N_14962);
and U15570 (N_15570,N_13849,N_14550);
and U15571 (N_15571,N_14657,N_14716);
nand U15572 (N_15572,N_14676,N_13933);
or U15573 (N_15573,N_14289,N_14129);
nand U15574 (N_15574,N_14035,N_13757);
xnor U15575 (N_15575,N_14324,N_14074);
and U15576 (N_15576,N_14331,N_14507);
xnor U15577 (N_15577,N_14703,N_14569);
xnor U15578 (N_15578,N_14421,N_13882);
or U15579 (N_15579,N_14334,N_14280);
or U15580 (N_15580,N_14172,N_13809);
nor U15581 (N_15581,N_14914,N_13847);
xnor U15582 (N_15582,N_14026,N_13951);
or U15583 (N_15583,N_14425,N_13858);
and U15584 (N_15584,N_13786,N_14620);
or U15585 (N_15585,N_14963,N_14068);
or U15586 (N_15586,N_14492,N_14384);
nand U15587 (N_15587,N_14804,N_14850);
or U15588 (N_15588,N_13952,N_13867);
xor U15589 (N_15589,N_14441,N_14379);
nand U15590 (N_15590,N_13993,N_13769);
nand U15591 (N_15591,N_14860,N_13754);
nand U15592 (N_15592,N_13957,N_14526);
and U15593 (N_15593,N_14780,N_14094);
nand U15594 (N_15594,N_14005,N_13969);
and U15595 (N_15595,N_14671,N_13945);
nor U15596 (N_15596,N_14460,N_14531);
nor U15597 (N_15597,N_14029,N_14734);
nor U15598 (N_15598,N_14255,N_14282);
or U15599 (N_15599,N_14883,N_14987);
nand U15600 (N_15600,N_14220,N_14820);
nor U15601 (N_15601,N_14617,N_14881);
xnor U15602 (N_15602,N_14041,N_13837);
xor U15603 (N_15603,N_14599,N_14924);
and U15604 (N_15604,N_13932,N_14926);
and U15605 (N_15605,N_13944,N_13924);
xor U15606 (N_15606,N_14012,N_14588);
or U15607 (N_15607,N_14284,N_13955);
and U15608 (N_15608,N_14775,N_13907);
nand U15609 (N_15609,N_14539,N_13898);
or U15610 (N_15610,N_14310,N_14705);
and U15611 (N_15611,N_14048,N_14534);
and U15612 (N_15612,N_14779,N_14696);
nand U15613 (N_15613,N_14301,N_14242);
nor U15614 (N_15614,N_14691,N_13800);
or U15615 (N_15615,N_14416,N_14664);
xor U15616 (N_15616,N_13893,N_14219);
nand U15617 (N_15617,N_14080,N_14662);
xnor U15618 (N_15618,N_14770,N_14141);
or U15619 (N_15619,N_13767,N_14090);
nand U15620 (N_15620,N_14177,N_14995);
and U15621 (N_15621,N_14380,N_14489);
or U15622 (N_15622,N_14683,N_14755);
nor U15623 (N_15623,N_14994,N_14237);
and U15624 (N_15624,N_13988,N_14006);
xnor U15625 (N_15625,N_13869,N_14454);
and U15626 (N_15626,N_13861,N_14580);
or U15627 (N_15627,N_14334,N_14778);
nand U15628 (N_15628,N_14930,N_14561);
nand U15629 (N_15629,N_14817,N_14027);
or U15630 (N_15630,N_14773,N_14100);
and U15631 (N_15631,N_14979,N_14390);
and U15632 (N_15632,N_13812,N_13939);
or U15633 (N_15633,N_14658,N_14258);
xor U15634 (N_15634,N_14888,N_14042);
and U15635 (N_15635,N_14979,N_14096);
nor U15636 (N_15636,N_13787,N_14872);
nand U15637 (N_15637,N_14457,N_14626);
or U15638 (N_15638,N_14578,N_14185);
or U15639 (N_15639,N_14325,N_14342);
and U15640 (N_15640,N_14586,N_14343);
nor U15641 (N_15641,N_14683,N_13800);
nor U15642 (N_15642,N_13851,N_14710);
and U15643 (N_15643,N_14322,N_14058);
or U15644 (N_15644,N_14320,N_14431);
nor U15645 (N_15645,N_14621,N_13879);
and U15646 (N_15646,N_14584,N_14558);
nand U15647 (N_15647,N_14431,N_14889);
nor U15648 (N_15648,N_14129,N_14769);
or U15649 (N_15649,N_14609,N_14616);
nor U15650 (N_15650,N_14826,N_14614);
nor U15651 (N_15651,N_14115,N_14156);
and U15652 (N_15652,N_13764,N_14867);
nand U15653 (N_15653,N_13883,N_14965);
nor U15654 (N_15654,N_13850,N_14231);
xnor U15655 (N_15655,N_13765,N_14193);
xor U15656 (N_15656,N_14246,N_14584);
or U15657 (N_15657,N_14011,N_13804);
nor U15658 (N_15658,N_14653,N_14605);
nand U15659 (N_15659,N_14532,N_14397);
and U15660 (N_15660,N_14366,N_14902);
or U15661 (N_15661,N_14337,N_14409);
nor U15662 (N_15662,N_14165,N_13872);
nand U15663 (N_15663,N_14779,N_14380);
and U15664 (N_15664,N_14548,N_14926);
nor U15665 (N_15665,N_13773,N_14846);
xnor U15666 (N_15666,N_13797,N_14530);
xnor U15667 (N_15667,N_13843,N_14891);
and U15668 (N_15668,N_14287,N_13799);
and U15669 (N_15669,N_13771,N_14526);
xnor U15670 (N_15670,N_14610,N_14141);
and U15671 (N_15671,N_14625,N_13781);
nor U15672 (N_15672,N_14750,N_13886);
nor U15673 (N_15673,N_14008,N_14671);
and U15674 (N_15674,N_13763,N_14658);
or U15675 (N_15675,N_13994,N_14996);
or U15676 (N_15676,N_14052,N_13902);
nor U15677 (N_15677,N_14459,N_13893);
nor U15678 (N_15678,N_14944,N_14557);
nand U15679 (N_15679,N_14571,N_13775);
nand U15680 (N_15680,N_14821,N_14680);
or U15681 (N_15681,N_14528,N_14071);
or U15682 (N_15682,N_14975,N_13891);
nand U15683 (N_15683,N_14530,N_13864);
or U15684 (N_15684,N_14645,N_13887);
nor U15685 (N_15685,N_14466,N_14789);
or U15686 (N_15686,N_13755,N_14554);
nand U15687 (N_15687,N_14749,N_14322);
xor U15688 (N_15688,N_14042,N_14517);
nor U15689 (N_15689,N_14999,N_14675);
or U15690 (N_15690,N_13812,N_14610);
xnor U15691 (N_15691,N_13957,N_14152);
nand U15692 (N_15692,N_14415,N_14861);
nor U15693 (N_15693,N_14566,N_14995);
nor U15694 (N_15694,N_14336,N_14590);
or U15695 (N_15695,N_14314,N_14361);
xnor U15696 (N_15696,N_14045,N_14991);
nor U15697 (N_15697,N_13758,N_13777);
nor U15698 (N_15698,N_14477,N_14663);
nor U15699 (N_15699,N_14426,N_14963);
and U15700 (N_15700,N_13985,N_14240);
or U15701 (N_15701,N_14031,N_14995);
nor U15702 (N_15702,N_14559,N_14095);
and U15703 (N_15703,N_13825,N_13900);
and U15704 (N_15704,N_14141,N_14990);
nand U15705 (N_15705,N_13781,N_13928);
xor U15706 (N_15706,N_13807,N_14032);
nor U15707 (N_15707,N_13907,N_14562);
or U15708 (N_15708,N_14080,N_14550);
nor U15709 (N_15709,N_14245,N_14637);
or U15710 (N_15710,N_14534,N_14751);
nor U15711 (N_15711,N_14298,N_13859);
or U15712 (N_15712,N_14312,N_14211);
nor U15713 (N_15713,N_14889,N_14258);
or U15714 (N_15714,N_14682,N_14911);
nor U15715 (N_15715,N_14732,N_13783);
nor U15716 (N_15716,N_13827,N_14180);
xnor U15717 (N_15717,N_14383,N_14660);
nor U15718 (N_15718,N_14520,N_14045);
nor U15719 (N_15719,N_14430,N_14064);
nor U15720 (N_15720,N_14576,N_13787);
nor U15721 (N_15721,N_13775,N_14708);
and U15722 (N_15722,N_14726,N_14277);
and U15723 (N_15723,N_14998,N_14643);
and U15724 (N_15724,N_14090,N_14931);
xor U15725 (N_15725,N_13767,N_14855);
xor U15726 (N_15726,N_13759,N_14202);
nand U15727 (N_15727,N_13906,N_13801);
xnor U15728 (N_15728,N_14206,N_14498);
and U15729 (N_15729,N_14715,N_13755);
nor U15730 (N_15730,N_14384,N_14959);
xor U15731 (N_15731,N_14105,N_14987);
nand U15732 (N_15732,N_14443,N_13764);
xor U15733 (N_15733,N_14846,N_14082);
nand U15734 (N_15734,N_14262,N_14192);
nor U15735 (N_15735,N_14373,N_13750);
or U15736 (N_15736,N_14591,N_14972);
and U15737 (N_15737,N_13897,N_14282);
or U15738 (N_15738,N_14989,N_14604);
or U15739 (N_15739,N_13777,N_13971);
xnor U15740 (N_15740,N_14959,N_14889);
nor U15741 (N_15741,N_14900,N_14633);
or U15742 (N_15742,N_14056,N_13928);
or U15743 (N_15743,N_14736,N_14973);
or U15744 (N_15744,N_13876,N_14840);
or U15745 (N_15745,N_14226,N_13990);
nor U15746 (N_15746,N_13988,N_14744);
nor U15747 (N_15747,N_14212,N_13798);
xor U15748 (N_15748,N_14746,N_14883);
xnor U15749 (N_15749,N_13999,N_14277);
nor U15750 (N_15750,N_14711,N_14990);
and U15751 (N_15751,N_14840,N_14068);
or U15752 (N_15752,N_14398,N_14182);
nand U15753 (N_15753,N_14141,N_14979);
nand U15754 (N_15754,N_14666,N_14392);
nand U15755 (N_15755,N_14506,N_14804);
or U15756 (N_15756,N_14210,N_14887);
nand U15757 (N_15757,N_14149,N_14559);
or U15758 (N_15758,N_14228,N_14902);
and U15759 (N_15759,N_14525,N_14388);
and U15760 (N_15760,N_14970,N_14152);
nor U15761 (N_15761,N_14030,N_14304);
nand U15762 (N_15762,N_14199,N_13951);
or U15763 (N_15763,N_14851,N_14178);
or U15764 (N_15764,N_14525,N_14451);
nand U15765 (N_15765,N_13918,N_14998);
nor U15766 (N_15766,N_14256,N_14490);
nor U15767 (N_15767,N_14802,N_13929);
and U15768 (N_15768,N_14062,N_14315);
or U15769 (N_15769,N_13989,N_14384);
nor U15770 (N_15770,N_14682,N_14843);
nand U15771 (N_15771,N_14977,N_13759);
or U15772 (N_15772,N_14531,N_14690);
nand U15773 (N_15773,N_14222,N_13802);
nor U15774 (N_15774,N_14589,N_13807);
nand U15775 (N_15775,N_14111,N_13816);
xor U15776 (N_15776,N_14791,N_14636);
and U15777 (N_15777,N_14971,N_13981);
and U15778 (N_15778,N_13841,N_14925);
nor U15779 (N_15779,N_14854,N_14964);
and U15780 (N_15780,N_14015,N_14126);
or U15781 (N_15781,N_14546,N_14133);
nand U15782 (N_15782,N_14851,N_14296);
or U15783 (N_15783,N_13793,N_14751);
nand U15784 (N_15784,N_13964,N_14496);
nor U15785 (N_15785,N_14103,N_14897);
and U15786 (N_15786,N_14868,N_14482);
xnor U15787 (N_15787,N_14699,N_14744);
nor U15788 (N_15788,N_14637,N_14276);
nand U15789 (N_15789,N_14592,N_14786);
and U15790 (N_15790,N_13929,N_14481);
and U15791 (N_15791,N_14143,N_14893);
or U15792 (N_15792,N_14257,N_14057);
nand U15793 (N_15793,N_14790,N_14009);
and U15794 (N_15794,N_13985,N_14063);
xnor U15795 (N_15795,N_13809,N_14096);
xor U15796 (N_15796,N_13891,N_13928);
and U15797 (N_15797,N_14269,N_13841);
nand U15798 (N_15798,N_14735,N_14764);
nor U15799 (N_15799,N_14777,N_14255);
xnor U15800 (N_15800,N_14302,N_14912);
nand U15801 (N_15801,N_14972,N_14259);
xor U15802 (N_15802,N_14701,N_13750);
xor U15803 (N_15803,N_14878,N_14807);
nor U15804 (N_15804,N_13756,N_14633);
nand U15805 (N_15805,N_14807,N_14799);
nand U15806 (N_15806,N_14976,N_13900);
nand U15807 (N_15807,N_14235,N_14951);
nand U15808 (N_15808,N_14448,N_14505);
nand U15809 (N_15809,N_14576,N_14355);
nand U15810 (N_15810,N_14098,N_14489);
xnor U15811 (N_15811,N_14183,N_14986);
nand U15812 (N_15812,N_14411,N_14852);
and U15813 (N_15813,N_14759,N_13804);
nor U15814 (N_15814,N_13978,N_13798);
nor U15815 (N_15815,N_14325,N_14102);
or U15816 (N_15816,N_14317,N_14468);
or U15817 (N_15817,N_14257,N_14242);
nor U15818 (N_15818,N_14395,N_14038);
nor U15819 (N_15819,N_14269,N_14792);
nand U15820 (N_15820,N_14386,N_14099);
or U15821 (N_15821,N_14047,N_14098);
nor U15822 (N_15822,N_14787,N_13757);
nand U15823 (N_15823,N_14090,N_14684);
xnor U15824 (N_15824,N_14842,N_13996);
and U15825 (N_15825,N_13752,N_13826);
xnor U15826 (N_15826,N_14321,N_14938);
nor U15827 (N_15827,N_14560,N_13829);
nand U15828 (N_15828,N_14991,N_13926);
nor U15829 (N_15829,N_14488,N_13780);
nor U15830 (N_15830,N_14481,N_14729);
nor U15831 (N_15831,N_14012,N_14479);
nor U15832 (N_15832,N_14844,N_14178);
or U15833 (N_15833,N_14911,N_14051);
xnor U15834 (N_15834,N_14917,N_13818);
and U15835 (N_15835,N_14791,N_14858);
nand U15836 (N_15836,N_14283,N_13807);
and U15837 (N_15837,N_14749,N_14487);
xnor U15838 (N_15838,N_14795,N_14929);
or U15839 (N_15839,N_14769,N_14906);
and U15840 (N_15840,N_14064,N_14522);
or U15841 (N_15841,N_14307,N_14579);
and U15842 (N_15842,N_13975,N_14263);
nor U15843 (N_15843,N_14855,N_13846);
nand U15844 (N_15844,N_14956,N_14869);
or U15845 (N_15845,N_14641,N_14388);
nand U15846 (N_15846,N_14836,N_14579);
xor U15847 (N_15847,N_14338,N_14111);
and U15848 (N_15848,N_13938,N_14274);
nand U15849 (N_15849,N_14334,N_14811);
and U15850 (N_15850,N_14500,N_14938);
xor U15851 (N_15851,N_14013,N_13857);
or U15852 (N_15852,N_14492,N_14934);
nor U15853 (N_15853,N_14524,N_14125);
nor U15854 (N_15854,N_14329,N_13857);
or U15855 (N_15855,N_14043,N_14662);
xor U15856 (N_15856,N_14171,N_13753);
nor U15857 (N_15857,N_14924,N_14210);
or U15858 (N_15858,N_14456,N_14521);
or U15859 (N_15859,N_14462,N_14606);
nand U15860 (N_15860,N_14075,N_13966);
xnor U15861 (N_15861,N_14070,N_14872);
xor U15862 (N_15862,N_14164,N_14869);
or U15863 (N_15863,N_14706,N_14146);
or U15864 (N_15864,N_14464,N_14604);
or U15865 (N_15865,N_14935,N_14809);
xnor U15866 (N_15866,N_14814,N_14518);
or U15867 (N_15867,N_14136,N_13807);
nand U15868 (N_15868,N_14395,N_14471);
xor U15869 (N_15869,N_13993,N_14816);
xnor U15870 (N_15870,N_13801,N_14707);
nor U15871 (N_15871,N_14813,N_14818);
and U15872 (N_15872,N_14919,N_14231);
or U15873 (N_15873,N_14238,N_14185);
nor U15874 (N_15874,N_14317,N_13911);
and U15875 (N_15875,N_13966,N_14206);
xnor U15876 (N_15876,N_14116,N_14484);
or U15877 (N_15877,N_14099,N_13974);
nor U15878 (N_15878,N_14733,N_13882);
nor U15879 (N_15879,N_14834,N_14084);
nor U15880 (N_15880,N_14904,N_14090);
xnor U15881 (N_15881,N_14590,N_14188);
and U15882 (N_15882,N_14573,N_13890);
nand U15883 (N_15883,N_14042,N_14048);
xnor U15884 (N_15884,N_14052,N_13897);
nor U15885 (N_15885,N_14315,N_14231);
and U15886 (N_15886,N_14524,N_14219);
nand U15887 (N_15887,N_14457,N_14190);
nand U15888 (N_15888,N_14754,N_14267);
xor U15889 (N_15889,N_14319,N_14778);
nand U15890 (N_15890,N_14811,N_14630);
nand U15891 (N_15891,N_14931,N_14166);
and U15892 (N_15892,N_13755,N_13761);
or U15893 (N_15893,N_13940,N_14408);
or U15894 (N_15894,N_14699,N_14265);
nand U15895 (N_15895,N_14108,N_14501);
and U15896 (N_15896,N_14957,N_14665);
and U15897 (N_15897,N_14607,N_14307);
nand U15898 (N_15898,N_14050,N_13822);
or U15899 (N_15899,N_14433,N_14739);
nand U15900 (N_15900,N_14397,N_13818);
or U15901 (N_15901,N_14334,N_14273);
or U15902 (N_15902,N_13961,N_14438);
or U15903 (N_15903,N_13794,N_14746);
nor U15904 (N_15904,N_14929,N_14882);
nor U15905 (N_15905,N_13757,N_14769);
nand U15906 (N_15906,N_14277,N_14211);
xnor U15907 (N_15907,N_14177,N_13869);
and U15908 (N_15908,N_14196,N_14667);
or U15909 (N_15909,N_14777,N_13951);
or U15910 (N_15910,N_14941,N_14971);
nor U15911 (N_15911,N_14902,N_14018);
nor U15912 (N_15912,N_14040,N_13832);
nor U15913 (N_15913,N_14273,N_14148);
nor U15914 (N_15914,N_14721,N_14613);
nand U15915 (N_15915,N_14319,N_14535);
or U15916 (N_15916,N_14764,N_14363);
xnor U15917 (N_15917,N_14650,N_13916);
or U15918 (N_15918,N_13829,N_14969);
nand U15919 (N_15919,N_14038,N_14927);
xor U15920 (N_15920,N_14923,N_14970);
xnor U15921 (N_15921,N_14500,N_14840);
nor U15922 (N_15922,N_13905,N_14819);
xnor U15923 (N_15923,N_14299,N_14755);
xnor U15924 (N_15924,N_14117,N_14355);
nand U15925 (N_15925,N_14425,N_14182);
or U15926 (N_15926,N_14848,N_13932);
or U15927 (N_15927,N_14671,N_14611);
nand U15928 (N_15928,N_13900,N_14308);
nor U15929 (N_15929,N_14765,N_14601);
nand U15930 (N_15930,N_14393,N_14664);
and U15931 (N_15931,N_14340,N_13920);
or U15932 (N_15932,N_14028,N_13862);
nand U15933 (N_15933,N_14342,N_14698);
or U15934 (N_15934,N_14482,N_14130);
and U15935 (N_15935,N_14215,N_14526);
nand U15936 (N_15936,N_14345,N_14929);
or U15937 (N_15937,N_14538,N_13825);
xor U15938 (N_15938,N_14390,N_14341);
nand U15939 (N_15939,N_13908,N_14422);
nand U15940 (N_15940,N_14570,N_14957);
nor U15941 (N_15941,N_14353,N_14616);
xnor U15942 (N_15942,N_14544,N_14705);
xnor U15943 (N_15943,N_14860,N_14423);
and U15944 (N_15944,N_14837,N_14211);
nand U15945 (N_15945,N_14917,N_13938);
and U15946 (N_15946,N_14420,N_14255);
xnor U15947 (N_15947,N_14214,N_14514);
nand U15948 (N_15948,N_14602,N_14909);
nand U15949 (N_15949,N_13809,N_14305);
nor U15950 (N_15950,N_14318,N_14760);
nor U15951 (N_15951,N_14057,N_14865);
nor U15952 (N_15952,N_14324,N_14050);
and U15953 (N_15953,N_13900,N_13990);
or U15954 (N_15954,N_14121,N_14853);
nor U15955 (N_15955,N_14253,N_14258);
nor U15956 (N_15956,N_14618,N_14859);
and U15957 (N_15957,N_13817,N_14861);
nor U15958 (N_15958,N_14738,N_14454);
or U15959 (N_15959,N_13871,N_13852);
xor U15960 (N_15960,N_13768,N_14525);
or U15961 (N_15961,N_14685,N_14106);
and U15962 (N_15962,N_14250,N_14770);
or U15963 (N_15963,N_14811,N_14886);
or U15964 (N_15964,N_14744,N_14223);
xnor U15965 (N_15965,N_14998,N_14242);
or U15966 (N_15966,N_14162,N_14575);
nand U15967 (N_15967,N_14741,N_14701);
and U15968 (N_15968,N_14810,N_14062);
nand U15969 (N_15969,N_13754,N_14879);
xor U15970 (N_15970,N_14085,N_14199);
nor U15971 (N_15971,N_14366,N_14942);
and U15972 (N_15972,N_14042,N_14038);
and U15973 (N_15973,N_13761,N_14674);
nor U15974 (N_15974,N_13949,N_14101);
and U15975 (N_15975,N_14722,N_14419);
xor U15976 (N_15976,N_13982,N_14937);
xor U15977 (N_15977,N_14848,N_14268);
nor U15978 (N_15978,N_14415,N_13836);
xor U15979 (N_15979,N_14079,N_14764);
or U15980 (N_15980,N_14606,N_14394);
nor U15981 (N_15981,N_14992,N_14182);
nand U15982 (N_15982,N_13765,N_14273);
nor U15983 (N_15983,N_14179,N_14125);
nand U15984 (N_15984,N_13925,N_13782);
xnor U15985 (N_15985,N_13852,N_14315);
xor U15986 (N_15986,N_14375,N_14177);
nor U15987 (N_15987,N_14490,N_14662);
nor U15988 (N_15988,N_14946,N_14839);
nand U15989 (N_15989,N_14315,N_14358);
xnor U15990 (N_15990,N_14698,N_14504);
nand U15991 (N_15991,N_14542,N_13990);
and U15992 (N_15992,N_14082,N_13777);
xor U15993 (N_15993,N_14033,N_13996);
or U15994 (N_15994,N_14743,N_14099);
and U15995 (N_15995,N_14192,N_14918);
or U15996 (N_15996,N_14137,N_14795);
nor U15997 (N_15997,N_13765,N_14829);
and U15998 (N_15998,N_14258,N_14625);
and U15999 (N_15999,N_14171,N_13766);
nand U16000 (N_16000,N_14082,N_14308);
or U16001 (N_16001,N_14460,N_13750);
and U16002 (N_16002,N_14974,N_14722);
and U16003 (N_16003,N_14574,N_14898);
or U16004 (N_16004,N_13840,N_14797);
nand U16005 (N_16005,N_14677,N_14831);
xor U16006 (N_16006,N_14412,N_13996);
xor U16007 (N_16007,N_13929,N_14532);
and U16008 (N_16008,N_14345,N_14977);
xor U16009 (N_16009,N_14944,N_14022);
xor U16010 (N_16010,N_14299,N_14729);
nand U16011 (N_16011,N_14396,N_14388);
nand U16012 (N_16012,N_14863,N_14594);
nand U16013 (N_16013,N_13902,N_14072);
xnor U16014 (N_16014,N_13785,N_14747);
xnor U16015 (N_16015,N_14684,N_13873);
nor U16016 (N_16016,N_13778,N_14048);
nor U16017 (N_16017,N_14823,N_14123);
xnor U16018 (N_16018,N_14927,N_14118);
nor U16019 (N_16019,N_14145,N_14423);
xnor U16020 (N_16020,N_14608,N_14716);
nand U16021 (N_16021,N_13801,N_13982);
and U16022 (N_16022,N_13866,N_13953);
nor U16023 (N_16023,N_13976,N_14578);
nor U16024 (N_16024,N_14877,N_14042);
or U16025 (N_16025,N_14078,N_14534);
and U16026 (N_16026,N_14086,N_14775);
nand U16027 (N_16027,N_14145,N_14178);
nor U16028 (N_16028,N_14461,N_14942);
nor U16029 (N_16029,N_14417,N_14833);
nand U16030 (N_16030,N_13897,N_14736);
nor U16031 (N_16031,N_13786,N_14827);
and U16032 (N_16032,N_14618,N_14085);
nor U16033 (N_16033,N_14244,N_14988);
or U16034 (N_16034,N_13904,N_14723);
and U16035 (N_16035,N_14220,N_14203);
nand U16036 (N_16036,N_13829,N_14042);
nor U16037 (N_16037,N_14202,N_14888);
or U16038 (N_16038,N_13995,N_14924);
nand U16039 (N_16039,N_14814,N_13951);
nand U16040 (N_16040,N_13773,N_14389);
nand U16041 (N_16041,N_14953,N_14671);
or U16042 (N_16042,N_13952,N_14675);
or U16043 (N_16043,N_14136,N_14998);
and U16044 (N_16044,N_14157,N_14828);
xor U16045 (N_16045,N_14305,N_14568);
or U16046 (N_16046,N_14197,N_14548);
or U16047 (N_16047,N_14521,N_14588);
nor U16048 (N_16048,N_14153,N_14276);
xor U16049 (N_16049,N_14884,N_14886);
nand U16050 (N_16050,N_14167,N_14622);
xor U16051 (N_16051,N_14591,N_14968);
and U16052 (N_16052,N_14432,N_13886);
and U16053 (N_16053,N_14773,N_14613);
xnor U16054 (N_16054,N_14729,N_13808);
nor U16055 (N_16055,N_14109,N_14823);
or U16056 (N_16056,N_14890,N_14813);
or U16057 (N_16057,N_14034,N_14252);
xnor U16058 (N_16058,N_14453,N_14197);
xnor U16059 (N_16059,N_14569,N_14328);
nand U16060 (N_16060,N_14881,N_14971);
nor U16061 (N_16061,N_14754,N_14814);
or U16062 (N_16062,N_14176,N_14904);
nor U16063 (N_16063,N_14746,N_14657);
and U16064 (N_16064,N_13926,N_13936);
xor U16065 (N_16065,N_14619,N_14322);
nand U16066 (N_16066,N_14436,N_14735);
nand U16067 (N_16067,N_13881,N_14185);
and U16068 (N_16068,N_14793,N_14351);
nand U16069 (N_16069,N_13978,N_13838);
or U16070 (N_16070,N_13924,N_14571);
or U16071 (N_16071,N_13848,N_14937);
and U16072 (N_16072,N_14963,N_14248);
and U16073 (N_16073,N_14646,N_14372);
nand U16074 (N_16074,N_14994,N_14041);
or U16075 (N_16075,N_14458,N_14083);
and U16076 (N_16076,N_14151,N_14275);
nor U16077 (N_16077,N_14717,N_14925);
xor U16078 (N_16078,N_14243,N_13881);
xnor U16079 (N_16079,N_14933,N_14597);
or U16080 (N_16080,N_14423,N_14637);
nor U16081 (N_16081,N_14413,N_14870);
nand U16082 (N_16082,N_14151,N_14527);
xor U16083 (N_16083,N_13883,N_14759);
nand U16084 (N_16084,N_14885,N_14414);
xnor U16085 (N_16085,N_14886,N_14129);
xnor U16086 (N_16086,N_14620,N_14873);
and U16087 (N_16087,N_14087,N_13926);
nor U16088 (N_16088,N_14690,N_14049);
nand U16089 (N_16089,N_14790,N_13973);
or U16090 (N_16090,N_14329,N_14875);
nand U16091 (N_16091,N_14177,N_14157);
and U16092 (N_16092,N_14123,N_13862);
nand U16093 (N_16093,N_14288,N_14204);
nand U16094 (N_16094,N_14280,N_13804);
nor U16095 (N_16095,N_14424,N_14890);
nor U16096 (N_16096,N_14889,N_14306);
and U16097 (N_16097,N_14904,N_13894);
and U16098 (N_16098,N_13960,N_14633);
nand U16099 (N_16099,N_14480,N_14850);
or U16100 (N_16100,N_13889,N_14909);
nand U16101 (N_16101,N_14994,N_14936);
xnor U16102 (N_16102,N_13982,N_14006);
and U16103 (N_16103,N_13915,N_14730);
xnor U16104 (N_16104,N_14007,N_14082);
nor U16105 (N_16105,N_14235,N_14077);
and U16106 (N_16106,N_14858,N_14704);
nand U16107 (N_16107,N_14589,N_14972);
nand U16108 (N_16108,N_14274,N_14599);
and U16109 (N_16109,N_14756,N_13865);
or U16110 (N_16110,N_14963,N_14448);
or U16111 (N_16111,N_14563,N_14016);
nand U16112 (N_16112,N_14585,N_14664);
xnor U16113 (N_16113,N_14592,N_14857);
and U16114 (N_16114,N_14692,N_13958);
and U16115 (N_16115,N_14627,N_13843);
or U16116 (N_16116,N_14061,N_14848);
or U16117 (N_16117,N_14347,N_14339);
xor U16118 (N_16118,N_14210,N_14068);
and U16119 (N_16119,N_14027,N_14212);
and U16120 (N_16120,N_14029,N_14861);
or U16121 (N_16121,N_14473,N_14394);
or U16122 (N_16122,N_14489,N_14432);
nand U16123 (N_16123,N_13891,N_14102);
and U16124 (N_16124,N_14708,N_14882);
and U16125 (N_16125,N_14899,N_14866);
nor U16126 (N_16126,N_13849,N_14925);
xnor U16127 (N_16127,N_14505,N_14526);
nor U16128 (N_16128,N_14945,N_14859);
xnor U16129 (N_16129,N_14309,N_13832);
nor U16130 (N_16130,N_13968,N_14865);
nand U16131 (N_16131,N_14707,N_13866);
or U16132 (N_16132,N_14923,N_14119);
nor U16133 (N_16133,N_14701,N_14191);
nand U16134 (N_16134,N_14333,N_14582);
nor U16135 (N_16135,N_13976,N_13908);
and U16136 (N_16136,N_14154,N_13984);
or U16137 (N_16137,N_14597,N_14999);
xnor U16138 (N_16138,N_14614,N_14529);
nor U16139 (N_16139,N_14615,N_14910);
nand U16140 (N_16140,N_14512,N_14310);
xor U16141 (N_16141,N_14811,N_14288);
and U16142 (N_16142,N_13908,N_14904);
or U16143 (N_16143,N_14569,N_13881);
nor U16144 (N_16144,N_14903,N_14506);
or U16145 (N_16145,N_14214,N_14817);
nor U16146 (N_16146,N_14976,N_13766);
nand U16147 (N_16147,N_13847,N_14255);
or U16148 (N_16148,N_14678,N_14182);
nor U16149 (N_16149,N_14798,N_14064);
xnor U16150 (N_16150,N_14145,N_14904);
and U16151 (N_16151,N_13923,N_13873);
xnor U16152 (N_16152,N_14353,N_13788);
nand U16153 (N_16153,N_14156,N_14047);
nor U16154 (N_16154,N_14662,N_14169);
or U16155 (N_16155,N_14410,N_14851);
xnor U16156 (N_16156,N_14941,N_14689);
or U16157 (N_16157,N_13858,N_14202);
xnor U16158 (N_16158,N_14817,N_14818);
and U16159 (N_16159,N_14904,N_13864);
and U16160 (N_16160,N_14085,N_14477);
xnor U16161 (N_16161,N_14820,N_14395);
nand U16162 (N_16162,N_14291,N_14043);
or U16163 (N_16163,N_14869,N_14207);
xor U16164 (N_16164,N_14976,N_14155);
xnor U16165 (N_16165,N_14300,N_14277);
nor U16166 (N_16166,N_13785,N_14767);
and U16167 (N_16167,N_14565,N_14516);
and U16168 (N_16168,N_14971,N_13838);
or U16169 (N_16169,N_14573,N_14643);
nor U16170 (N_16170,N_13816,N_14466);
nor U16171 (N_16171,N_14568,N_13958);
nand U16172 (N_16172,N_14324,N_14449);
xnor U16173 (N_16173,N_14726,N_14266);
and U16174 (N_16174,N_14620,N_13789);
and U16175 (N_16175,N_14785,N_14923);
and U16176 (N_16176,N_13930,N_14553);
or U16177 (N_16177,N_13799,N_13982);
or U16178 (N_16178,N_13865,N_14125);
or U16179 (N_16179,N_13805,N_13991);
and U16180 (N_16180,N_14862,N_14010);
nor U16181 (N_16181,N_14615,N_14302);
or U16182 (N_16182,N_14377,N_13979);
xnor U16183 (N_16183,N_14097,N_13915);
nor U16184 (N_16184,N_14323,N_14842);
or U16185 (N_16185,N_14767,N_13946);
nand U16186 (N_16186,N_13848,N_14800);
xnor U16187 (N_16187,N_14008,N_14382);
nand U16188 (N_16188,N_13883,N_14539);
nand U16189 (N_16189,N_14705,N_14242);
xor U16190 (N_16190,N_14815,N_13922);
and U16191 (N_16191,N_14547,N_14668);
nand U16192 (N_16192,N_14442,N_13907);
xnor U16193 (N_16193,N_14333,N_14593);
or U16194 (N_16194,N_13963,N_13950);
nand U16195 (N_16195,N_14618,N_13906);
xnor U16196 (N_16196,N_14424,N_13785);
nor U16197 (N_16197,N_13820,N_14349);
and U16198 (N_16198,N_13925,N_14400);
nor U16199 (N_16199,N_14909,N_14347);
or U16200 (N_16200,N_14610,N_14274);
and U16201 (N_16201,N_14145,N_14945);
and U16202 (N_16202,N_14586,N_14511);
nand U16203 (N_16203,N_13806,N_14646);
or U16204 (N_16204,N_14007,N_14562);
or U16205 (N_16205,N_13834,N_14152);
xor U16206 (N_16206,N_14316,N_14304);
nand U16207 (N_16207,N_13939,N_14342);
nand U16208 (N_16208,N_14916,N_14300);
or U16209 (N_16209,N_14534,N_14720);
xor U16210 (N_16210,N_14173,N_14014);
or U16211 (N_16211,N_13820,N_14874);
xnor U16212 (N_16212,N_14663,N_14769);
nor U16213 (N_16213,N_13902,N_14529);
nand U16214 (N_16214,N_14616,N_14416);
or U16215 (N_16215,N_14480,N_14820);
and U16216 (N_16216,N_14832,N_14129);
or U16217 (N_16217,N_14389,N_14797);
xnor U16218 (N_16218,N_14548,N_14303);
or U16219 (N_16219,N_14944,N_14513);
and U16220 (N_16220,N_14733,N_14951);
nand U16221 (N_16221,N_14316,N_14683);
xor U16222 (N_16222,N_14955,N_14123);
nand U16223 (N_16223,N_13985,N_14722);
nor U16224 (N_16224,N_14765,N_13984);
nand U16225 (N_16225,N_14675,N_14172);
or U16226 (N_16226,N_14066,N_14571);
nor U16227 (N_16227,N_14063,N_14105);
xnor U16228 (N_16228,N_14233,N_14167);
and U16229 (N_16229,N_14298,N_14601);
or U16230 (N_16230,N_14786,N_13987);
nand U16231 (N_16231,N_14141,N_14101);
and U16232 (N_16232,N_13841,N_14220);
nor U16233 (N_16233,N_14577,N_14299);
xor U16234 (N_16234,N_14615,N_13752);
or U16235 (N_16235,N_14188,N_14824);
nor U16236 (N_16236,N_13800,N_14641);
nor U16237 (N_16237,N_14345,N_14119);
xnor U16238 (N_16238,N_13775,N_14424);
xnor U16239 (N_16239,N_13776,N_14174);
and U16240 (N_16240,N_14106,N_14743);
nand U16241 (N_16241,N_14516,N_14760);
or U16242 (N_16242,N_14077,N_13758);
xnor U16243 (N_16243,N_14188,N_14432);
nand U16244 (N_16244,N_14712,N_14175);
nand U16245 (N_16245,N_13936,N_14336);
nand U16246 (N_16246,N_14846,N_14792);
xor U16247 (N_16247,N_14076,N_14061);
and U16248 (N_16248,N_14662,N_13968);
nor U16249 (N_16249,N_14685,N_13989);
and U16250 (N_16250,N_15928,N_15005);
nor U16251 (N_16251,N_15430,N_15596);
or U16252 (N_16252,N_16011,N_15177);
nand U16253 (N_16253,N_15066,N_15132);
xnor U16254 (N_16254,N_16130,N_15585);
or U16255 (N_16255,N_15803,N_15749);
or U16256 (N_16256,N_15047,N_15074);
nand U16257 (N_16257,N_16024,N_15082);
nor U16258 (N_16258,N_16199,N_15506);
or U16259 (N_16259,N_16154,N_16073);
or U16260 (N_16260,N_15703,N_15198);
nor U16261 (N_16261,N_15744,N_15060);
or U16262 (N_16262,N_15178,N_15913);
nor U16263 (N_16263,N_15428,N_15118);
xor U16264 (N_16264,N_15455,N_15248);
xor U16265 (N_16265,N_15834,N_15383);
and U16266 (N_16266,N_16075,N_15784);
or U16267 (N_16267,N_15173,N_15948);
and U16268 (N_16268,N_15999,N_15136);
nor U16269 (N_16269,N_15688,N_15564);
or U16270 (N_16270,N_15826,N_15634);
nor U16271 (N_16271,N_16122,N_15462);
or U16272 (N_16272,N_15276,N_15465);
or U16273 (N_16273,N_15116,N_15985);
nand U16274 (N_16274,N_15336,N_16184);
and U16275 (N_16275,N_15451,N_15864);
xnor U16276 (N_16276,N_15840,N_15930);
xnor U16277 (N_16277,N_15499,N_15095);
nand U16278 (N_16278,N_15482,N_15642);
or U16279 (N_16279,N_15282,N_15500);
nor U16280 (N_16280,N_16091,N_15837);
and U16281 (N_16281,N_15824,N_16242);
nand U16282 (N_16282,N_15423,N_16236);
or U16283 (N_16283,N_16038,N_16004);
nor U16284 (N_16284,N_15606,N_16089);
and U16285 (N_16285,N_15682,N_15615);
xor U16286 (N_16286,N_15502,N_15216);
and U16287 (N_16287,N_15994,N_15043);
nand U16288 (N_16288,N_16027,N_15353);
xnor U16289 (N_16289,N_15631,N_15644);
xor U16290 (N_16290,N_16243,N_15001);
nand U16291 (N_16291,N_15846,N_15998);
or U16292 (N_16292,N_15341,N_15097);
and U16293 (N_16293,N_15681,N_16115);
nor U16294 (N_16294,N_16202,N_15275);
and U16295 (N_16295,N_15504,N_15203);
nor U16296 (N_16296,N_16097,N_15664);
and U16297 (N_16297,N_15626,N_15153);
xnor U16298 (N_16298,N_15567,N_15947);
nor U16299 (N_16299,N_16132,N_16066);
and U16300 (N_16300,N_15384,N_15781);
or U16301 (N_16301,N_15167,N_15478);
xnor U16302 (N_16302,N_15022,N_15603);
or U16303 (N_16303,N_16082,N_16120);
and U16304 (N_16304,N_15378,N_15432);
or U16305 (N_16305,N_16214,N_15185);
nand U16306 (N_16306,N_15550,N_15356);
xnor U16307 (N_16307,N_15100,N_15842);
and U16308 (N_16308,N_15918,N_15814);
nand U16309 (N_16309,N_15474,N_15157);
nor U16310 (N_16310,N_15054,N_16197);
xor U16311 (N_16311,N_15010,N_15140);
or U16312 (N_16312,N_15458,N_15106);
nor U16313 (N_16313,N_15878,N_15014);
nor U16314 (N_16314,N_16131,N_15058);
nand U16315 (N_16315,N_15900,N_15121);
nand U16316 (N_16316,N_15646,N_15373);
nand U16317 (N_16317,N_15069,N_15623);
nand U16318 (N_16318,N_15907,N_15475);
nand U16319 (N_16319,N_15126,N_15723);
and U16320 (N_16320,N_15484,N_15397);
nor U16321 (N_16321,N_16167,N_16051);
nor U16322 (N_16322,N_15130,N_15419);
nand U16323 (N_16323,N_15041,N_15827);
or U16324 (N_16324,N_15344,N_15571);
nor U16325 (N_16325,N_15717,N_16030);
or U16326 (N_16326,N_15169,N_15141);
and U16327 (N_16327,N_15368,N_15332);
xor U16328 (N_16328,N_15679,N_16116);
nor U16329 (N_16329,N_15329,N_16060);
nor U16330 (N_16330,N_15525,N_15122);
nand U16331 (N_16331,N_15135,N_15694);
or U16332 (N_16332,N_15162,N_15779);
and U16333 (N_16333,N_15796,N_15745);
nand U16334 (N_16334,N_15736,N_15156);
nand U16335 (N_16335,N_15922,N_16233);
nand U16336 (N_16336,N_15547,N_16149);
nor U16337 (N_16337,N_15188,N_15676);
xnor U16338 (N_16338,N_15070,N_15269);
nand U16339 (N_16339,N_15242,N_15758);
nand U16340 (N_16340,N_15017,N_15446);
xnor U16341 (N_16341,N_15243,N_15398);
nor U16342 (N_16342,N_15290,N_15608);
nor U16343 (N_16343,N_15230,N_15975);
nor U16344 (N_16344,N_15856,N_15422);
and U16345 (N_16345,N_15649,N_15782);
nand U16346 (N_16346,N_15027,N_15955);
nand U16347 (N_16347,N_15754,N_15711);
xor U16348 (N_16348,N_15841,N_15285);
nor U16349 (N_16349,N_15390,N_15809);
or U16350 (N_16350,N_15175,N_15035);
nor U16351 (N_16351,N_15743,N_15239);
or U16352 (N_16352,N_15435,N_15150);
nor U16353 (N_16353,N_15487,N_15407);
and U16354 (N_16354,N_15024,N_15787);
nor U16355 (N_16355,N_15697,N_15920);
nor U16356 (N_16356,N_16138,N_16205);
and U16357 (N_16357,N_15892,N_15042);
and U16358 (N_16358,N_15110,N_15252);
xor U16359 (N_16359,N_15944,N_15850);
nor U16360 (N_16360,N_16071,N_15541);
nand U16361 (N_16361,N_16007,N_15746);
xnor U16362 (N_16362,N_16204,N_15854);
nand U16363 (N_16363,N_16191,N_16156);
or U16364 (N_16364,N_16019,N_15418);
or U16365 (N_16365,N_15219,N_15543);
nor U16366 (N_16366,N_15466,N_15450);
nand U16367 (N_16367,N_16222,N_16195);
xnor U16368 (N_16368,N_15993,N_16244);
nor U16369 (N_16369,N_15086,N_15965);
or U16370 (N_16370,N_15729,N_15545);
or U16371 (N_16371,N_16045,N_15414);
nor U16372 (N_16372,N_15443,N_15469);
and U16373 (N_16373,N_15555,N_15293);
xor U16374 (N_16374,N_15897,N_16145);
or U16375 (N_16375,N_16106,N_15817);
xor U16376 (N_16376,N_15361,N_15348);
nand U16377 (N_16377,N_16163,N_15514);
and U16378 (N_16378,N_16128,N_15233);
and U16379 (N_16379,N_16144,N_15884);
nand U16380 (N_16380,N_15958,N_15762);
or U16381 (N_16381,N_15895,N_15025);
and U16382 (N_16382,N_16157,N_15454);
nor U16383 (N_16383,N_16117,N_16014);
nand U16384 (N_16384,N_15532,N_16186);
nor U16385 (N_16385,N_15191,N_16052);
nand U16386 (N_16386,N_16234,N_15189);
nor U16387 (N_16387,N_15160,N_15148);
or U16388 (N_16388,N_15513,N_15765);
or U16389 (N_16389,N_15180,N_15379);
nand U16390 (N_16390,N_15342,N_15053);
xnor U16391 (N_16391,N_15785,N_16118);
nor U16392 (N_16392,N_15804,N_15587);
nor U16393 (N_16393,N_15404,N_15166);
xor U16394 (N_16394,N_16241,N_15675);
nor U16395 (N_16395,N_16054,N_15117);
nand U16396 (N_16396,N_15128,N_16101);
or U16397 (N_16397,N_15727,N_15096);
nor U16398 (N_16398,N_15839,N_15464);
xnor U16399 (N_16399,N_15205,N_15769);
or U16400 (N_16400,N_16048,N_15406);
nor U16401 (N_16401,N_15125,N_15877);
nand U16402 (N_16402,N_15701,N_15509);
nand U16403 (N_16403,N_15124,N_15660);
or U16404 (N_16404,N_15441,N_16183);
nor U16405 (N_16405,N_16136,N_15569);
xor U16406 (N_16406,N_16239,N_16168);
and U16407 (N_16407,N_16068,N_15733);
xor U16408 (N_16408,N_15393,N_15992);
and U16409 (N_16409,N_15164,N_15260);
and U16410 (N_16410,N_15105,N_15562);
nor U16411 (N_16411,N_15088,N_15534);
nand U16412 (N_16412,N_15168,N_16245);
nor U16413 (N_16413,N_15935,N_15287);
or U16414 (N_16414,N_15305,N_16160);
nand U16415 (N_16415,N_16246,N_15415);
and U16416 (N_16416,N_15819,N_15737);
and U16417 (N_16417,N_16047,N_15020);
xor U16418 (N_16418,N_16077,N_16067);
or U16419 (N_16419,N_15732,N_15387);
xnor U16420 (N_16420,N_15146,N_15671);
xnor U16421 (N_16421,N_15716,N_15927);
xor U16422 (N_16422,N_15031,N_16166);
xnor U16423 (N_16423,N_16172,N_15740);
nand U16424 (N_16424,N_15349,N_15119);
nand U16425 (N_16425,N_15951,N_16194);
and U16426 (N_16426,N_16200,N_15581);
nand U16427 (N_16427,N_15715,N_15616);
or U16428 (N_16428,N_15019,N_15748);
nand U16429 (N_16429,N_16232,N_15656);
nand U16430 (N_16430,N_16176,N_15849);
and U16431 (N_16431,N_15246,N_15793);
xnor U16432 (N_16432,N_15971,N_15797);
nand U16433 (N_16433,N_15577,N_15926);
and U16434 (N_16434,N_15392,N_15327);
or U16435 (N_16435,N_15409,N_15396);
xnor U16436 (N_16436,N_15625,N_15771);
or U16437 (N_16437,N_15565,N_15347);
and U16438 (N_16438,N_15859,N_15181);
or U16439 (N_16439,N_15560,N_15059);
and U16440 (N_16440,N_15250,N_16190);
nor U16441 (N_16441,N_15657,N_15906);
xor U16442 (N_16442,N_15395,N_15786);
nor U16443 (N_16443,N_15068,N_15568);
nor U16444 (N_16444,N_16020,N_15557);
nand U16445 (N_16445,N_15956,N_15145);
nor U16446 (N_16446,N_15843,N_15923);
nand U16447 (N_16447,N_15983,N_16201);
nand U16448 (N_16448,N_16148,N_15519);
nor U16449 (N_16449,N_15790,N_15322);
nand U16450 (N_16450,N_16065,N_16080);
xnor U16451 (N_16451,N_15328,N_16098);
xnor U16452 (N_16452,N_15820,N_16013);
nand U16453 (N_16453,N_16248,N_15801);
or U16454 (N_16454,N_15516,N_16000);
and U16455 (N_16455,N_16018,N_15990);
and U16456 (N_16456,N_15885,N_15719);
or U16457 (N_16457,N_16162,N_15071);
and U16458 (N_16458,N_16100,N_15868);
and U16459 (N_16459,N_15278,N_15987);
nand U16460 (N_16460,N_15352,N_15741);
nor U16461 (N_16461,N_15115,N_15385);
xor U16462 (N_16462,N_15594,N_15083);
xnor U16463 (N_16463,N_15369,N_15072);
nand U16464 (N_16464,N_16240,N_15908);
nor U16465 (N_16465,N_16035,N_16108);
nor U16466 (N_16466,N_15202,N_15034);
nand U16467 (N_16467,N_15274,N_15770);
nor U16468 (N_16468,N_16203,N_16057);
nor U16469 (N_16469,N_15092,N_16212);
or U16470 (N_16470,N_15860,N_15183);
and U16471 (N_16471,N_15380,N_15959);
nand U16472 (N_16472,N_15261,N_15537);
or U16473 (N_16473,N_16179,N_15492);
nand U16474 (N_16474,N_15111,N_15315);
nand U16475 (N_16475,N_15238,N_15773);
nand U16476 (N_16476,N_15190,N_15755);
nand U16477 (N_16477,N_15747,N_15237);
nor U16478 (N_16478,N_15381,N_15978);
xor U16479 (N_16479,N_16093,N_15280);
or U16480 (N_16480,N_15942,N_15389);
nor U16481 (N_16481,N_15997,N_15641);
xnor U16482 (N_16482,N_15970,N_15004);
nand U16483 (N_16483,N_15912,N_15777);
nor U16484 (N_16484,N_15039,N_16139);
and U16485 (N_16485,N_15628,N_15257);
and U16486 (N_16486,N_15915,N_15038);
nand U16487 (N_16487,N_15220,N_15447);
nor U16488 (N_16488,N_15444,N_15154);
nand U16489 (N_16489,N_15200,N_15600);
nor U16490 (N_16490,N_15090,N_15187);
nand U16491 (N_16491,N_15221,N_15386);
and U16492 (N_16492,N_16042,N_15120);
xor U16493 (N_16493,N_15972,N_15033);
xnor U16494 (N_16494,N_15916,N_16229);
or U16495 (N_16495,N_16211,N_15476);
or U16496 (N_16496,N_16095,N_15601);
and U16497 (N_16497,N_15873,N_15832);
nand U16498 (N_16498,N_15835,N_16188);
xnor U16499 (N_16499,N_15789,N_15807);
nand U16500 (N_16500,N_15296,N_15686);
nand U16501 (N_16501,N_15377,N_15340);
xor U16502 (N_16502,N_15667,N_15388);
nand U16503 (N_16503,N_15354,N_15515);
nand U16504 (N_16504,N_15522,N_15831);
nor U16505 (N_16505,N_15210,N_15573);
and U16506 (N_16506,N_16143,N_15056);
nor U16507 (N_16507,N_15412,N_15000);
or U16508 (N_16508,N_15776,N_15979);
xor U16509 (N_16509,N_15351,N_16076);
or U16510 (N_16510,N_15687,N_15330);
and U16511 (N_16511,N_15247,N_15981);
nor U16512 (N_16512,N_15241,N_15855);
nand U16513 (N_16513,N_15575,N_15822);
and U16514 (N_16514,N_15498,N_15886);
and U16515 (N_16515,N_15629,N_15339);
nor U16516 (N_16516,N_15151,N_15234);
nand U16517 (N_16517,N_15761,N_16113);
nor U16518 (N_16518,N_15866,N_15880);
or U16519 (N_16519,N_15325,N_15662);
nand U16520 (N_16520,N_16181,N_15961);
nand U16521 (N_16521,N_15805,N_16125);
nand U16522 (N_16522,N_15689,N_15052);
nand U16523 (N_16523,N_15791,N_16146);
or U16524 (N_16524,N_15604,N_15778);
nand U16525 (N_16525,N_15417,N_15311);
nand U16526 (N_16526,N_15477,N_15029);
nand U16527 (N_16527,N_16009,N_15991);
nand U16528 (N_16528,N_15520,N_15936);
or U16529 (N_16529,N_15374,N_15182);
nand U16530 (N_16530,N_15273,N_16196);
nand U16531 (N_16531,N_16056,N_15730);
nand U16532 (N_16532,N_15962,N_15062);
or U16533 (N_16533,N_15830,N_15268);
or U16534 (N_16534,N_15867,N_15529);
nor U16535 (N_16535,N_15910,N_16088);
nand U16536 (N_16536,N_15888,N_15810);
nand U16537 (N_16537,N_15574,N_16006);
nor U16538 (N_16538,N_15133,N_15207);
xor U16539 (N_16539,N_16126,N_15724);
nor U16540 (N_16540,N_15833,N_15802);
xor U16541 (N_16541,N_15931,N_15538);
nand U16542 (N_16542,N_16026,N_15933);
or U16543 (N_16543,N_15693,N_15792);
nor U16544 (N_16544,N_16141,N_15301);
nor U16545 (N_16545,N_15459,N_16170);
nand U16546 (N_16546,N_16237,N_16221);
nor U16547 (N_16547,N_15813,N_15588);
xnor U16548 (N_16548,N_15319,N_15708);
and U16549 (N_16549,N_15067,N_15431);
nor U16550 (N_16550,N_16001,N_15750);
nand U16551 (N_16551,N_15570,N_15613);
xor U16552 (N_16552,N_15045,N_15760);
nand U16553 (N_16553,N_15087,N_15359);
and U16554 (N_16554,N_15172,N_16079);
or U16555 (N_16555,N_15486,N_15030);
xnor U16556 (N_16556,N_15986,N_16022);
nand U16557 (N_16557,N_15980,N_16090);
nand U16558 (N_16558,N_15528,N_15424);
xnor U16559 (N_16559,N_15277,N_15317);
or U16560 (N_16560,N_15905,N_16010);
nor U16561 (N_16561,N_15114,N_15799);
nand U16562 (N_16562,N_15310,N_15222);
and U16563 (N_16563,N_16210,N_15511);
or U16564 (N_16564,N_16028,N_15139);
xor U16565 (N_16565,N_15851,N_15583);
nor U16566 (N_16566,N_15919,N_15094);
or U16567 (N_16567,N_15470,N_15382);
or U16568 (N_16568,N_15195,N_15403);
nor U16569 (N_16569,N_15367,N_15292);
xor U16570 (N_16570,N_15394,N_15411);
nand U16571 (N_16571,N_15943,N_15279);
and U16572 (N_16572,N_15627,N_15206);
and U16573 (N_16573,N_15940,N_15527);
nand U16574 (N_16574,N_16185,N_15084);
nor U16575 (N_16575,N_15874,N_15245);
nand U16576 (N_16576,N_16213,N_15147);
nor U16577 (N_16577,N_15018,N_15479);
and U16578 (N_16578,N_16074,N_15009);
xnor U16579 (N_16579,N_15300,N_15966);
and U16580 (N_16580,N_15635,N_15607);
xor U16581 (N_16581,N_15680,N_16174);
nand U16582 (N_16582,N_16062,N_15491);
or U16583 (N_16583,N_15298,N_15003);
and U16584 (N_16584,N_15938,N_16033);
and U16585 (N_16585,N_15853,N_15774);
nand U16586 (N_16586,N_15700,N_15413);
nor U16587 (N_16587,N_15112,N_16050);
nor U16588 (N_16588,N_15165,N_15847);
or U16589 (N_16589,N_15609,N_15218);
nand U16590 (N_16590,N_15127,N_15463);
nand U16591 (N_16591,N_15610,N_15669);
nor U16592 (N_16592,N_15879,N_15767);
or U16593 (N_16593,N_15297,N_15093);
and U16594 (N_16594,N_15370,N_15224);
or U16595 (N_16595,N_16153,N_15870);
nor U16596 (N_16596,N_16164,N_15193);
xor U16597 (N_16597,N_15652,N_16096);
and U16598 (N_16598,N_15705,N_15063);
or U16599 (N_16599,N_15896,N_16182);
xnor U16600 (N_16600,N_15651,N_15064);
nand U16601 (N_16601,N_15002,N_15579);
xnor U16602 (N_16602,N_15284,N_15924);
xor U16603 (N_16603,N_15932,N_15756);
xor U16604 (N_16604,N_15848,N_15324);
nor U16605 (N_16605,N_16142,N_15974);
xor U16606 (N_16606,N_16111,N_15505);
or U16607 (N_16607,N_15442,N_15670);
nor U16608 (N_16608,N_15592,N_15371);
nand U16609 (N_16609,N_15089,N_15350);
nand U16610 (N_16610,N_15326,N_16005);
nand U16611 (N_16611,N_15286,N_15973);
xor U16612 (N_16612,N_16220,N_15338);
or U16613 (N_16613,N_15254,N_15137);
xor U16614 (N_16614,N_15333,N_15345);
nand U16615 (N_16615,N_16029,N_16147);
xnor U16616 (N_16616,N_15037,N_15898);
xnor U16617 (N_16617,N_16171,N_15901);
and U16618 (N_16618,N_15952,N_15129);
xnor U16619 (N_16619,N_15057,N_16114);
nand U16620 (N_16620,N_15739,N_15876);
nor U16621 (N_16621,N_15863,N_16086);
nand U16622 (N_16622,N_15967,N_15170);
or U16623 (N_16623,N_15134,N_15065);
nand U16624 (N_16624,N_16208,N_15964);
or U16625 (N_16625,N_15391,N_15512);
nand U16626 (N_16626,N_15934,N_15457);
nand U16627 (N_16627,N_15098,N_16046);
xnor U16628 (N_16628,N_15375,N_16044);
nor U16629 (N_16629,N_15204,N_15303);
or U16630 (N_16630,N_16023,N_15818);
xor U16631 (N_16631,N_15757,N_15533);
xor U16632 (N_16632,N_16127,N_15426);
nand U16633 (N_16633,N_15438,N_15914);
and U16634 (N_16634,N_15678,N_15421);
and U16635 (N_16635,N_15698,N_15542);
nor U16636 (N_16636,N_15085,N_15073);
or U16637 (N_16637,N_15427,N_15862);
nand U16638 (N_16638,N_15323,N_16133);
and U16639 (N_16639,N_15535,N_15903);
and U16640 (N_16640,N_15531,N_16135);
xor U16641 (N_16641,N_15561,N_15256);
xnor U16642 (N_16642,N_15639,N_15695);
nor U16643 (N_16643,N_15696,N_16227);
or U16644 (N_16644,N_15471,N_15401);
xor U16645 (N_16645,N_15467,N_16215);
xor U16646 (N_16646,N_15163,N_15954);
xor U16647 (N_16647,N_15016,N_15706);
nand U16648 (N_16648,N_15517,N_15365);
nand U16649 (N_16649,N_15075,N_15677);
nand U16650 (N_16650,N_15044,N_15364);
and U16651 (N_16651,N_16103,N_15823);
xor U16652 (N_16652,N_15871,N_15416);
nand U16653 (N_16653,N_15960,N_15977);
nand U16654 (N_16654,N_15963,N_15857);
and U16655 (N_16655,N_15355,N_15449);
or U16656 (N_16656,N_15232,N_15215);
xnor U16657 (N_16657,N_15726,N_15598);
and U16658 (N_16658,N_15262,N_15825);
nand U16659 (N_16659,N_16040,N_15138);
and U16660 (N_16660,N_15889,N_15473);
and U16661 (N_16661,N_16175,N_15586);
xor U16662 (N_16662,N_15614,N_15720);
xor U16663 (N_16663,N_16206,N_15713);
nor U16664 (N_16664,N_15882,N_15654);
nor U16665 (N_16665,N_15108,N_15161);
and U16666 (N_16666,N_15887,N_15271);
or U16667 (N_16667,N_16155,N_15131);
and U16668 (N_16668,N_15081,N_15690);
xnor U16669 (N_16669,N_15618,N_15214);
nor U16670 (N_16670,N_16003,N_16017);
or U16671 (N_16671,N_15702,N_15728);
and U16672 (N_16672,N_15731,N_15015);
and U16673 (N_16673,N_15780,N_16032);
nand U16674 (N_16674,N_15872,N_15530);
or U16675 (N_16675,N_15925,N_15314);
nor U16676 (N_16676,N_15308,N_15225);
and U16677 (N_16677,N_15620,N_15171);
or U16678 (N_16678,N_15196,N_16031);
nand U16679 (N_16679,N_15299,N_15468);
nor U16680 (N_16680,N_15794,N_15643);
xnor U16681 (N_16681,N_15048,N_16224);
or U16682 (N_16682,N_16121,N_15590);
and U16683 (N_16683,N_15307,N_15102);
and U16684 (N_16684,N_15869,N_15968);
nand U16685 (N_16685,N_15852,N_16231);
or U16686 (N_16686,N_15798,N_15521);
or U16687 (N_16687,N_15313,N_15602);
nor U16688 (N_16688,N_16161,N_15209);
xor U16689 (N_16689,N_15036,N_15544);
or U16690 (N_16690,N_15448,N_15496);
or U16691 (N_16691,N_15249,N_15023);
xor U16692 (N_16692,N_16078,N_15665);
nor U16693 (N_16693,N_15433,N_15306);
and U16694 (N_16694,N_15244,N_15937);
nand U16695 (N_16695,N_15434,N_15772);
or U16696 (N_16696,N_15346,N_15211);
and U16697 (N_16697,N_15712,N_15400);
nand U16698 (N_16698,N_16151,N_15865);
xor U16699 (N_16699,N_16226,N_15946);
or U16700 (N_16700,N_15672,N_15674);
and U16701 (N_16701,N_15360,N_15704);
or U16702 (N_16702,N_16123,N_16134);
xor U16703 (N_16703,N_15768,N_15572);
xnor U16704 (N_16704,N_15316,N_15563);
or U16705 (N_16705,N_15483,N_15402);
or U16706 (N_16706,N_15929,N_15595);
xnor U16707 (N_16707,N_15061,N_15107);
and U16708 (N_16708,N_16247,N_15472);
and U16709 (N_16709,N_15692,N_15751);
nand U16710 (N_16710,N_15331,N_16217);
or U16711 (N_16711,N_15497,N_15647);
and U16712 (N_16712,N_15815,N_15995);
nand U16713 (N_16713,N_15357,N_15201);
nor U16714 (N_16714,N_15227,N_15845);
nand U16715 (N_16715,N_15718,N_15372);
nor U16716 (N_16716,N_16228,N_15123);
or U16717 (N_16717,N_15405,N_15939);
nand U16718 (N_16718,N_15640,N_16053);
xnor U16719 (N_16719,N_15155,N_15578);
or U16720 (N_16720,N_15055,N_16002);
or U16721 (N_16721,N_16049,N_15524);
and U16722 (N_16722,N_15101,N_16209);
nand U16723 (N_16723,N_15988,N_15309);
nor U16724 (N_16724,N_16219,N_15883);
and U16725 (N_16725,N_15078,N_15742);
and U16726 (N_16726,N_15838,N_15891);
and U16727 (N_16727,N_15673,N_15894);
and U16728 (N_16728,N_15582,N_15645);
nand U16729 (N_16729,N_15861,N_15358);
nand U16730 (N_16730,N_15811,N_15179);
nor U16731 (N_16731,N_15683,N_15622);
or U16732 (N_16732,N_15028,N_15829);
nor U16733 (N_16733,N_15553,N_15080);
or U16734 (N_16734,N_15461,N_15709);
nand U16735 (N_16735,N_16015,N_16218);
xor U16736 (N_16736,N_15546,N_15240);
nand U16737 (N_16737,N_16092,N_15366);
or U16738 (N_16738,N_15440,N_16058);
nor U16739 (N_16739,N_15337,N_15593);
or U16740 (N_16740,N_15808,N_15235);
and U16741 (N_16741,N_15548,N_16055);
and U16742 (N_16742,N_15911,N_15691);
nor U16743 (N_16743,N_15812,N_15109);
and U16744 (N_16744,N_15103,N_15489);
nand U16745 (N_16745,N_15552,N_15143);
or U16746 (N_16746,N_15456,N_15549);
nand U16747 (N_16747,N_15788,N_15295);
xnor U16748 (N_16748,N_16129,N_15420);
nand U16749 (N_16749,N_15821,N_15011);
nor U16750 (N_16750,N_15079,N_15759);
nand U16751 (N_16751,N_15253,N_15226);
and U16752 (N_16752,N_16238,N_15599);
xnor U16753 (N_16753,N_16225,N_16070);
or U16754 (N_16754,N_15899,N_16137);
nand U16755 (N_16755,N_15738,N_15026);
xor U16756 (N_16756,N_15653,N_15255);
or U16757 (N_16757,N_15485,N_15638);
or U16758 (N_16758,N_16193,N_15208);
and U16759 (N_16759,N_15184,N_15707);
xor U16760 (N_16760,N_15764,N_15013);
nand U16761 (N_16761,N_15659,N_15158);
and U16762 (N_16762,N_15725,N_15251);
or U16763 (N_16763,N_16230,N_16102);
xor U16764 (N_16764,N_15149,N_15194);
or U16765 (N_16765,N_15710,N_15229);
or U16766 (N_16766,N_15334,N_15558);
nor U16767 (N_16767,N_15540,N_16081);
nor U16768 (N_16768,N_15142,N_15775);
xnor U16769 (N_16769,N_15893,N_15091);
xnor U16770 (N_16770,N_15989,N_15984);
or U16771 (N_16771,N_15763,N_15668);
nor U16772 (N_16772,N_15945,N_16140);
nand U16773 (N_16773,N_16107,N_15289);
xnor U16774 (N_16774,N_15828,N_15663);
and U16775 (N_16775,N_15554,N_16150);
nand U16776 (N_16776,N_16192,N_16152);
nand U16777 (N_16777,N_15566,N_15611);
and U16778 (N_16778,N_15144,N_15766);
nand U16779 (N_16779,N_15283,N_15559);
and U16780 (N_16780,N_15050,N_16094);
nand U16781 (N_16781,N_15881,N_15518);
or U16782 (N_16782,N_16064,N_15077);
and U16783 (N_16783,N_15488,N_16061);
nor U16784 (N_16784,N_16083,N_15605);
xnor U16785 (N_16785,N_15152,N_15051);
or U16786 (N_16786,N_16124,N_15722);
nor U16787 (N_16787,N_15648,N_16119);
and U16788 (N_16788,N_15969,N_15957);
xor U16789 (N_16789,N_15174,N_15376);
or U16790 (N_16790,N_15452,N_15949);
and U16791 (N_16791,N_16087,N_15320);
nand U16792 (N_16792,N_16039,N_15267);
and U16793 (N_16793,N_16235,N_15584);
and U16794 (N_16794,N_15399,N_15258);
and U16795 (N_16795,N_16034,N_15721);
and U16796 (N_16796,N_15633,N_16178);
and U16797 (N_16797,N_15032,N_15858);
nand U16798 (N_16798,N_16072,N_16159);
nand U16799 (N_16799,N_15806,N_15264);
xor U16800 (N_16800,N_15637,N_15176);
nand U16801 (N_16801,N_15021,N_15113);
and U16802 (N_16802,N_15410,N_15982);
nor U16803 (N_16803,N_15270,N_15236);
nor U16804 (N_16804,N_15186,N_15321);
and U16805 (N_16805,N_16037,N_16173);
nand U16806 (N_16806,N_15589,N_15429);
and U16807 (N_16807,N_15650,N_15630);
or U16808 (N_16808,N_15917,N_16198);
nand U16809 (N_16809,N_16249,N_15281);
and U16810 (N_16810,N_15734,N_15658);
nand U16811 (N_16811,N_15523,N_15192);
or U16812 (N_16812,N_15266,N_15875);
nor U16813 (N_16813,N_15304,N_15199);
nor U16814 (N_16814,N_15576,N_15212);
and U16815 (N_16815,N_16012,N_15909);
or U16816 (N_16816,N_16187,N_15294);
and U16817 (N_16817,N_15526,N_15460);
xnor U16818 (N_16818,N_15617,N_15950);
xor U16819 (N_16819,N_15921,N_15508);
nand U16820 (N_16820,N_15481,N_15503);
xor U16821 (N_16821,N_15213,N_15104);
and U16822 (N_16822,N_15490,N_15159);
nand U16823 (N_16823,N_15445,N_15265);
xor U16824 (N_16824,N_15501,N_16105);
and U16825 (N_16825,N_15844,N_16112);
and U16826 (N_16826,N_15291,N_15362);
nor U16827 (N_16827,N_16169,N_15636);
or U16828 (N_16828,N_15580,N_16165);
or U16829 (N_16829,N_15539,N_15288);
nand U16830 (N_16830,N_15507,N_15996);
nor U16831 (N_16831,N_15453,N_15439);
xnor U16832 (N_16832,N_15228,N_15335);
nand U16833 (N_16833,N_15655,N_15495);
xnor U16834 (N_16834,N_15753,N_15597);
or U16835 (N_16835,N_16021,N_15621);
nor U16836 (N_16836,N_15318,N_16069);
xor U16837 (N_16837,N_15800,N_15661);
nor U16838 (N_16838,N_15591,N_15231);
nand U16839 (N_16839,N_16025,N_16043);
and U16840 (N_16840,N_16085,N_16216);
and U16841 (N_16841,N_15049,N_16099);
nand U16842 (N_16842,N_15312,N_15836);
and U16843 (N_16843,N_15619,N_15510);
or U16844 (N_16844,N_15890,N_16207);
nand U16845 (N_16845,N_15272,N_15480);
nand U16846 (N_16846,N_15556,N_16084);
and U16847 (N_16847,N_15735,N_15436);
xnor U16848 (N_16848,N_15223,N_15494);
nor U16849 (N_16849,N_15752,N_15536);
and U16850 (N_16850,N_15046,N_15699);
nand U16851 (N_16851,N_15006,N_15040);
xnor U16852 (N_16852,N_15953,N_15343);
nor U16853 (N_16853,N_15012,N_15684);
or U16854 (N_16854,N_16223,N_15666);
and U16855 (N_16855,N_15783,N_15624);
and U16856 (N_16856,N_16109,N_15904);
xor U16857 (N_16857,N_16110,N_15551);
xor U16858 (N_16858,N_15259,N_16041);
xnor U16859 (N_16859,N_15976,N_15197);
or U16860 (N_16860,N_15076,N_15302);
and U16861 (N_16861,N_15714,N_15493);
nor U16862 (N_16862,N_15685,N_16189);
and U16863 (N_16863,N_15437,N_16008);
and U16864 (N_16864,N_15263,N_15007);
and U16865 (N_16865,N_16177,N_16036);
nand U16866 (N_16866,N_16158,N_15816);
nand U16867 (N_16867,N_15217,N_15612);
nand U16868 (N_16868,N_16016,N_15408);
xnor U16869 (N_16869,N_16063,N_16104);
xor U16870 (N_16870,N_16059,N_16180);
and U16871 (N_16871,N_15363,N_15099);
nand U16872 (N_16872,N_15795,N_15902);
nor U16873 (N_16873,N_15632,N_15941);
and U16874 (N_16874,N_15425,N_15008);
nand U16875 (N_16875,N_15672,N_15472);
nor U16876 (N_16876,N_16113,N_15252);
nand U16877 (N_16877,N_15357,N_15118);
or U16878 (N_16878,N_15438,N_15326);
and U16879 (N_16879,N_16011,N_15252);
or U16880 (N_16880,N_16234,N_15687);
nor U16881 (N_16881,N_15305,N_15314);
nand U16882 (N_16882,N_15573,N_15575);
nor U16883 (N_16883,N_15173,N_16176);
and U16884 (N_16884,N_15795,N_15456);
nor U16885 (N_16885,N_16200,N_15903);
nor U16886 (N_16886,N_16180,N_16227);
nand U16887 (N_16887,N_16249,N_15575);
and U16888 (N_16888,N_15261,N_15525);
nand U16889 (N_16889,N_16058,N_15630);
or U16890 (N_16890,N_15818,N_15154);
xor U16891 (N_16891,N_15704,N_15531);
or U16892 (N_16892,N_15601,N_15196);
nor U16893 (N_16893,N_15381,N_16094);
nor U16894 (N_16894,N_15994,N_15804);
nand U16895 (N_16895,N_15512,N_15772);
and U16896 (N_16896,N_15409,N_15929);
or U16897 (N_16897,N_16123,N_15848);
or U16898 (N_16898,N_15833,N_15340);
nand U16899 (N_16899,N_15216,N_15391);
nand U16900 (N_16900,N_16205,N_16012);
xor U16901 (N_16901,N_16241,N_15558);
nor U16902 (N_16902,N_15103,N_15261);
xnor U16903 (N_16903,N_15641,N_15924);
or U16904 (N_16904,N_15464,N_15884);
xor U16905 (N_16905,N_16156,N_16142);
xor U16906 (N_16906,N_15634,N_15065);
and U16907 (N_16907,N_15154,N_15242);
nor U16908 (N_16908,N_15596,N_15609);
and U16909 (N_16909,N_16136,N_16065);
nor U16910 (N_16910,N_15261,N_15437);
nand U16911 (N_16911,N_15469,N_16209);
nand U16912 (N_16912,N_15614,N_16001);
and U16913 (N_16913,N_15058,N_15076);
nand U16914 (N_16914,N_15409,N_15890);
xnor U16915 (N_16915,N_15311,N_15200);
nand U16916 (N_16916,N_15238,N_15918);
and U16917 (N_16917,N_15208,N_15107);
xnor U16918 (N_16918,N_16058,N_15032);
nor U16919 (N_16919,N_15147,N_15195);
xnor U16920 (N_16920,N_15792,N_15869);
and U16921 (N_16921,N_15849,N_15876);
or U16922 (N_16922,N_15649,N_16026);
nor U16923 (N_16923,N_15731,N_16064);
xor U16924 (N_16924,N_15717,N_16059);
xor U16925 (N_16925,N_15329,N_15528);
and U16926 (N_16926,N_15435,N_16013);
nand U16927 (N_16927,N_15649,N_15560);
nor U16928 (N_16928,N_15177,N_15302);
xor U16929 (N_16929,N_16189,N_15624);
xor U16930 (N_16930,N_15672,N_15256);
nor U16931 (N_16931,N_16092,N_15548);
and U16932 (N_16932,N_15596,N_16186);
or U16933 (N_16933,N_15802,N_15791);
xor U16934 (N_16934,N_15392,N_16172);
xnor U16935 (N_16935,N_15287,N_15993);
or U16936 (N_16936,N_15816,N_15374);
nand U16937 (N_16937,N_16060,N_15507);
or U16938 (N_16938,N_15998,N_15611);
or U16939 (N_16939,N_15152,N_15594);
nor U16940 (N_16940,N_15454,N_16113);
nand U16941 (N_16941,N_15124,N_15048);
nand U16942 (N_16942,N_15087,N_15000);
nand U16943 (N_16943,N_15063,N_15278);
xor U16944 (N_16944,N_15678,N_16169);
nor U16945 (N_16945,N_15410,N_16137);
or U16946 (N_16946,N_15429,N_15450);
xnor U16947 (N_16947,N_16018,N_15855);
nor U16948 (N_16948,N_15966,N_15307);
nand U16949 (N_16949,N_16048,N_15008);
xor U16950 (N_16950,N_15530,N_15227);
nand U16951 (N_16951,N_15974,N_16007);
nand U16952 (N_16952,N_15932,N_15677);
nor U16953 (N_16953,N_15022,N_15458);
nor U16954 (N_16954,N_16196,N_15590);
nor U16955 (N_16955,N_15787,N_16206);
and U16956 (N_16956,N_15136,N_16086);
or U16957 (N_16957,N_15672,N_15486);
nand U16958 (N_16958,N_15355,N_15789);
xnor U16959 (N_16959,N_16163,N_16207);
xor U16960 (N_16960,N_15549,N_16151);
nand U16961 (N_16961,N_15003,N_15018);
and U16962 (N_16962,N_15667,N_15608);
nor U16963 (N_16963,N_15181,N_15756);
xnor U16964 (N_16964,N_16197,N_16165);
nor U16965 (N_16965,N_15742,N_15699);
nand U16966 (N_16966,N_15682,N_15870);
and U16967 (N_16967,N_15337,N_15045);
nand U16968 (N_16968,N_16239,N_15900);
nand U16969 (N_16969,N_15994,N_16150);
xnor U16970 (N_16970,N_16229,N_15818);
xor U16971 (N_16971,N_15326,N_16019);
and U16972 (N_16972,N_15475,N_15858);
and U16973 (N_16973,N_15794,N_15339);
xor U16974 (N_16974,N_15036,N_15447);
nor U16975 (N_16975,N_15451,N_15525);
or U16976 (N_16976,N_15599,N_15237);
nor U16977 (N_16977,N_15969,N_15935);
or U16978 (N_16978,N_15331,N_15727);
or U16979 (N_16979,N_15687,N_15710);
xor U16980 (N_16980,N_15442,N_15911);
and U16981 (N_16981,N_15275,N_15777);
nor U16982 (N_16982,N_15395,N_15149);
or U16983 (N_16983,N_15443,N_16122);
or U16984 (N_16984,N_15312,N_15876);
nand U16985 (N_16985,N_15017,N_15090);
or U16986 (N_16986,N_15396,N_16221);
nor U16987 (N_16987,N_15721,N_15727);
xor U16988 (N_16988,N_15687,N_15482);
nor U16989 (N_16989,N_16173,N_15088);
or U16990 (N_16990,N_15521,N_16228);
xnor U16991 (N_16991,N_15181,N_15676);
or U16992 (N_16992,N_15062,N_15937);
or U16993 (N_16993,N_16094,N_15871);
xor U16994 (N_16994,N_15236,N_15366);
nor U16995 (N_16995,N_15730,N_16104);
xor U16996 (N_16996,N_15846,N_15360);
nand U16997 (N_16997,N_16092,N_16156);
xor U16998 (N_16998,N_15679,N_15779);
and U16999 (N_16999,N_16068,N_16009);
or U17000 (N_17000,N_16116,N_15503);
and U17001 (N_17001,N_15111,N_15044);
nand U17002 (N_17002,N_15539,N_15706);
and U17003 (N_17003,N_15125,N_15963);
xnor U17004 (N_17004,N_16122,N_15032);
or U17005 (N_17005,N_15028,N_15440);
xor U17006 (N_17006,N_15988,N_15867);
and U17007 (N_17007,N_15180,N_15157);
nor U17008 (N_17008,N_15192,N_15718);
xor U17009 (N_17009,N_16157,N_15758);
nand U17010 (N_17010,N_15880,N_16029);
nand U17011 (N_17011,N_15491,N_15730);
nand U17012 (N_17012,N_15273,N_16050);
nand U17013 (N_17013,N_15351,N_15251);
or U17014 (N_17014,N_15301,N_15166);
or U17015 (N_17015,N_16063,N_16246);
and U17016 (N_17016,N_15466,N_15821);
nor U17017 (N_17017,N_15754,N_15782);
and U17018 (N_17018,N_15910,N_15839);
nor U17019 (N_17019,N_15975,N_16141);
nor U17020 (N_17020,N_15456,N_15840);
or U17021 (N_17021,N_16174,N_15878);
xor U17022 (N_17022,N_15174,N_15699);
nand U17023 (N_17023,N_15640,N_15209);
nor U17024 (N_17024,N_15842,N_15692);
and U17025 (N_17025,N_15917,N_15303);
or U17026 (N_17026,N_15112,N_15861);
nor U17027 (N_17027,N_16128,N_15329);
nand U17028 (N_17028,N_15707,N_15053);
and U17029 (N_17029,N_16137,N_15032);
or U17030 (N_17030,N_15906,N_16174);
nand U17031 (N_17031,N_15022,N_15788);
xor U17032 (N_17032,N_15394,N_15168);
nor U17033 (N_17033,N_16244,N_15460);
or U17034 (N_17034,N_16229,N_15281);
nand U17035 (N_17035,N_16077,N_16160);
nand U17036 (N_17036,N_15165,N_16013);
nand U17037 (N_17037,N_16202,N_16064);
nand U17038 (N_17038,N_15954,N_15097);
nand U17039 (N_17039,N_15126,N_16146);
xor U17040 (N_17040,N_15113,N_15747);
and U17041 (N_17041,N_15195,N_16150);
xnor U17042 (N_17042,N_15627,N_16052);
nor U17043 (N_17043,N_16061,N_15988);
and U17044 (N_17044,N_16167,N_15258);
nand U17045 (N_17045,N_15718,N_15920);
or U17046 (N_17046,N_15654,N_15438);
nor U17047 (N_17047,N_15718,N_15464);
xor U17048 (N_17048,N_15078,N_16226);
and U17049 (N_17049,N_15654,N_15640);
or U17050 (N_17050,N_15103,N_16079);
or U17051 (N_17051,N_15374,N_16115);
xor U17052 (N_17052,N_15037,N_15210);
nand U17053 (N_17053,N_15739,N_15941);
or U17054 (N_17054,N_15442,N_15785);
nand U17055 (N_17055,N_15164,N_16191);
or U17056 (N_17056,N_15711,N_15237);
or U17057 (N_17057,N_15660,N_16167);
nor U17058 (N_17058,N_16229,N_15052);
nand U17059 (N_17059,N_16014,N_15374);
nor U17060 (N_17060,N_15757,N_15926);
nand U17061 (N_17061,N_15062,N_15477);
nand U17062 (N_17062,N_15196,N_15251);
xor U17063 (N_17063,N_15857,N_15777);
nand U17064 (N_17064,N_15103,N_15122);
nand U17065 (N_17065,N_15048,N_15121);
or U17066 (N_17066,N_15767,N_16207);
nor U17067 (N_17067,N_15202,N_15409);
nor U17068 (N_17068,N_16052,N_15194);
and U17069 (N_17069,N_15245,N_15768);
and U17070 (N_17070,N_15702,N_15130);
and U17071 (N_17071,N_15288,N_15412);
or U17072 (N_17072,N_15016,N_15147);
xor U17073 (N_17073,N_15232,N_15908);
xor U17074 (N_17074,N_15478,N_15942);
or U17075 (N_17075,N_16171,N_15494);
or U17076 (N_17076,N_15705,N_15890);
xor U17077 (N_17077,N_15847,N_15831);
or U17078 (N_17078,N_16077,N_16050);
nand U17079 (N_17079,N_15806,N_15455);
or U17080 (N_17080,N_16115,N_16011);
and U17081 (N_17081,N_15567,N_15042);
and U17082 (N_17082,N_15096,N_15212);
xor U17083 (N_17083,N_15005,N_15511);
nand U17084 (N_17084,N_16042,N_16052);
xnor U17085 (N_17085,N_15725,N_15310);
and U17086 (N_17086,N_16035,N_15888);
nand U17087 (N_17087,N_15035,N_15946);
nor U17088 (N_17088,N_15346,N_15073);
nor U17089 (N_17089,N_15373,N_15846);
and U17090 (N_17090,N_16244,N_15347);
nor U17091 (N_17091,N_16148,N_15370);
nand U17092 (N_17092,N_15260,N_15473);
nand U17093 (N_17093,N_15957,N_15664);
nor U17094 (N_17094,N_16019,N_15857);
nand U17095 (N_17095,N_15452,N_15793);
or U17096 (N_17096,N_15961,N_15051);
nand U17097 (N_17097,N_15735,N_15344);
nand U17098 (N_17098,N_16055,N_15137);
and U17099 (N_17099,N_15080,N_16064);
xor U17100 (N_17100,N_16105,N_15415);
and U17101 (N_17101,N_15465,N_15079);
or U17102 (N_17102,N_15401,N_15461);
xnor U17103 (N_17103,N_15604,N_15520);
and U17104 (N_17104,N_15920,N_15863);
nand U17105 (N_17105,N_15294,N_16052);
nand U17106 (N_17106,N_15158,N_15741);
xnor U17107 (N_17107,N_15539,N_16110);
xor U17108 (N_17108,N_15725,N_15878);
xor U17109 (N_17109,N_15314,N_15829);
nor U17110 (N_17110,N_15066,N_16078);
nand U17111 (N_17111,N_15959,N_15939);
and U17112 (N_17112,N_15425,N_15788);
and U17113 (N_17113,N_15759,N_16139);
or U17114 (N_17114,N_15887,N_15600);
and U17115 (N_17115,N_15142,N_15167);
xor U17116 (N_17116,N_16217,N_16048);
nand U17117 (N_17117,N_15562,N_15592);
or U17118 (N_17118,N_15000,N_16000);
nor U17119 (N_17119,N_15948,N_15599);
or U17120 (N_17120,N_15410,N_15032);
xnor U17121 (N_17121,N_15105,N_15175);
nand U17122 (N_17122,N_15826,N_15441);
nand U17123 (N_17123,N_15857,N_15691);
nand U17124 (N_17124,N_15205,N_16104);
and U17125 (N_17125,N_15224,N_16016);
and U17126 (N_17126,N_15033,N_15336);
nor U17127 (N_17127,N_15734,N_16152);
and U17128 (N_17128,N_16118,N_15042);
or U17129 (N_17129,N_15982,N_15100);
or U17130 (N_17130,N_16089,N_15995);
or U17131 (N_17131,N_15650,N_15137);
and U17132 (N_17132,N_15260,N_15188);
nand U17133 (N_17133,N_15736,N_15068);
nand U17134 (N_17134,N_15267,N_16224);
and U17135 (N_17135,N_15155,N_15330);
nor U17136 (N_17136,N_15171,N_15320);
and U17137 (N_17137,N_15918,N_15866);
nor U17138 (N_17138,N_16161,N_15680);
xnor U17139 (N_17139,N_15952,N_15541);
or U17140 (N_17140,N_16143,N_16135);
and U17141 (N_17141,N_15325,N_15699);
or U17142 (N_17142,N_15365,N_16036);
or U17143 (N_17143,N_15735,N_16041);
xor U17144 (N_17144,N_15677,N_15610);
xor U17145 (N_17145,N_15909,N_15404);
and U17146 (N_17146,N_15108,N_15530);
nand U17147 (N_17147,N_15661,N_15854);
nand U17148 (N_17148,N_15718,N_15831);
nor U17149 (N_17149,N_15717,N_15190);
nand U17150 (N_17150,N_15574,N_16240);
nor U17151 (N_17151,N_15970,N_15684);
xor U17152 (N_17152,N_15484,N_15448);
or U17153 (N_17153,N_15265,N_15149);
or U17154 (N_17154,N_15678,N_15687);
xor U17155 (N_17155,N_16176,N_15007);
xor U17156 (N_17156,N_15435,N_15388);
nand U17157 (N_17157,N_16095,N_15884);
or U17158 (N_17158,N_15027,N_15021);
or U17159 (N_17159,N_16118,N_16045);
nand U17160 (N_17160,N_15055,N_15251);
xor U17161 (N_17161,N_15763,N_15137);
nor U17162 (N_17162,N_15761,N_15058);
or U17163 (N_17163,N_15581,N_15693);
nand U17164 (N_17164,N_15557,N_15211);
or U17165 (N_17165,N_15934,N_15452);
and U17166 (N_17166,N_15836,N_16248);
nor U17167 (N_17167,N_15222,N_15758);
and U17168 (N_17168,N_15751,N_15618);
nor U17169 (N_17169,N_15342,N_15742);
xnor U17170 (N_17170,N_15522,N_16112);
or U17171 (N_17171,N_16132,N_15156);
nor U17172 (N_17172,N_16170,N_15423);
nor U17173 (N_17173,N_16203,N_15654);
nand U17174 (N_17174,N_15650,N_15471);
xnor U17175 (N_17175,N_15108,N_15607);
and U17176 (N_17176,N_15640,N_16054);
nor U17177 (N_17177,N_16173,N_16127);
nand U17178 (N_17178,N_15500,N_16125);
nand U17179 (N_17179,N_16167,N_15935);
nand U17180 (N_17180,N_16074,N_15157);
nand U17181 (N_17181,N_15446,N_15395);
xnor U17182 (N_17182,N_15747,N_15622);
and U17183 (N_17183,N_16214,N_16012);
and U17184 (N_17184,N_15181,N_16160);
nor U17185 (N_17185,N_15140,N_15837);
nor U17186 (N_17186,N_15020,N_15498);
or U17187 (N_17187,N_15632,N_15063);
nand U17188 (N_17188,N_16135,N_15247);
or U17189 (N_17189,N_15845,N_15112);
xnor U17190 (N_17190,N_15684,N_15022);
or U17191 (N_17191,N_15268,N_15220);
or U17192 (N_17192,N_15442,N_16092);
or U17193 (N_17193,N_15133,N_15372);
xnor U17194 (N_17194,N_15345,N_16132);
nor U17195 (N_17195,N_15459,N_15344);
nand U17196 (N_17196,N_15489,N_15288);
nor U17197 (N_17197,N_16226,N_16101);
nand U17198 (N_17198,N_15271,N_16173);
and U17199 (N_17199,N_15813,N_15198);
nand U17200 (N_17200,N_15528,N_16183);
and U17201 (N_17201,N_15757,N_15238);
nand U17202 (N_17202,N_16021,N_15938);
nand U17203 (N_17203,N_15312,N_16069);
xnor U17204 (N_17204,N_15009,N_15620);
and U17205 (N_17205,N_15039,N_15053);
nand U17206 (N_17206,N_15165,N_15274);
and U17207 (N_17207,N_15634,N_15951);
xnor U17208 (N_17208,N_15990,N_15123);
nor U17209 (N_17209,N_15656,N_15713);
nor U17210 (N_17210,N_15936,N_16135);
nor U17211 (N_17211,N_15323,N_15049);
xnor U17212 (N_17212,N_15900,N_16139);
nor U17213 (N_17213,N_15999,N_15368);
xnor U17214 (N_17214,N_15989,N_16159);
and U17215 (N_17215,N_15257,N_15963);
or U17216 (N_17216,N_16057,N_15664);
nor U17217 (N_17217,N_16197,N_15310);
or U17218 (N_17218,N_15934,N_15004);
or U17219 (N_17219,N_15094,N_15206);
or U17220 (N_17220,N_15118,N_15431);
nand U17221 (N_17221,N_15058,N_15583);
nand U17222 (N_17222,N_15967,N_15834);
xor U17223 (N_17223,N_15820,N_15147);
or U17224 (N_17224,N_15420,N_15709);
and U17225 (N_17225,N_15290,N_15308);
nand U17226 (N_17226,N_15310,N_15000);
xor U17227 (N_17227,N_15985,N_16054);
or U17228 (N_17228,N_15081,N_15574);
or U17229 (N_17229,N_15118,N_15784);
or U17230 (N_17230,N_16163,N_16142);
nor U17231 (N_17231,N_15735,N_15853);
and U17232 (N_17232,N_15770,N_15031);
or U17233 (N_17233,N_15698,N_15931);
or U17234 (N_17234,N_16000,N_15878);
or U17235 (N_17235,N_15794,N_16108);
nand U17236 (N_17236,N_15579,N_15041);
and U17237 (N_17237,N_15118,N_15264);
nor U17238 (N_17238,N_15046,N_15360);
nand U17239 (N_17239,N_16204,N_15808);
xor U17240 (N_17240,N_15602,N_15326);
or U17241 (N_17241,N_16055,N_15037);
or U17242 (N_17242,N_15954,N_15025);
nor U17243 (N_17243,N_16079,N_15769);
nand U17244 (N_17244,N_15109,N_15882);
xor U17245 (N_17245,N_16091,N_15287);
or U17246 (N_17246,N_16206,N_15223);
xnor U17247 (N_17247,N_15249,N_15791);
xor U17248 (N_17248,N_16065,N_15190);
and U17249 (N_17249,N_15671,N_15300);
nand U17250 (N_17250,N_15828,N_16188);
nor U17251 (N_17251,N_15464,N_15170);
and U17252 (N_17252,N_15850,N_15009);
or U17253 (N_17253,N_16201,N_15974);
nand U17254 (N_17254,N_16022,N_16010);
nand U17255 (N_17255,N_15749,N_15661);
and U17256 (N_17256,N_15234,N_15795);
or U17257 (N_17257,N_15252,N_15196);
nor U17258 (N_17258,N_15751,N_15587);
nand U17259 (N_17259,N_15808,N_15554);
and U17260 (N_17260,N_15995,N_15172);
nand U17261 (N_17261,N_15618,N_15386);
xnor U17262 (N_17262,N_15875,N_15704);
or U17263 (N_17263,N_15028,N_15204);
nand U17264 (N_17264,N_15206,N_15375);
and U17265 (N_17265,N_15191,N_15221);
xor U17266 (N_17266,N_15534,N_15260);
xor U17267 (N_17267,N_15226,N_16033);
or U17268 (N_17268,N_15958,N_15431);
nor U17269 (N_17269,N_15734,N_15977);
nor U17270 (N_17270,N_15190,N_15258);
and U17271 (N_17271,N_15702,N_15499);
nor U17272 (N_17272,N_15613,N_15574);
and U17273 (N_17273,N_15262,N_15145);
nand U17274 (N_17274,N_15144,N_16234);
and U17275 (N_17275,N_15930,N_15369);
and U17276 (N_17276,N_15794,N_15759);
or U17277 (N_17277,N_15377,N_15474);
nor U17278 (N_17278,N_15855,N_16065);
xor U17279 (N_17279,N_16011,N_15856);
nand U17280 (N_17280,N_15526,N_15317);
or U17281 (N_17281,N_15969,N_16059);
and U17282 (N_17282,N_15857,N_16187);
and U17283 (N_17283,N_15377,N_15273);
nor U17284 (N_17284,N_15085,N_16131);
nor U17285 (N_17285,N_16120,N_15776);
and U17286 (N_17286,N_16061,N_16204);
nand U17287 (N_17287,N_15106,N_16157);
xor U17288 (N_17288,N_16076,N_15352);
xnor U17289 (N_17289,N_15721,N_15276);
nor U17290 (N_17290,N_15144,N_15288);
xnor U17291 (N_17291,N_15111,N_15895);
nor U17292 (N_17292,N_15972,N_15966);
and U17293 (N_17293,N_15978,N_15649);
xor U17294 (N_17294,N_16003,N_15232);
xnor U17295 (N_17295,N_15740,N_15227);
nand U17296 (N_17296,N_15259,N_15750);
nand U17297 (N_17297,N_15240,N_16013);
and U17298 (N_17298,N_15530,N_16145);
and U17299 (N_17299,N_15343,N_16084);
nand U17300 (N_17300,N_15748,N_15800);
nand U17301 (N_17301,N_15753,N_15400);
nand U17302 (N_17302,N_15783,N_15518);
nand U17303 (N_17303,N_15662,N_15579);
xor U17304 (N_17304,N_15400,N_15093);
and U17305 (N_17305,N_16033,N_15455);
xnor U17306 (N_17306,N_15570,N_15412);
nand U17307 (N_17307,N_15540,N_15748);
and U17308 (N_17308,N_15961,N_15249);
and U17309 (N_17309,N_15256,N_15493);
nor U17310 (N_17310,N_15640,N_16190);
nand U17311 (N_17311,N_15654,N_15309);
or U17312 (N_17312,N_15077,N_15641);
or U17313 (N_17313,N_15355,N_15866);
nand U17314 (N_17314,N_15782,N_16153);
or U17315 (N_17315,N_15343,N_15387);
xnor U17316 (N_17316,N_15636,N_15610);
xnor U17317 (N_17317,N_15549,N_15377);
nand U17318 (N_17318,N_15050,N_15269);
xnor U17319 (N_17319,N_15799,N_15397);
and U17320 (N_17320,N_15619,N_16007);
xnor U17321 (N_17321,N_15512,N_16196);
nand U17322 (N_17322,N_16061,N_15733);
nand U17323 (N_17323,N_16167,N_16106);
nand U17324 (N_17324,N_16116,N_16002);
nand U17325 (N_17325,N_16223,N_15806);
nor U17326 (N_17326,N_15884,N_15967);
or U17327 (N_17327,N_15768,N_16041);
nand U17328 (N_17328,N_15179,N_15356);
or U17329 (N_17329,N_15733,N_15993);
and U17330 (N_17330,N_15190,N_15548);
xor U17331 (N_17331,N_16165,N_15989);
nor U17332 (N_17332,N_15465,N_15263);
nor U17333 (N_17333,N_15215,N_15776);
and U17334 (N_17334,N_16044,N_16168);
and U17335 (N_17335,N_16050,N_15818);
xnor U17336 (N_17336,N_15136,N_16208);
or U17337 (N_17337,N_15166,N_16089);
nand U17338 (N_17338,N_15993,N_15054);
and U17339 (N_17339,N_15908,N_15502);
nand U17340 (N_17340,N_16196,N_15881);
nor U17341 (N_17341,N_15711,N_15031);
and U17342 (N_17342,N_16221,N_15116);
nor U17343 (N_17343,N_16129,N_15898);
nand U17344 (N_17344,N_15885,N_15672);
and U17345 (N_17345,N_15653,N_15195);
and U17346 (N_17346,N_15446,N_15746);
and U17347 (N_17347,N_16206,N_15256);
xnor U17348 (N_17348,N_15579,N_15540);
nand U17349 (N_17349,N_15135,N_15201);
xnor U17350 (N_17350,N_16166,N_15601);
and U17351 (N_17351,N_16092,N_15343);
nor U17352 (N_17352,N_15699,N_15134);
and U17353 (N_17353,N_15118,N_15872);
and U17354 (N_17354,N_15702,N_15245);
or U17355 (N_17355,N_16202,N_15073);
nor U17356 (N_17356,N_16060,N_15967);
or U17357 (N_17357,N_16061,N_16079);
or U17358 (N_17358,N_15321,N_15482);
nor U17359 (N_17359,N_15636,N_15124);
nand U17360 (N_17360,N_15791,N_15887);
xnor U17361 (N_17361,N_15829,N_15676);
xor U17362 (N_17362,N_16019,N_15100);
and U17363 (N_17363,N_15175,N_15469);
nand U17364 (N_17364,N_15163,N_15466);
nand U17365 (N_17365,N_15705,N_15162);
xnor U17366 (N_17366,N_15853,N_15824);
xnor U17367 (N_17367,N_15070,N_16142);
and U17368 (N_17368,N_15986,N_15775);
nand U17369 (N_17369,N_16174,N_16134);
and U17370 (N_17370,N_15768,N_16179);
xor U17371 (N_17371,N_15194,N_15230);
nor U17372 (N_17372,N_15505,N_15484);
nor U17373 (N_17373,N_16105,N_15292);
or U17374 (N_17374,N_15529,N_15540);
and U17375 (N_17375,N_15408,N_15208);
and U17376 (N_17376,N_15824,N_15203);
nand U17377 (N_17377,N_15550,N_15334);
nor U17378 (N_17378,N_16095,N_15474);
xor U17379 (N_17379,N_15141,N_15560);
or U17380 (N_17380,N_15705,N_15964);
nand U17381 (N_17381,N_15702,N_15461);
nand U17382 (N_17382,N_15042,N_16085);
xor U17383 (N_17383,N_15756,N_15711);
nor U17384 (N_17384,N_15403,N_15166);
nor U17385 (N_17385,N_15152,N_15379);
xor U17386 (N_17386,N_16115,N_15017);
and U17387 (N_17387,N_15552,N_15876);
nor U17388 (N_17388,N_15578,N_15506);
and U17389 (N_17389,N_15720,N_15531);
xor U17390 (N_17390,N_15142,N_15865);
or U17391 (N_17391,N_15056,N_15162);
xor U17392 (N_17392,N_16088,N_15656);
nor U17393 (N_17393,N_16142,N_15458);
nor U17394 (N_17394,N_16108,N_16153);
and U17395 (N_17395,N_15860,N_15845);
xnor U17396 (N_17396,N_16106,N_15590);
xor U17397 (N_17397,N_15722,N_15610);
xor U17398 (N_17398,N_15097,N_15616);
xor U17399 (N_17399,N_15131,N_16072);
or U17400 (N_17400,N_15022,N_15080);
and U17401 (N_17401,N_15391,N_16229);
or U17402 (N_17402,N_15283,N_15372);
nand U17403 (N_17403,N_16159,N_15524);
or U17404 (N_17404,N_15527,N_15421);
or U17405 (N_17405,N_16231,N_15762);
nor U17406 (N_17406,N_15346,N_15632);
nor U17407 (N_17407,N_15347,N_15741);
or U17408 (N_17408,N_15081,N_15757);
xnor U17409 (N_17409,N_16171,N_16249);
nand U17410 (N_17410,N_15534,N_15588);
and U17411 (N_17411,N_15788,N_15582);
xor U17412 (N_17412,N_15881,N_15379);
nor U17413 (N_17413,N_15885,N_16075);
xnor U17414 (N_17414,N_15699,N_15676);
and U17415 (N_17415,N_15168,N_15332);
nor U17416 (N_17416,N_15872,N_15063);
nor U17417 (N_17417,N_15082,N_15163);
nor U17418 (N_17418,N_15806,N_15943);
nand U17419 (N_17419,N_15343,N_15188);
nor U17420 (N_17420,N_16133,N_15951);
and U17421 (N_17421,N_16194,N_15391);
or U17422 (N_17422,N_16220,N_15623);
xnor U17423 (N_17423,N_15661,N_15123);
xor U17424 (N_17424,N_15181,N_15763);
xnor U17425 (N_17425,N_15673,N_15603);
xor U17426 (N_17426,N_16126,N_16238);
nor U17427 (N_17427,N_15142,N_16094);
nand U17428 (N_17428,N_16039,N_15813);
xor U17429 (N_17429,N_15879,N_15811);
or U17430 (N_17430,N_15895,N_15934);
or U17431 (N_17431,N_15379,N_15582);
nor U17432 (N_17432,N_15855,N_15688);
or U17433 (N_17433,N_15587,N_15894);
or U17434 (N_17434,N_15658,N_15992);
nand U17435 (N_17435,N_15236,N_15010);
and U17436 (N_17436,N_15266,N_15957);
nand U17437 (N_17437,N_15037,N_15943);
nand U17438 (N_17438,N_15498,N_16106);
or U17439 (N_17439,N_15520,N_16159);
or U17440 (N_17440,N_15382,N_16201);
xor U17441 (N_17441,N_15334,N_15275);
or U17442 (N_17442,N_15947,N_15654);
nand U17443 (N_17443,N_15689,N_15988);
and U17444 (N_17444,N_16059,N_15126);
nand U17445 (N_17445,N_16145,N_15247);
xor U17446 (N_17446,N_15830,N_15677);
or U17447 (N_17447,N_15294,N_15720);
nor U17448 (N_17448,N_15991,N_15499);
nor U17449 (N_17449,N_15567,N_16072);
and U17450 (N_17450,N_15340,N_16023);
or U17451 (N_17451,N_15681,N_15236);
nor U17452 (N_17452,N_16193,N_15114);
and U17453 (N_17453,N_16148,N_15731);
and U17454 (N_17454,N_15040,N_15728);
nand U17455 (N_17455,N_15370,N_16168);
or U17456 (N_17456,N_16220,N_15397);
nor U17457 (N_17457,N_15116,N_15159);
and U17458 (N_17458,N_15988,N_15027);
xor U17459 (N_17459,N_16225,N_15964);
nor U17460 (N_17460,N_15811,N_16128);
xor U17461 (N_17461,N_15756,N_16039);
nand U17462 (N_17462,N_15882,N_15556);
nor U17463 (N_17463,N_16110,N_15274);
xor U17464 (N_17464,N_15608,N_15315);
and U17465 (N_17465,N_15663,N_16088);
nor U17466 (N_17466,N_15360,N_15612);
and U17467 (N_17467,N_15148,N_15322);
nand U17468 (N_17468,N_15935,N_15643);
nand U17469 (N_17469,N_15700,N_15415);
and U17470 (N_17470,N_15690,N_15247);
xnor U17471 (N_17471,N_15561,N_15476);
or U17472 (N_17472,N_15369,N_16172);
and U17473 (N_17473,N_15030,N_15018);
nand U17474 (N_17474,N_16002,N_15286);
xor U17475 (N_17475,N_15093,N_15210);
xnor U17476 (N_17476,N_16030,N_15197);
or U17477 (N_17477,N_15343,N_15191);
nand U17478 (N_17478,N_15633,N_16173);
or U17479 (N_17479,N_15555,N_15089);
nand U17480 (N_17480,N_15821,N_15327);
xor U17481 (N_17481,N_15614,N_16066);
or U17482 (N_17482,N_15883,N_15131);
or U17483 (N_17483,N_15517,N_15068);
nand U17484 (N_17484,N_15543,N_15283);
and U17485 (N_17485,N_15188,N_16242);
nand U17486 (N_17486,N_15520,N_16010);
xor U17487 (N_17487,N_16048,N_15556);
nand U17488 (N_17488,N_15330,N_15778);
or U17489 (N_17489,N_15119,N_15491);
xnor U17490 (N_17490,N_15213,N_15752);
nand U17491 (N_17491,N_15770,N_16139);
or U17492 (N_17492,N_15586,N_15576);
or U17493 (N_17493,N_16008,N_15898);
and U17494 (N_17494,N_16233,N_16002);
or U17495 (N_17495,N_16218,N_15111);
nor U17496 (N_17496,N_15798,N_15236);
and U17497 (N_17497,N_15431,N_15979);
and U17498 (N_17498,N_15773,N_16123);
and U17499 (N_17499,N_15452,N_15296);
nand U17500 (N_17500,N_16320,N_16876);
nor U17501 (N_17501,N_16616,N_17000);
xor U17502 (N_17502,N_16689,N_16659);
or U17503 (N_17503,N_16934,N_17482);
or U17504 (N_17504,N_16845,N_17167);
or U17505 (N_17505,N_16313,N_16351);
nor U17506 (N_17506,N_16858,N_16681);
or U17507 (N_17507,N_16540,N_16725);
xor U17508 (N_17508,N_16478,N_16477);
or U17509 (N_17509,N_17194,N_17499);
nand U17510 (N_17510,N_16953,N_16877);
nand U17511 (N_17511,N_17258,N_16976);
xnor U17512 (N_17512,N_16864,N_16278);
xnor U17513 (N_17513,N_17048,N_17139);
and U17514 (N_17514,N_16622,N_17283);
or U17515 (N_17515,N_16441,N_16504);
or U17516 (N_17516,N_17109,N_17134);
and U17517 (N_17517,N_16492,N_17398);
nor U17518 (N_17518,N_16870,N_16533);
nor U17519 (N_17519,N_17219,N_17494);
nor U17520 (N_17520,N_16792,N_17433);
or U17521 (N_17521,N_17376,N_16642);
and U17522 (N_17522,N_16577,N_17133);
nand U17523 (N_17523,N_16493,N_16471);
or U17524 (N_17524,N_16400,N_16502);
nor U17525 (N_17525,N_16838,N_16826);
xor U17526 (N_17526,N_16458,N_16824);
nand U17527 (N_17527,N_16348,N_17047);
and U17528 (N_17528,N_17187,N_17483);
and U17529 (N_17529,N_17214,N_17141);
xnor U17530 (N_17530,N_17299,N_16366);
xnor U17531 (N_17531,N_16703,N_16254);
nand U17532 (N_17532,N_16835,N_16747);
and U17533 (N_17533,N_16874,N_17424);
and U17534 (N_17534,N_16639,N_17367);
and U17535 (N_17535,N_16701,N_16602);
nand U17536 (N_17536,N_16630,N_16500);
nor U17537 (N_17537,N_16572,N_16300);
or U17538 (N_17538,N_16849,N_16922);
or U17539 (N_17539,N_16463,N_17381);
nor U17540 (N_17540,N_17215,N_16940);
or U17541 (N_17541,N_17051,N_17274);
or U17542 (N_17542,N_17041,N_16442);
nor U17543 (N_17543,N_17369,N_16267);
and U17544 (N_17544,N_17289,N_17106);
nor U17545 (N_17545,N_16556,N_17119);
or U17546 (N_17546,N_17102,N_17476);
nor U17547 (N_17547,N_17067,N_16529);
nand U17548 (N_17548,N_17082,N_16739);
nand U17549 (N_17549,N_16633,N_17240);
nor U17550 (N_17550,N_16299,N_16863);
or U17551 (N_17551,N_16880,N_17216);
xor U17552 (N_17552,N_17011,N_16503);
and U17553 (N_17553,N_16798,N_16936);
nor U17554 (N_17554,N_17479,N_17189);
nor U17555 (N_17555,N_17073,N_16872);
xor U17556 (N_17556,N_16855,N_16354);
and U17557 (N_17557,N_17374,N_16722);
nor U17558 (N_17558,N_17137,N_16718);
nor U17559 (N_17559,N_16697,N_16549);
and U17560 (N_17560,N_16668,N_17411);
or U17561 (N_17561,N_17322,N_16850);
nor U17562 (N_17562,N_17326,N_16303);
nor U17563 (N_17563,N_16468,N_17400);
and U17564 (N_17564,N_17370,N_16357);
and U17565 (N_17565,N_17265,N_16494);
nor U17566 (N_17566,N_16524,N_17066);
and U17567 (N_17567,N_16565,N_17111);
or U17568 (N_17568,N_17026,N_16388);
nand U17569 (N_17569,N_16707,N_17282);
and U17570 (N_17570,N_16818,N_17454);
nand U17571 (N_17571,N_17426,N_16617);
or U17572 (N_17572,N_17457,N_17484);
or U17573 (N_17573,N_17065,N_17419);
or U17574 (N_17574,N_16520,N_17081);
and U17575 (N_17575,N_16347,N_17035);
xor U17576 (N_17576,N_16250,N_17447);
nand U17577 (N_17577,N_16365,N_17290);
or U17578 (N_17578,N_17347,N_16614);
nand U17579 (N_17579,N_16414,N_16544);
or U17580 (N_17580,N_16484,N_16685);
and U17581 (N_17581,N_16277,N_17199);
nor U17582 (N_17582,N_16930,N_16412);
nand U17583 (N_17583,N_16432,N_16293);
nand U17584 (N_17584,N_17249,N_17425);
xnor U17585 (N_17585,N_16905,N_16771);
xor U17586 (N_17586,N_16355,N_17163);
and U17587 (N_17587,N_16803,N_16329);
or U17588 (N_17588,N_17180,N_16954);
and U17589 (N_17589,N_16931,N_17383);
nor U17590 (N_17590,N_17360,N_17182);
nor U17591 (N_17591,N_16909,N_16558);
and U17592 (N_17592,N_17059,N_17352);
nor U17593 (N_17593,N_16919,N_17105);
and U17594 (N_17594,N_16847,N_17197);
xor U17595 (N_17595,N_16264,N_16944);
nand U17596 (N_17596,N_17008,N_17452);
and U17597 (N_17597,N_16638,N_16595);
and U17598 (N_17598,N_16472,N_17293);
and U17599 (N_17599,N_17122,N_17003);
or U17600 (N_17600,N_16433,N_16274);
xnor U17601 (N_17601,N_16531,N_16843);
xor U17602 (N_17602,N_16415,N_17377);
and U17603 (N_17603,N_16822,N_16457);
nand U17604 (N_17604,N_17331,N_17438);
or U17605 (N_17605,N_17110,N_17328);
nor U17606 (N_17606,N_17112,N_16810);
xor U17607 (N_17607,N_16527,N_17344);
nor U17608 (N_17608,N_17224,N_16596);
xor U17609 (N_17609,N_17034,N_17399);
xnor U17610 (N_17610,N_16435,N_17261);
or U17611 (N_17611,N_17267,N_16383);
nand U17612 (N_17612,N_16997,N_17028);
or U17613 (N_17613,N_17001,N_17055);
nor U17614 (N_17614,N_16839,N_17121);
nor U17615 (N_17615,N_16598,N_16330);
or U17616 (N_17616,N_17190,N_16555);
or U17617 (N_17617,N_17470,N_17253);
and U17618 (N_17618,N_17286,N_16653);
and U17619 (N_17619,N_17225,N_16604);
and U17620 (N_17620,N_16754,N_17116);
nand U17621 (N_17621,N_16889,N_16903);
nand U17622 (N_17622,N_17157,N_16927);
nand U17623 (N_17623,N_17031,N_17246);
and U17624 (N_17624,N_17464,N_17467);
xnor U17625 (N_17625,N_16446,N_16311);
xor U17626 (N_17626,N_16346,N_17304);
nor U17627 (N_17627,N_17229,N_17206);
xor U17628 (N_17628,N_16842,N_16761);
xnor U17629 (N_17629,N_17485,N_16466);
or U17630 (N_17630,N_16994,N_17168);
xor U17631 (N_17631,N_17451,N_17096);
and U17632 (N_17632,N_16546,N_16717);
and U17633 (N_17633,N_17118,N_16356);
xor U17634 (N_17634,N_16450,N_17404);
nand U17635 (N_17635,N_16482,N_16542);
xor U17636 (N_17636,N_16791,N_17029);
nand U17637 (N_17637,N_16436,N_17223);
and U17638 (N_17638,N_16916,N_17150);
and U17639 (N_17639,N_16698,N_17439);
or U17640 (N_17640,N_16424,N_16692);
xor U17641 (N_17641,N_16812,N_16519);
nor U17642 (N_17642,N_16343,N_16779);
nand U17643 (N_17643,N_17456,N_17227);
nand U17644 (N_17644,N_17459,N_17414);
and U17645 (N_17645,N_17138,N_17444);
xnor U17646 (N_17646,N_16406,N_17366);
nor U17647 (N_17647,N_16339,N_16262);
xnor U17648 (N_17648,N_17062,N_16308);
nor U17649 (N_17649,N_17016,N_17221);
nand U17650 (N_17650,N_16738,N_16663);
or U17651 (N_17651,N_16852,N_16497);
and U17652 (N_17652,N_16404,N_17329);
and U17653 (N_17653,N_16635,N_16714);
nor U17654 (N_17654,N_16597,N_17292);
or U17655 (N_17655,N_17027,N_16397);
or U17656 (N_17656,N_17358,N_16841);
and U17657 (N_17657,N_17045,N_17443);
nand U17658 (N_17658,N_16280,N_16765);
nand U17659 (N_17659,N_16475,N_16378);
nor U17660 (N_17660,N_17135,N_16372);
nor U17661 (N_17661,N_17114,N_17303);
and U17662 (N_17662,N_16766,N_16933);
nor U17663 (N_17663,N_16677,N_16547);
nand U17664 (N_17664,N_17146,N_16946);
or U17665 (N_17665,N_16434,N_17204);
nor U17666 (N_17666,N_16734,N_16797);
or U17667 (N_17667,N_16521,N_16594);
nand U17668 (N_17668,N_16586,N_16788);
and U17669 (N_17669,N_16831,N_16921);
or U17670 (N_17670,N_17236,N_16370);
and U17671 (N_17671,N_17394,N_16900);
or U17672 (N_17672,N_17429,N_17402);
or U17673 (N_17673,N_16266,N_17418);
and U17674 (N_17674,N_17038,N_17480);
or U17675 (N_17675,N_16669,N_17353);
xor U17676 (N_17676,N_16608,N_17013);
nor U17677 (N_17677,N_16525,N_16918);
nand U17678 (N_17678,N_16288,N_16580);
and U17679 (N_17679,N_16548,N_16999);
and U17680 (N_17680,N_16759,N_17237);
nor U17681 (N_17681,N_17491,N_16823);
nor U17682 (N_17682,N_17022,N_16671);
nand U17683 (N_17683,N_17203,N_16682);
and U17684 (N_17684,N_17173,N_16440);
nand U17685 (N_17685,N_17251,N_16570);
xnor U17686 (N_17686,N_17448,N_16750);
nand U17687 (N_17687,N_17427,N_16592);
or U17688 (N_17688,N_17256,N_17019);
nand U17689 (N_17689,N_16950,N_17211);
and U17690 (N_17690,N_16537,N_16958);
xnor U17691 (N_17691,N_16702,N_17291);
nor U17692 (N_17692,N_16272,N_16951);
and U17693 (N_17693,N_16382,N_16904);
nand U17694 (N_17694,N_17333,N_16509);
or U17695 (N_17695,N_17487,N_16449);
nand U17696 (N_17696,N_17222,N_17496);
nand U17697 (N_17697,N_17044,N_17159);
xnor U17698 (N_17698,N_16584,N_16768);
and U17699 (N_17699,N_16643,N_17162);
or U17700 (N_17700,N_17126,N_16680);
nor U17701 (N_17701,N_16938,N_16964);
xor U17702 (N_17702,N_17198,N_17341);
nand U17703 (N_17703,N_16840,N_16676);
nand U17704 (N_17704,N_16460,N_17263);
xnor U17705 (N_17705,N_17275,N_16695);
and U17706 (N_17706,N_17243,N_16967);
xor U17707 (N_17707,N_16706,N_16295);
nand U17708 (N_17708,N_16395,N_16470);
nand U17709 (N_17709,N_16796,N_16683);
xor U17710 (N_17710,N_16777,N_16998);
xor U17711 (N_17711,N_16389,N_17170);
xor U17712 (N_17712,N_16741,N_17294);
or U17713 (N_17713,N_17355,N_16691);
xor U17714 (N_17714,N_16983,N_16658);
nand U17715 (N_17715,N_16793,N_17490);
nor U17716 (N_17716,N_16960,N_17030);
or U17717 (N_17717,N_16917,N_17239);
or U17718 (N_17718,N_17437,N_17339);
and U17719 (N_17719,N_16336,N_17010);
xnor U17720 (N_17720,N_17405,N_17270);
and U17721 (N_17721,N_17099,N_16730);
xnor U17722 (N_17722,N_16405,N_17469);
nor U17723 (N_17723,N_16379,N_16882);
xor U17724 (N_17724,N_16416,N_17155);
xnor U17725 (N_17725,N_16952,N_16618);
or U17726 (N_17726,N_17080,N_17193);
nor U17727 (N_17727,N_17205,N_17196);
xor U17728 (N_17728,N_16417,N_16528);
or U17729 (N_17729,N_16422,N_17321);
xor U17730 (N_17730,N_16495,N_17040);
and U17731 (N_17731,N_16310,N_17363);
or U17732 (N_17732,N_17200,N_16773);
and U17733 (N_17733,N_16569,N_16915);
or U17734 (N_17734,N_17435,N_17131);
nand U17735 (N_17735,N_16323,N_16965);
xor U17736 (N_17736,N_17273,N_16720);
nand U17737 (N_17737,N_17072,N_16923);
nor U17738 (N_17738,N_16846,N_16265);
nand U17739 (N_17739,N_17287,N_16612);
and U17740 (N_17740,N_16552,N_17348);
nor U17741 (N_17741,N_17086,N_16955);
nand U17742 (N_17742,N_17091,N_17475);
nand U17743 (N_17743,N_16376,N_16333);
nand U17744 (N_17744,N_16772,N_17497);
xor U17745 (N_17745,N_16794,N_16814);
nand U17746 (N_17746,N_16253,N_16786);
xnor U17747 (N_17747,N_16884,N_16342);
xor U17748 (N_17748,N_17075,N_17201);
and U17749 (N_17749,N_16309,N_16898);
or U17750 (N_17750,N_17334,N_16710);
and U17751 (N_17751,N_16939,N_17492);
nand U17752 (N_17752,N_17488,N_16575);
nand U17753 (N_17753,N_17486,N_17218);
or U17754 (N_17754,N_17115,N_16957);
nor U17755 (N_17755,N_17407,N_16636);
and U17756 (N_17756,N_16578,N_17281);
nand U17757 (N_17757,N_17154,N_17254);
and U17758 (N_17758,N_17087,N_16709);
xnor U17759 (N_17759,N_16410,N_16486);
xnor U17760 (N_17760,N_16666,N_17186);
or U17761 (N_17761,N_17395,N_17242);
nor U17762 (N_17762,N_16473,N_17093);
nor U17763 (N_17763,N_17002,N_17174);
or U17764 (N_17764,N_17060,N_16775);
or U17765 (N_17765,N_17350,N_16438);
or U17766 (N_17766,N_17185,N_17177);
xor U17767 (N_17767,N_16276,N_16752);
xnor U17768 (N_17768,N_17101,N_17365);
nand U17769 (N_17769,N_17313,N_16538);
or U17770 (N_17770,N_16968,N_16590);
nand U17771 (N_17771,N_16326,N_16606);
nand U17772 (N_17772,N_16297,N_17233);
xor U17773 (N_17773,N_17058,N_16862);
or U17774 (N_17774,N_16984,N_17160);
xor U17775 (N_17775,N_17018,N_16711);
nor U17776 (N_17776,N_16920,N_16325);
xnor U17777 (N_17777,N_16479,N_17311);
or U17778 (N_17778,N_16543,N_16615);
and U17779 (N_17779,N_16801,N_17409);
nor U17780 (N_17780,N_17129,N_16769);
or U17781 (N_17781,N_16985,N_16631);
and U17782 (N_17782,N_16854,N_16421);
nand U17783 (N_17783,N_16411,N_16251);
and U17784 (N_17784,N_16755,N_16361);
and U17785 (N_17785,N_16970,N_16894);
or U17786 (N_17786,N_16273,N_17285);
nand U17787 (N_17787,N_16398,N_16380);
nand U17788 (N_17788,N_17017,N_16319);
and U17789 (N_17789,N_17455,N_16439);
and U17790 (N_17790,N_17410,N_17465);
and U17791 (N_17791,N_16526,N_16514);
xor U17792 (N_17792,N_17226,N_16474);
or U17793 (N_17793,N_17310,N_17458);
nor U17794 (N_17794,N_16275,N_16559);
nor U17795 (N_17795,N_16760,N_17009);
nor U17796 (N_17796,N_16879,N_17025);
xor U17797 (N_17797,N_16576,N_17235);
and U17798 (N_17798,N_17388,N_16252);
and U17799 (N_17799,N_16665,N_17295);
nor U17800 (N_17800,N_17463,N_17006);
or U17801 (N_17801,N_16423,N_17493);
xnor U17802 (N_17802,N_16799,N_16829);
nand U17803 (N_17803,N_16599,N_16358);
nor U17804 (N_17804,N_16719,N_17104);
and U17805 (N_17805,N_17308,N_16536);
or U17806 (N_17806,N_17166,N_16969);
or U17807 (N_17807,N_17092,N_16662);
nand U17808 (N_17808,N_16499,N_16802);
nor U17809 (N_17809,N_16393,N_16981);
nand U17810 (N_17810,N_16991,N_16651);
and U17811 (N_17811,N_16886,N_17271);
xor U17812 (N_17812,N_17332,N_17349);
nand U17813 (N_17813,N_17357,N_16591);
nor U17814 (N_17814,N_17181,N_17387);
xor U17815 (N_17815,N_17098,N_16974);
or U17816 (N_17816,N_16451,N_16385);
or U17817 (N_17817,N_16749,N_16906);
nand U17818 (N_17818,N_16770,N_17207);
and U17819 (N_17819,N_17440,N_16430);
or U17820 (N_17820,N_17037,N_16688);
xor U17821 (N_17821,N_17004,N_17151);
or U17822 (N_17822,N_17191,N_16407);
xor U17823 (N_17823,N_17397,N_17472);
nand U17824 (N_17824,N_16285,N_16391);
nor U17825 (N_17825,N_16571,N_17176);
and U17826 (N_17826,N_16568,N_17054);
nand U17827 (N_17827,N_16522,N_16744);
nor U17828 (N_17828,N_16805,N_16255);
nor U17829 (N_17829,N_16743,N_16650);
and U17830 (N_17830,N_16827,N_16627);
nor U17831 (N_17831,N_17036,N_16327);
nand U17832 (N_17832,N_17130,N_16490);
and U17833 (N_17833,N_16312,N_16541);
xnor U17834 (N_17834,N_17453,N_16640);
nand U17835 (N_17835,N_16896,N_16881);
xor U17836 (N_17836,N_16532,N_16634);
xor U17837 (N_17837,N_16269,N_16800);
xnor U17838 (N_17838,N_16481,N_16787);
xor U17839 (N_17839,N_16649,N_16992);
or U17840 (N_17840,N_16456,N_16485);
nor U17841 (N_17841,N_16892,N_16294);
nor U17842 (N_17842,N_17183,N_17232);
and U17843 (N_17843,N_16956,N_16573);
nand U17844 (N_17844,N_16943,N_16270);
nand U17845 (N_17845,N_16563,N_17172);
nand U17846 (N_17846,N_16632,N_16712);
nor U17847 (N_17847,N_17390,N_16767);
nand U17848 (N_17848,N_17147,N_16513);
and U17849 (N_17849,N_16619,N_16982);
xor U17850 (N_17850,N_17095,N_17158);
or U17851 (N_17851,N_17033,N_16554);
and U17852 (N_17852,N_16780,N_16304);
nor U17853 (N_17853,N_16963,N_16748);
nor U17854 (N_17854,N_16447,N_17372);
or U17855 (N_17855,N_17354,N_16834);
and U17856 (N_17856,N_16871,N_16891);
and U17857 (N_17857,N_16505,N_16753);
nand U17858 (N_17858,N_16989,N_16789);
nor U17859 (N_17859,N_16652,N_16966);
or U17860 (N_17860,N_17257,N_16721);
nand U17861 (N_17861,N_16693,N_16925);
or U17862 (N_17862,N_17462,N_16910);
and U17863 (N_17863,N_16444,N_16736);
nand U17864 (N_17864,N_16282,N_16353);
xnor U17865 (N_17865,N_16687,N_16828);
xor U17866 (N_17866,N_17343,N_16972);
or U17867 (N_17867,N_17077,N_17247);
nor U17868 (N_17868,N_16907,N_17260);
and U17869 (N_17869,N_16567,N_17132);
and U17870 (N_17870,N_17188,N_16785);
and U17871 (N_17871,N_17415,N_16757);
nor U17872 (N_17872,N_16291,N_16959);
or U17873 (N_17873,N_16851,N_16784);
nor U17874 (N_17874,N_16945,N_16716);
nand U17875 (N_17875,N_17244,N_16815);
nand U17876 (N_17876,N_16674,N_16811);
nor U17877 (N_17877,N_17391,N_16661);
and U17878 (N_17878,N_17268,N_16419);
nor U17879 (N_17879,N_17074,N_16374);
or U17880 (N_17880,N_17171,N_17128);
nand U17881 (N_17881,N_16489,N_16724);
and U17882 (N_17882,N_17406,N_16335);
or U17883 (N_17883,N_17069,N_17148);
nand U17884 (N_17884,N_16625,N_16301);
xor U17885 (N_17885,N_16629,N_16700);
nand U17886 (N_17886,N_16646,N_16545);
or U17887 (N_17887,N_16947,N_16641);
and U17888 (N_17888,N_16427,N_16699);
and U17889 (N_17889,N_17327,N_16403);
and U17890 (N_17890,N_16445,N_16515);
and U17891 (N_17891,N_16742,N_16993);
nand U17892 (N_17892,N_16733,N_16428);
nor U17893 (N_17893,N_16279,N_16885);
and U17894 (N_17894,N_17124,N_16402);
or U17895 (N_17895,N_16732,N_16924);
or U17896 (N_17896,N_17428,N_16860);
or U17897 (N_17897,N_16307,N_17248);
nand U17898 (N_17898,N_16868,N_16807);
nand U17899 (N_17899,N_16941,N_16324);
nor U17900 (N_17900,N_16283,N_17085);
nand U17901 (N_17901,N_16901,N_17245);
and U17902 (N_17902,N_16836,N_16867);
or U17903 (N_17903,N_16715,N_17269);
xnor U17904 (N_17904,N_17061,N_16830);
nor U17905 (N_17905,N_16648,N_16620);
or U17906 (N_17906,N_16413,N_17434);
or U17907 (N_17907,N_16292,N_17449);
or U17908 (N_17908,N_16534,N_16564);
nand U17909 (N_17909,N_16942,N_17234);
nor U17910 (N_17910,N_16281,N_16332);
nor U17911 (N_17911,N_17259,N_17323);
and U17912 (N_17912,N_17319,N_16655);
nand U17913 (N_17913,N_16461,N_16588);
xnor U17914 (N_17914,N_16360,N_16574);
and U17915 (N_17915,N_17078,N_16298);
nor U17916 (N_17916,N_16675,N_17468);
nand U17917 (N_17917,N_16696,N_17403);
and U17918 (N_17918,N_16888,N_17345);
nand U17919 (N_17919,N_16988,N_16401);
nand U17920 (N_17920,N_17117,N_17314);
xor U17921 (N_17921,N_17279,N_16913);
or U17922 (N_17922,N_16350,N_17142);
and U17923 (N_17923,N_16607,N_16809);
and U17924 (N_17924,N_16795,N_16337);
nand U17925 (N_17925,N_17231,N_17384);
or U17926 (N_17926,N_17301,N_17143);
xor U17927 (N_17927,N_17043,N_16464);
nand U17928 (N_17928,N_17436,N_17368);
nand U17929 (N_17929,N_16409,N_17379);
and U17930 (N_17930,N_16510,N_16883);
xor U17931 (N_17931,N_16609,N_17315);
or U17932 (N_17932,N_16377,N_17446);
or U17933 (N_17933,N_17431,N_16420);
or U17934 (N_17934,N_16853,N_16837);
nand U17935 (N_17935,N_17380,N_16816);
or U17936 (N_17936,N_16581,N_16425);
nor U17937 (N_17937,N_16454,N_16390);
nand U17938 (N_17938,N_17152,N_16507);
and U17939 (N_17939,N_16605,N_17416);
or U17940 (N_17940,N_17298,N_17307);
or U17941 (N_17941,N_16394,N_17495);
nor U17942 (N_17942,N_17103,N_17277);
and U17943 (N_17943,N_17209,N_17378);
xnor U17944 (N_17944,N_16990,N_16987);
and U17945 (N_17945,N_17318,N_16287);
xor U17946 (N_17946,N_17325,N_16705);
nand U17947 (N_17947,N_16518,N_17389);
or U17948 (N_17948,N_16271,N_16352);
or U17949 (N_17949,N_17050,N_16911);
nor U17950 (N_17950,N_17169,N_17007);
xnor U17951 (N_17951,N_17335,N_17309);
and U17952 (N_17952,N_16654,N_16316);
nor U17953 (N_17953,N_16873,N_16399);
nand U17954 (N_17954,N_16935,N_17213);
and U17955 (N_17955,N_16535,N_16364);
xor U17956 (N_17956,N_16670,N_16745);
nor U17957 (N_17957,N_16603,N_16465);
nor U17958 (N_17958,N_16322,N_16448);
or U17959 (N_17959,N_17014,N_16344);
xnor U17960 (N_17960,N_16928,N_16418);
or U17961 (N_17961,N_16937,N_17250);
xnor U17962 (N_17962,N_17430,N_16341);
and U17963 (N_17963,N_16367,N_16926);
or U17964 (N_17964,N_16763,N_16686);
and U17965 (N_17965,N_17153,N_16708);
nor U17966 (N_17966,N_16516,N_17441);
or U17967 (N_17967,N_17362,N_16306);
and U17968 (N_17968,N_16704,N_17413);
nand U17969 (N_17969,N_17108,N_16808);
or U17970 (N_17970,N_17471,N_17412);
nand U17971 (N_17971,N_16317,N_16645);
or U17972 (N_17972,N_16857,N_16462);
nand U17973 (N_17973,N_16684,N_17276);
nand U17974 (N_17974,N_17120,N_16305);
nand U17975 (N_17975,N_17097,N_16289);
or U17976 (N_17976,N_16469,N_16813);
and U17977 (N_17977,N_17220,N_17076);
and U17978 (N_17978,N_17032,N_17094);
nor U17979 (N_17979,N_16539,N_16751);
xor U17980 (N_17980,N_16561,N_16914);
xor U17981 (N_17981,N_16261,N_16756);
or U17982 (N_17982,N_16601,N_17336);
nor U17983 (N_17983,N_16560,N_17442);
nor U17984 (N_17984,N_17052,N_16455);
nand U17985 (N_17985,N_16980,N_17042);
or U17986 (N_17986,N_17208,N_16369);
and U17987 (N_17987,N_17064,N_16723);
nor U17988 (N_17988,N_17421,N_17342);
or U17989 (N_17989,N_16728,N_17113);
or U17990 (N_17990,N_16562,N_16978);
xor U17991 (N_17991,N_17288,N_16694);
and U17992 (N_17992,N_17338,N_17356);
xnor U17993 (N_17993,N_17324,N_16817);
nor U17994 (N_17994,N_16897,N_16727);
xor U17995 (N_17995,N_17423,N_16583);
nor U17996 (N_17996,N_17161,N_16340);
xnor U17997 (N_17997,N_17450,N_17070);
and U17998 (N_17998,N_16713,N_16673);
xor U17999 (N_17999,N_17156,N_17088);
or U18000 (N_18000,N_17473,N_16731);
nand U18001 (N_18001,N_16511,N_17386);
nand U18002 (N_18002,N_17175,N_17192);
and U18003 (N_18003,N_17140,N_16762);
nor U18004 (N_18004,N_16856,N_16820);
nor U18005 (N_18005,N_16375,N_16579);
and U18006 (N_18006,N_16825,N_16523);
xnor U18007 (N_18007,N_17477,N_17179);
or U18008 (N_18008,N_16426,N_16286);
or U18009 (N_18009,N_17393,N_16318);
nor U18010 (N_18010,N_17401,N_17005);
xnor U18011 (N_18011,N_17015,N_16656);
and U18012 (N_18012,N_16263,N_16869);
and U18013 (N_18013,N_17195,N_17306);
nand U18014 (N_18014,N_17417,N_16557);
and U18015 (N_18015,N_16334,N_16975);
nand U18016 (N_18016,N_17053,N_16783);
and U18017 (N_18017,N_17012,N_16302);
nor U18018 (N_18018,N_16315,N_16387);
nand U18019 (N_18019,N_17305,N_17364);
nor U18020 (N_18020,N_16961,N_16624);
and U18021 (N_18021,N_16566,N_16833);
nand U18022 (N_18022,N_17125,N_16774);
xnor U18023 (N_18023,N_16726,N_16256);
nor U18024 (N_18024,N_17297,N_16290);
nor U18025 (N_18025,N_17280,N_17252);
nand U18026 (N_18026,N_16610,N_17498);
xnor U18027 (N_18027,N_17210,N_17144);
or U18028 (N_18028,N_16506,N_16806);
or U18029 (N_18029,N_17024,N_16740);
nand U18030 (N_18030,N_16517,N_16363);
nand U18031 (N_18031,N_17296,N_16296);
and U18032 (N_18032,N_16977,N_17184);
nand U18033 (N_18033,N_17089,N_17278);
xor U18034 (N_18034,N_17461,N_16623);
xor U18035 (N_18035,N_17164,N_17090);
nor U18036 (N_18036,N_17100,N_17478);
and U18037 (N_18037,N_16258,N_16866);
or U18038 (N_18038,N_16467,N_16496);
nand U18039 (N_18039,N_17255,N_16314);
nand U18040 (N_18040,N_17136,N_16512);
and U18041 (N_18041,N_16657,N_17241);
xnor U18042 (N_18042,N_17481,N_16501);
xnor U18043 (N_18043,N_16979,N_16908);
and U18044 (N_18044,N_17408,N_16328);
nor U18045 (N_18045,N_17340,N_17084);
or U18046 (N_18046,N_17083,N_16986);
or U18047 (N_18047,N_17422,N_16371);
nor U18048 (N_18048,N_16392,N_16284);
nand U18049 (N_18049,N_17432,N_16488);
or U18050 (N_18050,N_16737,N_16593);
or U18051 (N_18051,N_17474,N_17021);
nor U18052 (N_18052,N_17330,N_16667);
nor U18053 (N_18053,N_16735,N_16764);
nand U18054 (N_18054,N_17489,N_17046);
nand U18055 (N_18055,N_17079,N_17302);
xor U18056 (N_18056,N_17165,N_17178);
nor U18057 (N_18057,N_16890,N_16628);
or U18058 (N_18058,N_16832,N_16859);
xnor U18059 (N_18059,N_17392,N_17262);
and U18060 (N_18060,N_17145,N_17445);
and U18061 (N_18061,N_16476,N_16259);
nand U18062 (N_18062,N_16368,N_16949);
or U18063 (N_18063,N_16758,N_17346);
nand U18064 (N_18064,N_17312,N_17202);
and U18065 (N_18065,N_17359,N_17071);
xnor U18066 (N_18066,N_16776,N_16948);
nand U18067 (N_18067,N_16600,N_16429);
nor U18068 (N_18068,N_16973,N_16902);
and U18069 (N_18069,N_16582,N_16257);
nand U18070 (N_18070,N_16452,N_16678);
and U18071 (N_18071,N_17068,N_17127);
or U18072 (N_18072,N_17337,N_16644);
and U18073 (N_18073,N_16491,N_16664);
nor U18074 (N_18074,N_16647,N_16878);
and U18075 (N_18075,N_16386,N_16585);
nor U18076 (N_18076,N_16895,N_16996);
or U18077 (N_18077,N_16359,N_16381);
nor U18078 (N_18078,N_17361,N_16821);
nor U18079 (N_18079,N_16932,N_17107);
nor U18080 (N_18080,N_16508,N_16453);
nor U18081 (N_18081,N_16861,N_17266);
nand U18082 (N_18082,N_16782,N_16971);
or U18083 (N_18083,N_16553,N_16995);
xor U18084 (N_18084,N_17317,N_17316);
nand U18085 (N_18085,N_16396,N_16690);
xor U18086 (N_18086,N_16865,N_17264);
nor U18087 (N_18087,N_16550,N_17212);
nand U18088 (N_18088,N_16443,N_16887);
and U18089 (N_18089,N_16530,N_16790);
and U18090 (N_18090,N_16679,N_17039);
or U18091 (N_18091,N_17284,N_16437);
nor U18092 (N_18092,N_16373,N_17063);
nand U18093 (N_18093,N_16637,N_16929);
and U18094 (N_18094,N_16331,N_16912);
nand U18095 (N_18095,N_17123,N_17460);
nor U18096 (N_18096,N_16459,N_16613);
and U18097 (N_18097,N_17385,N_16551);
and U18098 (N_18098,N_16844,N_17371);
nor U18099 (N_18099,N_16498,N_16781);
and U18100 (N_18100,N_16626,N_17320);
xnor U18101 (N_18101,N_16483,N_16321);
nor U18102 (N_18102,N_17057,N_16408);
nand U18103 (N_18103,N_16899,N_17373);
nand U18104 (N_18104,N_16338,N_17149);
xor U18105 (N_18105,N_17238,N_17217);
nor U18106 (N_18106,N_17020,N_16384);
and U18107 (N_18107,N_16819,N_16746);
xor U18108 (N_18108,N_17049,N_16480);
and U18109 (N_18109,N_16962,N_17351);
nor U18110 (N_18110,N_16660,N_17396);
or U18111 (N_18111,N_17382,N_17228);
or U18112 (N_18112,N_17375,N_17420);
nand U18113 (N_18113,N_16587,N_16611);
nor U18114 (N_18114,N_16621,N_17023);
and U18115 (N_18115,N_17056,N_17272);
nor U18116 (N_18116,N_16848,N_16349);
xor U18117 (N_18117,N_16487,N_17466);
or U18118 (N_18118,N_16875,N_16672);
or U18119 (N_18119,N_17230,N_16362);
and U18120 (N_18120,N_17300,N_16260);
nand U18121 (N_18121,N_16589,N_16804);
xnor U18122 (N_18122,N_16431,N_16893);
nor U18123 (N_18123,N_16345,N_16729);
nand U18124 (N_18124,N_16268,N_16778);
nor U18125 (N_18125,N_17339,N_17480);
or U18126 (N_18126,N_16812,N_16681);
nor U18127 (N_18127,N_16295,N_16883);
nand U18128 (N_18128,N_16600,N_17234);
nand U18129 (N_18129,N_16260,N_16618);
nand U18130 (N_18130,N_17209,N_17310);
nor U18131 (N_18131,N_17206,N_16979);
nor U18132 (N_18132,N_16982,N_16374);
nand U18133 (N_18133,N_16264,N_16552);
or U18134 (N_18134,N_17377,N_17254);
and U18135 (N_18135,N_17294,N_16614);
nor U18136 (N_18136,N_17046,N_16349);
and U18137 (N_18137,N_17059,N_16519);
or U18138 (N_18138,N_17430,N_17057);
and U18139 (N_18139,N_16392,N_16527);
or U18140 (N_18140,N_16636,N_17087);
or U18141 (N_18141,N_16511,N_16950);
nor U18142 (N_18142,N_16487,N_16548);
nor U18143 (N_18143,N_17221,N_16725);
or U18144 (N_18144,N_16568,N_16628);
xnor U18145 (N_18145,N_16389,N_17304);
or U18146 (N_18146,N_17468,N_16906);
xnor U18147 (N_18147,N_16296,N_16644);
nand U18148 (N_18148,N_16576,N_17294);
nand U18149 (N_18149,N_16885,N_16980);
nand U18150 (N_18150,N_16488,N_16890);
xnor U18151 (N_18151,N_17286,N_17045);
xnor U18152 (N_18152,N_16485,N_17139);
or U18153 (N_18153,N_17250,N_17377);
and U18154 (N_18154,N_16820,N_16763);
nand U18155 (N_18155,N_16504,N_16414);
or U18156 (N_18156,N_17286,N_16659);
xor U18157 (N_18157,N_17052,N_16732);
nor U18158 (N_18158,N_17364,N_16773);
xor U18159 (N_18159,N_16764,N_16539);
or U18160 (N_18160,N_16451,N_16804);
and U18161 (N_18161,N_17179,N_17497);
xnor U18162 (N_18162,N_17343,N_16913);
xnor U18163 (N_18163,N_17204,N_16828);
and U18164 (N_18164,N_16590,N_16454);
nand U18165 (N_18165,N_16320,N_16910);
xor U18166 (N_18166,N_16824,N_16599);
nor U18167 (N_18167,N_17212,N_16909);
and U18168 (N_18168,N_17095,N_17309);
nor U18169 (N_18169,N_17013,N_17443);
or U18170 (N_18170,N_16746,N_16571);
nor U18171 (N_18171,N_16789,N_17487);
or U18172 (N_18172,N_17458,N_16615);
and U18173 (N_18173,N_16852,N_16722);
and U18174 (N_18174,N_16987,N_17180);
nand U18175 (N_18175,N_16717,N_16813);
and U18176 (N_18176,N_17134,N_16659);
or U18177 (N_18177,N_17011,N_17037);
and U18178 (N_18178,N_17240,N_16509);
xnor U18179 (N_18179,N_16307,N_17384);
or U18180 (N_18180,N_17405,N_17065);
xor U18181 (N_18181,N_17136,N_16893);
nor U18182 (N_18182,N_17376,N_17473);
or U18183 (N_18183,N_17227,N_16925);
nor U18184 (N_18184,N_17374,N_17243);
and U18185 (N_18185,N_17435,N_17026);
or U18186 (N_18186,N_17461,N_16274);
and U18187 (N_18187,N_16840,N_16687);
nor U18188 (N_18188,N_17314,N_17210);
and U18189 (N_18189,N_16322,N_16726);
or U18190 (N_18190,N_16892,N_16517);
xor U18191 (N_18191,N_17460,N_17445);
nor U18192 (N_18192,N_16359,N_17247);
nand U18193 (N_18193,N_16312,N_17205);
and U18194 (N_18194,N_16379,N_16573);
xnor U18195 (N_18195,N_17488,N_16642);
nand U18196 (N_18196,N_16805,N_16948);
or U18197 (N_18197,N_16760,N_16412);
nor U18198 (N_18198,N_17430,N_16364);
xor U18199 (N_18199,N_17226,N_16564);
and U18200 (N_18200,N_16304,N_17291);
or U18201 (N_18201,N_16332,N_17208);
nand U18202 (N_18202,N_17141,N_16411);
or U18203 (N_18203,N_17469,N_16611);
nand U18204 (N_18204,N_17449,N_16772);
xnor U18205 (N_18205,N_17387,N_17477);
xnor U18206 (N_18206,N_17403,N_16269);
nand U18207 (N_18207,N_16738,N_17194);
xnor U18208 (N_18208,N_17123,N_16273);
or U18209 (N_18209,N_17092,N_16651);
nand U18210 (N_18210,N_17094,N_16973);
or U18211 (N_18211,N_17216,N_16543);
nor U18212 (N_18212,N_16893,N_17475);
xnor U18213 (N_18213,N_16996,N_17258);
nand U18214 (N_18214,N_16704,N_17484);
nor U18215 (N_18215,N_16947,N_16256);
nand U18216 (N_18216,N_17005,N_16371);
xnor U18217 (N_18217,N_16957,N_16628);
nor U18218 (N_18218,N_16567,N_16907);
or U18219 (N_18219,N_16311,N_16350);
nand U18220 (N_18220,N_16790,N_16735);
xor U18221 (N_18221,N_16350,N_16556);
nor U18222 (N_18222,N_16961,N_16448);
and U18223 (N_18223,N_16528,N_17399);
nor U18224 (N_18224,N_16998,N_17266);
nor U18225 (N_18225,N_17068,N_17293);
or U18226 (N_18226,N_17135,N_17202);
or U18227 (N_18227,N_17222,N_16365);
nand U18228 (N_18228,N_16785,N_16935);
or U18229 (N_18229,N_16576,N_16266);
nand U18230 (N_18230,N_17059,N_16379);
and U18231 (N_18231,N_16997,N_16485);
nor U18232 (N_18232,N_16481,N_16676);
or U18233 (N_18233,N_16832,N_17130);
and U18234 (N_18234,N_16827,N_17182);
or U18235 (N_18235,N_16691,N_17497);
nor U18236 (N_18236,N_16565,N_16804);
nor U18237 (N_18237,N_16291,N_16566);
xor U18238 (N_18238,N_16633,N_16640);
nor U18239 (N_18239,N_16636,N_17143);
or U18240 (N_18240,N_16823,N_17381);
xnor U18241 (N_18241,N_16888,N_17253);
nor U18242 (N_18242,N_16855,N_16719);
and U18243 (N_18243,N_17115,N_17037);
xnor U18244 (N_18244,N_17215,N_17263);
or U18245 (N_18245,N_17353,N_16894);
nor U18246 (N_18246,N_16513,N_17302);
or U18247 (N_18247,N_17266,N_16854);
nand U18248 (N_18248,N_16821,N_16373);
and U18249 (N_18249,N_17055,N_17395);
nand U18250 (N_18250,N_17233,N_16960);
nor U18251 (N_18251,N_16799,N_17193);
xor U18252 (N_18252,N_17190,N_17200);
and U18253 (N_18253,N_16504,N_17174);
nor U18254 (N_18254,N_16686,N_17291);
nor U18255 (N_18255,N_16768,N_17297);
nor U18256 (N_18256,N_16743,N_16696);
nand U18257 (N_18257,N_17009,N_16973);
xor U18258 (N_18258,N_17161,N_17316);
and U18259 (N_18259,N_16712,N_16662);
nand U18260 (N_18260,N_16400,N_17231);
nand U18261 (N_18261,N_16702,N_17329);
nand U18262 (N_18262,N_16323,N_16581);
and U18263 (N_18263,N_17005,N_16819);
xnor U18264 (N_18264,N_16927,N_16761);
nor U18265 (N_18265,N_17114,N_16954);
nor U18266 (N_18266,N_17348,N_16850);
or U18267 (N_18267,N_16387,N_16648);
xor U18268 (N_18268,N_17421,N_17407);
and U18269 (N_18269,N_17480,N_17217);
nor U18270 (N_18270,N_16459,N_16454);
nor U18271 (N_18271,N_17144,N_17493);
or U18272 (N_18272,N_16570,N_16909);
nand U18273 (N_18273,N_16299,N_16845);
nand U18274 (N_18274,N_16738,N_17299);
or U18275 (N_18275,N_17190,N_16983);
xnor U18276 (N_18276,N_17372,N_17159);
nor U18277 (N_18277,N_17164,N_16744);
nand U18278 (N_18278,N_17356,N_16303);
nand U18279 (N_18279,N_16276,N_16961);
or U18280 (N_18280,N_17440,N_17362);
or U18281 (N_18281,N_17295,N_16885);
and U18282 (N_18282,N_16274,N_17065);
nand U18283 (N_18283,N_16754,N_16544);
or U18284 (N_18284,N_17336,N_16326);
nor U18285 (N_18285,N_17178,N_16851);
nand U18286 (N_18286,N_16632,N_17002);
xor U18287 (N_18287,N_17401,N_16740);
xnor U18288 (N_18288,N_17159,N_17469);
nand U18289 (N_18289,N_17092,N_16253);
nand U18290 (N_18290,N_16995,N_17077);
nand U18291 (N_18291,N_16784,N_17399);
xor U18292 (N_18292,N_17349,N_16259);
nand U18293 (N_18293,N_16890,N_17105);
nand U18294 (N_18294,N_16787,N_16477);
nand U18295 (N_18295,N_16658,N_16432);
nand U18296 (N_18296,N_16934,N_16619);
and U18297 (N_18297,N_16283,N_16365);
xnor U18298 (N_18298,N_16881,N_16570);
and U18299 (N_18299,N_16654,N_17165);
nand U18300 (N_18300,N_16702,N_16369);
nand U18301 (N_18301,N_16451,N_17084);
xnor U18302 (N_18302,N_16718,N_16260);
nand U18303 (N_18303,N_16535,N_16284);
nor U18304 (N_18304,N_17471,N_16894);
nor U18305 (N_18305,N_16636,N_17132);
nor U18306 (N_18306,N_17392,N_16471);
or U18307 (N_18307,N_16371,N_16260);
nand U18308 (N_18308,N_17304,N_16440);
nor U18309 (N_18309,N_16570,N_16624);
xnor U18310 (N_18310,N_16975,N_17340);
nand U18311 (N_18311,N_17114,N_17307);
or U18312 (N_18312,N_17169,N_16432);
xnor U18313 (N_18313,N_16821,N_16511);
and U18314 (N_18314,N_16370,N_16256);
and U18315 (N_18315,N_17334,N_16412);
xnor U18316 (N_18316,N_16634,N_16826);
nand U18317 (N_18317,N_16649,N_16605);
nor U18318 (N_18318,N_16690,N_17276);
or U18319 (N_18319,N_16431,N_16822);
xnor U18320 (N_18320,N_16719,N_17083);
or U18321 (N_18321,N_16526,N_16370);
or U18322 (N_18322,N_17089,N_16606);
or U18323 (N_18323,N_17034,N_16776);
nor U18324 (N_18324,N_16631,N_17474);
and U18325 (N_18325,N_16471,N_17205);
nor U18326 (N_18326,N_17062,N_16755);
nor U18327 (N_18327,N_17178,N_17434);
xnor U18328 (N_18328,N_16792,N_16826);
xor U18329 (N_18329,N_16938,N_17328);
or U18330 (N_18330,N_17325,N_16446);
and U18331 (N_18331,N_17205,N_16964);
and U18332 (N_18332,N_16290,N_16565);
xor U18333 (N_18333,N_17218,N_17018);
and U18334 (N_18334,N_16376,N_17106);
nor U18335 (N_18335,N_16255,N_16848);
xnor U18336 (N_18336,N_16299,N_16316);
or U18337 (N_18337,N_16439,N_16415);
xnor U18338 (N_18338,N_16846,N_17269);
nor U18339 (N_18339,N_16746,N_16818);
nor U18340 (N_18340,N_16332,N_17006);
nor U18341 (N_18341,N_17481,N_16583);
nor U18342 (N_18342,N_16601,N_16820);
or U18343 (N_18343,N_17428,N_17087);
nand U18344 (N_18344,N_16372,N_17321);
or U18345 (N_18345,N_16882,N_16862);
and U18346 (N_18346,N_17261,N_16496);
and U18347 (N_18347,N_17107,N_16344);
nand U18348 (N_18348,N_17368,N_16926);
nand U18349 (N_18349,N_17074,N_16713);
nor U18350 (N_18350,N_17477,N_16400);
nor U18351 (N_18351,N_16775,N_16511);
nand U18352 (N_18352,N_17478,N_16552);
nor U18353 (N_18353,N_16627,N_16974);
nor U18354 (N_18354,N_17051,N_17021);
or U18355 (N_18355,N_16891,N_17308);
and U18356 (N_18356,N_16733,N_16574);
or U18357 (N_18357,N_16311,N_17395);
xor U18358 (N_18358,N_16892,N_17068);
or U18359 (N_18359,N_16904,N_16575);
and U18360 (N_18360,N_16390,N_16459);
xor U18361 (N_18361,N_16281,N_17122);
xnor U18362 (N_18362,N_17133,N_16568);
nor U18363 (N_18363,N_16694,N_17320);
xor U18364 (N_18364,N_17028,N_16853);
nand U18365 (N_18365,N_16273,N_16483);
nor U18366 (N_18366,N_16796,N_16515);
and U18367 (N_18367,N_16829,N_16884);
xor U18368 (N_18368,N_16791,N_17448);
or U18369 (N_18369,N_17405,N_16958);
or U18370 (N_18370,N_16906,N_16831);
or U18371 (N_18371,N_16556,N_16817);
nand U18372 (N_18372,N_16947,N_17397);
nor U18373 (N_18373,N_16831,N_17163);
or U18374 (N_18374,N_16700,N_16890);
nor U18375 (N_18375,N_17497,N_17006);
or U18376 (N_18376,N_16899,N_16443);
or U18377 (N_18377,N_16451,N_16345);
and U18378 (N_18378,N_16557,N_17230);
nor U18379 (N_18379,N_16475,N_16417);
and U18380 (N_18380,N_16750,N_17092);
nand U18381 (N_18381,N_17177,N_16725);
and U18382 (N_18382,N_17253,N_17180);
and U18383 (N_18383,N_16304,N_17068);
or U18384 (N_18384,N_16902,N_16769);
xnor U18385 (N_18385,N_17237,N_17225);
nor U18386 (N_18386,N_16311,N_17476);
or U18387 (N_18387,N_16466,N_16952);
and U18388 (N_18388,N_16961,N_16685);
and U18389 (N_18389,N_16455,N_16548);
and U18390 (N_18390,N_16307,N_16797);
or U18391 (N_18391,N_16794,N_17124);
nand U18392 (N_18392,N_17009,N_16695);
or U18393 (N_18393,N_17353,N_16847);
nand U18394 (N_18394,N_17205,N_16628);
nor U18395 (N_18395,N_17058,N_17170);
xnor U18396 (N_18396,N_16557,N_17221);
or U18397 (N_18397,N_17320,N_17028);
nand U18398 (N_18398,N_16787,N_17013);
xnor U18399 (N_18399,N_17110,N_17311);
nor U18400 (N_18400,N_16581,N_16893);
xor U18401 (N_18401,N_16879,N_17091);
xnor U18402 (N_18402,N_16810,N_16688);
and U18403 (N_18403,N_17164,N_17392);
nor U18404 (N_18404,N_17130,N_16556);
nor U18405 (N_18405,N_16611,N_16255);
and U18406 (N_18406,N_17371,N_16647);
nor U18407 (N_18407,N_16627,N_16671);
and U18408 (N_18408,N_16449,N_17422);
nor U18409 (N_18409,N_16466,N_16971);
and U18410 (N_18410,N_16986,N_17209);
nand U18411 (N_18411,N_16269,N_17321);
xor U18412 (N_18412,N_17326,N_16653);
nand U18413 (N_18413,N_17333,N_17055);
and U18414 (N_18414,N_16423,N_17465);
xnor U18415 (N_18415,N_17447,N_16398);
and U18416 (N_18416,N_17042,N_16675);
and U18417 (N_18417,N_17260,N_17304);
or U18418 (N_18418,N_16833,N_17372);
nand U18419 (N_18419,N_16549,N_17456);
nand U18420 (N_18420,N_16914,N_16411);
nand U18421 (N_18421,N_16803,N_17283);
xnor U18422 (N_18422,N_16969,N_17228);
xor U18423 (N_18423,N_16986,N_17467);
nand U18424 (N_18424,N_16569,N_16897);
nand U18425 (N_18425,N_16661,N_17149);
xnor U18426 (N_18426,N_16673,N_17011);
xor U18427 (N_18427,N_17056,N_16592);
and U18428 (N_18428,N_16701,N_16962);
xnor U18429 (N_18429,N_16358,N_16408);
and U18430 (N_18430,N_17107,N_16451);
nor U18431 (N_18431,N_17359,N_16521);
and U18432 (N_18432,N_16482,N_16933);
nand U18433 (N_18433,N_16558,N_16859);
and U18434 (N_18434,N_16502,N_16256);
nor U18435 (N_18435,N_16509,N_16366);
nand U18436 (N_18436,N_16640,N_16848);
xnor U18437 (N_18437,N_16728,N_16522);
xor U18438 (N_18438,N_16652,N_16390);
nand U18439 (N_18439,N_17187,N_16631);
nand U18440 (N_18440,N_16928,N_16451);
nand U18441 (N_18441,N_16795,N_16735);
xor U18442 (N_18442,N_17158,N_17325);
xor U18443 (N_18443,N_16498,N_16268);
and U18444 (N_18444,N_17306,N_16341);
nor U18445 (N_18445,N_16410,N_16651);
or U18446 (N_18446,N_16842,N_17322);
or U18447 (N_18447,N_16633,N_17279);
or U18448 (N_18448,N_16373,N_16840);
xnor U18449 (N_18449,N_16399,N_17092);
nand U18450 (N_18450,N_17005,N_16350);
or U18451 (N_18451,N_16748,N_17021);
and U18452 (N_18452,N_17177,N_16880);
or U18453 (N_18453,N_16329,N_17079);
and U18454 (N_18454,N_16259,N_16780);
or U18455 (N_18455,N_16924,N_16939);
nor U18456 (N_18456,N_16978,N_17374);
nand U18457 (N_18457,N_16589,N_17374);
or U18458 (N_18458,N_16628,N_16844);
or U18459 (N_18459,N_17468,N_16697);
xor U18460 (N_18460,N_17476,N_16958);
xnor U18461 (N_18461,N_17489,N_16415);
nand U18462 (N_18462,N_17220,N_17336);
xnor U18463 (N_18463,N_17118,N_16299);
nand U18464 (N_18464,N_16860,N_17459);
nor U18465 (N_18465,N_17311,N_16269);
and U18466 (N_18466,N_17292,N_17249);
nor U18467 (N_18467,N_17149,N_16460);
nand U18468 (N_18468,N_17067,N_17237);
nand U18469 (N_18469,N_16545,N_17496);
nand U18470 (N_18470,N_16924,N_16694);
nor U18471 (N_18471,N_17034,N_16804);
nand U18472 (N_18472,N_17488,N_16783);
nor U18473 (N_18473,N_16436,N_16698);
or U18474 (N_18474,N_16596,N_17272);
and U18475 (N_18475,N_16499,N_16718);
nand U18476 (N_18476,N_16747,N_16263);
nand U18477 (N_18477,N_16532,N_16594);
or U18478 (N_18478,N_17191,N_17456);
nand U18479 (N_18479,N_17129,N_16680);
xnor U18480 (N_18480,N_17379,N_16794);
or U18481 (N_18481,N_16897,N_17098);
and U18482 (N_18482,N_16543,N_17177);
xnor U18483 (N_18483,N_16625,N_16806);
nand U18484 (N_18484,N_16905,N_16412);
and U18485 (N_18485,N_16767,N_17026);
and U18486 (N_18486,N_16825,N_17005);
nand U18487 (N_18487,N_17266,N_17005);
nor U18488 (N_18488,N_16467,N_16850);
or U18489 (N_18489,N_17019,N_17044);
and U18490 (N_18490,N_17429,N_16622);
xnor U18491 (N_18491,N_16447,N_16534);
and U18492 (N_18492,N_16271,N_16832);
and U18493 (N_18493,N_17201,N_16735);
nand U18494 (N_18494,N_17391,N_16873);
xor U18495 (N_18495,N_16544,N_16410);
nor U18496 (N_18496,N_16447,N_16561);
and U18497 (N_18497,N_17431,N_17133);
nand U18498 (N_18498,N_16362,N_16568);
or U18499 (N_18499,N_16730,N_16947);
or U18500 (N_18500,N_16462,N_17273);
xnor U18501 (N_18501,N_16587,N_17239);
nor U18502 (N_18502,N_17027,N_16709);
and U18503 (N_18503,N_17144,N_17019);
and U18504 (N_18504,N_16365,N_16580);
and U18505 (N_18505,N_17179,N_16821);
nor U18506 (N_18506,N_16443,N_17353);
nor U18507 (N_18507,N_16292,N_16766);
nand U18508 (N_18508,N_17419,N_17468);
and U18509 (N_18509,N_16626,N_17469);
nand U18510 (N_18510,N_16547,N_16398);
nor U18511 (N_18511,N_16370,N_16318);
xor U18512 (N_18512,N_16655,N_16560);
or U18513 (N_18513,N_17302,N_17043);
or U18514 (N_18514,N_17485,N_17142);
nor U18515 (N_18515,N_17429,N_16438);
nor U18516 (N_18516,N_16786,N_16956);
nor U18517 (N_18517,N_17197,N_17044);
xor U18518 (N_18518,N_16583,N_16440);
and U18519 (N_18519,N_16682,N_16605);
nor U18520 (N_18520,N_16762,N_17056);
and U18521 (N_18521,N_17122,N_16390);
nand U18522 (N_18522,N_17131,N_17106);
and U18523 (N_18523,N_17009,N_17394);
and U18524 (N_18524,N_17148,N_16685);
xor U18525 (N_18525,N_16697,N_16685);
xnor U18526 (N_18526,N_16766,N_17274);
nor U18527 (N_18527,N_17057,N_16564);
and U18528 (N_18528,N_17394,N_16459);
or U18529 (N_18529,N_16617,N_17303);
nand U18530 (N_18530,N_17248,N_16291);
and U18531 (N_18531,N_16925,N_17304);
or U18532 (N_18532,N_16274,N_16904);
or U18533 (N_18533,N_17428,N_16689);
nand U18534 (N_18534,N_17316,N_17121);
or U18535 (N_18535,N_16986,N_16711);
or U18536 (N_18536,N_16308,N_16578);
nor U18537 (N_18537,N_17239,N_16428);
and U18538 (N_18538,N_17208,N_16709);
and U18539 (N_18539,N_16919,N_17232);
xnor U18540 (N_18540,N_16644,N_17006);
nand U18541 (N_18541,N_17113,N_17084);
or U18542 (N_18542,N_17422,N_17365);
nand U18543 (N_18543,N_16659,N_16807);
xnor U18544 (N_18544,N_16364,N_16302);
nand U18545 (N_18545,N_17168,N_17458);
or U18546 (N_18546,N_16285,N_16945);
nor U18547 (N_18547,N_16585,N_16652);
and U18548 (N_18548,N_17385,N_17156);
nand U18549 (N_18549,N_16912,N_16383);
and U18550 (N_18550,N_17432,N_16408);
nand U18551 (N_18551,N_16736,N_16836);
or U18552 (N_18552,N_16784,N_16342);
nor U18553 (N_18553,N_16832,N_16576);
nor U18554 (N_18554,N_16944,N_16364);
nand U18555 (N_18555,N_16820,N_16911);
and U18556 (N_18556,N_17073,N_17161);
or U18557 (N_18557,N_16704,N_16709);
and U18558 (N_18558,N_16279,N_16739);
or U18559 (N_18559,N_16410,N_17139);
or U18560 (N_18560,N_16445,N_17321);
or U18561 (N_18561,N_16549,N_16428);
nand U18562 (N_18562,N_17234,N_17246);
nor U18563 (N_18563,N_16418,N_17036);
or U18564 (N_18564,N_16469,N_17244);
or U18565 (N_18565,N_17131,N_16960);
and U18566 (N_18566,N_17086,N_17259);
and U18567 (N_18567,N_16597,N_17355);
or U18568 (N_18568,N_16795,N_17286);
or U18569 (N_18569,N_17396,N_16407);
and U18570 (N_18570,N_16644,N_16970);
xor U18571 (N_18571,N_16749,N_17214);
xor U18572 (N_18572,N_17342,N_17318);
nand U18573 (N_18573,N_17377,N_16632);
nand U18574 (N_18574,N_16392,N_16272);
nand U18575 (N_18575,N_17403,N_16501);
or U18576 (N_18576,N_17185,N_16814);
xor U18577 (N_18577,N_17189,N_17190);
nor U18578 (N_18578,N_16630,N_16822);
xnor U18579 (N_18579,N_16488,N_16275);
nand U18580 (N_18580,N_16357,N_16375);
nor U18581 (N_18581,N_17015,N_16979);
nand U18582 (N_18582,N_16599,N_17477);
nand U18583 (N_18583,N_17393,N_16543);
or U18584 (N_18584,N_17113,N_16609);
nand U18585 (N_18585,N_17269,N_17235);
and U18586 (N_18586,N_16476,N_16732);
or U18587 (N_18587,N_17350,N_16408);
nand U18588 (N_18588,N_17345,N_17461);
xnor U18589 (N_18589,N_16882,N_16469);
or U18590 (N_18590,N_16914,N_17451);
and U18591 (N_18591,N_17078,N_16619);
xor U18592 (N_18592,N_17305,N_17333);
and U18593 (N_18593,N_16459,N_17188);
xor U18594 (N_18594,N_16571,N_17474);
nand U18595 (N_18595,N_17019,N_16921);
or U18596 (N_18596,N_17005,N_16697);
nand U18597 (N_18597,N_16389,N_17365);
xnor U18598 (N_18598,N_16909,N_16672);
xnor U18599 (N_18599,N_16767,N_16819);
or U18600 (N_18600,N_17161,N_16599);
xor U18601 (N_18601,N_16970,N_16397);
xnor U18602 (N_18602,N_17190,N_16900);
xnor U18603 (N_18603,N_16499,N_16385);
or U18604 (N_18604,N_17303,N_16696);
and U18605 (N_18605,N_16313,N_16935);
nand U18606 (N_18606,N_16911,N_16788);
or U18607 (N_18607,N_16530,N_16420);
nand U18608 (N_18608,N_16833,N_17154);
or U18609 (N_18609,N_16357,N_16976);
nand U18610 (N_18610,N_16954,N_17363);
or U18611 (N_18611,N_16887,N_16716);
nand U18612 (N_18612,N_16823,N_16513);
or U18613 (N_18613,N_17044,N_16499);
nor U18614 (N_18614,N_16417,N_17011);
xor U18615 (N_18615,N_16839,N_17012);
and U18616 (N_18616,N_16929,N_16778);
nor U18617 (N_18617,N_17269,N_16866);
xnor U18618 (N_18618,N_16250,N_16666);
and U18619 (N_18619,N_16780,N_17107);
nor U18620 (N_18620,N_16291,N_16712);
xor U18621 (N_18621,N_17003,N_17172);
nor U18622 (N_18622,N_16871,N_16389);
xnor U18623 (N_18623,N_16733,N_16876);
and U18624 (N_18624,N_16964,N_17165);
nor U18625 (N_18625,N_16733,N_17057);
nor U18626 (N_18626,N_16322,N_16911);
xnor U18627 (N_18627,N_16962,N_16776);
xor U18628 (N_18628,N_16415,N_17200);
or U18629 (N_18629,N_16291,N_17076);
nand U18630 (N_18630,N_16344,N_16952);
xnor U18631 (N_18631,N_16570,N_16441);
or U18632 (N_18632,N_16477,N_16278);
or U18633 (N_18633,N_16898,N_17436);
xnor U18634 (N_18634,N_17086,N_16715);
or U18635 (N_18635,N_17036,N_16802);
nand U18636 (N_18636,N_16612,N_16571);
nand U18637 (N_18637,N_16962,N_16835);
xor U18638 (N_18638,N_16424,N_17186);
and U18639 (N_18639,N_16395,N_17231);
or U18640 (N_18640,N_16799,N_17471);
and U18641 (N_18641,N_16965,N_16302);
or U18642 (N_18642,N_17256,N_17240);
xnor U18643 (N_18643,N_17039,N_16929);
nor U18644 (N_18644,N_16326,N_16546);
or U18645 (N_18645,N_17311,N_17072);
xor U18646 (N_18646,N_16579,N_16378);
or U18647 (N_18647,N_16523,N_16921);
or U18648 (N_18648,N_16479,N_16323);
nor U18649 (N_18649,N_16864,N_17243);
nand U18650 (N_18650,N_16295,N_17227);
or U18651 (N_18651,N_16513,N_17290);
nand U18652 (N_18652,N_16519,N_17185);
nand U18653 (N_18653,N_17257,N_17371);
nand U18654 (N_18654,N_17285,N_17198);
nor U18655 (N_18655,N_17446,N_16552);
nor U18656 (N_18656,N_17472,N_16939);
and U18657 (N_18657,N_16386,N_16937);
nor U18658 (N_18658,N_17011,N_16563);
xnor U18659 (N_18659,N_16687,N_17440);
or U18660 (N_18660,N_17061,N_16685);
or U18661 (N_18661,N_16339,N_16345);
nand U18662 (N_18662,N_17413,N_16446);
or U18663 (N_18663,N_17400,N_17176);
xor U18664 (N_18664,N_17463,N_16640);
and U18665 (N_18665,N_17446,N_17150);
nand U18666 (N_18666,N_16519,N_17115);
nor U18667 (N_18667,N_16339,N_16471);
or U18668 (N_18668,N_17305,N_17313);
and U18669 (N_18669,N_17164,N_17238);
xor U18670 (N_18670,N_16758,N_17231);
nor U18671 (N_18671,N_16504,N_17006);
nor U18672 (N_18672,N_16286,N_16642);
or U18673 (N_18673,N_16806,N_17052);
xor U18674 (N_18674,N_17001,N_16685);
or U18675 (N_18675,N_17316,N_16498);
or U18676 (N_18676,N_16663,N_16586);
and U18677 (N_18677,N_16753,N_17339);
or U18678 (N_18678,N_17098,N_17163);
nor U18679 (N_18679,N_17181,N_16745);
and U18680 (N_18680,N_17027,N_16952);
nor U18681 (N_18681,N_17266,N_16544);
nand U18682 (N_18682,N_17459,N_16267);
xnor U18683 (N_18683,N_16752,N_16924);
or U18684 (N_18684,N_17408,N_16388);
and U18685 (N_18685,N_17404,N_17037);
and U18686 (N_18686,N_16402,N_17214);
or U18687 (N_18687,N_17187,N_17165);
nand U18688 (N_18688,N_16405,N_16850);
nor U18689 (N_18689,N_16980,N_17322);
xnor U18690 (N_18690,N_17464,N_17476);
nand U18691 (N_18691,N_16498,N_16477);
and U18692 (N_18692,N_16746,N_16749);
nand U18693 (N_18693,N_17270,N_17375);
xnor U18694 (N_18694,N_16435,N_16318);
and U18695 (N_18695,N_17397,N_17019);
nor U18696 (N_18696,N_16654,N_17279);
or U18697 (N_18697,N_17103,N_17399);
nor U18698 (N_18698,N_16982,N_17479);
and U18699 (N_18699,N_16449,N_17305);
xnor U18700 (N_18700,N_17006,N_16345);
and U18701 (N_18701,N_16320,N_16646);
or U18702 (N_18702,N_17036,N_16999);
or U18703 (N_18703,N_16365,N_17485);
nand U18704 (N_18704,N_17162,N_17397);
and U18705 (N_18705,N_16914,N_16927);
or U18706 (N_18706,N_16626,N_16937);
xnor U18707 (N_18707,N_17239,N_16448);
xnor U18708 (N_18708,N_17097,N_16467);
xnor U18709 (N_18709,N_17163,N_16674);
and U18710 (N_18710,N_16729,N_17178);
and U18711 (N_18711,N_16706,N_16661);
xor U18712 (N_18712,N_17219,N_16690);
nor U18713 (N_18713,N_16988,N_16365);
or U18714 (N_18714,N_16773,N_17412);
xnor U18715 (N_18715,N_16961,N_17462);
or U18716 (N_18716,N_16786,N_17149);
or U18717 (N_18717,N_16985,N_16729);
xor U18718 (N_18718,N_16805,N_16430);
or U18719 (N_18719,N_16897,N_16592);
xnor U18720 (N_18720,N_17295,N_17347);
or U18721 (N_18721,N_17045,N_16956);
or U18722 (N_18722,N_17231,N_16287);
xor U18723 (N_18723,N_16734,N_16832);
xnor U18724 (N_18724,N_16367,N_16554);
or U18725 (N_18725,N_17445,N_17334);
nand U18726 (N_18726,N_17324,N_17422);
or U18727 (N_18727,N_17379,N_17003);
xnor U18728 (N_18728,N_16927,N_16506);
nand U18729 (N_18729,N_16779,N_16451);
nor U18730 (N_18730,N_17297,N_16806);
and U18731 (N_18731,N_16440,N_16556);
nand U18732 (N_18732,N_17472,N_17082);
xor U18733 (N_18733,N_16902,N_16262);
xor U18734 (N_18734,N_16251,N_17076);
nor U18735 (N_18735,N_16294,N_16497);
xor U18736 (N_18736,N_16870,N_16889);
nand U18737 (N_18737,N_16821,N_16719);
or U18738 (N_18738,N_16605,N_16866);
and U18739 (N_18739,N_16714,N_17142);
nor U18740 (N_18740,N_17050,N_17444);
nand U18741 (N_18741,N_16328,N_17338);
and U18742 (N_18742,N_16616,N_17120);
nor U18743 (N_18743,N_16700,N_16534);
or U18744 (N_18744,N_16776,N_17164);
nand U18745 (N_18745,N_16533,N_16346);
xnor U18746 (N_18746,N_16913,N_17253);
nor U18747 (N_18747,N_16536,N_16445);
nor U18748 (N_18748,N_16731,N_16275);
nand U18749 (N_18749,N_16276,N_17301);
nor U18750 (N_18750,N_17970,N_17943);
nor U18751 (N_18751,N_17641,N_17590);
nor U18752 (N_18752,N_17861,N_18055);
nor U18753 (N_18753,N_17586,N_18463);
nor U18754 (N_18754,N_18267,N_18490);
nand U18755 (N_18755,N_18618,N_18241);
xnor U18756 (N_18756,N_17840,N_18140);
nand U18757 (N_18757,N_18624,N_18204);
nor U18758 (N_18758,N_18654,N_18659);
and U18759 (N_18759,N_17953,N_18308);
xor U18760 (N_18760,N_17775,N_17524);
nor U18761 (N_18761,N_18538,N_17695);
or U18762 (N_18762,N_18337,N_17838);
or U18763 (N_18763,N_18260,N_18229);
nor U18764 (N_18764,N_18275,N_17661);
and U18765 (N_18765,N_18284,N_18533);
and U18766 (N_18766,N_17922,N_18161);
nand U18767 (N_18767,N_18147,N_18743);
and U18768 (N_18768,N_18468,N_18334);
and U18769 (N_18769,N_17761,N_17688);
nor U18770 (N_18770,N_18655,N_18052);
or U18771 (N_18771,N_18724,N_18678);
xor U18772 (N_18772,N_17843,N_17879);
and U18773 (N_18773,N_18303,N_18113);
and U18774 (N_18774,N_17981,N_18461);
or U18775 (N_18775,N_17842,N_18549);
nor U18776 (N_18776,N_18142,N_17785);
nand U18777 (N_18777,N_18374,N_18112);
xnor U18778 (N_18778,N_18395,N_17573);
and U18779 (N_18779,N_17741,N_18180);
nor U18780 (N_18780,N_18477,N_18561);
xor U18781 (N_18781,N_18368,N_18221);
nor U18782 (N_18782,N_18686,N_17992);
or U18783 (N_18783,N_18351,N_17856);
and U18784 (N_18784,N_18746,N_17979);
xor U18785 (N_18785,N_18247,N_18721);
nor U18786 (N_18786,N_17958,N_18710);
and U18787 (N_18787,N_18285,N_17753);
nand U18788 (N_18788,N_18125,N_17938);
or U18789 (N_18789,N_18700,N_17621);
xor U18790 (N_18790,N_17703,N_18290);
and U18791 (N_18791,N_18223,N_18390);
or U18792 (N_18792,N_17694,N_17522);
nand U18793 (N_18793,N_18656,N_18363);
nor U18794 (N_18794,N_18118,N_17528);
and U18795 (N_18795,N_18551,N_17850);
nand U18796 (N_18796,N_18109,N_18547);
nor U18797 (N_18797,N_18070,N_17831);
and U18798 (N_18798,N_17950,N_18075);
or U18799 (N_18799,N_17713,N_18697);
xnor U18800 (N_18800,N_18729,N_18122);
and U18801 (N_18801,N_17540,N_17719);
nor U18802 (N_18802,N_18625,N_17585);
xor U18803 (N_18803,N_18029,N_18505);
nor U18804 (N_18804,N_17518,N_18708);
nor U18805 (N_18805,N_17508,N_17639);
or U18806 (N_18806,N_18545,N_17886);
and U18807 (N_18807,N_18025,N_17935);
nor U18808 (N_18808,N_17776,N_18424);
nand U18809 (N_18809,N_18471,N_18536);
or U18810 (N_18810,N_18610,N_17803);
nand U18811 (N_18811,N_17570,N_17902);
and U18812 (N_18812,N_18230,N_17867);
nand U18813 (N_18813,N_18612,N_17564);
xnor U18814 (N_18814,N_18018,N_18513);
nor U18815 (N_18815,N_18420,N_18234);
or U18816 (N_18816,N_17788,N_18094);
or U18817 (N_18817,N_17920,N_17746);
nand U18818 (N_18818,N_18263,N_17821);
and U18819 (N_18819,N_18085,N_18379);
or U18820 (N_18820,N_18535,N_18623);
or U18821 (N_18821,N_17516,N_18728);
nand U18822 (N_18822,N_18309,N_18346);
nand U18823 (N_18823,N_18064,N_18311);
and U18824 (N_18824,N_18130,N_17651);
or U18825 (N_18825,N_18205,N_17536);
or U18826 (N_18826,N_17642,N_18392);
and U18827 (N_18827,N_18009,N_17934);
nand U18828 (N_18828,N_17998,N_18176);
nand U18829 (N_18829,N_18145,N_18193);
xor U18830 (N_18830,N_18149,N_18671);
nor U18831 (N_18831,N_18555,N_18341);
or U18832 (N_18832,N_18053,N_17875);
nand U18833 (N_18833,N_17672,N_17566);
nand U18834 (N_18834,N_18670,N_17957);
nor U18835 (N_18835,N_17822,N_17510);
nand U18836 (N_18836,N_17645,N_17533);
and U18837 (N_18837,N_17773,N_18388);
nand U18838 (N_18838,N_18160,N_18736);
nand U18839 (N_18839,N_17725,N_18570);
or U18840 (N_18840,N_17544,N_18277);
and U18841 (N_18841,N_17655,N_17954);
or U18842 (N_18842,N_18375,N_18480);
nand U18843 (N_18843,N_18329,N_18298);
nor U18844 (N_18844,N_18074,N_18279);
nor U18845 (N_18845,N_17567,N_18579);
nand U18846 (N_18846,N_17561,N_18523);
nor U18847 (N_18847,N_17638,N_18376);
xnor U18848 (N_18848,N_18508,N_17738);
nor U18849 (N_18849,N_18104,N_17534);
nand U18850 (N_18850,N_18034,N_17551);
and U18851 (N_18851,N_18199,N_18464);
nor U18852 (N_18852,N_17808,N_18521);
xnor U18853 (N_18853,N_17600,N_17909);
and U18854 (N_18854,N_18627,N_18296);
xnor U18855 (N_18855,N_18639,N_18097);
nand U18856 (N_18856,N_18099,N_17851);
and U18857 (N_18857,N_17568,N_18294);
nand U18858 (N_18858,N_18599,N_18172);
xor U18859 (N_18859,N_18013,N_18428);
nand U18860 (N_18860,N_18592,N_17878);
and U18861 (N_18861,N_18493,N_18417);
or U18862 (N_18862,N_17759,N_18015);
nand U18863 (N_18863,N_18137,N_17976);
xnor U18864 (N_18864,N_18169,N_18452);
xnor U18865 (N_18865,N_18411,N_17668);
nor U18866 (N_18866,N_18698,N_17974);
xnor U18867 (N_18867,N_18462,N_17809);
nor U18868 (N_18868,N_18032,N_17597);
and U18869 (N_18869,N_17774,N_17825);
nand U18870 (N_18870,N_18295,N_18061);
xor U18871 (N_18871,N_18072,N_18119);
nor U18872 (N_18872,N_17892,N_17519);
and U18873 (N_18873,N_18430,N_18382);
nor U18874 (N_18874,N_18709,N_17982);
nand U18875 (N_18875,N_18386,N_18384);
or U18876 (N_18876,N_17891,N_18083);
and U18877 (N_18877,N_17849,N_18620);
nand U18878 (N_18878,N_17936,N_17735);
and U18879 (N_18879,N_18281,N_17669);
or U18880 (N_18880,N_18225,N_18722);
nand U18881 (N_18881,N_17880,N_18092);
or U18882 (N_18882,N_18051,N_17572);
or U18883 (N_18883,N_17846,N_17824);
xnor U18884 (N_18884,N_18011,N_17557);
nand U18885 (N_18885,N_17752,N_18177);
nand U18886 (N_18886,N_18262,N_17975);
xnor U18887 (N_18887,N_17833,N_17720);
nor U18888 (N_18888,N_18343,N_17614);
nand U18889 (N_18889,N_18259,N_17545);
nand U18890 (N_18890,N_18103,N_17962);
or U18891 (N_18891,N_18187,N_17576);
and U18892 (N_18892,N_17917,N_17784);
xnor U18893 (N_18893,N_18695,N_17529);
nor U18894 (N_18894,N_17659,N_18614);
or U18895 (N_18895,N_18682,N_18544);
and U18896 (N_18896,N_17717,N_18664);
or U18897 (N_18897,N_18691,N_17733);
nor U18898 (N_18898,N_18421,N_17637);
nor U18899 (N_18899,N_18398,N_18492);
nand U18900 (N_18900,N_18110,N_17754);
or U18901 (N_18901,N_17684,N_18423);
and U18902 (N_18902,N_18242,N_17852);
or U18903 (N_18903,N_17799,N_18058);
nor U18904 (N_18904,N_17829,N_18283);
and U18905 (N_18905,N_18338,N_18220);
and U18906 (N_18906,N_18453,N_18603);
and U18907 (N_18907,N_17689,N_17865);
and U18908 (N_18908,N_18228,N_17818);
xor U18909 (N_18909,N_18484,N_18393);
or U18910 (N_18910,N_18391,N_17952);
and U18911 (N_18911,N_17928,N_17523);
nor U18912 (N_18912,N_18261,N_17966);
nand U18913 (N_18913,N_18543,N_17514);
xor U18914 (N_18914,N_17630,N_17647);
xnor U18915 (N_18915,N_17571,N_17884);
nor U18916 (N_18916,N_18323,N_18626);
nor U18917 (N_18917,N_17827,N_18278);
nor U18918 (N_18918,N_18235,N_18608);
and U18919 (N_18919,N_18433,N_17959);
nor U18920 (N_18920,N_18226,N_18353);
nor U18921 (N_18921,N_17742,N_17805);
nor U18922 (N_18922,N_17780,N_18036);
nand U18923 (N_18923,N_17743,N_17736);
nor U18924 (N_18924,N_18106,N_18183);
nor U18925 (N_18925,N_18657,N_18280);
and U18926 (N_18926,N_18550,N_18131);
xor U18927 (N_18927,N_18356,N_17667);
or U18928 (N_18928,N_18159,N_18287);
nor U18929 (N_18929,N_18429,N_17705);
xor U18930 (N_18930,N_18560,N_17580);
nand U18931 (N_18931,N_18256,N_18566);
xor U18932 (N_18932,N_17648,N_18587);
and U18933 (N_18933,N_17628,N_18595);
or U18934 (N_18934,N_17558,N_17766);
nand U18935 (N_18935,N_18641,N_17758);
nor U18936 (N_18936,N_17757,N_17912);
or U18937 (N_18937,N_18213,N_18745);
xnor U18938 (N_18938,N_18252,N_18450);
or U18939 (N_18939,N_18040,N_18344);
nor U18940 (N_18940,N_18556,N_18133);
nand U18941 (N_18941,N_17673,N_18589);
or U18942 (N_18942,N_17560,N_18668);
nor U18943 (N_18943,N_18330,N_18258);
or U18944 (N_18944,N_18369,N_17587);
and U18945 (N_18945,N_17726,N_17960);
nand U18946 (N_18946,N_18292,N_18380);
nor U18947 (N_18947,N_18076,N_17947);
and U18948 (N_18948,N_18073,N_18186);
or U18949 (N_18949,N_18482,N_17665);
nand U18950 (N_18950,N_18370,N_17714);
xor U18951 (N_18951,N_18266,N_17916);
xnor U18952 (N_18952,N_17539,N_18470);
and U18953 (N_18953,N_18397,N_17697);
xnor U18954 (N_18954,N_18683,N_17887);
and U18955 (N_18955,N_18504,N_18321);
xnor U18956 (N_18956,N_18496,N_18658);
xor U18957 (N_18957,N_17677,N_18095);
nand U18958 (N_18958,N_17834,N_18748);
or U18959 (N_18959,N_17986,N_17881);
xor U18960 (N_18960,N_18647,N_18518);
nor U18961 (N_18961,N_18232,N_18030);
xnor U18962 (N_18962,N_18552,N_17893);
or U18963 (N_18963,N_17712,N_17800);
or U18964 (N_18964,N_17595,N_17543);
nor U18965 (N_18965,N_17857,N_18738);
or U18966 (N_18966,N_18134,N_18043);
nand U18967 (N_18967,N_17807,N_18439);
nor U18968 (N_18968,N_17617,N_17964);
or U18969 (N_18969,N_18066,N_18609);
nand U18970 (N_18970,N_17955,N_18690);
and U18971 (N_18971,N_18002,N_18243);
nor U18972 (N_18972,N_18527,N_18102);
nor U18973 (N_18973,N_18486,N_18387);
and U18974 (N_18974,N_18385,N_18336);
and U18975 (N_18975,N_17579,N_18063);
and U18976 (N_18976,N_18707,N_17888);
nor U18977 (N_18977,N_17961,N_18081);
nand U18978 (N_18978,N_17599,N_17940);
or U18979 (N_18979,N_18182,N_17869);
nand U18980 (N_18980,N_18617,N_17899);
nor U18981 (N_18981,N_18675,N_18444);
nand U18982 (N_18982,N_18004,N_17941);
or U18983 (N_18983,N_18373,N_18202);
and U18984 (N_18984,N_18568,N_18189);
nor U18985 (N_18985,N_17509,N_17820);
nor U18986 (N_18986,N_17619,N_18636);
and U18987 (N_18987,N_18737,N_18209);
nor U18988 (N_18988,N_18162,N_17721);
and U18989 (N_18989,N_18231,N_18715);
nor U18990 (N_18990,N_17797,N_17565);
or U18991 (N_18991,N_18522,N_18151);
nor U18992 (N_18992,N_17606,N_18567);
nand U18993 (N_18993,N_17882,N_17744);
xnor U18994 (N_18994,N_18537,N_18196);
and U18995 (N_18995,N_18600,N_18315);
nand U18996 (N_18996,N_17646,N_18157);
and U18997 (N_18997,N_18512,N_17636);
nor U18998 (N_18998,N_17872,N_18335);
or U18999 (N_18999,N_17795,N_18179);
xor U19000 (N_19000,N_17601,N_17730);
or U19001 (N_19001,N_18489,N_18185);
or U19002 (N_19002,N_18451,N_18141);
nor U19003 (N_19003,N_17520,N_17501);
nor U19004 (N_19004,N_18057,N_17983);
and U19005 (N_19005,N_18101,N_18306);
and U19006 (N_19006,N_17620,N_17790);
nand U19007 (N_19007,N_17613,N_18272);
nor U19008 (N_19008,N_18704,N_17683);
or U19009 (N_19009,N_18622,N_17789);
xor U19010 (N_19010,N_18476,N_18687);
and U19011 (N_19011,N_17811,N_17512);
xnor U19012 (N_19012,N_17608,N_18498);
or U19013 (N_19013,N_18509,N_18465);
xor U19014 (N_19014,N_18514,N_18553);
and U19015 (N_19015,N_17830,N_17678);
and U19016 (N_19016,N_17546,N_18297);
nor U19017 (N_19017,N_17542,N_17710);
nor U19018 (N_19018,N_17696,N_18328);
and U19019 (N_19019,N_18100,N_18449);
or U19020 (N_19020,N_18676,N_17691);
nand U19021 (N_19021,N_18605,N_17762);
or U19022 (N_19022,N_17749,N_18249);
nand U19023 (N_19023,N_18046,N_18607);
nand U19024 (N_19024,N_18679,N_18405);
nor U19025 (N_19025,N_17836,N_18250);
and U19026 (N_19026,N_17709,N_17552);
xnor U19027 (N_19027,N_18293,N_18717);
and U19028 (N_19028,N_18733,N_17903);
or U19029 (N_19029,N_18497,N_18559);
xor U19030 (N_19030,N_18028,N_17883);
nand U19031 (N_19031,N_18383,N_17679);
or U19032 (N_19032,N_18271,N_17685);
and U19033 (N_19033,N_17837,N_17716);
nand U19034 (N_19034,N_17594,N_18431);
and U19035 (N_19035,N_17707,N_18662);
nor U19036 (N_19036,N_17708,N_17793);
nor U19037 (N_19037,N_17589,N_17658);
nor U19038 (N_19038,N_17819,N_18720);
xnor U19039 (N_19039,N_18558,N_17698);
xnor U19040 (N_19040,N_17755,N_17578);
and U19041 (N_19041,N_18005,N_18744);
nand U19042 (N_19042,N_17817,N_18197);
nor U19043 (N_19043,N_18467,N_18019);
nand U19044 (N_19044,N_18239,N_18472);
and U19045 (N_19045,N_17871,N_17898);
or U19046 (N_19046,N_18584,N_17631);
nand U19047 (N_19047,N_17907,N_18577);
and U19048 (N_19048,N_18153,N_17972);
nand U19049 (N_19049,N_17693,N_18727);
or U19050 (N_19050,N_18093,N_17905);
nand U19051 (N_19051,N_18143,N_18646);
nor U19052 (N_19052,N_18020,N_17993);
and U19053 (N_19053,N_18152,N_18396);
xnor U19054 (N_19054,N_18590,N_18166);
and U19055 (N_19055,N_17791,N_18065);
nand U19056 (N_19056,N_17618,N_18500);
xnor U19057 (N_19057,N_17999,N_18460);
xnor U19058 (N_19058,N_18310,N_17692);
nand U19059 (N_19059,N_18546,N_18680);
and U19060 (N_19060,N_18079,N_18517);
and U19061 (N_19061,N_17581,N_18684);
xnor U19062 (N_19062,N_18615,N_18479);
nor U19063 (N_19063,N_18254,N_17503);
and U19064 (N_19064,N_17554,N_17745);
nor U19065 (N_19065,N_18454,N_18007);
and U19066 (N_19066,N_18069,N_18441);
xnor U19067 (N_19067,N_18583,N_18701);
nor U19068 (N_19068,N_17847,N_17656);
nor U19069 (N_19069,N_18339,N_17575);
xor U19070 (N_19070,N_18006,N_18115);
xor U19071 (N_19071,N_17796,N_17666);
or U19072 (N_19072,N_17990,N_17681);
and U19073 (N_19073,N_18510,N_18206);
and U19074 (N_19074,N_18173,N_18619);
nor U19075 (N_19075,N_17911,N_17676);
xor U19076 (N_19076,N_18148,N_18731);
and U19077 (N_19077,N_17945,N_18473);
and U19078 (N_19078,N_17663,N_18457);
and U19079 (N_19079,N_18437,N_17813);
nand U19080 (N_19080,N_18352,N_18163);
or U19081 (N_19081,N_18693,N_18082);
and U19082 (N_19082,N_18154,N_18347);
nor U19083 (N_19083,N_17783,N_18077);
or U19084 (N_19084,N_17627,N_18406);
nor U19085 (N_19085,N_17591,N_18361);
or U19086 (N_19086,N_17980,N_18714);
xor U19087 (N_19087,N_18650,N_18672);
nor U19088 (N_19088,N_17779,N_18132);
or U19089 (N_19089,N_18503,N_18067);
nor U19090 (N_19090,N_18024,N_18367);
and U19091 (N_19091,N_18240,N_17701);
nor U19092 (N_19092,N_18144,N_17702);
and U19093 (N_19093,N_18696,N_18105);
nor U19094 (N_19094,N_17946,N_18635);
or U19095 (N_19095,N_18569,N_17967);
or U19096 (N_19096,N_18107,N_17812);
and U19097 (N_19097,N_17640,N_17728);
nor U19098 (N_19098,N_17996,N_18416);
or U19099 (N_19099,N_17722,N_18371);
or U19100 (N_19100,N_17505,N_18192);
xor U19101 (N_19101,N_18021,N_18571);
nand U19102 (N_19102,N_17772,N_17866);
nand U19103 (N_19103,N_18060,N_17860);
nand U19104 (N_19104,N_17874,N_18435);
or U19105 (N_19105,N_17547,N_18319);
nand U19106 (N_19106,N_18087,N_17863);
or U19107 (N_19107,N_17930,N_18528);
nor U19108 (N_19108,N_17626,N_18312);
xor U19109 (N_19109,N_17751,N_17848);
nand U19110 (N_19110,N_17854,N_18171);
and U19111 (N_19111,N_18524,N_18120);
nand U19112 (N_19112,N_18129,N_18591);
and U19113 (N_19113,N_17632,N_17984);
nand U19114 (N_19114,N_18224,N_18730);
xor U19115 (N_19115,N_17802,N_18372);
xor U19116 (N_19116,N_17969,N_18487);
or U19117 (N_19117,N_18410,N_18348);
xnor U19118 (N_19118,N_18214,N_17515);
xnor U19119 (N_19119,N_18349,N_18170);
or U19120 (N_19120,N_18354,N_17937);
xor U19121 (N_19121,N_18364,N_18529);
nand U19122 (N_19122,N_17908,N_18459);
nor U19123 (N_19123,N_17674,N_17914);
nor U19124 (N_19124,N_18652,N_17616);
nand U19125 (N_19125,N_18314,N_18359);
nor U19126 (N_19126,N_17664,N_18282);
nand U19127 (N_19127,N_18026,N_18155);
xnor U19128 (N_19128,N_17569,N_17765);
and U19129 (N_19129,N_18150,N_18685);
or U19130 (N_19130,N_18702,N_18366);
nand U19131 (N_19131,N_18474,N_18404);
nor U19132 (N_19132,N_18041,N_17901);
or U19133 (N_19133,N_17657,N_18207);
xnor U19134 (N_19134,N_18201,N_18488);
and U19135 (N_19135,N_17926,N_17506);
xor U19136 (N_19136,N_18270,N_18723);
xor U19137 (N_19137,N_17770,N_18236);
or U19138 (N_19138,N_18403,N_17718);
nor U19139 (N_19139,N_17971,N_18059);
nor U19140 (N_19140,N_18276,N_18594);
nor U19141 (N_19141,N_17949,N_18578);
nand U19142 (N_19142,N_18016,N_18212);
xor U19143 (N_19143,N_18313,N_18237);
or U19144 (N_19144,N_18017,N_18634);
and U19145 (N_19145,N_17801,N_18531);
xor U19146 (N_19146,N_18126,N_17624);
and U19147 (N_19147,N_18322,N_18644);
nor U19148 (N_19148,N_18222,N_18638);
or U19149 (N_19149,N_18300,N_18432);
and U19150 (N_19150,N_18084,N_18211);
nor U19151 (N_19151,N_17792,N_18741);
or U19152 (N_19152,N_17781,N_18649);
nand U19153 (N_19153,N_18665,N_18502);
nor U19154 (N_19154,N_17731,N_17931);
xnor U19155 (N_19155,N_17649,N_17704);
and U19156 (N_19156,N_17629,N_18495);
or U19157 (N_19157,N_18062,N_18557);
xnor U19158 (N_19158,N_17517,N_17988);
and U19159 (N_19159,N_18711,N_18585);
and U19160 (N_19160,N_17997,N_18673);
and U19161 (N_19161,N_18168,N_17804);
and U19162 (N_19162,N_18588,N_18190);
and U19163 (N_19163,N_17826,N_18540);
or U19164 (N_19164,N_18056,N_17635);
nand U19165 (N_19165,N_18245,N_17526);
nand U19166 (N_19166,N_17844,N_18394);
and U19167 (N_19167,N_18291,N_18705);
and U19168 (N_19168,N_18340,N_18191);
or U19169 (N_19169,N_17611,N_18400);
nor U19170 (N_19170,N_17913,N_18001);
nand U19171 (N_19171,N_17723,N_17690);
xnor U19172 (N_19172,N_17652,N_18307);
nand U19173 (N_19173,N_18541,N_17845);
xor U19174 (N_19174,N_17769,N_17915);
nor U19175 (N_19175,N_17634,N_17607);
nand U19176 (N_19176,N_17864,N_18175);
nor U19177 (N_19177,N_18613,N_17747);
xnor U19178 (N_19178,N_18726,N_18516);
nor U19179 (N_19179,N_18358,N_17994);
or U19180 (N_19180,N_17732,N_18640);
nor U19181 (N_19181,N_18038,N_18506);
and U19182 (N_19182,N_18299,N_17633);
nor U19183 (N_19183,N_18629,N_18507);
xnor U19184 (N_19184,N_17987,N_18088);
nor U19185 (N_19185,N_17748,N_17615);
nand U19186 (N_19186,N_18269,N_18739);
nand U19187 (N_19187,N_17859,N_18653);
and U19188 (N_19188,N_18611,N_18688);
or U19189 (N_19189,N_18203,N_17711);
or U19190 (N_19190,N_18520,N_18326);
nor U19191 (N_19191,N_18478,N_17625);
nor U19192 (N_19192,N_18572,N_17923);
xor U19193 (N_19193,N_18712,N_17686);
xor U19194 (N_19194,N_18289,N_17927);
xnor U19195 (N_19195,N_17680,N_17858);
nor U19196 (N_19196,N_17729,N_17504);
nand U19197 (N_19197,N_17548,N_18469);
nand U19198 (N_19198,N_18581,N_18286);
or U19199 (N_19199,N_18445,N_17868);
nand U19200 (N_19200,N_17556,N_18677);
nand U19201 (N_19201,N_18216,N_17995);
and U19202 (N_19202,N_17577,N_18381);
xor U19203 (N_19203,N_17574,N_18481);
or U19204 (N_19204,N_18035,N_18045);
xor U19205 (N_19205,N_18436,N_17963);
or U19206 (N_19206,N_17653,N_18357);
nor U19207 (N_19207,N_17918,N_17610);
or U19208 (N_19208,N_18548,N_18438);
nor U19209 (N_19209,N_18117,N_18174);
nor U19210 (N_19210,N_18458,N_18606);
or U19211 (N_19211,N_18532,N_18325);
xor U19212 (N_19212,N_17675,N_18123);
nor U19213 (N_19213,N_18633,N_17734);
nand U19214 (N_19214,N_17562,N_18345);
xor U19215 (N_19215,N_18217,N_18719);
nand U19216 (N_19216,N_18494,N_17876);
and U19217 (N_19217,N_17764,N_18248);
and U19218 (N_19218,N_18331,N_18023);
nor U19219 (N_19219,N_18257,N_18033);
nand U19220 (N_19220,N_18539,N_17596);
nor U19221 (N_19221,N_18651,N_17900);
and U19222 (N_19222,N_17737,N_17550);
nand U19223 (N_19223,N_17782,N_18596);
xor U19224 (N_19224,N_17910,N_18342);
nand U19225 (N_19225,N_18184,N_18574);
or U19226 (N_19226,N_18573,N_18426);
xnor U19227 (N_19227,N_18740,N_17604);
nor U19228 (N_19228,N_18499,N_18068);
xor U19229 (N_19229,N_18320,N_18027);
xnor U19230 (N_19230,N_18455,N_17740);
and U19231 (N_19231,N_18412,N_18318);
nand U19232 (N_19232,N_17985,N_17767);
and U19233 (N_19233,N_18542,N_18227);
and U19234 (N_19234,N_17989,N_18165);
nand U19235 (N_19235,N_18194,N_18415);
xnor U19236 (N_19236,N_18602,N_17760);
and U19237 (N_19237,N_17538,N_18317);
or U19238 (N_19238,N_18604,N_18660);
or U19239 (N_19239,N_18418,N_18219);
or U19240 (N_19240,N_18402,N_18111);
nand U19241 (N_19241,N_17870,N_18138);
and U19242 (N_19242,N_18526,N_18554);
and U19243 (N_19243,N_17592,N_17602);
xnor U19244 (N_19244,N_18050,N_18188);
or U19245 (N_19245,N_17877,N_18408);
nand U19246 (N_19246,N_17527,N_17816);
nor U19247 (N_19247,N_17682,N_18401);
nand U19248 (N_19248,N_18265,N_17890);
nand U19249 (N_19249,N_18483,N_17612);
and U19250 (N_19250,N_17549,N_17814);
or U19251 (N_19251,N_17806,N_17777);
and U19252 (N_19252,N_18098,N_18689);
or U19253 (N_19253,N_17724,N_18389);
nor U19254 (N_19254,N_18139,N_17644);
and U19255 (N_19255,N_18598,N_18749);
nand U19256 (N_19256,N_18316,N_17660);
and U19257 (N_19257,N_18442,N_17978);
xnor U19258 (N_19258,N_17933,N_17853);
and U19259 (N_19259,N_18674,N_17786);
nand U19260 (N_19260,N_18049,N_18515);
nor U19261 (N_19261,N_18008,N_17921);
nor U19262 (N_19262,N_18511,N_18501);
and U19263 (N_19263,N_17977,N_18666);
and U19264 (N_19264,N_18648,N_17895);
or U19265 (N_19265,N_17991,N_17559);
and U19266 (N_19266,N_17839,N_18443);
xnor U19267 (N_19267,N_17896,N_18114);
nor U19268 (N_19268,N_18440,N_18425);
nor U19269 (N_19269,N_18593,N_17798);
or U19270 (N_19270,N_18246,N_18564);
xnor U19271 (N_19271,N_18663,N_18350);
nand U19272 (N_19272,N_17555,N_17885);
nand U19273 (N_19273,N_18399,N_18096);
nor U19274 (N_19274,N_18365,N_17951);
xor U19275 (N_19275,N_17906,N_17904);
or U19276 (N_19276,N_18333,N_18378);
or U19277 (N_19277,N_17794,N_18218);
xor U19278 (N_19278,N_17944,N_17521);
and U19279 (N_19279,N_18667,N_17932);
and U19280 (N_19280,N_17815,N_17507);
and U19281 (N_19281,N_18732,N_18661);
xnor U19282 (N_19282,N_17699,N_18014);
nand U19283 (N_19283,N_18012,N_18718);
nor U19284 (N_19284,N_17778,N_17919);
and U19285 (N_19285,N_18047,N_17873);
nand U19286 (N_19286,N_18268,N_18244);
or U19287 (N_19287,N_18210,N_18124);
or U19288 (N_19288,N_18706,N_18238);
and U19289 (N_19289,N_17541,N_17968);
nand U19290 (N_19290,N_17700,N_17750);
xnor U19291 (N_19291,N_18642,N_18645);
nand U19292 (N_19292,N_18000,N_18108);
nor U19293 (N_19293,N_18360,N_18447);
or U19294 (N_19294,N_17828,N_17553);
and U19295 (N_19295,N_17650,N_17810);
and U19296 (N_19296,N_18562,N_18301);
and U19297 (N_19297,N_17835,N_18534);
nor U19298 (N_19298,N_18576,N_18485);
or U19299 (N_19299,N_17855,N_18409);
or U19300 (N_19300,N_17841,N_18586);
xnor U19301 (N_19301,N_18288,N_17588);
and U19302 (N_19302,N_17535,N_18616);
xor U19303 (N_19303,N_18327,N_17925);
nand U19304 (N_19304,N_17513,N_18699);
or U19305 (N_19305,N_17739,N_17706);
nor U19306 (N_19306,N_18044,N_18669);
xnor U19307 (N_19307,N_18621,N_18734);
nor U19308 (N_19308,N_18377,N_18198);
and U19309 (N_19309,N_17862,N_18010);
or U19310 (N_19310,N_18195,N_17662);
or U19311 (N_19311,N_18264,N_17525);
and U19312 (N_19312,N_18446,N_18273);
nand U19313 (N_19313,N_18200,N_17532);
nor U19314 (N_19314,N_17832,N_18601);
xnor U19315 (N_19315,N_17942,N_18630);
or U19316 (N_19316,N_18692,N_18178);
xnor U19317 (N_19317,N_18054,N_18434);
and U19318 (N_19318,N_18091,N_18215);
xor U19319 (N_19319,N_18694,N_18031);
nor U19320 (N_19320,N_18089,N_18039);
or U19321 (N_19321,N_18407,N_17511);
nand U19322 (N_19322,N_18637,N_17500);
and U19323 (N_19323,N_18164,N_18048);
xnor U19324 (N_19324,N_17756,N_17531);
xor U19325 (N_19325,N_18681,N_18156);
xor U19326 (N_19326,N_17889,N_18582);
nor U19327 (N_19327,N_17502,N_18419);
nand U19328 (N_19328,N_18116,N_17973);
xor U19329 (N_19329,N_17563,N_18233);
or U19330 (N_19330,N_18597,N_18071);
and U19331 (N_19331,N_18078,N_17768);
nor U19332 (N_19332,N_17582,N_18563);
nor U19333 (N_19333,N_17583,N_18090);
nand U19334 (N_19334,N_18146,N_18362);
or U19335 (N_19335,N_18003,N_18037);
xnor U19336 (N_19336,N_17727,N_17603);
nand U19337 (N_19337,N_17609,N_18135);
nand U19338 (N_19338,N_18080,N_18302);
xor U19339 (N_19339,N_18631,N_17894);
xnor U19340 (N_19340,N_17598,N_18448);
nor U19341 (N_19341,N_18713,N_17771);
nand U19342 (N_19342,N_17593,N_18475);
or U19343 (N_19343,N_17897,N_17622);
xor U19344 (N_19344,N_17715,N_17671);
or U19345 (N_19345,N_18355,N_17537);
and U19346 (N_19346,N_17687,N_17763);
or U19347 (N_19347,N_18128,N_18456);
nor U19348 (N_19348,N_18427,N_17929);
nand U19349 (N_19349,N_18274,N_18305);
xor U19350 (N_19350,N_18575,N_18158);
or U19351 (N_19351,N_18332,N_18167);
or U19352 (N_19352,N_18525,N_17823);
nor U19353 (N_19353,N_18643,N_18580);
nand U19354 (N_19354,N_18324,N_18466);
nand U19355 (N_19355,N_18208,N_18121);
and U19356 (N_19356,N_18086,N_18127);
and U19357 (N_19357,N_17965,N_18042);
and U19358 (N_19358,N_18735,N_17623);
or U19359 (N_19359,N_18742,N_17939);
xnor U19360 (N_19360,N_17605,N_18022);
or U19361 (N_19361,N_18703,N_17787);
xnor U19362 (N_19362,N_17643,N_18628);
and U19363 (N_19363,N_18251,N_17670);
and U19364 (N_19364,N_18422,N_17530);
nand U19365 (N_19365,N_17924,N_18530);
nor U19366 (N_19366,N_18632,N_18519);
nand U19367 (N_19367,N_18255,N_17948);
nor U19368 (N_19368,N_18565,N_18747);
and U19369 (N_19369,N_18414,N_18253);
nand U19370 (N_19370,N_18716,N_18491);
or U19371 (N_19371,N_17654,N_18413);
nor U19372 (N_19372,N_18304,N_17584);
nor U19373 (N_19373,N_18136,N_17956);
and U19374 (N_19374,N_18725,N_18181);
xnor U19375 (N_19375,N_18159,N_18510);
nor U19376 (N_19376,N_18654,N_18266);
nand U19377 (N_19377,N_18254,N_17578);
and U19378 (N_19378,N_18172,N_18269);
nand U19379 (N_19379,N_17890,N_18156);
or U19380 (N_19380,N_17817,N_18456);
and U19381 (N_19381,N_17658,N_17577);
and U19382 (N_19382,N_18593,N_17914);
xnor U19383 (N_19383,N_17964,N_18615);
nand U19384 (N_19384,N_18086,N_17870);
or U19385 (N_19385,N_18622,N_17689);
xnor U19386 (N_19386,N_17813,N_17977);
nor U19387 (N_19387,N_18365,N_18033);
nand U19388 (N_19388,N_18251,N_17882);
nand U19389 (N_19389,N_18320,N_18463);
nor U19390 (N_19390,N_17946,N_17921);
nor U19391 (N_19391,N_18662,N_18040);
or U19392 (N_19392,N_18553,N_18344);
xor U19393 (N_19393,N_18385,N_17600);
nor U19394 (N_19394,N_18341,N_18633);
or U19395 (N_19395,N_18194,N_18146);
nor U19396 (N_19396,N_17837,N_17766);
xor U19397 (N_19397,N_18640,N_18052);
or U19398 (N_19398,N_17975,N_18147);
xnor U19399 (N_19399,N_17978,N_17777);
nor U19400 (N_19400,N_18181,N_18019);
or U19401 (N_19401,N_17666,N_17831);
nand U19402 (N_19402,N_18244,N_18661);
nor U19403 (N_19403,N_18633,N_18026);
nand U19404 (N_19404,N_18215,N_18370);
nor U19405 (N_19405,N_18746,N_18544);
xor U19406 (N_19406,N_18311,N_18361);
nand U19407 (N_19407,N_17681,N_17895);
nand U19408 (N_19408,N_17588,N_18106);
or U19409 (N_19409,N_17737,N_18121);
or U19410 (N_19410,N_17945,N_18249);
nor U19411 (N_19411,N_18219,N_18075);
nor U19412 (N_19412,N_17858,N_18561);
or U19413 (N_19413,N_17699,N_18570);
nor U19414 (N_19414,N_18355,N_18547);
or U19415 (N_19415,N_17744,N_18701);
or U19416 (N_19416,N_18539,N_18370);
nor U19417 (N_19417,N_18583,N_17612);
or U19418 (N_19418,N_18489,N_18623);
xnor U19419 (N_19419,N_18003,N_17775);
nor U19420 (N_19420,N_17827,N_18440);
or U19421 (N_19421,N_17988,N_18109);
nor U19422 (N_19422,N_18737,N_18265);
nor U19423 (N_19423,N_18556,N_18451);
nor U19424 (N_19424,N_17676,N_17632);
xor U19425 (N_19425,N_17600,N_18203);
xnor U19426 (N_19426,N_18288,N_17531);
nand U19427 (N_19427,N_17917,N_18349);
or U19428 (N_19428,N_17993,N_18597);
xnor U19429 (N_19429,N_18355,N_18047);
xnor U19430 (N_19430,N_18442,N_18103);
or U19431 (N_19431,N_17793,N_17754);
or U19432 (N_19432,N_18279,N_17522);
nand U19433 (N_19433,N_18605,N_18343);
or U19434 (N_19434,N_17730,N_17807);
and U19435 (N_19435,N_18324,N_18265);
nand U19436 (N_19436,N_17932,N_18221);
or U19437 (N_19437,N_18425,N_18083);
xnor U19438 (N_19438,N_18199,N_18262);
and U19439 (N_19439,N_18019,N_17717);
nand U19440 (N_19440,N_17749,N_17769);
xnor U19441 (N_19441,N_17732,N_18010);
or U19442 (N_19442,N_17716,N_18721);
and U19443 (N_19443,N_18672,N_17784);
xnor U19444 (N_19444,N_18288,N_17775);
nand U19445 (N_19445,N_17930,N_18217);
or U19446 (N_19446,N_17948,N_18408);
and U19447 (N_19447,N_17588,N_17807);
or U19448 (N_19448,N_18305,N_18159);
nand U19449 (N_19449,N_18587,N_18742);
or U19450 (N_19450,N_18370,N_17675);
or U19451 (N_19451,N_18561,N_17818);
xor U19452 (N_19452,N_18099,N_17895);
nand U19453 (N_19453,N_17832,N_17991);
xor U19454 (N_19454,N_18016,N_18267);
nor U19455 (N_19455,N_17526,N_17549);
xnor U19456 (N_19456,N_17578,N_18395);
nor U19457 (N_19457,N_18053,N_18698);
xor U19458 (N_19458,N_18299,N_18640);
or U19459 (N_19459,N_17721,N_18312);
or U19460 (N_19460,N_17944,N_18176);
or U19461 (N_19461,N_18270,N_18160);
xor U19462 (N_19462,N_17809,N_17841);
or U19463 (N_19463,N_18743,N_18236);
or U19464 (N_19464,N_18623,N_18687);
xnor U19465 (N_19465,N_17763,N_18084);
xnor U19466 (N_19466,N_18644,N_18615);
xor U19467 (N_19467,N_18471,N_17759);
nor U19468 (N_19468,N_18053,N_17710);
and U19469 (N_19469,N_18169,N_17812);
nor U19470 (N_19470,N_17912,N_18410);
nand U19471 (N_19471,N_18117,N_18033);
and U19472 (N_19472,N_17561,N_18733);
nand U19473 (N_19473,N_17895,N_18509);
nand U19474 (N_19474,N_17839,N_18738);
and U19475 (N_19475,N_18304,N_17826);
nor U19476 (N_19476,N_18012,N_18081);
nand U19477 (N_19477,N_18531,N_18668);
nand U19478 (N_19478,N_18611,N_18525);
and U19479 (N_19479,N_18443,N_18446);
or U19480 (N_19480,N_18566,N_17860);
xor U19481 (N_19481,N_18051,N_17509);
nor U19482 (N_19482,N_17646,N_18228);
xnor U19483 (N_19483,N_18235,N_17719);
and U19484 (N_19484,N_17748,N_17862);
nor U19485 (N_19485,N_18514,N_18471);
or U19486 (N_19486,N_17501,N_18548);
or U19487 (N_19487,N_17625,N_18231);
xnor U19488 (N_19488,N_17668,N_17533);
nand U19489 (N_19489,N_17765,N_17972);
nand U19490 (N_19490,N_18243,N_18544);
xnor U19491 (N_19491,N_17582,N_18346);
and U19492 (N_19492,N_17543,N_18540);
xor U19493 (N_19493,N_17505,N_17585);
and U19494 (N_19494,N_17911,N_18400);
and U19495 (N_19495,N_18723,N_18180);
xor U19496 (N_19496,N_18411,N_17540);
nor U19497 (N_19497,N_17636,N_18317);
xor U19498 (N_19498,N_18424,N_18318);
xnor U19499 (N_19499,N_18085,N_18136);
and U19500 (N_19500,N_18530,N_17543);
nand U19501 (N_19501,N_18187,N_17679);
xor U19502 (N_19502,N_17866,N_18496);
and U19503 (N_19503,N_17680,N_18025);
nand U19504 (N_19504,N_17557,N_17982);
nor U19505 (N_19505,N_18304,N_18586);
xnor U19506 (N_19506,N_17512,N_17948);
or U19507 (N_19507,N_18352,N_18095);
nor U19508 (N_19508,N_17861,N_17834);
and U19509 (N_19509,N_17662,N_17803);
nor U19510 (N_19510,N_18129,N_18582);
and U19511 (N_19511,N_17673,N_17803);
and U19512 (N_19512,N_17501,N_18264);
or U19513 (N_19513,N_18742,N_18700);
xnor U19514 (N_19514,N_18518,N_18612);
xor U19515 (N_19515,N_17670,N_17900);
and U19516 (N_19516,N_18018,N_17637);
xor U19517 (N_19517,N_18442,N_17740);
xnor U19518 (N_19518,N_17597,N_17895);
nor U19519 (N_19519,N_18034,N_17666);
xor U19520 (N_19520,N_17774,N_18498);
and U19521 (N_19521,N_18139,N_18295);
xnor U19522 (N_19522,N_18022,N_17524);
and U19523 (N_19523,N_18463,N_18650);
or U19524 (N_19524,N_17990,N_18180);
nand U19525 (N_19525,N_18714,N_18224);
and U19526 (N_19526,N_17927,N_18119);
and U19527 (N_19527,N_18721,N_17750);
and U19528 (N_19528,N_17996,N_18632);
nand U19529 (N_19529,N_18381,N_18544);
nand U19530 (N_19530,N_17679,N_17968);
xor U19531 (N_19531,N_18233,N_17671);
and U19532 (N_19532,N_18128,N_17529);
and U19533 (N_19533,N_18225,N_17786);
nand U19534 (N_19534,N_18743,N_17624);
nor U19535 (N_19535,N_18347,N_18710);
and U19536 (N_19536,N_17913,N_18605);
nand U19537 (N_19537,N_18657,N_17700);
nand U19538 (N_19538,N_17979,N_18226);
xnor U19539 (N_19539,N_18553,N_18724);
nor U19540 (N_19540,N_18144,N_18567);
nor U19541 (N_19541,N_18703,N_18202);
xnor U19542 (N_19542,N_18215,N_18548);
nand U19543 (N_19543,N_18610,N_17800);
and U19544 (N_19544,N_18202,N_17697);
nor U19545 (N_19545,N_17662,N_18219);
nand U19546 (N_19546,N_17984,N_18231);
nand U19547 (N_19547,N_17956,N_18517);
and U19548 (N_19548,N_18091,N_17760);
nor U19549 (N_19549,N_18673,N_18229);
and U19550 (N_19550,N_17962,N_17533);
or U19551 (N_19551,N_18521,N_18061);
or U19552 (N_19552,N_18279,N_17981);
nor U19553 (N_19553,N_18612,N_17633);
and U19554 (N_19554,N_18724,N_18614);
xnor U19555 (N_19555,N_18130,N_18514);
xnor U19556 (N_19556,N_18096,N_18031);
nand U19557 (N_19557,N_17617,N_18552);
nand U19558 (N_19558,N_17666,N_18450);
and U19559 (N_19559,N_17989,N_18421);
or U19560 (N_19560,N_18298,N_18584);
nor U19561 (N_19561,N_17582,N_17660);
nand U19562 (N_19562,N_18211,N_18625);
nor U19563 (N_19563,N_18698,N_18262);
nor U19564 (N_19564,N_18098,N_18446);
xor U19565 (N_19565,N_17820,N_18701);
xnor U19566 (N_19566,N_18606,N_17983);
nor U19567 (N_19567,N_17618,N_17540);
nor U19568 (N_19568,N_17731,N_18117);
and U19569 (N_19569,N_18327,N_17582);
xnor U19570 (N_19570,N_18086,N_17573);
nor U19571 (N_19571,N_18321,N_18457);
and U19572 (N_19572,N_18243,N_18238);
nand U19573 (N_19573,N_18237,N_18668);
nor U19574 (N_19574,N_18240,N_17583);
and U19575 (N_19575,N_18711,N_18023);
or U19576 (N_19576,N_17520,N_17682);
nor U19577 (N_19577,N_18081,N_17512);
xnor U19578 (N_19578,N_18272,N_17749);
xor U19579 (N_19579,N_18072,N_18356);
xor U19580 (N_19580,N_17949,N_18003);
xnor U19581 (N_19581,N_18475,N_17950);
and U19582 (N_19582,N_18005,N_17859);
nor U19583 (N_19583,N_18438,N_17840);
nor U19584 (N_19584,N_18543,N_18104);
xor U19585 (N_19585,N_17533,N_18000);
xnor U19586 (N_19586,N_18258,N_18530);
and U19587 (N_19587,N_17513,N_18429);
xor U19588 (N_19588,N_18458,N_17655);
nor U19589 (N_19589,N_18559,N_18430);
and U19590 (N_19590,N_18526,N_18345);
xor U19591 (N_19591,N_17593,N_17574);
or U19592 (N_19592,N_18264,N_18294);
nand U19593 (N_19593,N_17781,N_17536);
and U19594 (N_19594,N_17597,N_18206);
and U19595 (N_19595,N_18708,N_18526);
xor U19596 (N_19596,N_18522,N_18441);
nor U19597 (N_19597,N_17616,N_18666);
nand U19598 (N_19598,N_17585,N_17705);
and U19599 (N_19599,N_18034,N_17668);
or U19600 (N_19600,N_18357,N_18583);
nand U19601 (N_19601,N_18672,N_18516);
nor U19602 (N_19602,N_17937,N_17912);
nand U19603 (N_19603,N_17720,N_18171);
xor U19604 (N_19604,N_17757,N_17615);
and U19605 (N_19605,N_18401,N_17967);
xnor U19606 (N_19606,N_17510,N_17675);
nand U19607 (N_19607,N_17728,N_17631);
and U19608 (N_19608,N_18409,N_18679);
nor U19609 (N_19609,N_17602,N_18320);
and U19610 (N_19610,N_18125,N_17519);
or U19611 (N_19611,N_17961,N_17787);
nand U19612 (N_19612,N_18653,N_18285);
nor U19613 (N_19613,N_17942,N_18566);
and U19614 (N_19614,N_17559,N_18683);
xor U19615 (N_19615,N_17787,N_18045);
nor U19616 (N_19616,N_18445,N_18243);
nand U19617 (N_19617,N_18069,N_17970);
xor U19618 (N_19618,N_18234,N_18083);
nand U19619 (N_19619,N_18305,N_17923);
xor U19620 (N_19620,N_18437,N_18328);
or U19621 (N_19621,N_17905,N_18311);
nand U19622 (N_19622,N_17992,N_18654);
or U19623 (N_19623,N_18194,N_18186);
and U19624 (N_19624,N_18606,N_17786);
or U19625 (N_19625,N_18045,N_18256);
nand U19626 (N_19626,N_18512,N_18361);
nor U19627 (N_19627,N_17680,N_18294);
nand U19628 (N_19628,N_17539,N_17508);
or U19629 (N_19629,N_18091,N_18720);
xor U19630 (N_19630,N_18689,N_17519);
or U19631 (N_19631,N_18717,N_18234);
and U19632 (N_19632,N_18087,N_18586);
nand U19633 (N_19633,N_18444,N_18414);
xor U19634 (N_19634,N_17708,N_18556);
nor U19635 (N_19635,N_17972,N_17741);
nand U19636 (N_19636,N_18048,N_18535);
nor U19637 (N_19637,N_18673,N_17681);
nor U19638 (N_19638,N_18093,N_17839);
and U19639 (N_19639,N_18276,N_18004);
xnor U19640 (N_19640,N_18025,N_18458);
nand U19641 (N_19641,N_17585,N_18218);
nand U19642 (N_19642,N_18247,N_18531);
xnor U19643 (N_19643,N_18597,N_17693);
nor U19644 (N_19644,N_17658,N_17716);
xor U19645 (N_19645,N_17667,N_18718);
or U19646 (N_19646,N_18365,N_17524);
or U19647 (N_19647,N_18609,N_18676);
xor U19648 (N_19648,N_18180,N_18335);
or U19649 (N_19649,N_18574,N_18134);
and U19650 (N_19650,N_18071,N_17527);
or U19651 (N_19651,N_18623,N_17846);
xnor U19652 (N_19652,N_18156,N_17815);
nor U19653 (N_19653,N_17571,N_18614);
nand U19654 (N_19654,N_18566,N_18627);
and U19655 (N_19655,N_18725,N_17709);
or U19656 (N_19656,N_18591,N_18186);
nand U19657 (N_19657,N_18238,N_17950);
and U19658 (N_19658,N_18151,N_17875);
nand U19659 (N_19659,N_18561,N_17559);
and U19660 (N_19660,N_17818,N_18555);
nand U19661 (N_19661,N_17859,N_17544);
or U19662 (N_19662,N_17742,N_17804);
nor U19663 (N_19663,N_17680,N_18521);
xnor U19664 (N_19664,N_18268,N_17944);
nand U19665 (N_19665,N_18243,N_18194);
nor U19666 (N_19666,N_17575,N_17996);
and U19667 (N_19667,N_17596,N_17869);
or U19668 (N_19668,N_17550,N_17637);
xor U19669 (N_19669,N_17544,N_17784);
nor U19670 (N_19670,N_18026,N_18411);
and U19671 (N_19671,N_17723,N_18440);
or U19672 (N_19672,N_17923,N_17963);
nor U19673 (N_19673,N_18081,N_18129);
nand U19674 (N_19674,N_18278,N_17521);
and U19675 (N_19675,N_17671,N_17962);
nor U19676 (N_19676,N_17666,N_18257);
or U19677 (N_19677,N_18225,N_17510);
or U19678 (N_19678,N_17945,N_17702);
or U19679 (N_19679,N_18437,N_17871);
and U19680 (N_19680,N_18306,N_18328);
nor U19681 (N_19681,N_18556,N_17574);
xor U19682 (N_19682,N_17644,N_18609);
nor U19683 (N_19683,N_18158,N_18286);
nor U19684 (N_19684,N_18726,N_17884);
and U19685 (N_19685,N_17749,N_18331);
xor U19686 (N_19686,N_18088,N_18646);
nor U19687 (N_19687,N_18275,N_18378);
xor U19688 (N_19688,N_18165,N_17555);
nand U19689 (N_19689,N_18324,N_18647);
nor U19690 (N_19690,N_17889,N_17965);
or U19691 (N_19691,N_18633,N_18611);
nand U19692 (N_19692,N_18173,N_18224);
nor U19693 (N_19693,N_17569,N_18545);
or U19694 (N_19694,N_18747,N_18145);
nor U19695 (N_19695,N_18399,N_18710);
nand U19696 (N_19696,N_18014,N_18467);
or U19697 (N_19697,N_17622,N_18462);
xor U19698 (N_19698,N_18074,N_17926);
or U19699 (N_19699,N_18544,N_18612);
nor U19700 (N_19700,N_18706,N_18418);
and U19701 (N_19701,N_18301,N_18088);
and U19702 (N_19702,N_17976,N_18057);
nand U19703 (N_19703,N_17982,N_17877);
and U19704 (N_19704,N_17545,N_18124);
or U19705 (N_19705,N_18188,N_17710);
nand U19706 (N_19706,N_17787,N_17594);
or U19707 (N_19707,N_17819,N_18161);
xor U19708 (N_19708,N_17638,N_17674);
nand U19709 (N_19709,N_17522,N_18638);
nor U19710 (N_19710,N_18225,N_18197);
or U19711 (N_19711,N_18107,N_18023);
nor U19712 (N_19712,N_18380,N_18421);
nor U19713 (N_19713,N_17983,N_17634);
nand U19714 (N_19714,N_18211,N_17875);
nand U19715 (N_19715,N_18321,N_17969);
nor U19716 (N_19716,N_18743,N_17680);
and U19717 (N_19717,N_17867,N_18473);
nor U19718 (N_19718,N_18679,N_17612);
and U19719 (N_19719,N_17790,N_18039);
nand U19720 (N_19720,N_17928,N_18327);
nor U19721 (N_19721,N_18044,N_18200);
and U19722 (N_19722,N_18569,N_18728);
xnor U19723 (N_19723,N_17850,N_18349);
and U19724 (N_19724,N_17810,N_18178);
or U19725 (N_19725,N_17740,N_18665);
nor U19726 (N_19726,N_17822,N_18156);
nor U19727 (N_19727,N_18594,N_18387);
or U19728 (N_19728,N_17846,N_17505);
nor U19729 (N_19729,N_18326,N_17590);
xor U19730 (N_19730,N_17558,N_17755);
and U19731 (N_19731,N_17961,N_17890);
and U19732 (N_19732,N_17856,N_18402);
nand U19733 (N_19733,N_18597,N_18344);
nor U19734 (N_19734,N_18335,N_18117);
nor U19735 (N_19735,N_18286,N_18538);
and U19736 (N_19736,N_17766,N_17737);
or U19737 (N_19737,N_18057,N_18254);
nand U19738 (N_19738,N_17685,N_18127);
or U19739 (N_19739,N_17998,N_18209);
nor U19740 (N_19740,N_17962,N_17522);
or U19741 (N_19741,N_17961,N_18167);
nand U19742 (N_19742,N_17846,N_18374);
or U19743 (N_19743,N_18407,N_17996);
nand U19744 (N_19744,N_17934,N_18442);
xnor U19745 (N_19745,N_18248,N_17682);
or U19746 (N_19746,N_18217,N_18667);
xor U19747 (N_19747,N_18255,N_18698);
xnor U19748 (N_19748,N_18036,N_18265);
and U19749 (N_19749,N_17924,N_18376);
nand U19750 (N_19750,N_18408,N_18503);
xnor U19751 (N_19751,N_18595,N_17747);
nor U19752 (N_19752,N_18104,N_17613);
nand U19753 (N_19753,N_18165,N_18241);
nand U19754 (N_19754,N_18095,N_18536);
or U19755 (N_19755,N_18672,N_17514);
nand U19756 (N_19756,N_17573,N_18088);
nor U19757 (N_19757,N_17926,N_18076);
and U19758 (N_19758,N_18200,N_17566);
xor U19759 (N_19759,N_18365,N_17539);
and U19760 (N_19760,N_17532,N_18366);
and U19761 (N_19761,N_18044,N_17534);
or U19762 (N_19762,N_18250,N_18445);
nand U19763 (N_19763,N_17571,N_17983);
nor U19764 (N_19764,N_18508,N_17541);
and U19765 (N_19765,N_17573,N_18369);
xnor U19766 (N_19766,N_17894,N_17581);
nand U19767 (N_19767,N_17955,N_18343);
and U19768 (N_19768,N_18198,N_18357);
nand U19769 (N_19769,N_18173,N_17575);
and U19770 (N_19770,N_18132,N_17618);
nand U19771 (N_19771,N_17957,N_17942);
xnor U19772 (N_19772,N_17679,N_17781);
xor U19773 (N_19773,N_18078,N_18261);
nand U19774 (N_19774,N_17778,N_18453);
or U19775 (N_19775,N_17506,N_18306);
or U19776 (N_19776,N_18016,N_17852);
nor U19777 (N_19777,N_17973,N_17813);
or U19778 (N_19778,N_18559,N_18148);
and U19779 (N_19779,N_17958,N_17913);
nand U19780 (N_19780,N_18075,N_18274);
and U19781 (N_19781,N_18394,N_18471);
and U19782 (N_19782,N_18432,N_18138);
nor U19783 (N_19783,N_18637,N_17503);
xor U19784 (N_19784,N_17838,N_18332);
xor U19785 (N_19785,N_17949,N_17959);
nand U19786 (N_19786,N_18229,N_17762);
or U19787 (N_19787,N_18182,N_17523);
xnor U19788 (N_19788,N_18663,N_17765);
xor U19789 (N_19789,N_17840,N_18517);
or U19790 (N_19790,N_18207,N_17543);
nor U19791 (N_19791,N_17774,N_18539);
and U19792 (N_19792,N_17535,N_18200);
xnor U19793 (N_19793,N_18703,N_18739);
or U19794 (N_19794,N_18148,N_18011);
or U19795 (N_19795,N_18156,N_17588);
xnor U19796 (N_19796,N_17948,N_18099);
or U19797 (N_19797,N_17946,N_18442);
xor U19798 (N_19798,N_18582,N_17681);
nand U19799 (N_19799,N_17934,N_17771);
nand U19800 (N_19800,N_18025,N_17991);
nand U19801 (N_19801,N_17558,N_18421);
nor U19802 (N_19802,N_18303,N_18492);
nor U19803 (N_19803,N_17782,N_18645);
or U19804 (N_19804,N_17912,N_17929);
or U19805 (N_19805,N_17912,N_18173);
xnor U19806 (N_19806,N_17854,N_17586);
nand U19807 (N_19807,N_17693,N_17844);
or U19808 (N_19808,N_18613,N_17573);
nand U19809 (N_19809,N_17888,N_17522);
nand U19810 (N_19810,N_18645,N_18251);
or U19811 (N_19811,N_18568,N_18740);
and U19812 (N_19812,N_17675,N_17724);
or U19813 (N_19813,N_17758,N_17565);
xor U19814 (N_19814,N_18340,N_17600);
nand U19815 (N_19815,N_17871,N_18352);
or U19816 (N_19816,N_18046,N_18137);
nand U19817 (N_19817,N_18557,N_17859);
xor U19818 (N_19818,N_17755,N_17869);
nor U19819 (N_19819,N_18582,N_18290);
nor U19820 (N_19820,N_18453,N_18314);
and U19821 (N_19821,N_18467,N_18096);
or U19822 (N_19822,N_17582,N_18040);
xnor U19823 (N_19823,N_18487,N_18233);
nand U19824 (N_19824,N_18604,N_17785);
xor U19825 (N_19825,N_17788,N_18544);
and U19826 (N_19826,N_18144,N_18697);
nor U19827 (N_19827,N_18571,N_18666);
nand U19828 (N_19828,N_18670,N_17945);
and U19829 (N_19829,N_18156,N_17869);
or U19830 (N_19830,N_18666,N_18720);
and U19831 (N_19831,N_18104,N_18156);
and U19832 (N_19832,N_17727,N_18527);
xnor U19833 (N_19833,N_18327,N_18145);
xor U19834 (N_19834,N_18210,N_18532);
nor U19835 (N_19835,N_17601,N_18350);
nand U19836 (N_19836,N_17905,N_17797);
nor U19837 (N_19837,N_17966,N_17601);
or U19838 (N_19838,N_17547,N_17512);
xor U19839 (N_19839,N_18410,N_18515);
nor U19840 (N_19840,N_18611,N_18717);
and U19841 (N_19841,N_17691,N_18387);
nand U19842 (N_19842,N_17613,N_17647);
xor U19843 (N_19843,N_18038,N_17567);
nand U19844 (N_19844,N_17557,N_18237);
nor U19845 (N_19845,N_18377,N_17561);
or U19846 (N_19846,N_18010,N_18556);
and U19847 (N_19847,N_17679,N_18318);
or U19848 (N_19848,N_18257,N_17730);
nand U19849 (N_19849,N_18008,N_18377);
and U19850 (N_19850,N_18257,N_18358);
or U19851 (N_19851,N_18470,N_18519);
nand U19852 (N_19852,N_18744,N_18322);
xor U19853 (N_19853,N_17737,N_17921);
and U19854 (N_19854,N_18052,N_18032);
xor U19855 (N_19855,N_17634,N_18721);
nor U19856 (N_19856,N_18721,N_18073);
xor U19857 (N_19857,N_18276,N_18484);
nand U19858 (N_19858,N_18460,N_18711);
xnor U19859 (N_19859,N_17855,N_18097);
xor U19860 (N_19860,N_17666,N_17878);
xor U19861 (N_19861,N_18450,N_18391);
nor U19862 (N_19862,N_18263,N_17627);
nor U19863 (N_19863,N_17733,N_17797);
xnor U19864 (N_19864,N_17669,N_17827);
or U19865 (N_19865,N_18068,N_17713);
nand U19866 (N_19866,N_17817,N_18305);
or U19867 (N_19867,N_18584,N_17957);
nand U19868 (N_19868,N_18285,N_18445);
xnor U19869 (N_19869,N_17623,N_18522);
nand U19870 (N_19870,N_17611,N_17793);
xnor U19871 (N_19871,N_18408,N_17908);
or U19872 (N_19872,N_17509,N_18420);
and U19873 (N_19873,N_18020,N_17996);
and U19874 (N_19874,N_18611,N_18576);
and U19875 (N_19875,N_17949,N_18702);
nand U19876 (N_19876,N_17631,N_18007);
and U19877 (N_19877,N_18037,N_17939);
nor U19878 (N_19878,N_18222,N_18629);
and U19879 (N_19879,N_17830,N_18581);
nor U19880 (N_19880,N_17787,N_18369);
xnor U19881 (N_19881,N_18083,N_17980);
nor U19882 (N_19882,N_18347,N_18307);
xnor U19883 (N_19883,N_17611,N_17522);
and U19884 (N_19884,N_18364,N_18286);
xor U19885 (N_19885,N_18556,N_17680);
xnor U19886 (N_19886,N_17841,N_18322);
and U19887 (N_19887,N_17733,N_17522);
nor U19888 (N_19888,N_17578,N_17640);
and U19889 (N_19889,N_18408,N_18166);
nor U19890 (N_19890,N_17912,N_18580);
xnor U19891 (N_19891,N_17998,N_18404);
and U19892 (N_19892,N_18500,N_18278);
and U19893 (N_19893,N_17679,N_18231);
xor U19894 (N_19894,N_18014,N_18401);
nand U19895 (N_19895,N_18476,N_18568);
nand U19896 (N_19896,N_18266,N_18515);
or U19897 (N_19897,N_18740,N_17746);
or U19898 (N_19898,N_17688,N_18311);
and U19899 (N_19899,N_17856,N_18282);
and U19900 (N_19900,N_17695,N_18151);
xor U19901 (N_19901,N_18380,N_18257);
or U19902 (N_19902,N_18182,N_18192);
nand U19903 (N_19903,N_18194,N_18209);
and U19904 (N_19904,N_18706,N_18332);
and U19905 (N_19905,N_17969,N_18666);
xnor U19906 (N_19906,N_17590,N_18677);
xnor U19907 (N_19907,N_18262,N_18358);
nand U19908 (N_19908,N_18719,N_18349);
nor U19909 (N_19909,N_18068,N_17829);
or U19910 (N_19910,N_17679,N_18572);
nor U19911 (N_19911,N_17640,N_17913);
nand U19912 (N_19912,N_18037,N_18544);
nand U19913 (N_19913,N_18565,N_18384);
or U19914 (N_19914,N_18361,N_18661);
and U19915 (N_19915,N_17917,N_18302);
or U19916 (N_19916,N_18220,N_18135);
nand U19917 (N_19917,N_18566,N_17588);
and U19918 (N_19918,N_18679,N_18083);
xnor U19919 (N_19919,N_18553,N_18085);
and U19920 (N_19920,N_18032,N_17988);
nand U19921 (N_19921,N_18579,N_18217);
nand U19922 (N_19922,N_17632,N_18284);
xor U19923 (N_19923,N_18330,N_17919);
nand U19924 (N_19924,N_18430,N_17549);
nand U19925 (N_19925,N_18213,N_18108);
nand U19926 (N_19926,N_18013,N_18719);
xnor U19927 (N_19927,N_17782,N_18393);
xor U19928 (N_19928,N_17995,N_17620);
and U19929 (N_19929,N_18224,N_17568);
and U19930 (N_19930,N_17508,N_18434);
and U19931 (N_19931,N_17564,N_18026);
and U19932 (N_19932,N_17626,N_17918);
nor U19933 (N_19933,N_17904,N_17705);
xnor U19934 (N_19934,N_18498,N_18440);
nand U19935 (N_19935,N_18551,N_18306);
and U19936 (N_19936,N_17595,N_18124);
xor U19937 (N_19937,N_18568,N_18342);
nand U19938 (N_19938,N_17918,N_17600);
and U19939 (N_19939,N_17609,N_17733);
and U19940 (N_19940,N_18494,N_17866);
and U19941 (N_19941,N_18577,N_17543);
or U19942 (N_19942,N_18303,N_18009);
xor U19943 (N_19943,N_17506,N_18235);
and U19944 (N_19944,N_17846,N_18093);
xnor U19945 (N_19945,N_17651,N_18388);
nand U19946 (N_19946,N_18618,N_18122);
and U19947 (N_19947,N_17963,N_18516);
and U19948 (N_19948,N_17593,N_18583);
or U19949 (N_19949,N_17902,N_18565);
nand U19950 (N_19950,N_18263,N_18124);
nand U19951 (N_19951,N_17625,N_18072);
and U19952 (N_19952,N_18628,N_18494);
or U19953 (N_19953,N_18381,N_17910);
or U19954 (N_19954,N_18254,N_18650);
nand U19955 (N_19955,N_18053,N_18670);
and U19956 (N_19956,N_18413,N_17515);
nand U19957 (N_19957,N_18747,N_18228);
nor U19958 (N_19958,N_17957,N_18391);
or U19959 (N_19959,N_17756,N_18728);
nand U19960 (N_19960,N_18476,N_17814);
or U19961 (N_19961,N_18315,N_17992);
nor U19962 (N_19962,N_18087,N_18001);
nor U19963 (N_19963,N_18649,N_18701);
or U19964 (N_19964,N_18068,N_18540);
xnor U19965 (N_19965,N_17900,N_17925);
xnor U19966 (N_19966,N_17527,N_18558);
xor U19967 (N_19967,N_18671,N_17726);
and U19968 (N_19968,N_17807,N_17557);
nand U19969 (N_19969,N_17620,N_18368);
nand U19970 (N_19970,N_18312,N_17524);
xor U19971 (N_19971,N_18500,N_18336);
nand U19972 (N_19972,N_18383,N_17762);
nor U19973 (N_19973,N_18198,N_18469);
nor U19974 (N_19974,N_18440,N_18136);
and U19975 (N_19975,N_18022,N_17567);
xor U19976 (N_19976,N_17521,N_17868);
xor U19977 (N_19977,N_17517,N_17657);
xor U19978 (N_19978,N_18683,N_18286);
and U19979 (N_19979,N_18610,N_18341);
xor U19980 (N_19980,N_17674,N_18676);
xor U19981 (N_19981,N_18313,N_18531);
nor U19982 (N_19982,N_18455,N_18418);
nand U19983 (N_19983,N_17704,N_18085);
nand U19984 (N_19984,N_17608,N_18624);
or U19985 (N_19985,N_17797,N_18495);
nor U19986 (N_19986,N_17761,N_18168);
nand U19987 (N_19987,N_18417,N_17649);
nand U19988 (N_19988,N_18598,N_17832);
xor U19989 (N_19989,N_18336,N_18014);
or U19990 (N_19990,N_17711,N_18067);
and U19991 (N_19991,N_18091,N_18337);
nor U19992 (N_19992,N_18467,N_18363);
or U19993 (N_19993,N_18490,N_17502);
xor U19994 (N_19994,N_18507,N_17917);
xnor U19995 (N_19995,N_17576,N_17893);
xnor U19996 (N_19996,N_18554,N_18416);
and U19997 (N_19997,N_18123,N_17563);
and U19998 (N_19998,N_18610,N_17759);
or U19999 (N_19999,N_17876,N_18501);
nand U20000 (N_20000,N_19052,N_19593);
nand U20001 (N_20001,N_19071,N_18900);
xor U20002 (N_20002,N_19365,N_19711);
nand U20003 (N_20003,N_19179,N_19286);
and U20004 (N_20004,N_19131,N_19962);
or U20005 (N_20005,N_19579,N_19808);
nor U20006 (N_20006,N_19033,N_19200);
nand U20007 (N_20007,N_19148,N_18753);
nand U20008 (N_20008,N_19235,N_19223);
nand U20009 (N_20009,N_19011,N_19116);
and U20010 (N_20010,N_19768,N_19991);
and U20011 (N_20011,N_18862,N_19161);
xnor U20012 (N_20012,N_19344,N_19598);
nor U20013 (N_20013,N_19631,N_19078);
or U20014 (N_20014,N_19121,N_18899);
or U20015 (N_20015,N_19426,N_19325);
xnor U20016 (N_20016,N_18907,N_18870);
xnor U20017 (N_20017,N_19602,N_19554);
and U20018 (N_20018,N_19105,N_19907);
or U20019 (N_20019,N_19735,N_19329);
or U20020 (N_20020,N_19122,N_19158);
or U20021 (N_20021,N_18782,N_19425);
or U20022 (N_20022,N_19212,N_19386);
or U20023 (N_20023,N_19516,N_19569);
and U20024 (N_20024,N_19731,N_19846);
or U20025 (N_20025,N_19421,N_19450);
nand U20026 (N_20026,N_19701,N_19043);
and U20027 (N_20027,N_19199,N_19376);
nor U20028 (N_20028,N_19065,N_19869);
nand U20029 (N_20029,N_19526,N_19612);
and U20030 (N_20030,N_18866,N_19480);
nor U20031 (N_20031,N_19015,N_18985);
nand U20032 (N_20032,N_18794,N_19936);
and U20033 (N_20033,N_18976,N_19639);
nand U20034 (N_20034,N_19081,N_19141);
nor U20035 (N_20035,N_18755,N_19397);
xor U20036 (N_20036,N_19427,N_19156);
nand U20037 (N_20037,N_19816,N_19620);
xor U20038 (N_20038,N_19658,N_18958);
nor U20039 (N_20039,N_19959,N_19811);
nor U20040 (N_20040,N_19479,N_19844);
nor U20041 (N_20041,N_18903,N_18892);
nand U20042 (N_20042,N_19398,N_19993);
xnor U20043 (N_20043,N_19171,N_18799);
nor U20044 (N_20044,N_19556,N_18959);
nor U20045 (N_20045,N_19027,N_19572);
or U20046 (N_20046,N_19010,N_19515);
xnor U20047 (N_20047,N_18857,N_19412);
nand U20048 (N_20048,N_19168,N_19111);
nor U20049 (N_20049,N_19989,N_19749);
xnor U20050 (N_20050,N_18843,N_18830);
and U20051 (N_20051,N_19361,N_18928);
or U20052 (N_20052,N_19674,N_19039);
and U20053 (N_20053,N_19667,N_19162);
and U20054 (N_20054,N_18954,N_19410);
nor U20055 (N_20055,N_19341,N_19436);
or U20056 (N_20056,N_19944,N_19401);
and U20057 (N_20057,N_18908,N_19964);
and U20058 (N_20058,N_18804,N_19560);
nand U20059 (N_20059,N_19134,N_19834);
and U20060 (N_20060,N_18953,N_19879);
nand U20061 (N_20061,N_19822,N_19885);
nor U20062 (N_20062,N_19153,N_19193);
nor U20063 (N_20063,N_19483,N_19845);
nand U20064 (N_20064,N_18921,N_19002);
and U20065 (N_20065,N_19752,N_19177);
nand U20066 (N_20066,N_19130,N_19695);
or U20067 (N_20067,N_19222,N_19088);
nand U20068 (N_20068,N_19032,N_19167);
and U20069 (N_20069,N_19256,N_19857);
nand U20070 (N_20070,N_19584,N_19404);
nor U20071 (N_20071,N_18896,N_19666);
or U20072 (N_20072,N_19353,N_19040);
or U20073 (N_20073,N_19917,N_19294);
xnor U20074 (N_20074,N_19688,N_19003);
or U20075 (N_20075,N_19916,N_18820);
or U20076 (N_20076,N_18826,N_19050);
nor U20077 (N_20077,N_19431,N_19679);
nor U20078 (N_20078,N_18929,N_18860);
or U20079 (N_20079,N_19607,N_19102);
and U20080 (N_20080,N_18955,N_19465);
and U20081 (N_20081,N_19823,N_19971);
xnor U20082 (N_20082,N_19859,N_18802);
nor U20083 (N_20083,N_18837,N_19313);
xor U20084 (N_20084,N_18939,N_19248);
and U20085 (N_20085,N_19301,N_19580);
nor U20086 (N_20086,N_18932,N_19908);
xnor U20087 (N_20087,N_19403,N_19255);
or U20088 (N_20088,N_19918,N_19746);
or U20089 (N_20089,N_19977,N_19541);
xnor U20090 (N_20090,N_18865,N_18834);
and U20091 (N_20091,N_19831,N_19174);
nand U20092 (N_20092,N_18871,N_18919);
nand U20093 (N_20093,N_19447,N_19750);
or U20094 (N_20094,N_19107,N_19778);
xnor U20095 (N_20095,N_19542,N_19502);
or U20096 (N_20096,N_19644,N_19910);
or U20097 (N_20097,N_19262,N_19187);
or U20098 (N_20098,N_19439,N_19098);
or U20099 (N_20099,N_19266,N_18788);
nand U20100 (N_20100,N_19460,N_19949);
nor U20101 (N_20101,N_19986,N_19407);
and U20102 (N_20102,N_19546,N_18855);
xnor U20103 (N_20103,N_19522,N_19478);
or U20104 (N_20104,N_19570,N_19780);
nor U20105 (N_20105,N_19549,N_19417);
xor U20106 (N_20106,N_19958,N_19020);
and U20107 (N_20107,N_19799,N_19180);
nor U20108 (N_20108,N_18867,N_19792);
or U20109 (N_20109,N_19878,N_19905);
and U20110 (N_20110,N_19416,N_18801);
and U20111 (N_20111,N_18877,N_19609);
nand U20112 (N_20112,N_19617,N_19893);
nand U20113 (N_20113,N_18938,N_18996);
xnor U20114 (N_20114,N_19477,N_19770);
and U20115 (N_20115,N_19796,N_19506);
nor U20116 (N_20116,N_19942,N_19614);
or U20117 (N_20117,N_19793,N_19628);
nand U20118 (N_20118,N_19079,N_19345);
and U20119 (N_20119,N_19095,N_19021);
or U20120 (N_20120,N_19292,N_18845);
nor U20121 (N_20121,N_18930,N_19448);
nand U20122 (N_20122,N_19623,N_19348);
and U20123 (N_20123,N_19832,N_19568);
or U20124 (N_20124,N_19629,N_19956);
and U20125 (N_20125,N_19794,N_18809);
nand U20126 (N_20126,N_19661,N_18993);
or U20127 (N_20127,N_19764,N_19928);
xnor U20128 (N_20128,N_18918,N_19709);
nor U20129 (N_20129,N_18934,N_19565);
nand U20130 (N_20130,N_19836,N_19847);
or U20131 (N_20131,N_18814,N_19449);
nand U20132 (N_20132,N_19160,N_19152);
nor U20133 (N_20133,N_19428,N_19108);
nand U20134 (N_20134,N_19529,N_19521);
and U20135 (N_20135,N_19599,N_18817);
xnor U20136 (N_20136,N_19797,N_19343);
nor U20137 (N_20137,N_19535,N_18940);
nand U20138 (N_20138,N_19539,N_19247);
or U20139 (N_20139,N_18758,N_19992);
nand U20140 (N_20140,N_19585,N_19897);
and U20141 (N_20141,N_19728,N_18931);
nor U20142 (N_20142,N_18835,N_19354);
and U20143 (N_20143,N_19024,N_18780);
and U20144 (N_20144,N_19699,N_19402);
and U20145 (N_20145,N_19821,N_19547);
xnor U20146 (N_20146,N_18840,N_19475);
xnor U20147 (N_20147,N_19967,N_19356);
and U20148 (N_20148,N_19605,N_19297);
nor U20149 (N_20149,N_19594,N_19181);
and U20150 (N_20150,N_19227,N_19038);
or U20151 (N_20151,N_19323,N_19707);
nand U20152 (N_20152,N_19611,N_18765);
and U20153 (N_20153,N_19007,N_19000);
and U20154 (N_20154,N_19637,N_19236);
and U20155 (N_20155,N_18973,N_19938);
xnor U20156 (N_20156,N_19159,N_19385);
xnor U20157 (N_20157,N_19525,N_18838);
nand U20158 (N_20158,N_19660,N_18991);
nand U20159 (N_20159,N_19948,N_19429);
and U20160 (N_20160,N_19953,N_19865);
nor U20161 (N_20161,N_19034,N_18989);
nor U20162 (N_20162,N_19716,N_18988);
nor U20163 (N_20163,N_19259,N_18791);
and U20164 (N_20164,N_19012,N_19538);
and U20165 (N_20165,N_19087,N_18997);
xor U20166 (N_20166,N_18948,N_19360);
nand U20167 (N_20167,N_18910,N_19451);
or U20168 (N_20168,N_19459,N_19984);
xor U20169 (N_20169,N_19619,N_19067);
and U20170 (N_20170,N_18844,N_18884);
or U20171 (N_20171,N_19837,N_19642);
xnor U20172 (N_20172,N_19053,N_18785);
xnor U20173 (N_20173,N_18767,N_19391);
and U20174 (N_20174,N_19943,N_19302);
or U20175 (N_20175,N_19476,N_19718);
nand U20176 (N_20176,N_19678,N_18813);
xnor U20177 (N_20177,N_19800,N_19801);
or U20178 (N_20178,N_19120,N_19265);
xnor U20179 (N_20179,N_19492,N_19693);
nor U20180 (N_20180,N_19576,N_19604);
nor U20181 (N_20181,N_19420,N_19858);
and U20182 (N_20182,N_19671,N_19315);
nor U20183 (N_20183,N_19934,N_19906);
xor U20184 (N_20184,N_19810,N_18912);
and U20185 (N_20185,N_19049,N_19328);
or U20186 (N_20186,N_19241,N_18972);
xor U20187 (N_20187,N_19068,N_19504);
nand U20188 (N_20188,N_18781,N_19980);
or U20189 (N_20189,N_19616,N_19875);
nand U20190 (N_20190,N_18949,N_19951);
nor U20191 (N_20191,N_19717,N_19567);
and U20192 (N_20192,N_19370,N_19820);
and U20193 (N_20193,N_19226,N_19714);
nand U20194 (N_20194,N_19291,N_19443);
or U20195 (N_20195,N_19895,N_19221);
xor U20196 (N_20196,N_18797,N_19840);
nor U20197 (N_20197,N_18787,N_19473);
and U20198 (N_20198,N_19287,N_19855);
or U20199 (N_20199,N_19048,N_19037);
nand U20200 (N_20200,N_18822,N_19972);
or U20201 (N_20201,N_19110,N_19084);
or U20202 (N_20202,N_19862,N_19779);
xor U20203 (N_20203,N_19016,N_19947);
and U20204 (N_20204,N_19999,N_19785);
nor U20205 (N_20205,N_18878,N_19471);
and U20206 (N_20206,N_19649,N_18823);
and U20207 (N_20207,N_19901,N_19374);
nor U20208 (N_20208,N_19829,N_19231);
nand U20209 (N_20209,N_19096,N_19381);
or U20210 (N_20210,N_19753,N_19319);
xnor U20211 (N_20211,N_19497,N_19268);
xnor U20212 (N_20212,N_19462,N_19830);
nor U20213 (N_20213,N_19932,N_19507);
nand U20214 (N_20214,N_19807,N_19969);
xnor U20215 (N_20215,N_19782,N_19633);
nand U20216 (N_20216,N_19940,N_19795);
or U20217 (N_20217,N_18764,N_19998);
nand U20218 (N_20218,N_19237,N_19101);
or U20219 (N_20219,N_19184,N_19406);
or U20220 (N_20220,N_19210,N_19994);
and U20221 (N_20221,N_18978,N_18786);
nand U20222 (N_20222,N_19233,N_19091);
nor U20223 (N_20223,N_19201,N_19727);
xnor U20224 (N_20224,N_19288,N_19380);
or U20225 (N_20225,N_19145,N_18987);
and U20226 (N_20226,N_19191,N_19045);
nor U20227 (N_20227,N_19518,N_19474);
xor U20228 (N_20228,N_19511,N_19119);
nor U20229 (N_20229,N_19335,N_19149);
xor U20230 (N_20230,N_19044,N_19009);
xor U20231 (N_20231,N_19132,N_19279);
nand U20232 (N_20232,N_19788,N_19269);
nor U20233 (N_20233,N_19890,N_18982);
nor U20234 (N_20234,N_19139,N_19115);
or U20235 (N_20235,N_19982,N_19787);
and U20236 (N_20236,N_19653,N_19305);
nand U20237 (N_20237,N_19519,N_19896);
xnor U20238 (N_20238,N_19157,N_19899);
or U20239 (N_20239,N_19379,N_18915);
nand U20240 (N_20240,N_19851,N_19528);
or U20241 (N_20241,N_18942,N_19777);
or U20242 (N_20242,N_19610,N_19500);
nor U20243 (N_20243,N_19996,N_19640);
nand U20244 (N_20244,N_19981,N_19164);
nor U20245 (N_20245,N_19469,N_19643);
nor U20246 (N_20246,N_19337,N_18760);
or U20247 (N_20247,N_19880,N_19888);
and U20248 (N_20248,N_19596,N_19487);
nand U20249 (N_20249,N_18812,N_19806);
nor U20250 (N_20250,N_18754,N_19347);
xor U20251 (N_20251,N_19662,N_19929);
or U20252 (N_20252,N_19244,N_19987);
and U20253 (N_20253,N_19850,N_18916);
nor U20254 (N_20254,N_18775,N_19627);
xor U20255 (N_20255,N_19466,N_19970);
nand U20256 (N_20256,N_18895,N_19083);
and U20257 (N_20257,N_18776,N_19383);
and U20258 (N_20258,N_19817,N_19220);
nand U20259 (N_20259,N_19126,N_19544);
nand U20260 (N_20260,N_19721,N_19127);
xor U20261 (N_20261,N_19188,N_19290);
and U20262 (N_20262,N_19868,N_19508);
nor U20263 (N_20263,N_19697,N_19713);
and U20264 (N_20264,N_19352,N_19151);
nor U20265 (N_20265,N_19976,N_19809);
xnor U20266 (N_20266,N_18861,N_19411);
or U20267 (N_20267,N_19505,N_19077);
or U20268 (N_20268,N_19258,N_19140);
and U20269 (N_20269,N_19514,N_19481);
nand U20270 (N_20270,N_19902,N_18879);
nor U20271 (N_20271,N_19317,N_19655);
xor U20272 (N_20272,N_18992,N_19968);
nor U20273 (N_20273,N_19589,N_19756);
nand U20274 (N_20274,N_19990,N_19424);
and U20275 (N_20275,N_19251,N_19591);
nand U20276 (N_20276,N_19457,N_19245);
or U20277 (N_20277,N_19493,N_19112);
or U20278 (N_20278,N_18924,N_19574);
or U20279 (N_20279,N_19921,N_18827);
nand U20280 (N_20280,N_19732,N_19853);
and U20281 (N_20281,N_19334,N_18890);
nand U20282 (N_20282,N_19710,N_19664);
xor U20283 (N_20283,N_19937,N_19960);
nor U20284 (N_20284,N_18925,N_19252);
xnor U20285 (N_20285,N_19138,N_19326);
and U20286 (N_20286,N_19961,N_19647);
nand U20287 (N_20287,N_19283,N_19057);
xnor U20288 (N_20288,N_18815,N_19239);
nor U20289 (N_20289,N_19856,N_18829);
and U20290 (N_20290,N_19310,N_19510);
or U20291 (N_20291,N_19914,N_18913);
or U20292 (N_20292,N_19240,N_19747);
nand U20293 (N_20293,N_19866,N_19503);
or U20294 (N_20294,N_19419,N_18839);
or U20295 (N_20295,N_19613,N_19042);
or U20296 (N_20296,N_19757,N_18808);
or U20297 (N_20297,N_18874,N_19440);
or U20298 (N_20298,N_19299,N_19592);
and U20299 (N_20299,N_19769,N_19881);
and U20300 (N_20300,N_18796,N_19722);
xor U20301 (N_20301,N_19074,N_19657);
xor U20302 (N_20302,N_19069,N_19267);
and U20303 (N_20303,N_19675,N_18784);
nor U20304 (N_20304,N_19690,N_19531);
or U20305 (N_20305,N_19553,N_18885);
xnor U20306 (N_20306,N_19520,N_19578);
xor U20307 (N_20307,N_19638,N_19295);
nand U20308 (N_20308,N_18811,N_19304);
nor U20309 (N_20309,N_18847,N_19147);
or U20310 (N_20310,N_19509,N_19125);
or U20311 (N_20311,N_18898,N_18995);
and U20312 (N_20312,N_19673,N_19312);
nor U20313 (N_20313,N_19733,N_19490);
nor U20314 (N_20314,N_19280,N_19729);
and U20315 (N_20315,N_19804,N_18828);
nand U20316 (N_20316,N_18963,N_18886);
and U20317 (N_20317,N_19708,N_19861);
xor U20318 (N_20318,N_19997,N_19583);
xor U20319 (N_20319,N_18858,N_19186);
and U20320 (N_20320,N_19367,N_19550);
xnor U20321 (N_20321,N_19155,N_18759);
nor U20322 (N_20322,N_18752,N_18937);
nand U20323 (N_20323,N_19561,N_19775);
xor U20324 (N_20324,N_19004,N_19537);
xor U20325 (N_20325,N_19877,N_19296);
xor U20326 (N_20326,N_19672,N_18970);
or U20327 (N_20327,N_19357,N_19724);
nand U20328 (N_20328,N_19072,N_19029);
nand U20329 (N_20329,N_19144,N_19172);
xor U20330 (N_20330,N_19333,N_19389);
nand U20331 (N_20331,N_19204,N_18831);
or U20332 (N_20332,N_18933,N_19253);
or U20333 (N_20333,N_19827,N_19046);
or U20334 (N_20334,N_19587,N_18936);
xor U20335 (N_20335,N_19725,N_18783);
xnor U20336 (N_20336,N_19985,N_19659);
or U20337 (N_20337,N_19499,N_18944);
xnor U20338 (N_20338,N_19826,N_19080);
nor U20339 (N_20339,N_19945,N_19109);
nand U20340 (N_20340,N_19931,N_19498);
and U20341 (N_20341,N_19636,N_18841);
xor U20342 (N_20342,N_19812,N_19263);
and U20343 (N_20343,N_19852,N_19285);
nor U20344 (N_20344,N_19470,N_18984);
xnor U20345 (N_20345,N_18872,N_19742);
nor U20346 (N_20346,N_18810,N_19308);
nand U20347 (N_20347,N_19104,N_19698);
or U20348 (N_20348,N_18751,N_19264);
or U20349 (N_20349,N_19645,N_19198);
xnor U20350 (N_20350,N_19791,N_19372);
or U20351 (N_20351,N_18961,N_19501);
nand U20352 (N_20352,N_19332,N_18920);
nand U20353 (N_20353,N_19117,N_19324);
nor U20354 (N_20354,N_19097,N_19755);
nor U20355 (N_20355,N_19339,N_18941);
xor U20356 (N_20356,N_19789,N_19496);
xnor U20357 (N_20357,N_18893,N_19702);
nor U20358 (N_20358,N_19113,N_19835);
xor U20359 (N_20359,N_19512,N_19955);
nand U20360 (N_20360,N_19103,N_19135);
nand U20361 (N_20361,N_18816,N_19618);
nor U20362 (N_20362,N_19208,N_19963);
xnor U20363 (N_20363,N_19723,N_18935);
nand U20364 (N_20364,N_19281,N_19663);
nor U20365 (N_20365,N_19382,N_19368);
and U20366 (N_20366,N_19058,N_18901);
nand U20367 (N_20367,N_19446,N_19726);
nand U20368 (N_20368,N_19458,N_19524);
and U20369 (N_20369,N_18882,N_19358);
xnor U20370 (N_20370,N_18968,N_19927);
or U20371 (N_20371,N_19298,N_19924);
nand U20372 (N_20372,N_19601,N_19196);
nor U20373 (N_20373,N_19118,N_19734);
and U20374 (N_20374,N_18821,N_19484);
xnor U20375 (N_20375,N_19558,N_19242);
nand U20376 (N_20376,N_18926,N_18869);
nor U20377 (N_20377,N_18960,N_19489);
or U20378 (N_20378,N_19185,N_19920);
and U20379 (N_20379,N_19133,N_19559);
and U20380 (N_20380,N_19912,N_19142);
or U20381 (N_20381,N_19232,N_18986);
nor U20382 (N_20382,N_19454,N_19586);
or U20383 (N_20383,N_19271,N_19941);
xnor U20384 (N_20384,N_19467,N_19300);
nor U20385 (N_20385,N_19387,N_19229);
nand U20386 (N_20386,N_19340,N_19774);
and U20387 (N_20387,N_19066,N_19218);
or U20388 (N_20388,N_19978,N_19552);
nor U20389 (N_20389,N_18965,N_19178);
nor U20390 (N_20390,N_19468,N_18777);
nor U20391 (N_20391,N_19163,N_19676);
xnor U20392 (N_20392,N_19798,N_19394);
and U20393 (N_20393,N_19277,N_19225);
nand U20394 (N_20394,N_19533,N_18876);
and U20395 (N_20395,N_19363,N_19923);
or U20396 (N_20396,N_18769,N_18763);
xor U20397 (N_20397,N_19683,N_19355);
nor U20398 (N_20398,N_18848,N_19939);
nand U20399 (N_20399,N_19254,N_19621);
nor U20400 (N_20400,N_18990,N_19189);
or U20401 (N_20401,N_18967,N_19434);
or U20402 (N_20402,N_19124,N_19327);
xnor U20403 (N_20403,N_19926,N_18979);
and U20404 (N_20404,N_19555,N_19925);
xnor U20405 (N_20405,N_18766,N_19100);
or U20406 (N_20406,N_18998,N_19595);
nand U20407 (N_20407,N_19014,N_19892);
xnor U20408 (N_20408,N_18945,N_18778);
and U20409 (N_20409,N_19170,N_18789);
xnor U20410 (N_20410,N_18883,N_19076);
and U20411 (N_20411,N_18887,N_19001);
or U20412 (N_20412,N_19534,N_19843);
nor U20413 (N_20413,N_18853,N_18951);
nand U20414 (N_20414,N_18807,N_19523);
nor U20415 (N_20415,N_19036,N_18761);
xnor U20416 (N_20416,N_18889,N_19128);
xnor U20417 (N_20417,N_18971,N_18897);
or U20418 (N_20418,N_19680,N_19687);
and U20419 (N_20419,N_19006,N_19838);
nand U20420 (N_20420,N_19965,N_19915);
and U20421 (N_20421,N_19754,N_19654);
nor U20422 (N_20422,N_19651,N_19681);
or U20423 (N_20423,N_19686,N_19712);
nor U20424 (N_20424,N_19331,N_19073);
xor U20425 (N_20425,N_19089,N_19703);
and U20426 (N_20426,N_19739,N_18854);
xnor U20427 (N_20427,N_18850,N_19209);
nand U20428 (N_20428,N_19759,N_19776);
nor U20429 (N_20429,N_19889,N_19070);
or U20430 (N_20430,N_19849,N_18792);
and U20431 (N_20431,N_19696,N_19023);
xor U20432 (N_20432,N_19626,N_19022);
nor U20433 (N_20433,N_18773,N_18793);
nor U20434 (N_20434,N_18980,N_18966);
nand U20435 (N_20435,N_19571,N_19824);
xor U20436 (N_20436,N_19872,N_19597);
and U20437 (N_20437,N_19129,N_19648);
or U20438 (N_20438,N_19581,N_19273);
nand U20439 (N_20439,N_19075,N_19551);
and U20440 (N_20440,N_18859,N_19195);
xnor U20441 (N_20441,N_19405,N_19995);
nor U20442 (N_20442,N_19543,N_19017);
xnor U20443 (N_20443,N_19026,N_19061);
and U20444 (N_20444,N_19123,N_19395);
or U20445 (N_20445,N_19922,N_19650);
nor U20446 (N_20446,N_19564,N_19876);
or U20447 (N_20447,N_19217,N_19311);
xnor U20448 (N_20448,N_19219,N_18962);
or U20449 (N_20449,N_19803,N_18969);
or U20450 (N_20450,N_19409,N_18891);
nor U20451 (N_20451,N_19455,N_19761);
xnor U20452 (N_20452,N_19445,N_19656);
nor U20453 (N_20453,N_19983,N_19143);
nand U20454 (N_20454,N_18833,N_19527);
or U20455 (N_20455,N_19874,N_19441);
and U20456 (N_20456,N_19634,N_19913);
nor U20457 (N_20457,N_19169,N_18803);
and U20458 (N_20458,N_19622,N_19632);
and U20459 (N_20459,N_19206,N_19919);
and U20460 (N_20460,N_19867,N_19275);
and U20461 (N_20461,N_19563,N_19668);
nand U20462 (N_20462,N_19346,N_18868);
and U20463 (N_20463,N_18863,N_19737);
or U20464 (N_20464,N_19842,N_19215);
nand U20465 (N_20465,N_19086,N_19582);
or U20466 (N_20466,N_19194,N_19099);
xnor U20467 (N_20467,N_19903,N_19056);
nand U20468 (N_20468,N_19975,N_19137);
nand U20469 (N_20469,N_19682,N_19979);
xnor U20470 (N_20470,N_18880,N_19270);
and U20471 (N_20471,N_19028,N_19399);
or U20472 (N_20472,N_19359,N_19371);
or U20473 (N_20473,N_19224,N_19307);
or U20474 (N_20474,N_19216,N_19444);
xor U20475 (N_20475,N_19373,N_19887);
and U20476 (N_20476,N_19408,N_19350);
or U20477 (N_20477,N_19884,N_19284);
nor U20478 (N_20478,N_19886,N_18851);
xnor U20479 (N_20479,N_19183,N_19772);
or U20480 (N_20480,N_19828,N_19548);
nand U20481 (N_20481,N_18762,N_19150);
nor U20482 (N_20482,N_19669,N_19430);
and U20483 (N_20483,N_19396,N_19362);
nor U20484 (N_20484,N_19815,N_19182);
nor U20485 (N_20485,N_19577,N_19854);
nor U20486 (N_20486,N_19494,N_19202);
nand U20487 (N_20487,N_18956,N_19615);
or U20488 (N_20488,N_18964,N_19093);
nand U20489 (N_20489,N_19745,N_19375);
and U20490 (N_20490,N_19719,N_19203);
and U20491 (N_20491,N_19625,N_19442);
nand U20492 (N_20492,N_18852,N_19760);
nor U20493 (N_20493,N_19624,N_19463);
nand U20494 (N_20494,N_19952,N_19894);
or U20495 (N_20495,N_18909,N_19390);
nand U20496 (N_20496,N_19306,N_19691);
and U20497 (N_20497,N_19019,N_19871);
nor U20498 (N_20498,N_18894,N_19435);
nor U20499 (N_20499,N_19684,N_19035);
nor U20500 (N_20500,N_19781,N_18943);
xnor U20501 (N_20501,N_18798,N_19720);
nand U20502 (N_20502,N_19635,N_18842);
and U20503 (N_20503,N_19532,N_19730);
xnor U20504 (N_20504,N_19758,N_19349);
and U20505 (N_20505,N_19818,N_19414);
nor U20506 (N_20506,N_19848,N_19909);
and U20507 (N_20507,N_19833,N_18950);
and U20508 (N_20508,N_19166,N_19031);
xnor U20509 (N_20509,N_18906,N_18750);
nand U20510 (N_20510,N_19173,N_19665);
or U20511 (N_20511,N_19064,N_19054);
or U20512 (N_20512,N_18957,N_19689);
nand U20513 (N_20513,N_19234,N_18819);
nor U20514 (N_20514,N_19641,N_18772);
xor U20515 (N_20515,N_19957,N_18947);
xor U20516 (N_20516,N_19646,N_19461);
and U20517 (N_20517,N_19566,N_19741);
or U20518 (N_20518,N_19805,N_19330);
nor U20519 (N_20519,N_19289,N_19018);
and U20520 (N_20520,N_19092,N_19243);
and U20521 (N_20521,N_19190,N_19762);
and U20522 (N_20522,N_19314,N_19767);
nor U20523 (N_20523,N_19763,N_18974);
nand U20524 (N_20524,N_18952,N_19214);
and U20525 (N_20525,N_19303,N_19973);
nor U20526 (N_20526,N_19706,N_19950);
nand U20527 (N_20527,N_19282,N_19085);
or U20528 (N_20528,N_19704,N_18832);
and U20529 (N_20529,N_19257,N_19738);
nand U20530 (N_20530,N_19751,N_19059);
nand U20531 (N_20531,N_19090,N_19744);
and U20532 (N_20532,N_19400,N_19213);
or U20533 (N_20533,N_19930,N_18805);
and U20534 (N_20534,N_19415,N_19211);
xnor U20535 (N_20535,N_19094,N_19904);
or U20536 (N_20536,N_19911,N_19860);
or U20537 (N_20537,N_19175,N_19486);
xnor U20538 (N_20538,N_18770,N_19630);
xor U20539 (N_20539,N_19205,N_19482);
and U20540 (N_20540,N_19773,N_19765);
or U20541 (N_20541,N_19230,N_19082);
or U20542 (N_20542,N_19495,N_18904);
and U20543 (N_20543,N_19743,N_19025);
nor U20544 (N_20544,N_19246,N_19320);
nor U20545 (N_20545,N_19005,N_19318);
nand U20546 (N_20546,N_19293,N_18846);
xor U20547 (N_20547,N_18790,N_19600);
or U20548 (N_20548,N_19974,N_18922);
and U20549 (N_20549,N_19393,N_19472);
xor U20550 (N_20550,N_18917,N_19608);
xor U20551 (N_20551,N_19545,N_19575);
and U20552 (N_20552,N_19736,N_19453);
xnor U20553 (N_20553,N_18994,N_19438);
or U20554 (N_20554,N_19418,N_19870);
nand U20555 (N_20555,N_19692,N_19197);
nand U20556 (N_20556,N_18771,N_19377);
nor U20557 (N_20557,N_19274,N_19250);
nand U20558 (N_20558,N_19055,N_18795);
xor U20559 (N_20559,N_19261,N_19891);
nor U20560 (N_20560,N_18757,N_19106);
or U20561 (N_20561,N_18774,N_19677);
nand U20562 (N_20562,N_19384,N_18946);
and U20563 (N_20563,N_18873,N_19452);
or U20564 (N_20564,N_19321,N_19063);
xor U20565 (N_20565,N_19378,N_19685);
xnor U20566 (N_20566,N_19694,N_18756);
and U20567 (N_20567,N_19988,N_19863);
or U20568 (N_20568,N_19748,N_19336);
nand U20569 (N_20569,N_19260,N_19898);
xor U20570 (N_20570,N_19338,N_19249);
or U20571 (N_20571,N_19041,N_19705);
nand U20572 (N_20572,N_19136,N_19051);
xnor U20573 (N_20573,N_19165,N_19008);
or U20574 (N_20574,N_19276,N_18983);
and U20575 (N_20575,N_18856,N_18902);
nand U20576 (N_20576,N_19491,N_18914);
nand U20577 (N_20577,N_19700,N_19517);
nand U20578 (N_20578,N_19456,N_18806);
nor U20579 (N_20579,N_19278,N_18836);
and U20580 (N_20580,N_19839,N_18977);
and U20581 (N_20581,N_19882,N_19228);
nand U20582 (N_20582,N_19652,N_19488);
nand U20583 (N_20583,N_19900,N_19883);
xor U20584 (N_20584,N_19933,N_19047);
nor U20585 (N_20585,N_19060,N_18881);
nor U20586 (N_20586,N_19841,N_19342);
or U20587 (N_20587,N_19013,N_18825);
nand U20588 (N_20588,N_19309,N_19366);
nand U20589 (N_20589,N_19207,N_18911);
nor U20590 (N_20590,N_19825,N_19766);
or U20591 (N_20591,N_19790,N_19670);
nand U20592 (N_20592,N_18818,N_19864);
nand U20593 (N_20593,N_19422,N_18927);
xnor U20594 (N_20594,N_19432,N_19437);
nor U20595 (N_20595,N_19176,N_19771);
nand U20596 (N_20596,N_19588,N_19485);
and U20597 (N_20597,N_19154,N_19935);
nand U20598 (N_20598,N_19590,N_18768);
and U20599 (N_20599,N_19784,N_19062);
xor U20600 (N_20600,N_19369,N_19322);
or U20601 (N_20601,N_19030,N_18875);
and U20602 (N_20602,N_19873,N_19814);
nand U20603 (N_20603,N_19413,N_19540);
xnor U20604 (N_20604,N_19813,N_19740);
nor U20605 (N_20605,N_18800,N_19573);
nor U20606 (N_20606,N_19786,N_19433);
nor U20607 (N_20607,N_19562,N_19715);
and U20608 (N_20608,N_19392,N_19423);
nor U20609 (N_20609,N_18981,N_18824);
or U20610 (N_20610,N_19530,N_18849);
nand U20611 (N_20611,N_19272,N_19819);
xnor U20612 (N_20612,N_18975,N_19966);
or U20613 (N_20613,N_18888,N_19946);
or U20614 (N_20614,N_19802,N_19783);
and U20615 (N_20615,N_19954,N_19316);
or U20616 (N_20616,N_19114,N_18779);
nand U20617 (N_20617,N_19238,N_18905);
nand U20618 (N_20618,N_19603,N_19557);
xor U20619 (N_20619,N_19351,N_18999);
nand U20620 (N_20620,N_19606,N_19388);
nor U20621 (N_20621,N_19464,N_19364);
nor U20622 (N_20622,N_19146,N_18923);
or U20623 (N_20623,N_19192,N_19513);
and U20624 (N_20624,N_18864,N_19536);
nand U20625 (N_20625,N_19225,N_19071);
or U20626 (N_20626,N_19408,N_19172);
or U20627 (N_20627,N_18921,N_19259);
xor U20628 (N_20628,N_19607,N_19161);
and U20629 (N_20629,N_19558,N_18764);
or U20630 (N_20630,N_19665,N_18795);
xnor U20631 (N_20631,N_19340,N_18914);
xor U20632 (N_20632,N_19602,N_18926);
xnor U20633 (N_20633,N_19610,N_19317);
nor U20634 (N_20634,N_19950,N_18991);
and U20635 (N_20635,N_19166,N_19271);
nand U20636 (N_20636,N_19546,N_19780);
nor U20637 (N_20637,N_18823,N_19619);
and U20638 (N_20638,N_19962,N_19398);
or U20639 (N_20639,N_19327,N_19965);
nor U20640 (N_20640,N_19836,N_18966);
or U20641 (N_20641,N_19707,N_19057);
or U20642 (N_20642,N_19165,N_19908);
and U20643 (N_20643,N_18888,N_18801);
nand U20644 (N_20644,N_19631,N_19701);
nand U20645 (N_20645,N_19710,N_18940);
nor U20646 (N_20646,N_19015,N_19080);
or U20647 (N_20647,N_19030,N_19260);
or U20648 (N_20648,N_19856,N_19378);
nand U20649 (N_20649,N_19430,N_19558);
nand U20650 (N_20650,N_18869,N_19348);
xnor U20651 (N_20651,N_18932,N_19268);
xor U20652 (N_20652,N_19788,N_19404);
xor U20653 (N_20653,N_18808,N_19149);
xnor U20654 (N_20654,N_19077,N_19382);
xor U20655 (N_20655,N_18974,N_18938);
or U20656 (N_20656,N_19332,N_18987);
nor U20657 (N_20657,N_19495,N_19272);
and U20658 (N_20658,N_19714,N_18896);
nand U20659 (N_20659,N_18785,N_18901);
xnor U20660 (N_20660,N_19699,N_19265);
or U20661 (N_20661,N_18756,N_18985);
nor U20662 (N_20662,N_19258,N_19501);
xor U20663 (N_20663,N_19325,N_18794);
xnor U20664 (N_20664,N_19340,N_18841);
and U20665 (N_20665,N_18873,N_19134);
and U20666 (N_20666,N_18897,N_19332);
or U20667 (N_20667,N_19629,N_19688);
or U20668 (N_20668,N_18930,N_19910);
xnor U20669 (N_20669,N_18877,N_19290);
and U20670 (N_20670,N_19584,N_19880);
xnor U20671 (N_20671,N_19771,N_19807);
nand U20672 (N_20672,N_19355,N_19363);
or U20673 (N_20673,N_19235,N_18804);
nand U20674 (N_20674,N_18916,N_19080);
or U20675 (N_20675,N_19081,N_19403);
xor U20676 (N_20676,N_19071,N_19373);
or U20677 (N_20677,N_18759,N_19822);
and U20678 (N_20678,N_19048,N_19406);
or U20679 (N_20679,N_19940,N_19086);
nor U20680 (N_20680,N_19541,N_18998);
xnor U20681 (N_20681,N_18878,N_18875);
or U20682 (N_20682,N_18905,N_19462);
nor U20683 (N_20683,N_19459,N_19075);
xnor U20684 (N_20684,N_18976,N_18883);
xnor U20685 (N_20685,N_19212,N_19076);
nand U20686 (N_20686,N_19648,N_19618);
xnor U20687 (N_20687,N_19678,N_19490);
nand U20688 (N_20688,N_19479,N_19044);
or U20689 (N_20689,N_19509,N_19165);
xnor U20690 (N_20690,N_19794,N_19896);
xor U20691 (N_20691,N_19518,N_19338);
nor U20692 (N_20692,N_19400,N_19138);
nand U20693 (N_20693,N_19696,N_18800);
nand U20694 (N_20694,N_19090,N_18984);
nand U20695 (N_20695,N_19826,N_19394);
nand U20696 (N_20696,N_19177,N_19458);
and U20697 (N_20697,N_18932,N_19784);
nor U20698 (N_20698,N_19059,N_19708);
and U20699 (N_20699,N_19959,N_19213);
xnor U20700 (N_20700,N_19197,N_18985);
nand U20701 (N_20701,N_18890,N_19058);
nand U20702 (N_20702,N_19165,N_19415);
nand U20703 (N_20703,N_19756,N_19274);
nor U20704 (N_20704,N_19899,N_19607);
and U20705 (N_20705,N_18969,N_19948);
nand U20706 (N_20706,N_19753,N_19325);
nor U20707 (N_20707,N_19297,N_19497);
nand U20708 (N_20708,N_18983,N_19662);
xnor U20709 (N_20709,N_19509,N_19487);
nand U20710 (N_20710,N_19385,N_18772);
and U20711 (N_20711,N_19248,N_19192);
nor U20712 (N_20712,N_19339,N_18865);
nand U20713 (N_20713,N_19294,N_19494);
nand U20714 (N_20714,N_19694,N_19913);
nand U20715 (N_20715,N_19413,N_19493);
and U20716 (N_20716,N_18954,N_19134);
or U20717 (N_20717,N_19949,N_19952);
xnor U20718 (N_20718,N_19103,N_19965);
or U20719 (N_20719,N_19178,N_19167);
nand U20720 (N_20720,N_19910,N_19013);
nor U20721 (N_20721,N_19629,N_19416);
and U20722 (N_20722,N_19563,N_18952);
and U20723 (N_20723,N_19297,N_19183);
xor U20724 (N_20724,N_19923,N_19978);
nand U20725 (N_20725,N_19845,N_18778);
or U20726 (N_20726,N_19227,N_19870);
nand U20727 (N_20727,N_19175,N_19385);
nand U20728 (N_20728,N_19659,N_19204);
and U20729 (N_20729,N_18952,N_19150);
or U20730 (N_20730,N_19691,N_18952);
and U20731 (N_20731,N_18864,N_19496);
xor U20732 (N_20732,N_19636,N_18767);
and U20733 (N_20733,N_19341,N_19666);
nor U20734 (N_20734,N_19769,N_19485);
or U20735 (N_20735,N_19602,N_19585);
or U20736 (N_20736,N_19738,N_18824);
and U20737 (N_20737,N_19950,N_19688);
nor U20738 (N_20738,N_19122,N_19537);
nand U20739 (N_20739,N_18925,N_19220);
xnor U20740 (N_20740,N_19128,N_19698);
and U20741 (N_20741,N_18907,N_19733);
nand U20742 (N_20742,N_19213,N_19612);
xnor U20743 (N_20743,N_19018,N_19619);
and U20744 (N_20744,N_18968,N_18800);
and U20745 (N_20745,N_19980,N_18871);
or U20746 (N_20746,N_18789,N_18828);
and U20747 (N_20747,N_19043,N_19516);
and U20748 (N_20748,N_19970,N_19874);
or U20749 (N_20749,N_19363,N_19896);
xnor U20750 (N_20750,N_19040,N_19525);
xor U20751 (N_20751,N_19160,N_19378);
nand U20752 (N_20752,N_19045,N_19882);
nor U20753 (N_20753,N_19605,N_19432);
nor U20754 (N_20754,N_19820,N_19638);
xnor U20755 (N_20755,N_18960,N_19019);
nand U20756 (N_20756,N_18908,N_18799);
and U20757 (N_20757,N_19884,N_19391);
and U20758 (N_20758,N_19935,N_19565);
or U20759 (N_20759,N_19163,N_19078);
nor U20760 (N_20760,N_19144,N_18840);
or U20761 (N_20761,N_19161,N_19203);
and U20762 (N_20762,N_19915,N_18875);
and U20763 (N_20763,N_19838,N_19437);
nor U20764 (N_20764,N_19534,N_19754);
nor U20765 (N_20765,N_19744,N_19394);
nor U20766 (N_20766,N_19418,N_19362);
and U20767 (N_20767,N_19139,N_19108);
nor U20768 (N_20768,N_19508,N_19340);
nor U20769 (N_20769,N_19849,N_19344);
or U20770 (N_20770,N_19601,N_19634);
or U20771 (N_20771,N_19505,N_19538);
xnor U20772 (N_20772,N_19974,N_19080);
and U20773 (N_20773,N_19299,N_19766);
nor U20774 (N_20774,N_19060,N_19933);
xor U20775 (N_20775,N_18760,N_18983);
and U20776 (N_20776,N_19549,N_19208);
nand U20777 (N_20777,N_19648,N_19470);
xnor U20778 (N_20778,N_19500,N_18777);
nor U20779 (N_20779,N_18923,N_19959);
or U20780 (N_20780,N_19841,N_19758);
or U20781 (N_20781,N_19543,N_19292);
or U20782 (N_20782,N_19001,N_19805);
xnor U20783 (N_20783,N_18963,N_18938);
xnor U20784 (N_20784,N_19218,N_19857);
nand U20785 (N_20785,N_19152,N_18895);
nand U20786 (N_20786,N_19816,N_19779);
or U20787 (N_20787,N_19881,N_19370);
nor U20788 (N_20788,N_19210,N_19639);
and U20789 (N_20789,N_19777,N_19036);
nand U20790 (N_20790,N_19219,N_19233);
nand U20791 (N_20791,N_19913,N_19547);
and U20792 (N_20792,N_18849,N_18887);
and U20793 (N_20793,N_19410,N_19343);
xor U20794 (N_20794,N_19573,N_18987);
nor U20795 (N_20795,N_19206,N_19503);
and U20796 (N_20796,N_18975,N_19314);
and U20797 (N_20797,N_19263,N_19866);
or U20798 (N_20798,N_19008,N_19062);
nand U20799 (N_20799,N_19008,N_19178);
or U20800 (N_20800,N_19314,N_19808);
or U20801 (N_20801,N_19370,N_19801);
xor U20802 (N_20802,N_19491,N_18942);
and U20803 (N_20803,N_19706,N_19001);
and U20804 (N_20804,N_18792,N_19894);
nand U20805 (N_20805,N_18939,N_19186);
and U20806 (N_20806,N_19730,N_19380);
and U20807 (N_20807,N_19620,N_19649);
nand U20808 (N_20808,N_19726,N_19486);
nand U20809 (N_20809,N_19239,N_19106);
and U20810 (N_20810,N_19287,N_19401);
or U20811 (N_20811,N_19237,N_18930);
xor U20812 (N_20812,N_19669,N_19784);
nor U20813 (N_20813,N_19108,N_19828);
xor U20814 (N_20814,N_19451,N_18916);
or U20815 (N_20815,N_19922,N_19110);
nand U20816 (N_20816,N_19370,N_19505);
nor U20817 (N_20817,N_19940,N_19342);
and U20818 (N_20818,N_19380,N_18767);
and U20819 (N_20819,N_19517,N_19762);
nor U20820 (N_20820,N_19024,N_19647);
and U20821 (N_20821,N_19245,N_19388);
nand U20822 (N_20822,N_19120,N_19898);
and U20823 (N_20823,N_19546,N_19886);
and U20824 (N_20824,N_18874,N_19628);
xnor U20825 (N_20825,N_19632,N_19157);
xnor U20826 (N_20826,N_19990,N_19855);
xnor U20827 (N_20827,N_19193,N_18876);
nand U20828 (N_20828,N_19430,N_19650);
and U20829 (N_20829,N_19681,N_19429);
xnor U20830 (N_20830,N_19474,N_19809);
nand U20831 (N_20831,N_18901,N_18860);
nor U20832 (N_20832,N_18964,N_19107);
or U20833 (N_20833,N_18828,N_19198);
xnor U20834 (N_20834,N_18840,N_19074);
nand U20835 (N_20835,N_19896,N_19378);
or U20836 (N_20836,N_19990,N_19103);
xnor U20837 (N_20837,N_18771,N_19851);
and U20838 (N_20838,N_18873,N_19492);
or U20839 (N_20839,N_19145,N_19210);
nor U20840 (N_20840,N_19735,N_18818);
nor U20841 (N_20841,N_19990,N_18763);
or U20842 (N_20842,N_19142,N_19303);
nand U20843 (N_20843,N_19391,N_19302);
nand U20844 (N_20844,N_19343,N_19333);
nand U20845 (N_20845,N_19393,N_19513);
nand U20846 (N_20846,N_19483,N_19935);
and U20847 (N_20847,N_18912,N_19771);
nor U20848 (N_20848,N_19517,N_19689);
nor U20849 (N_20849,N_19430,N_19803);
and U20850 (N_20850,N_19325,N_19090);
xnor U20851 (N_20851,N_19393,N_19674);
nor U20852 (N_20852,N_19581,N_19089);
nand U20853 (N_20853,N_19096,N_18910);
nor U20854 (N_20854,N_19793,N_19471);
xor U20855 (N_20855,N_19195,N_18903);
and U20856 (N_20856,N_19356,N_19629);
nand U20857 (N_20857,N_19063,N_19797);
and U20858 (N_20858,N_19851,N_19381);
or U20859 (N_20859,N_19668,N_19310);
nand U20860 (N_20860,N_19001,N_19772);
nor U20861 (N_20861,N_19747,N_18889);
nand U20862 (N_20862,N_18881,N_19070);
and U20863 (N_20863,N_19362,N_18945);
xnor U20864 (N_20864,N_19502,N_19629);
xnor U20865 (N_20865,N_19160,N_19214);
and U20866 (N_20866,N_18913,N_19894);
or U20867 (N_20867,N_19191,N_19223);
xor U20868 (N_20868,N_19897,N_19630);
or U20869 (N_20869,N_18887,N_19446);
xor U20870 (N_20870,N_19659,N_19554);
xnor U20871 (N_20871,N_19591,N_19910);
nand U20872 (N_20872,N_19915,N_19055);
or U20873 (N_20873,N_19376,N_19370);
or U20874 (N_20874,N_19653,N_19696);
nor U20875 (N_20875,N_19020,N_19110);
or U20876 (N_20876,N_19411,N_19037);
and U20877 (N_20877,N_19456,N_19514);
nand U20878 (N_20878,N_19292,N_18967);
xnor U20879 (N_20879,N_19111,N_19621);
nand U20880 (N_20880,N_18779,N_18987);
nand U20881 (N_20881,N_19794,N_18888);
and U20882 (N_20882,N_19298,N_19986);
nand U20883 (N_20883,N_19822,N_18873);
xnor U20884 (N_20884,N_19391,N_19055);
nand U20885 (N_20885,N_19620,N_18827);
xor U20886 (N_20886,N_18989,N_19505);
nand U20887 (N_20887,N_19363,N_19826);
and U20888 (N_20888,N_19900,N_19241);
nor U20889 (N_20889,N_19229,N_19747);
and U20890 (N_20890,N_19559,N_19643);
nor U20891 (N_20891,N_19673,N_19756);
or U20892 (N_20892,N_19973,N_19465);
and U20893 (N_20893,N_19369,N_19986);
xor U20894 (N_20894,N_19903,N_18998);
nor U20895 (N_20895,N_19754,N_19418);
and U20896 (N_20896,N_19307,N_19834);
nand U20897 (N_20897,N_19752,N_19769);
nor U20898 (N_20898,N_18905,N_18765);
nand U20899 (N_20899,N_19803,N_19668);
xor U20900 (N_20900,N_19780,N_18874);
and U20901 (N_20901,N_19108,N_19590);
and U20902 (N_20902,N_19732,N_18898);
nor U20903 (N_20903,N_19484,N_19453);
and U20904 (N_20904,N_19449,N_19696);
xor U20905 (N_20905,N_19105,N_19224);
and U20906 (N_20906,N_19976,N_19587);
xor U20907 (N_20907,N_19356,N_19343);
nand U20908 (N_20908,N_18763,N_19790);
nor U20909 (N_20909,N_19737,N_18992);
and U20910 (N_20910,N_19856,N_18810);
nor U20911 (N_20911,N_19032,N_18913);
xor U20912 (N_20912,N_19718,N_19885);
nor U20913 (N_20913,N_19892,N_19662);
and U20914 (N_20914,N_19828,N_19713);
xnor U20915 (N_20915,N_18920,N_19121);
nand U20916 (N_20916,N_19571,N_18805);
nor U20917 (N_20917,N_19084,N_19912);
or U20918 (N_20918,N_19617,N_18792);
nor U20919 (N_20919,N_18880,N_18851);
and U20920 (N_20920,N_19485,N_19665);
nor U20921 (N_20921,N_19563,N_18957);
and U20922 (N_20922,N_18959,N_19247);
or U20923 (N_20923,N_19188,N_19551);
xor U20924 (N_20924,N_19172,N_19272);
and U20925 (N_20925,N_19488,N_19572);
or U20926 (N_20926,N_18976,N_19891);
and U20927 (N_20927,N_19810,N_19285);
nand U20928 (N_20928,N_19279,N_19620);
nand U20929 (N_20929,N_19507,N_19013);
xor U20930 (N_20930,N_19126,N_18891);
nor U20931 (N_20931,N_19830,N_18856);
or U20932 (N_20932,N_19014,N_19638);
nor U20933 (N_20933,N_19828,N_19629);
xnor U20934 (N_20934,N_18876,N_19552);
or U20935 (N_20935,N_19662,N_19898);
nand U20936 (N_20936,N_19193,N_19063);
or U20937 (N_20937,N_19748,N_18826);
and U20938 (N_20938,N_18940,N_19079);
or U20939 (N_20939,N_18769,N_18967);
xor U20940 (N_20940,N_19783,N_18851);
nand U20941 (N_20941,N_19160,N_18962);
xor U20942 (N_20942,N_19179,N_18918);
nand U20943 (N_20943,N_18888,N_19111);
and U20944 (N_20944,N_19826,N_19856);
nor U20945 (N_20945,N_19993,N_18834);
and U20946 (N_20946,N_19651,N_19467);
xnor U20947 (N_20947,N_19382,N_19784);
nor U20948 (N_20948,N_18906,N_19772);
xnor U20949 (N_20949,N_19729,N_19370);
nor U20950 (N_20950,N_19441,N_19544);
and U20951 (N_20951,N_19125,N_19257);
and U20952 (N_20952,N_19763,N_18968);
and U20953 (N_20953,N_19259,N_19266);
nand U20954 (N_20954,N_19029,N_19122);
and U20955 (N_20955,N_19998,N_19241);
or U20956 (N_20956,N_18862,N_19696);
and U20957 (N_20957,N_19491,N_19621);
nand U20958 (N_20958,N_19091,N_19402);
and U20959 (N_20959,N_18862,N_18909);
nand U20960 (N_20960,N_19227,N_19468);
and U20961 (N_20961,N_19532,N_19528);
and U20962 (N_20962,N_18836,N_19722);
nor U20963 (N_20963,N_18906,N_19526);
nor U20964 (N_20964,N_19065,N_19915);
or U20965 (N_20965,N_19168,N_19761);
nand U20966 (N_20966,N_19013,N_18791);
xnor U20967 (N_20967,N_19071,N_19994);
xnor U20968 (N_20968,N_19667,N_19109);
nor U20969 (N_20969,N_19572,N_19826);
nand U20970 (N_20970,N_19645,N_19129);
or U20971 (N_20971,N_19111,N_18910);
xnor U20972 (N_20972,N_19028,N_19152);
nand U20973 (N_20973,N_19263,N_19050);
nand U20974 (N_20974,N_19341,N_19285);
nor U20975 (N_20975,N_19699,N_19805);
xnor U20976 (N_20976,N_19426,N_19856);
nand U20977 (N_20977,N_19134,N_19887);
and U20978 (N_20978,N_19529,N_19359);
nor U20979 (N_20979,N_19220,N_19550);
or U20980 (N_20980,N_19031,N_18928);
xnor U20981 (N_20981,N_19228,N_19071);
xor U20982 (N_20982,N_19422,N_19428);
or U20983 (N_20983,N_19238,N_19155);
or U20984 (N_20984,N_19651,N_19931);
nand U20985 (N_20985,N_19691,N_19073);
and U20986 (N_20986,N_19136,N_18787);
nand U20987 (N_20987,N_19699,N_19217);
nor U20988 (N_20988,N_19877,N_19624);
nor U20989 (N_20989,N_19577,N_19940);
nor U20990 (N_20990,N_19790,N_18779);
nor U20991 (N_20991,N_19128,N_18875);
nor U20992 (N_20992,N_19482,N_19934);
nor U20993 (N_20993,N_18953,N_19258);
nor U20994 (N_20994,N_19321,N_19563);
xor U20995 (N_20995,N_19270,N_19662);
or U20996 (N_20996,N_19595,N_19112);
nor U20997 (N_20997,N_18769,N_19213);
xnor U20998 (N_20998,N_18826,N_19468);
nand U20999 (N_20999,N_18864,N_19208);
xor U21000 (N_21000,N_19463,N_19807);
xor U21001 (N_21001,N_19550,N_19219);
xor U21002 (N_21002,N_19889,N_19100);
nor U21003 (N_21003,N_19110,N_19060);
or U21004 (N_21004,N_19438,N_19504);
and U21005 (N_21005,N_19163,N_19450);
or U21006 (N_21006,N_19417,N_19209);
nand U21007 (N_21007,N_18970,N_19295);
and U21008 (N_21008,N_19284,N_18758);
xor U21009 (N_21009,N_19438,N_19829);
nor U21010 (N_21010,N_19378,N_19572);
and U21011 (N_21011,N_19032,N_19667);
nor U21012 (N_21012,N_19601,N_19869);
nor U21013 (N_21013,N_19203,N_19669);
xor U21014 (N_21014,N_19391,N_18762);
and U21015 (N_21015,N_19590,N_19988);
nor U21016 (N_21016,N_19251,N_19723);
xnor U21017 (N_21017,N_19860,N_19692);
or U21018 (N_21018,N_19599,N_18955);
nor U21019 (N_21019,N_19643,N_19562);
xnor U21020 (N_21020,N_18878,N_19300);
or U21021 (N_21021,N_19468,N_19038);
xor U21022 (N_21022,N_19947,N_19883);
xor U21023 (N_21023,N_19780,N_19447);
or U21024 (N_21024,N_19045,N_19954);
xnor U21025 (N_21025,N_19049,N_19144);
and U21026 (N_21026,N_19845,N_19380);
nor U21027 (N_21027,N_18779,N_19682);
nor U21028 (N_21028,N_19400,N_19407);
and U21029 (N_21029,N_18988,N_19884);
and U21030 (N_21030,N_18839,N_19278);
and U21031 (N_21031,N_19609,N_19735);
nor U21032 (N_21032,N_19107,N_19804);
xor U21033 (N_21033,N_19832,N_19116);
nor U21034 (N_21034,N_19852,N_19026);
xor U21035 (N_21035,N_19381,N_19983);
xnor U21036 (N_21036,N_19458,N_19359);
nor U21037 (N_21037,N_19214,N_19226);
xor U21038 (N_21038,N_18929,N_19420);
nor U21039 (N_21039,N_19042,N_19829);
nand U21040 (N_21040,N_19561,N_19587);
and U21041 (N_21041,N_19144,N_19335);
or U21042 (N_21042,N_19123,N_19366);
or U21043 (N_21043,N_19337,N_19507);
xnor U21044 (N_21044,N_19255,N_19801);
nor U21045 (N_21045,N_19609,N_19286);
nor U21046 (N_21046,N_18880,N_19123);
and U21047 (N_21047,N_19952,N_19109);
nand U21048 (N_21048,N_19240,N_19580);
nand U21049 (N_21049,N_18978,N_19088);
nand U21050 (N_21050,N_18931,N_19450);
nor U21051 (N_21051,N_18899,N_19389);
nor U21052 (N_21052,N_19329,N_19778);
xnor U21053 (N_21053,N_19269,N_19989);
and U21054 (N_21054,N_19764,N_18848);
xor U21055 (N_21055,N_18987,N_19578);
and U21056 (N_21056,N_19080,N_19815);
nor U21057 (N_21057,N_18911,N_19365);
and U21058 (N_21058,N_19533,N_19547);
and U21059 (N_21059,N_19360,N_19904);
or U21060 (N_21060,N_19556,N_19208);
xnor U21061 (N_21061,N_18875,N_19820);
nor U21062 (N_21062,N_19243,N_18911);
or U21063 (N_21063,N_19614,N_18834);
and U21064 (N_21064,N_19396,N_19454);
xor U21065 (N_21065,N_19200,N_19393);
nor U21066 (N_21066,N_19448,N_19263);
xnor U21067 (N_21067,N_19237,N_19856);
nor U21068 (N_21068,N_19872,N_18883);
nand U21069 (N_21069,N_19624,N_18839);
nand U21070 (N_21070,N_19563,N_19376);
nand U21071 (N_21071,N_19374,N_19315);
nand U21072 (N_21072,N_18965,N_19640);
xnor U21073 (N_21073,N_19407,N_19013);
and U21074 (N_21074,N_19245,N_19100);
nand U21075 (N_21075,N_19498,N_19602);
and U21076 (N_21076,N_19419,N_19062);
or U21077 (N_21077,N_19913,N_19910);
nor U21078 (N_21078,N_19271,N_19449);
nand U21079 (N_21079,N_19739,N_19537);
xor U21080 (N_21080,N_19581,N_19073);
nor U21081 (N_21081,N_19382,N_18887);
nor U21082 (N_21082,N_19326,N_19757);
or U21083 (N_21083,N_18985,N_19791);
and U21084 (N_21084,N_19336,N_19466);
or U21085 (N_21085,N_19902,N_19316);
nor U21086 (N_21086,N_19356,N_18779);
nor U21087 (N_21087,N_18845,N_19914);
nor U21088 (N_21088,N_18915,N_18772);
xor U21089 (N_21089,N_19574,N_19077);
nand U21090 (N_21090,N_18908,N_19528);
or U21091 (N_21091,N_19192,N_19282);
nand U21092 (N_21092,N_19253,N_19028);
nand U21093 (N_21093,N_19071,N_19333);
or U21094 (N_21094,N_19822,N_19971);
nor U21095 (N_21095,N_19674,N_19111);
xnor U21096 (N_21096,N_19746,N_19498);
nand U21097 (N_21097,N_19938,N_19263);
xnor U21098 (N_21098,N_19833,N_19337);
and U21099 (N_21099,N_19412,N_19748);
nand U21100 (N_21100,N_19148,N_19862);
xnor U21101 (N_21101,N_19701,N_19859);
and U21102 (N_21102,N_19392,N_18854);
or U21103 (N_21103,N_19072,N_19537);
nor U21104 (N_21104,N_19450,N_19098);
or U21105 (N_21105,N_19623,N_18799);
nor U21106 (N_21106,N_19075,N_19176);
and U21107 (N_21107,N_19662,N_19627);
or U21108 (N_21108,N_18913,N_19769);
or U21109 (N_21109,N_18948,N_19818);
and U21110 (N_21110,N_19203,N_19882);
and U21111 (N_21111,N_19707,N_19640);
or U21112 (N_21112,N_18802,N_19646);
and U21113 (N_21113,N_19927,N_19096);
or U21114 (N_21114,N_18991,N_19759);
or U21115 (N_21115,N_19068,N_19320);
xor U21116 (N_21116,N_19645,N_19475);
and U21117 (N_21117,N_18955,N_19339);
and U21118 (N_21118,N_19157,N_19802);
nor U21119 (N_21119,N_19068,N_19156);
and U21120 (N_21120,N_19905,N_19422);
xnor U21121 (N_21121,N_19125,N_19068);
and U21122 (N_21122,N_19400,N_19109);
nor U21123 (N_21123,N_18845,N_19009);
or U21124 (N_21124,N_19626,N_19593);
nor U21125 (N_21125,N_19881,N_19337);
xnor U21126 (N_21126,N_19290,N_19544);
nand U21127 (N_21127,N_18855,N_19712);
nor U21128 (N_21128,N_18926,N_19634);
nand U21129 (N_21129,N_19645,N_19271);
nor U21130 (N_21130,N_19906,N_19668);
nand U21131 (N_21131,N_19882,N_19728);
and U21132 (N_21132,N_18892,N_19033);
and U21133 (N_21133,N_19559,N_19147);
and U21134 (N_21134,N_19942,N_19517);
nand U21135 (N_21135,N_19356,N_19702);
xor U21136 (N_21136,N_19750,N_19504);
or U21137 (N_21137,N_19065,N_19149);
xnor U21138 (N_21138,N_19658,N_19315);
and U21139 (N_21139,N_19700,N_19156);
and U21140 (N_21140,N_18912,N_19741);
or U21141 (N_21141,N_19580,N_19555);
and U21142 (N_21142,N_19238,N_19867);
nand U21143 (N_21143,N_19504,N_18853);
nand U21144 (N_21144,N_19466,N_19469);
xor U21145 (N_21145,N_19095,N_19357);
or U21146 (N_21146,N_19533,N_18769);
or U21147 (N_21147,N_19122,N_18941);
nor U21148 (N_21148,N_18994,N_19160);
or U21149 (N_21149,N_19763,N_18909);
or U21150 (N_21150,N_19458,N_18864);
xor U21151 (N_21151,N_19353,N_19951);
nand U21152 (N_21152,N_18935,N_19907);
nor U21153 (N_21153,N_19231,N_19790);
xor U21154 (N_21154,N_19984,N_19374);
and U21155 (N_21155,N_19667,N_18784);
or U21156 (N_21156,N_19765,N_19546);
and U21157 (N_21157,N_19953,N_19405);
and U21158 (N_21158,N_18796,N_19954);
nor U21159 (N_21159,N_19942,N_19255);
or U21160 (N_21160,N_19507,N_18770);
nand U21161 (N_21161,N_19631,N_19330);
and U21162 (N_21162,N_19324,N_19463);
nand U21163 (N_21163,N_19324,N_19464);
and U21164 (N_21164,N_19207,N_19363);
nor U21165 (N_21165,N_18762,N_19722);
and U21166 (N_21166,N_19464,N_19982);
nand U21167 (N_21167,N_19051,N_18765);
nor U21168 (N_21168,N_19753,N_19892);
nand U21169 (N_21169,N_19518,N_19423);
or U21170 (N_21170,N_19184,N_19057);
nand U21171 (N_21171,N_18917,N_18808);
or U21172 (N_21172,N_19327,N_19125);
nor U21173 (N_21173,N_19895,N_19773);
and U21174 (N_21174,N_19692,N_19281);
nand U21175 (N_21175,N_19594,N_18921);
nand U21176 (N_21176,N_18960,N_19571);
nand U21177 (N_21177,N_18864,N_19639);
or U21178 (N_21178,N_19302,N_19072);
nor U21179 (N_21179,N_19510,N_18904);
nand U21180 (N_21180,N_18858,N_19792);
or U21181 (N_21181,N_19843,N_19846);
nand U21182 (N_21182,N_19677,N_19817);
xor U21183 (N_21183,N_19927,N_19080);
and U21184 (N_21184,N_19045,N_19770);
and U21185 (N_21185,N_19348,N_19011);
and U21186 (N_21186,N_19630,N_18810);
nand U21187 (N_21187,N_19206,N_19322);
xnor U21188 (N_21188,N_19588,N_19566);
nor U21189 (N_21189,N_19133,N_19643);
and U21190 (N_21190,N_19352,N_18874);
xnor U21191 (N_21191,N_19515,N_19993);
or U21192 (N_21192,N_19756,N_18857);
and U21193 (N_21193,N_19879,N_19696);
nor U21194 (N_21194,N_19563,N_19045);
and U21195 (N_21195,N_18983,N_19193);
and U21196 (N_21196,N_18801,N_19256);
xor U21197 (N_21197,N_19345,N_19860);
and U21198 (N_21198,N_19651,N_19097);
nand U21199 (N_21199,N_18936,N_19776);
or U21200 (N_21200,N_18856,N_19319);
nor U21201 (N_21201,N_19924,N_19398);
nor U21202 (N_21202,N_19762,N_19457);
xnor U21203 (N_21203,N_19212,N_19278);
nand U21204 (N_21204,N_19665,N_19765);
or U21205 (N_21205,N_19930,N_19357);
xor U21206 (N_21206,N_18827,N_19445);
or U21207 (N_21207,N_19721,N_19292);
and U21208 (N_21208,N_19437,N_19205);
nand U21209 (N_21209,N_19878,N_19448);
nand U21210 (N_21210,N_18779,N_19899);
xnor U21211 (N_21211,N_19696,N_19263);
and U21212 (N_21212,N_19501,N_19017);
xor U21213 (N_21213,N_19793,N_19925);
or U21214 (N_21214,N_19203,N_19614);
xor U21215 (N_21215,N_19396,N_19584);
and U21216 (N_21216,N_18764,N_18790);
and U21217 (N_21217,N_18760,N_18926);
or U21218 (N_21218,N_19310,N_19590);
xor U21219 (N_21219,N_19425,N_19036);
and U21220 (N_21220,N_19275,N_19747);
nor U21221 (N_21221,N_19100,N_18910);
nand U21222 (N_21222,N_19976,N_19485);
xor U21223 (N_21223,N_19861,N_19383);
xnor U21224 (N_21224,N_19718,N_19618);
or U21225 (N_21225,N_19807,N_19122);
or U21226 (N_21226,N_19529,N_19322);
or U21227 (N_21227,N_19595,N_19807);
xor U21228 (N_21228,N_19292,N_19603);
or U21229 (N_21229,N_19897,N_19948);
or U21230 (N_21230,N_19010,N_19044);
or U21231 (N_21231,N_19703,N_19476);
and U21232 (N_21232,N_19608,N_19988);
or U21233 (N_21233,N_19098,N_18935);
and U21234 (N_21234,N_19251,N_19641);
nor U21235 (N_21235,N_19697,N_19019);
and U21236 (N_21236,N_19615,N_19906);
nand U21237 (N_21237,N_19243,N_19780);
nand U21238 (N_21238,N_19758,N_19446);
nor U21239 (N_21239,N_19015,N_18810);
or U21240 (N_21240,N_18907,N_18885);
nor U21241 (N_21241,N_19753,N_19109);
and U21242 (N_21242,N_19424,N_19275);
or U21243 (N_21243,N_19391,N_19078);
xnor U21244 (N_21244,N_19806,N_19959);
or U21245 (N_21245,N_19497,N_18946);
and U21246 (N_21246,N_19686,N_19884);
and U21247 (N_21247,N_19212,N_19587);
and U21248 (N_21248,N_19439,N_19145);
nand U21249 (N_21249,N_18858,N_18818);
and U21250 (N_21250,N_21052,N_20964);
or U21251 (N_21251,N_20565,N_20749);
nor U21252 (N_21252,N_20954,N_20935);
or U21253 (N_21253,N_21203,N_20645);
and U21254 (N_21254,N_20280,N_20063);
nor U21255 (N_21255,N_21104,N_21219);
or U21256 (N_21256,N_20884,N_20201);
xnor U21257 (N_21257,N_20829,N_20497);
nor U21258 (N_21258,N_20109,N_21140);
nand U21259 (N_21259,N_20902,N_20222);
xor U21260 (N_21260,N_20499,N_21167);
and U21261 (N_21261,N_20786,N_20694);
nand U21262 (N_21262,N_21247,N_20721);
nor U21263 (N_21263,N_21188,N_20292);
or U21264 (N_21264,N_20197,N_20287);
nor U21265 (N_21265,N_20804,N_21003);
xor U21266 (N_21266,N_20479,N_20074);
xor U21267 (N_21267,N_20324,N_20315);
or U21268 (N_21268,N_20569,N_20370);
nor U21269 (N_21269,N_20367,N_20757);
and U21270 (N_21270,N_20088,N_20971);
xnor U21271 (N_21271,N_20910,N_20758);
and U21272 (N_21272,N_21205,N_20769);
xnor U21273 (N_21273,N_20234,N_20007);
xor U21274 (N_21274,N_20493,N_20768);
nor U21275 (N_21275,N_20520,N_20089);
xor U21276 (N_21276,N_20422,N_20306);
xor U21277 (N_21277,N_20153,N_20257);
and U21278 (N_21278,N_20115,N_20242);
nor U21279 (N_21279,N_20177,N_20340);
and U21280 (N_21280,N_20724,N_21149);
nor U21281 (N_21281,N_21183,N_20219);
and U21282 (N_21282,N_20097,N_20094);
or U21283 (N_21283,N_20132,N_21084);
nor U21284 (N_21284,N_20398,N_20502);
xnor U21285 (N_21285,N_20859,N_21064);
xor U21286 (N_21286,N_21120,N_20464);
and U21287 (N_21287,N_20393,N_20707);
and U21288 (N_21288,N_20833,N_21193);
nor U21289 (N_21289,N_21077,N_21006);
nor U21290 (N_21290,N_20861,N_20245);
or U21291 (N_21291,N_21156,N_20547);
nor U21292 (N_21292,N_20686,N_20874);
nand U21293 (N_21293,N_20380,N_20791);
xor U21294 (N_21294,N_20086,N_20326);
nor U21295 (N_21295,N_20276,N_20171);
or U21296 (N_21296,N_20400,N_20210);
nand U21297 (N_21297,N_20933,N_20535);
nor U21298 (N_21298,N_20920,N_20545);
xor U21299 (N_21299,N_20266,N_21039);
and U21300 (N_21300,N_20173,N_20608);
nor U21301 (N_21301,N_20461,N_20390);
or U21302 (N_21302,N_20442,N_20636);
nor U21303 (N_21303,N_21143,N_21015);
nor U21304 (N_21304,N_20033,N_20947);
xnor U21305 (N_21305,N_21030,N_20144);
and U21306 (N_21306,N_20555,N_20263);
or U21307 (N_21307,N_20277,N_20489);
nor U21308 (N_21308,N_21046,N_20426);
or U21309 (N_21309,N_21029,N_20695);
nor U21310 (N_21310,N_20381,N_20647);
and U21311 (N_21311,N_20262,N_20925);
and U21312 (N_21312,N_21108,N_21142);
or U21313 (N_21313,N_20844,N_20514);
or U21314 (N_21314,N_20800,N_20581);
xnor U21315 (N_21315,N_21199,N_20830);
xnor U21316 (N_21316,N_21150,N_20548);
nor U21317 (N_21317,N_20043,N_20612);
nand U21318 (N_21318,N_20665,N_20605);
and U21319 (N_21319,N_20602,N_21189);
nor U21320 (N_21320,N_21169,N_20772);
nor U21321 (N_21321,N_21034,N_21095);
and U21322 (N_21322,N_20477,N_20842);
and U21323 (N_21323,N_20092,N_20737);
and U21324 (N_21324,N_20738,N_20813);
nor U21325 (N_21325,N_21002,N_20190);
nand U21326 (N_21326,N_20078,N_20974);
nor U21327 (N_21327,N_20530,N_21222);
xor U21328 (N_21328,N_21135,N_20396);
nor U21329 (N_21329,N_20147,N_21014);
nand U21330 (N_21330,N_20610,N_20876);
and U21331 (N_21331,N_20207,N_21026);
nor U21332 (N_21332,N_20484,N_20658);
xnor U21333 (N_21333,N_21066,N_20471);
and U21334 (N_21334,N_20538,N_20453);
nor U21335 (N_21335,N_20918,N_20194);
or U21336 (N_21336,N_20973,N_20812);
nor U21337 (N_21337,N_20205,N_20577);
or U21338 (N_21338,N_20771,N_20354);
nor U21339 (N_21339,N_20717,N_20452);
nor U21340 (N_21340,N_20766,N_20533);
and U21341 (N_21341,N_20650,N_21195);
or U21342 (N_21342,N_20914,N_20170);
xor U21343 (N_21343,N_20655,N_20268);
xnor U21344 (N_21344,N_20022,N_20403);
nand U21345 (N_21345,N_20251,N_20901);
or U21346 (N_21346,N_20810,N_20590);
nor U21347 (N_21347,N_20120,N_20591);
nand U21348 (N_21348,N_20875,N_20013);
and U21349 (N_21349,N_20437,N_20822);
nor U21350 (N_21350,N_20241,N_20832);
nand U21351 (N_21351,N_20006,N_20085);
nor U21352 (N_21352,N_20880,N_21214);
nand U21353 (N_21353,N_20139,N_21249);
nand U21354 (N_21354,N_20339,N_20248);
nor U21355 (N_21355,N_20575,N_20274);
nand U21356 (N_21356,N_20388,N_20482);
and U21357 (N_21357,N_20728,N_20365);
or U21358 (N_21358,N_20269,N_21005);
or U21359 (N_21359,N_20077,N_20035);
xor U21360 (N_21360,N_20767,N_20878);
nand U21361 (N_21361,N_20010,N_20183);
nand U21362 (N_21362,N_20056,N_21239);
or U21363 (N_21363,N_20179,N_20322);
nor U21364 (N_21364,N_20950,N_21109);
xor U21365 (N_21365,N_20617,N_21098);
xnor U21366 (N_21366,N_20927,N_20379);
nor U21367 (N_21367,N_21102,N_20506);
nor U21368 (N_21368,N_20250,N_21232);
xnor U21369 (N_21369,N_21168,N_21117);
nand U21370 (N_21370,N_21107,N_21067);
nand U21371 (N_21371,N_20188,N_21136);
or U21372 (N_21372,N_21160,N_20126);
or U21373 (N_21373,N_20977,N_20095);
nand U21374 (N_21374,N_20220,N_21151);
or U21375 (N_21375,N_20849,N_20116);
nand U21376 (N_21376,N_21073,N_20318);
xnor U21377 (N_21377,N_20402,N_20818);
xnor U21378 (N_21378,N_20456,N_20510);
nor U21379 (N_21379,N_20331,N_20049);
and U21380 (N_21380,N_21091,N_21134);
and U21381 (N_21381,N_20106,N_20785);
nor U21382 (N_21382,N_20748,N_20899);
nand U21383 (N_21383,N_20395,N_20789);
nor U21384 (N_21384,N_20713,N_20890);
xor U21385 (N_21385,N_20991,N_20125);
or U21386 (N_21386,N_20540,N_20620);
nand U21387 (N_21387,N_20962,N_20199);
or U21388 (N_21388,N_20570,N_21027);
or U21389 (N_21389,N_20671,N_20467);
xnor U21390 (N_21390,N_20451,N_20258);
nand U21391 (N_21391,N_21206,N_20681);
xnor U21392 (N_21392,N_21041,N_20413);
nor U21393 (N_21393,N_20421,N_21191);
and U21394 (N_21394,N_21180,N_20029);
nor U21395 (N_21395,N_20983,N_20600);
or U21396 (N_21396,N_20037,N_20682);
xnor U21397 (N_21397,N_20433,N_20752);
xnor U21398 (N_21398,N_20486,N_20019);
and U21399 (N_21399,N_20811,N_20601);
or U21400 (N_21400,N_20819,N_20892);
and U21401 (N_21401,N_20736,N_20993);
xnor U21402 (N_21402,N_20643,N_20182);
xor U21403 (N_21403,N_21124,N_20491);
nor U21404 (N_21404,N_21105,N_21157);
nand U21405 (N_21405,N_21125,N_20239);
and U21406 (N_21406,N_20701,N_20465);
or U21407 (N_21407,N_20543,N_20689);
nor U21408 (N_21408,N_21246,N_20852);
xor U21409 (N_21409,N_21159,N_20012);
or U21410 (N_21410,N_20755,N_20666);
and U21411 (N_21411,N_20953,N_20944);
xor U21412 (N_21412,N_20366,N_20314);
xor U21413 (N_21413,N_20517,N_20709);
nor U21414 (N_21414,N_20524,N_20378);
nor U21415 (N_21415,N_20123,N_20165);
nand U21416 (N_21416,N_20934,N_20928);
and U21417 (N_21417,N_20310,N_20989);
nand U21418 (N_21418,N_20494,N_20026);
nor U21419 (N_21419,N_20630,N_20857);
or U21420 (N_21420,N_20943,N_20956);
xnor U21421 (N_21421,N_20196,N_21099);
nand U21422 (N_21422,N_20705,N_20972);
nor U21423 (N_21423,N_20990,N_20181);
nand U21424 (N_21424,N_20615,N_20386);
nor U21425 (N_21425,N_20138,N_20834);
nor U21426 (N_21426,N_20803,N_20428);
and U21427 (N_21427,N_20688,N_20368);
nor U21428 (N_21428,N_20317,N_20279);
xnor U21429 (N_21429,N_20148,N_20759);
nor U21430 (N_21430,N_20434,N_20392);
nand U21431 (N_21431,N_20516,N_20742);
nor U21432 (N_21432,N_20754,N_21208);
and U21433 (N_21433,N_20572,N_20741);
nor U21434 (N_21434,N_20995,N_20770);
nand U21435 (N_21435,N_21139,N_20492);
xor U21436 (N_21436,N_20566,N_21241);
xnor U21437 (N_21437,N_20198,N_20394);
nor U21438 (N_21438,N_20230,N_20678);
or U21439 (N_21439,N_20090,N_20312);
nor U21440 (N_21440,N_20599,N_20435);
or U21441 (N_21441,N_20903,N_20141);
and U21442 (N_21442,N_21050,N_20327);
xnor U21443 (N_21443,N_20161,N_20202);
nand U21444 (N_21444,N_20356,N_20409);
nor U21445 (N_21445,N_20556,N_20909);
nand U21446 (N_21446,N_20333,N_20416);
or U21447 (N_21447,N_20628,N_20782);
nor U21448 (N_21448,N_20850,N_21076);
nor U21449 (N_21449,N_20837,N_20487);
nand U21450 (N_21450,N_20417,N_20679);
nor U21451 (N_21451,N_20443,N_20329);
and U21452 (N_21452,N_20146,N_20374);
and U21453 (N_21453,N_21049,N_20363);
nor U21454 (N_21454,N_20805,N_20659);
xnor U21455 (N_21455,N_21154,N_21047);
xnor U21456 (N_21456,N_21106,N_20233);
and U21457 (N_21457,N_20906,N_21235);
nand U21458 (N_21458,N_20911,N_21025);
nor U21459 (N_21459,N_20457,N_20031);
xnor U21460 (N_21460,N_20128,N_20072);
nand U21461 (N_21461,N_20328,N_20050);
xnor U21462 (N_21462,N_20613,N_20235);
and U21463 (N_21463,N_20725,N_20440);
nor U21464 (N_21464,N_21080,N_20981);
nor U21465 (N_21465,N_21146,N_20481);
xnor U21466 (N_21466,N_21162,N_20136);
or U21467 (N_21467,N_20382,N_20041);
or U21468 (N_21468,N_20727,N_20024);
xor U21469 (N_21469,N_20240,N_20345);
and U21470 (N_21470,N_20206,N_21111);
nor U21471 (N_21471,N_21007,N_20814);
and U21472 (N_21472,N_20025,N_21115);
xor U21473 (N_21473,N_20895,N_20868);
xor U21474 (N_21474,N_21114,N_21051);
xnor U21475 (N_21475,N_21213,N_21122);
and U21476 (N_21476,N_20042,N_20664);
and U21477 (N_21477,N_20508,N_20756);
and U21478 (N_21478,N_20593,N_20711);
or U21479 (N_21479,N_20885,N_20323);
xor U21480 (N_21480,N_20054,N_20015);
xor U21481 (N_21481,N_20835,N_20377);
and U21482 (N_21482,N_20618,N_20271);
nand U21483 (N_21483,N_21129,N_21230);
or U21484 (N_21484,N_20101,N_21012);
and U21485 (N_21485,N_20255,N_20411);
xnor U21486 (N_21486,N_20924,N_20635);
xnor U21487 (N_21487,N_20912,N_20296);
nand U21488 (N_21488,N_20735,N_21017);
nand U21489 (N_21489,N_20642,N_20632);
or U21490 (N_21490,N_20557,N_20361);
or U21491 (N_21491,N_21155,N_21031);
or U21492 (N_21492,N_20096,N_20004);
and U21493 (N_21493,N_20761,N_20383);
nor U21494 (N_21494,N_21116,N_21190);
and U21495 (N_21495,N_20949,N_20750);
and U21496 (N_21496,N_20866,N_21089);
nand U21497 (N_21497,N_20896,N_20936);
xor U21498 (N_21498,N_20163,N_20794);
nand U21499 (N_21499,N_20714,N_21164);
nor U21500 (N_21500,N_20285,N_20424);
xor U21501 (N_21501,N_20619,N_20751);
or U21502 (N_21502,N_20629,N_21023);
xnor U21503 (N_21503,N_20114,N_20763);
or U21504 (N_21504,N_20131,N_20825);
xor U21505 (N_21505,N_20313,N_20208);
or U21506 (N_21506,N_20069,N_20355);
and U21507 (N_21507,N_20897,N_20888);
and U21508 (N_21508,N_20656,N_20661);
xnor U21509 (N_21509,N_20001,N_21185);
or U21510 (N_21510,N_20213,N_21210);
and U21511 (N_21511,N_20305,N_20552);
or U21512 (N_21512,N_21209,N_20343);
or U21513 (N_21513,N_20980,N_20055);
xnor U21514 (N_21514,N_20851,N_20444);
xnor U21515 (N_21515,N_20856,N_20445);
xnor U21516 (N_21516,N_21224,N_20308);
xor U21517 (N_21517,N_20799,N_20284);
and U21518 (N_21518,N_20715,N_20275);
xnor U21519 (N_21519,N_20446,N_20747);
or U21520 (N_21520,N_20554,N_20061);
or U21521 (N_21521,N_20321,N_21075);
nand U21522 (N_21522,N_20224,N_21128);
or U21523 (N_21523,N_20137,N_20553);
and U21524 (N_21524,N_20261,N_20108);
and U21525 (N_21525,N_20838,N_20332);
nand U21526 (N_21526,N_21038,N_20963);
or U21527 (N_21527,N_21090,N_20567);
nor U21528 (N_21528,N_20702,N_20423);
xnor U21529 (N_21529,N_20959,N_20587);
xor U21530 (N_21530,N_20623,N_21171);
and U21531 (N_21531,N_20607,N_20631);
nand U21532 (N_21532,N_20145,N_21141);
xnor U21533 (N_21533,N_20621,N_21245);
and U21534 (N_21534,N_20889,N_20293);
nand U21535 (N_21535,N_21081,N_20073);
xnor U21536 (N_21536,N_20160,N_20438);
nor U21537 (N_21537,N_20149,N_20930);
nor U21538 (N_21538,N_21145,N_21240);
nor U21539 (N_21539,N_20410,N_21220);
or U21540 (N_21540,N_20706,N_20578);
nand U21541 (N_21541,N_21083,N_20586);
nand U21542 (N_21542,N_21086,N_21087);
nand U21543 (N_21543,N_20873,N_20534);
and U21544 (N_21544,N_20961,N_20948);
and U21545 (N_21545,N_20674,N_20064);
or U21546 (N_21546,N_20560,N_20187);
or U21547 (N_21547,N_21223,N_20564);
xnor U21548 (N_21548,N_20614,N_20121);
and U21549 (N_21549,N_21035,N_20773);
nor U21550 (N_21550,N_21072,N_20667);
and U21551 (N_21551,N_20532,N_20931);
and U21552 (N_21552,N_20683,N_20823);
xor U21553 (N_21553,N_20412,N_20519);
or U21554 (N_21554,N_20300,N_20639);
xnor U21555 (N_21555,N_20191,N_20303);
nor U21556 (N_21556,N_21178,N_20062);
nand U21557 (N_21557,N_20908,N_20836);
or U21558 (N_21558,N_20152,N_21096);
and U21559 (N_21559,N_21060,N_21217);
or U21560 (N_21560,N_20937,N_21194);
and U21561 (N_21561,N_20060,N_20133);
xnor U21562 (N_21562,N_20790,N_20309);
nor U21563 (N_21563,N_20371,N_20893);
xor U21564 (N_21564,N_20625,N_20831);
or U21565 (N_21565,N_20017,N_20164);
nand U21566 (N_21566,N_20307,N_20458);
and U21567 (N_21567,N_20244,N_20192);
nor U21568 (N_21568,N_20518,N_20883);
or U21569 (N_21569,N_21053,N_20325);
nand U21570 (N_21570,N_20525,N_20845);
or U21571 (N_21571,N_20460,N_20140);
nor U21572 (N_21572,N_20783,N_20969);
nand U21573 (N_21573,N_21018,N_20929);
or U21574 (N_21574,N_21056,N_20166);
nor U21575 (N_21575,N_21123,N_20020);
and U21576 (N_21576,N_20051,N_20375);
or U21577 (N_21577,N_20942,N_20404);
and U21578 (N_21578,N_20111,N_21158);
nand U21579 (N_21579,N_20172,N_20117);
xnor U21580 (N_21580,N_20670,N_20626);
xnor U21581 (N_21581,N_20917,N_20316);
and U21582 (N_21582,N_20743,N_20746);
nor U21583 (N_21583,N_20507,N_20023);
nand U21584 (N_21584,N_20719,N_20870);
nor U21585 (N_21585,N_20387,N_21013);
nand U21586 (N_21586,N_20082,N_20846);
nor U21587 (N_21587,N_20466,N_20021);
or U21588 (N_21588,N_20504,N_20124);
nand U21589 (N_21589,N_20588,N_21042);
or U21590 (N_21590,N_20765,N_20008);
nor U21591 (N_21591,N_21048,N_21061);
and U21592 (N_21592,N_20018,N_21244);
nor U21593 (N_21593,N_20227,N_21071);
nor U21594 (N_21594,N_20462,N_20604);
nor U21595 (N_21595,N_20544,N_20776);
xnor U21596 (N_21596,N_20399,N_20690);
xnor U21597 (N_21597,N_20176,N_20817);
or U21598 (N_21598,N_20301,N_20186);
nand U21599 (N_21599,N_20351,N_20523);
xor U21600 (N_21600,N_21130,N_20985);
nor U21601 (N_21601,N_20596,N_21062);
nor U21602 (N_21602,N_20968,N_20648);
nand U21603 (N_21603,N_20359,N_20155);
nand U21604 (N_21604,N_20231,N_20988);
xnor U21605 (N_21605,N_20685,N_20036);
or U21606 (N_21606,N_21182,N_20463);
nor U21607 (N_21607,N_21100,N_20039);
nand U21608 (N_21608,N_21074,N_20254);
and U21609 (N_21609,N_20958,N_21103);
nor U21610 (N_21610,N_20966,N_20887);
nor U21611 (N_21611,N_20295,N_20000);
xnor U21612 (N_21612,N_20574,N_20536);
nor U21613 (N_21613,N_21175,N_20729);
nand U21614 (N_21614,N_20784,N_20449);
xor U21615 (N_21615,N_20011,N_20406);
nand U21616 (N_21616,N_20360,N_20084);
nand U21617 (N_21617,N_20606,N_20853);
or U21618 (N_21618,N_20143,N_20304);
and U21619 (N_21619,N_20986,N_20067);
xnor U21620 (N_21620,N_20718,N_20175);
nand U21621 (N_21621,N_20478,N_20075);
or U21622 (N_21622,N_20796,N_20372);
nand U21623 (N_21623,N_20527,N_21144);
or U21624 (N_21624,N_20653,N_20112);
and U21625 (N_21625,N_20640,N_21163);
xor U21626 (N_21626,N_20641,N_21192);
nand U21627 (N_21627,N_20298,N_20916);
and U21628 (N_21628,N_21044,N_20488);
nand U21629 (N_21629,N_20157,N_20228);
xor U21630 (N_21630,N_20158,N_20703);
or U21631 (N_21631,N_20282,N_20824);
and U21632 (N_21632,N_20730,N_20521);
or U21633 (N_21633,N_20698,N_20739);
or U21634 (N_21634,N_20162,N_20104);
or U21635 (N_21635,N_20470,N_20038);
xor U21636 (N_21636,N_20483,N_20130);
and U21637 (N_21637,N_20216,N_20081);
and U21638 (N_21638,N_20855,N_21079);
and U21639 (N_21639,N_20265,N_21058);
nor U21640 (N_21640,N_20068,N_20408);
or U21641 (N_21641,N_20091,N_20236);
nand U21642 (N_21642,N_20319,N_20997);
nor U21643 (N_21643,N_21069,N_20014);
or U21644 (N_21644,N_20215,N_21132);
or U21645 (N_21645,N_21233,N_21166);
nand U21646 (N_21646,N_21028,N_20259);
nand U21647 (N_21647,N_20221,N_20882);
and U21648 (N_21648,N_20195,N_21112);
nor U21649 (N_21649,N_20649,N_20419);
nand U21650 (N_21650,N_20563,N_20003);
nor U21651 (N_21651,N_20102,N_20745);
and U21652 (N_21652,N_21137,N_20294);
nor U21653 (N_21653,N_20592,N_20529);
nand U21654 (N_21654,N_20218,N_20005);
nand U21655 (N_21655,N_20841,N_20979);
xor U21656 (N_21656,N_20778,N_21138);
xor U21657 (N_21657,N_20212,N_20657);
xor U21658 (N_21658,N_20211,N_20344);
nand U21659 (N_21659,N_20740,N_20346);
and U21660 (N_21660,N_20447,N_21211);
or U21661 (N_21661,N_21101,N_21054);
and U21662 (N_21662,N_20414,N_20469);
nor U21663 (N_21663,N_21020,N_20193);
nor U21664 (N_21664,N_20032,N_20809);
nand U21665 (N_21665,N_20900,N_21187);
xnor U21666 (N_21666,N_20352,N_20203);
xor U21667 (N_21667,N_20053,N_20229);
xor U21668 (N_21668,N_20941,N_20511);
and U21669 (N_21669,N_21177,N_20722);
nor U21670 (N_21670,N_20762,N_20270);
nand U21671 (N_21671,N_20663,N_20744);
nor U21672 (N_21672,N_20712,N_20699);
nor U21673 (N_21673,N_20816,N_20357);
or U21674 (N_21674,N_20495,N_21127);
nor U21675 (N_21675,N_20700,N_21225);
xnor U21676 (N_21676,N_20975,N_20335);
and U21677 (N_21677,N_20802,N_20877);
and U21678 (N_21678,N_20611,N_20862);
or U21679 (N_21679,N_20168,N_20052);
nor U21680 (N_21680,N_20180,N_20687);
and U21681 (N_21681,N_20531,N_20350);
nor U21682 (N_21682,N_20839,N_20040);
and U21683 (N_21683,N_20099,N_21088);
nand U21684 (N_21684,N_20797,N_21238);
and U21685 (N_21685,N_20637,N_20500);
or U21686 (N_21686,N_20764,N_20891);
or U21687 (N_21687,N_20957,N_20238);
xnor U21688 (N_21688,N_20217,N_20945);
or U21689 (N_21689,N_20485,N_20589);
xor U21690 (N_21690,N_20726,N_20573);
nor U21691 (N_21691,N_20840,N_20723);
and U21692 (N_21692,N_21068,N_20616);
xnor U21693 (N_21693,N_20118,N_20919);
xnor U21694 (N_21694,N_20439,N_20496);
and U21695 (N_21695,N_20503,N_20473);
or U21696 (N_21696,N_20644,N_20528);
nand U21697 (N_21697,N_20076,N_21032);
nor U21698 (N_21698,N_21218,N_21198);
or U21699 (N_21699,N_20474,N_21063);
nor U21700 (N_21700,N_20184,N_20336);
and U21701 (N_21701,N_21043,N_20634);
xor U21702 (N_21702,N_20537,N_20448);
nand U21703 (N_21703,N_20156,N_21022);
nor U21704 (N_21704,N_20708,N_20734);
and U21705 (N_21705,N_20376,N_20358);
nand U21706 (N_21706,N_20872,N_21172);
or U21707 (N_21707,N_20455,N_20710);
nand U21708 (N_21708,N_20843,N_20505);
xor U21709 (N_21709,N_20260,N_20167);
nand U21710 (N_21710,N_20996,N_20334);
xor U21711 (N_21711,N_20509,N_20119);
and U21712 (N_21712,N_20684,N_20777);
and U21713 (N_21713,N_20169,N_20283);
nor U21714 (N_21714,N_20580,N_20070);
nor U21715 (N_21715,N_20369,N_21152);
and U21716 (N_21716,N_20058,N_20820);
and U21717 (N_21717,N_20952,N_21059);
or U21718 (N_21718,N_20110,N_20512);
nand U21719 (N_21719,N_20174,N_21227);
or U21720 (N_21720,N_20583,N_20341);
nand U21721 (N_21721,N_20364,N_21196);
xor U21722 (N_21722,N_20597,N_20429);
and U21723 (N_21723,N_20865,N_21174);
nor U21724 (N_21724,N_20871,N_21165);
nand U21725 (N_21725,N_20122,N_20526);
nor U21726 (N_21726,N_20603,N_21045);
and U21727 (N_21727,N_20472,N_20047);
nand U21728 (N_21728,N_20427,N_20951);
nor U21729 (N_21729,N_21037,N_20232);
and U21730 (N_21730,N_20297,N_20965);
or U21731 (N_21731,N_20609,N_20189);
nand U21732 (N_21732,N_20894,N_20562);
xnor U21733 (N_21733,N_21131,N_20848);
nand U21734 (N_21734,N_20881,N_20559);
nand U21735 (N_21735,N_21176,N_20584);
xnor U21736 (N_21736,N_21236,N_20913);
or U21737 (N_21737,N_20792,N_21082);
nor U21738 (N_21738,N_21173,N_20498);
and U21739 (N_21739,N_20127,N_21004);
nand U21740 (N_21740,N_20200,N_20978);
nand U21741 (N_21741,N_20045,N_21226);
nor U21742 (N_21742,N_20693,N_20113);
nor U21743 (N_21743,N_20080,N_20342);
or U21744 (N_21744,N_20940,N_20281);
nor U21745 (N_21745,N_21040,N_20436);
and U21746 (N_21746,N_21181,N_20828);
nand U21747 (N_21747,N_20549,N_20987);
or U21748 (N_21748,N_20256,N_20454);
or U21749 (N_21749,N_20278,N_20932);
nand U21750 (N_21750,N_20904,N_20672);
or U21751 (N_21751,N_20093,N_20697);
nand U21752 (N_21752,N_20353,N_20286);
xnor U21753 (N_21753,N_20252,N_20807);
or U21754 (N_21754,N_20384,N_20267);
nor U21755 (N_21755,N_21008,N_21121);
or U21756 (N_21756,N_21113,N_20338);
xor U21757 (N_21757,N_20801,N_20795);
nand U21758 (N_21758,N_20652,N_20134);
nand U21759 (N_21759,N_20431,N_20154);
nand U21760 (N_21760,N_20984,N_20490);
xnor U21761 (N_21761,N_20405,N_20009);
and U21762 (N_21762,N_20753,N_20774);
or U21763 (N_21763,N_20311,N_20716);
nor U21764 (N_21764,N_21207,N_20967);
or U21765 (N_21765,N_20915,N_20209);
xnor U21766 (N_21766,N_20468,N_20373);
nand U21767 (N_21767,N_20151,N_20733);
or U21768 (N_21768,N_20420,N_21170);
and U21769 (N_21769,N_20860,N_21234);
and U21770 (N_21770,N_20598,N_20083);
xnor U21771 (N_21771,N_21216,N_20407);
xnor U21772 (N_21772,N_20480,N_21016);
nand U21773 (N_21773,N_21057,N_21179);
xnor U21774 (N_21774,N_21000,N_21200);
nor U21775 (N_21775,N_20624,N_20561);
or U21776 (N_21776,N_20105,N_20976);
or U21777 (N_21777,N_20551,N_20898);
xor U21778 (N_21778,N_20815,N_21148);
xor U21779 (N_21779,N_20185,N_20223);
nand U21780 (N_21780,N_20243,N_21237);
and U21781 (N_21781,N_21184,N_20389);
xor U21782 (N_21782,N_20854,N_20775);
and U21783 (N_21783,N_20946,N_20677);
nor U21784 (N_21784,N_20226,N_20907);
nand U21785 (N_21785,N_20288,N_20430);
nor U21786 (N_21786,N_21110,N_20087);
or U21787 (N_21787,N_20142,N_20237);
xnor U21788 (N_21788,N_20576,N_20970);
nand U21789 (N_21789,N_20886,N_20135);
nor U21790 (N_21790,N_20289,N_21186);
xor U21791 (N_21791,N_20781,N_21094);
nor U21792 (N_21792,N_20249,N_20348);
nor U21793 (N_21793,N_20654,N_20059);
or U21794 (N_21794,N_20827,N_20863);
nand U21795 (N_21795,N_20542,N_20760);
xor U21796 (N_21796,N_20302,N_20676);
xor U21797 (N_21797,N_21065,N_20669);
and U21798 (N_21798,N_20204,N_20926);
nor U21799 (N_21799,N_20905,N_21248);
nand U21800 (N_21800,N_20675,N_21229);
nand U21801 (N_21801,N_20585,N_20362);
or U21802 (N_21802,N_20476,N_20214);
nor U21803 (N_21803,N_20982,N_20673);
and U21804 (N_21804,N_20779,N_20065);
nand U21805 (N_21805,N_20441,N_21118);
nor U21806 (N_21806,N_20066,N_20071);
nor U21807 (N_21807,N_20079,N_21243);
nand U21808 (N_21808,N_21093,N_20028);
nand U21809 (N_21809,N_20696,N_21228);
xnor U21810 (N_21810,N_20869,N_20299);
xor U21811 (N_21811,N_20272,N_21133);
nor U21812 (N_21812,N_20691,N_21212);
xor U21813 (N_21813,N_20558,N_20178);
nor U21814 (N_21814,N_20513,N_20680);
nor U21815 (N_21815,N_20879,N_21215);
nor U21816 (N_21816,N_21197,N_20633);
or U21817 (N_21817,N_20798,N_20720);
nand U21818 (N_21818,N_21078,N_20418);
nor U21819 (N_21819,N_21085,N_20546);
or U21820 (N_21820,N_21153,N_21019);
or U21821 (N_21821,N_20867,N_21097);
nor U21822 (N_21822,N_20450,N_20550);
nand U21823 (N_21823,N_20034,N_20541);
nand U21824 (N_21824,N_21033,N_20046);
or U21825 (N_21825,N_20103,N_20291);
nand U21826 (N_21826,N_20992,N_20246);
nand U21827 (N_21827,N_20100,N_20595);
nor U21828 (N_21828,N_20150,N_21092);
and U21829 (N_21829,N_20858,N_20571);
and U21830 (N_21830,N_20627,N_20501);
or U21831 (N_21831,N_21001,N_20660);
or U21832 (N_21832,N_20826,N_21201);
and U21833 (N_21833,N_20337,N_20048);
and U21834 (N_21834,N_20921,N_21055);
nand U21835 (N_21835,N_21009,N_21161);
or U21836 (N_21836,N_20044,N_20385);
nor U21837 (N_21837,N_20347,N_20646);
xnor U21838 (N_21838,N_20998,N_20847);
nor U21839 (N_21839,N_20397,N_20582);
xnor U21840 (N_21840,N_20425,N_20568);
nor U21841 (N_21841,N_21204,N_20273);
nand U21842 (N_21842,N_20401,N_20994);
nor U21843 (N_21843,N_20732,N_20030);
nand U21844 (N_21844,N_20821,N_20622);
nor U21845 (N_21845,N_21036,N_20432);
xor U21846 (N_21846,N_20922,N_20864);
nor U21847 (N_21847,N_20806,N_20539);
nor U21848 (N_21848,N_20522,N_20638);
xor U21849 (N_21849,N_20159,N_21119);
and U21850 (N_21850,N_20129,N_21147);
nand U21851 (N_21851,N_20594,N_20264);
nor U21852 (N_21852,N_20923,N_20668);
or U21853 (N_21853,N_20955,N_21202);
nor U21854 (N_21854,N_20787,N_20939);
xnor U21855 (N_21855,N_21242,N_21231);
or U21856 (N_21856,N_20016,N_20780);
or U21857 (N_21857,N_20731,N_21010);
xnor U21858 (N_21858,N_20225,N_20253);
nor U21859 (N_21859,N_20027,N_21024);
and U21860 (N_21860,N_20391,N_20002);
or U21861 (N_21861,N_20459,N_20475);
xor U21862 (N_21862,N_20290,N_20579);
xnor U21863 (N_21863,N_20320,N_20247);
or U21864 (N_21864,N_20960,N_20793);
nor U21865 (N_21865,N_20415,N_20788);
and U21866 (N_21866,N_20349,N_20651);
or U21867 (N_21867,N_20808,N_21126);
xor U21868 (N_21868,N_20330,N_21011);
nand U21869 (N_21869,N_21021,N_20057);
xor U21870 (N_21870,N_20098,N_20938);
or U21871 (N_21871,N_20515,N_20662);
xor U21872 (N_21872,N_20704,N_20692);
xnor U21873 (N_21873,N_20999,N_21221);
nor U21874 (N_21874,N_20107,N_21070);
or U21875 (N_21875,N_20333,N_21128);
or U21876 (N_21876,N_20688,N_20823);
or U21877 (N_21877,N_20965,N_20086);
or U21878 (N_21878,N_20383,N_20578);
and U21879 (N_21879,N_20626,N_20497);
nand U21880 (N_21880,N_20083,N_20635);
xor U21881 (N_21881,N_21122,N_20269);
and U21882 (N_21882,N_21070,N_21078);
xnor U21883 (N_21883,N_20699,N_20569);
nor U21884 (N_21884,N_20819,N_20981);
and U21885 (N_21885,N_20042,N_21123);
or U21886 (N_21886,N_20876,N_20100);
xor U21887 (N_21887,N_20223,N_20459);
xor U21888 (N_21888,N_21014,N_20788);
or U21889 (N_21889,N_20980,N_21016);
and U21890 (N_21890,N_20276,N_20110);
nor U21891 (N_21891,N_20048,N_20933);
nand U21892 (N_21892,N_20476,N_20262);
xnor U21893 (N_21893,N_20053,N_21042);
or U21894 (N_21894,N_20240,N_20919);
and U21895 (N_21895,N_20582,N_20495);
nor U21896 (N_21896,N_20609,N_20993);
xor U21897 (N_21897,N_20834,N_20238);
nor U21898 (N_21898,N_20733,N_20723);
nand U21899 (N_21899,N_20064,N_20145);
or U21900 (N_21900,N_20485,N_20491);
nand U21901 (N_21901,N_21023,N_20599);
and U21902 (N_21902,N_20311,N_20435);
or U21903 (N_21903,N_20457,N_20040);
xnor U21904 (N_21904,N_20895,N_20905);
nor U21905 (N_21905,N_20099,N_20594);
or U21906 (N_21906,N_20823,N_21126);
nand U21907 (N_21907,N_20429,N_20230);
nand U21908 (N_21908,N_20862,N_20394);
and U21909 (N_21909,N_21089,N_20817);
xor U21910 (N_21910,N_20315,N_20248);
nand U21911 (N_21911,N_20309,N_20443);
nor U21912 (N_21912,N_21136,N_20336);
or U21913 (N_21913,N_20346,N_20958);
and U21914 (N_21914,N_20773,N_20838);
xor U21915 (N_21915,N_20936,N_20712);
nor U21916 (N_21916,N_20328,N_20940);
xor U21917 (N_21917,N_20874,N_20858);
nand U21918 (N_21918,N_20501,N_20849);
nand U21919 (N_21919,N_20907,N_20437);
or U21920 (N_21920,N_20171,N_20462);
or U21921 (N_21921,N_20273,N_20467);
xor U21922 (N_21922,N_20370,N_21044);
nor U21923 (N_21923,N_20751,N_20825);
or U21924 (N_21924,N_20494,N_20387);
nor U21925 (N_21925,N_20048,N_21157);
nor U21926 (N_21926,N_20048,N_20173);
xnor U21927 (N_21927,N_20448,N_20819);
and U21928 (N_21928,N_20337,N_20003);
nand U21929 (N_21929,N_20054,N_21116);
and U21930 (N_21930,N_20947,N_20030);
or U21931 (N_21931,N_20949,N_20369);
nand U21932 (N_21932,N_20746,N_20436);
and U21933 (N_21933,N_21249,N_20155);
nand U21934 (N_21934,N_21084,N_20577);
nor U21935 (N_21935,N_20891,N_20926);
and U21936 (N_21936,N_20898,N_20003);
and U21937 (N_21937,N_20128,N_20655);
and U21938 (N_21938,N_20399,N_20432);
or U21939 (N_21939,N_21084,N_21076);
and U21940 (N_21940,N_20775,N_20021);
and U21941 (N_21941,N_21059,N_20368);
nor U21942 (N_21942,N_21136,N_20908);
and U21943 (N_21943,N_20024,N_20579);
and U21944 (N_21944,N_20710,N_20635);
nor U21945 (N_21945,N_21077,N_20402);
and U21946 (N_21946,N_20982,N_20776);
nor U21947 (N_21947,N_20897,N_20782);
nand U21948 (N_21948,N_20214,N_20207);
nor U21949 (N_21949,N_21032,N_20166);
or U21950 (N_21950,N_20921,N_20017);
nand U21951 (N_21951,N_20158,N_20351);
nand U21952 (N_21952,N_21181,N_21241);
or U21953 (N_21953,N_20233,N_20349);
nand U21954 (N_21954,N_21229,N_20411);
nand U21955 (N_21955,N_21171,N_20417);
nor U21956 (N_21956,N_20365,N_20393);
nand U21957 (N_21957,N_20146,N_21022);
nand U21958 (N_21958,N_20753,N_20572);
nand U21959 (N_21959,N_20116,N_20636);
xnor U21960 (N_21960,N_21219,N_21135);
or U21961 (N_21961,N_20125,N_20090);
nor U21962 (N_21962,N_21206,N_20954);
xnor U21963 (N_21963,N_20232,N_20161);
nand U21964 (N_21964,N_20197,N_20927);
xor U21965 (N_21965,N_21171,N_20099);
and U21966 (N_21966,N_20694,N_20343);
and U21967 (N_21967,N_20267,N_20953);
xor U21968 (N_21968,N_20454,N_20115);
or U21969 (N_21969,N_20049,N_21009);
or U21970 (N_21970,N_21074,N_20875);
and U21971 (N_21971,N_20296,N_20193);
nor U21972 (N_21972,N_20132,N_20352);
and U21973 (N_21973,N_21147,N_21077);
or U21974 (N_21974,N_20907,N_20939);
xnor U21975 (N_21975,N_20342,N_20556);
and U21976 (N_21976,N_20955,N_20644);
xor U21977 (N_21977,N_20766,N_20026);
and U21978 (N_21978,N_21033,N_20977);
nor U21979 (N_21979,N_20184,N_20127);
xnor U21980 (N_21980,N_20237,N_20666);
nand U21981 (N_21981,N_21042,N_20940);
nor U21982 (N_21982,N_20423,N_20289);
or U21983 (N_21983,N_20252,N_21185);
nand U21984 (N_21984,N_20865,N_21223);
xor U21985 (N_21985,N_20522,N_20889);
xor U21986 (N_21986,N_21042,N_21150);
nand U21987 (N_21987,N_20858,N_20523);
xnor U21988 (N_21988,N_20550,N_21095);
or U21989 (N_21989,N_20485,N_20137);
nand U21990 (N_21990,N_20844,N_21150);
nand U21991 (N_21991,N_20800,N_20515);
or U21992 (N_21992,N_20092,N_20536);
xnor U21993 (N_21993,N_20775,N_20487);
nand U21994 (N_21994,N_20470,N_20364);
nand U21995 (N_21995,N_20588,N_20767);
or U21996 (N_21996,N_20644,N_20293);
nor U21997 (N_21997,N_20334,N_20795);
nor U21998 (N_21998,N_20216,N_20982);
or U21999 (N_21999,N_20886,N_20709);
nor U22000 (N_22000,N_20739,N_20582);
nor U22001 (N_22001,N_20976,N_20999);
and U22002 (N_22002,N_20969,N_20852);
or U22003 (N_22003,N_20411,N_20652);
nor U22004 (N_22004,N_21102,N_20034);
or U22005 (N_22005,N_20585,N_20242);
nand U22006 (N_22006,N_21047,N_20630);
nor U22007 (N_22007,N_20554,N_20071);
xor U22008 (N_22008,N_21159,N_20835);
xor U22009 (N_22009,N_20660,N_20904);
xnor U22010 (N_22010,N_20829,N_20678);
nor U22011 (N_22011,N_21092,N_20575);
and U22012 (N_22012,N_20307,N_20839);
nand U22013 (N_22013,N_20511,N_20256);
xor U22014 (N_22014,N_20876,N_20874);
nand U22015 (N_22015,N_20777,N_20755);
and U22016 (N_22016,N_20798,N_20195);
xor U22017 (N_22017,N_21032,N_20606);
xor U22018 (N_22018,N_20420,N_20070);
nand U22019 (N_22019,N_21015,N_21152);
or U22020 (N_22020,N_20257,N_21156);
nand U22021 (N_22021,N_20511,N_20043);
or U22022 (N_22022,N_20300,N_20766);
xnor U22023 (N_22023,N_21146,N_20383);
nor U22024 (N_22024,N_20244,N_20753);
and U22025 (N_22025,N_20764,N_20546);
nor U22026 (N_22026,N_20939,N_20000);
nor U22027 (N_22027,N_20594,N_21245);
or U22028 (N_22028,N_20445,N_20179);
nand U22029 (N_22029,N_21225,N_20666);
and U22030 (N_22030,N_20602,N_20393);
nand U22031 (N_22031,N_20499,N_20452);
xor U22032 (N_22032,N_20944,N_20554);
or U22033 (N_22033,N_20828,N_20685);
xor U22034 (N_22034,N_20901,N_20710);
xnor U22035 (N_22035,N_21196,N_20691);
nand U22036 (N_22036,N_20537,N_20617);
or U22037 (N_22037,N_20215,N_20874);
or U22038 (N_22038,N_20647,N_21049);
xnor U22039 (N_22039,N_20221,N_20512);
xnor U22040 (N_22040,N_21184,N_20802);
or U22041 (N_22041,N_20091,N_20010);
or U22042 (N_22042,N_20028,N_20128);
nor U22043 (N_22043,N_21099,N_20419);
xor U22044 (N_22044,N_21061,N_20681);
xor U22045 (N_22045,N_20791,N_21175);
or U22046 (N_22046,N_20884,N_20618);
nand U22047 (N_22047,N_20049,N_20583);
and U22048 (N_22048,N_21175,N_20351);
or U22049 (N_22049,N_20829,N_20609);
nor U22050 (N_22050,N_20073,N_20601);
and U22051 (N_22051,N_21040,N_20804);
nor U22052 (N_22052,N_21046,N_20524);
nor U22053 (N_22053,N_20441,N_20069);
and U22054 (N_22054,N_20054,N_20485);
and U22055 (N_22055,N_20692,N_20001);
nand U22056 (N_22056,N_20062,N_20749);
nor U22057 (N_22057,N_20842,N_21160);
nor U22058 (N_22058,N_20645,N_20749);
and U22059 (N_22059,N_20437,N_20720);
and U22060 (N_22060,N_20340,N_20383);
and U22061 (N_22061,N_20904,N_21177);
or U22062 (N_22062,N_20491,N_20068);
xor U22063 (N_22063,N_20918,N_21067);
nor U22064 (N_22064,N_20597,N_20149);
and U22065 (N_22065,N_20133,N_20930);
xnor U22066 (N_22066,N_20175,N_20274);
xnor U22067 (N_22067,N_21199,N_20465);
and U22068 (N_22068,N_20531,N_20797);
or U22069 (N_22069,N_20584,N_20395);
nor U22070 (N_22070,N_20263,N_20864);
and U22071 (N_22071,N_20769,N_20333);
nor U22072 (N_22072,N_20076,N_21243);
xnor U22073 (N_22073,N_21112,N_20485);
xnor U22074 (N_22074,N_20219,N_21052);
nor U22075 (N_22075,N_20050,N_20329);
and U22076 (N_22076,N_21072,N_20378);
and U22077 (N_22077,N_21048,N_20158);
xnor U22078 (N_22078,N_20769,N_20364);
or U22079 (N_22079,N_21049,N_20665);
or U22080 (N_22080,N_20409,N_20505);
nor U22081 (N_22081,N_21003,N_21033);
nor U22082 (N_22082,N_20568,N_20935);
nor U22083 (N_22083,N_20601,N_20733);
nor U22084 (N_22084,N_20176,N_20882);
xnor U22085 (N_22085,N_20876,N_20748);
xor U22086 (N_22086,N_20448,N_20208);
nand U22087 (N_22087,N_21195,N_21043);
xnor U22088 (N_22088,N_21006,N_20321);
xnor U22089 (N_22089,N_20257,N_20513);
or U22090 (N_22090,N_20683,N_20348);
nand U22091 (N_22091,N_20365,N_21047);
or U22092 (N_22092,N_20376,N_21025);
xor U22093 (N_22093,N_21224,N_20539);
and U22094 (N_22094,N_20414,N_20666);
xor U22095 (N_22095,N_20315,N_20096);
nor U22096 (N_22096,N_20742,N_20508);
nand U22097 (N_22097,N_20076,N_20664);
and U22098 (N_22098,N_20881,N_20140);
or U22099 (N_22099,N_20774,N_20821);
nor U22100 (N_22100,N_20197,N_20060);
nor U22101 (N_22101,N_20237,N_20646);
nor U22102 (N_22102,N_20162,N_20117);
and U22103 (N_22103,N_20769,N_20669);
or U22104 (N_22104,N_20036,N_20357);
and U22105 (N_22105,N_20065,N_20637);
xnor U22106 (N_22106,N_21086,N_21138);
or U22107 (N_22107,N_21079,N_21177);
xor U22108 (N_22108,N_20815,N_20368);
nand U22109 (N_22109,N_20311,N_20117);
nand U22110 (N_22110,N_20752,N_21001);
xor U22111 (N_22111,N_20646,N_20980);
or U22112 (N_22112,N_20302,N_20926);
or U22113 (N_22113,N_21221,N_20781);
xor U22114 (N_22114,N_20620,N_20392);
or U22115 (N_22115,N_20593,N_20386);
or U22116 (N_22116,N_20265,N_20375);
nand U22117 (N_22117,N_20258,N_20735);
or U22118 (N_22118,N_20119,N_20482);
nand U22119 (N_22119,N_20048,N_20788);
or U22120 (N_22120,N_21083,N_20696);
and U22121 (N_22121,N_20087,N_20567);
nor U22122 (N_22122,N_20168,N_20829);
nand U22123 (N_22123,N_20318,N_20575);
or U22124 (N_22124,N_20805,N_20314);
and U22125 (N_22125,N_21102,N_20075);
xor U22126 (N_22126,N_20960,N_20067);
or U22127 (N_22127,N_20764,N_20498);
xnor U22128 (N_22128,N_20210,N_20611);
and U22129 (N_22129,N_20874,N_20044);
xnor U22130 (N_22130,N_20224,N_21155);
xnor U22131 (N_22131,N_20286,N_20058);
nand U22132 (N_22132,N_21113,N_21086);
and U22133 (N_22133,N_20995,N_20454);
nand U22134 (N_22134,N_20014,N_20807);
nor U22135 (N_22135,N_20370,N_20065);
nand U22136 (N_22136,N_21238,N_21002);
xor U22137 (N_22137,N_21107,N_20973);
xnor U22138 (N_22138,N_20473,N_20812);
nand U22139 (N_22139,N_21169,N_20843);
and U22140 (N_22140,N_20791,N_20505);
nand U22141 (N_22141,N_20599,N_20057);
or U22142 (N_22142,N_20874,N_20742);
or U22143 (N_22143,N_20037,N_20325);
and U22144 (N_22144,N_20368,N_20976);
nor U22145 (N_22145,N_20060,N_20372);
nor U22146 (N_22146,N_20209,N_20588);
and U22147 (N_22147,N_20807,N_20272);
nor U22148 (N_22148,N_20767,N_21011);
and U22149 (N_22149,N_20444,N_20533);
or U22150 (N_22150,N_20432,N_21173);
xor U22151 (N_22151,N_20388,N_20308);
nor U22152 (N_22152,N_20023,N_20888);
and U22153 (N_22153,N_20242,N_21236);
and U22154 (N_22154,N_20828,N_20467);
or U22155 (N_22155,N_21201,N_20979);
nor U22156 (N_22156,N_21088,N_20921);
nand U22157 (N_22157,N_21223,N_20643);
or U22158 (N_22158,N_20358,N_21028);
nand U22159 (N_22159,N_20937,N_20021);
xor U22160 (N_22160,N_20706,N_20674);
nand U22161 (N_22161,N_20275,N_20661);
nor U22162 (N_22162,N_20169,N_20563);
xnor U22163 (N_22163,N_20660,N_20085);
or U22164 (N_22164,N_20967,N_20541);
and U22165 (N_22165,N_21196,N_20156);
and U22166 (N_22166,N_21123,N_20268);
xnor U22167 (N_22167,N_20755,N_20530);
or U22168 (N_22168,N_20103,N_20437);
xnor U22169 (N_22169,N_20577,N_20673);
and U22170 (N_22170,N_20094,N_20175);
nand U22171 (N_22171,N_20488,N_20719);
xor U22172 (N_22172,N_21137,N_20827);
and U22173 (N_22173,N_20720,N_20612);
xnor U22174 (N_22174,N_20005,N_20156);
nand U22175 (N_22175,N_20934,N_20105);
and U22176 (N_22176,N_20581,N_20021);
nor U22177 (N_22177,N_20105,N_20860);
or U22178 (N_22178,N_21201,N_21008);
and U22179 (N_22179,N_21066,N_20228);
or U22180 (N_22180,N_21221,N_20037);
nor U22181 (N_22181,N_20434,N_20967);
xnor U22182 (N_22182,N_21162,N_20826);
and U22183 (N_22183,N_20568,N_20327);
and U22184 (N_22184,N_20946,N_21208);
or U22185 (N_22185,N_20998,N_20338);
nand U22186 (N_22186,N_20506,N_20579);
nand U22187 (N_22187,N_21225,N_20373);
nand U22188 (N_22188,N_20756,N_20136);
nor U22189 (N_22189,N_20320,N_20184);
nand U22190 (N_22190,N_20193,N_20908);
and U22191 (N_22191,N_20807,N_20039);
nand U22192 (N_22192,N_20063,N_20106);
or U22193 (N_22193,N_20408,N_20098);
or U22194 (N_22194,N_20545,N_20547);
or U22195 (N_22195,N_21211,N_20139);
or U22196 (N_22196,N_20357,N_20660);
and U22197 (N_22197,N_20129,N_21101);
or U22198 (N_22198,N_20229,N_21249);
or U22199 (N_22199,N_20703,N_21171);
or U22200 (N_22200,N_20627,N_20440);
nor U22201 (N_22201,N_21085,N_20985);
and U22202 (N_22202,N_20183,N_20240);
xor U22203 (N_22203,N_20062,N_21225);
and U22204 (N_22204,N_21245,N_20756);
nor U22205 (N_22205,N_20188,N_20013);
nand U22206 (N_22206,N_21224,N_20117);
nor U22207 (N_22207,N_20069,N_20433);
nand U22208 (N_22208,N_20610,N_20160);
nand U22209 (N_22209,N_20136,N_20420);
xor U22210 (N_22210,N_20988,N_20670);
or U22211 (N_22211,N_20504,N_21158);
nor U22212 (N_22212,N_20618,N_20564);
and U22213 (N_22213,N_20062,N_21235);
and U22214 (N_22214,N_20562,N_20516);
nor U22215 (N_22215,N_21106,N_20461);
xnor U22216 (N_22216,N_20685,N_20197);
or U22217 (N_22217,N_20882,N_20018);
nor U22218 (N_22218,N_21055,N_20091);
xnor U22219 (N_22219,N_21047,N_20401);
and U22220 (N_22220,N_21156,N_20222);
or U22221 (N_22221,N_20243,N_20598);
xnor U22222 (N_22222,N_20625,N_20608);
nand U22223 (N_22223,N_20325,N_20657);
nor U22224 (N_22224,N_20971,N_20564);
xor U22225 (N_22225,N_20852,N_20494);
nor U22226 (N_22226,N_20243,N_20265);
and U22227 (N_22227,N_20839,N_20572);
xnor U22228 (N_22228,N_20027,N_20511);
nor U22229 (N_22229,N_20254,N_20173);
xor U22230 (N_22230,N_20624,N_20676);
nand U22231 (N_22231,N_20153,N_21039);
or U22232 (N_22232,N_20688,N_21194);
and U22233 (N_22233,N_20224,N_20804);
or U22234 (N_22234,N_21101,N_20712);
nor U22235 (N_22235,N_21098,N_21160);
and U22236 (N_22236,N_20746,N_21154);
xnor U22237 (N_22237,N_20595,N_20245);
nand U22238 (N_22238,N_20458,N_20531);
xor U22239 (N_22239,N_20348,N_20984);
and U22240 (N_22240,N_20599,N_20899);
or U22241 (N_22241,N_20708,N_20079);
or U22242 (N_22242,N_21233,N_20616);
and U22243 (N_22243,N_20968,N_20601);
and U22244 (N_22244,N_20844,N_20030);
nor U22245 (N_22245,N_21113,N_20186);
nor U22246 (N_22246,N_21145,N_20381);
and U22247 (N_22247,N_20152,N_20767);
or U22248 (N_22248,N_20101,N_20647);
nand U22249 (N_22249,N_21027,N_20790);
or U22250 (N_22250,N_20117,N_20188);
nand U22251 (N_22251,N_20377,N_20305);
or U22252 (N_22252,N_20287,N_21152);
xnor U22253 (N_22253,N_20864,N_20776);
nor U22254 (N_22254,N_20878,N_20834);
nand U22255 (N_22255,N_20242,N_20854);
nand U22256 (N_22256,N_20583,N_20520);
and U22257 (N_22257,N_20077,N_20675);
xor U22258 (N_22258,N_21169,N_20547);
xor U22259 (N_22259,N_20461,N_20028);
and U22260 (N_22260,N_20768,N_20961);
nor U22261 (N_22261,N_20240,N_20632);
or U22262 (N_22262,N_21184,N_20028);
and U22263 (N_22263,N_20120,N_20316);
xor U22264 (N_22264,N_20824,N_20349);
nand U22265 (N_22265,N_21173,N_21134);
nand U22266 (N_22266,N_20664,N_20996);
xor U22267 (N_22267,N_21045,N_21144);
and U22268 (N_22268,N_20981,N_20239);
and U22269 (N_22269,N_20706,N_20317);
xnor U22270 (N_22270,N_20594,N_20377);
and U22271 (N_22271,N_20683,N_20954);
and U22272 (N_22272,N_20050,N_20092);
xnor U22273 (N_22273,N_20533,N_21098);
or U22274 (N_22274,N_20377,N_20593);
xor U22275 (N_22275,N_20416,N_20291);
xor U22276 (N_22276,N_20922,N_20127);
nor U22277 (N_22277,N_20191,N_21148);
xnor U22278 (N_22278,N_20967,N_20972);
xor U22279 (N_22279,N_20155,N_20848);
nand U22280 (N_22280,N_20364,N_20301);
and U22281 (N_22281,N_20197,N_20819);
xor U22282 (N_22282,N_20573,N_20992);
and U22283 (N_22283,N_20035,N_20239);
or U22284 (N_22284,N_20308,N_20608);
nand U22285 (N_22285,N_20738,N_21231);
nor U22286 (N_22286,N_20423,N_20092);
or U22287 (N_22287,N_20294,N_20979);
nor U22288 (N_22288,N_21050,N_20431);
xnor U22289 (N_22289,N_20411,N_20338);
xnor U22290 (N_22290,N_21045,N_20978);
nand U22291 (N_22291,N_20580,N_20160);
nor U22292 (N_22292,N_21150,N_21154);
xnor U22293 (N_22293,N_21176,N_20142);
or U22294 (N_22294,N_21059,N_20528);
and U22295 (N_22295,N_20206,N_20281);
or U22296 (N_22296,N_20861,N_20149);
nor U22297 (N_22297,N_20855,N_20284);
xor U22298 (N_22298,N_21117,N_20103);
nand U22299 (N_22299,N_21195,N_20862);
xor U22300 (N_22300,N_20882,N_20975);
or U22301 (N_22301,N_20349,N_20327);
nor U22302 (N_22302,N_21052,N_20957);
xor U22303 (N_22303,N_20214,N_21011);
nand U22304 (N_22304,N_21019,N_20088);
xnor U22305 (N_22305,N_20610,N_21106);
and U22306 (N_22306,N_20950,N_20637);
and U22307 (N_22307,N_20627,N_20165);
nor U22308 (N_22308,N_20877,N_21052);
nor U22309 (N_22309,N_21089,N_20194);
nand U22310 (N_22310,N_21155,N_21136);
nor U22311 (N_22311,N_20636,N_20315);
nor U22312 (N_22312,N_20838,N_20915);
or U22313 (N_22313,N_20709,N_20130);
or U22314 (N_22314,N_20176,N_20071);
or U22315 (N_22315,N_21085,N_21113);
or U22316 (N_22316,N_21153,N_20001);
xor U22317 (N_22317,N_20784,N_20882);
or U22318 (N_22318,N_20162,N_20089);
and U22319 (N_22319,N_20454,N_20887);
nor U22320 (N_22320,N_20036,N_20870);
xnor U22321 (N_22321,N_20283,N_20322);
nand U22322 (N_22322,N_20118,N_20897);
and U22323 (N_22323,N_21084,N_20110);
or U22324 (N_22324,N_20331,N_20066);
nor U22325 (N_22325,N_20628,N_20899);
xor U22326 (N_22326,N_20361,N_20694);
nand U22327 (N_22327,N_20495,N_20510);
nand U22328 (N_22328,N_20506,N_20335);
nand U22329 (N_22329,N_20306,N_20305);
or U22330 (N_22330,N_20949,N_20839);
or U22331 (N_22331,N_20671,N_20979);
xor U22332 (N_22332,N_20670,N_21092);
nor U22333 (N_22333,N_20610,N_21010);
xnor U22334 (N_22334,N_20833,N_20595);
nand U22335 (N_22335,N_21245,N_20870);
xor U22336 (N_22336,N_20997,N_20657);
nor U22337 (N_22337,N_20825,N_20114);
xor U22338 (N_22338,N_20154,N_20450);
and U22339 (N_22339,N_20111,N_20509);
nand U22340 (N_22340,N_20755,N_21150);
nor U22341 (N_22341,N_20949,N_20164);
and U22342 (N_22342,N_20012,N_20421);
and U22343 (N_22343,N_20589,N_20206);
xnor U22344 (N_22344,N_20587,N_20297);
nor U22345 (N_22345,N_20380,N_20979);
and U22346 (N_22346,N_21150,N_20606);
and U22347 (N_22347,N_20052,N_20572);
or U22348 (N_22348,N_20471,N_20876);
nand U22349 (N_22349,N_20093,N_20149);
xnor U22350 (N_22350,N_20487,N_20812);
and U22351 (N_22351,N_20621,N_21136);
or U22352 (N_22352,N_21162,N_21219);
xnor U22353 (N_22353,N_21247,N_20730);
or U22354 (N_22354,N_21161,N_20700);
nor U22355 (N_22355,N_21104,N_20504);
xor U22356 (N_22356,N_21041,N_21035);
or U22357 (N_22357,N_20309,N_20678);
or U22358 (N_22358,N_20299,N_20080);
or U22359 (N_22359,N_20165,N_20182);
or U22360 (N_22360,N_20238,N_20409);
xor U22361 (N_22361,N_21155,N_20477);
nor U22362 (N_22362,N_20887,N_20494);
nand U22363 (N_22363,N_20452,N_21166);
and U22364 (N_22364,N_20910,N_21183);
nor U22365 (N_22365,N_20945,N_21070);
or U22366 (N_22366,N_20025,N_20044);
or U22367 (N_22367,N_20622,N_20372);
xor U22368 (N_22368,N_21190,N_20278);
nand U22369 (N_22369,N_21032,N_20396);
and U22370 (N_22370,N_21244,N_21066);
nor U22371 (N_22371,N_21222,N_20171);
nand U22372 (N_22372,N_20247,N_20719);
xnor U22373 (N_22373,N_20484,N_21205);
or U22374 (N_22374,N_21060,N_20652);
nand U22375 (N_22375,N_20018,N_20707);
nand U22376 (N_22376,N_20585,N_21112);
or U22377 (N_22377,N_20118,N_20080);
or U22378 (N_22378,N_21001,N_21040);
nor U22379 (N_22379,N_20142,N_20830);
and U22380 (N_22380,N_21087,N_20437);
or U22381 (N_22381,N_20220,N_20230);
or U22382 (N_22382,N_20288,N_20066);
or U22383 (N_22383,N_20777,N_20010);
or U22384 (N_22384,N_20800,N_20770);
or U22385 (N_22385,N_20685,N_20248);
nor U22386 (N_22386,N_21168,N_20775);
and U22387 (N_22387,N_21044,N_21081);
and U22388 (N_22388,N_20636,N_20924);
xnor U22389 (N_22389,N_21206,N_20154);
xnor U22390 (N_22390,N_20753,N_21024);
nor U22391 (N_22391,N_20653,N_21008);
nand U22392 (N_22392,N_20708,N_20656);
and U22393 (N_22393,N_21014,N_20561);
or U22394 (N_22394,N_20812,N_20711);
xnor U22395 (N_22395,N_21105,N_20131);
nor U22396 (N_22396,N_20525,N_21033);
and U22397 (N_22397,N_20228,N_20267);
and U22398 (N_22398,N_20141,N_20933);
xnor U22399 (N_22399,N_20680,N_20345);
nor U22400 (N_22400,N_20869,N_20373);
xor U22401 (N_22401,N_21150,N_21003);
or U22402 (N_22402,N_20792,N_20697);
and U22403 (N_22403,N_21217,N_20061);
nand U22404 (N_22404,N_20300,N_20644);
xor U22405 (N_22405,N_21108,N_20640);
or U22406 (N_22406,N_20090,N_21126);
nand U22407 (N_22407,N_21069,N_20324);
nor U22408 (N_22408,N_20396,N_20181);
nand U22409 (N_22409,N_20253,N_21091);
or U22410 (N_22410,N_21233,N_20300);
xor U22411 (N_22411,N_20788,N_20454);
nor U22412 (N_22412,N_20361,N_21017);
or U22413 (N_22413,N_20107,N_20316);
xor U22414 (N_22414,N_20425,N_21051);
or U22415 (N_22415,N_20920,N_20187);
xnor U22416 (N_22416,N_20218,N_21129);
nand U22417 (N_22417,N_20703,N_20267);
xor U22418 (N_22418,N_21119,N_21185);
nor U22419 (N_22419,N_20433,N_20420);
xor U22420 (N_22420,N_20020,N_20310);
or U22421 (N_22421,N_21153,N_20749);
or U22422 (N_22422,N_20543,N_20497);
and U22423 (N_22423,N_20497,N_21091);
nand U22424 (N_22424,N_20155,N_20989);
or U22425 (N_22425,N_20696,N_20543);
nor U22426 (N_22426,N_20785,N_20079);
and U22427 (N_22427,N_20742,N_20861);
nor U22428 (N_22428,N_20481,N_21112);
nand U22429 (N_22429,N_20540,N_20950);
nor U22430 (N_22430,N_20406,N_21227);
or U22431 (N_22431,N_20420,N_20058);
xor U22432 (N_22432,N_20767,N_20899);
xnor U22433 (N_22433,N_20270,N_21049);
and U22434 (N_22434,N_21178,N_20012);
or U22435 (N_22435,N_21006,N_20587);
nand U22436 (N_22436,N_20076,N_20955);
nor U22437 (N_22437,N_20147,N_20180);
xor U22438 (N_22438,N_20426,N_20345);
and U22439 (N_22439,N_21084,N_20595);
and U22440 (N_22440,N_20799,N_20450);
xnor U22441 (N_22441,N_20453,N_20887);
and U22442 (N_22442,N_20624,N_20447);
and U22443 (N_22443,N_20231,N_20024);
and U22444 (N_22444,N_21064,N_20298);
and U22445 (N_22445,N_20444,N_20653);
or U22446 (N_22446,N_20747,N_20705);
nand U22447 (N_22447,N_20435,N_20717);
xnor U22448 (N_22448,N_21128,N_21146);
and U22449 (N_22449,N_20381,N_21153);
xnor U22450 (N_22450,N_20013,N_20850);
nor U22451 (N_22451,N_21025,N_20396);
nor U22452 (N_22452,N_21202,N_21018);
nor U22453 (N_22453,N_20773,N_20453);
nor U22454 (N_22454,N_20233,N_20879);
xnor U22455 (N_22455,N_20557,N_20324);
or U22456 (N_22456,N_20411,N_20251);
nand U22457 (N_22457,N_20886,N_21102);
xnor U22458 (N_22458,N_20033,N_20531);
nand U22459 (N_22459,N_20706,N_20928);
nor U22460 (N_22460,N_20501,N_21175);
nand U22461 (N_22461,N_20497,N_21219);
or U22462 (N_22462,N_21009,N_20482);
or U22463 (N_22463,N_20548,N_20190);
nand U22464 (N_22464,N_20730,N_21082);
nand U22465 (N_22465,N_20807,N_20161);
or U22466 (N_22466,N_20040,N_20804);
or U22467 (N_22467,N_21134,N_20220);
xnor U22468 (N_22468,N_20466,N_20358);
and U22469 (N_22469,N_21036,N_20831);
or U22470 (N_22470,N_20502,N_20211);
nor U22471 (N_22471,N_21226,N_20235);
and U22472 (N_22472,N_20169,N_21230);
nand U22473 (N_22473,N_20245,N_20241);
and U22474 (N_22474,N_20434,N_21037);
or U22475 (N_22475,N_20949,N_21247);
nor U22476 (N_22476,N_20552,N_20867);
and U22477 (N_22477,N_20655,N_20692);
or U22478 (N_22478,N_20366,N_21109);
nor U22479 (N_22479,N_20109,N_20639);
and U22480 (N_22480,N_20942,N_21021);
and U22481 (N_22481,N_20102,N_20132);
nand U22482 (N_22482,N_20348,N_20339);
nand U22483 (N_22483,N_20334,N_20640);
nor U22484 (N_22484,N_20267,N_20485);
and U22485 (N_22485,N_20087,N_21146);
and U22486 (N_22486,N_20705,N_20288);
nand U22487 (N_22487,N_20976,N_20166);
xor U22488 (N_22488,N_20409,N_20135);
and U22489 (N_22489,N_20805,N_20646);
or U22490 (N_22490,N_20313,N_20789);
nand U22491 (N_22491,N_20251,N_20008);
xor U22492 (N_22492,N_20464,N_20479);
or U22493 (N_22493,N_20039,N_21162);
or U22494 (N_22494,N_20482,N_20464);
nand U22495 (N_22495,N_20226,N_20884);
nor U22496 (N_22496,N_20096,N_21144);
and U22497 (N_22497,N_20705,N_20679);
or U22498 (N_22498,N_20742,N_20065);
xor U22499 (N_22499,N_20113,N_20158);
and U22500 (N_22500,N_22450,N_21719);
nor U22501 (N_22501,N_21460,N_22289);
nor U22502 (N_22502,N_21931,N_21273);
nor U22503 (N_22503,N_21283,N_21937);
nand U22504 (N_22504,N_21718,N_21311);
xnor U22505 (N_22505,N_22108,N_21899);
or U22506 (N_22506,N_22118,N_21877);
or U22507 (N_22507,N_21280,N_21717);
or U22508 (N_22508,N_22447,N_22451);
xor U22509 (N_22509,N_21782,N_22199);
or U22510 (N_22510,N_21855,N_21513);
or U22511 (N_22511,N_21825,N_22381);
and U22512 (N_22512,N_22055,N_22375);
and U22513 (N_22513,N_21888,N_21408);
nor U22514 (N_22514,N_22245,N_21765);
or U22515 (N_22515,N_22133,N_22126);
xnor U22516 (N_22516,N_22013,N_22311);
and U22517 (N_22517,N_22112,N_21594);
and U22518 (N_22518,N_21482,N_21954);
nand U22519 (N_22519,N_21308,N_22073);
nand U22520 (N_22520,N_21788,N_22164);
xnor U22521 (N_22521,N_21777,N_22281);
and U22522 (N_22522,N_21382,N_22001);
or U22523 (N_22523,N_21442,N_21412);
and U22524 (N_22524,N_21720,N_22490);
nor U22525 (N_22525,N_21810,N_21560);
and U22526 (N_22526,N_21912,N_22215);
xnor U22527 (N_22527,N_21252,N_22337);
nand U22528 (N_22528,N_21686,N_22338);
nand U22529 (N_22529,N_22363,N_22256);
xnor U22530 (N_22530,N_22440,N_22237);
nor U22531 (N_22531,N_21292,N_22177);
nor U22532 (N_22532,N_22260,N_21301);
nand U22533 (N_22533,N_21813,N_21354);
nand U22534 (N_22534,N_22343,N_21550);
xnor U22535 (N_22535,N_21724,N_21812);
and U22536 (N_22536,N_22057,N_21380);
xnor U22537 (N_22537,N_22089,N_22261);
nor U22538 (N_22538,N_21994,N_22077);
or U22539 (N_22539,N_22472,N_21956);
or U22540 (N_22540,N_21447,N_21590);
and U22541 (N_22541,N_22029,N_21650);
nor U22542 (N_22542,N_21584,N_22161);
and U22543 (N_22543,N_22146,N_21974);
nand U22544 (N_22544,N_22230,N_22022);
xnor U22545 (N_22545,N_21572,N_21741);
and U22546 (N_22546,N_21330,N_22178);
or U22547 (N_22547,N_21573,N_21869);
and U22548 (N_22548,N_22279,N_21499);
xnor U22549 (N_22549,N_22188,N_22005);
nand U22550 (N_22550,N_21346,N_22492);
and U22551 (N_22551,N_22259,N_22132);
xnor U22552 (N_22552,N_22393,N_22438);
nor U22553 (N_22553,N_22266,N_21522);
or U22554 (N_22554,N_22402,N_21404);
or U22555 (N_22555,N_21933,N_21856);
nand U22556 (N_22556,N_21335,N_21608);
nand U22557 (N_22557,N_22020,N_21520);
xor U22558 (N_22558,N_22332,N_21387);
xor U22559 (N_22559,N_22234,N_21631);
and U22560 (N_22560,N_21474,N_21348);
and U22561 (N_22561,N_21427,N_21998);
or U22562 (N_22562,N_21434,N_21898);
and U22563 (N_22563,N_21776,N_21675);
and U22564 (N_22564,N_21701,N_21975);
xnor U22565 (N_22565,N_22187,N_21599);
and U22566 (N_22566,N_21481,N_21309);
and U22567 (N_22567,N_21723,N_21706);
or U22568 (N_22568,N_22464,N_21725);
or U22569 (N_22569,N_21655,N_21555);
or U22570 (N_22570,N_21430,N_22114);
nor U22571 (N_22571,N_21388,N_21862);
and U22572 (N_22572,N_21909,N_22340);
or U22573 (N_22573,N_21532,N_21523);
or U22574 (N_22574,N_21269,N_22427);
or U22575 (N_22575,N_22488,N_21548);
nor U22576 (N_22576,N_22086,N_22479);
or U22577 (N_22577,N_22449,N_21685);
nand U22578 (N_22578,N_21250,N_21504);
nor U22579 (N_22579,N_21903,N_22244);
xnor U22580 (N_22580,N_22262,N_21907);
nand U22581 (N_22581,N_21964,N_21942);
nor U22582 (N_22582,N_21754,N_22342);
and U22583 (N_22583,N_22064,N_21350);
and U22584 (N_22584,N_21727,N_21651);
or U22585 (N_22585,N_22452,N_22165);
nor U22586 (N_22586,N_21817,N_21772);
nand U22587 (N_22587,N_21323,N_21470);
nor U22588 (N_22588,N_21298,N_21882);
nand U22589 (N_22589,N_21977,N_21875);
and U22590 (N_22590,N_22496,N_21670);
or U22591 (N_22591,N_21566,N_22380);
xor U22592 (N_22592,N_21258,N_21829);
and U22593 (N_22593,N_21413,N_22068);
or U22594 (N_22594,N_21688,N_22305);
and U22595 (N_22595,N_22208,N_22459);
nor U22596 (N_22596,N_22127,N_21652);
and U22597 (N_22597,N_21624,N_22128);
nor U22598 (N_22598,N_21785,N_21851);
and U22599 (N_22599,N_21338,N_22044);
and U22600 (N_22600,N_22238,N_21614);
nand U22601 (N_22601,N_21393,N_22214);
nor U22602 (N_22602,N_21664,N_21733);
nand U22603 (N_22603,N_21973,N_22168);
nor U22604 (N_22604,N_21697,N_21285);
xor U22605 (N_22605,N_22009,N_21756);
xnor U22606 (N_22606,N_21692,N_22019);
and U22607 (N_22607,N_22329,N_22333);
or U22608 (N_22608,N_22475,N_21517);
xor U22609 (N_22609,N_21618,N_21487);
and U22610 (N_22610,N_21431,N_22288);
nand U22611 (N_22611,N_21696,N_21498);
or U22612 (N_22612,N_22360,N_22220);
and U22613 (N_22613,N_21578,N_22499);
nand U22614 (N_22614,N_22071,N_21911);
and U22615 (N_22615,N_21834,N_21366);
nor U22616 (N_22616,N_21627,N_22415);
and U22617 (N_22617,N_22207,N_21360);
and U22618 (N_22618,N_21472,N_21589);
or U22619 (N_22619,N_21748,N_21489);
or U22620 (N_22620,N_21604,N_21377);
xor U22621 (N_22621,N_22198,N_21728);
nand U22622 (N_22622,N_21508,N_21503);
nor U22623 (N_22623,N_22455,N_22115);
xor U22624 (N_22624,N_21780,N_22372);
and U22625 (N_22625,N_21970,N_22028);
or U22626 (N_22626,N_22474,N_21957);
xnor U22627 (N_22627,N_22000,N_21385);
nor U22628 (N_22628,N_21809,N_21617);
nand U22629 (N_22629,N_22058,N_21750);
xor U22630 (N_22630,N_21488,N_21633);
or U22631 (N_22631,N_22246,N_22378);
xor U22632 (N_22632,N_21967,N_21923);
xnor U22633 (N_22633,N_21887,N_21337);
nand U22634 (N_22634,N_22320,N_22181);
and U22635 (N_22635,N_21564,N_21559);
nand U22636 (N_22636,N_21713,N_22122);
and U22637 (N_22637,N_21403,N_21804);
or U22638 (N_22638,N_21781,N_21894);
xor U22639 (N_22639,N_21831,N_21846);
nor U22640 (N_22640,N_21268,N_21893);
and U22641 (N_22641,N_22497,N_22352);
and U22642 (N_22642,N_21310,N_22139);
nand U22643 (N_22643,N_22038,N_21859);
or U22644 (N_22644,N_21658,N_22142);
and U22645 (N_22645,N_22345,N_21251);
nor U22646 (N_22646,N_22152,N_21902);
nand U22647 (N_22647,N_22042,N_21542);
and U22648 (N_22648,N_22463,N_21928);
nand U22649 (N_22649,N_22151,N_21419);
or U22650 (N_22650,N_22141,N_22160);
xnor U22651 (N_22651,N_22027,N_21418);
nor U22652 (N_22652,N_21300,N_21867);
or U22653 (N_22653,N_22222,N_21468);
nand U22654 (N_22654,N_21556,N_21635);
and U22655 (N_22655,N_22493,N_21277);
xnor U22656 (N_22656,N_21653,N_21314);
or U22657 (N_22657,N_21986,N_22206);
nand U22658 (N_22658,N_21381,N_21730);
or U22659 (N_22659,N_21798,N_21569);
and U22660 (N_22660,N_22482,N_21477);
nand U22661 (N_22661,N_22078,N_22460);
and U22662 (N_22662,N_21553,N_21575);
nor U22663 (N_22663,N_21443,N_21265);
or U22664 (N_22664,N_22148,N_21913);
nand U22665 (N_22665,N_21509,N_21270);
xnor U22666 (N_22666,N_21819,N_22006);
and U22667 (N_22667,N_22418,N_21878);
xnor U22668 (N_22668,N_21726,N_21996);
nor U22669 (N_22669,N_21676,N_22030);
xor U22670 (N_22670,N_22051,N_21304);
nand U22671 (N_22671,N_22173,N_22365);
or U22672 (N_22672,N_21552,N_21716);
xnor U22673 (N_22673,N_22185,N_22346);
and U22674 (N_22674,N_22322,N_22087);
nor U22675 (N_22675,N_22095,N_21699);
or U22676 (N_22676,N_21574,N_22016);
or U22677 (N_22677,N_21332,N_21511);
and U22678 (N_22678,N_21557,N_21389);
nand U22679 (N_22679,N_22473,N_21497);
nand U22680 (N_22680,N_21592,N_22159);
nor U22681 (N_22681,N_21839,N_22062);
and U22682 (N_22682,N_21405,N_22075);
nand U22683 (N_22683,N_22248,N_21462);
nand U22684 (N_22684,N_21806,N_21944);
or U22685 (N_22685,N_21990,N_21634);
xnor U22686 (N_22686,N_22403,N_21612);
xor U22687 (N_22687,N_21355,N_21491);
nand U22688 (N_22688,N_21565,N_21929);
nor U22689 (N_22689,N_21345,N_22123);
xnor U22690 (N_22690,N_21734,N_22102);
or U22691 (N_22691,N_21274,N_21784);
and U22692 (N_22692,N_21885,N_22325);
nor U22693 (N_22693,N_21968,N_22134);
and U22694 (N_22694,N_22221,N_21392);
nor U22695 (N_22695,N_21845,N_21663);
nor U22696 (N_22696,N_21526,N_21591);
nand U22697 (N_22697,N_21561,N_21527);
xnor U22698 (N_22698,N_21879,N_22462);
xnor U22699 (N_22699,N_21950,N_21953);
xor U22700 (N_22700,N_22357,N_22179);
nand U22701 (N_22701,N_22034,N_21373);
nor U22702 (N_22702,N_21638,N_21399);
nand U22703 (N_22703,N_22258,N_21991);
nor U22704 (N_22704,N_21985,N_21883);
xor U22705 (N_22705,N_21786,N_21948);
nand U22706 (N_22706,N_21336,N_21865);
nor U22707 (N_22707,N_21828,N_21826);
nor U22708 (N_22708,N_21476,N_22251);
or U22709 (N_22709,N_21352,N_21537);
or U22710 (N_22710,N_21600,N_21854);
xnor U22711 (N_22711,N_21293,N_21266);
nand U22712 (N_22712,N_22196,N_22439);
xor U22713 (N_22713,N_21965,N_22436);
nor U22714 (N_22714,N_21630,N_22094);
nand U22715 (N_22715,N_22454,N_21836);
nor U22716 (N_22716,N_22053,N_22025);
xnor U22717 (N_22717,N_22153,N_21708);
nor U22718 (N_22718,N_21414,N_21820);
or U22719 (N_22719,N_21762,N_21299);
nand U22720 (N_22720,N_22136,N_22303);
nand U22721 (N_22721,N_21282,N_21496);
or U22722 (N_22722,N_22377,N_22280);
nand U22723 (N_22723,N_21347,N_21473);
and U22724 (N_22724,N_21945,N_21666);
xor U22725 (N_22725,N_21607,N_21936);
nor U22726 (N_22726,N_21409,N_22236);
nand U22727 (N_22727,N_22219,N_22318);
xnor U22728 (N_22728,N_22400,N_21778);
xor U22729 (N_22729,N_22107,N_22045);
nor U22730 (N_22730,N_21823,N_22444);
and U22731 (N_22731,N_22176,N_22110);
xor U22732 (N_22732,N_22106,N_22171);
or U22733 (N_22733,N_21534,N_21976);
nand U22734 (N_22734,N_21621,N_21326);
or U22735 (N_22735,N_22056,N_21712);
xor U22736 (N_22736,N_22366,N_21689);
and U22737 (N_22737,N_21832,N_22186);
or U22738 (N_22738,N_22046,N_22384);
or U22739 (N_22739,N_22412,N_22494);
nor U22740 (N_22740,N_21288,N_21458);
nor U22741 (N_22741,N_22465,N_22074);
or U22742 (N_22742,N_21475,N_22469);
nor U22743 (N_22743,N_21735,N_22278);
nor U22744 (N_22744,N_22461,N_21359);
nand U22745 (N_22745,N_21428,N_21917);
nand U22746 (N_22746,N_22167,N_22379);
nand U22747 (N_22747,N_21463,N_21294);
and U22748 (N_22748,N_21276,N_21671);
and U22749 (N_22749,N_21992,N_22374);
or U22750 (N_22750,N_22401,N_21597);
nor U22751 (N_22751,N_21822,N_21924);
nand U22752 (N_22752,N_21988,N_22286);
and U22753 (N_22753,N_21915,N_22209);
or U22754 (N_22754,N_22104,N_21512);
and U22755 (N_22755,N_21690,N_21400);
xnor U22756 (N_22756,N_22388,N_22033);
nand U22757 (N_22757,N_21921,N_22390);
or U22758 (N_22758,N_21800,N_21925);
nand U22759 (N_22759,N_22323,N_22267);
nand U22760 (N_22760,N_22232,N_21943);
nand U22761 (N_22761,N_21629,N_22295);
nand U22762 (N_22762,N_21455,N_21637);
and U22763 (N_22763,N_22495,N_21922);
or U22764 (N_22764,N_22011,N_21383);
nor U22765 (N_22765,N_21742,N_21320);
or U22766 (N_22766,N_22275,N_21640);
nand U22767 (N_22767,N_21585,N_21744);
nand U22768 (N_22768,N_21279,N_22297);
nand U22769 (N_22769,N_21371,N_21540);
and U22770 (N_22770,N_21372,N_21884);
and U22771 (N_22771,N_22096,N_22347);
nand U22772 (N_22772,N_22334,N_22240);
or U22773 (N_22773,N_22026,N_21480);
or U22774 (N_22774,N_21551,N_22098);
nand U22775 (N_22775,N_21702,N_21278);
or U22776 (N_22776,N_22483,N_21598);
nor U22777 (N_22777,N_21313,N_22394);
nand U22778 (N_22778,N_22399,N_22067);
nor U22779 (N_22779,N_21467,N_22478);
nand U22780 (N_22780,N_21426,N_21287);
nand U22781 (N_22781,N_21451,N_21626);
or U22782 (N_22782,N_21303,N_22480);
nor U22783 (N_22783,N_21502,N_21824);
nor U22784 (N_22784,N_21642,N_21681);
or U22785 (N_22785,N_21615,N_21619);
or U22786 (N_22786,N_21456,N_21721);
xor U22787 (N_22787,N_22210,N_21500);
or U22788 (N_22788,N_22428,N_21581);
nand U22789 (N_22789,N_22316,N_22012);
nor U22790 (N_22790,N_22231,N_21580);
and U22791 (N_22791,N_22306,N_21745);
xnor U22792 (N_22792,N_22111,N_21789);
or U22793 (N_22793,N_22154,N_21654);
nor U22794 (N_22794,N_21763,N_21448);
xnor U22795 (N_22795,N_21764,N_21889);
nor U22796 (N_22796,N_21466,N_21835);
nor U22797 (N_22797,N_22109,N_22117);
or U22798 (N_22798,N_21325,N_22298);
nor U22799 (N_22799,N_21940,N_21356);
xor U22800 (N_22800,N_21732,N_21683);
nand U22801 (N_22801,N_22330,N_22191);
and U22802 (N_22802,N_22489,N_21432);
and U22803 (N_22803,N_22430,N_22113);
xnor U22804 (N_22804,N_21868,N_22140);
or U22805 (N_22805,N_22359,N_22476);
nand U22806 (N_22806,N_21286,N_21871);
nor U22807 (N_22807,N_21770,N_21562);
xnor U22808 (N_22808,N_21773,N_21648);
or U22809 (N_22809,N_21257,N_21679);
or U22810 (N_22810,N_22253,N_22395);
xor U22811 (N_22811,N_21863,N_21351);
nor U22812 (N_22812,N_21886,N_21441);
and U22813 (N_22813,N_21736,N_21814);
nor U22814 (N_22814,N_22069,N_22131);
xor U22815 (N_22815,N_21622,N_21774);
nor U22816 (N_22816,N_22304,N_21691);
or U22817 (N_22817,N_21368,N_22054);
or U22818 (N_22818,N_21394,N_21340);
xor U22819 (N_22819,N_22409,N_22484);
and U22820 (N_22820,N_21905,N_22018);
nor U22821 (N_22821,N_21980,N_22119);
or U22822 (N_22822,N_21792,N_22211);
and U22823 (N_22823,N_22383,N_22202);
xor U22824 (N_22824,N_21535,N_21844);
nor U22825 (N_22825,N_21367,N_22097);
or U22826 (N_22826,N_21757,N_22195);
and U22827 (N_22827,N_21486,N_22060);
nand U22828 (N_22828,N_21932,N_22021);
xnor U22829 (N_22829,N_22170,N_21541);
or U22830 (N_22830,N_21495,N_21677);
nand U22831 (N_22831,N_21331,N_21737);
and U22832 (N_22832,N_21319,N_21505);
and U22833 (N_22833,N_21935,N_22437);
xor U22834 (N_22834,N_21661,N_21904);
and U22835 (N_22835,N_22453,N_21853);
and U22836 (N_22836,N_21946,N_21445);
and U22837 (N_22837,N_21563,N_21843);
nand U22838 (N_22838,N_22043,N_21914);
nand U22839 (N_22839,N_21593,N_21892);
nand U22840 (N_22840,N_21860,N_22326);
xnor U22841 (N_22841,N_22156,N_22235);
and U22842 (N_22842,N_21729,N_21465);
nand U22843 (N_22843,N_21791,N_21861);
nor U22844 (N_22844,N_22413,N_22270);
xor U22845 (N_22845,N_21739,N_21398);
and U22846 (N_22846,N_21391,N_21628);
xnor U22847 (N_22847,N_21406,N_22143);
nor U22848 (N_22848,N_21411,N_22242);
nand U22849 (N_22849,N_21874,N_22189);
nand U22850 (N_22850,N_22371,N_22446);
and U22851 (N_22851,N_22432,N_21515);
nand U22852 (N_22852,N_22405,N_21710);
and U22853 (N_22853,N_21849,N_22082);
xnor U22854 (N_22854,N_21769,N_21571);
or U22855 (N_22855,N_22424,N_22302);
nand U22856 (N_22856,N_21587,N_21672);
xor U22857 (N_22857,N_21811,N_22217);
xor U22858 (N_22858,N_21687,N_21866);
nor U22859 (N_22859,N_21848,N_21751);
nand U22860 (N_22860,N_21646,N_22024);
or U22861 (N_22861,N_21343,N_21521);
nor U22862 (N_22862,N_21318,N_22085);
nand U22863 (N_22863,N_22312,N_22150);
or U22864 (N_22864,N_22169,N_22088);
or U22865 (N_22865,N_22174,N_21795);
and U22866 (N_22866,N_21362,N_21760);
or U22867 (N_22867,N_22397,N_22081);
xnor U22868 (N_22868,N_22285,N_22434);
and U22869 (N_22869,N_22335,N_21524);
xor U22870 (N_22870,N_22373,N_21281);
nor U22871 (N_22871,N_22435,N_21349);
nand U22872 (N_22872,N_21386,N_21966);
nor U22873 (N_22873,N_21963,N_21930);
and U22874 (N_22874,N_22367,N_21514);
nand U22875 (N_22875,N_21852,N_21987);
and U22876 (N_22876,N_21410,N_21955);
xor U22877 (N_22877,N_21595,N_21494);
nor U22878 (N_22878,N_21972,N_21461);
nor U22879 (N_22879,N_22105,N_22162);
or U22880 (N_22880,N_22369,N_21397);
and U22881 (N_22881,N_22282,N_22183);
nand U22882 (N_22882,N_21596,N_21457);
or U22883 (N_22883,N_22124,N_22315);
nand U22884 (N_22884,N_21433,N_21890);
and U22885 (N_22885,N_21401,N_22052);
nor U22886 (N_22886,N_22203,N_21827);
xnor U22887 (N_22887,N_22300,N_21421);
or U22888 (N_22888,N_22149,N_22442);
nor U22889 (N_22889,N_22125,N_22041);
and U22890 (N_22890,N_21850,N_22339);
or U22891 (N_22891,N_21339,N_21983);
nor U22892 (N_22892,N_22036,N_21808);
xnor U22893 (N_22893,N_21993,N_22184);
and U22894 (N_22894,N_21544,N_21938);
xnor U22895 (N_22895,N_22299,N_22370);
nand U22896 (N_22896,N_21284,N_21793);
nor U22897 (N_22897,N_21695,N_21324);
and U22898 (N_22898,N_22396,N_22080);
and U22899 (N_22899,N_22091,N_22227);
or U22900 (N_22900,N_22129,N_22048);
or U22901 (N_22901,N_22182,N_22003);
xnor U22902 (N_22902,N_21603,N_22099);
nand U22903 (N_22903,N_21342,N_21538);
nand U22904 (N_22904,N_21816,N_21478);
nor U22905 (N_22905,N_21361,N_21771);
xnor U22906 (N_22906,N_21830,N_22361);
nand U22907 (N_22907,N_22145,N_22100);
or U22908 (N_22908,N_21821,N_22348);
or U22909 (N_22909,N_21805,N_22355);
and U22910 (N_22910,N_22175,N_21753);
or U22911 (N_22911,N_22284,N_22336);
nand U22912 (N_22912,N_21799,N_21295);
xnor U22913 (N_22913,N_21801,N_21643);
and U22914 (N_22914,N_21424,N_21711);
and U22915 (N_22915,N_22172,N_21605);
xnor U22916 (N_22916,N_21506,N_22283);
and U22917 (N_22917,N_21897,N_22121);
nand U22918 (N_22918,N_22101,N_21507);
xnor U22919 (N_22919,N_21369,N_21297);
and U22920 (N_22920,N_21900,N_21315);
and U22921 (N_22921,N_22408,N_21375);
xnor U22922 (N_22922,N_21864,N_21895);
nor U22923 (N_22923,N_21947,N_22276);
nand U22924 (N_22924,N_22090,N_22201);
nor U22925 (N_22925,N_21978,N_22471);
and U22926 (N_22926,N_22116,N_22155);
nand U22927 (N_22927,N_21305,N_22213);
nand U22928 (N_22928,N_21841,N_21317);
or U22929 (N_22929,N_22414,N_21379);
nor U22930 (N_22930,N_21546,N_21700);
nor U22931 (N_22931,N_22243,N_21962);
and U22932 (N_22932,N_21601,N_22263);
and U22933 (N_22933,N_22007,N_22002);
nand U22934 (N_22934,N_22228,N_21370);
xor U22935 (N_22935,N_21531,N_21396);
nor U22936 (N_22936,N_21668,N_21636);
and U22937 (N_22937,N_21549,N_22406);
and U22938 (N_22938,N_21847,N_21838);
and U22939 (N_22939,N_21632,N_21260);
xnor U22940 (N_22940,N_22037,N_22032);
nand U22941 (N_22941,N_21684,N_22274);
and U22942 (N_22942,N_21464,N_21759);
or U22943 (N_22943,N_22010,N_22314);
nor U22944 (N_22944,N_22239,N_21704);
xor U22945 (N_22945,N_21602,N_22225);
nor U22946 (N_22946,N_21390,N_22130);
nand U22947 (N_22947,N_21450,N_22456);
nand U22948 (N_22948,N_21678,N_22192);
and U22949 (N_22949,N_21960,N_21749);
xnor U22950 (N_22950,N_21334,N_22392);
nand U22951 (N_22951,N_21952,N_22387);
xnor U22952 (N_22952,N_22040,N_21436);
or U22953 (N_22953,N_22050,N_21459);
and U22954 (N_22954,N_22420,N_22218);
nand U22955 (N_22955,N_22470,N_21896);
and U22956 (N_22956,N_21981,N_21610);
xnor U22957 (N_22957,N_21576,N_21698);
and U22958 (N_22958,N_22180,N_21919);
and U22959 (N_22959,N_22431,N_21803);
nand U22960 (N_22960,N_21918,N_21645);
nor U22961 (N_22961,N_22204,N_21705);
nand U22962 (N_22962,N_22331,N_22223);
xnor U22963 (N_22963,N_21870,N_21586);
or U22964 (N_22964,N_22233,N_21920);
and U22965 (N_22965,N_22035,N_21767);
or U22966 (N_22966,N_22294,N_22458);
and U22967 (N_22967,N_21583,N_21490);
nor U22968 (N_22968,N_22349,N_22076);
nor U22969 (N_22969,N_21395,N_21543);
nor U22970 (N_22970,N_22317,N_22324);
xor U22971 (N_22971,N_22354,N_21858);
or U22972 (N_22972,N_21766,N_22350);
nor U22973 (N_22973,N_21402,N_21358);
and U22974 (N_22974,N_21302,N_21989);
nor U22975 (N_22975,N_21471,N_21949);
nor U22976 (N_22976,N_21255,N_21329);
and U22977 (N_22977,N_22356,N_22015);
or U22978 (N_22978,N_21483,N_21916);
and U22979 (N_22979,N_22072,N_21876);
xor U22980 (N_22980,N_21623,N_21840);
nand U22981 (N_22981,N_22481,N_22092);
xor U22982 (N_22982,N_22008,N_21364);
nor U22983 (N_22983,N_22419,N_21709);
or U22984 (N_22984,N_21694,N_22407);
or U22985 (N_22985,N_21665,N_21452);
and U22986 (N_22986,N_22065,N_22466);
and U22987 (N_22987,N_21908,N_22120);
and U22988 (N_22988,N_21272,N_22047);
and U22989 (N_22989,N_21797,N_22252);
nor U22990 (N_22990,N_21755,N_21941);
and U22991 (N_22991,N_21253,N_21647);
and U22992 (N_22992,N_21363,N_22190);
or U22993 (N_22993,N_22287,N_22158);
nor U22994 (N_22994,N_22014,N_22426);
nand U22995 (N_22995,N_21365,N_22327);
nor U22996 (N_22996,N_21384,N_21926);
or U22997 (N_22997,N_21656,N_21775);
or U22998 (N_22998,N_22273,N_22468);
nand U22999 (N_22999,N_22376,N_22429);
xor U23000 (N_23000,N_21423,N_22486);
xnor U23001 (N_23001,N_21558,N_21842);
and U23002 (N_23002,N_21446,N_21620);
xnor U23003 (N_23003,N_21625,N_21525);
xnor U23004 (N_23004,N_21256,N_21995);
nand U23005 (N_23005,N_21644,N_21416);
xnor U23006 (N_23006,N_22059,N_21485);
nor U23007 (N_23007,N_22061,N_21740);
nor U23008 (N_23008,N_21554,N_21743);
nor U23009 (N_23009,N_21731,N_21417);
nand U23010 (N_23010,N_22353,N_22467);
and U23011 (N_23011,N_21790,N_22385);
or U23012 (N_23012,N_22250,N_22039);
nand U23013 (N_23013,N_21873,N_22157);
nor U23014 (N_23014,N_21703,N_21818);
nand U23015 (N_23015,N_22457,N_21881);
nor U23016 (N_23016,N_22448,N_22255);
nor U23017 (N_23017,N_21880,N_21588);
or U23018 (N_23018,N_22103,N_21307);
nor U23019 (N_23019,N_21752,N_22277);
xnor U23020 (N_23020,N_21693,N_21682);
or U23021 (N_23021,N_21312,N_21783);
xnor U23022 (N_23022,N_22200,N_22272);
nor U23023 (N_23023,N_22066,N_22309);
and U23024 (N_23024,N_21261,N_22249);
xor U23025 (N_23025,N_22487,N_21439);
or U23026 (N_23026,N_22194,N_22477);
nor U23027 (N_23027,N_22310,N_21707);
and U23028 (N_23028,N_22368,N_22319);
and U23029 (N_23029,N_22386,N_21997);
and U23030 (N_23030,N_22358,N_22328);
nand U23031 (N_23031,N_21833,N_21415);
nand U23032 (N_23032,N_21961,N_22254);
and U23033 (N_23033,N_22389,N_22084);
and U23034 (N_23034,N_21420,N_21802);
and U23035 (N_23035,N_22144,N_22093);
nor U23036 (N_23036,N_21906,N_21747);
or U23037 (N_23037,N_22307,N_21714);
and U23038 (N_23038,N_22441,N_21259);
and U23039 (N_23039,N_22265,N_22163);
xnor U23040 (N_23040,N_21639,N_21971);
or U23041 (N_23041,N_21984,N_22166);
xnor U23042 (N_23042,N_21289,N_21577);
xor U23043 (N_23043,N_22296,N_21582);
or U23044 (N_23044,N_21758,N_22229);
nor U23045 (N_23045,N_21999,N_21533);
and U23046 (N_23046,N_21787,N_21738);
and U23047 (N_23047,N_21568,N_21939);
nor U23048 (N_23048,N_21761,N_21910);
and U23049 (N_23049,N_21982,N_21667);
and U23050 (N_23050,N_21437,N_22351);
and U23051 (N_23051,N_21901,N_22017);
nor U23052 (N_23052,N_22137,N_22301);
or U23053 (N_23053,N_21969,N_21492);
and U23054 (N_23054,N_21341,N_22498);
and U23055 (N_23055,N_21254,N_22321);
nand U23056 (N_23056,N_22308,N_21449);
or U23057 (N_23057,N_21479,N_21794);
and U23058 (N_23058,N_21609,N_22147);
and U23059 (N_23059,N_22226,N_21951);
nor U23060 (N_23060,N_21570,N_22290);
and U23061 (N_23061,N_22364,N_21333);
nor U23062 (N_23062,N_21606,N_22271);
xor U23063 (N_23063,N_21353,N_22070);
and U23064 (N_23064,N_21616,N_22031);
and U23065 (N_23065,N_22391,N_22224);
or U23066 (N_23066,N_22443,N_21267);
or U23067 (N_23067,N_21807,N_21872);
or U23068 (N_23068,N_21611,N_22247);
nor U23069 (N_23069,N_21407,N_22291);
and U23070 (N_23070,N_21530,N_22264);
xor U23071 (N_23071,N_22293,N_21641);
nand U23072 (N_23072,N_21680,N_21528);
or U23073 (N_23073,N_21715,N_22425);
nor U23074 (N_23074,N_21422,N_21429);
nand U23075 (N_23075,N_22138,N_21263);
or U23076 (N_23076,N_21673,N_22341);
nor U23077 (N_23077,N_21453,N_22216);
and U23078 (N_23078,N_21516,N_21316);
and U23079 (N_23079,N_22205,N_21321);
and U23080 (N_23080,N_21438,N_21322);
and U23081 (N_23081,N_22417,N_21484);
or U23082 (N_23082,N_22193,N_22362);
xor U23083 (N_23083,N_21501,N_21435);
or U23084 (N_23084,N_21440,N_21979);
and U23085 (N_23085,N_22433,N_21327);
or U23086 (N_23086,N_21469,N_21746);
nand U23087 (N_23087,N_21328,N_21796);
or U23088 (N_23088,N_21374,N_21547);
xnor U23089 (N_23089,N_21425,N_21657);
nand U23090 (N_23090,N_21271,N_21510);
xor U23091 (N_23091,N_21649,N_21545);
nand U23092 (N_23092,N_21722,N_21376);
and U23093 (N_23093,N_21857,N_22049);
nand U23094 (N_23094,N_22423,N_22212);
nand U23095 (N_23095,N_21296,N_22257);
or U23096 (N_23096,N_21306,N_22410);
and U23097 (N_23097,N_22404,N_22135);
and U23098 (N_23098,N_22023,N_22269);
and U23099 (N_23099,N_21378,N_21669);
or U23100 (N_23100,N_22268,N_21674);
and U23101 (N_23101,N_22411,N_22313);
or U23102 (N_23102,N_22445,N_22004);
xor U23103 (N_23103,N_21934,N_21567);
and U23104 (N_23104,N_21659,N_22241);
xor U23105 (N_23105,N_21579,N_22292);
nand U23106 (N_23106,N_21444,N_21959);
xnor U23107 (N_23107,N_21662,N_21275);
xnor U23108 (N_23108,N_22083,N_21927);
or U23109 (N_23109,N_22422,N_22491);
nand U23110 (N_23110,N_21815,N_22344);
and U23111 (N_23111,N_22063,N_21518);
or U23112 (N_23112,N_21837,N_21613);
xor U23113 (N_23113,N_21344,N_21779);
nor U23114 (N_23114,N_22079,N_22421);
nor U23115 (N_23115,N_21529,N_22398);
xor U23116 (N_23116,N_21262,N_22197);
nand U23117 (N_23117,N_21539,N_21768);
xnor U23118 (N_23118,N_21357,N_21264);
xnor U23119 (N_23119,N_21290,N_21660);
and U23120 (N_23120,N_22382,N_21891);
nand U23121 (N_23121,N_21519,N_21493);
xor U23122 (N_23122,N_22416,N_21536);
or U23123 (N_23123,N_22485,N_21291);
nor U23124 (N_23124,N_21958,N_21454);
or U23125 (N_23125,N_21468,N_22234);
nor U23126 (N_23126,N_21606,N_22467);
xor U23127 (N_23127,N_21368,N_21717);
xnor U23128 (N_23128,N_21606,N_21867);
or U23129 (N_23129,N_21999,N_22420);
xor U23130 (N_23130,N_21702,N_21369);
xnor U23131 (N_23131,N_21684,N_21809);
or U23132 (N_23132,N_21530,N_22466);
nor U23133 (N_23133,N_21568,N_22231);
or U23134 (N_23134,N_21386,N_21368);
xor U23135 (N_23135,N_22387,N_22381);
nor U23136 (N_23136,N_21701,N_21973);
nor U23137 (N_23137,N_22498,N_21686);
xor U23138 (N_23138,N_22435,N_22051);
and U23139 (N_23139,N_22056,N_21403);
nor U23140 (N_23140,N_21600,N_22219);
and U23141 (N_23141,N_21655,N_21757);
nor U23142 (N_23142,N_22216,N_21903);
or U23143 (N_23143,N_21617,N_21535);
nand U23144 (N_23144,N_21576,N_22261);
nand U23145 (N_23145,N_21904,N_22476);
and U23146 (N_23146,N_21363,N_21366);
xor U23147 (N_23147,N_21427,N_21721);
and U23148 (N_23148,N_22457,N_21406);
xor U23149 (N_23149,N_21890,N_21642);
nand U23150 (N_23150,N_22489,N_21433);
nand U23151 (N_23151,N_21966,N_21611);
and U23152 (N_23152,N_21878,N_21406);
or U23153 (N_23153,N_21302,N_21741);
and U23154 (N_23154,N_22024,N_22328);
xnor U23155 (N_23155,N_21339,N_22246);
nor U23156 (N_23156,N_22077,N_21871);
nand U23157 (N_23157,N_22297,N_22124);
nand U23158 (N_23158,N_21538,N_21609);
or U23159 (N_23159,N_21847,N_22383);
xnor U23160 (N_23160,N_22319,N_21962);
xor U23161 (N_23161,N_22445,N_21391);
xnor U23162 (N_23162,N_22089,N_22181);
xnor U23163 (N_23163,N_21946,N_22243);
nor U23164 (N_23164,N_21900,N_21814);
nor U23165 (N_23165,N_21484,N_22250);
xor U23166 (N_23166,N_21540,N_22171);
and U23167 (N_23167,N_21509,N_21857);
nand U23168 (N_23168,N_21385,N_22314);
or U23169 (N_23169,N_22009,N_21412);
nand U23170 (N_23170,N_21993,N_21540);
nand U23171 (N_23171,N_22385,N_21630);
nand U23172 (N_23172,N_21686,N_22263);
or U23173 (N_23173,N_21482,N_21789);
or U23174 (N_23174,N_21540,N_21729);
xor U23175 (N_23175,N_21995,N_22080);
nand U23176 (N_23176,N_21877,N_22149);
xnor U23177 (N_23177,N_21519,N_22351);
nor U23178 (N_23178,N_22098,N_22378);
and U23179 (N_23179,N_21861,N_22043);
nand U23180 (N_23180,N_21955,N_22483);
nor U23181 (N_23181,N_22440,N_21540);
or U23182 (N_23182,N_21806,N_22093);
or U23183 (N_23183,N_21942,N_21532);
or U23184 (N_23184,N_22054,N_22349);
nand U23185 (N_23185,N_21855,N_22169);
xnor U23186 (N_23186,N_21884,N_21476);
or U23187 (N_23187,N_21912,N_21417);
or U23188 (N_23188,N_21624,N_21993);
nand U23189 (N_23189,N_22298,N_21281);
or U23190 (N_23190,N_22180,N_21588);
xnor U23191 (N_23191,N_22411,N_22176);
and U23192 (N_23192,N_21888,N_22429);
nor U23193 (N_23193,N_22042,N_21707);
or U23194 (N_23194,N_22460,N_22330);
xor U23195 (N_23195,N_21863,N_21297);
xnor U23196 (N_23196,N_21341,N_22244);
and U23197 (N_23197,N_21810,N_21791);
or U23198 (N_23198,N_22080,N_21448);
nand U23199 (N_23199,N_21383,N_21979);
or U23200 (N_23200,N_21888,N_22340);
xor U23201 (N_23201,N_21627,N_22285);
and U23202 (N_23202,N_21487,N_22010);
nor U23203 (N_23203,N_22491,N_21385);
nor U23204 (N_23204,N_22027,N_22494);
nand U23205 (N_23205,N_21438,N_21768);
nor U23206 (N_23206,N_21697,N_21857);
nor U23207 (N_23207,N_22392,N_22029);
nand U23208 (N_23208,N_21692,N_21586);
and U23209 (N_23209,N_21252,N_21478);
or U23210 (N_23210,N_22338,N_21549);
or U23211 (N_23211,N_22176,N_21464);
nand U23212 (N_23212,N_22412,N_22489);
nor U23213 (N_23213,N_21737,N_21299);
nand U23214 (N_23214,N_21266,N_22289);
nand U23215 (N_23215,N_22307,N_22051);
or U23216 (N_23216,N_21727,N_21646);
nor U23217 (N_23217,N_21347,N_21507);
and U23218 (N_23218,N_21398,N_22150);
nor U23219 (N_23219,N_21862,N_21356);
or U23220 (N_23220,N_22263,N_21279);
xor U23221 (N_23221,N_22249,N_22385);
and U23222 (N_23222,N_21511,N_21390);
or U23223 (N_23223,N_21774,N_22246);
nand U23224 (N_23224,N_21545,N_22123);
nand U23225 (N_23225,N_21494,N_22378);
or U23226 (N_23226,N_21637,N_21953);
xnor U23227 (N_23227,N_22256,N_22188);
nor U23228 (N_23228,N_21953,N_21721);
or U23229 (N_23229,N_21462,N_21483);
nor U23230 (N_23230,N_21289,N_21462);
xnor U23231 (N_23231,N_21637,N_21464);
or U23232 (N_23232,N_21649,N_21739);
and U23233 (N_23233,N_22497,N_21332);
and U23234 (N_23234,N_21932,N_21613);
and U23235 (N_23235,N_21869,N_22029);
or U23236 (N_23236,N_21718,N_21669);
nor U23237 (N_23237,N_21341,N_21580);
xor U23238 (N_23238,N_21938,N_21716);
xnor U23239 (N_23239,N_22000,N_22379);
and U23240 (N_23240,N_22112,N_21402);
and U23241 (N_23241,N_21261,N_21820);
nor U23242 (N_23242,N_21597,N_21471);
nor U23243 (N_23243,N_22055,N_22393);
nand U23244 (N_23244,N_22228,N_21997);
nor U23245 (N_23245,N_21792,N_21808);
or U23246 (N_23246,N_22069,N_21924);
nand U23247 (N_23247,N_21451,N_21996);
nor U23248 (N_23248,N_21630,N_22359);
nor U23249 (N_23249,N_21880,N_22072);
nor U23250 (N_23250,N_21288,N_22309);
nand U23251 (N_23251,N_21884,N_21913);
xor U23252 (N_23252,N_21825,N_21363);
nor U23253 (N_23253,N_22173,N_22487);
nand U23254 (N_23254,N_22241,N_21725);
xnor U23255 (N_23255,N_22032,N_22169);
nand U23256 (N_23256,N_21641,N_21541);
nand U23257 (N_23257,N_22001,N_22433);
xnor U23258 (N_23258,N_21780,N_21794);
xor U23259 (N_23259,N_22209,N_21464);
nand U23260 (N_23260,N_21552,N_21687);
xnor U23261 (N_23261,N_21365,N_22283);
nor U23262 (N_23262,N_21351,N_21430);
xor U23263 (N_23263,N_22076,N_21843);
or U23264 (N_23264,N_21662,N_22450);
or U23265 (N_23265,N_21643,N_21945);
nor U23266 (N_23266,N_22496,N_21666);
and U23267 (N_23267,N_22273,N_21913);
and U23268 (N_23268,N_21822,N_22292);
and U23269 (N_23269,N_21863,N_21584);
or U23270 (N_23270,N_22351,N_21425);
and U23271 (N_23271,N_21541,N_21624);
nand U23272 (N_23272,N_21632,N_22244);
or U23273 (N_23273,N_21779,N_21595);
nor U23274 (N_23274,N_21522,N_22189);
and U23275 (N_23275,N_22264,N_22340);
or U23276 (N_23276,N_21954,N_21933);
xnor U23277 (N_23277,N_21402,N_21348);
or U23278 (N_23278,N_21800,N_21707);
or U23279 (N_23279,N_22450,N_22131);
nor U23280 (N_23280,N_21947,N_21630);
and U23281 (N_23281,N_22335,N_22310);
nor U23282 (N_23282,N_22251,N_21724);
and U23283 (N_23283,N_21381,N_21452);
nand U23284 (N_23284,N_21705,N_21793);
nand U23285 (N_23285,N_22025,N_21508);
xor U23286 (N_23286,N_22427,N_21886);
nand U23287 (N_23287,N_21281,N_22142);
nand U23288 (N_23288,N_22135,N_21469);
or U23289 (N_23289,N_21806,N_22047);
or U23290 (N_23290,N_21933,N_21992);
xor U23291 (N_23291,N_21896,N_21936);
or U23292 (N_23292,N_21539,N_21945);
nand U23293 (N_23293,N_21548,N_21709);
nand U23294 (N_23294,N_21682,N_22098);
nor U23295 (N_23295,N_21312,N_21271);
or U23296 (N_23296,N_22374,N_22386);
or U23297 (N_23297,N_22450,N_21511);
and U23298 (N_23298,N_21634,N_22246);
and U23299 (N_23299,N_21288,N_21918);
and U23300 (N_23300,N_21460,N_22316);
or U23301 (N_23301,N_21558,N_21942);
or U23302 (N_23302,N_22262,N_21978);
and U23303 (N_23303,N_22412,N_21621);
and U23304 (N_23304,N_21917,N_21548);
or U23305 (N_23305,N_22414,N_21755);
nor U23306 (N_23306,N_21933,N_21447);
xor U23307 (N_23307,N_21290,N_21339);
nand U23308 (N_23308,N_21940,N_21474);
or U23309 (N_23309,N_22249,N_21727);
xnor U23310 (N_23310,N_21791,N_21813);
nand U23311 (N_23311,N_21534,N_21889);
nand U23312 (N_23312,N_22008,N_21923);
nand U23313 (N_23313,N_21270,N_21295);
xor U23314 (N_23314,N_21945,N_21490);
xnor U23315 (N_23315,N_22049,N_21647);
or U23316 (N_23316,N_21777,N_21707);
nor U23317 (N_23317,N_21519,N_21618);
nor U23318 (N_23318,N_21555,N_21552);
and U23319 (N_23319,N_22262,N_21601);
and U23320 (N_23320,N_21963,N_22057);
and U23321 (N_23321,N_21333,N_22040);
xor U23322 (N_23322,N_21939,N_21702);
and U23323 (N_23323,N_21457,N_21310);
xnor U23324 (N_23324,N_21350,N_22405);
xor U23325 (N_23325,N_22020,N_22445);
xor U23326 (N_23326,N_22090,N_21846);
and U23327 (N_23327,N_22006,N_21749);
and U23328 (N_23328,N_21421,N_21401);
nor U23329 (N_23329,N_21731,N_21332);
nand U23330 (N_23330,N_21330,N_21517);
xor U23331 (N_23331,N_21550,N_21892);
or U23332 (N_23332,N_21871,N_21847);
nor U23333 (N_23333,N_21907,N_21381);
or U23334 (N_23334,N_22340,N_22075);
nand U23335 (N_23335,N_21391,N_22429);
nand U23336 (N_23336,N_21986,N_21874);
xor U23337 (N_23337,N_21427,N_21351);
nand U23338 (N_23338,N_21545,N_21273);
nand U23339 (N_23339,N_21530,N_22419);
nor U23340 (N_23340,N_22237,N_22341);
nor U23341 (N_23341,N_21254,N_21275);
or U23342 (N_23342,N_21443,N_22154);
or U23343 (N_23343,N_21437,N_21773);
xnor U23344 (N_23344,N_22313,N_22115);
or U23345 (N_23345,N_21811,N_22446);
or U23346 (N_23346,N_21842,N_21796);
or U23347 (N_23347,N_21263,N_21606);
and U23348 (N_23348,N_22019,N_22036);
xnor U23349 (N_23349,N_21920,N_21482);
xnor U23350 (N_23350,N_21890,N_21270);
xnor U23351 (N_23351,N_21272,N_21880);
xnor U23352 (N_23352,N_21849,N_22283);
nand U23353 (N_23353,N_21577,N_21698);
nor U23354 (N_23354,N_21676,N_21427);
nand U23355 (N_23355,N_21711,N_22022);
nor U23356 (N_23356,N_22488,N_21956);
xor U23357 (N_23357,N_21935,N_22377);
nor U23358 (N_23358,N_21420,N_21956);
or U23359 (N_23359,N_21586,N_22366);
and U23360 (N_23360,N_21810,N_21602);
or U23361 (N_23361,N_22012,N_21942);
and U23362 (N_23362,N_21576,N_22013);
xnor U23363 (N_23363,N_21295,N_21534);
or U23364 (N_23364,N_22486,N_21917);
xnor U23365 (N_23365,N_21325,N_21838);
and U23366 (N_23366,N_21719,N_22335);
nor U23367 (N_23367,N_21884,N_21595);
xor U23368 (N_23368,N_21857,N_21778);
nand U23369 (N_23369,N_21932,N_21717);
and U23370 (N_23370,N_21584,N_22427);
nand U23371 (N_23371,N_22402,N_22035);
nor U23372 (N_23372,N_22400,N_21515);
or U23373 (N_23373,N_21916,N_22449);
or U23374 (N_23374,N_22333,N_21532);
nand U23375 (N_23375,N_21879,N_21636);
xor U23376 (N_23376,N_21605,N_22447);
and U23377 (N_23377,N_21730,N_21738);
and U23378 (N_23378,N_22423,N_21886);
or U23379 (N_23379,N_21296,N_21349);
xnor U23380 (N_23380,N_21653,N_21844);
nor U23381 (N_23381,N_22311,N_22388);
nor U23382 (N_23382,N_22010,N_22268);
nand U23383 (N_23383,N_21660,N_21395);
and U23384 (N_23384,N_21674,N_21578);
or U23385 (N_23385,N_21522,N_21867);
nor U23386 (N_23386,N_22287,N_21630);
nor U23387 (N_23387,N_22216,N_22377);
and U23388 (N_23388,N_21532,N_21356);
xnor U23389 (N_23389,N_22338,N_22013);
xor U23390 (N_23390,N_21761,N_21370);
or U23391 (N_23391,N_22307,N_21282);
or U23392 (N_23392,N_22344,N_22416);
nand U23393 (N_23393,N_21610,N_21644);
or U23394 (N_23394,N_22493,N_21492);
nor U23395 (N_23395,N_21687,N_21558);
nand U23396 (N_23396,N_21879,N_21347);
nor U23397 (N_23397,N_22055,N_21901);
nor U23398 (N_23398,N_21987,N_22154);
and U23399 (N_23399,N_21315,N_22076);
nand U23400 (N_23400,N_21709,N_22128);
and U23401 (N_23401,N_21893,N_21712);
xor U23402 (N_23402,N_22344,N_22401);
or U23403 (N_23403,N_21301,N_21468);
or U23404 (N_23404,N_21253,N_21487);
and U23405 (N_23405,N_21541,N_21422);
nand U23406 (N_23406,N_21875,N_22229);
nor U23407 (N_23407,N_22241,N_22232);
xor U23408 (N_23408,N_21382,N_21835);
or U23409 (N_23409,N_21750,N_22489);
xnor U23410 (N_23410,N_21731,N_21581);
nand U23411 (N_23411,N_22126,N_21713);
and U23412 (N_23412,N_22126,N_21627);
or U23413 (N_23413,N_22010,N_22393);
and U23414 (N_23414,N_22285,N_21623);
xor U23415 (N_23415,N_21925,N_21755);
or U23416 (N_23416,N_22122,N_21368);
nand U23417 (N_23417,N_21509,N_22476);
xor U23418 (N_23418,N_21956,N_21755);
nor U23419 (N_23419,N_21940,N_21505);
nand U23420 (N_23420,N_22205,N_21524);
xnor U23421 (N_23421,N_22335,N_21491);
and U23422 (N_23422,N_21313,N_22102);
xnor U23423 (N_23423,N_21937,N_21671);
nor U23424 (N_23424,N_21399,N_21501);
and U23425 (N_23425,N_21648,N_22416);
nand U23426 (N_23426,N_22414,N_21677);
nand U23427 (N_23427,N_21704,N_22250);
nand U23428 (N_23428,N_21479,N_21877);
or U23429 (N_23429,N_21515,N_22389);
nor U23430 (N_23430,N_22208,N_21769);
and U23431 (N_23431,N_21875,N_21375);
or U23432 (N_23432,N_21864,N_21957);
xor U23433 (N_23433,N_21990,N_21510);
xor U23434 (N_23434,N_22112,N_21730);
and U23435 (N_23435,N_21599,N_21397);
or U23436 (N_23436,N_21895,N_21512);
and U23437 (N_23437,N_21715,N_21496);
xnor U23438 (N_23438,N_21288,N_21407);
xor U23439 (N_23439,N_21428,N_21271);
nor U23440 (N_23440,N_21909,N_21444);
or U23441 (N_23441,N_22420,N_21473);
nand U23442 (N_23442,N_22316,N_22470);
or U23443 (N_23443,N_21354,N_21412);
and U23444 (N_23444,N_21721,N_21285);
xor U23445 (N_23445,N_21359,N_22150);
xor U23446 (N_23446,N_21444,N_22474);
nor U23447 (N_23447,N_22017,N_21512);
nor U23448 (N_23448,N_21390,N_21319);
xnor U23449 (N_23449,N_21458,N_21597);
or U23450 (N_23450,N_21661,N_21361);
or U23451 (N_23451,N_21300,N_21652);
or U23452 (N_23452,N_22351,N_21723);
and U23453 (N_23453,N_22392,N_21648);
and U23454 (N_23454,N_21832,N_21346);
nor U23455 (N_23455,N_22238,N_22222);
nand U23456 (N_23456,N_21387,N_21420);
or U23457 (N_23457,N_21853,N_21981);
xor U23458 (N_23458,N_21820,N_21844);
nor U23459 (N_23459,N_22203,N_21472);
nand U23460 (N_23460,N_22369,N_22263);
nand U23461 (N_23461,N_21725,N_22436);
or U23462 (N_23462,N_22113,N_22293);
or U23463 (N_23463,N_22241,N_21680);
nand U23464 (N_23464,N_22481,N_21629);
nor U23465 (N_23465,N_21877,N_22024);
or U23466 (N_23466,N_21368,N_22353);
nand U23467 (N_23467,N_21542,N_21498);
or U23468 (N_23468,N_21662,N_21844);
nand U23469 (N_23469,N_22370,N_22493);
xor U23470 (N_23470,N_21812,N_22486);
and U23471 (N_23471,N_22042,N_22056);
or U23472 (N_23472,N_21610,N_22086);
or U23473 (N_23473,N_22103,N_21448);
nand U23474 (N_23474,N_21737,N_22108);
xor U23475 (N_23475,N_21894,N_21390);
nor U23476 (N_23476,N_21450,N_21842);
xnor U23477 (N_23477,N_21884,N_22168);
or U23478 (N_23478,N_21474,N_21761);
nor U23479 (N_23479,N_21327,N_22333);
or U23480 (N_23480,N_21771,N_22405);
nor U23481 (N_23481,N_21521,N_22097);
xor U23482 (N_23482,N_21457,N_21665);
nand U23483 (N_23483,N_21254,N_21346);
or U23484 (N_23484,N_22453,N_22362);
or U23485 (N_23485,N_21966,N_22174);
or U23486 (N_23486,N_22271,N_22380);
xnor U23487 (N_23487,N_22023,N_21966);
xnor U23488 (N_23488,N_21887,N_21664);
nor U23489 (N_23489,N_22040,N_22295);
or U23490 (N_23490,N_21588,N_21270);
nand U23491 (N_23491,N_21728,N_22452);
xor U23492 (N_23492,N_21987,N_22456);
nor U23493 (N_23493,N_21816,N_22484);
nor U23494 (N_23494,N_22377,N_22287);
and U23495 (N_23495,N_21894,N_22233);
nand U23496 (N_23496,N_21743,N_21581);
nand U23497 (N_23497,N_22316,N_22396);
xor U23498 (N_23498,N_21987,N_21942);
or U23499 (N_23499,N_21634,N_21982);
nand U23500 (N_23500,N_21722,N_21498);
nand U23501 (N_23501,N_22023,N_22070);
xor U23502 (N_23502,N_21713,N_21954);
and U23503 (N_23503,N_21340,N_21783);
xnor U23504 (N_23504,N_21327,N_22366);
xor U23505 (N_23505,N_21273,N_22183);
and U23506 (N_23506,N_21943,N_22338);
or U23507 (N_23507,N_22173,N_22026);
xnor U23508 (N_23508,N_22344,N_22268);
nor U23509 (N_23509,N_22309,N_22239);
and U23510 (N_23510,N_22455,N_21694);
nor U23511 (N_23511,N_22013,N_22196);
nand U23512 (N_23512,N_22139,N_21462);
nand U23513 (N_23513,N_21696,N_22160);
nor U23514 (N_23514,N_22128,N_22437);
nand U23515 (N_23515,N_21497,N_21907);
nor U23516 (N_23516,N_21749,N_21643);
and U23517 (N_23517,N_22113,N_22408);
nor U23518 (N_23518,N_22225,N_21364);
or U23519 (N_23519,N_21981,N_22013);
nand U23520 (N_23520,N_22317,N_21921);
nand U23521 (N_23521,N_22296,N_21794);
and U23522 (N_23522,N_21526,N_21403);
nand U23523 (N_23523,N_22027,N_22149);
xnor U23524 (N_23524,N_22202,N_22352);
nor U23525 (N_23525,N_22111,N_21803);
nor U23526 (N_23526,N_22027,N_21866);
and U23527 (N_23527,N_21559,N_21876);
and U23528 (N_23528,N_22454,N_21806);
or U23529 (N_23529,N_22011,N_22254);
xor U23530 (N_23530,N_21802,N_22316);
xor U23531 (N_23531,N_21946,N_21974);
xor U23532 (N_23532,N_22266,N_22198);
xnor U23533 (N_23533,N_21436,N_21589);
nand U23534 (N_23534,N_21616,N_21396);
and U23535 (N_23535,N_21800,N_22317);
xor U23536 (N_23536,N_22344,N_22393);
nand U23537 (N_23537,N_21539,N_21781);
nand U23538 (N_23538,N_22098,N_22152);
and U23539 (N_23539,N_21317,N_22023);
nor U23540 (N_23540,N_21454,N_21575);
and U23541 (N_23541,N_21726,N_21684);
nor U23542 (N_23542,N_22280,N_21586);
xnor U23543 (N_23543,N_21579,N_22459);
and U23544 (N_23544,N_21538,N_21371);
nand U23545 (N_23545,N_21800,N_21256);
nand U23546 (N_23546,N_22034,N_21530);
nor U23547 (N_23547,N_21946,N_21581);
and U23548 (N_23548,N_21677,N_22072);
or U23549 (N_23549,N_22096,N_21761);
nand U23550 (N_23550,N_21868,N_22262);
nor U23551 (N_23551,N_22007,N_22326);
nor U23552 (N_23552,N_21807,N_21551);
or U23553 (N_23553,N_21815,N_21888);
xor U23554 (N_23554,N_22180,N_22482);
xor U23555 (N_23555,N_21383,N_22412);
and U23556 (N_23556,N_21327,N_21515);
xor U23557 (N_23557,N_21742,N_21905);
nor U23558 (N_23558,N_21963,N_21638);
or U23559 (N_23559,N_21548,N_22343);
nand U23560 (N_23560,N_22143,N_21259);
and U23561 (N_23561,N_21446,N_21365);
and U23562 (N_23562,N_21587,N_21886);
nand U23563 (N_23563,N_22489,N_21288);
xor U23564 (N_23564,N_21832,N_21943);
or U23565 (N_23565,N_21275,N_21475);
and U23566 (N_23566,N_22485,N_21316);
nor U23567 (N_23567,N_21846,N_21839);
or U23568 (N_23568,N_21722,N_21806);
xor U23569 (N_23569,N_22269,N_22200);
nor U23570 (N_23570,N_21667,N_22328);
nand U23571 (N_23571,N_21678,N_21547);
nor U23572 (N_23572,N_22309,N_21649);
xor U23573 (N_23573,N_22221,N_21747);
nor U23574 (N_23574,N_22466,N_21831);
xnor U23575 (N_23575,N_22320,N_21709);
nand U23576 (N_23576,N_21420,N_22185);
nand U23577 (N_23577,N_21955,N_21476);
or U23578 (N_23578,N_22116,N_21820);
nand U23579 (N_23579,N_21809,N_22250);
or U23580 (N_23580,N_21784,N_21825);
and U23581 (N_23581,N_21265,N_21901);
or U23582 (N_23582,N_22091,N_21447);
nor U23583 (N_23583,N_22136,N_21970);
xor U23584 (N_23584,N_21560,N_21324);
xor U23585 (N_23585,N_22236,N_21399);
or U23586 (N_23586,N_21549,N_21823);
and U23587 (N_23587,N_21611,N_22006);
xor U23588 (N_23588,N_21685,N_21309);
or U23589 (N_23589,N_21882,N_21563);
nor U23590 (N_23590,N_22313,N_21418);
xnor U23591 (N_23591,N_21720,N_21432);
nand U23592 (N_23592,N_22056,N_22111);
and U23593 (N_23593,N_22496,N_21385);
nor U23594 (N_23594,N_21479,N_21375);
xor U23595 (N_23595,N_21581,N_22210);
and U23596 (N_23596,N_21555,N_21357);
xnor U23597 (N_23597,N_21864,N_21460);
nor U23598 (N_23598,N_22469,N_22275);
nand U23599 (N_23599,N_22325,N_21975);
and U23600 (N_23600,N_21582,N_21580);
xor U23601 (N_23601,N_22245,N_21584);
or U23602 (N_23602,N_22012,N_22318);
nand U23603 (N_23603,N_22483,N_22236);
nor U23604 (N_23604,N_21663,N_21767);
or U23605 (N_23605,N_21343,N_22040);
nand U23606 (N_23606,N_22256,N_21520);
or U23607 (N_23607,N_22131,N_21573);
or U23608 (N_23608,N_21772,N_21901);
nor U23609 (N_23609,N_22357,N_22139);
and U23610 (N_23610,N_21827,N_22441);
nand U23611 (N_23611,N_22317,N_22481);
nand U23612 (N_23612,N_22208,N_22042);
or U23613 (N_23613,N_21416,N_22137);
or U23614 (N_23614,N_21608,N_21833);
and U23615 (N_23615,N_21513,N_22198);
or U23616 (N_23616,N_21532,N_21479);
and U23617 (N_23617,N_21836,N_21979);
nor U23618 (N_23618,N_22104,N_21646);
nor U23619 (N_23619,N_21997,N_21413);
nand U23620 (N_23620,N_22493,N_21286);
or U23621 (N_23621,N_21563,N_21395);
nor U23622 (N_23622,N_21755,N_21852);
xor U23623 (N_23623,N_21760,N_21908);
or U23624 (N_23624,N_22394,N_21794);
nor U23625 (N_23625,N_22157,N_21416);
nand U23626 (N_23626,N_21406,N_22215);
xnor U23627 (N_23627,N_21956,N_22286);
nor U23628 (N_23628,N_22022,N_22111);
and U23629 (N_23629,N_21457,N_22252);
xnor U23630 (N_23630,N_22332,N_22021);
nor U23631 (N_23631,N_21424,N_22373);
nand U23632 (N_23632,N_22027,N_21923);
xor U23633 (N_23633,N_21747,N_22297);
or U23634 (N_23634,N_21822,N_21896);
nor U23635 (N_23635,N_22001,N_21687);
and U23636 (N_23636,N_21798,N_21431);
nor U23637 (N_23637,N_22115,N_21944);
or U23638 (N_23638,N_22117,N_21938);
nor U23639 (N_23639,N_21351,N_22497);
or U23640 (N_23640,N_21275,N_21551);
xor U23641 (N_23641,N_22001,N_21926);
and U23642 (N_23642,N_22231,N_21422);
or U23643 (N_23643,N_21610,N_21972);
nor U23644 (N_23644,N_21333,N_22150);
nand U23645 (N_23645,N_21852,N_22304);
xor U23646 (N_23646,N_21250,N_21263);
and U23647 (N_23647,N_22451,N_22109);
nand U23648 (N_23648,N_22054,N_21321);
nand U23649 (N_23649,N_22193,N_21318);
nor U23650 (N_23650,N_21747,N_21848);
and U23651 (N_23651,N_22098,N_21861);
nand U23652 (N_23652,N_22185,N_21857);
xnor U23653 (N_23653,N_21717,N_22426);
or U23654 (N_23654,N_22126,N_21814);
nand U23655 (N_23655,N_22204,N_22008);
nand U23656 (N_23656,N_22288,N_21997);
and U23657 (N_23657,N_22024,N_22173);
nand U23658 (N_23658,N_21793,N_22065);
or U23659 (N_23659,N_22457,N_21964);
and U23660 (N_23660,N_21326,N_22176);
nand U23661 (N_23661,N_22373,N_21318);
xnor U23662 (N_23662,N_21867,N_22092);
or U23663 (N_23663,N_22309,N_21720);
nor U23664 (N_23664,N_22393,N_21484);
and U23665 (N_23665,N_21375,N_21315);
xnor U23666 (N_23666,N_21977,N_22143);
and U23667 (N_23667,N_21577,N_22113);
or U23668 (N_23668,N_22271,N_21920);
nand U23669 (N_23669,N_22154,N_21493);
nand U23670 (N_23670,N_21979,N_21921);
nor U23671 (N_23671,N_21951,N_21593);
nor U23672 (N_23672,N_21624,N_21389);
nor U23673 (N_23673,N_21828,N_22026);
xor U23674 (N_23674,N_22015,N_22084);
and U23675 (N_23675,N_22229,N_21595);
or U23676 (N_23676,N_22411,N_21366);
xor U23677 (N_23677,N_21828,N_21707);
or U23678 (N_23678,N_21605,N_21548);
xnor U23679 (N_23679,N_21537,N_21367);
and U23680 (N_23680,N_21719,N_21434);
nand U23681 (N_23681,N_21405,N_21476);
nand U23682 (N_23682,N_22225,N_21974);
or U23683 (N_23683,N_22360,N_21588);
and U23684 (N_23684,N_21826,N_21701);
or U23685 (N_23685,N_21839,N_22198);
xor U23686 (N_23686,N_21476,N_22194);
nand U23687 (N_23687,N_21535,N_21771);
xor U23688 (N_23688,N_21605,N_22059);
or U23689 (N_23689,N_21940,N_21633);
xor U23690 (N_23690,N_21758,N_21785);
xnor U23691 (N_23691,N_21648,N_21678);
and U23692 (N_23692,N_21696,N_21564);
xor U23693 (N_23693,N_22046,N_22325);
and U23694 (N_23694,N_21302,N_21449);
or U23695 (N_23695,N_21633,N_22121);
xor U23696 (N_23696,N_21995,N_22351);
or U23697 (N_23697,N_21615,N_21638);
and U23698 (N_23698,N_21868,N_21513);
nor U23699 (N_23699,N_21784,N_22078);
nand U23700 (N_23700,N_21628,N_22135);
nor U23701 (N_23701,N_22294,N_21769);
xor U23702 (N_23702,N_21635,N_21557);
xor U23703 (N_23703,N_22365,N_22447);
xor U23704 (N_23704,N_22198,N_22067);
xnor U23705 (N_23705,N_22102,N_21986);
nor U23706 (N_23706,N_21586,N_21354);
and U23707 (N_23707,N_21479,N_22225);
nand U23708 (N_23708,N_21709,N_21893);
nand U23709 (N_23709,N_22316,N_21968);
nand U23710 (N_23710,N_21882,N_22373);
and U23711 (N_23711,N_21865,N_21700);
nand U23712 (N_23712,N_21763,N_22240);
nor U23713 (N_23713,N_22180,N_21580);
or U23714 (N_23714,N_21719,N_22427);
nor U23715 (N_23715,N_22024,N_21963);
xor U23716 (N_23716,N_22102,N_22469);
nand U23717 (N_23717,N_22209,N_22158);
and U23718 (N_23718,N_22297,N_21731);
xnor U23719 (N_23719,N_21805,N_21511);
nor U23720 (N_23720,N_21970,N_21575);
nand U23721 (N_23721,N_21965,N_21327);
or U23722 (N_23722,N_21379,N_21294);
or U23723 (N_23723,N_22414,N_21689);
xnor U23724 (N_23724,N_21991,N_22206);
and U23725 (N_23725,N_21767,N_22145);
or U23726 (N_23726,N_22241,N_22292);
nor U23727 (N_23727,N_22153,N_22262);
and U23728 (N_23728,N_22176,N_22437);
xor U23729 (N_23729,N_22365,N_21386);
xnor U23730 (N_23730,N_22449,N_21572);
or U23731 (N_23731,N_22012,N_22246);
xnor U23732 (N_23732,N_21386,N_21970);
xnor U23733 (N_23733,N_22028,N_21772);
or U23734 (N_23734,N_22064,N_22014);
and U23735 (N_23735,N_21475,N_22022);
nand U23736 (N_23736,N_21912,N_21575);
or U23737 (N_23737,N_21898,N_22233);
xor U23738 (N_23738,N_21332,N_22357);
nand U23739 (N_23739,N_22177,N_21324);
and U23740 (N_23740,N_21409,N_22343);
nand U23741 (N_23741,N_21746,N_22292);
or U23742 (N_23742,N_22127,N_21552);
nand U23743 (N_23743,N_22263,N_21658);
nand U23744 (N_23744,N_21422,N_22423);
nor U23745 (N_23745,N_22215,N_22286);
or U23746 (N_23746,N_21775,N_21702);
and U23747 (N_23747,N_21874,N_21763);
and U23748 (N_23748,N_22049,N_22316);
and U23749 (N_23749,N_21815,N_22024);
nor U23750 (N_23750,N_22814,N_23178);
nand U23751 (N_23751,N_22561,N_23592);
xor U23752 (N_23752,N_22826,N_23033);
xor U23753 (N_23753,N_23399,N_23478);
xnor U23754 (N_23754,N_22860,N_23097);
xnor U23755 (N_23755,N_23749,N_22861);
and U23756 (N_23756,N_23093,N_23320);
xor U23757 (N_23757,N_23070,N_23725);
and U23758 (N_23758,N_23104,N_23356);
and U23759 (N_23759,N_22889,N_23305);
and U23760 (N_23760,N_23148,N_22977);
nand U23761 (N_23761,N_22936,N_23415);
xor U23762 (N_23762,N_23105,N_22575);
nand U23763 (N_23763,N_22985,N_22953);
nor U23764 (N_23764,N_23522,N_23740);
nand U23765 (N_23765,N_22836,N_23298);
nand U23766 (N_23766,N_23466,N_22669);
nand U23767 (N_23767,N_23184,N_22552);
and U23768 (N_23768,N_22980,N_22941);
nor U23769 (N_23769,N_23718,N_22940);
nand U23770 (N_23770,N_23677,N_22984);
nor U23771 (N_23771,N_22998,N_22511);
and U23772 (N_23772,N_22965,N_23712);
nor U23773 (N_23773,N_23682,N_23265);
nor U23774 (N_23774,N_23433,N_22642);
or U23775 (N_23775,N_22793,N_22791);
nor U23776 (N_23776,N_23479,N_22920);
and U23777 (N_23777,N_23678,N_23338);
nor U23778 (N_23778,N_22990,N_23539);
xor U23779 (N_23779,N_23542,N_22877);
or U23780 (N_23780,N_22858,N_23568);
xor U23781 (N_23781,N_23620,N_23589);
xnor U23782 (N_23782,N_22755,N_23458);
or U23783 (N_23783,N_22570,N_23680);
nand U23784 (N_23784,N_23556,N_23639);
nand U23785 (N_23785,N_22677,N_23003);
xnor U23786 (N_23786,N_22944,N_23333);
nand U23787 (N_23787,N_23497,N_22875);
nor U23788 (N_23788,N_23714,N_23100);
and U23789 (N_23789,N_23444,N_23624);
xor U23790 (N_23790,N_22686,N_22651);
nor U23791 (N_23791,N_23613,N_22942);
xor U23792 (N_23792,N_22528,N_22750);
and U23793 (N_23793,N_22892,N_22736);
or U23794 (N_23794,N_22547,N_23622);
nand U23795 (N_23795,N_23741,N_23660);
xnor U23796 (N_23796,N_23641,N_22807);
or U23797 (N_23797,N_23135,N_22572);
and U23798 (N_23798,N_22979,N_23482);
nor U23799 (N_23799,N_23061,N_23745);
nand U23800 (N_23800,N_23658,N_23189);
and U23801 (N_23801,N_22598,N_22630);
or U23802 (N_23802,N_23457,N_22662);
nor U23803 (N_23803,N_23101,N_23566);
nor U23804 (N_23804,N_22676,N_23552);
and U23805 (N_23805,N_23309,N_22742);
xor U23806 (N_23806,N_22830,N_23180);
nand U23807 (N_23807,N_23359,N_23448);
nand U23808 (N_23808,N_22696,N_23087);
xor U23809 (N_23809,N_23263,N_22746);
and U23810 (N_23810,N_22524,N_22852);
or U23811 (N_23811,N_22579,N_23285);
or U23812 (N_23812,N_23232,N_23160);
or U23813 (N_23813,N_23273,N_22612);
nor U23814 (N_23814,N_23260,N_23605);
and U23815 (N_23815,N_23630,N_23106);
nand U23816 (N_23816,N_22603,N_23102);
and U23817 (N_23817,N_23084,N_23591);
xnor U23818 (N_23818,N_23029,N_23256);
xor U23819 (N_23819,N_23158,N_23242);
or U23820 (N_23820,N_23570,N_22619);
or U23821 (N_23821,N_23673,N_23295);
xnor U23822 (N_23822,N_23372,N_23430);
or U23823 (N_23823,N_23472,N_23137);
nor U23824 (N_23824,N_23109,N_22683);
nor U23825 (N_23825,N_22799,N_23512);
and U23826 (N_23826,N_22681,N_23058);
and U23827 (N_23827,N_22781,N_22695);
nor U23828 (N_23828,N_23253,N_23411);
nand U23829 (N_23829,N_23728,N_22749);
nand U23830 (N_23830,N_22866,N_23549);
and U23831 (N_23831,N_23202,N_22777);
or U23832 (N_23832,N_23557,N_23145);
or U23833 (N_23833,N_22548,N_23516);
nor U23834 (N_23834,N_23244,N_23737);
xor U23835 (N_23835,N_23386,N_23590);
nor U23836 (N_23836,N_23593,N_22650);
and U23837 (N_23837,N_23354,N_22805);
nor U23838 (N_23838,N_23079,N_22520);
or U23839 (N_23839,N_23429,N_23417);
xnor U23840 (N_23840,N_22706,N_23606);
or U23841 (N_23841,N_23318,N_23648);
nand U23842 (N_23842,N_23390,N_23743);
and U23843 (N_23843,N_23609,N_22752);
or U23844 (N_23844,N_22559,N_23396);
and U23845 (N_23845,N_23428,N_23443);
nand U23846 (N_23846,N_22823,N_22949);
xnor U23847 (N_23847,N_23272,N_23629);
and U23848 (N_23848,N_23200,N_23492);
or U23849 (N_23849,N_22933,N_23564);
nand U23850 (N_23850,N_23048,N_23530);
nand U23851 (N_23851,N_22978,N_23614);
nor U23852 (N_23852,N_22734,N_23695);
or U23853 (N_23853,N_22756,N_23579);
nor U23854 (N_23854,N_23481,N_22664);
xor U23855 (N_23855,N_22809,N_23451);
nand U23856 (N_23856,N_23014,N_22928);
or U23857 (N_23857,N_23550,N_23240);
nor U23858 (N_23858,N_23423,N_22813);
xnor U23859 (N_23859,N_22899,N_22989);
or U23860 (N_23860,N_23360,N_23267);
or U23861 (N_23861,N_23005,N_23581);
and U23862 (N_23862,N_23604,N_23308);
nor U23863 (N_23863,N_23069,N_23221);
nand U23864 (N_23864,N_22895,N_22788);
nor U23865 (N_23865,N_22568,N_23602);
nand U23866 (N_23866,N_23529,N_22615);
nand U23867 (N_23867,N_22613,N_22586);
xor U23868 (N_23868,N_23111,N_23340);
nor U23869 (N_23869,N_22567,N_22714);
or U23870 (N_23870,N_22689,N_22710);
nand U23871 (N_23871,N_22810,N_22565);
or U23872 (N_23872,N_23616,N_22842);
and U23873 (N_23873,N_22956,N_23282);
and U23874 (N_23874,N_22685,N_23045);
nand U23875 (N_23875,N_22735,N_23508);
or U23876 (N_23876,N_22782,N_23526);
xor U23877 (N_23877,N_23450,N_22691);
or U23878 (N_23878,N_23726,N_22825);
nand U23879 (N_23879,N_22578,N_22897);
nor U23880 (N_23880,N_23537,N_23352);
xor U23881 (N_23881,N_23693,N_23531);
or U23882 (N_23882,N_22702,N_23357);
xnor U23883 (N_23883,N_22566,N_23075);
and U23884 (N_23884,N_22549,N_23153);
and U23885 (N_23885,N_23435,N_23012);
or U23886 (N_23886,N_23652,N_23043);
or U23887 (N_23887,N_23215,N_23599);
nand U23888 (N_23888,N_23204,N_23144);
xnor U23889 (N_23889,N_22886,N_22994);
xnor U23890 (N_23890,N_23013,N_22607);
xor U23891 (N_23891,N_23057,N_23133);
or U23892 (N_23892,N_23747,N_22937);
or U23893 (N_23893,N_22917,N_22509);
and U23894 (N_23894,N_23621,N_23656);
or U23895 (N_23895,N_23227,N_22964);
xor U23896 (N_23896,N_22656,N_23649);
nor U23897 (N_23897,N_23494,N_22649);
nand U23898 (N_23898,N_22804,N_22754);
and U23899 (N_23899,N_23170,N_23578);
nand U23900 (N_23900,N_23096,N_23703);
or U23901 (N_23901,N_22594,N_23683);
xnor U23902 (N_23902,N_23329,N_23163);
nor U23903 (N_23903,N_22851,N_23248);
xnor U23904 (N_23904,N_22792,N_23518);
nand U23905 (N_23905,N_22828,N_22611);
nor U23906 (N_23906,N_23032,N_23021);
nor U23907 (N_23907,N_22834,N_23730);
nand U23908 (N_23908,N_23380,N_23532);
xor U23909 (N_23909,N_22536,N_23619);
nor U23910 (N_23910,N_23146,N_22883);
nor U23911 (N_23911,N_23638,N_23555);
xor U23912 (N_23912,N_22762,N_23073);
or U23913 (N_23913,N_23488,N_22694);
nand U23914 (N_23914,N_23464,N_22508);
nor U23915 (N_23915,N_22577,N_23724);
nor U23916 (N_23916,N_23572,N_23646);
and U23917 (N_23917,N_22801,N_23696);
nor U23918 (N_23918,N_23065,N_22705);
nand U23919 (N_23919,N_22906,N_22692);
nor U23920 (N_23920,N_23662,N_22512);
and U23921 (N_23921,N_23027,N_23195);
or U23922 (N_23922,N_22768,N_23562);
or U23923 (N_23923,N_23299,N_23569);
xnor U23924 (N_23924,N_22622,N_23262);
or U23925 (N_23925,N_23213,N_22505);
xnor U23926 (N_23926,N_22583,N_22724);
and U23927 (N_23927,N_23210,N_22659);
and U23928 (N_23928,N_23344,N_23300);
or U23929 (N_23929,N_23664,N_22885);
nand U23930 (N_23930,N_23729,N_23580);
nand U23931 (N_23931,N_23085,N_23040);
nor U23932 (N_23932,N_22966,N_23047);
and U23933 (N_23933,N_22789,N_23402);
or U23934 (N_23934,N_23440,N_23617);
or U23935 (N_23935,N_23187,N_23534);
nor U23936 (N_23936,N_23306,N_22618);
or U23937 (N_23937,N_23296,N_22873);
nand U23938 (N_23938,N_22541,N_23667);
xnor U23939 (N_23939,N_23369,N_23672);
xor U23940 (N_23940,N_22787,N_23155);
nor U23941 (N_23941,N_23080,N_22982);
and U23942 (N_23942,N_23001,N_22704);
xnor U23943 (N_23943,N_22740,N_23293);
nand U23944 (N_23944,N_22832,N_22995);
nand U23945 (N_23945,N_22530,N_22760);
and U23946 (N_23946,N_22876,N_23182);
nand U23947 (N_23947,N_22916,N_22816);
nand U23948 (N_23948,N_23722,N_22716);
or U23949 (N_23949,N_22766,N_23548);
nor U23950 (N_23950,N_22723,N_22569);
nor U23951 (N_23951,N_22661,N_22514);
nor U23952 (N_23952,N_23422,N_23460);
nor U23953 (N_23953,N_23496,N_23067);
and U23954 (N_23954,N_22688,N_22926);
and U23955 (N_23955,N_22532,N_23661);
nor U23956 (N_23956,N_22904,N_22913);
and U23957 (N_23957,N_22881,N_22604);
and U23958 (N_23958,N_23050,N_23268);
nor U23959 (N_23959,N_23387,N_23463);
nand U23960 (N_23960,N_23337,N_23132);
xnor U23961 (N_23961,N_23536,N_23071);
nand U23962 (N_23962,N_23301,N_23162);
or U23963 (N_23963,N_23596,N_23082);
xnor U23964 (N_23964,N_22890,N_22846);
and U23965 (N_23965,N_22727,N_22674);
or U23966 (N_23966,N_23078,N_23136);
xnor U23967 (N_23967,N_23194,N_22961);
nand U23968 (N_23968,N_22925,N_22513);
xor U23969 (N_23969,N_22999,N_23684);
and U23970 (N_23970,N_22856,N_22741);
nand U23971 (N_23971,N_23595,N_23710);
xor U23972 (N_23972,N_22790,N_23108);
or U23973 (N_23973,N_22693,N_22812);
and U23974 (N_23974,N_22555,N_23343);
nor U23975 (N_23975,N_23503,N_23310);
nor U23976 (N_23976,N_23023,N_22535);
nand U23977 (N_23977,N_22930,N_23420);
or U23978 (N_23978,N_23654,N_22628);
nor U23979 (N_23979,N_23666,N_23511);
xnor U23980 (N_23980,N_23236,N_23607);
xor U23981 (N_23981,N_22921,N_23383);
and U23982 (N_23982,N_22655,N_22867);
and U23983 (N_23983,N_23164,N_22663);
nor U23984 (N_23984,N_22845,N_22821);
and U23985 (N_23985,N_23375,N_23404);
and U23986 (N_23986,N_22901,N_22601);
nand U23987 (N_23987,N_23312,N_23247);
nand U23988 (N_23988,N_23188,N_23241);
or U23989 (N_23989,N_22647,N_23528);
or U23990 (N_23990,N_23363,N_22597);
nor U23991 (N_23991,N_23089,N_23510);
xor U23992 (N_23992,N_23706,N_22785);
nor U23993 (N_23993,N_22700,N_23668);
or U23994 (N_23994,N_23651,N_23545);
or U23995 (N_23995,N_23063,N_23019);
or U23996 (N_23996,N_23222,N_23351);
nand U23997 (N_23997,N_23576,N_23112);
nor U23998 (N_23998,N_22841,N_23243);
and U23999 (N_23999,N_22773,N_23092);
and U24000 (N_24000,N_23231,N_23487);
nor U24001 (N_24001,N_22938,N_23348);
xnor U24002 (N_24002,N_23173,N_23117);
nand U24003 (N_24003,N_23535,N_23397);
nor U24004 (N_24004,N_23470,N_22522);
nor U24005 (N_24005,N_23465,N_22955);
or U24006 (N_24006,N_23558,N_22697);
and U24007 (N_24007,N_23167,N_23626);
and U24008 (N_24008,N_23199,N_22639);
or U24009 (N_24009,N_23563,N_23409);
nor U24010 (N_24010,N_23715,N_23594);
nor U24011 (N_24011,N_23115,N_23573);
or U24012 (N_24012,N_23467,N_23501);
nand U24013 (N_24013,N_22797,N_23254);
or U24014 (N_24014,N_22739,N_23395);
xor U24015 (N_24015,N_23313,N_22786);
nand U24016 (N_24016,N_23468,N_22592);
or U24017 (N_24017,N_23201,N_22620);
or U24018 (N_24018,N_23461,N_22951);
and U24019 (N_24019,N_23230,N_22991);
and U24020 (N_24020,N_23723,N_23413);
and U24021 (N_24021,N_22726,N_22629);
xor U24022 (N_24022,N_23653,N_23280);
or U24023 (N_24023,N_23125,N_23416);
xor U24024 (N_24024,N_23203,N_23447);
xor U24025 (N_24025,N_23322,N_23220);
or U24026 (N_24026,N_23315,N_23017);
or U24027 (N_24027,N_22753,N_23509);
or U24028 (N_24028,N_23317,N_23355);
xnor U24029 (N_24029,N_22835,N_23471);
and U24030 (N_24030,N_22775,N_23062);
and U24031 (N_24031,N_23191,N_23186);
and U24032 (N_24032,N_22800,N_23636);
nor U24033 (N_24033,N_22763,N_23700);
or U24034 (N_24034,N_22997,N_23176);
nand U24035 (N_24035,N_22969,N_23676);
or U24036 (N_24036,N_23052,N_23055);
xnor U24037 (N_24037,N_22665,N_23190);
nor U24038 (N_24038,N_23025,N_23418);
nor U24039 (N_24039,N_23250,N_22679);
and U24040 (N_24040,N_22822,N_23367);
and U24041 (N_24041,N_23456,N_23291);
xnor U24042 (N_24042,N_23547,N_22546);
nand U24043 (N_24043,N_23628,N_23328);
nor U24044 (N_24044,N_22887,N_23165);
xor U24045 (N_24045,N_23600,N_22634);
nand U24046 (N_24046,N_23088,N_23037);
nor U24047 (N_24047,N_23571,N_23459);
or U24048 (N_24048,N_23127,N_23228);
nand U24049 (N_24049,N_22854,N_22931);
xnor U24050 (N_24050,N_23053,N_22986);
nor U24051 (N_24051,N_23270,N_23292);
xor U24052 (N_24052,N_23261,N_23642);
nor U24053 (N_24053,N_23437,N_22888);
nor U24054 (N_24054,N_23401,N_22914);
xnor U24055 (N_24055,N_22682,N_22948);
xor U24056 (N_24056,N_23166,N_23121);
or U24057 (N_24057,N_22588,N_23587);
and U24058 (N_24058,N_23392,N_23517);
and U24059 (N_24059,N_23708,N_22987);
or U24060 (N_24060,N_23640,N_23655);
and U24061 (N_24061,N_22593,N_22668);
xnor U24062 (N_24062,N_22880,N_23533);
nand U24063 (N_24063,N_23098,N_23632);
nand U24064 (N_24064,N_22958,N_22529);
xnor U24065 (N_24065,N_23634,N_23326);
xnor U24066 (N_24066,N_23103,N_23245);
nand U24067 (N_24067,N_23704,N_22929);
nand U24068 (N_24068,N_22780,N_23284);
nand U24069 (N_24069,N_23076,N_23008);
or U24070 (N_24070,N_22616,N_23018);
and U24071 (N_24071,N_22924,N_23434);
or U24072 (N_24072,N_23685,N_23505);
or U24073 (N_24073,N_23659,N_23427);
xor U24074 (N_24074,N_22729,N_23424);
nor U24075 (N_24075,N_22684,N_23026);
and U24076 (N_24076,N_23675,N_23431);
nand U24077 (N_24077,N_22507,N_23670);
nor U24078 (N_24078,N_23567,N_22640);
nor U24079 (N_24079,N_23279,N_22701);
xnor U24080 (N_24080,N_23142,N_23206);
nor U24081 (N_24081,N_23381,N_23152);
xor U24082 (N_24082,N_23633,N_22523);
and U24083 (N_24083,N_22837,N_22621);
or U24084 (N_24084,N_22759,N_22855);
nor U24085 (N_24085,N_22556,N_22962);
xor U24086 (N_24086,N_23623,N_23691);
nand U24087 (N_24087,N_23453,N_22945);
nor U24088 (N_24088,N_23469,N_23277);
nor U24089 (N_24089,N_22932,N_22974);
nor U24090 (N_24090,N_23699,N_23303);
and U24091 (N_24091,N_23311,N_22747);
or U24092 (N_24092,N_22707,N_22703);
nand U24093 (N_24093,N_22590,N_22839);
or U24094 (N_24094,N_22779,N_22770);
and U24095 (N_24095,N_22973,N_22527);
or U24096 (N_24096,N_23702,N_22796);
nand U24097 (N_24097,N_23538,N_23185);
nand U24098 (N_24098,N_22908,N_23376);
xor U24099 (N_24099,N_22859,N_23504);
and U24100 (N_24100,N_23218,N_23031);
nand U24101 (N_24101,N_22952,N_22554);
or U24102 (N_24102,N_23156,N_22582);
nor U24103 (N_24103,N_23056,N_22719);
xnor U24104 (N_24104,N_22539,N_23233);
nor U24105 (N_24105,N_23412,N_23034);
and U24106 (N_24106,N_23574,N_22981);
nand U24107 (N_24107,N_22819,N_23251);
or U24108 (N_24108,N_22660,N_22580);
nand U24109 (N_24109,N_23332,N_23224);
and U24110 (N_24110,N_22690,N_23389);
xnor U24111 (N_24111,N_23319,N_22820);
xnor U24112 (N_24112,N_23382,N_22843);
nor U24113 (N_24113,N_22874,N_23257);
and U24114 (N_24114,N_22894,N_22672);
and U24115 (N_24115,N_22960,N_22784);
or U24116 (N_24116,N_22503,N_23197);
and U24117 (N_24117,N_23283,N_23582);
xnor U24118 (N_24118,N_23588,N_23400);
or U24119 (N_24119,N_23287,N_23364);
and U24120 (N_24120,N_23339,N_23362);
xor U24121 (N_24121,N_22817,N_22811);
and U24122 (N_24122,N_22738,N_22648);
xnor U24123 (N_24123,N_22840,N_23631);
nor U24124 (N_24124,N_23738,N_23225);
nand U24125 (N_24125,N_23368,N_22946);
or U24126 (N_24126,N_23114,N_23095);
nand U24127 (N_24127,N_22896,N_22833);
or U24128 (N_24128,N_22870,N_23347);
or U24129 (N_24129,N_23583,N_23502);
nand U24130 (N_24130,N_23331,N_23341);
or U24131 (N_24131,N_23216,N_23692);
and U24132 (N_24132,N_23346,N_22538);
nand U24133 (N_24133,N_23543,N_22993);
xor U24134 (N_24134,N_22708,N_23110);
nand U24135 (N_24135,N_22608,N_23499);
or U24136 (N_24136,N_23325,N_23748);
or U24137 (N_24137,N_23011,N_23697);
nand U24138 (N_24138,N_23246,N_22614);
nand U24139 (N_24139,N_23377,N_23081);
nor U24140 (N_24140,N_22517,N_22776);
xnor U24141 (N_24141,N_22687,N_23374);
xnor U24142 (N_24142,N_22605,N_23371);
and U24143 (N_24143,N_23120,N_23419);
and U24144 (N_24144,N_23403,N_23689);
nand U24145 (N_24145,N_23577,N_22518);
xnor U24146 (N_24146,N_22943,N_23235);
or U24147 (N_24147,N_23441,N_23015);
or U24148 (N_24148,N_23159,N_22627);
or U24149 (N_24149,N_22778,N_23006);
or U24150 (N_24150,N_23480,N_22502);
or U24151 (N_24151,N_22666,N_23681);
or U24152 (N_24152,N_22927,N_23615);
nor U24153 (N_24153,N_23131,N_22774);
nand U24154 (N_24154,N_23211,N_22562);
nand U24155 (N_24155,N_23414,N_23330);
or U24156 (N_24156,N_22996,N_23177);
or U24157 (N_24157,N_22862,N_23736);
nand U24158 (N_24158,N_23183,N_22519);
and U24159 (N_24159,N_22632,N_23735);
and U24160 (N_24160,N_23426,N_22879);
nand U24161 (N_24161,N_23205,N_23407);
or U24162 (N_24162,N_23669,N_23719);
nor U24163 (N_24163,N_23671,N_22783);
nor U24164 (N_24164,N_22950,N_23147);
nor U24165 (N_24165,N_22715,N_23687);
and U24166 (N_24166,N_22911,N_22652);
and U24167 (N_24167,N_23234,N_22954);
and U24168 (N_24168,N_22806,N_22882);
nor U24169 (N_24169,N_22847,N_23514);
or U24170 (N_24170,N_23525,N_22543);
nor U24171 (N_24171,N_22803,N_22721);
xnor U24172 (N_24172,N_23515,N_22553);
xor U24173 (N_24173,N_23122,N_23314);
nand U24174 (N_24174,N_23643,N_22970);
nand U24175 (N_24175,N_23408,N_23091);
nand U24176 (N_24176,N_22560,N_22902);
or U24177 (N_24177,N_23172,N_23610);
nor U24178 (N_24178,N_23139,N_23732);
nand U24179 (N_24179,N_23321,N_23004);
nand U24180 (N_24180,N_22678,N_22872);
and U24181 (N_24181,N_23546,N_23174);
xnor U24182 (N_24182,N_22827,N_23000);
nor U24183 (N_24183,N_22959,N_22534);
and U24184 (N_24184,N_23255,N_23193);
nand U24185 (N_24185,N_23405,N_23495);
xor U24186 (N_24186,N_22574,N_22891);
nor U24187 (N_24187,N_23690,N_23727);
and U24188 (N_24188,N_23289,N_23214);
nand U24189 (N_24189,N_23039,N_22844);
nor U24190 (N_24190,N_22849,N_22521);
xnor U24191 (N_24191,N_23157,N_23198);
xnor U24192 (N_24192,N_23625,N_22798);
nor U24193 (N_24193,N_23462,N_22657);
and U24194 (N_24194,N_23711,N_22884);
xnor U24195 (N_24195,N_22531,N_23421);
nor U24196 (N_24196,N_23541,N_23384);
and U24197 (N_24197,N_23490,N_23540);
or U24198 (N_24198,N_23009,N_23278);
nor U24199 (N_24199,N_22915,N_22646);
and U24200 (N_24200,N_22900,N_23028);
and U24201 (N_24201,N_22767,N_22635);
and U24202 (N_24202,N_23288,N_22935);
and U24203 (N_24203,N_22626,N_23140);
nor U24204 (N_24204,N_22699,N_22510);
xor U24205 (N_24205,N_23559,N_23698);
and U24206 (N_24206,N_22500,N_23281);
nor U24207 (N_24207,N_22863,N_23324);
xor U24208 (N_24208,N_23138,N_22525);
and U24209 (N_24209,N_23143,N_23679);
or U24210 (N_24210,N_23597,N_22831);
nand U24211 (N_24211,N_23438,N_23406);
or U24212 (N_24212,N_22641,N_22624);
or U24213 (N_24213,N_23523,N_23474);
and U24214 (N_24214,N_23030,N_22599);
xnor U24215 (N_24215,N_23500,N_22963);
nor U24216 (N_24216,N_22838,N_23196);
or U24217 (N_24217,N_23051,N_22595);
nand U24218 (N_24218,N_23713,N_22713);
nand U24219 (N_24219,N_23665,N_23192);
and U24220 (N_24220,N_22898,N_23521);
xor U24221 (N_24221,N_23650,N_22636);
xnor U24222 (N_24222,N_22585,N_22829);
nand U24223 (N_24223,N_23393,N_22732);
and U24224 (N_24224,N_23618,N_22564);
nor U24225 (N_24225,N_23686,N_23601);
and U24226 (N_24226,N_23739,N_23020);
nor U24227 (N_24227,N_23335,N_23113);
nor U24228 (N_24228,N_22922,N_22712);
xor U24229 (N_24229,N_23394,N_23388);
xnor U24230 (N_24230,N_22623,N_23130);
xor U24231 (N_24231,N_23060,N_23452);
nand U24232 (N_24232,N_23551,N_22976);
nand U24233 (N_24233,N_23066,N_22745);
or U24234 (N_24234,N_22865,N_23608);
nor U24235 (N_24235,N_23002,N_23223);
and U24236 (N_24236,N_22818,N_22557);
xor U24237 (N_24237,N_23022,N_22912);
and U24238 (N_24238,N_22737,N_22542);
and U24239 (N_24239,N_22516,N_23627);
nor U24240 (N_24240,N_23154,N_22589);
nor U24241 (N_24241,N_23454,N_23358);
and U24242 (N_24242,N_23519,N_22526);
and U24243 (N_24243,N_23436,N_22540);
or U24244 (N_24244,N_22654,N_23327);
or U24245 (N_24245,N_22905,N_23286);
nand U24246 (N_24246,N_22871,N_22957);
xor U24247 (N_24247,N_22673,N_23483);
nor U24248 (N_24248,N_23128,N_23720);
or U24249 (N_24249,N_23209,N_22633);
and U24250 (N_24250,N_23425,N_22558);
and U24251 (N_24251,N_22864,N_23391);
nor U24252 (N_24252,N_22971,N_23378);
and U24253 (N_24253,N_23099,N_22617);
xor U24254 (N_24254,N_23717,N_22625);
or U24255 (N_24255,N_23129,N_23258);
nor U24256 (N_24256,N_22645,N_22658);
nor U24257 (N_24257,N_23252,N_23442);
or U24258 (N_24258,N_23524,N_22637);
nor U24259 (N_24259,N_22923,N_23561);
nor U24260 (N_24260,N_22918,N_23598);
nand U24261 (N_24261,N_23635,N_22751);
and U24262 (N_24262,N_23644,N_23705);
and U24263 (N_24263,N_23016,N_23647);
and U24264 (N_24264,N_22711,N_23151);
and U24265 (N_24265,N_22850,N_22550);
or U24266 (N_24266,N_23297,N_23637);
nand U24267 (N_24267,N_22769,N_23035);
xor U24268 (N_24268,N_23119,N_23554);
and U24269 (N_24269,N_22764,N_22644);
and U24270 (N_24270,N_23074,N_23237);
and U24271 (N_24271,N_23379,N_23150);
nand U24272 (N_24272,N_23072,N_23049);
nand U24273 (N_24273,N_23226,N_22600);
xor U24274 (N_24274,N_22609,N_23350);
or U24275 (N_24275,N_23365,N_23731);
nand U24276 (N_24276,N_22545,N_23373);
xnor U24277 (N_24277,N_22533,N_23219);
or U24278 (N_24278,N_23271,N_22504);
nand U24279 (N_24279,N_22758,N_22544);
xor U24280 (N_24280,N_23249,N_23432);
nor U24281 (N_24281,N_23044,N_22506);
nand U24282 (N_24282,N_23645,N_23473);
nand U24283 (N_24283,N_23007,N_23349);
nor U24284 (N_24284,N_22733,N_23038);
nor U24285 (N_24285,N_23439,N_22709);
nor U24286 (N_24286,N_22670,N_23746);
and U24287 (N_24287,N_22537,N_23477);
nor U24288 (N_24288,N_23498,N_23489);
nand U24289 (N_24289,N_23116,N_23212);
nand U24290 (N_24290,N_23316,N_23274);
xnor U24291 (N_24291,N_22910,N_22815);
nor U24292 (N_24292,N_23449,N_23694);
xnor U24293 (N_24293,N_23208,N_23611);
nor U24294 (N_24294,N_23259,N_23553);
nor U24295 (N_24295,N_23484,N_23304);
and U24296 (N_24296,N_23323,N_23124);
nor U24297 (N_24297,N_22748,N_22731);
nor U24298 (N_24298,N_22967,N_23493);
nor U24299 (N_24299,N_23544,N_23294);
nand U24300 (N_24300,N_23342,N_23169);
and U24301 (N_24301,N_23476,N_23290);
nand U24302 (N_24302,N_23239,N_23036);
or U24303 (N_24303,N_23560,N_22571);
and U24304 (N_24304,N_23054,N_23094);
nor U24305 (N_24305,N_23485,N_22744);
xnor U24306 (N_24306,N_22853,N_23024);
nor U24307 (N_24307,N_23361,N_23475);
nand U24308 (N_24308,N_23302,N_22730);
and U24309 (N_24309,N_23709,N_23068);
nor U24310 (N_24310,N_23266,N_23445);
or U24311 (N_24311,N_23042,N_23275);
or U24312 (N_24312,N_23086,N_22718);
and U24313 (N_24313,N_22638,N_22857);
nor U24314 (N_24314,N_22725,N_23520);
nor U24315 (N_24315,N_23134,N_22765);
nand U24316 (N_24316,N_23276,N_22743);
nor U24317 (N_24317,N_23171,N_22771);
and U24318 (N_24318,N_23175,N_23688);
or U24319 (N_24319,N_22761,N_23584);
and U24320 (N_24320,N_22675,N_23733);
or U24321 (N_24321,N_23336,N_23657);
xnor U24322 (N_24322,N_22975,N_23410);
nor U24323 (N_24323,N_22972,N_22757);
or U24324 (N_24324,N_23366,N_23744);
nor U24325 (N_24325,N_22643,N_22992);
and U24326 (N_24326,N_22878,N_22795);
and U24327 (N_24327,N_23345,N_22903);
nand U24328 (N_24328,N_23181,N_23064);
or U24329 (N_24329,N_22722,N_23179);
xor U24330 (N_24330,N_22576,N_23491);
nand U24331 (N_24331,N_22794,N_23126);
nor U24332 (N_24332,N_23385,N_22606);
and U24333 (N_24333,N_23742,N_22893);
or U24334 (N_24334,N_23565,N_23149);
nand U24335 (N_24335,N_22667,N_23217);
xor U24336 (N_24336,N_23507,N_23586);
and U24337 (N_24337,N_22808,N_23446);
nand U24338 (N_24338,N_23168,N_22581);
and U24339 (N_24339,N_23707,N_22563);
or U24340 (N_24340,N_22983,N_22720);
xnor U24341 (N_24341,N_23207,N_22802);
nand U24342 (N_24342,N_22653,N_23716);
nor U24343 (N_24343,N_23506,N_22988);
or U24344 (N_24344,N_22848,N_22717);
nor U24345 (N_24345,N_22631,N_23486);
nor U24346 (N_24346,N_22584,N_22551);
nand U24347 (N_24347,N_22501,N_23141);
and U24348 (N_24348,N_23334,N_22869);
and U24349 (N_24349,N_22947,N_22824);
nand U24350 (N_24350,N_22919,N_23046);
nor U24351 (N_24351,N_23513,N_23238);
and U24352 (N_24352,N_22515,N_22610);
and U24353 (N_24353,N_22587,N_23585);
nand U24354 (N_24354,N_23575,N_23701);
and U24355 (N_24355,N_22591,N_23118);
nand U24356 (N_24356,N_23010,N_23353);
and U24357 (N_24357,N_23527,N_22772);
nand U24358 (N_24358,N_23721,N_23307);
xor U24359 (N_24359,N_23264,N_22602);
and U24360 (N_24360,N_22728,N_22968);
xnor U24361 (N_24361,N_23090,N_22573);
and U24362 (N_24362,N_23398,N_22907);
or U24363 (N_24363,N_23734,N_23229);
xor U24364 (N_24364,N_23123,N_23455);
nand U24365 (N_24365,N_22671,N_23041);
or U24366 (N_24366,N_23077,N_23107);
and U24367 (N_24367,N_23269,N_23161);
nand U24368 (N_24368,N_22680,N_23612);
or U24369 (N_24369,N_23083,N_22934);
nor U24370 (N_24370,N_22909,N_23370);
nand U24371 (N_24371,N_23674,N_23603);
nor U24372 (N_24372,N_23059,N_22939);
xor U24373 (N_24373,N_23663,N_22596);
xor U24374 (N_24374,N_22698,N_22868);
xor U24375 (N_24375,N_22795,N_23697);
nor U24376 (N_24376,N_22537,N_22744);
nor U24377 (N_24377,N_23404,N_23411);
nand U24378 (N_24378,N_22619,N_23402);
or U24379 (N_24379,N_23313,N_22758);
and U24380 (N_24380,N_22500,N_22724);
xnor U24381 (N_24381,N_22835,N_23510);
nor U24382 (N_24382,N_23119,N_23176);
or U24383 (N_24383,N_22551,N_22678);
or U24384 (N_24384,N_23184,N_23252);
or U24385 (N_24385,N_23560,N_23318);
or U24386 (N_24386,N_23436,N_23610);
xnor U24387 (N_24387,N_22831,N_23641);
or U24388 (N_24388,N_23584,N_23269);
nand U24389 (N_24389,N_23714,N_23666);
nand U24390 (N_24390,N_23234,N_22968);
xnor U24391 (N_24391,N_22715,N_22954);
xor U24392 (N_24392,N_22957,N_23634);
and U24393 (N_24393,N_23469,N_23452);
and U24394 (N_24394,N_23733,N_23588);
nand U24395 (N_24395,N_22907,N_22630);
or U24396 (N_24396,N_22912,N_23046);
nand U24397 (N_24397,N_23278,N_23532);
xnor U24398 (N_24398,N_22709,N_23364);
or U24399 (N_24399,N_23185,N_23097);
and U24400 (N_24400,N_22885,N_22816);
nor U24401 (N_24401,N_23364,N_23390);
xnor U24402 (N_24402,N_23612,N_22897);
or U24403 (N_24403,N_23290,N_22819);
nand U24404 (N_24404,N_22779,N_23161);
nand U24405 (N_24405,N_22671,N_23648);
nand U24406 (N_24406,N_22771,N_23116);
nor U24407 (N_24407,N_23308,N_22782);
nand U24408 (N_24408,N_23009,N_22748);
nand U24409 (N_24409,N_22870,N_23365);
or U24410 (N_24410,N_23241,N_23087);
nor U24411 (N_24411,N_23489,N_22784);
nand U24412 (N_24412,N_23276,N_23619);
xor U24413 (N_24413,N_23574,N_22647);
xor U24414 (N_24414,N_23236,N_22696);
or U24415 (N_24415,N_23458,N_23144);
or U24416 (N_24416,N_23131,N_23492);
nand U24417 (N_24417,N_23140,N_23644);
or U24418 (N_24418,N_23128,N_22855);
or U24419 (N_24419,N_23148,N_22534);
nor U24420 (N_24420,N_23359,N_22710);
xor U24421 (N_24421,N_23170,N_23332);
and U24422 (N_24422,N_23213,N_23662);
nor U24423 (N_24423,N_23336,N_23094);
xor U24424 (N_24424,N_23083,N_23049);
nor U24425 (N_24425,N_22781,N_23057);
nand U24426 (N_24426,N_23068,N_23396);
and U24427 (N_24427,N_23011,N_23517);
and U24428 (N_24428,N_23370,N_23593);
and U24429 (N_24429,N_22860,N_22751);
nor U24430 (N_24430,N_22567,N_23574);
nand U24431 (N_24431,N_23309,N_23213);
or U24432 (N_24432,N_23146,N_23107);
nand U24433 (N_24433,N_23677,N_23698);
and U24434 (N_24434,N_23683,N_22761);
and U24435 (N_24435,N_23711,N_22618);
and U24436 (N_24436,N_23288,N_23036);
xor U24437 (N_24437,N_23012,N_23446);
and U24438 (N_24438,N_23210,N_23000);
or U24439 (N_24439,N_22629,N_23055);
nor U24440 (N_24440,N_22592,N_22665);
xor U24441 (N_24441,N_23227,N_22656);
nand U24442 (N_24442,N_22586,N_22798);
nand U24443 (N_24443,N_22658,N_23161);
nor U24444 (N_24444,N_23683,N_22809);
nand U24445 (N_24445,N_22968,N_23468);
nor U24446 (N_24446,N_23228,N_23595);
nor U24447 (N_24447,N_22559,N_22742);
or U24448 (N_24448,N_22732,N_22754);
and U24449 (N_24449,N_22993,N_23672);
nand U24450 (N_24450,N_22556,N_23268);
and U24451 (N_24451,N_22913,N_23110);
nand U24452 (N_24452,N_22872,N_22803);
and U24453 (N_24453,N_23625,N_23408);
or U24454 (N_24454,N_23243,N_23733);
and U24455 (N_24455,N_23052,N_23334);
nor U24456 (N_24456,N_22680,N_22898);
nand U24457 (N_24457,N_23325,N_22744);
nor U24458 (N_24458,N_23321,N_22644);
nor U24459 (N_24459,N_22792,N_23423);
or U24460 (N_24460,N_22621,N_22940);
nor U24461 (N_24461,N_23438,N_23054);
xnor U24462 (N_24462,N_22545,N_22571);
nor U24463 (N_24463,N_23572,N_23494);
and U24464 (N_24464,N_23089,N_22582);
nor U24465 (N_24465,N_23285,N_23735);
nor U24466 (N_24466,N_22783,N_22704);
or U24467 (N_24467,N_23218,N_22574);
nand U24468 (N_24468,N_22539,N_23601);
xor U24469 (N_24469,N_22809,N_23000);
and U24470 (N_24470,N_23243,N_22810);
and U24471 (N_24471,N_22975,N_23481);
or U24472 (N_24472,N_23551,N_23608);
nor U24473 (N_24473,N_23508,N_22962);
xor U24474 (N_24474,N_23717,N_23656);
or U24475 (N_24475,N_22519,N_22547);
nor U24476 (N_24476,N_23687,N_23078);
nand U24477 (N_24477,N_22681,N_22510);
nor U24478 (N_24478,N_23404,N_23696);
nand U24479 (N_24479,N_22747,N_23317);
or U24480 (N_24480,N_23349,N_23280);
and U24481 (N_24481,N_22852,N_23644);
and U24482 (N_24482,N_22913,N_23722);
nand U24483 (N_24483,N_23112,N_23082);
or U24484 (N_24484,N_23152,N_23423);
nand U24485 (N_24485,N_23522,N_23552);
xnor U24486 (N_24486,N_23214,N_23475);
xor U24487 (N_24487,N_23731,N_23268);
nand U24488 (N_24488,N_22932,N_22825);
nand U24489 (N_24489,N_22674,N_23609);
and U24490 (N_24490,N_23157,N_22719);
xnor U24491 (N_24491,N_22878,N_23485);
and U24492 (N_24492,N_22878,N_23529);
or U24493 (N_24493,N_23272,N_23208);
nand U24494 (N_24494,N_23195,N_23592);
xnor U24495 (N_24495,N_22939,N_22518);
and U24496 (N_24496,N_23539,N_23111);
nor U24497 (N_24497,N_22992,N_23168);
nor U24498 (N_24498,N_22928,N_22840);
or U24499 (N_24499,N_23543,N_22771);
xor U24500 (N_24500,N_22517,N_23628);
nand U24501 (N_24501,N_23485,N_23368);
nand U24502 (N_24502,N_22660,N_22683);
and U24503 (N_24503,N_23001,N_22582);
and U24504 (N_24504,N_23475,N_22759);
or U24505 (N_24505,N_22964,N_22794);
xnor U24506 (N_24506,N_22641,N_23261);
and U24507 (N_24507,N_22745,N_22678);
nor U24508 (N_24508,N_23667,N_23016);
xnor U24509 (N_24509,N_23593,N_22827);
nand U24510 (N_24510,N_23574,N_23582);
xnor U24511 (N_24511,N_23487,N_23606);
nand U24512 (N_24512,N_23590,N_23322);
xor U24513 (N_24513,N_23250,N_22637);
nand U24514 (N_24514,N_23292,N_23088);
xor U24515 (N_24515,N_22786,N_23214);
and U24516 (N_24516,N_22791,N_23054);
and U24517 (N_24517,N_23408,N_23704);
and U24518 (N_24518,N_22778,N_22723);
xnor U24519 (N_24519,N_23447,N_22505);
and U24520 (N_24520,N_23572,N_23593);
xnor U24521 (N_24521,N_23313,N_23495);
nor U24522 (N_24522,N_23028,N_23424);
nand U24523 (N_24523,N_22687,N_23288);
xor U24524 (N_24524,N_23505,N_23510);
nand U24525 (N_24525,N_22551,N_22992);
nand U24526 (N_24526,N_23364,N_23016);
xnor U24527 (N_24527,N_23303,N_22885);
xnor U24528 (N_24528,N_23666,N_22686);
nand U24529 (N_24529,N_22765,N_22968);
nand U24530 (N_24530,N_22543,N_22730);
nor U24531 (N_24531,N_23378,N_23704);
xor U24532 (N_24532,N_22619,N_23739);
nand U24533 (N_24533,N_22596,N_23418);
xnor U24534 (N_24534,N_22979,N_22927);
or U24535 (N_24535,N_23128,N_23424);
and U24536 (N_24536,N_23054,N_22631);
nor U24537 (N_24537,N_23115,N_23510);
xor U24538 (N_24538,N_22586,N_22660);
xor U24539 (N_24539,N_23047,N_22548);
nand U24540 (N_24540,N_23073,N_22652);
nor U24541 (N_24541,N_22912,N_23179);
and U24542 (N_24542,N_22936,N_23623);
and U24543 (N_24543,N_23464,N_22795);
or U24544 (N_24544,N_23207,N_22722);
or U24545 (N_24545,N_23539,N_22866);
or U24546 (N_24546,N_23655,N_23630);
and U24547 (N_24547,N_22502,N_23550);
or U24548 (N_24548,N_22686,N_23146);
and U24549 (N_24549,N_23595,N_23548);
nor U24550 (N_24550,N_23669,N_22796);
xnor U24551 (N_24551,N_22665,N_22548);
xor U24552 (N_24552,N_22686,N_23493);
xor U24553 (N_24553,N_23443,N_23210);
and U24554 (N_24554,N_23551,N_23705);
nor U24555 (N_24555,N_23413,N_23117);
nor U24556 (N_24556,N_22662,N_23051);
nand U24557 (N_24557,N_23167,N_22950);
nand U24558 (N_24558,N_23175,N_22872);
nor U24559 (N_24559,N_22844,N_23360);
nor U24560 (N_24560,N_22650,N_23267);
nor U24561 (N_24561,N_22865,N_22666);
and U24562 (N_24562,N_23575,N_23622);
xor U24563 (N_24563,N_23442,N_23448);
nor U24564 (N_24564,N_22784,N_22755);
and U24565 (N_24565,N_22886,N_23446);
nand U24566 (N_24566,N_23466,N_23041);
nand U24567 (N_24567,N_22805,N_22884);
nor U24568 (N_24568,N_23200,N_22853);
or U24569 (N_24569,N_22854,N_22781);
and U24570 (N_24570,N_23556,N_23497);
nand U24571 (N_24571,N_23583,N_22840);
nor U24572 (N_24572,N_23426,N_23252);
or U24573 (N_24573,N_23482,N_23566);
xnor U24574 (N_24574,N_22869,N_22509);
or U24575 (N_24575,N_22670,N_23512);
nand U24576 (N_24576,N_22544,N_23230);
and U24577 (N_24577,N_22756,N_23472);
xor U24578 (N_24578,N_23699,N_23454);
and U24579 (N_24579,N_22736,N_23204);
or U24580 (N_24580,N_23578,N_23420);
or U24581 (N_24581,N_23145,N_22650);
or U24582 (N_24582,N_23673,N_23210);
nor U24583 (N_24583,N_23052,N_23701);
or U24584 (N_24584,N_23596,N_23261);
and U24585 (N_24585,N_23484,N_22622);
nand U24586 (N_24586,N_22688,N_22906);
nor U24587 (N_24587,N_22660,N_22771);
and U24588 (N_24588,N_23207,N_22597);
and U24589 (N_24589,N_23441,N_23612);
or U24590 (N_24590,N_22910,N_22583);
or U24591 (N_24591,N_22952,N_23411);
or U24592 (N_24592,N_23637,N_22588);
nor U24593 (N_24593,N_23006,N_22900);
xor U24594 (N_24594,N_22506,N_23149);
and U24595 (N_24595,N_23327,N_22868);
or U24596 (N_24596,N_23552,N_22576);
nor U24597 (N_24597,N_23169,N_23657);
or U24598 (N_24598,N_23655,N_22913);
and U24599 (N_24599,N_23224,N_22761);
nor U24600 (N_24600,N_23034,N_23410);
and U24601 (N_24601,N_23450,N_23008);
nand U24602 (N_24602,N_22935,N_22927);
xor U24603 (N_24603,N_22617,N_23705);
nand U24604 (N_24604,N_23299,N_22908);
or U24605 (N_24605,N_22529,N_23575);
nor U24606 (N_24606,N_22937,N_23199);
nand U24607 (N_24607,N_23257,N_23350);
xnor U24608 (N_24608,N_23703,N_22723);
nand U24609 (N_24609,N_22866,N_22500);
or U24610 (N_24610,N_22706,N_22513);
and U24611 (N_24611,N_23303,N_22570);
nand U24612 (N_24612,N_22759,N_23338);
or U24613 (N_24613,N_23520,N_23054);
nor U24614 (N_24614,N_23737,N_23327);
or U24615 (N_24615,N_23497,N_23063);
or U24616 (N_24616,N_22539,N_23651);
or U24617 (N_24617,N_23366,N_23469);
xnor U24618 (N_24618,N_23182,N_22754);
xnor U24619 (N_24619,N_23419,N_22617);
and U24620 (N_24620,N_22928,N_23310);
xnor U24621 (N_24621,N_23572,N_22792);
nor U24622 (N_24622,N_23628,N_23525);
nor U24623 (N_24623,N_22768,N_22992);
and U24624 (N_24624,N_22504,N_23301);
and U24625 (N_24625,N_22523,N_22693);
nor U24626 (N_24626,N_22544,N_23643);
nand U24627 (N_24627,N_23469,N_23505);
or U24628 (N_24628,N_22892,N_22754);
nor U24629 (N_24629,N_22818,N_23729);
nand U24630 (N_24630,N_23738,N_23385);
nand U24631 (N_24631,N_22702,N_23291);
and U24632 (N_24632,N_23592,N_22961);
and U24633 (N_24633,N_22537,N_23707);
and U24634 (N_24634,N_23118,N_22688);
and U24635 (N_24635,N_22815,N_23506);
nor U24636 (N_24636,N_23069,N_23480);
nor U24637 (N_24637,N_22957,N_22654);
and U24638 (N_24638,N_23688,N_22849);
and U24639 (N_24639,N_23580,N_22908);
xor U24640 (N_24640,N_23391,N_23498);
or U24641 (N_24641,N_23649,N_23701);
and U24642 (N_24642,N_23058,N_22928);
or U24643 (N_24643,N_23270,N_23336);
xor U24644 (N_24644,N_23440,N_22513);
and U24645 (N_24645,N_23692,N_22515);
and U24646 (N_24646,N_23280,N_23564);
nor U24647 (N_24647,N_23188,N_23284);
and U24648 (N_24648,N_23223,N_23694);
xnor U24649 (N_24649,N_22857,N_23624);
nor U24650 (N_24650,N_22653,N_23692);
and U24651 (N_24651,N_23116,N_23479);
xor U24652 (N_24652,N_22875,N_23427);
or U24653 (N_24653,N_23720,N_23354);
nand U24654 (N_24654,N_23158,N_22734);
and U24655 (N_24655,N_22841,N_23484);
nand U24656 (N_24656,N_23246,N_23018);
or U24657 (N_24657,N_23451,N_22841);
and U24658 (N_24658,N_22636,N_22731);
and U24659 (N_24659,N_23541,N_23481);
or U24660 (N_24660,N_23294,N_22681);
nand U24661 (N_24661,N_22954,N_22822);
or U24662 (N_24662,N_23543,N_22741);
or U24663 (N_24663,N_23490,N_23555);
nand U24664 (N_24664,N_23023,N_22858);
xor U24665 (N_24665,N_22580,N_23582);
nor U24666 (N_24666,N_23457,N_23095);
xnor U24667 (N_24667,N_23495,N_22903);
or U24668 (N_24668,N_23274,N_22949);
nor U24669 (N_24669,N_23242,N_23093);
nand U24670 (N_24670,N_22829,N_23416);
or U24671 (N_24671,N_22801,N_23365);
nand U24672 (N_24672,N_23593,N_22646);
and U24673 (N_24673,N_23369,N_23741);
and U24674 (N_24674,N_22647,N_23567);
nor U24675 (N_24675,N_22609,N_23108);
and U24676 (N_24676,N_23238,N_23598);
nand U24677 (N_24677,N_22716,N_23171);
xor U24678 (N_24678,N_22632,N_23608);
or U24679 (N_24679,N_22593,N_22748);
and U24680 (N_24680,N_22839,N_23468);
and U24681 (N_24681,N_22671,N_22798);
xnor U24682 (N_24682,N_22851,N_22970);
nor U24683 (N_24683,N_23668,N_23199);
xnor U24684 (N_24684,N_23431,N_22651);
or U24685 (N_24685,N_23199,N_23747);
nor U24686 (N_24686,N_23562,N_23166);
or U24687 (N_24687,N_23194,N_22618);
and U24688 (N_24688,N_22845,N_23567);
or U24689 (N_24689,N_22888,N_23412);
nor U24690 (N_24690,N_22696,N_22718);
or U24691 (N_24691,N_22970,N_23727);
and U24692 (N_24692,N_22657,N_23338);
nor U24693 (N_24693,N_22501,N_23716);
nor U24694 (N_24694,N_23726,N_23098);
nor U24695 (N_24695,N_23551,N_22891);
nand U24696 (N_24696,N_23239,N_23157);
and U24697 (N_24697,N_23372,N_23182);
nor U24698 (N_24698,N_23696,N_22886);
nand U24699 (N_24699,N_22598,N_23220);
nor U24700 (N_24700,N_22883,N_23684);
nand U24701 (N_24701,N_22607,N_23300);
nor U24702 (N_24702,N_23363,N_22939);
and U24703 (N_24703,N_22700,N_22948);
and U24704 (N_24704,N_22959,N_22645);
and U24705 (N_24705,N_23675,N_23707);
and U24706 (N_24706,N_23669,N_23562);
or U24707 (N_24707,N_23557,N_23180);
and U24708 (N_24708,N_23028,N_22689);
and U24709 (N_24709,N_23609,N_22756);
nand U24710 (N_24710,N_22865,N_23300);
nand U24711 (N_24711,N_22762,N_22912);
nor U24712 (N_24712,N_23156,N_23332);
xnor U24713 (N_24713,N_22920,N_23543);
xnor U24714 (N_24714,N_22544,N_23066);
nand U24715 (N_24715,N_23124,N_22877);
nand U24716 (N_24716,N_22604,N_23594);
xnor U24717 (N_24717,N_23674,N_22930);
nand U24718 (N_24718,N_23659,N_23579);
nand U24719 (N_24719,N_23408,N_23295);
nor U24720 (N_24720,N_22644,N_22513);
nor U24721 (N_24721,N_22720,N_23529);
nor U24722 (N_24722,N_22667,N_23169);
or U24723 (N_24723,N_23104,N_23734);
and U24724 (N_24724,N_23328,N_22783);
or U24725 (N_24725,N_23706,N_23525);
or U24726 (N_24726,N_23709,N_23126);
or U24727 (N_24727,N_23486,N_23389);
or U24728 (N_24728,N_22836,N_23172);
and U24729 (N_24729,N_22710,N_23024);
or U24730 (N_24730,N_23341,N_23194);
or U24731 (N_24731,N_23614,N_23148);
nor U24732 (N_24732,N_22973,N_23443);
xor U24733 (N_24733,N_23366,N_23631);
nand U24734 (N_24734,N_23073,N_22587);
nand U24735 (N_24735,N_23303,N_23735);
nor U24736 (N_24736,N_23309,N_23340);
and U24737 (N_24737,N_23350,N_23185);
nand U24738 (N_24738,N_23430,N_23231);
or U24739 (N_24739,N_22572,N_22515);
nand U24740 (N_24740,N_23422,N_23436);
nor U24741 (N_24741,N_22980,N_22567);
or U24742 (N_24742,N_23208,N_23446);
and U24743 (N_24743,N_23396,N_22888);
and U24744 (N_24744,N_22610,N_22589);
nand U24745 (N_24745,N_23490,N_22766);
and U24746 (N_24746,N_22536,N_23711);
nor U24747 (N_24747,N_23317,N_23390);
and U24748 (N_24748,N_22617,N_23449);
xnor U24749 (N_24749,N_22795,N_23552);
and U24750 (N_24750,N_23603,N_23524);
and U24751 (N_24751,N_23414,N_22691);
or U24752 (N_24752,N_23027,N_23476);
and U24753 (N_24753,N_23747,N_23602);
or U24754 (N_24754,N_23455,N_23026);
xor U24755 (N_24755,N_23310,N_22748);
nand U24756 (N_24756,N_22595,N_22614);
nand U24757 (N_24757,N_23155,N_22956);
and U24758 (N_24758,N_22523,N_22733);
nor U24759 (N_24759,N_23086,N_23604);
or U24760 (N_24760,N_22859,N_23418);
nor U24761 (N_24761,N_23249,N_23189);
or U24762 (N_24762,N_23218,N_22779);
nand U24763 (N_24763,N_23364,N_23310);
or U24764 (N_24764,N_23649,N_23194);
nand U24765 (N_24765,N_22768,N_23135);
nor U24766 (N_24766,N_23156,N_22567);
nor U24767 (N_24767,N_23367,N_23511);
and U24768 (N_24768,N_23228,N_22882);
or U24769 (N_24769,N_22765,N_22744);
nand U24770 (N_24770,N_23181,N_23464);
xnor U24771 (N_24771,N_23013,N_22916);
nor U24772 (N_24772,N_22950,N_22942);
nor U24773 (N_24773,N_22702,N_23597);
nor U24774 (N_24774,N_22575,N_23435);
and U24775 (N_24775,N_23716,N_23558);
nand U24776 (N_24776,N_22505,N_23587);
nor U24777 (N_24777,N_22997,N_23501);
and U24778 (N_24778,N_23477,N_22742);
xnor U24779 (N_24779,N_23502,N_22953);
nand U24780 (N_24780,N_23671,N_22512);
or U24781 (N_24781,N_22529,N_23719);
nand U24782 (N_24782,N_22830,N_23507);
or U24783 (N_24783,N_22954,N_22607);
nand U24784 (N_24784,N_23495,N_23326);
or U24785 (N_24785,N_23685,N_23074);
or U24786 (N_24786,N_23589,N_23069);
nor U24787 (N_24787,N_22664,N_23690);
or U24788 (N_24788,N_22985,N_22840);
xnor U24789 (N_24789,N_22756,N_23567);
and U24790 (N_24790,N_23317,N_23460);
and U24791 (N_24791,N_23288,N_22756);
and U24792 (N_24792,N_23511,N_22558);
xnor U24793 (N_24793,N_23097,N_22866);
nand U24794 (N_24794,N_23635,N_22526);
xnor U24795 (N_24795,N_22723,N_22806);
nand U24796 (N_24796,N_22625,N_22936);
nand U24797 (N_24797,N_23568,N_23249);
and U24798 (N_24798,N_23543,N_23659);
and U24799 (N_24799,N_23375,N_23133);
or U24800 (N_24800,N_22719,N_23683);
xnor U24801 (N_24801,N_23127,N_22638);
or U24802 (N_24802,N_23530,N_23142);
nand U24803 (N_24803,N_22797,N_22668);
nand U24804 (N_24804,N_23257,N_23537);
or U24805 (N_24805,N_23508,N_23462);
and U24806 (N_24806,N_22598,N_23140);
xnor U24807 (N_24807,N_22707,N_23046);
or U24808 (N_24808,N_23747,N_22869);
and U24809 (N_24809,N_23149,N_22719);
and U24810 (N_24810,N_22829,N_23088);
nand U24811 (N_24811,N_23644,N_22901);
and U24812 (N_24812,N_22722,N_23268);
nor U24813 (N_24813,N_23119,N_22910);
nand U24814 (N_24814,N_23211,N_23586);
and U24815 (N_24815,N_23646,N_23585);
nand U24816 (N_24816,N_23198,N_22683);
or U24817 (N_24817,N_23428,N_23141);
or U24818 (N_24818,N_23110,N_22612);
or U24819 (N_24819,N_22514,N_22779);
xor U24820 (N_24820,N_23226,N_23743);
or U24821 (N_24821,N_23291,N_23121);
nor U24822 (N_24822,N_23588,N_22852);
nand U24823 (N_24823,N_23471,N_23528);
nand U24824 (N_24824,N_23411,N_23498);
nand U24825 (N_24825,N_23099,N_23103);
nor U24826 (N_24826,N_23581,N_22889);
nor U24827 (N_24827,N_22910,N_23527);
nand U24828 (N_24828,N_23464,N_23008);
or U24829 (N_24829,N_22721,N_23271);
nor U24830 (N_24830,N_23102,N_23668);
nand U24831 (N_24831,N_23588,N_23316);
nand U24832 (N_24832,N_23091,N_23426);
and U24833 (N_24833,N_22712,N_22716);
nand U24834 (N_24834,N_23165,N_23249);
nor U24835 (N_24835,N_22700,N_23532);
nor U24836 (N_24836,N_23164,N_22858);
and U24837 (N_24837,N_22625,N_22779);
nor U24838 (N_24838,N_23642,N_23737);
nand U24839 (N_24839,N_22643,N_22817);
nand U24840 (N_24840,N_23692,N_23106);
nor U24841 (N_24841,N_23116,N_23567);
and U24842 (N_24842,N_22593,N_23580);
nand U24843 (N_24843,N_22994,N_22611);
and U24844 (N_24844,N_23373,N_22979);
nand U24845 (N_24845,N_22839,N_22909);
xor U24846 (N_24846,N_23542,N_22643);
and U24847 (N_24847,N_23089,N_23445);
nand U24848 (N_24848,N_23044,N_23629);
xor U24849 (N_24849,N_23133,N_23289);
and U24850 (N_24850,N_22992,N_22912);
and U24851 (N_24851,N_23076,N_23150);
and U24852 (N_24852,N_23617,N_22595);
nor U24853 (N_24853,N_22886,N_22572);
xnor U24854 (N_24854,N_23175,N_23365);
or U24855 (N_24855,N_23329,N_23102);
nor U24856 (N_24856,N_22643,N_23631);
or U24857 (N_24857,N_22727,N_23214);
and U24858 (N_24858,N_23749,N_23440);
xnor U24859 (N_24859,N_22921,N_22866);
nand U24860 (N_24860,N_22599,N_22716);
nor U24861 (N_24861,N_23387,N_23633);
nand U24862 (N_24862,N_23135,N_23339);
nor U24863 (N_24863,N_23300,N_23679);
nor U24864 (N_24864,N_22941,N_22614);
and U24865 (N_24865,N_22898,N_22796);
and U24866 (N_24866,N_23163,N_22716);
nand U24867 (N_24867,N_22998,N_23727);
nor U24868 (N_24868,N_23433,N_22933);
nand U24869 (N_24869,N_23037,N_23130);
and U24870 (N_24870,N_22576,N_22960);
nor U24871 (N_24871,N_23098,N_23434);
and U24872 (N_24872,N_23115,N_23022);
xnor U24873 (N_24873,N_22578,N_23135);
or U24874 (N_24874,N_22914,N_23318);
nand U24875 (N_24875,N_22716,N_23336);
and U24876 (N_24876,N_22640,N_22555);
nand U24877 (N_24877,N_22527,N_23593);
nor U24878 (N_24878,N_22675,N_23705);
and U24879 (N_24879,N_22861,N_23089);
or U24880 (N_24880,N_23077,N_23402);
and U24881 (N_24881,N_22573,N_22812);
nand U24882 (N_24882,N_22969,N_22776);
or U24883 (N_24883,N_23578,N_23163);
and U24884 (N_24884,N_23210,N_22507);
nor U24885 (N_24885,N_23206,N_23006);
nor U24886 (N_24886,N_23024,N_23635);
and U24887 (N_24887,N_23028,N_23665);
or U24888 (N_24888,N_23623,N_23626);
nor U24889 (N_24889,N_23266,N_23147);
nor U24890 (N_24890,N_23063,N_23387);
nor U24891 (N_24891,N_22967,N_23519);
nand U24892 (N_24892,N_23473,N_23365);
nor U24893 (N_24893,N_22754,N_22715);
or U24894 (N_24894,N_23647,N_22576);
and U24895 (N_24895,N_22816,N_23487);
nor U24896 (N_24896,N_23212,N_22648);
or U24897 (N_24897,N_22997,N_23452);
nand U24898 (N_24898,N_23320,N_23188);
nor U24899 (N_24899,N_22520,N_22768);
and U24900 (N_24900,N_22842,N_22807);
or U24901 (N_24901,N_23065,N_22587);
xnor U24902 (N_24902,N_22621,N_22988);
nor U24903 (N_24903,N_22985,N_23458);
nand U24904 (N_24904,N_23575,N_22576);
nand U24905 (N_24905,N_23537,N_23171);
nor U24906 (N_24906,N_22591,N_22720);
xor U24907 (N_24907,N_23645,N_23050);
and U24908 (N_24908,N_22686,N_22530);
nor U24909 (N_24909,N_22756,N_23090);
or U24910 (N_24910,N_23117,N_23116);
xor U24911 (N_24911,N_23504,N_23234);
nand U24912 (N_24912,N_23184,N_23063);
nand U24913 (N_24913,N_23046,N_23126);
nor U24914 (N_24914,N_22571,N_22792);
nand U24915 (N_24915,N_22724,N_23192);
nor U24916 (N_24916,N_23594,N_22528);
nand U24917 (N_24917,N_23487,N_23152);
nand U24918 (N_24918,N_22580,N_23585);
nor U24919 (N_24919,N_23238,N_22821);
nor U24920 (N_24920,N_22866,N_23141);
nor U24921 (N_24921,N_23468,N_22746);
and U24922 (N_24922,N_22523,N_22647);
nand U24923 (N_24923,N_22864,N_23726);
nand U24924 (N_24924,N_23126,N_22876);
nor U24925 (N_24925,N_23240,N_22912);
nand U24926 (N_24926,N_23453,N_23685);
nand U24927 (N_24927,N_22938,N_23456);
nor U24928 (N_24928,N_22515,N_22571);
and U24929 (N_24929,N_23403,N_23286);
nand U24930 (N_24930,N_22712,N_22928);
xnor U24931 (N_24931,N_23591,N_22540);
and U24932 (N_24932,N_23305,N_23438);
or U24933 (N_24933,N_23628,N_22801);
or U24934 (N_24934,N_23329,N_23504);
xnor U24935 (N_24935,N_22685,N_23002);
nand U24936 (N_24936,N_23220,N_23561);
and U24937 (N_24937,N_23149,N_22633);
xnor U24938 (N_24938,N_22717,N_22574);
xnor U24939 (N_24939,N_22944,N_22514);
nor U24940 (N_24940,N_23542,N_22546);
nand U24941 (N_24941,N_23373,N_23379);
or U24942 (N_24942,N_23333,N_22958);
and U24943 (N_24943,N_23204,N_22819);
nand U24944 (N_24944,N_23485,N_22756);
xor U24945 (N_24945,N_23255,N_23157);
nor U24946 (N_24946,N_22986,N_22944);
and U24947 (N_24947,N_23727,N_23552);
or U24948 (N_24948,N_23037,N_23739);
nand U24949 (N_24949,N_23587,N_22739);
xnor U24950 (N_24950,N_23507,N_22795);
xnor U24951 (N_24951,N_23224,N_23272);
and U24952 (N_24952,N_23730,N_22826);
and U24953 (N_24953,N_23113,N_23470);
xor U24954 (N_24954,N_22783,N_23413);
or U24955 (N_24955,N_22801,N_22683);
nor U24956 (N_24956,N_23078,N_23172);
xnor U24957 (N_24957,N_23167,N_22906);
and U24958 (N_24958,N_22985,N_23045);
or U24959 (N_24959,N_23526,N_23206);
and U24960 (N_24960,N_23719,N_22791);
nor U24961 (N_24961,N_22728,N_22737);
nand U24962 (N_24962,N_23564,N_23008);
nor U24963 (N_24963,N_22506,N_23230);
xnor U24964 (N_24964,N_23355,N_23087);
xor U24965 (N_24965,N_22735,N_22587);
nand U24966 (N_24966,N_22654,N_22930);
and U24967 (N_24967,N_23463,N_22854);
nand U24968 (N_24968,N_23415,N_23619);
or U24969 (N_24969,N_22727,N_23721);
and U24970 (N_24970,N_23527,N_23323);
nand U24971 (N_24971,N_23423,N_22635);
nand U24972 (N_24972,N_23198,N_22889);
xor U24973 (N_24973,N_22915,N_22781);
nor U24974 (N_24974,N_22955,N_22500);
xor U24975 (N_24975,N_23570,N_23531);
or U24976 (N_24976,N_23290,N_22866);
or U24977 (N_24977,N_23423,N_23061);
xnor U24978 (N_24978,N_23277,N_23502);
xor U24979 (N_24979,N_23456,N_22698);
or U24980 (N_24980,N_22555,N_23269);
xor U24981 (N_24981,N_23737,N_22603);
and U24982 (N_24982,N_23622,N_23081);
nor U24983 (N_24983,N_22587,N_22780);
or U24984 (N_24984,N_23532,N_22714);
or U24985 (N_24985,N_22930,N_23134);
or U24986 (N_24986,N_23212,N_23079);
or U24987 (N_24987,N_23665,N_23253);
or U24988 (N_24988,N_22766,N_22633);
nand U24989 (N_24989,N_23146,N_23603);
and U24990 (N_24990,N_22562,N_23107);
nand U24991 (N_24991,N_22932,N_23166);
and U24992 (N_24992,N_23698,N_23077);
xor U24993 (N_24993,N_22621,N_22636);
nand U24994 (N_24994,N_23273,N_23429);
xnor U24995 (N_24995,N_23517,N_23655);
nor U24996 (N_24996,N_23539,N_22566);
or U24997 (N_24997,N_23294,N_23096);
xnor U24998 (N_24998,N_23091,N_22961);
or U24999 (N_24999,N_23176,N_22669);
or UO_0 (O_0,N_24208,N_24963);
xnor UO_1 (O_1,N_24368,N_24906);
xor UO_2 (O_2,N_24572,N_24456);
and UO_3 (O_3,N_23996,N_23957);
nand UO_4 (O_4,N_24950,N_24130);
and UO_5 (O_5,N_24201,N_24378);
xnor UO_6 (O_6,N_24432,N_23910);
nand UO_7 (O_7,N_24257,N_24487);
nor UO_8 (O_8,N_24956,N_24347);
or UO_9 (O_9,N_24069,N_24611);
or UO_10 (O_10,N_24073,N_24612);
nand UO_11 (O_11,N_24031,N_24655);
and UO_12 (O_12,N_24892,N_24515);
or UO_13 (O_13,N_23900,N_23809);
nand UO_14 (O_14,N_24014,N_24436);
nand UO_15 (O_15,N_24348,N_23822);
nand UO_16 (O_16,N_23935,N_24163);
xnor UO_17 (O_17,N_23816,N_24986);
xnor UO_18 (O_18,N_24443,N_24643);
and UO_19 (O_19,N_24565,N_24067);
nand UO_20 (O_20,N_24949,N_24769);
or UO_21 (O_21,N_24918,N_23912);
or UO_22 (O_22,N_24004,N_23986);
nand UO_23 (O_23,N_24016,N_24283);
and UO_24 (O_24,N_23922,N_24756);
nand UO_25 (O_25,N_24260,N_24496);
or UO_26 (O_26,N_24092,N_24736);
or UO_27 (O_27,N_24838,N_24581);
or UO_28 (O_28,N_24191,N_24000);
nand UO_29 (O_29,N_24763,N_24328);
and UO_30 (O_30,N_24250,N_24122);
xnor UO_31 (O_31,N_24789,N_24154);
nor UO_32 (O_32,N_23752,N_24697);
nor UO_33 (O_33,N_24526,N_23997);
nand UO_34 (O_34,N_23792,N_24959);
xor UO_35 (O_35,N_24110,N_24290);
and UO_36 (O_36,N_24943,N_24404);
nor UO_37 (O_37,N_24678,N_23949);
xor UO_38 (O_38,N_24089,N_24304);
and UO_39 (O_39,N_24844,N_23806);
and UO_40 (O_40,N_24808,N_24142);
xnor UO_41 (O_41,N_24141,N_24822);
or UO_42 (O_42,N_24783,N_24277);
nor UO_43 (O_43,N_23911,N_24753);
and UO_44 (O_44,N_24026,N_24811);
xnor UO_45 (O_45,N_24477,N_24075);
nand UO_46 (O_46,N_24781,N_24005);
nand UO_47 (O_47,N_24019,N_24746);
xnor UO_48 (O_48,N_24398,N_24412);
nor UO_49 (O_49,N_24859,N_24561);
or UO_50 (O_50,N_24941,N_24936);
nand UO_51 (O_51,N_23772,N_23812);
nor UO_52 (O_52,N_24103,N_24536);
or UO_53 (O_53,N_24274,N_24706);
nor UO_54 (O_54,N_24704,N_24939);
or UO_55 (O_55,N_23895,N_24902);
or UO_56 (O_56,N_24206,N_24869);
or UO_57 (O_57,N_24938,N_24500);
xnor UO_58 (O_58,N_23976,N_24241);
nand UO_59 (O_59,N_24270,N_24013);
xnor UO_60 (O_60,N_24900,N_23914);
nor UO_61 (O_61,N_24463,N_23800);
nand UO_62 (O_62,N_23953,N_24948);
and UO_63 (O_63,N_24856,N_24128);
nand UO_64 (O_64,N_23784,N_24374);
nor UO_65 (O_65,N_23825,N_24217);
nand UO_66 (O_66,N_24689,N_24007);
and UO_67 (O_67,N_24155,N_24478);
nand UO_68 (O_68,N_24768,N_23968);
or UO_69 (O_69,N_24778,N_24578);
and UO_70 (O_70,N_24717,N_24659);
or UO_71 (O_71,N_24628,N_24006);
nand UO_72 (O_72,N_24440,N_24299);
xor UO_73 (O_73,N_24731,N_23937);
or UO_74 (O_74,N_24958,N_24457);
or UO_75 (O_75,N_24406,N_24445);
nor UO_76 (O_76,N_23942,N_24125);
or UO_77 (O_77,N_24624,N_24197);
xnor UO_78 (O_78,N_24329,N_24589);
nand UO_79 (O_79,N_24660,N_24316);
or UO_80 (O_80,N_24084,N_24411);
xor UO_81 (O_81,N_24512,N_24805);
nor UO_82 (O_82,N_24326,N_24592);
or UO_83 (O_83,N_23853,N_24567);
or UO_84 (O_84,N_24271,N_24887);
xnor UO_85 (O_85,N_24181,N_23920);
nor UO_86 (O_86,N_24204,N_23793);
and UO_87 (O_87,N_24306,N_24606);
and UO_88 (O_88,N_24139,N_23835);
or UO_89 (O_89,N_24910,N_24280);
nand UO_90 (O_90,N_24189,N_24102);
xnor UO_91 (O_91,N_24766,N_23995);
nor UO_92 (O_92,N_24192,N_23850);
nand UO_93 (O_93,N_24894,N_23764);
nor UO_94 (O_94,N_23971,N_24977);
nand UO_95 (O_95,N_24227,N_24131);
xor UO_96 (O_96,N_23844,N_24570);
nand UO_97 (O_97,N_23828,N_24331);
or UO_98 (O_98,N_24523,N_24203);
and UO_99 (O_99,N_24134,N_23903);
or UO_100 (O_100,N_24807,N_24816);
xor UO_101 (O_101,N_23964,N_23901);
or UO_102 (O_102,N_24249,N_23882);
nand UO_103 (O_103,N_24981,N_24866);
nand UO_104 (O_104,N_24247,N_24119);
nor UO_105 (O_105,N_24978,N_24549);
or UO_106 (O_106,N_24458,N_24730);
xnor UO_107 (O_107,N_24202,N_24662);
xor UO_108 (O_108,N_24051,N_24022);
xnor UO_109 (O_109,N_24373,N_24895);
nand UO_110 (O_110,N_24547,N_24771);
nand UO_111 (O_111,N_24556,N_23821);
xor UO_112 (O_112,N_24738,N_24244);
xnor UO_113 (O_113,N_24988,N_24175);
nand UO_114 (O_114,N_23928,N_23872);
nand UO_115 (O_115,N_23939,N_24231);
nor UO_116 (O_116,N_24307,N_23795);
nor UO_117 (O_117,N_24312,N_24147);
and UO_118 (O_118,N_24148,N_24464);
and UO_119 (O_119,N_24205,N_24799);
nand UO_120 (O_120,N_24101,N_24944);
nand UO_121 (O_121,N_23857,N_24777);
nand UO_122 (O_122,N_24124,N_24982);
or UO_123 (O_123,N_24210,N_24710);
xnor UO_124 (O_124,N_24743,N_24994);
nand UO_125 (O_125,N_23803,N_24359);
nor UO_126 (O_126,N_23948,N_24330);
or UO_127 (O_127,N_24713,N_24546);
and UO_128 (O_128,N_24390,N_23779);
nand UO_129 (O_129,N_23931,N_23819);
and UO_130 (O_130,N_24946,N_24577);
and UO_131 (O_131,N_24955,N_24970);
nor UO_132 (O_132,N_23785,N_24094);
nand UO_133 (O_133,N_23962,N_24603);
nor UO_134 (O_134,N_24183,N_24248);
nand UO_135 (O_135,N_24828,N_23781);
or UO_136 (O_136,N_24648,N_23909);
and UO_137 (O_137,N_24468,N_24700);
or UO_138 (O_138,N_24922,N_23786);
xor UO_139 (O_139,N_24645,N_24976);
xor UO_140 (O_140,N_23755,N_24166);
xor UO_141 (O_141,N_23992,N_23831);
and UO_142 (O_142,N_24372,N_24538);
and UO_143 (O_143,N_23990,N_24225);
or UO_144 (O_144,N_24725,N_24379);
nor UO_145 (O_145,N_24078,N_24173);
nor UO_146 (O_146,N_24465,N_24727);
and UO_147 (O_147,N_24888,N_24834);
and UO_148 (O_148,N_24772,N_24211);
xnor UO_149 (O_149,N_24246,N_24542);
nand UO_150 (O_150,N_24493,N_24968);
nand UO_151 (O_151,N_23769,N_24703);
xnor UO_152 (O_152,N_24399,N_24522);
or UO_153 (O_153,N_24886,N_24284);
and UO_154 (O_154,N_24190,N_24149);
nand UO_155 (O_155,N_24055,N_24971);
or UO_156 (O_156,N_24126,N_24198);
nor UO_157 (O_157,N_24448,N_23908);
xnor UO_158 (O_158,N_23972,N_24692);
nor UO_159 (O_159,N_24511,N_24282);
nand UO_160 (O_160,N_24414,N_24626);
xnor UO_161 (O_161,N_24845,N_24063);
or UO_162 (O_162,N_24686,N_24791);
xor UO_163 (O_163,N_24025,N_24762);
xnor UO_164 (O_164,N_24721,N_23840);
or UO_165 (O_165,N_24947,N_24786);
nor UO_166 (O_166,N_24891,N_24951);
nand UO_167 (O_167,N_23789,N_24999);
or UO_168 (O_168,N_24759,N_23930);
nor UO_169 (O_169,N_24165,N_24296);
or UO_170 (O_170,N_24381,N_24983);
xor UO_171 (O_171,N_24884,N_23974);
and UO_172 (O_172,N_24524,N_23805);
and UO_173 (O_173,N_24669,N_24683);
nor UO_174 (O_174,N_24230,N_24953);
nand UO_175 (O_175,N_24355,N_23940);
nand UO_176 (O_176,N_24898,N_24521);
or UO_177 (O_177,N_24042,N_24600);
or UO_178 (O_178,N_23843,N_24528);
xnor UO_179 (O_179,N_24705,N_24897);
xor UO_180 (O_180,N_24054,N_24694);
or UO_181 (O_181,N_24853,N_24661);
and UO_182 (O_182,N_24543,N_23938);
nand UO_183 (O_183,N_23936,N_24403);
xor UO_184 (O_184,N_24377,N_24009);
and UO_185 (O_185,N_24868,N_24819);
xor UO_186 (O_186,N_23780,N_23775);
xnor UO_187 (O_187,N_23902,N_24472);
and UO_188 (O_188,N_23788,N_24150);
and UO_189 (O_189,N_24485,N_24494);
nand UO_190 (O_190,N_24752,N_24962);
and UO_191 (O_191,N_23998,N_24106);
xor UO_192 (O_192,N_24264,N_23907);
or UO_193 (O_193,N_23878,N_23876);
and UO_194 (O_194,N_24687,N_23979);
xnor UO_195 (O_195,N_24785,N_23776);
xor UO_196 (O_196,N_24323,N_24532);
or UO_197 (O_197,N_24407,N_24251);
xnor UO_198 (O_198,N_24666,N_23967);
nand UO_199 (O_199,N_24975,N_24876);
nand UO_200 (O_200,N_24402,N_23873);
xor UO_201 (O_201,N_24276,N_24665);
or UO_202 (O_202,N_24254,N_23801);
or UO_203 (O_203,N_23827,N_24739);
xnor UO_204 (O_204,N_24095,N_24568);
and UO_205 (O_205,N_24972,N_23982);
or UO_206 (O_206,N_23863,N_24114);
nor UO_207 (O_207,N_24934,N_24028);
or UO_208 (O_208,N_23871,N_24823);
and UO_209 (O_209,N_24174,N_24991);
nor UO_210 (O_210,N_24901,N_24112);
or UO_211 (O_211,N_24245,N_23924);
and UO_212 (O_212,N_23770,N_24942);
nor UO_213 (O_213,N_24180,N_24560);
xnor UO_214 (O_214,N_24072,N_24057);
or UO_215 (O_215,N_24680,N_24920);
and UO_216 (O_216,N_24671,N_24608);
xor UO_217 (O_217,N_24300,N_24928);
xnor UO_218 (O_218,N_24872,N_23848);
and UO_219 (O_219,N_24881,N_24423);
or UO_220 (O_220,N_24926,N_24917);
nand UO_221 (O_221,N_24641,N_24010);
or UO_222 (O_222,N_24497,N_24930);
xnor UO_223 (O_223,N_23799,N_24837);
nand UO_224 (O_224,N_24744,N_23919);
or UO_225 (O_225,N_24614,N_24363);
xor UO_226 (O_226,N_24745,N_24143);
and UO_227 (O_227,N_24599,N_24594);
and UO_228 (O_228,N_23888,N_24815);
and UO_229 (O_229,N_24818,N_24564);
nand UO_230 (O_230,N_24236,N_24784);
xor UO_231 (O_231,N_23796,N_23790);
nor UO_232 (O_232,N_23927,N_24722);
nand UO_233 (O_233,N_24921,N_24961);
or UO_234 (O_234,N_24220,N_24366);
and UO_235 (O_235,N_24430,N_24548);
and UO_236 (O_236,N_24076,N_24332);
xnor UO_237 (O_237,N_24302,N_24215);
nor UO_238 (O_238,N_24890,N_24408);
or UO_239 (O_239,N_24663,N_23759);
xor UO_240 (O_240,N_24840,N_23947);
xnor UO_241 (O_241,N_24442,N_24885);
xnor UO_242 (O_242,N_24158,N_24672);
or UO_243 (O_243,N_24322,N_24481);
xor UO_244 (O_244,N_23832,N_24966);
and UO_245 (O_245,N_24848,N_24261);
or UO_246 (O_246,N_23866,N_23933);
nor UO_247 (O_247,N_24118,N_24169);
nand UO_248 (O_248,N_23950,N_24291);
nor UO_249 (O_249,N_24576,N_23960);
nand UO_250 (O_250,N_24882,N_23894);
nand UO_251 (O_251,N_23926,N_24317);
xnor UO_252 (O_252,N_24446,N_24151);
or UO_253 (O_253,N_24698,N_24957);
or UO_254 (O_254,N_24038,N_24188);
xor UO_255 (O_255,N_23988,N_24896);
and UO_256 (O_256,N_24630,N_24364);
xnor UO_257 (O_257,N_24207,N_23774);
nor UO_258 (O_258,N_24193,N_23859);
and UO_259 (O_259,N_24653,N_24679);
or UO_260 (O_260,N_24266,N_24221);
xnor UO_261 (O_261,N_24985,N_24135);
and UO_262 (O_262,N_24501,N_24431);
xor UO_263 (O_263,N_24804,N_24466);
nand UO_264 (O_264,N_24369,N_23750);
nor UO_265 (O_265,N_24450,N_24066);
or UO_266 (O_266,N_24758,N_24021);
nor UO_267 (O_267,N_24664,N_24699);
and UO_268 (O_268,N_24232,N_24311);
xnor UO_269 (O_269,N_23946,N_23861);
or UO_270 (O_270,N_23887,N_24839);
xnor UO_271 (O_271,N_24488,N_24422);
nand UO_272 (O_272,N_24824,N_24087);
and UO_273 (O_273,N_24562,N_24167);
or UO_274 (O_274,N_24842,N_24638);
or UO_275 (O_275,N_23983,N_24011);
nand UO_276 (O_276,N_24670,N_24827);
nor UO_277 (O_277,N_24437,N_24340);
xor UO_278 (O_278,N_24305,N_24269);
nand UO_279 (O_279,N_24631,N_24486);
and UO_280 (O_280,N_24289,N_24989);
xor UO_281 (O_281,N_24609,N_24105);
xor UO_282 (O_282,N_24161,N_24677);
nand UO_283 (O_283,N_23757,N_24144);
and UO_284 (O_284,N_23952,N_23762);
or UO_285 (O_285,N_24234,N_24243);
and UO_286 (O_286,N_23753,N_24854);
and UO_287 (O_287,N_24857,N_24362);
or UO_288 (O_288,N_24111,N_24413);
nor UO_289 (O_289,N_24726,N_24252);
nor UO_290 (O_290,N_24790,N_23767);
nor UO_291 (O_291,N_23991,N_24908);
nor UO_292 (O_292,N_24199,N_24865);
xnor UO_293 (O_293,N_24438,N_24779);
xor UO_294 (O_294,N_24925,N_24048);
or UO_295 (O_295,N_24580,N_23833);
nor UO_296 (O_296,N_24187,N_24761);
and UO_297 (O_297,N_24964,N_24176);
and UO_298 (O_298,N_24195,N_24081);
nor UO_299 (O_299,N_23879,N_23855);
nand UO_300 (O_300,N_24850,N_24843);
nor UO_301 (O_301,N_24097,N_24474);
nand UO_302 (O_302,N_24099,N_24219);
or UO_303 (O_303,N_23754,N_24965);
nor UO_304 (O_304,N_24426,N_24419);
nor UO_305 (O_305,N_24350,N_24405);
nor UO_306 (O_306,N_24987,N_24079);
nand UO_307 (O_307,N_24821,N_24121);
xnor UO_308 (O_308,N_24382,N_23883);
or UO_309 (O_309,N_24336,N_24002);
nand UO_310 (O_310,N_24421,N_24080);
xor UO_311 (O_311,N_24554,N_24851);
or UO_312 (O_312,N_23847,N_24702);
xnor UO_313 (O_313,N_24574,N_24428);
nand UO_314 (O_314,N_24186,N_24831);
and UO_315 (O_315,N_24877,N_24914);
xnor UO_316 (O_316,N_24642,N_24749);
nor UO_317 (O_317,N_24091,N_24708);
nor UO_318 (O_318,N_23944,N_24637);
and UO_319 (O_319,N_23791,N_24658);
or UO_320 (O_320,N_24682,N_24846);
nand UO_321 (O_321,N_24303,N_24903);
or UO_322 (O_322,N_24058,N_23815);
and UO_323 (O_323,N_24632,N_24935);
xnor UO_324 (O_324,N_24153,N_24878);
xor UO_325 (O_325,N_24253,N_24294);
or UO_326 (O_326,N_24770,N_23985);
or UO_327 (O_327,N_23771,N_24598);
and UO_328 (O_328,N_24633,N_24397);
xnor UO_329 (O_329,N_24904,N_24588);
nand UO_330 (O_330,N_24849,N_23765);
xor UO_331 (O_331,N_24222,N_24455);
or UO_332 (O_332,N_24425,N_23808);
nand UO_333 (O_333,N_24082,N_24674);
and UO_334 (O_334,N_24342,N_24714);
nor UO_335 (O_335,N_24287,N_24992);
nor UO_336 (O_336,N_24590,N_24919);
or UO_337 (O_337,N_23989,N_24056);
nor UO_338 (O_338,N_24410,N_23858);
or UO_339 (O_339,N_24471,N_24343);
nand UO_340 (O_340,N_24960,N_23963);
nand UO_341 (O_341,N_23834,N_24858);
or UO_342 (O_342,N_24695,N_24035);
or UO_343 (O_343,N_24707,N_24467);
or UO_344 (O_344,N_24320,N_23925);
nand UO_345 (O_345,N_23778,N_24718);
and UO_346 (O_346,N_24810,N_24997);
xor UO_347 (O_347,N_24803,N_24751);
and UO_348 (O_348,N_24820,N_23885);
xnor UO_349 (O_349,N_24755,N_24484);
and UO_350 (O_350,N_24052,N_24313);
or UO_351 (O_351,N_24218,N_24324);
xor UO_352 (O_352,N_24979,N_24108);
nor UO_353 (O_353,N_24575,N_24156);
xor UO_354 (O_354,N_24389,N_24529);
or UO_355 (O_355,N_24242,N_24654);
or UO_356 (O_356,N_23923,N_24813);
nor UO_357 (O_357,N_24059,N_23987);
or UO_358 (O_358,N_24875,N_24229);
nand UO_359 (O_359,N_24506,N_24841);
and UO_360 (O_360,N_24420,N_24646);
nor UO_361 (O_361,N_24889,N_24764);
nand UO_362 (O_362,N_23849,N_24863);
nor UO_363 (O_363,N_24912,N_24375);
nor UO_364 (O_364,N_24476,N_24527);
and UO_365 (O_365,N_23917,N_24003);
xor UO_366 (O_366,N_23802,N_24117);
nand UO_367 (O_367,N_24760,N_24507);
nor UO_368 (O_368,N_24498,N_24138);
nand UO_369 (O_369,N_24675,N_23896);
and UO_370 (O_370,N_24774,N_24335);
or UO_371 (O_371,N_24281,N_24435);
nand UO_372 (O_372,N_24179,N_24071);
nor UO_373 (O_373,N_24809,N_24415);
xnor UO_374 (O_374,N_24974,N_24899);
nand UO_375 (O_375,N_23869,N_24927);
nand UO_376 (O_376,N_24288,N_24530);
or UO_377 (O_377,N_24929,N_24107);
or UO_378 (O_378,N_23804,N_24395);
nand UO_379 (O_379,N_24239,N_24667);
and UO_380 (O_380,N_24285,N_24321);
or UO_381 (O_381,N_24510,N_23941);
nor UO_382 (O_382,N_24386,N_23813);
nand UO_383 (O_383,N_24053,N_24757);
nand UO_384 (O_384,N_24490,N_24693);
nor UO_385 (O_385,N_24644,N_23980);
nand UO_386 (O_386,N_23905,N_23814);
or UO_387 (O_387,N_23824,N_24194);
nor UO_388 (O_388,N_24635,N_24060);
and UO_389 (O_389,N_24470,N_23958);
xor UO_390 (O_390,N_23773,N_24684);
and UO_391 (O_391,N_24544,N_24657);
nor UO_392 (O_392,N_24040,N_24074);
xor UO_393 (O_393,N_24712,N_23811);
and UO_394 (O_394,N_24595,N_23890);
xnor UO_395 (O_395,N_24649,N_23761);
nor UO_396 (O_396,N_24940,N_23893);
nor UO_397 (O_397,N_23838,N_24238);
nor UO_398 (O_398,N_24380,N_23932);
and UO_399 (O_399,N_24826,N_24127);
xor UO_400 (O_400,N_24618,N_24298);
nand UO_401 (O_401,N_24715,N_23826);
or UO_402 (O_402,N_24518,N_24874);
nor UO_403 (O_403,N_23934,N_24113);
and UO_404 (O_404,N_23841,N_24909);
nand UO_405 (O_405,N_24093,N_24213);
xor UO_406 (O_406,N_24333,N_24650);
nand UO_407 (O_407,N_24475,N_24424);
xnor UO_408 (O_408,N_24171,N_24376);
nand UO_409 (O_409,N_24393,N_24237);
xor UO_410 (O_410,N_24732,N_24685);
or UO_411 (O_411,N_23867,N_24370);
or UO_412 (O_412,N_24429,N_24491);
and UO_413 (O_413,N_23999,N_24800);
nand UO_414 (O_414,N_24133,N_23830);
nand UO_415 (O_415,N_24371,N_24226);
nor UO_416 (O_416,N_24719,N_24045);
nor UO_417 (O_417,N_24352,N_24137);
xor UO_418 (O_418,N_23884,N_24172);
and UO_419 (O_419,N_24505,N_24583);
xnor UO_420 (O_420,N_24473,N_24096);
nand UO_421 (O_421,N_24020,N_24318);
nor UO_422 (O_422,N_24109,N_24338);
xor UO_423 (O_423,N_24434,N_24571);
nor UO_424 (O_424,N_24339,N_23794);
nand UO_425 (O_425,N_24798,N_24587);
xnor UO_426 (O_426,N_23943,N_24923);
xnor UO_427 (O_427,N_23929,N_24400);
or UO_428 (O_428,N_24152,N_23981);
nor UO_429 (O_429,N_24295,N_24579);
nor UO_430 (O_430,N_23961,N_24479);
or UO_431 (O_431,N_24100,N_24676);
or UO_432 (O_432,N_24651,N_24535);
and UO_433 (O_433,N_24534,N_24796);
or UO_434 (O_434,N_24459,N_24065);
xor UO_435 (O_435,N_24622,N_24301);
nand UO_436 (O_436,N_24835,N_24584);
and UO_437 (O_437,N_24337,N_24417);
or UO_438 (O_438,N_24036,N_23892);
and UO_439 (O_439,N_23766,N_24852);
nor UO_440 (O_440,N_23860,N_24867);
nor UO_441 (O_441,N_24272,N_24267);
and UO_442 (O_442,N_24984,N_24085);
nor UO_443 (O_443,N_24995,N_24748);
nor UO_444 (O_444,N_23783,N_24775);
nor UO_445 (O_445,N_24990,N_24862);
and UO_446 (O_446,N_24688,N_24433);
nor UO_447 (O_447,N_24050,N_23763);
and UO_448 (O_448,N_24325,N_24569);
nand UO_449 (O_449,N_24504,N_23823);
and UO_450 (O_450,N_24508,N_23846);
or UO_451 (O_451,N_24652,N_23852);
or UO_452 (O_452,N_24742,N_24754);
or UO_453 (O_453,N_24619,N_24737);
and UO_454 (O_454,N_24444,N_24023);
nand UO_455 (O_455,N_24345,N_23856);
or UO_456 (O_456,N_23874,N_24427);
nand UO_457 (O_457,N_24351,N_24701);
or UO_458 (O_458,N_24709,N_23868);
and UO_459 (O_459,N_24309,N_24392);
and UO_460 (O_460,N_24519,N_24613);
nor UO_461 (O_461,N_24344,N_24178);
and UO_462 (O_462,N_24461,N_23756);
nor UO_463 (O_463,N_24394,N_23906);
nand UO_464 (O_464,N_24315,N_23984);
nand UO_465 (O_465,N_24354,N_23918);
nand UO_466 (O_466,N_24033,N_23751);
and UO_467 (O_467,N_24711,N_24604);
or UO_468 (O_468,N_24537,N_24747);
nor UO_469 (O_469,N_24911,N_24454);
and UO_470 (O_470,N_24157,N_23817);
and UO_471 (O_471,N_24334,N_24555);
or UO_472 (O_472,N_24557,N_24690);
nor UO_473 (O_473,N_24932,N_24639);
nor UO_474 (O_474,N_23854,N_24275);
or UO_475 (O_475,N_24314,N_24520);
nor UO_476 (O_476,N_24625,N_24830);
and UO_477 (O_477,N_24001,N_24032);
xnor UO_478 (O_478,N_24610,N_24802);
and UO_479 (O_479,N_24541,N_23836);
and UO_480 (O_480,N_24883,N_23886);
nand UO_481 (O_481,N_24453,N_24279);
nand UO_482 (O_482,N_24924,N_24952);
xor UO_483 (O_483,N_24441,N_24046);
and UO_484 (O_484,N_24795,N_23969);
and UO_485 (O_485,N_24495,N_24164);
nor UO_486 (O_486,N_24224,N_24787);
nor UO_487 (O_487,N_24409,N_24559);
and UO_488 (O_488,N_24765,N_24558);
xor UO_489 (O_489,N_24933,N_23818);
xnor UO_490 (O_490,N_23777,N_24525);
and UO_491 (O_491,N_24341,N_23977);
and UO_492 (O_492,N_24513,N_24353);
or UO_493 (O_493,N_23956,N_24621);
and UO_494 (O_494,N_24634,N_24469);
and UO_495 (O_495,N_24460,N_23898);
nor UO_496 (O_496,N_24793,N_24483);
xnor UO_497 (O_497,N_23797,N_24871);
or UO_498 (O_498,N_24954,N_24360);
nor UO_499 (O_499,N_23954,N_23965);
xnor UO_500 (O_500,N_24265,N_24767);
and UO_501 (O_501,N_24083,N_24502);
xnor UO_502 (O_502,N_24729,N_24061);
or UO_503 (O_503,N_24880,N_24357);
nor UO_504 (O_504,N_23966,N_24077);
nor UO_505 (O_505,N_24836,N_24829);
nand UO_506 (O_506,N_24531,N_24723);
nand UO_507 (O_507,N_24860,N_24566);
nor UO_508 (O_508,N_23782,N_24773);
or UO_509 (O_509,N_24160,N_24017);
or UO_510 (O_510,N_24514,N_24893);
and UO_511 (O_511,N_24636,N_24273);
xnor UO_512 (O_512,N_24586,N_24041);
or UO_513 (O_513,N_23845,N_24627);
nand UO_514 (O_514,N_24136,N_24049);
or UO_515 (O_515,N_23837,N_24550);
or UO_516 (O_516,N_24696,N_24367);
or UO_517 (O_517,N_24623,N_24553);
nand UO_518 (O_518,N_24673,N_23820);
xnor UO_519 (O_519,N_24597,N_24235);
nand UO_520 (O_520,N_24482,N_24263);
or UO_521 (O_521,N_24735,N_24733);
and UO_522 (O_522,N_24905,N_23973);
and UO_523 (O_523,N_23916,N_24750);
nor UO_524 (O_524,N_24517,N_24044);
xnor UO_525 (O_525,N_24573,N_24788);
or UO_526 (O_526,N_24825,N_24551);
xor UO_527 (O_527,N_24015,N_23945);
or UO_528 (O_528,N_24212,N_24451);
and UO_529 (O_529,N_23881,N_23870);
xor UO_530 (O_530,N_24396,N_24262);
nand UO_531 (O_531,N_24024,N_23807);
nand UO_532 (O_532,N_24993,N_24064);
xnor UO_533 (O_533,N_24447,N_24310);
nand UO_534 (O_534,N_24255,N_24387);
nand UO_535 (O_535,N_24915,N_24668);
xnor UO_536 (O_536,N_24391,N_24278);
nand UO_537 (O_537,N_24120,N_23865);
or UO_538 (O_538,N_24418,N_24563);
xnor UO_539 (O_539,N_24129,N_24170);
and UO_540 (O_540,N_23829,N_24741);
nor UO_541 (O_541,N_24104,N_24792);
xnor UO_542 (O_542,N_24293,N_24401);
nand UO_543 (O_543,N_24146,N_23959);
and UO_544 (O_544,N_24913,N_24797);
nand UO_545 (O_545,N_24346,N_24185);
or UO_546 (O_546,N_24907,N_24980);
and UO_547 (O_547,N_23810,N_24214);
nand UO_548 (O_548,N_24159,N_24365);
nand UO_549 (O_549,N_24140,N_24591);
nand UO_550 (O_550,N_24832,N_24062);
nand UO_551 (O_551,N_24596,N_24817);
nor UO_552 (O_552,N_23875,N_23955);
nor UO_553 (O_553,N_24740,N_24216);
nand UO_554 (O_554,N_24184,N_24008);
nor UO_555 (O_555,N_24384,N_24916);
nor UO_556 (O_556,N_24640,N_24540);
nor UO_557 (O_557,N_24782,N_24601);
nand UO_558 (O_558,N_24196,N_24240);
nand UO_559 (O_559,N_24388,N_24728);
nor UO_560 (O_560,N_24292,N_24545);
and UO_561 (O_561,N_24088,N_24582);
nand UO_562 (O_562,N_23864,N_23787);
nor UO_563 (O_563,N_24070,N_24132);
or UO_564 (O_564,N_24681,N_24356);
or UO_565 (O_565,N_24931,N_24873);
xor UO_566 (O_566,N_23891,N_24012);
nand UO_567 (O_567,N_24098,N_24029);
nor UO_568 (O_568,N_24620,N_24027);
xnor UO_569 (O_569,N_23851,N_24452);
and UO_570 (O_570,N_24996,N_23842);
xor UO_571 (O_571,N_24615,N_24861);
nand UO_572 (O_572,N_24607,N_24776);
nor UO_573 (O_573,N_24030,N_24492);
xor UO_574 (O_574,N_24794,N_24086);
or UO_575 (O_575,N_24268,N_24539);
xor UO_576 (O_576,N_23904,N_24967);
or UO_577 (O_577,N_24720,N_24864);
xnor UO_578 (O_578,N_24358,N_24937);
nor UO_579 (O_579,N_24945,N_24177);
and UO_580 (O_580,N_24585,N_24258);
nand UO_581 (O_581,N_24647,N_24724);
xnor UO_582 (O_582,N_24383,N_24047);
nand UO_583 (O_583,N_24605,N_23970);
or UO_584 (O_584,N_24209,N_24039);
nor UO_585 (O_585,N_24998,N_24516);
or UO_586 (O_586,N_24462,N_24503);
and UO_587 (O_587,N_23915,N_23889);
nor UO_588 (O_588,N_24439,N_23877);
nand UO_589 (O_589,N_24806,N_24449);
and UO_590 (O_590,N_24616,N_24043);
and UO_591 (O_591,N_23899,N_23768);
nor UO_592 (O_592,N_24145,N_23994);
nand UO_593 (O_593,N_24870,N_23862);
nor UO_594 (O_594,N_24879,N_24416);
nand UO_595 (O_595,N_24814,N_24327);
and UO_596 (O_596,N_24812,N_24533);
xor UO_597 (O_597,N_23993,N_24847);
nand UO_598 (O_598,N_24090,N_24162);
nor UO_599 (O_599,N_24361,N_24801);
nor UO_600 (O_600,N_23978,N_24552);
xor UO_601 (O_601,N_24308,N_24656);
or UO_602 (O_602,N_24973,N_23897);
or UO_603 (O_603,N_23921,N_23975);
nor UO_604 (O_604,N_24123,N_24833);
nand UO_605 (O_605,N_24034,N_24780);
xnor UO_606 (O_606,N_24168,N_24499);
nor UO_607 (O_607,N_24259,N_24385);
or UO_608 (O_608,N_24716,N_23798);
nand UO_609 (O_609,N_24509,N_23880);
or UO_610 (O_610,N_24297,N_23758);
and UO_611 (O_611,N_24116,N_24319);
nand UO_612 (O_612,N_24286,N_23913);
nor UO_613 (O_613,N_24691,N_24200);
nor UO_614 (O_614,N_24593,N_24617);
nand UO_615 (O_615,N_24115,N_23760);
xnor UO_616 (O_616,N_24480,N_24602);
xnor UO_617 (O_617,N_24068,N_24018);
nor UO_618 (O_618,N_24228,N_24037);
or UO_619 (O_619,N_24855,N_24629);
nand UO_620 (O_620,N_24969,N_24182);
nor UO_621 (O_621,N_24489,N_24734);
and UO_622 (O_622,N_24349,N_23839);
nand UO_623 (O_623,N_24223,N_23951);
nor UO_624 (O_624,N_24233,N_24256);
and UO_625 (O_625,N_23906,N_24872);
or UO_626 (O_626,N_24028,N_23805);
nand UO_627 (O_627,N_24686,N_23875);
nor UO_628 (O_628,N_23894,N_23767);
or UO_629 (O_629,N_24514,N_24531);
nor UO_630 (O_630,N_24856,N_24607);
and UO_631 (O_631,N_24979,N_23753);
xnor UO_632 (O_632,N_24178,N_24359);
or UO_633 (O_633,N_24711,N_24597);
or UO_634 (O_634,N_24580,N_24967);
xnor UO_635 (O_635,N_24542,N_24341);
nand UO_636 (O_636,N_24324,N_24568);
and UO_637 (O_637,N_24884,N_23976);
or UO_638 (O_638,N_23801,N_24474);
and UO_639 (O_639,N_24226,N_24130);
xor UO_640 (O_640,N_24349,N_24045);
nor UO_641 (O_641,N_24063,N_24483);
nor UO_642 (O_642,N_23757,N_24426);
xor UO_643 (O_643,N_24018,N_24382);
nand UO_644 (O_644,N_24649,N_24632);
and UO_645 (O_645,N_24914,N_24329);
or UO_646 (O_646,N_24004,N_24372);
and UO_647 (O_647,N_24379,N_24734);
or UO_648 (O_648,N_23854,N_24245);
nand UO_649 (O_649,N_24135,N_23869);
nor UO_650 (O_650,N_24008,N_24682);
nor UO_651 (O_651,N_24694,N_24584);
xor UO_652 (O_652,N_24690,N_23993);
or UO_653 (O_653,N_24878,N_24423);
or UO_654 (O_654,N_24536,N_23943);
nand UO_655 (O_655,N_24597,N_23977);
or UO_656 (O_656,N_24433,N_23941);
or UO_657 (O_657,N_23775,N_23925);
xnor UO_658 (O_658,N_24943,N_24137);
or UO_659 (O_659,N_24911,N_23835);
nand UO_660 (O_660,N_24242,N_23914);
xor UO_661 (O_661,N_23815,N_23988);
xnor UO_662 (O_662,N_24776,N_24529);
and UO_663 (O_663,N_24928,N_24037);
or UO_664 (O_664,N_24125,N_24853);
and UO_665 (O_665,N_24532,N_24832);
xor UO_666 (O_666,N_23770,N_24790);
nand UO_667 (O_667,N_24387,N_23979);
xnor UO_668 (O_668,N_24437,N_24739);
or UO_669 (O_669,N_23933,N_24007);
xor UO_670 (O_670,N_23972,N_24429);
xor UO_671 (O_671,N_24393,N_24482);
nor UO_672 (O_672,N_24422,N_24345);
xor UO_673 (O_673,N_24382,N_24772);
nand UO_674 (O_674,N_24302,N_24677);
nand UO_675 (O_675,N_24572,N_24524);
nand UO_676 (O_676,N_24119,N_24251);
nor UO_677 (O_677,N_24986,N_24633);
or UO_678 (O_678,N_24671,N_24221);
and UO_679 (O_679,N_23852,N_24236);
and UO_680 (O_680,N_24308,N_24860);
or UO_681 (O_681,N_24495,N_24412);
or UO_682 (O_682,N_24709,N_24224);
and UO_683 (O_683,N_24762,N_24073);
nand UO_684 (O_684,N_23957,N_24720);
nor UO_685 (O_685,N_24394,N_24633);
nand UO_686 (O_686,N_24904,N_24815);
nand UO_687 (O_687,N_24179,N_24388);
xor UO_688 (O_688,N_24672,N_24942);
nor UO_689 (O_689,N_23831,N_24880);
and UO_690 (O_690,N_23930,N_24754);
and UO_691 (O_691,N_24037,N_24651);
or UO_692 (O_692,N_23895,N_24042);
nor UO_693 (O_693,N_24169,N_24605);
xnor UO_694 (O_694,N_24144,N_24249);
and UO_695 (O_695,N_23934,N_23945);
nand UO_696 (O_696,N_24697,N_24966);
and UO_697 (O_697,N_23769,N_24859);
xor UO_698 (O_698,N_24416,N_23909);
nor UO_699 (O_699,N_24312,N_24219);
xor UO_700 (O_700,N_24960,N_23811);
nand UO_701 (O_701,N_24251,N_23840);
or UO_702 (O_702,N_24409,N_23852);
or UO_703 (O_703,N_24250,N_24681);
or UO_704 (O_704,N_24058,N_24004);
nand UO_705 (O_705,N_24385,N_23986);
xnor UO_706 (O_706,N_24598,N_24278);
and UO_707 (O_707,N_24125,N_24366);
xor UO_708 (O_708,N_24938,N_23812);
nand UO_709 (O_709,N_24544,N_24595);
and UO_710 (O_710,N_24395,N_24426);
nand UO_711 (O_711,N_24681,N_24877);
nand UO_712 (O_712,N_24613,N_24620);
nor UO_713 (O_713,N_24643,N_24285);
nor UO_714 (O_714,N_24235,N_23854);
nor UO_715 (O_715,N_23865,N_24246);
nand UO_716 (O_716,N_23945,N_24244);
nand UO_717 (O_717,N_24076,N_23782);
and UO_718 (O_718,N_24391,N_24904);
nor UO_719 (O_719,N_24877,N_24380);
or UO_720 (O_720,N_23955,N_23828);
nor UO_721 (O_721,N_23979,N_24090);
and UO_722 (O_722,N_24731,N_23978);
and UO_723 (O_723,N_24589,N_24114);
xnor UO_724 (O_724,N_24247,N_24848);
xor UO_725 (O_725,N_23972,N_23852);
nor UO_726 (O_726,N_23774,N_24125);
nand UO_727 (O_727,N_24996,N_23903);
nand UO_728 (O_728,N_23932,N_24411);
nor UO_729 (O_729,N_23792,N_24482);
nand UO_730 (O_730,N_24373,N_24390);
xor UO_731 (O_731,N_23801,N_24517);
xnor UO_732 (O_732,N_24272,N_24489);
or UO_733 (O_733,N_23974,N_24714);
or UO_734 (O_734,N_24048,N_24690);
nor UO_735 (O_735,N_23829,N_24423);
nand UO_736 (O_736,N_24778,N_24725);
or UO_737 (O_737,N_24143,N_24533);
or UO_738 (O_738,N_24937,N_24424);
xnor UO_739 (O_739,N_24850,N_23902);
nor UO_740 (O_740,N_24157,N_24930);
nor UO_741 (O_741,N_24110,N_24557);
xor UO_742 (O_742,N_24876,N_24672);
or UO_743 (O_743,N_24448,N_24677);
nor UO_744 (O_744,N_24114,N_24948);
nor UO_745 (O_745,N_24541,N_24744);
xnor UO_746 (O_746,N_24887,N_24610);
nand UO_747 (O_747,N_24787,N_24979);
and UO_748 (O_748,N_24190,N_24263);
and UO_749 (O_749,N_24024,N_24055);
nand UO_750 (O_750,N_24613,N_24415);
or UO_751 (O_751,N_24090,N_23783);
xor UO_752 (O_752,N_24671,N_24679);
nand UO_753 (O_753,N_23768,N_24113);
or UO_754 (O_754,N_24567,N_23994);
xnor UO_755 (O_755,N_24356,N_24755);
nor UO_756 (O_756,N_24077,N_23870);
nor UO_757 (O_757,N_24457,N_24004);
nor UO_758 (O_758,N_24554,N_24158);
nand UO_759 (O_759,N_24251,N_24998);
nand UO_760 (O_760,N_23806,N_23804);
and UO_761 (O_761,N_24319,N_24362);
xnor UO_762 (O_762,N_23969,N_24689);
nand UO_763 (O_763,N_24390,N_24430);
nor UO_764 (O_764,N_24979,N_24211);
or UO_765 (O_765,N_24977,N_23818);
and UO_766 (O_766,N_24247,N_23883);
or UO_767 (O_767,N_24096,N_23969);
nor UO_768 (O_768,N_24180,N_24923);
nand UO_769 (O_769,N_23851,N_23940);
nand UO_770 (O_770,N_24735,N_24119);
nand UO_771 (O_771,N_23838,N_24244);
nand UO_772 (O_772,N_24804,N_24281);
xor UO_773 (O_773,N_23899,N_24789);
nor UO_774 (O_774,N_24274,N_23905);
and UO_775 (O_775,N_24410,N_24366);
nand UO_776 (O_776,N_23966,N_24384);
or UO_777 (O_777,N_24657,N_24456);
and UO_778 (O_778,N_24246,N_24412);
nor UO_779 (O_779,N_24481,N_24229);
xnor UO_780 (O_780,N_24614,N_24354);
xor UO_781 (O_781,N_24380,N_24108);
or UO_782 (O_782,N_24531,N_23960);
xor UO_783 (O_783,N_23836,N_24411);
nand UO_784 (O_784,N_24062,N_23927);
nand UO_785 (O_785,N_24224,N_24245);
or UO_786 (O_786,N_24061,N_24270);
or UO_787 (O_787,N_24134,N_24917);
and UO_788 (O_788,N_23779,N_24699);
and UO_789 (O_789,N_24805,N_24029);
nor UO_790 (O_790,N_24198,N_24424);
or UO_791 (O_791,N_24540,N_24795);
xor UO_792 (O_792,N_24637,N_24896);
and UO_793 (O_793,N_24615,N_24127);
xnor UO_794 (O_794,N_24493,N_24547);
xnor UO_795 (O_795,N_24266,N_23879);
nand UO_796 (O_796,N_24500,N_24202);
nor UO_797 (O_797,N_23826,N_24935);
and UO_798 (O_798,N_23777,N_24222);
xnor UO_799 (O_799,N_24416,N_24064);
xor UO_800 (O_800,N_24325,N_24269);
and UO_801 (O_801,N_24007,N_23944);
and UO_802 (O_802,N_24236,N_24211);
or UO_803 (O_803,N_23860,N_24600);
nor UO_804 (O_804,N_24919,N_24666);
or UO_805 (O_805,N_24053,N_23972);
or UO_806 (O_806,N_24869,N_24490);
xor UO_807 (O_807,N_24859,N_23940);
xor UO_808 (O_808,N_23785,N_23926);
nor UO_809 (O_809,N_24271,N_24682);
nand UO_810 (O_810,N_24370,N_24802);
or UO_811 (O_811,N_24492,N_24897);
xor UO_812 (O_812,N_24176,N_24589);
nor UO_813 (O_813,N_24310,N_24852);
nand UO_814 (O_814,N_23784,N_24488);
xnor UO_815 (O_815,N_23805,N_24965);
xor UO_816 (O_816,N_24546,N_24917);
and UO_817 (O_817,N_24799,N_24342);
xnor UO_818 (O_818,N_23945,N_24928);
xor UO_819 (O_819,N_24239,N_24072);
and UO_820 (O_820,N_23832,N_24423);
or UO_821 (O_821,N_24643,N_24909);
nor UO_822 (O_822,N_24072,N_23914);
xnor UO_823 (O_823,N_24788,N_24256);
or UO_824 (O_824,N_23909,N_24674);
or UO_825 (O_825,N_24207,N_24313);
nor UO_826 (O_826,N_24597,N_24391);
and UO_827 (O_827,N_24605,N_24664);
nor UO_828 (O_828,N_23834,N_24721);
and UO_829 (O_829,N_24958,N_24892);
or UO_830 (O_830,N_24248,N_24030);
xor UO_831 (O_831,N_23789,N_24534);
nor UO_832 (O_832,N_24418,N_24823);
nand UO_833 (O_833,N_24447,N_24945);
or UO_834 (O_834,N_24656,N_24590);
or UO_835 (O_835,N_24263,N_24598);
or UO_836 (O_836,N_23874,N_24598);
or UO_837 (O_837,N_24562,N_23862);
nor UO_838 (O_838,N_24786,N_24662);
nand UO_839 (O_839,N_24660,N_24181);
and UO_840 (O_840,N_24382,N_24471);
nor UO_841 (O_841,N_24542,N_24989);
nand UO_842 (O_842,N_23946,N_23950);
nor UO_843 (O_843,N_24976,N_24691);
nand UO_844 (O_844,N_24830,N_24701);
or UO_845 (O_845,N_24166,N_23850);
nor UO_846 (O_846,N_24964,N_23933);
and UO_847 (O_847,N_24384,N_24593);
xnor UO_848 (O_848,N_23872,N_24407);
and UO_849 (O_849,N_24030,N_24295);
and UO_850 (O_850,N_24356,N_24100);
nor UO_851 (O_851,N_24859,N_24785);
or UO_852 (O_852,N_24178,N_24828);
xor UO_853 (O_853,N_24766,N_24729);
xnor UO_854 (O_854,N_24713,N_24302);
and UO_855 (O_855,N_24864,N_24968);
nand UO_856 (O_856,N_23920,N_24340);
nor UO_857 (O_857,N_24308,N_23838);
or UO_858 (O_858,N_24107,N_23978);
xor UO_859 (O_859,N_24640,N_23802);
or UO_860 (O_860,N_23889,N_24174);
nor UO_861 (O_861,N_23974,N_23853);
and UO_862 (O_862,N_24227,N_23949);
nor UO_863 (O_863,N_24586,N_24855);
and UO_864 (O_864,N_24453,N_24365);
nor UO_865 (O_865,N_23788,N_24711);
nand UO_866 (O_866,N_24572,N_24141);
nand UO_867 (O_867,N_24456,N_24279);
nand UO_868 (O_868,N_24440,N_24537);
or UO_869 (O_869,N_24098,N_24873);
or UO_870 (O_870,N_24221,N_24030);
nand UO_871 (O_871,N_24551,N_24693);
xor UO_872 (O_872,N_23870,N_24590);
and UO_873 (O_873,N_24062,N_24859);
nand UO_874 (O_874,N_24295,N_24370);
and UO_875 (O_875,N_24888,N_24537);
or UO_876 (O_876,N_24812,N_24695);
nand UO_877 (O_877,N_24459,N_23811);
xnor UO_878 (O_878,N_24655,N_24346);
and UO_879 (O_879,N_24799,N_24547);
nor UO_880 (O_880,N_24801,N_24048);
nor UO_881 (O_881,N_23860,N_23893);
nand UO_882 (O_882,N_23888,N_24717);
nand UO_883 (O_883,N_24526,N_24910);
xor UO_884 (O_884,N_24918,N_24217);
nor UO_885 (O_885,N_24208,N_24065);
or UO_886 (O_886,N_24744,N_24415);
xor UO_887 (O_887,N_24068,N_24481);
and UO_888 (O_888,N_24666,N_24929);
or UO_889 (O_889,N_24538,N_24603);
nand UO_890 (O_890,N_24258,N_24724);
and UO_891 (O_891,N_24014,N_24466);
nand UO_892 (O_892,N_24590,N_24479);
nand UO_893 (O_893,N_23864,N_24706);
and UO_894 (O_894,N_24402,N_24159);
or UO_895 (O_895,N_24126,N_24271);
xnor UO_896 (O_896,N_23943,N_24282);
and UO_897 (O_897,N_24760,N_24553);
and UO_898 (O_898,N_24619,N_23880);
nor UO_899 (O_899,N_24409,N_24061);
and UO_900 (O_900,N_24486,N_23922);
and UO_901 (O_901,N_24596,N_24318);
and UO_902 (O_902,N_24997,N_24427);
and UO_903 (O_903,N_24737,N_23957);
and UO_904 (O_904,N_24168,N_24975);
nor UO_905 (O_905,N_24051,N_23852);
nor UO_906 (O_906,N_24830,N_24390);
xor UO_907 (O_907,N_23960,N_24574);
nand UO_908 (O_908,N_23872,N_23975);
nor UO_909 (O_909,N_23814,N_24410);
xnor UO_910 (O_910,N_24730,N_24925);
xor UO_911 (O_911,N_23972,N_24725);
nor UO_912 (O_912,N_24747,N_24249);
nand UO_913 (O_913,N_24839,N_24883);
nand UO_914 (O_914,N_24736,N_23944);
nand UO_915 (O_915,N_24418,N_24394);
nand UO_916 (O_916,N_24814,N_24951);
xnor UO_917 (O_917,N_24369,N_24674);
nor UO_918 (O_918,N_23852,N_23990);
nor UO_919 (O_919,N_23767,N_24330);
and UO_920 (O_920,N_24070,N_24217);
and UO_921 (O_921,N_24149,N_23897);
and UO_922 (O_922,N_24724,N_24921);
and UO_923 (O_923,N_24099,N_24002);
or UO_924 (O_924,N_23850,N_24554);
or UO_925 (O_925,N_24902,N_24514);
and UO_926 (O_926,N_24129,N_24939);
xnor UO_927 (O_927,N_23886,N_24079);
nor UO_928 (O_928,N_24893,N_24506);
or UO_929 (O_929,N_23869,N_24953);
xor UO_930 (O_930,N_24731,N_24977);
nand UO_931 (O_931,N_24952,N_24435);
nand UO_932 (O_932,N_24886,N_24815);
nand UO_933 (O_933,N_24469,N_24100);
nand UO_934 (O_934,N_24492,N_24337);
and UO_935 (O_935,N_24445,N_24743);
or UO_936 (O_936,N_24990,N_24541);
nor UO_937 (O_937,N_24614,N_24740);
nor UO_938 (O_938,N_24050,N_23976);
or UO_939 (O_939,N_24826,N_24386);
nand UO_940 (O_940,N_23788,N_23855);
or UO_941 (O_941,N_23956,N_24193);
xor UO_942 (O_942,N_24879,N_23825);
xor UO_943 (O_943,N_24330,N_24588);
nor UO_944 (O_944,N_24180,N_23846);
nand UO_945 (O_945,N_23884,N_23764);
xor UO_946 (O_946,N_24110,N_24778);
xor UO_947 (O_947,N_24997,N_24419);
or UO_948 (O_948,N_24425,N_23959);
and UO_949 (O_949,N_24209,N_24278);
nand UO_950 (O_950,N_24712,N_24341);
nand UO_951 (O_951,N_24790,N_24069);
xnor UO_952 (O_952,N_24443,N_24211);
nand UO_953 (O_953,N_24648,N_24815);
nor UO_954 (O_954,N_24479,N_24968);
nor UO_955 (O_955,N_24384,N_24545);
xnor UO_956 (O_956,N_24186,N_24690);
and UO_957 (O_957,N_24170,N_23756);
and UO_958 (O_958,N_24027,N_24212);
nor UO_959 (O_959,N_23916,N_24449);
or UO_960 (O_960,N_24495,N_24278);
and UO_961 (O_961,N_24261,N_24080);
and UO_962 (O_962,N_24243,N_24466);
and UO_963 (O_963,N_24621,N_24720);
or UO_964 (O_964,N_23824,N_24465);
nor UO_965 (O_965,N_24618,N_23867);
nand UO_966 (O_966,N_24309,N_24320);
nor UO_967 (O_967,N_24547,N_24608);
xnor UO_968 (O_968,N_24661,N_24039);
and UO_969 (O_969,N_24610,N_23767);
nor UO_970 (O_970,N_24299,N_23951);
or UO_971 (O_971,N_23914,N_24922);
nor UO_972 (O_972,N_23853,N_24865);
nand UO_973 (O_973,N_24052,N_24750);
xor UO_974 (O_974,N_24040,N_24140);
or UO_975 (O_975,N_24210,N_23860);
nor UO_976 (O_976,N_24379,N_24060);
nor UO_977 (O_977,N_24044,N_24476);
xnor UO_978 (O_978,N_24248,N_24718);
xnor UO_979 (O_979,N_23823,N_24464);
nand UO_980 (O_980,N_24418,N_24970);
nor UO_981 (O_981,N_24222,N_23831);
and UO_982 (O_982,N_24878,N_24885);
xnor UO_983 (O_983,N_24877,N_24805);
nor UO_984 (O_984,N_24056,N_24652);
nand UO_985 (O_985,N_23922,N_24863);
nor UO_986 (O_986,N_24281,N_24030);
nand UO_987 (O_987,N_23921,N_24795);
nand UO_988 (O_988,N_23954,N_24087);
xor UO_989 (O_989,N_23861,N_24746);
nor UO_990 (O_990,N_24986,N_24453);
nand UO_991 (O_991,N_23847,N_23765);
nand UO_992 (O_992,N_23905,N_24977);
or UO_993 (O_993,N_24450,N_23872);
nand UO_994 (O_994,N_23911,N_24162);
and UO_995 (O_995,N_24460,N_24380);
nor UO_996 (O_996,N_24317,N_23919);
nor UO_997 (O_997,N_24862,N_24622);
and UO_998 (O_998,N_24462,N_24303);
nand UO_999 (O_999,N_24157,N_24752);
nor UO_1000 (O_1000,N_24306,N_24709);
nor UO_1001 (O_1001,N_23776,N_24239);
nor UO_1002 (O_1002,N_24693,N_24591);
xor UO_1003 (O_1003,N_24700,N_24491);
nand UO_1004 (O_1004,N_24007,N_24201);
nand UO_1005 (O_1005,N_24013,N_23985);
xnor UO_1006 (O_1006,N_24686,N_23965);
and UO_1007 (O_1007,N_24089,N_24807);
or UO_1008 (O_1008,N_24742,N_24388);
or UO_1009 (O_1009,N_23936,N_24598);
xor UO_1010 (O_1010,N_24684,N_24552);
nor UO_1011 (O_1011,N_24742,N_24736);
xnor UO_1012 (O_1012,N_24655,N_23822);
and UO_1013 (O_1013,N_24559,N_24427);
and UO_1014 (O_1014,N_24045,N_24765);
or UO_1015 (O_1015,N_24953,N_23960);
nor UO_1016 (O_1016,N_24062,N_24142);
or UO_1017 (O_1017,N_24191,N_24507);
xnor UO_1018 (O_1018,N_23810,N_24707);
xor UO_1019 (O_1019,N_24903,N_24370);
and UO_1020 (O_1020,N_24299,N_24156);
xnor UO_1021 (O_1021,N_24030,N_24472);
nand UO_1022 (O_1022,N_24880,N_24719);
xor UO_1023 (O_1023,N_24159,N_24291);
xnor UO_1024 (O_1024,N_24146,N_24689);
xor UO_1025 (O_1025,N_24040,N_24413);
nor UO_1026 (O_1026,N_24284,N_24656);
xnor UO_1027 (O_1027,N_24018,N_24991);
or UO_1028 (O_1028,N_24568,N_24193);
and UO_1029 (O_1029,N_24194,N_24317);
xor UO_1030 (O_1030,N_23872,N_23762);
or UO_1031 (O_1031,N_24725,N_24227);
xnor UO_1032 (O_1032,N_24181,N_24139);
nand UO_1033 (O_1033,N_24456,N_23949);
and UO_1034 (O_1034,N_24177,N_23935);
xor UO_1035 (O_1035,N_24481,N_23972);
and UO_1036 (O_1036,N_24104,N_24065);
or UO_1037 (O_1037,N_24468,N_24089);
xor UO_1038 (O_1038,N_24326,N_24324);
and UO_1039 (O_1039,N_24001,N_24652);
or UO_1040 (O_1040,N_24763,N_24033);
or UO_1041 (O_1041,N_24332,N_24042);
and UO_1042 (O_1042,N_24511,N_24929);
nor UO_1043 (O_1043,N_24721,N_24612);
xor UO_1044 (O_1044,N_24791,N_24353);
nor UO_1045 (O_1045,N_24967,N_24789);
nand UO_1046 (O_1046,N_24407,N_23832);
or UO_1047 (O_1047,N_24630,N_23997);
and UO_1048 (O_1048,N_23878,N_24698);
or UO_1049 (O_1049,N_24340,N_24401);
nor UO_1050 (O_1050,N_24245,N_24797);
nor UO_1051 (O_1051,N_24104,N_24062);
and UO_1052 (O_1052,N_24556,N_24452);
xnor UO_1053 (O_1053,N_24755,N_23971);
or UO_1054 (O_1054,N_24772,N_24881);
nand UO_1055 (O_1055,N_24822,N_24423);
nand UO_1056 (O_1056,N_24479,N_23866);
or UO_1057 (O_1057,N_23980,N_23834);
xor UO_1058 (O_1058,N_24125,N_23807);
xnor UO_1059 (O_1059,N_24310,N_24915);
nand UO_1060 (O_1060,N_24100,N_24592);
nor UO_1061 (O_1061,N_24163,N_24485);
xor UO_1062 (O_1062,N_24963,N_24227);
or UO_1063 (O_1063,N_23803,N_24636);
or UO_1064 (O_1064,N_24760,N_24991);
nor UO_1065 (O_1065,N_24249,N_24154);
xnor UO_1066 (O_1066,N_24511,N_24321);
nand UO_1067 (O_1067,N_24886,N_24539);
and UO_1068 (O_1068,N_23848,N_23782);
xnor UO_1069 (O_1069,N_23792,N_24848);
and UO_1070 (O_1070,N_24713,N_24277);
xor UO_1071 (O_1071,N_23974,N_24974);
xor UO_1072 (O_1072,N_24748,N_24931);
or UO_1073 (O_1073,N_23915,N_24753);
and UO_1074 (O_1074,N_24411,N_23868);
and UO_1075 (O_1075,N_24032,N_24234);
and UO_1076 (O_1076,N_23933,N_24681);
xor UO_1077 (O_1077,N_24874,N_24442);
xnor UO_1078 (O_1078,N_24747,N_24470);
xor UO_1079 (O_1079,N_24704,N_24245);
or UO_1080 (O_1080,N_24098,N_23908);
nand UO_1081 (O_1081,N_24845,N_23954);
nor UO_1082 (O_1082,N_24097,N_24023);
and UO_1083 (O_1083,N_24478,N_24436);
and UO_1084 (O_1084,N_23899,N_24495);
or UO_1085 (O_1085,N_24063,N_24077);
nor UO_1086 (O_1086,N_24606,N_24917);
or UO_1087 (O_1087,N_24275,N_23908);
nand UO_1088 (O_1088,N_24686,N_24298);
and UO_1089 (O_1089,N_24092,N_24381);
nand UO_1090 (O_1090,N_24826,N_24909);
or UO_1091 (O_1091,N_24171,N_23904);
nor UO_1092 (O_1092,N_23783,N_23936);
nand UO_1093 (O_1093,N_24489,N_24090);
and UO_1094 (O_1094,N_24531,N_24556);
nor UO_1095 (O_1095,N_23993,N_24319);
xor UO_1096 (O_1096,N_23848,N_24177);
and UO_1097 (O_1097,N_24512,N_24832);
and UO_1098 (O_1098,N_24620,N_23868);
nand UO_1099 (O_1099,N_23872,N_24902);
nand UO_1100 (O_1100,N_23860,N_24640);
or UO_1101 (O_1101,N_24596,N_24088);
and UO_1102 (O_1102,N_23923,N_24972);
nand UO_1103 (O_1103,N_23835,N_24696);
nand UO_1104 (O_1104,N_24513,N_23806);
or UO_1105 (O_1105,N_24958,N_24606);
and UO_1106 (O_1106,N_24979,N_24083);
and UO_1107 (O_1107,N_23753,N_24138);
or UO_1108 (O_1108,N_23933,N_24036);
or UO_1109 (O_1109,N_24422,N_24758);
nand UO_1110 (O_1110,N_24715,N_24869);
nor UO_1111 (O_1111,N_24032,N_24089);
or UO_1112 (O_1112,N_24299,N_24119);
xnor UO_1113 (O_1113,N_24316,N_23935);
and UO_1114 (O_1114,N_23896,N_24770);
or UO_1115 (O_1115,N_23792,N_24029);
or UO_1116 (O_1116,N_23780,N_23897);
nor UO_1117 (O_1117,N_24265,N_24481);
xnor UO_1118 (O_1118,N_24808,N_24375);
or UO_1119 (O_1119,N_24799,N_24773);
and UO_1120 (O_1120,N_23993,N_24520);
nand UO_1121 (O_1121,N_23847,N_24622);
and UO_1122 (O_1122,N_24618,N_24241);
nand UO_1123 (O_1123,N_24713,N_24759);
or UO_1124 (O_1124,N_24433,N_24631);
or UO_1125 (O_1125,N_23967,N_24406);
or UO_1126 (O_1126,N_24476,N_23760);
xor UO_1127 (O_1127,N_24748,N_24195);
xor UO_1128 (O_1128,N_24631,N_24019);
nor UO_1129 (O_1129,N_23861,N_24589);
or UO_1130 (O_1130,N_24295,N_24731);
nor UO_1131 (O_1131,N_24027,N_23809);
nor UO_1132 (O_1132,N_23861,N_23987);
or UO_1133 (O_1133,N_23985,N_24318);
nor UO_1134 (O_1134,N_24314,N_24969);
nand UO_1135 (O_1135,N_24150,N_24710);
nor UO_1136 (O_1136,N_24983,N_23849);
nand UO_1137 (O_1137,N_24556,N_24701);
xor UO_1138 (O_1138,N_24748,N_24632);
xnor UO_1139 (O_1139,N_24442,N_24557);
and UO_1140 (O_1140,N_24167,N_24945);
xor UO_1141 (O_1141,N_24976,N_24914);
xor UO_1142 (O_1142,N_24716,N_24935);
or UO_1143 (O_1143,N_24867,N_24079);
nor UO_1144 (O_1144,N_24598,N_24836);
nand UO_1145 (O_1145,N_24687,N_24555);
or UO_1146 (O_1146,N_24811,N_24415);
or UO_1147 (O_1147,N_24373,N_24915);
xnor UO_1148 (O_1148,N_24719,N_24666);
nor UO_1149 (O_1149,N_24014,N_24840);
nor UO_1150 (O_1150,N_24530,N_24406);
and UO_1151 (O_1151,N_24597,N_24684);
nor UO_1152 (O_1152,N_24935,N_24363);
xnor UO_1153 (O_1153,N_24003,N_23863);
xnor UO_1154 (O_1154,N_24542,N_24956);
or UO_1155 (O_1155,N_24101,N_24442);
and UO_1156 (O_1156,N_23876,N_24446);
and UO_1157 (O_1157,N_23758,N_23753);
nor UO_1158 (O_1158,N_24568,N_24660);
nor UO_1159 (O_1159,N_24118,N_23960);
or UO_1160 (O_1160,N_24633,N_24912);
or UO_1161 (O_1161,N_23901,N_24293);
nand UO_1162 (O_1162,N_23789,N_23815);
and UO_1163 (O_1163,N_24205,N_23900);
xnor UO_1164 (O_1164,N_24141,N_24398);
nand UO_1165 (O_1165,N_24878,N_24109);
and UO_1166 (O_1166,N_24527,N_24239);
nand UO_1167 (O_1167,N_23900,N_23876);
and UO_1168 (O_1168,N_24061,N_24003);
xor UO_1169 (O_1169,N_24997,N_24769);
xnor UO_1170 (O_1170,N_23986,N_24158);
and UO_1171 (O_1171,N_24749,N_24016);
xor UO_1172 (O_1172,N_24431,N_24322);
xor UO_1173 (O_1173,N_24010,N_24459);
nand UO_1174 (O_1174,N_23995,N_23922);
nor UO_1175 (O_1175,N_24408,N_24592);
xor UO_1176 (O_1176,N_24083,N_24854);
nor UO_1177 (O_1177,N_24700,N_24997);
xor UO_1178 (O_1178,N_24768,N_23817);
nor UO_1179 (O_1179,N_24357,N_24846);
nor UO_1180 (O_1180,N_24290,N_24942);
nor UO_1181 (O_1181,N_24835,N_23843);
and UO_1182 (O_1182,N_24868,N_24763);
and UO_1183 (O_1183,N_24620,N_24444);
nand UO_1184 (O_1184,N_24743,N_24374);
or UO_1185 (O_1185,N_24756,N_24916);
nor UO_1186 (O_1186,N_24188,N_23807);
nor UO_1187 (O_1187,N_24740,N_24055);
nand UO_1188 (O_1188,N_24693,N_24386);
nor UO_1189 (O_1189,N_24835,N_24347);
or UO_1190 (O_1190,N_23792,N_24736);
nand UO_1191 (O_1191,N_24396,N_23775);
and UO_1192 (O_1192,N_23816,N_24209);
xor UO_1193 (O_1193,N_24745,N_24493);
or UO_1194 (O_1194,N_24052,N_23764);
nor UO_1195 (O_1195,N_24935,N_24792);
or UO_1196 (O_1196,N_24720,N_24045);
nand UO_1197 (O_1197,N_24845,N_24268);
or UO_1198 (O_1198,N_24033,N_24897);
or UO_1199 (O_1199,N_23876,N_24230);
nand UO_1200 (O_1200,N_23803,N_24905);
nor UO_1201 (O_1201,N_24056,N_24383);
and UO_1202 (O_1202,N_24373,N_24104);
xnor UO_1203 (O_1203,N_24567,N_24223);
nor UO_1204 (O_1204,N_24996,N_24400);
xor UO_1205 (O_1205,N_24316,N_23909);
and UO_1206 (O_1206,N_24413,N_24763);
xnor UO_1207 (O_1207,N_24817,N_24795);
or UO_1208 (O_1208,N_24486,N_23813);
and UO_1209 (O_1209,N_24528,N_24237);
nor UO_1210 (O_1210,N_24130,N_24690);
nor UO_1211 (O_1211,N_24021,N_24594);
nor UO_1212 (O_1212,N_24828,N_24022);
or UO_1213 (O_1213,N_24900,N_23930);
xnor UO_1214 (O_1214,N_24188,N_23820);
or UO_1215 (O_1215,N_24861,N_24831);
or UO_1216 (O_1216,N_24220,N_24824);
and UO_1217 (O_1217,N_24579,N_24673);
nor UO_1218 (O_1218,N_23750,N_23859);
nand UO_1219 (O_1219,N_24579,N_24948);
nor UO_1220 (O_1220,N_24094,N_24007);
and UO_1221 (O_1221,N_24389,N_24891);
or UO_1222 (O_1222,N_23906,N_24923);
nor UO_1223 (O_1223,N_24780,N_24666);
xor UO_1224 (O_1224,N_24454,N_23908);
nand UO_1225 (O_1225,N_24494,N_24840);
nand UO_1226 (O_1226,N_24257,N_24340);
nand UO_1227 (O_1227,N_24193,N_23840);
or UO_1228 (O_1228,N_24273,N_24835);
xnor UO_1229 (O_1229,N_23937,N_23916);
xor UO_1230 (O_1230,N_23762,N_24029);
nor UO_1231 (O_1231,N_24242,N_23871);
nor UO_1232 (O_1232,N_24186,N_24194);
or UO_1233 (O_1233,N_24341,N_24726);
and UO_1234 (O_1234,N_24153,N_24081);
and UO_1235 (O_1235,N_24726,N_24574);
xor UO_1236 (O_1236,N_24089,N_24404);
or UO_1237 (O_1237,N_24732,N_23957);
nor UO_1238 (O_1238,N_24544,N_23966);
or UO_1239 (O_1239,N_24639,N_24409);
or UO_1240 (O_1240,N_24171,N_24913);
nand UO_1241 (O_1241,N_24798,N_24991);
nand UO_1242 (O_1242,N_24083,N_23772);
and UO_1243 (O_1243,N_23754,N_24834);
and UO_1244 (O_1244,N_24160,N_24655);
nor UO_1245 (O_1245,N_24835,N_23912);
and UO_1246 (O_1246,N_24488,N_23819);
nor UO_1247 (O_1247,N_24337,N_24197);
or UO_1248 (O_1248,N_24029,N_24558);
or UO_1249 (O_1249,N_24727,N_24857);
and UO_1250 (O_1250,N_23920,N_24782);
nand UO_1251 (O_1251,N_24938,N_24764);
or UO_1252 (O_1252,N_24934,N_23876);
and UO_1253 (O_1253,N_23887,N_24538);
nand UO_1254 (O_1254,N_24852,N_24744);
xor UO_1255 (O_1255,N_23997,N_24031);
and UO_1256 (O_1256,N_24426,N_24879);
or UO_1257 (O_1257,N_24837,N_24357);
xor UO_1258 (O_1258,N_24417,N_24520);
xor UO_1259 (O_1259,N_24918,N_23925);
nand UO_1260 (O_1260,N_24908,N_23751);
and UO_1261 (O_1261,N_24008,N_24776);
xor UO_1262 (O_1262,N_24707,N_23946);
and UO_1263 (O_1263,N_24446,N_24448);
and UO_1264 (O_1264,N_24150,N_24049);
xnor UO_1265 (O_1265,N_24028,N_24208);
xnor UO_1266 (O_1266,N_24879,N_24754);
and UO_1267 (O_1267,N_24382,N_24746);
nor UO_1268 (O_1268,N_23824,N_24920);
nor UO_1269 (O_1269,N_24763,N_23915);
or UO_1270 (O_1270,N_24522,N_24557);
nor UO_1271 (O_1271,N_24452,N_24838);
nand UO_1272 (O_1272,N_24927,N_24513);
nand UO_1273 (O_1273,N_24588,N_24088);
nor UO_1274 (O_1274,N_24190,N_24059);
or UO_1275 (O_1275,N_24502,N_23770);
xor UO_1276 (O_1276,N_23871,N_23901);
or UO_1277 (O_1277,N_24705,N_23867);
or UO_1278 (O_1278,N_24104,N_24796);
xor UO_1279 (O_1279,N_23820,N_24493);
nand UO_1280 (O_1280,N_24877,N_23757);
nand UO_1281 (O_1281,N_24919,N_24499);
nand UO_1282 (O_1282,N_23809,N_23794);
xor UO_1283 (O_1283,N_23986,N_24261);
xor UO_1284 (O_1284,N_24329,N_24523);
xnor UO_1285 (O_1285,N_24144,N_24022);
nand UO_1286 (O_1286,N_23982,N_24185);
xnor UO_1287 (O_1287,N_24824,N_23940);
nor UO_1288 (O_1288,N_24500,N_24984);
or UO_1289 (O_1289,N_24728,N_24921);
xnor UO_1290 (O_1290,N_24198,N_24106);
nor UO_1291 (O_1291,N_24310,N_24690);
xnor UO_1292 (O_1292,N_24558,N_24384);
nand UO_1293 (O_1293,N_24677,N_24050);
and UO_1294 (O_1294,N_23771,N_24271);
nand UO_1295 (O_1295,N_24099,N_24133);
and UO_1296 (O_1296,N_24801,N_23828);
nand UO_1297 (O_1297,N_24717,N_23912);
and UO_1298 (O_1298,N_24289,N_24486);
or UO_1299 (O_1299,N_24904,N_24554);
nand UO_1300 (O_1300,N_23953,N_23751);
or UO_1301 (O_1301,N_24089,N_24388);
nand UO_1302 (O_1302,N_24214,N_24261);
nand UO_1303 (O_1303,N_24055,N_24461);
nor UO_1304 (O_1304,N_24905,N_24965);
nor UO_1305 (O_1305,N_23947,N_24908);
or UO_1306 (O_1306,N_23800,N_24030);
nand UO_1307 (O_1307,N_24539,N_24117);
xor UO_1308 (O_1308,N_24109,N_24176);
nor UO_1309 (O_1309,N_24360,N_23839);
or UO_1310 (O_1310,N_24938,N_23910);
or UO_1311 (O_1311,N_24976,N_24995);
or UO_1312 (O_1312,N_24908,N_24287);
nor UO_1313 (O_1313,N_24450,N_24832);
nor UO_1314 (O_1314,N_24175,N_23967);
or UO_1315 (O_1315,N_23948,N_24739);
xor UO_1316 (O_1316,N_24009,N_24159);
nand UO_1317 (O_1317,N_23992,N_24911);
or UO_1318 (O_1318,N_24282,N_23837);
nor UO_1319 (O_1319,N_24412,N_24368);
nand UO_1320 (O_1320,N_24435,N_24840);
nor UO_1321 (O_1321,N_24135,N_24854);
xor UO_1322 (O_1322,N_23762,N_24714);
and UO_1323 (O_1323,N_24368,N_24863);
or UO_1324 (O_1324,N_24711,N_24494);
or UO_1325 (O_1325,N_24625,N_24463);
xor UO_1326 (O_1326,N_24756,N_24677);
or UO_1327 (O_1327,N_24951,N_24532);
nand UO_1328 (O_1328,N_24849,N_24009);
nor UO_1329 (O_1329,N_24784,N_24755);
nand UO_1330 (O_1330,N_23773,N_24330);
xnor UO_1331 (O_1331,N_24321,N_24497);
and UO_1332 (O_1332,N_24388,N_23825);
or UO_1333 (O_1333,N_24629,N_24545);
nor UO_1334 (O_1334,N_24447,N_24789);
xnor UO_1335 (O_1335,N_24134,N_23960);
or UO_1336 (O_1336,N_24826,N_24321);
or UO_1337 (O_1337,N_24974,N_24901);
xor UO_1338 (O_1338,N_24147,N_24431);
nor UO_1339 (O_1339,N_24268,N_24837);
nor UO_1340 (O_1340,N_24336,N_24263);
nand UO_1341 (O_1341,N_23796,N_23826);
nand UO_1342 (O_1342,N_24620,N_24675);
or UO_1343 (O_1343,N_24664,N_24833);
or UO_1344 (O_1344,N_24561,N_24037);
and UO_1345 (O_1345,N_24038,N_24577);
or UO_1346 (O_1346,N_24844,N_23912);
nor UO_1347 (O_1347,N_24731,N_24523);
and UO_1348 (O_1348,N_24655,N_24470);
and UO_1349 (O_1349,N_23975,N_24470);
xnor UO_1350 (O_1350,N_24825,N_23803);
or UO_1351 (O_1351,N_24350,N_24566);
or UO_1352 (O_1352,N_24422,N_24279);
and UO_1353 (O_1353,N_23908,N_24446);
or UO_1354 (O_1354,N_24394,N_24380);
nand UO_1355 (O_1355,N_24782,N_24266);
xnor UO_1356 (O_1356,N_23962,N_24436);
and UO_1357 (O_1357,N_24246,N_24642);
nor UO_1358 (O_1358,N_24000,N_24645);
xor UO_1359 (O_1359,N_24269,N_24137);
and UO_1360 (O_1360,N_24101,N_24322);
or UO_1361 (O_1361,N_23920,N_24319);
nor UO_1362 (O_1362,N_24446,N_24020);
nand UO_1363 (O_1363,N_24474,N_23974);
or UO_1364 (O_1364,N_24372,N_23994);
or UO_1365 (O_1365,N_23927,N_24002);
nand UO_1366 (O_1366,N_24614,N_24508);
nor UO_1367 (O_1367,N_24278,N_24258);
xnor UO_1368 (O_1368,N_24771,N_23877);
nand UO_1369 (O_1369,N_24334,N_24455);
or UO_1370 (O_1370,N_23940,N_24174);
xor UO_1371 (O_1371,N_24001,N_24799);
and UO_1372 (O_1372,N_24504,N_24356);
and UO_1373 (O_1373,N_23917,N_24200);
xor UO_1374 (O_1374,N_24590,N_24244);
xnor UO_1375 (O_1375,N_24694,N_23972);
nor UO_1376 (O_1376,N_23877,N_24498);
nor UO_1377 (O_1377,N_24637,N_24845);
nand UO_1378 (O_1378,N_23780,N_24683);
or UO_1379 (O_1379,N_24200,N_23926);
nand UO_1380 (O_1380,N_24844,N_24049);
and UO_1381 (O_1381,N_24000,N_24524);
or UO_1382 (O_1382,N_24693,N_24801);
nand UO_1383 (O_1383,N_24810,N_24964);
or UO_1384 (O_1384,N_24962,N_24928);
xor UO_1385 (O_1385,N_24544,N_24190);
nand UO_1386 (O_1386,N_23940,N_24727);
xnor UO_1387 (O_1387,N_24469,N_23854);
xor UO_1388 (O_1388,N_24891,N_23814);
xnor UO_1389 (O_1389,N_24052,N_24323);
xor UO_1390 (O_1390,N_24219,N_23757);
or UO_1391 (O_1391,N_23966,N_24613);
xnor UO_1392 (O_1392,N_24671,N_23976);
and UO_1393 (O_1393,N_23951,N_23784);
nor UO_1394 (O_1394,N_24797,N_24590);
and UO_1395 (O_1395,N_24315,N_24464);
nand UO_1396 (O_1396,N_24987,N_23843);
nand UO_1397 (O_1397,N_23948,N_23810);
nor UO_1398 (O_1398,N_24881,N_24613);
nor UO_1399 (O_1399,N_23950,N_24059);
nand UO_1400 (O_1400,N_24496,N_24619);
and UO_1401 (O_1401,N_24557,N_24940);
nand UO_1402 (O_1402,N_24736,N_24050);
and UO_1403 (O_1403,N_23943,N_24802);
nand UO_1404 (O_1404,N_24898,N_24793);
and UO_1405 (O_1405,N_24694,N_24988);
xnor UO_1406 (O_1406,N_23898,N_23915);
and UO_1407 (O_1407,N_24315,N_24076);
nand UO_1408 (O_1408,N_23914,N_24572);
nor UO_1409 (O_1409,N_24754,N_24063);
nand UO_1410 (O_1410,N_24082,N_23979);
xor UO_1411 (O_1411,N_24803,N_24824);
xor UO_1412 (O_1412,N_23890,N_24662);
nand UO_1413 (O_1413,N_23795,N_24887);
xnor UO_1414 (O_1414,N_23761,N_24388);
xor UO_1415 (O_1415,N_24084,N_23771);
and UO_1416 (O_1416,N_24098,N_23847);
xor UO_1417 (O_1417,N_24275,N_23946);
or UO_1418 (O_1418,N_24598,N_24238);
xnor UO_1419 (O_1419,N_24137,N_23993);
xnor UO_1420 (O_1420,N_23786,N_24426);
xor UO_1421 (O_1421,N_24440,N_24347);
nand UO_1422 (O_1422,N_24355,N_23896);
nand UO_1423 (O_1423,N_24364,N_24500);
nand UO_1424 (O_1424,N_23881,N_24772);
and UO_1425 (O_1425,N_24039,N_23863);
and UO_1426 (O_1426,N_24253,N_24692);
and UO_1427 (O_1427,N_24425,N_24888);
nor UO_1428 (O_1428,N_24382,N_24722);
and UO_1429 (O_1429,N_24466,N_24290);
xnor UO_1430 (O_1430,N_24017,N_24040);
or UO_1431 (O_1431,N_24020,N_24631);
and UO_1432 (O_1432,N_23995,N_24408);
or UO_1433 (O_1433,N_24866,N_23806);
nand UO_1434 (O_1434,N_24194,N_24025);
or UO_1435 (O_1435,N_24381,N_24314);
nor UO_1436 (O_1436,N_24651,N_24974);
nand UO_1437 (O_1437,N_24304,N_24760);
nor UO_1438 (O_1438,N_24885,N_24054);
nor UO_1439 (O_1439,N_24362,N_24899);
xor UO_1440 (O_1440,N_23837,N_24210);
and UO_1441 (O_1441,N_23946,N_24146);
nor UO_1442 (O_1442,N_24746,N_24665);
and UO_1443 (O_1443,N_24099,N_24629);
nor UO_1444 (O_1444,N_23765,N_24201);
xnor UO_1445 (O_1445,N_23788,N_24689);
or UO_1446 (O_1446,N_24572,N_24878);
nor UO_1447 (O_1447,N_23889,N_24254);
xnor UO_1448 (O_1448,N_24945,N_23872);
and UO_1449 (O_1449,N_24927,N_24505);
or UO_1450 (O_1450,N_24318,N_24506);
or UO_1451 (O_1451,N_23994,N_24439);
xor UO_1452 (O_1452,N_24595,N_24586);
nor UO_1453 (O_1453,N_23967,N_23782);
nand UO_1454 (O_1454,N_24460,N_24396);
and UO_1455 (O_1455,N_24679,N_24794);
xnor UO_1456 (O_1456,N_24251,N_23812);
nand UO_1457 (O_1457,N_24452,N_23754);
and UO_1458 (O_1458,N_24565,N_24654);
nand UO_1459 (O_1459,N_23764,N_24696);
nand UO_1460 (O_1460,N_24171,N_24121);
nor UO_1461 (O_1461,N_24367,N_24071);
xnor UO_1462 (O_1462,N_24783,N_24486);
nor UO_1463 (O_1463,N_23806,N_23977);
xor UO_1464 (O_1464,N_24431,N_24878);
nand UO_1465 (O_1465,N_24572,N_24765);
or UO_1466 (O_1466,N_24453,N_24029);
nor UO_1467 (O_1467,N_24120,N_24411);
nor UO_1468 (O_1468,N_24194,N_24326);
or UO_1469 (O_1469,N_24780,N_24822);
xor UO_1470 (O_1470,N_24631,N_24272);
and UO_1471 (O_1471,N_24567,N_24741);
xor UO_1472 (O_1472,N_24278,N_24288);
and UO_1473 (O_1473,N_24350,N_24596);
nor UO_1474 (O_1474,N_24849,N_24395);
or UO_1475 (O_1475,N_24531,N_23900);
nand UO_1476 (O_1476,N_24715,N_24849);
nand UO_1477 (O_1477,N_24261,N_24700);
and UO_1478 (O_1478,N_23807,N_23971);
or UO_1479 (O_1479,N_24459,N_24609);
nand UO_1480 (O_1480,N_24909,N_24142);
xnor UO_1481 (O_1481,N_24006,N_24265);
nor UO_1482 (O_1482,N_24789,N_24774);
nand UO_1483 (O_1483,N_24923,N_24718);
xor UO_1484 (O_1484,N_24975,N_24029);
nand UO_1485 (O_1485,N_24284,N_24388);
nand UO_1486 (O_1486,N_23868,N_24787);
or UO_1487 (O_1487,N_23937,N_24223);
and UO_1488 (O_1488,N_24590,N_24959);
and UO_1489 (O_1489,N_24727,N_23889);
and UO_1490 (O_1490,N_24597,N_24607);
or UO_1491 (O_1491,N_23841,N_24771);
nand UO_1492 (O_1492,N_23995,N_24676);
and UO_1493 (O_1493,N_23845,N_24662);
and UO_1494 (O_1494,N_24442,N_23864);
xor UO_1495 (O_1495,N_24435,N_24471);
or UO_1496 (O_1496,N_24824,N_23924);
nand UO_1497 (O_1497,N_24337,N_24356);
and UO_1498 (O_1498,N_24122,N_24189);
or UO_1499 (O_1499,N_24438,N_23941);
and UO_1500 (O_1500,N_23872,N_24940);
xnor UO_1501 (O_1501,N_24847,N_24526);
xor UO_1502 (O_1502,N_24815,N_23915);
nor UO_1503 (O_1503,N_23866,N_24420);
nand UO_1504 (O_1504,N_23755,N_24165);
nand UO_1505 (O_1505,N_24090,N_24777);
nor UO_1506 (O_1506,N_23884,N_24314);
and UO_1507 (O_1507,N_24339,N_24158);
or UO_1508 (O_1508,N_24956,N_24623);
nand UO_1509 (O_1509,N_24683,N_24232);
nor UO_1510 (O_1510,N_24301,N_24552);
nand UO_1511 (O_1511,N_24510,N_23768);
xnor UO_1512 (O_1512,N_24378,N_24492);
xnor UO_1513 (O_1513,N_24595,N_24842);
nor UO_1514 (O_1514,N_24349,N_24738);
xor UO_1515 (O_1515,N_24435,N_24269);
nor UO_1516 (O_1516,N_24177,N_24996);
or UO_1517 (O_1517,N_23846,N_24558);
and UO_1518 (O_1518,N_24907,N_24556);
xor UO_1519 (O_1519,N_24529,N_24442);
nor UO_1520 (O_1520,N_24152,N_24378);
and UO_1521 (O_1521,N_24940,N_24430);
nand UO_1522 (O_1522,N_24958,N_24916);
xnor UO_1523 (O_1523,N_24134,N_24910);
and UO_1524 (O_1524,N_24356,N_24730);
and UO_1525 (O_1525,N_24975,N_24719);
nor UO_1526 (O_1526,N_24411,N_24064);
or UO_1527 (O_1527,N_24865,N_24275);
nand UO_1528 (O_1528,N_24997,N_24295);
and UO_1529 (O_1529,N_23887,N_24363);
nor UO_1530 (O_1530,N_24633,N_24874);
and UO_1531 (O_1531,N_23810,N_24893);
and UO_1532 (O_1532,N_24732,N_24502);
or UO_1533 (O_1533,N_24432,N_23823);
xnor UO_1534 (O_1534,N_24757,N_24952);
or UO_1535 (O_1535,N_24830,N_24946);
and UO_1536 (O_1536,N_24259,N_24365);
nor UO_1537 (O_1537,N_23965,N_24038);
and UO_1538 (O_1538,N_24603,N_24267);
nand UO_1539 (O_1539,N_24019,N_23823);
or UO_1540 (O_1540,N_24835,N_23973);
and UO_1541 (O_1541,N_24248,N_24570);
xor UO_1542 (O_1542,N_24334,N_24773);
nand UO_1543 (O_1543,N_24286,N_24214);
xnor UO_1544 (O_1544,N_24897,N_24603);
nor UO_1545 (O_1545,N_24030,N_24165);
nor UO_1546 (O_1546,N_24479,N_24218);
nor UO_1547 (O_1547,N_23793,N_24593);
nand UO_1548 (O_1548,N_24035,N_23796);
and UO_1549 (O_1549,N_23943,N_24297);
xor UO_1550 (O_1550,N_24097,N_24525);
nor UO_1551 (O_1551,N_24235,N_24795);
or UO_1552 (O_1552,N_24017,N_24016);
and UO_1553 (O_1553,N_23985,N_24868);
and UO_1554 (O_1554,N_24434,N_24136);
nand UO_1555 (O_1555,N_24728,N_24314);
and UO_1556 (O_1556,N_24896,N_24679);
nor UO_1557 (O_1557,N_24007,N_23907);
and UO_1558 (O_1558,N_24821,N_24151);
or UO_1559 (O_1559,N_24397,N_24880);
nor UO_1560 (O_1560,N_23857,N_24724);
xnor UO_1561 (O_1561,N_24171,N_24079);
nor UO_1562 (O_1562,N_24111,N_24311);
nor UO_1563 (O_1563,N_23995,N_24271);
and UO_1564 (O_1564,N_24622,N_24092);
nand UO_1565 (O_1565,N_24859,N_24897);
nand UO_1566 (O_1566,N_24318,N_23864);
nand UO_1567 (O_1567,N_24733,N_24655);
and UO_1568 (O_1568,N_24567,N_24155);
or UO_1569 (O_1569,N_23909,N_24476);
nor UO_1570 (O_1570,N_24970,N_24774);
and UO_1571 (O_1571,N_24647,N_23908);
and UO_1572 (O_1572,N_24161,N_24986);
nand UO_1573 (O_1573,N_24252,N_24850);
and UO_1574 (O_1574,N_23868,N_24868);
xor UO_1575 (O_1575,N_24273,N_24456);
and UO_1576 (O_1576,N_23895,N_24951);
nand UO_1577 (O_1577,N_24794,N_24435);
or UO_1578 (O_1578,N_24333,N_23826);
or UO_1579 (O_1579,N_24952,N_24059);
nand UO_1580 (O_1580,N_23887,N_24895);
and UO_1581 (O_1581,N_24650,N_24986);
nor UO_1582 (O_1582,N_24214,N_24440);
xnor UO_1583 (O_1583,N_24236,N_24270);
and UO_1584 (O_1584,N_23778,N_24286);
nand UO_1585 (O_1585,N_24239,N_23759);
and UO_1586 (O_1586,N_24731,N_24080);
nand UO_1587 (O_1587,N_24391,N_24971);
and UO_1588 (O_1588,N_24971,N_23986);
and UO_1589 (O_1589,N_24947,N_24849);
and UO_1590 (O_1590,N_24167,N_23774);
nor UO_1591 (O_1591,N_24070,N_23783);
and UO_1592 (O_1592,N_24475,N_23920);
nor UO_1593 (O_1593,N_24851,N_24977);
nor UO_1594 (O_1594,N_24184,N_24798);
nand UO_1595 (O_1595,N_24031,N_24867);
or UO_1596 (O_1596,N_24105,N_24035);
xnor UO_1597 (O_1597,N_24054,N_24538);
and UO_1598 (O_1598,N_23994,N_24649);
xnor UO_1599 (O_1599,N_24261,N_24331);
nand UO_1600 (O_1600,N_24398,N_24467);
nor UO_1601 (O_1601,N_23751,N_24570);
nor UO_1602 (O_1602,N_24324,N_24180);
nand UO_1603 (O_1603,N_23878,N_23836);
nand UO_1604 (O_1604,N_23848,N_24508);
and UO_1605 (O_1605,N_24534,N_24150);
nor UO_1606 (O_1606,N_24949,N_24169);
or UO_1607 (O_1607,N_24510,N_24271);
nor UO_1608 (O_1608,N_23787,N_23812);
and UO_1609 (O_1609,N_24027,N_24608);
nor UO_1610 (O_1610,N_24741,N_23759);
nand UO_1611 (O_1611,N_24492,N_24972);
and UO_1612 (O_1612,N_24935,N_24676);
or UO_1613 (O_1613,N_24339,N_24924);
xor UO_1614 (O_1614,N_24675,N_24563);
nor UO_1615 (O_1615,N_24304,N_24632);
xor UO_1616 (O_1616,N_24051,N_24034);
xnor UO_1617 (O_1617,N_24951,N_24618);
xor UO_1618 (O_1618,N_23826,N_23786);
nor UO_1619 (O_1619,N_24767,N_24497);
xnor UO_1620 (O_1620,N_23805,N_23777);
nand UO_1621 (O_1621,N_24953,N_24023);
or UO_1622 (O_1622,N_24585,N_23986);
and UO_1623 (O_1623,N_23755,N_24546);
nor UO_1624 (O_1624,N_23981,N_24896);
xnor UO_1625 (O_1625,N_24492,N_24464);
or UO_1626 (O_1626,N_24722,N_24631);
nor UO_1627 (O_1627,N_24074,N_24033);
and UO_1628 (O_1628,N_24474,N_24867);
xnor UO_1629 (O_1629,N_24863,N_24225);
nand UO_1630 (O_1630,N_24264,N_24173);
xnor UO_1631 (O_1631,N_24480,N_24114);
and UO_1632 (O_1632,N_24493,N_23834);
nand UO_1633 (O_1633,N_24170,N_24186);
xor UO_1634 (O_1634,N_24558,N_24934);
nand UO_1635 (O_1635,N_24850,N_24897);
or UO_1636 (O_1636,N_23922,N_24538);
or UO_1637 (O_1637,N_23848,N_23924);
or UO_1638 (O_1638,N_24797,N_24074);
nand UO_1639 (O_1639,N_24883,N_24738);
xor UO_1640 (O_1640,N_24167,N_24116);
and UO_1641 (O_1641,N_23887,N_23820);
nand UO_1642 (O_1642,N_24832,N_24501);
xnor UO_1643 (O_1643,N_24991,N_24393);
and UO_1644 (O_1644,N_24395,N_24839);
xor UO_1645 (O_1645,N_24234,N_23921);
or UO_1646 (O_1646,N_24059,N_24462);
or UO_1647 (O_1647,N_23796,N_24051);
nand UO_1648 (O_1648,N_24227,N_23957);
and UO_1649 (O_1649,N_24219,N_24747);
nand UO_1650 (O_1650,N_24094,N_23895);
nor UO_1651 (O_1651,N_24954,N_24553);
and UO_1652 (O_1652,N_24180,N_24622);
and UO_1653 (O_1653,N_24830,N_24715);
nand UO_1654 (O_1654,N_23821,N_24189);
xor UO_1655 (O_1655,N_23807,N_24012);
or UO_1656 (O_1656,N_23785,N_23943);
or UO_1657 (O_1657,N_23998,N_24386);
or UO_1658 (O_1658,N_23845,N_24303);
and UO_1659 (O_1659,N_23936,N_24138);
xor UO_1660 (O_1660,N_24426,N_24066);
and UO_1661 (O_1661,N_24714,N_24887);
and UO_1662 (O_1662,N_24586,N_24133);
or UO_1663 (O_1663,N_24910,N_24051);
xor UO_1664 (O_1664,N_24297,N_24232);
nor UO_1665 (O_1665,N_24306,N_24222);
or UO_1666 (O_1666,N_24537,N_24602);
nand UO_1667 (O_1667,N_24801,N_24982);
nor UO_1668 (O_1668,N_24288,N_24800);
nor UO_1669 (O_1669,N_24912,N_24703);
nand UO_1670 (O_1670,N_23925,N_24789);
nand UO_1671 (O_1671,N_24939,N_24249);
or UO_1672 (O_1672,N_24265,N_24355);
and UO_1673 (O_1673,N_24510,N_24358);
xnor UO_1674 (O_1674,N_24770,N_24079);
and UO_1675 (O_1675,N_24460,N_24704);
and UO_1676 (O_1676,N_24493,N_23758);
nand UO_1677 (O_1677,N_23851,N_24521);
and UO_1678 (O_1678,N_23815,N_23934);
and UO_1679 (O_1679,N_24192,N_24234);
and UO_1680 (O_1680,N_24262,N_24336);
nand UO_1681 (O_1681,N_24262,N_24083);
or UO_1682 (O_1682,N_24339,N_24181);
nor UO_1683 (O_1683,N_24195,N_24355);
nor UO_1684 (O_1684,N_24319,N_24942);
nor UO_1685 (O_1685,N_23753,N_24347);
xnor UO_1686 (O_1686,N_23954,N_24147);
nor UO_1687 (O_1687,N_24984,N_24808);
nand UO_1688 (O_1688,N_24691,N_24867);
or UO_1689 (O_1689,N_24033,N_24101);
or UO_1690 (O_1690,N_24206,N_23942);
or UO_1691 (O_1691,N_24476,N_24739);
nand UO_1692 (O_1692,N_24413,N_23822);
xor UO_1693 (O_1693,N_23867,N_24830);
xor UO_1694 (O_1694,N_24493,N_24927);
or UO_1695 (O_1695,N_24032,N_24829);
xnor UO_1696 (O_1696,N_24909,N_24076);
nand UO_1697 (O_1697,N_23958,N_24766);
nand UO_1698 (O_1698,N_24969,N_24468);
nand UO_1699 (O_1699,N_23917,N_24261);
nor UO_1700 (O_1700,N_23850,N_24845);
nor UO_1701 (O_1701,N_24429,N_24336);
nor UO_1702 (O_1702,N_23944,N_24290);
or UO_1703 (O_1703,N_24957,N_24192);
nand UO_1704 (O_1704,N_24374,N_24292);
and UO_1705 (O_1705,N_23807,N_24986);
and UO_1706 (O_1706,N_24410,N_23850);
and UO_1707 (O_1707,N_24834,N_24311);
and UO_1708 (O_1708,N_24873,N_24491);
and UO_1709 (O_1709,N_24992,N_24515);
and UO_1710 (O_1710,N_24436,N_24571);
and UO_1711 (O_1711,N_24355,N_24296);
nand UO_1712 (O_1712,N_23863,N_24246);
nand UO_1713 (O_1713,N_24227,N_24498);
and UO_1714 (O_1714,N_24864,N_24170);
or UO_1715 (O_1715,N_24430,N_23827);
nand UO_1716 (O_1716,N_24817,N_23774);
nand UO_1717 (O_1717,N_24665,N_24769);
xnor UO_1718 (O_1718,N_23829,N_24793);
xnor UO_1719 (O_1719,N_24265,N_24905);
xor UO_1720 (O_1720,N_24962,N_23921);
or UO_1721 (O_1721,N_23944,N_24941);
or UO_1722 (O_1722,N_23963,N_24480);
nor UO_1723 (O_1723,N_24214,N_24289);
nand UO_1724 (O_1724,N_24241,N_24033);
nor UO_1725 (O_1725,N_24635,N_24142);
nand UO_1726 (O_1726,N_24725,N_24665);
nor UO_1727 (O_1727,N_24166,N_23856);
and UO_1728 (O_1728,N_24759,N_23803);
nand UO_1729 (O_1729,N_24478,N_24970);
nand UO_1730 (O_1730,N_24953,N_24532);
nand UO_1731 (O_1731,N_23933,N_24770);
and UO_1732 (O_1732,N_24333,N_24311);
and UO_1733 (O_1733,N_24029,N_24032);
and UO_1734 (O_1734,N_24681,N_24579);
nor UO_1735 (O_1735,N_24334,N_23803);
nand UO_1736 (O_1736,N_23921,N_24853);
nor UO_1737 (O_1737,N_24243,N_24632);
and UO_1738 (O_1738,N_24025,N_24901);
nor UO_1739 (O_1739,N_23848,N_24890);
and UO_1740 (O_1740,N_24221,N_24002);
xnor UO_1741 (O_1741,N_24525,N_24408);
xnor UO_1742 (O_1742,N_24090,N_24723);
nor UO_1743 (O_1743,N_24555,N_23916);
or UO_1744 (O_1744,N_24644,N_24158);
nor UO_1745 (O_1745,N_24933,N_24803);
nor UO_1746 (O_1746,N_24657,N_24954);
xor UO_1747 (O_1747,N_24562,N_23998);
nor UO_1748 (O_1748,N_24251,N_23887);
nor UO_1749 (O_1749,N_24661,N_24288);
and UO_1750 (O_1750,N_24199,N_24510);
nor UO_1751 (O_1751,N_24577,N_23785);
xnor UO_1752 (O_1752,N_24937,N_24135);
xor UO_1753 (O_1753,N_24364,N_23763);
xor UO_1754 (O_1754,N_24711,N_24201);
or UO_1755 (O_1755,N_24882,N_23961);
xnor UO_1756 (O_1756,N_24489,N_23974);
xor UO_1757 (O_1757,N_23809,N_23926);
xnor UO_1758 (O_1758,N_23920,N_24894);
or UO_1759 (O_1759,N_24603,N_24783);
nand UO_1760 (O_1760,N_24426,N_24212);
nand UO_1761 (O_1761,N_24996,N_24071);
and UO_1762 (O_1762,N_24011,N_24749);
nor UO_1763 (O_1763,N_24912,N_23989);
or UO_1764 (O_1764,N_24417,N_24513);
nand UO_1765 (O_1765,N_24955,N_24492);
and UO_1766 (O_1766,N_23815,N_23856);
nand UO_1767 (O_1767,N_24940,N_24622);
xor UO_1768 (O_1768,N_24412,N_24148);
or UO_1769 (O_1769,N_24940,N_24388);
nand UO_1770 (O_1770,N_24284,N_24340);
and UO_1771 (O_1771,N_23803,N_24422);
xnor UO_1772 (O_1772,N_24512,N_24069);
nand UO_1773 (O_1773,N_24726,N_24048);
nand UO_1774 (O_1774,N_24702,N_23929);
nand UO_1775 (O_1775,N_24799,N_24181);
xor UO_1776 (O_1776,N_24617,N_24203);
or UO_1777 (O_1777,N_24665,N_23935);
nor UO_1778 (O_1778,N_23958,N_24402);
xnor UO_1779 (O_1779,N_24588,N_24162);
xor UO_1780 (O_1780,N_24431,N_23833);
nand UO_1781 (O_1781,N_24739,N_24897);
or UO_1782 (O_1782,N_24250,N_24892);
and UO_1783 (O_1783,N_24705,N_24662);
xor UO_1784 (O_1784,N_24465,N_24422);
xnor UO_1785 (O_1785,N_24442,N_24173);
or UO_1786 (O_1786,N_23938,N_24250);
nand UO_1787 (O_1787,N_24977,N_24757);
nor UO_1788 (O_1788,N_24471,N_24260);
xnor UO_1789 (O_1789,N_24629,N_24506);
nor UO_1790 (O_1790,N_23767,N_24281);
nor UO_1791 (O_1791,N_24274,N_24339);
and UO_1792 (O_1792,N_24221,N_24679);
or UO_1793 (O_1793,N_24939,N_24994);
nand UO_1794 (O_1794,N_23919,N_24933);
and UO_1795 (O_1795,N_24537,N_24343);
nor UO_1796 (O_1796,N_23980,N_24217);
xor UO_1797 (O_1797,N_24226,N_24727);
or UO_1798 (O_1798,N_23899,N_24815);
or UO_1799 (O_1799,N_24362,N_24652);
nor UO_1800 (O_1800,N_24466,N_24470);
nand UO_1801 (O_1801,N_24788,N_24266);
nand UO_1802 (O_1802,N_24278,N_24624);
and UO_1803 (O_1803,N_24087,N_24254);
nor UO_1804 (O_1804,N_24781,N_24838);
and UO_1805 (O_1805,N_24964,N_23921);
or UO_1806 (O_1806,N_23784,N_24653);
nor UO_1807 (O_1807,N_24161,N_24296);
nand UO_1808 (O_1808,N_24544,N_24572);
xor UO_1809 (O_1809,N_23900,N_24982);
xor UO_1810 (O_1810,N_24379,N_24233);
nor UO_1811 (O_1811,N_24136,N_24725);
xnor UO_1812 (O_1812,N_24565,N_23879);
and UO_1813 (O_1813,N_24919,N_24273);
or UO_1814 (O_1814,N_24965,N_24859);
and UO_1815 (O_1815,N_23831,N_24601);
nand UO_1816 (O_1816,N_23810,N_23828);
and UO_1817 (O_1817,N_24150,N_23960);
nor UO_1818 (O_1818,N_24580,N_24260);
or UO_1819 (O_1819,N_24853,N_24649);
or UO_1820 (O_1820,N_24010,N_23925);
or UO_1821 (O_1821,N_24830,N_24661);
nand UO_1822 (O_1822,N_24531,N_24468);
and UO_1823 (O_1823,N_23762,N_24484);
or UO_1824 (O_1824,N_24801,N_24354);
nor UO_1825 (O_1825,N_24155,N_24948);
xor UO_1826 (O_1826,N_24101,N_23915);
or UO_1827 (O_1827,N_23982,N_23767);
and UO_1828 (O_1828,N_24113,N_23930);
nand UO_1829 (O_1829,N_24149,N_24654);
nor UO_1830 (O_1830,N_24714,N_24856);
nand UO_1831 (O_1831,N_24553,N_24251);
or UO_1832 (O_1832,N_24297,N_24671);
xor UO_1833 (O_1833,N_23791,N_24582);
nor UO_1834 (O_1834,N_24561,N_24990);
xor UO_1835 (O_1835,N_24750,N_24935);
and UO_1836 (O_1836,N_24026,N_24991);
nor UO_1837 (O_1837,N_24145,N_24407);
and UO_1838 (O_1838,N_24769,N_24798);
nor UO_1839 (O_1839,N_24365,N_24465);
or UO_1840 (O_1840,N_23943,N_24584);
and UO_1841 (O_1841,N_24003,N_24629);
nand UO_1842 (O_1842,N_24298,N_23955);
nand UO_1843 (O_1843,N_24872,N_24128);
and UO_1844 (O_1844,N_24284,N_24911);
nor UO_1845 (O_1845,N_24856,N_24402);
or UO_1846 (O_1846,N_24159,N_24121);
and UO_1847 (O_1847,N_24928,N_24106);
or UO_1848 (O_1848,N_24014,N_24194);
and UO_1849 (O_1849,N_24312,N_24953);
and UO_1850 (O_1850,N_24884,N_24752);
nor UO_1851 (O_1851,N_24985,N_24292);
and UO_1852 (O_1852,N_24053,N_24075);
nor UO_1853 (O_1853,N_24979,N_23948);
nand UO_1854 (O_1854,N_24888,N_24590);
and UO_1855 (O_1855,N_24400,N_24554);
nand UO_1856 (O_1856,N_24234,N_24373);
or UO_1857 (O_1857,N_24780,N_23976);
nor UO_1858 (O_1858,N_24024,N_24506);
and UO_1859 (O_1859,N_24234,N_24408);
nor UO_1860 (O_1860,N_24382,N_24914);
and UO_1861 (O_1861,N_23931,N_24587);
or UO_1862 (O_1862,N_23767,N_24661);
and UO_1863 (O_1863,N_23905,N_24512);
and UO_1864 (O_1864,N_24352,N_24628);
xnor UO_1865 (O_1865,N_23805,N_23793);
xnor UO_1866 (O_1866,N_24538,N_24277);
nand UO_1867 (O_1867,N_24800,N_24883);
or UO_1868 (O_1868,N_24173,N_23950);
and UO_1869 (O_1869,N_24808,N_24649);
or UO_1870 (O_1870,N_24642,N_24801);
nor UO_1871 (O_1871,N_24951,N_24759);
and UO_1872 (O_1872,N_24703,N_24613);
xor UO_1873 (O_1873,N_24659,N_23911);
and UO_1874 (O_1874,N_24593,N_24976);
xor UO_1875 (O_1875,N_24953,N_24696);
nor UO_1876 (O_1876,N_24609,N_24566);
or UO_1877 (O_1877,N_24160,N_24600);
or UO_1878 (O_1878,N_23937,N_24259);
xor UO_1879 (O_1879,N_23938,N_23859);
or UO_1880 (O_1880,N_24892,N_24577);
or UO_1881 (O_1881,N_24818,N_24593);
xnor UO_1882 (O_1882,N_24479,N_23896);
or UO_1883 (O_1883,N_24619,N_24385);
nand UO_1884 (O_1884,N_24922,N_24728);
xnor UO_1885 (O_1885,N_23970,N_24502);
nand UO_1886 (O_1886,N_24579,N_24263);
nor UO_1887 (O_1887,N_24706,N_24660);
or UO_1888 (O_1888,N_24670,N_24045);
and UO_1889 (O_1889,N_24245,N_24078);
nand UO_1890 (O_1890,N_24329,N_24988);
and UO_1891 (O_1891,N_24532,N_24735);
or UO_1892 (O_1892,N_24877,N_24911);
nor UO_1893 (O_1893,N_24580,N_24472);
xor UO_1894 (O_1894,N_24856,N_23925);
and UO_1895 (O_1895,N_24361,N_24444);
or UO_1896 (O_1896,N_24205,N_24971);
or UO_1897 (O_1897,N_23813,N_24189);
and UO_1898 (O_1898,N_24059,N_24052);
nand UO_1899 (O_1899,N_23782,N_24691);
xnor UO_1900 (O_1900,N_24442,N_24542);
nor UO_1901 (O_1901,N_23905,N_24306);
nand UO_1902 (O_1902,N_24890,N_23948);
and UO_1903 (O_1903,N_24628,N_23890);
nand UO_1904 (O_1904,N_23818,N_23928);
nand UO_1905 (O_1905,N_23915,N_24861);
and UO_1906 (O_1906,N_24767,N_24424);
and UO_1907 (O_1907,N_24558,N_24449);
nand UO_1908 (O_1908,N_24935,N_24346);
xor UO_1909 (O_1909,N_24957,N_23985);
nor UO_1910 (O_1910,N_24238,N_24153);
nand UO_1911 (O_1911,N_24253,N_24395);
and UO_1912 (O_1912,N_24972,N_23877);
and UO_1913 (O_1913,N_24466,N_24703);
xor UO_1914 (O_1914,N_24322,N_24246);
or UO_1915 (O_1915,N_24261,N_23791);
nand UO_1916 (O_1916,N_24949,N_24260);
xor UO_1917 (O_1917,N_24000,N_24977);
or UO_1918 (O_1918,N_24807,N_24013);
xor UO_1919 (O_1919,N_24775,N_23842);
or UO_1920 (O_1920,N_24968,N_24820);
nand UO_1921 (O_1921,N_23910,N_24237);
or UO_1922 (O_1922,N_24296,N_24802);
and UO_1923 (O_1923,N_24231,N_24923);
or UO_1924 (O_1924,N_24355,N_24224);
nand UO_1925 (O_1925,N_24397,N_24456);
nor UO_1926 (O_1926,N_24215,N_23898);
nand UO_1927 (O_1927,N_23938,N_24012);
nor UO_1928 (O_1928,N_23855,N_23881);
or UO_1929 (O_1929,N_24342,N_23893);
or UO_1930 (O_1930,N_24434,N_24575);
and UO_1931 (O_1931,N_24116,N_24969);
or UO_1932 (O_1932,N_24651,N_23823);
nor UO_1933 (O_1933,N_23823,N_24799);
or UO_1934 (O_1934,N_24393,N_24415);
xor UO_1935 (O_1935,N_24343,N_24574);
or UO_1936 (O_1936,N_24578,N_24872);
nor UO_1937 (O_1937,N_24640,N_24648);
xor UO_1938 (O_1938,N_24881,N_24237);
nor UO_1939 (O_1939,N_24893,N_24430);
nand UO_1940 (O_1940,N_24858,N_24708);
nand UO_1941 (O_1941,N_24877,N_24459);
nor UO_1942 (O_1942,N_23978,N_24856);
or UO_1943 (O_1943,N_23920,N_24271);
or UO_1944 (O_1944,N_24355,N_23787);
and UO_1945 (O_1945,N_24157,N_24089);
nor UO_1946 (O_1946,N_24044,N_24956);
nor UO_1947 (O_1947,N_24803,N_24148);
or UO_1948 (O_1948,N_24426,N_24307);
xor UO_1949 (O_1949,N_24491,N_24480);
nand UO_1950 (O_1950,N_23804,N_24064);
or UO_1951 (O_1951,N_24100,N_24529);
xnor UO_1952 (O_1952,N_24946,N_24110);
xor UO_1953 (O_1953,N_24398,N_24943);
nand UO_1954 (O_1954,N_24687,N_24202);
xnor UO_1955 (O_1955,N_24029,N_24867);
xnor UO_1956 (O_1956,N_24331,N_24051);
nand UO_1957 (O_1957,N_24722,N_23875);
or UO_1958 (O_1958,N_24106,N_23990);
nand UO_1959 (O_1959,N_24097,N_24748);
or UO_1960 (O_1960,N_24065,N_24806);
nor UO_1961 (O_1961,N_24327,N_24733);
nor UO_1962 (O_1962,N_24933,N_24210);
xor UO_1963 (O_1963,N_24683,N_23846);
nor UO_1964 (O_1964,N_23925,N_24991);
or UO_1965 (O_1965,N_23979,N_24258);
nand UO_1966 (O_1966,N_24610,N_24015);
nand UO_1967 (O_1967,N_23948,N_24291);
and UO_1968 (O_1968,N_24370,N_24604);
nor UO_1969 (O_1969,N_23752,N_24489);
or UO_1970 (O_1970,N_24240,N_24763);
nor UO_1971 (O_1971,N_24499,N_23848);
and UO_1972 (O_1972,N_24093,N_24752);
and UO_1973 (O_1973,N_24398,N_24171);
nor UO_1974 (O_1974,N_23754,N_24364);
nand UO_1975 (O_1975,N_24380,N_23837);
or UO_1976 (O_1976,N_24954,N_24206);
nor UO_1977 (O_1977,N_24545,N_24572);
nor UO_1978 (O_1978,N_24519,N_23924);
nand UO_1979 (O_1979,N_24642,N_24517);
nand UO_1980 (O_1980,N_24726,N_24633);
nor UO_1981 (O_1981,N_24479,N_24741);
xnor UO_1982 (O_1982,N_24208,N_24567);
or UO_1983 (O_1983,N_24446,N_24123);
nand UO_1984 (O_1984,N_24431,N_23880);
nand UO_1985 (O_1985,N_24199,N_24740);
and UO_1986 (O_1986,N_23798,N_24039);
and UO_1987 (O_1987,N_24975,N_24228);
xnor UO_1988 (O_1988,N_24207,N_24012);
or UO_1989 (O_1989,N_24127,N_24976);
and UO_1990 (O_1990,N_24780,N_24841);
nor UO_1991 (O_1991,N_24395,N_23970);
xor UO_1992 (O_1992,N_24163,N_24322);
and UO_1993 (O_1993,N_24991,N_23912);
nand UO_1994 (O_1994,N_24724,N_23788);
nor UO_1995 (O_1995,N_23915,N_24091);
nor UO_1996 (O_1996,N_24676,N_24089);
xor UO_1997 (O_1997,N_24189,N_23992);
nor UO_1998 (O_1998,N_24878,N_23995);
or UO_1999 (O_1999,N_24983,N_23959);
or UO_2000 (O_2000,N_24467,N_24000);
nor UO_2001 (O_2001,N_24190,N_24568);
xnor UO_2002 (O_2002,N_24675,N_24880);
and UO_2003 (O_2003,N_24081,N_24549);
nand UO_2004 (O_2004,N_24734,N_24481);
xnor UO_2005 (O_2005,N_24450,N_24253);
nand UO_2006 (O_2006,N_24920,N_24309);
nand UO_2007 (O_2007,N_24931,N_24841);
or UO_2008 (O_2008,N_24326,N_24331);
and UO_2009 (O_2009,N_24886,N_24655);
nand UO_2010 (O_2010,N_24868,N_24691);
nand UO_2011 (O_2011,N_24054,N_24874);
or UO_2012 (O_2012,N_24239,N_24027);
nor UO_2013 (O_2013,N_24696,N_24209);
and UO_2014 (O_2014,N_24257,N_23874);
xor UO_2015 (O_2015,N_24050,N_24995);
xor UO_2016 (O_2016,N_23792,N_24942);
xnor UO_2017 (O_2017,N_23868,N_24216);
nand UO_2018 (O_2018,N_24164,N_24726);
nand UO_2019 (O_2019,N_24689,N_23846);
nor UO_2020 (O_2020,N_24360,N_24463);
nor UO_2021 (O_2021,N_24901,N_24471);
or UO_2022 (O_2022,N_24648,N_23814);
or UO_2023 (O_2023,N_24816,N_24808);
nor UO_2024 (O_2024,N_24992,N_23781);
xor UO_2025 (O_2025,N_24984,N_24309);
or UO_2026 (O_2026,N_24637,N_24113);
or UO_2027 (O_2027,N_24642,N_24513);
or UO_2028 (O_2028,N_23971,N_23999);
nor UO_2029 (O_2029,N_23776,N_24857);
or UO_2030 (O_2030,N_24655,N_24587);
nand UO_2031 (O_2031,N_23827,N_23804);
or UO_2032 (O_2032,N_24978,N_24134);
and UO_2033 (O_2033,N_23934,N_24544);
xnor UO_2034 (O_2034,N_24060,N_23818);
nand UO_2035 (O_2035,N_24839,N_24264);
and UO_2036 (O_2036,N_24458,N_24516);
nand UO_2037 (O_2037,N_24302,N_24094);
or UO_2038 (O_2038,N_24617,N_23913);
nor UO_2039 (O_2039,N_24952,N_24284);
nor UO_2040 (O_2040,N_24636,N_24974);
xnor UO_2041 (O_2041,N_24500,N_24793);
or UO_2042 (O_2042,N_23790,N_24668);
nand UO_2043 (O_2043,N_24069,N_24049);
and UO_2044 (O_2044,N_24281,N_24911);
xor UO_2045 (O_2045,N_24885,N_23829);
or UO_2046 (O_2046,N_24541,N_24903);
xnor UO_2047 (O_2047,N_24884,N_24985);
and UO_2048 (O_2048,N_24267,N_24438);
xor UO_2049 (O_2049,N_24140,N_23816);
xnor UO_2050 (O_2050,N_24526,N_24705);
xor UO_2051 (O_2051,N_24284,N_24359);
nor UO_2052 (O_2052,N_24145,N_23917);
and UO_2053 (O_2053,N_23847,N_24236);
xnor UO_2054 (O_2054,N_24236,N_23931);
nand UO_2055 (O_2055,N_24792,N_23755);
or UO_2056 (O_2056,N_24313,N_24239);
xor UO_2057 (O_2057,N_24271,N_23945);
or UO_2058 (O_2058,N_23967,N_23934);
and UO_2059 (O_2059,N_23948,N_24934);
and UO_2060 (O_2060,N_24183,N_24301);
nor UO_2061 (O_2061,N_24838,N_24603);
xnor UO_2062 (O_2062,N_24091,N_24088);
or UO_2063 (O_2063,N_24378,N_24796);
nand UO_2064 (O_2064,N_24189,N_24247);
nand UO_2065 (O_2065,N_24032,N_23984);
nor UO_2066 (O_2066,N_24705,N_24098);
nand UO_2067 (O_2067,N_24615,N_23791);
nand UO_2068 (O_2068,N_24044,N_24901);
xor UO_2069 (O_2069,N_23961,N_24254);
or UO_2070 (O_2070,N_24410,N_24739);
and UO_2071 (O_2071,N_24541,N_24992);
or UO_2072 (O_2072,N_24460,N_23842);
xnor UO_2073 (O_2073,N_24421,N_24060);
or UO_2074 (O_2074,N_24903,N_24557);
and UO_2075 (O_2075,N_24031,N_24143);
nor UO_2076 (O_2076,N_24950,N_23978);
or UO_2077 (O_2077,N_24291,N_24604);
and UO_2078 (O_2078,N_24066,N_24575);
or UO_2079 (O_2079,N_24993,N_24929);
and UO_2080 (O_2080,N_24809,N_24045);
xnor UO_2081 (O_2081,N_24649,N_23932);
xnor UO_2082 (O_2082,N_24095,N_24611);
xnor UO_2083 (O_2083,N_23851,N_24270);
xnor UO_2084 (O_2084,N_24024,N_24146);
or UO_2085 (O_2085,N_24478,N_23837);
nor UO_2086 (O_2086,N_24679,N_24244);
nand UO_2087 (O_2087,N_24866,N_24351);
nand UO_2088 (O_2088,N_24100,N_23983);
or UO_2089 (O_2089,N_24836,N_24687);
xor UO_2090 (O_2090,N_24364,N_23894);
nand UO_2091 (O_2091,N_23947,N_24735);
and UO_2092 (O_2092,N_23781,N_24006);
or UO_2093 (O_2093,N_24596,N_24246);
nand UO_2094 (O_2094,N_23816,N_24531);
or UO_2095 (O_2095,N_24318,N_24034);
and UO_2096 (O_2096,N_24242,N_23951);
xnor UO_2097 (O_2097,N_24236,N_24279);
nand UO_2098 (O_2098,N_24357,N_24545);
xor UO_2099 (O_2099,N_24124,N_24710);
nand UO_2100 (O_2100,N_24435,N_24161);
xnor UO_2101 (O_2101,N_24989,N_23954);
xnor UO_2102 (O_2102,N_24973,N_24057);
xor UO_2103 (O_2103,N_23779,N_24055);
xor UO_2104 (O_2104,N_24231,N_24493);
nand UO_2105 (O_2105,N_24071,N_24642);
xnor UO_2106 (O_2106,N_24541,N_23957);
or UO_2107 (O_2107,N_23853,N_23800);
nand UO_2108 (O_2108,N_23997,N_24250);
and UO_2109 (O_2109,N_24708,N_24212);
nand UO_2110 (O_2110,N_24435,N_24916);
nor UO_2111 (O_2111,N_23821,N_24127);
nand UO_2112 (O_2112,N_24244,N_23925);
or UO_2113 (O_2113,N_24366,N_24072);
nor UO_2114 (O_2114,N_24079,N_24677);
or UO_2115 (O_2115,N_24303,N_23843);
or UO_2116 (O_2116,N_24588,N_24304);
and UO_2117 (O_2117,N_24431,N_24493);
nor UO_2118 (O_2118,N_24038,N_24960);
or UO_2119 (O_2119,N_24833,N_24886);
xnor UO_2120 (O_2120,N_24502,N_24066);
and UO_2121 (O_2121,N_24709,N_24560);
xnor UO_2122 (O_2122,N_24547,N_24682);
nand UO_2123 (O_2123,N_24800,N_23789);
nand UO_2124 (O_2124,N_24963,N_24281);
xnor UO_2125 (O_2125,N_24426,N_24711);
nor UO_2126 (O_2126,N_24670,N_24566);
xor UO_2127 (O_2127,N_24597,N_24277);
and UO_2128 (O_2128,N_24810,N_24395);
nand UO_2129 (O_2129,N_24991,N_24577);
nor UO_2130 (O_2130,N_24078,N_24460);
xor UO_2131 (O_2131,N_24954,N_24982);
nor UO_2132 (O_2132,N_24168,N_24382);
xor UO_2133 (O_2133,N_24378,N_24523);
nand UO_2134 (O_2134,N_24657,N_24575);
or UO_2135 (O_2135,N_23852,N_24318);
or UO_2136 (O_2136,N_24510,N_24193);
or UO_2137 (O_2137,N_24342,N_24401);
nand UO_2138 (O_2138,N_23826,N_24456);
nor UO_2139 (O_2139,N_24855,N_23806);
xor UO_2140 (O_2140,N_24602,N_24076);
nor UO_2141 (O_2141,N_24382,N_23875);
and UO_2142 (O_2142,N_24737,N_23869);
or UO_2143 (O_2143,N_24339,N_23968);
xor UO_2144 (O_2144,N_24622,N_24972);
or UO_2145 (O_2145,N_24694,N_24585);
xnor UO_2146 (O_2146,N_24284,N_23906);
nand UO_2147 (O_2147,N_24020,N_24751);
nand UO_2148 (O_2148,N_24981,N_24103);
xor UO_2149 (O_2149,N_24389,N_24275);
nand UO_2150 (O_2150,N_24940,N_24919);
nand UO_2151 (O_2151,N_23841,N_24219);
nand UO_2152 (O_2152,N_23907,N_24207);
or UO_2153 (O_2153,N_24269,N_24161);
xor UO_2154 (O_2154,N_24269,N_23868);
nor UO_2155 (O_2155,N_23925,N_24280);
xnor UO_2156 (O_2156,N_24100,N_24378);
xnor UO_2157 (O_2157,N_24256,N_24374);
and UO_2158 (O_2158,N_23915,N_24668);
or UO_2159 (O_2159,N_23763,N_23830);
or UO_2160 (O_2160,N_24744,N_23926);
or UO_2161 (O_2161,N_23781,N_23799);
or UO_2162 (O_2162,N_24118,N_24404);
or UO_2163 (O_2163,N_24779,N_24474);
and UO_2164 (O_2164,N_24049,N_24307);
nor UO_2165 (O_2165,N_24998,N_24896);
and UO_2166 (O_2166,N_23900,N_23919);
or UO_2167 (O_2167,N_24591,N_24365);
nor UO_2168 (O_2168,N_23804,N_24199);
xnor UO_2169 (O_2169,N_24917,N_24815);
or UO_2170 (O_2170,N_24720,N_24470);
or UO_2171 (O_2171,N_24565,N_24535);
xnor UO_2172 (O_2172,N_23825,N_24939);
and UO_2173 (O_2173,N_24487,N_23995);
or UO_2174 (O_2174,N_24324,N_24533);
xor UO_2175 (O_2175,N_23928,N_24348);
xnor UO_2176 (O_2176,N_23849,N_24779);
and UO_2177 (O_2177,N_24342,N_24372);
or UO_2178 (O_2178,N_24693,N_24324);
and UO_2179 (O_2179,N_23980,N_24252);
nand UO_2180 (O_2180,N_24721,N_24221);
nor UO_2181 (O_2181,N_23874,N_24364);
or UO_2182 (O_2182,N_24853,N_24861);
nor UO_2183 (O_2183,N_23780,N_24963);
xor UO_2184 (O_2184,N_24949,N_24622);
and UO_2185 (O_2185,N_24331,N_24888);
or UO_2186 (O_2186,N_24099,N_24486);
and UO_2187 (O_2187,N_24696,N_24364);
and UO_2188 (O_2188,N_24746,N_24620);
nor UO_2189 (O_2189,N_24998,N_24823);
nand UO_2190 (O_2190,N_24822,N_24173);
nor UO_2191 (O_2191,N_23926,N_24384);
nand UO_2192 (O_2192,N_24591,N_24914);
or UO_2193 (O_2193,N_24823,N_24083);
or UO_2194 (O_2194,N_23934,N_24134);
nor UO_2195 (O_2195,N_24220,N_24608);
and UO_2196 (O_2196,N_24255,N_24296);
nor UO_2197 (O_2197,N_24940,N_24378);
nor UO_2198 (O_2198,N_24957,N_23765);
and UO_2199 (O_2199,N_24082,N_24596);
or UO_2200 (O_2200,N_24630,N_23798);
or UO_2201 (O_2201,N_24084,N_24993);
nand UO_2202 (O_2202,N_24569,N_24813);
nand UO_2203 (O_2203,N_24896,N_23793);
or UO_2204 (O_2204,N_24865,N_24959);
nand UO_2205 (O_2205,N_24944,N_24530);
nand UO_2206 (O_2206,N_23760,N_24947);
xnor UO_2207 (O_2207,N_23869,N_24046);
nand UO_2208 (O_2208,N_23887,N_23836);
and UO_2209 (O_2209,N_24922,N_24490);
nand UO_2210 (O_2210,N_23820,N_23770);
nor UO_2211 (O_2211,N_24751,N_24242);
nand UO_2212 (O_2212,N_24641,N_24758);
nand UO_2213 (O_2213,N_24575,N_24834);
nor UO_2214 (O_2214,N_24721,N_24469);
or UO_2215 (O_2215,N_24705,N_24575);
or UO_2216 (O_2216,N_24294,N_24275);
or UO_2217 (O_2217,N_23975,N_23877);
and UO_2218 (O_2218,N_24589,N_23789);
or UO_2219 (O_2219,N_24920,N_24006);
and UO_2220 (O_2220,N_24754,N_24141);
nor UO_2221 (O_2221,N_24394,N_24756);
xnor UO_2222 (O_2222,N_23923,N_24441);
xnor UO_2223 (O_2223,N_24708,N_24405);
nor UO_2224 (O_2224,N_24421,N_24122);
and UO_2225 (O_2225,N_24508,N_24671);
nor UO_2226 (O_2226,N_24393,N_24278);
nor UO_2227 (O_2227,N_24101,N_24287);
nand UO_2228 (O_2228,N_24662,N_24493);
and UO_2229 (O_2229,N_24578,N_23969);
and UO_2230 (O_2230,N_23849,N_24674);
and UO_2231 (O_2231,N_24570,N_24346);
nand UO_2232 (O_2232,N_24359,N_24009);
xor UO_2233 (O_2233,N_24381,N_24923);
nand UO_2234 (O_2234,N_23810,N_24314);
and UO_2235 (O_2235,N_24556,N_24662);
and UO_2236 (O_2236,N_24384,N_24143);
or UO_2237 (O_2237,N_24626,N_24909);
nand UO_2238 (O_2238,N_24118,N_23837);
and UO_2239 (O_2239,N_23894,N_23997);
and UO_2240 (O_2240,N_23794,N_24326);
nor UO_2241 (O_2241,N_23973,N_24747);
or UO_2242 (O_2242,N_24749,N_24529);
and UO_2243 (O_2243,N_24117,N_24345);
nor UO_2244 (O_2244,N_24580,N_24009);
xnor UO_2245 (O_2245,N_24848,N_24339);
or UO_2246 (O_2246,N_24460,N_24090);
xnor UO_2247 (O_2247,N_24136,N_24632);
or UO_2248 (O_2248,N_24319,N_23801);
xor UO_2249 (O_2249,N_24792,N_24312);
nor UO_2250 (O_2250,N_24228,N_23751);
and UO_2251 (O_2251,N_24111,N_23804);
nor UO_2252 (O_2252,N_24926,N_24684);
xor UO_2253 (O_2253,N_24650,N_24779);
and UO_2254 (O_2254,N_24737,N_24476);
nand UO_2255 (O_2255,N_24010,N_23805);
nor UO_2256 (O_2256,N_24125,N_24920);
nand UO_2257 (O_2257,N_23794,N_23928);
and UO_2258 (O_2258,N_24858,N_24292);
and UO_2259 (O_2259,N_24696,N_24695);
nand UO_2260 (O_2260,N_23906,N_23767);
xnor UO_2261 (O_2261,N_24762,N_24253);
and UO_2262 (O_2262,N_24160,N_24615);
xor UO_2263 (O_2263,N_24292,N_24120);
xor UO_2264 (O_2264,N_24147,N_24800);
nand UO_2265 (O_2265,N_24404,N_24346);
or UO_2266 (O_2266,N_23958,N_24135);
nand UO_2267 (O_2267,N_24496,N_23951);
and UO_2268 (O_2268,N_24074,N_24846);
and UO_2269 (O_2269,N_23846,N_23844);
and UO_2270 (O_2270,N_23986,N_24319);
or UO_2271 (O_2271,N_24476,N_24263);
xor UO_2272 (O_2272,N_23806,N_24109);
nor UO_2273 (O_2273,N_24032,N_23957);
and UO_2274 (O_2274,N_24846,N_24485);
nor UO_2275 (O_2275,N_24227,N_24488);
or UO_2276 (O_2276,N_24785,N_24610);
xnor UO_2277 (O_2277,N_24237,N_24640);
nand UO_2278 (O_2278,N_24927,N_24509);
or UO_2279 (O_2279,N_24508,N_24028);
or UO_2280 (O_2280,N_24177,N_24450);
nor UO_2281 (O_2281,N_24843,N_23828);
and UO_2282 (O_2282,N_24425,N_24465);
xor UO_2283 (O_2283,N_24116,N_24831);
nor UO_2284 (O_2284,N_24360,N_23768);
nand UO_2285 (O_2285,N_24029,N_24686);
nand UO_2286 (O_2286,N_24719,N_24477);
or UO_2287 (O_2287,N_24613,N_24119);
or UO_2288 (O_2288,N_24555,N_24639);
nand UO_2289 (O_2289,N_23881,N_24387);
or UO_2290 (O_2290,N_24934,N_24748);
xor UO_2291 (O_2291,N_24224,N_24150);
or UO_2292 (O_2292,N_24594,N_24419);
nor UO_2293 (O_2293,N_24208,N_24563);
xnor UO_2294 (O_2294,N_24688,N_24565);
nand UO_2295 (O_2295,N_24928,N_23750);
and UO_2296 (O_2296,N_24015,N_23785);
xnor UO_2297 (O_2297,N_23837,N_24946);
nor UO_2298 (O_2298,N_24705,N_24126);
and UO_2299 (O_2299,N_24687,N_24608);
or UO_2300 (O_2300,N_24992,N_24031);
nor UO_2301 (O_2301,N_24772,N_24336);
xor UO_2302 (O_2302,N_24457,N_24416);
nor UO_2303 (O_2303,N_24729,N_24450);
nor UO_2304 (O_2304,N_23916,N_23950);
nor UO_2305 (O_2305,N_23832,N_24104);
nand UO_2306 (O_2306,N_24165,N_24402);
and UO_2307 (O_2307,N_24534,N_23879);
nand UO_2308 (O_2308,N_24017,N_24501);
nor UO_2309 (O_2309,N_23761,N_23983);
nor UO_2310 (O_2310,N_24417,N_24819);
xnor UO_2311 (O_2311,N_24253,N_24848);
nand UO_2312 (O_2312,N_24806,N_24195);
and UO_2313 (O_2313,N_24941,N_24237);
nand UO_2314 (O_2314,N_24649,N_24792);
xnor UO_2315 (O_2315,N_24803,N_24663);
and UO_2316 (O_2316,N_24736,N_23897);
xor UO_2317 (O_2317,N_23813,N_24573);
nand UO_2318 (O_2318,N_23964,N_24641);
nand UO_2319 (O_2319,N_23810,N_24772);
nand UO_2320 (O_2320,N_24401,N_24055);
nor UO_2321 (O_2321,N_24675,N_24674);
nand UO_2322 (O_2322,N_24040,N_24312);
and UO_2323 (O_2323,N_23953,N_24078);
and UO_2324 (O_2324,N_24928,N_24284);
and UO_2325 (O_2325,N_24134,N_23917);
or UO_2326 (O_2326,N_24543,N_24367);
and UO_2327 (O_2327,N_24331,N_24467);
and UO_2328 (O_2328,N_24479,N_23906);
and UO_2329 (O_2329,N_24877,N_24105);
and UO_2330 (O_2330,N_23862,N_24849);
nor UO_2331 (O_2331,N_24638,N_24870);
or UO_2332 (O_2332,N_24071,N_24439);
or UO_2333 (O_2333,N_24632,N_24081);
nand UO_2334 (O_2334,N_24614,N_24772);
or UO_2335 (O_2335,N_23802,N_24379);
or UO_2336 (O_2336,N_24914,N_24477);
nor UO_2337 (O_2337,N_24782,N_24065);
xnor UO_2338 (O_2338,N_24363,N_24107);
nand UO_2339 (O_2339,N_24301,N_24973);
xnor UO_2340 (O_2340,N_24742,N_24277);
and UO_2341 (O_2341,N_24914,N_24804);
nor UO_2342 (O_2342,N_24956,N_24660);
or UO_2343 (O_2343,N_24923,N_24328);
and UO_2344 (O_2344,N_24300,N_24630);
and UO_2345 (O_2345,N_24176,N_24976);
nor UO_2346 (O_2346,N_24398,N_24697);
or UO_2347 (O_2347,N_23922,N_23794);
xnor UO_2348 (O_2348,N_24806,N_24752);
xor UO_2349 (O_2349,N_24503,N_23957);
or UO_2350 (O_2350,N_23917,N_23841);
or UO_2351 (O_2351,N_23978,N_24450);
nor UO_2352 (O_2352,N_24354,N_24120);
nand UO_2353 (O_2353,N_24619,N_23943);
and UO_2354 (O_2354,N_24771,N_24650);
nor UO_2355 (O_2355,N_23922,N_24150);
nor UO_2356 (O_2356,N_24194,N_24643);
or UO_2357 (O_2357,N_24574,N_24718);
and UO_2358 (O_2358,N_24638,N_24280);
or UO_2359 (O_2359,N_24796,N_24759);
xnor UO_2360 (O_2360,N_24068,N_23774);
xor UO_2361 (O_2361,N_24735,N_24663);
nand UO_2362 (O_2362,N_24077,N_24796);
xnor UO_2363 (O_2363,N_24096,N_24687);
nand UO_2364 (O_2364,N_24627,N_24140);
nor UO_2365 (O_2365,N_24633,N_24111);
or UO_2366 (O_2366,N_23873,N_24135);
and UO_2367 (O_2367,N_24896,N_24454);
nor UO_2368 (O_2368,N_23902,N_24377);
xor UO_2369 (O_2369,N_24132,N_23992);
and UO_2370 (O_2370,N_24068,N_24066);
nand UO_2371 (O_2371,N_24612,N_24936);
nand UO_2372 (O_2372,N_24818,N_24258);
nor UO_2373 (O_2373,N_24959,N_24893);
xnor UO_2374 (O_2374,N_23799,N_24582);
xnor UO_2375 (O_2375,N_24696,N_24551);
or UO_2376 (O_2376,N_23947,N_24108);
xor UO_2377 (O_2377,N_24356,N_24761);
or UO_2378 (O_2378,N_23911,N_23968);
nor UO_2379 (O_2379,N_23916,N_23976);
nor UO_2380 (O_2380,N_23954,N_24792);
xor UO_2381 (O_2381,N_24698,N_24274);
nor UO_2382 (O_2382,N_24129,N_24639);
and UO_2383 (O_2383,N_24831,N_23837);
nand UO_2384 (O_2384,N_23875,N_24435);
and UO_2385 (O_2385,N_24024,N_24372);
or UO_2386 (O_2386,N_24608,N_24015);
or UO_2387 (O_2387,N_24016,N_24314);
and UO_2388 (O_2388,N_24990,N_24076);
nor UO_2389 (O_2389,N_24915,N_24335);
and UO_2390 (O_2390,N_24880,N_24029);
nor UO_2391 (O_2391,N_24026,N_24885);
nand UO_2392 (O_2392,N_24416,N_24407);
nand UO_2393 (O_2393,N_24944,N_24378);
and UO_2394 (O_2394,N_24421,N_24791);
or UO_2395 (O_2395,N_24625,N_23906);
nor UO_2396 (O_2396,N_24243,N_24246);
nor UO_2397 (O_2397,N_24958,N_24529);
and UO_2398 (O_2398,N_24748,N_24749);
and UO_2399 (O_2399,N_24133,N_23862);
nand UO_2400 (O_2400,N_24688,N_24879);
xnor UO_2401 (O_2401,N_24356,N_24089);
and UO_2402 (O_2402,N_24213,N_24746);
nor UO_2403 (O_2403,N_24144,N_23777);
xnor UO_2404 (O_2404,N_24098,N_23776);
or UO_2405 (O_2405,N_23913,N_23990);
nor UO_2406 (O_2406,N_24869,N_24809);
nor UO_2407 (O_2407,N_23874,N_23783);
xor UO_2408 (O_2408,N_24955,N_24128);
or UO_2409 (O_2409,N_24117,N_24494);
nand UO_2410 (O_2410,N_24659,N_23782);
nor UO_2411 (O_2411,N_23998,N_24803);
nand UO_2412 (O_2412,N_23939,N_24587);
nor UO_2413 (O_2413,N_24023,N_24049);
nand UO_2414 (O_2414,N_24472,N_23877);
or UO_2415 (O_2415,N_24784,N_24868);
nor UO_2416 (O_2416,N_24726,N_23787);
nor UO_2417 (O_2417,N_24447,N_24087);
xor UO_2418 (O_2418,N_23879,N_24286);
nand UO_2419 (O_2419,N_24402,N_24699);
xor UO_2420 (O_2420,N_24660,N_24271);
nor UO_2421 (O_2421,N_23864,N_23860);
nand UO_2422 (O_2422,N_24357,N_23901);
nand UO_2423 (O_2423,N_24609,N_24985);
nor UO_2424 (O_2424,N_24824,N_24644);
and UO_2425 (O_2425,N_24823,N_24438);
or UO_2426 (O_2426,N_24124,N_24663);
or UO_2427 (O_2427,N_24474,N_24511);
nand UO_2428 (O_2428,N_24379,N_23921);
nand UO_2429 (O_2429,N_24513,N_24856);
nand UO_2430 (O_2430,N_24615,N_24063);
xnor UO_2431 (O_2431,N_24917,N_24008);
and UO_2432 (O_2432,N_24912,N_23994);
nand UO_2433 (O_2433,N_24021,N_24097);
xnor UO_2434 (O_2434,N_23883,N_24585);
or UO_2435 (O_2435,N_23971,N_23792);
or UO_2436 (O_2436,N_24785,N_24458);
nor UO_2437 (O_2437,N_24470,N_24590);
or UO_2438 (O_2438,N_24937,N_24766);
nand UO_2439 (O_2439,N_23814,N_24693);
and UO_2440 (O_2440,N_24369,N_24030);
xnor UO_2441 (O_2441,N_24854,N_24540);
and UO_2442 (O_2442,N_24684,N_24475);
xnor UO_2443 (O_2443,N_24264,N_24983);
and UO_2444 (O_2444,N_24112,N_24687);
nor UO_2445 (O_2445,N_24962,N_24974);
and UO_2446 (O_2446,N_24374,N_24086);
xnor UO_2447 (O_2447,N_24790,N_24606);
or UO_2448 (O_2448,N_24651,N_24049);
nand UO_2449 (O_2449,N_23974,N_24638);
and UO_2450 (O_2450,N_24082,N_23877);
and UO_2451 (O_2451,N_23855,N_24331);
nand UO_2452 (O_2452,N_24294,N_24185);
nand UO_2453 (O_2453,N_23865,N_23978);
nor UO_2454 (O_2454,N_24494,N_24381);
and UO_2455 (O_2455,N_24616,N_24848);
nand UO_2456 (O_2456,N_24978,N_24981);
or UO_2457 (O_2457,N_24245,N_24347);
nand UO_2458 (O_2458,N_24118,N_24082);
or UO_2459 (O_2459,N_24696,N_24805);
nand UO_2460 (O_2460,N_24477,N_24166);
xnor UO_2461 (O_2461,N_24440,N_23843);
and UO_2462 (O_2462,N_23785,N_24583);
nand UO_2463 (O_2463,N_24446,N_24565);
nand UO_2464 (O_2464,N_23828,N_24731);
nand UO_2465 (O_2465,N_24365,N_24032);
or UO_2466 (O_2466,N_23851,N_24656);
nand UO_2467 (O_2467,N_24316,N_24629);
and UO_2468 (O_2468,N_24633,N_24908);
or UO_2469 (O_2469,N_24776,N_24492);
nor UO_2470 (O_2470,N_24512,N_24825);
nor UO_2471 (O_2471,N_24795,N_24988);
or UO_2472 (O_2472,N_23889,N_24224);
xnor UO_2473 (O_2473,N_24621,N_24742);
nor UO_2474 (O_2474,N_24478,N_24966);
nand UO_2475 (O_2475,N_24984,N_23884);
nand UO_2476 (O_2476,N_24246,N_24435);
or UO_2477 (O_2477,N_24987,N_24292);
and UO_2478 (O_2478,N_24077,N_23948);
nor UO_2479 (O_2479,N_23871,N_24398);
nand UO_2480 (O_2480,N_24514,N_24191);
nand UO_2481 (O_2481,N_23876,N_24372);
xor UO_2482 (O_2482,N_24521,N_24616);
and UO_2483 (O_2483,N_24835,N_24170);
or UO_2484 (O_2484,N_24978,N_24550);
nand UO_2485 (O_2485,N_23904,N_23790);
nand UO_2486 (O_2486,N_24880,N_24942);
or UO_2487 (O_2487,N_24464,N_24419);
nor UO_2488 (O_2488,N_24861,N_24049);
nor UO_2489 (O_2489,N_24879,N_24383);
or UO_2490 (O_2490,N_24736,N_24952);
nand UO_2491 (O_2491,N_23829,N_24050);
nand UO_2492 (O_2492,N_24004,N_24879);
or UO_2493 (O_2493,N_24356,N_24743);
or UO_2494 (O_2494,N_24665,N_24312);
or UO_2495 (O_2495,N_23915,N_24544);
nor UO_2496 (O_2496,N_23925,N_24243);
and UO_2497 (O_2497,N_24217,N_24369);
nand UO_2498 (O_2498,N_23764,N_24901);
nand UO_2499 (O_2499,N_24146,N_24910);
and UO_2500 (O_2500,N_24080,N_24375);
and UO_2501 (O_2501,N_24091,N_24587);
or UO_2502 (O_2502,N_23845,N_23931);
or UO_2503 (O_2503,N_24435,N_23762);
nand UO_2504 (O_2504,N_24806,N_23864);
or UO_2505 (O_2505,N_24046,N_23966);
xor UO_2506 (O_2506,N_23945,N_24716);
nand UO_2507 (O_2507,N_24188,N_24496);
and UO_2508 (O_2508,N_24626,N_24751);
and UO_2509 (O_2509,N_24403,N_24028);
nand UO_2510 (O_2510,N_24003,N_24544);
and UO_2511 (O_2511,N_24026,N_24303);
and UO_2512 (O_2512,N_24802,N_24416);
nand UO_2513 (O_2513,N_23886,N_24396);
nand UO_2514 (O_2514,N_24883,N_24489);
or UO_2515 (O_2515,N_24484,N_24615);
and UO_2516 (O_2516,N_24730,N_24580);
or UO_2517 (O_2517,N_24775,N_24081);
nand UO_2518 (O_2518,N_24171,N_24563);
nand UO_2519 (O_2519,N_23944,N_23987);
and UO_2520 (O_2520,N_24375,N_24469);
or UO_2521 (O_2521,N_24933,N_24714);
nand UO_2522 (O_2522,N_24781,N_23935);
and UO_2523 (O_2523,N_24606,N_24932);
nor UO_2524 (O_2524,N_24455,N_24263);
or UO_2525 (O_2525,N_24556,N_24467);
or UO_2526 (O_2526,N_24949,N_24771);
nand UO_2527 (O_2527,N_24631,N_24979);
xor UO_2528 (O_2528,N_24816,N_24263);
xor UO_2529 (O_2529,N_24044,N_24527);
and UO_2530 (O_2530,N_23994,N_23781);
and UO_2531 (O_2531,N_24062,N_24402);
nand UO_2532 (O_2532,N_24145,N_24991);
or UO_2533 (O_2533,N_23904,N_24416);
and UO_2534 (O_2534,N_24602,N_24501);
or UO_2535 (O_2535,N_24604,N_24645);
xnor UO_2536 (O_2536,N_24947,N_24130);
nand UO_2537 (O_2537,N_24046,N_23891);
or UO_2538 (O_2538,N_24614,N_24842);
nand UO_2539 (O_2539,N_24835,N_24792);
nor UO_2540 (O_2540,N_24539,N_24692);
nand UO_2541 (O_2541,N_24792,N_23784);
nor UO_2542 (O_2542,N_24396,N_24522);
and UO_2543 (O_2543,N_24660,N_23981);
and UO_2544 (O_2544,N_24564,N_24773);
nand UO_2545 (O_2545,N_23776,N_24053);
or UO_2546 (O_2546,N_24136,N_24554);
or UO_2547 (O_2547,N_24955,N_24745);
nor UO_2548 (O_2548,N_23940,N_24478);
nand UO_2549 (O_2549,N_24622,N_24978);
or UO_2550 (O_2550,N_24386,N_23959);
and UO_2551 (O_2551,N_23832,N_24837);
or UO_2552 (O_2552,N_24365,N_24047);
or UO_2553 (O_2553,N_23894,N_24624);
and UO_2554 (O_2554,N_23879,N_24199);
and UO_2555 (O_2555,N_24068,N_24132);
xnor UO_2556 (O_2556,N_24053,N_24693);
and UO_2557 (O_2557,N_24062,N_24263);
nand UO_2558 (O_2558,N_24942,N_24902);
xor UO_2559 (O_2559,N_24306,N_23961);
nor UO_2560 (O_2560,N_24216,N_24809);
nand UO_2561 (O_2561,N_23786,N_23791);
nand UO_2562 (O_2562,N_24219,N_24509);
or UO_2563 (O_2563,N_24461,N_24322);
nand UO_2564 (O_2564,N_24719,N_24284);
nor UO_2565 (O_2565,N_24590,N_24365);
nor UO_2566 (O_2566,N_24073,N_24453);
nand UO_2567 (O_2567,N_23796,N_24743);
nand UO_2568 (O_2568,N_24000,N_24260);
nor UO_2569 (O_2569,N_23851,N_23868);
xor UO_2570 (O_2570,N_24981,N_24824);
or UO_2571 (O_2571,N_24935,N_23809);
and UO_2572 (O_2572,N_23934,N_23900);
and UO_2573 (O_2573,N_24474,N_24707);
nand UO_2574 (O_2574,N_24939,N_24727);
xor UO_2575 (O_2575,N_23918,N_24501);
or UO_2576 (O_2576,N_24593,N_24344);
or UO_2577 (O_2577,N_24586,N_23788);
nand UO_2578 (O_2578,N_24716,N_24687);
nand UO_2579 (O_2579,N_24542,N_24959);
xor UO_2580 (O_2580,N_24336,N_24480);
or UO_2581 (O_2581,N_23829,N_24062);
nor UO_2582 (O_2582,N_24665,N_24585);
nor UO_2583 (O_2583,N_24123,N_24723);
xnor UO_2584 (O_2584,N_24966,N_24595);
and UO_2585 (O_2585,N_24272,N_24343);
or UO_2586 (O_2586,N_24534,N_24242);
or UO_2587 (O_2587,N_24518,N_24371);
nor UO_2588 (O_2588,N_24173,N_24025);
or UO_2589 (O_2589,N_24944,N_23796);
xor UO_2590 (O_2590,N_23961,N_24338);
nand UO_2591 (O_2591,N_23874,N_24602);
or UO_2592 (O_2592,N_24434,N_24061);
nor UO_2593 (O_2593,N_24601,N_24875);
and UO_2594 (O_2594,N_23841,N_24784);
or UO_2595 (O_2595,N_24602,N_24316);
nor UO_2596 (O_2596,N_24382,N_24973);
or UO_2597 (O_2597,N_24114,N_24570);
xor UO_2598 (O_2598,N_24415,N_24932);
or UO_2599 (O_2599,N_24857,N_24077);
xor UO_2600 (O_2600,N_24439,N_24010);
nand UO_2601 (O_2601,N_24366,N_23766);
xor UO_2602 (O_2602,N_23840,N_24962);
xor UO_2603 (O_2603,N_24860,N_23884);
nand UO_2604 (O_2604,N_24451,N_24928);
or UO_2605 (O_2605,N_24223,N_23901);
nand UO_2606 (O_2606,N_24628,N_24924);
nand UO_2607 (O_2607,N_24805,N_24698);
xor UO_2608 (O_2608,N_24785,N_24581);
xor UO_2609 (O_2609,N_24834,N_24617);
and UO_2610 (O_2610,N_23947,N_24801);
nand UO_2611 (O_2611,N_24129,N_24297);
and UO_2612 (O_2612,N_24565,N_24963);
nor UO_2613 (O_2613,N_24638,N_24592);
nand UO_2614 (O_2614,N_23944,N_24963);
and UO_2615 (O_2615,N_24198,N_23973);
nand UO_2616 (O_2616,N_24058,N_24145);
or UO_2617 (O_2617,N_24902,N_24633);
nand UO_2618 (O_2618,N_24352,N_24057);
xor UO_2619 (O_2619,N_24593,N_24174);
or UO_2620 (O_2620,N_24036,N_24232);
or UO_2621 (O_2621,N_24343,N_24659);
or UO_2622 (O_2622,N_23931,N_24181);
xnor UO_2623 (O_2623,N_24444,N_24316);
or UO_2624 (O_2624,N_24644,N_24467);
nor UO_2625 (O_2625,N_24460,N_23871);
and UO_2626 (O_2626,N_24081,N_24731);
or UO_2627 (O_2627,N_24370,N_24139);
or UO_2628 (O_2628,N_24074,N_24813);
or UO_2629 (O_2629,N_24570,N_24496);
or UO_2630 (O_2630,N_24074,N_24614);
xor UO_2631 (O_2631,N_24685,N_23877);
and UO_2632 (O_2632,N_24581,N_24351);
nand UO_2633 (O_2633,N_24799,N_23891);
and UO_2634 (O_2634,N_24620,N_24186);
nand UO_2635 (O_2635,N_24866,N_24025);
nand UO_2636 (O_2636,N_24673,N_24159);
and UO_2637 (O_2637,N_24440,N_24304);
xnor UO_2638 (O_2638,N_23899,N_24425);
nand UO_2639 (O_2639,N_24457,N_24594);
xnor UO_2640 (O_2640,N_24106,N_24301);
or UO_2641 (O_2641,N_23992,N_24458);
nand UO_2642 (O_2642,N_23882,N_24122);
or UO_2643 (O_2643,N_24566,N_24175);
or UO_2644 (O_2644,N_24647,N_24825);
or UO_2645 (O_2645,N_24729,N_23818);
nand UO_2646 (O_2646,N_24658,N_24745);
nand UO_2647 (O_2647,N_24161,N_24102);
and UO_2648 (O_2648,N_23978,N_24320);
xnor UO_2649 (O_2649,N_24013,N_24760);
nand UO_2650 (O_2650,N_23826,N_24205);
nand UO_2651 (O_2651,N_24701,N_24445);
nand UO_2652 (O_2652,N_23955,N_24528);
or UO_2653 (O_2653,N_24607,N_24512);
xor UO_2654 (O_2654,N_24164,N_23950);
and UO_2655 (O_2655,N_24634,N_23756);
and UO_2656 (O_2656,N_23836,N_24775);
and UO_2657 (O_2657,N_24769,N_24577);
nor UO_2658 (O_2658,N_24356,N_24919);
or UO_2659 (O_2659,N_24534,N_24923);
nand UO_2660 (O_2660,N_24255,N_23917);
nor UO_2661 (O_2661,N_24017,N_24483);
or UO_2662 (O_2662,N_23835,N_24980);
and UO_2663 (O_2663,N_24475,N_24770);
xor UO_2664 (O_2664,N_23853,N_24872);
nor UO_2665 (O_2665,N_24976,N_23917);
or UO_2666 (O_2666,N_24053,N_23806);
nor UO_2667 (O_2667,N_24016,N_24476);
nor UO_2668 (O_2668,N_24190,N_24629);
nand UO_2669 (O_2669,N_24183,N_24493);
nor UO_2670 (O_2670,N_24813,N_24005);
and UO_2671 (O_2671,N_23914,N_24834);
or UO_2672 (O_2672,N_24143,N_24896);
or UO_2673 (O_2673,N_24043,N_24059);
and UO_2674 (O_2674,N_24751,N_24618);
and UO_2675 (O_2675,N_24959,N_24726);
or UO_2676 (O_2676,N_23875,N_24698);
or UO_2677 (O_2677,N_23807,N_24539);
or UO_2678 (O_2678,N_24479,N_24952);
and UO_2679 (O_2679,N_24388,N_24158);
xor UO_2680 (O_2680,N_24686,N_23871);
xnor UO_2681 (O_2681,N_24384,N_24490);
nor UO_2682 (O_2682,N_24883,N_23848);
and UO_2683 (O_2683,N_23967,N_23891);
or UO_2684 (O_2684,N_24602,N_24692);
nor UO_2685 (O_2685,N_24904,N_23822);
and UO_2686 (O_2686,N_23816,N_24610);
and UO_2687 (O_2687,N_24079,N_24866);
xnor UO_2688 (O_2688,N_24454,N_24635);
xnor UO_2689 (O_2689,N_24705,N_24239);
nand UO_2690 (O_2690,N_24090,N_24771);
nor UO_2691 (O_2691,N_24705,N_24857);
or UO_2692 (O_2692,N_24618,N_24648);
or UO_2693 (O_2693,N_23858,N_24969);
nor UO_2694 (O_2694,N_24261,N_24505);
nand UO_2695 (O_2695,N_24229,N_24453);
or UO_2696 (O_2696,N_24746,N_24050);
nor UO_2697 (O_2697,N_23931,N_24984);
or UO_2698 (O_2698,N_24840,N_24388);
nand UO_2699 (O_2699,N_23780,N_24879);
nor UO_2700 (O_2700,N_24247,N_23790);
and UO_2701 (O_2701,N_24815,N_23951);
or UO_2702 (O_2702,N_23805,N_24069);
xor UO_2703 (O_2703,N_24492,N_23767);
nand UO_2704 (O_2704,N_24160,N_24385);
nand UO_2705 (O_2705,N_24929,N_24025);
xor UO_2706 (O_2706,N_23963,N_24736);
nor UO_2707 (O_2707,N_24112,N_24199);
and UO_2708 (O_2708,N_24656,N_23896);
xnor UO_2709 (O_2709,N_24535,N_24219);
nor UO_2710 (O_2710,N_24926,N_23822);
and UO_2711 (O_2711,N_24674,N_23914);
xor UO_2712 (O_2712,N_24455,N_24461);
nand UO_2713 (O_2713,N_24952,N_24272);
nand UO_2714 (O_2714,N_24587,N_23774);
and UO_2715 (O_2715,N_24596,N_24707);
or UO_2716 (O_2716,N_24720,N_24020);
or UO_2717 (O_2717,N_24499,N_23876);
nor UO_2718 (O_2718,N_23939,N_24348);
and UO_2719 (O_2719,N_24811,N_24550);
nor UO_2720 (O_2720,N_24182,N_24601);
nor UO_2721 (O_2721,N_24948,N_24733);
and UO_2722 (O_2722,N_24237,N_24159);
and UO_2723 (O_2723,N_24196,N_24749);
and UO_2724 (O_2724,N_24501,N_24872);
and UO_2725 (O_2725,N_24134,N_24860);
or UO_2726 (O_2726,N_23758,N_24370);
nor UO_2727 (O_2727,N_24784,N_24126);
or UO_2728 (O_2728,N_23923,N_23821);
nor UO_2729 (O_2729,N_23967,N_24197);
nor UO_2730 (O_2730,N_23950,N_24753);
nor UO_2731 (O_2731,N_24727,N_24440);
nand UO_2732 (O_2732,N_24230,N_24839);
nor UO_2733 (O_2733,N_24039,N_24566);
xor UO_2734 (O_2734,N_23930,N_24057);
xnor UO_2735 (O_2735,N_24541,N_24735);
nand UO_2736 (O_2736,N_24252,N_24815);
xnor UO_2737 (O_2737,N_24672,N_24985);
nor UO_2738 (O_2738,N_24629,N_24744);
or UO_2739 (O_2739,N_24247,N_24851);
or UO_2740 (O_2740,N_24030,N_24703);
or UO_2741 (O_2741,N_23868,N_23912);
or UO_2742 (O_2742,N_23816,N_24548);
and UO_2743 (O_2743,N_24007,N_24740);
nand UO_2744 (O_2744,N_24631,N_23975);
or UO_2745 (O_2745,N_24855,N_24738);
nor UO_2746 (O_2746,N_24280,N_24275);
nand UO_2747 (O_2747,N_24506,N_24619);
and UO_2748 (O_2748,N_24322,N_24992);
and UO_2749 (O_2749,N_24189,N_24275);
and UO_2750 (O_2750,N_23781,N_24999);
xor UO_2751 (O_2751,N_23982,N_24063);
nand UO_2752 (O_2752,N_24252,N_24218);
or UO_2753 (O_2753,N_23956,N_24582);
or UO_2754 (O_2754,N_24055,N_24449);
or UO_2755 (O_2755,N_23995,N_24716);
xor UO_2756 (O_2756,N_24556,N_24972);
or UO_2757 (O_2757,N_24556,N_24666);
xor UO_2758 (O_2758,N_23996,N_24392);
and UO_2759 (O_2759,N_24764,N_24645);
xor UO_2760 (O_2760,N_23908,N_24631);
nor UO_2761 (O_2761,N_24891,N_23880);
nor UO_2762 (O_2762,N_23890,N_24284);
nand UO_2763 (O_2763,N_24541,N_24889);
or UO_2764 (O_2764,N_23893,N_24541);
or UO_2765 (O_2765,N_24440,N_23880);
and UO_2766 (O_2766,N_23938,N_24680);
and UO_2767 (O_2767,N_23834,N_24109);
nor UO_2768 (O_2768,N_23961,N_24126);
and UO_2769 (O_2769,N_24413,N_23805);
xnor UO_2770 (O_2770,N_24979,N_23768);
xor UO_2771 (O_2771,N_23994,N_24109);
nor UO_2772 (O_2772,N_24381,N_24818);
nor UO_2773 (O_2773,N_24228,N_24752);
or UO_2774 (O_2774,N_24091,N_24160);
xor UO_2775 (O_2775,N_23978,N_23775);
nor UO_2776 (O_2776,N_23815,N_24220);
nor UO_2777 (O_2777,N_24194,N_24310);
nand UO_2778 (O_2778,N_24784,N_23889);
nand UO_2779 (O_2779,N_24239,N_24699);
or UO_2780 (O_2780,N_24462,N_24154);
or UO_2781 (O_2781,N_24347,N_24708);
and UO_2782 (O_2782,N_24441,N_23782);
xnor UO_2783 (O_2783,N_24158,N_24981);
xnor UO_2784 (O_2784,N_24935,N_24989);
or UO_2785 (O_2785,N_24435,N_24579);
xor UO_2786 (O_2786,N_24129,N_24289);
and UO_2787 (O_2787,N_24800,N_24323);
nand UO_2788 (O_2788,N_24630,N_24602);
nor UO_2789 (O_2789,N_23968,N_23947);
nor UO_2790 (O_2790,N_24905,N_24107);
and UO_2791 (O_2791,N_24462,N_24074);
xor UO_2792 (O_2792,N_24960,N_24432);
and UO_2793 (O_2793,N_24521,N_23889);
nand UO_2794 (O_2794,N_24557,N_24335);
or UO_2795 (O_2795,N_24422,N_24311);
and UO_2796 (O_2796,N_23982,N_24437);
nor UO_2797 (O_2797,N_24772,N_24267);
xnor UO_2798 (O_2798,N_24739,N_24237);
xnor UO_2799 (O_2799,N_24945,N_24890);
xor UO_2800 (O_2800,N_24171,N_24680);
nand UO_2801 (O_2801,N_24063,N_24241);
xor UO_2802 (O_2802,N_24922,N_24259);
nor UO_2803 (O_2803,N_23785,N_24975);
and UO_2804 (O_2804,N_24768,N_24041);
nand UO_2805 (O_2805,N_24837,N_24557);
xor UO_2806 (O_2806,N_24781,N_24664);
nor UO_2807 (O_2807,N_23807,N_23967);
nor UO_2808 (O_2808,N_23892,N_24778);
nand UO_2809 (O_2809,N_24503,N_24720);
xor UO_2810 (O_2810,N_23755,N_23839);
nand UO_2811 (O_2811,N_24073,N_24205);
nand UO_2812 (O_2812,N_24049,N_23916);
nand UO_2813 (O_2813,N_24780,N_23824);
or UO_2814 (O_2814,N_24393,N_23957);
nand UO_2815 (O_2815,N_24969,N_24894);
and UO_2816 (O_2816,N_24669,N_24658);
xnor UO_2817 (O_2817,N_24409,N_24432);
nand UO_2818 (O_2818,N_24269,N_24966);
and UO_2819 (O_2819,N_24622,N_24716);
nand UO_2820 (O_2820,N_23984,N_24662);
and UO_2821 (O_2821,N_24367,N_24887);
xnor UO_2822 (O_2822,N_23959,N_24212);
or UO_2823 (O_2823,N_24558,N_24215);
or UO_2824 (O_2824,N_24209,N_24561);
xor UO_2825 (O_2825,N_24836,N_23830);
nand UO_2826 (O_2826,N_24899,N_23887);
nand UO_2827 (O_2827,N_23861,N_24645);
or UO_2828 (O_2828,N_24999,N_24058);
xnor UO_2829 (O_2829,N_24147,N_24674);
xnor UO_2830 (O_2830,N_24405,N_24557);
nand UO_2831 (O_2831,N_23881,N_24469);
nand UO_2832 (O_2832,N_24723,N_24917);
nand UO_2833 (O_2833,N_24068,N_23846);
or UO_2834 (O_2834,N_24370,N_24185);
or UO_2835 (O_2835,N_23903,N_24845);
xor UO_2836 (O_2836,N_24611,N_24991);
nor UO_2837 (O_2837,N_23854,N_24798);
and UO_2838 (O_2838,N_24589,N_24501);
xor UO_2839 (O_2839,N_24830,N_23889);
xnor UO_2840 (O_2840,N_24600,N_24374);
and UO_2841 (O_2841,N_24567,N_24548);
xnor UO_2842 (O_2842,N_24156,N_24419);
nand UO_2843 (O_2843,N_24387,N_24936);
nand UO_2844 (O_2844,N_24103,N_24031);
and UO_2845 (O_2845,N_24929,N_24293);
and UO_2846 (O_2846,N_24761,N_24154);
nor UO_2847 (O_2847,N_24994,N_24081);
nor UO_2848 (O_2848,N_24328,N_24924);
nor UO_2849 (O_2849,N_24808,N_24117);
nand UO_2850 (O_2850,N_24624,N_24897);
nor UO_2851 (O_2851,N_24555,N_23889);
and UO_2852 (O_2852,N_24951,N_24059);
xnor UO_2853 (O_2853,N_23982,N_24051);
nand UO_2854 (O_2854,N_24054,N_24087);
or UO_2855 (O_2855,N_23935,N_24990);
nor UO_2856 (O_2856,N_24494,N_23893);
nor UO_2857 (O_2857,N_24280,N_24375);
nand UO_2858 (O_2858,N_24116,N_24247);
nand UO_2859 (O_2859,N_24837,N_24637);
or UO_2860 (O_2860,N_24260,N_24181);
nor UO_2861 (O_2861,N_24540,N_23796);
nor UO_2862 (O_2862,N_23986,N_24348);
and UO_2863 (O_2863,N_24856,N_24997);
and UO_2864 (O_2864,N_24099,N_24607);
or UO_2865 (O_2865,N_24206,N_23956);
and UO_2866 (O_2866,N_23835,N_24449);
nand UO_2867 (O_2867,N_24843,N_24828);
or UO_2868 (O_2868,N_23820,N_24892);
nor UO_2869 (O_2869,N_24008,N_24371);
or UO_2870 (O_2870,N_24013,N_24921);
or UO_2871 (O_2871,N_24011,N_24354);
or UO_2872 (O_2872,N_24685,N_24125);
and UO_2873 (O_2873,N_24718,N_24959);
or UO_2874 (O_2874,N_23933,N_23794);
xor UO_2875 (O_2875,N_23996,N_24063);
or UO_2876 (O_2876,N_24208,N_24607);
and UO_2877 (O_2877,N_24291,N_24962);
nand UO_2878 (O_2878,N_24639,N_24087);
nor UO_2879 (O_2879,N_24337,N_24265);
and UO_2880 (O_2880,N_23758,N_24116);
and UO_2881 (O_2881,N_24479,N_24977);
xnor UO_2882 (O_2882,N_23929,N_24742);
xnor UO_2883 (O_2883,N_24108,N_24118);
and UO_2884 (O_2884,N_24436,N_24668);
xor UO_2885 (O_2885,N_24195,N_24202);
nand UO_2886 (O_2886,N_24067,N_23835);
nor UO_2887 (O_2887,N_24037,N_24946);
xor UO_2888 (O_2888,N_23778,N_24377);
and UO_2889 (O_2889,N_24894,N_24956);
xnor UO_2890 (O_2890,N_24523,N_24817);
or UO_2891 (O_2891,N_23961,N_23806);
xnor UO_2892 (O_2892,N_24757,N_24046);
nor UO_2893 (O_2893,N_24408,N_23903);
and UO_2894 (O_2894,N_24141,N_24958);
nor UO_2895 (O_2895,N_24156,N_24304);
nor UO_2896 (O_2896,N_24217,N_23908);
nor UO_2897 (O_2897,N_24448,N_24369);
nor UO_2898 (O_2898,N_24383,N_23911);
nand UO_2899 (O_2899,N_24934,N_24935);
or UO_2900 (O_2900,N_24546,N_23880);
nor UO_2901 (O_2901,N_24929,N_23864);
nor UO_2902 (O_2902,N_24282,N_23980);
nor UO_2903 (O_2903,N_24054,N_24303);
nand UO_2904 (O_2904,N_23935,N_23878);
nand UO_2905 (O_2905,N_24395,N_23844);
or UO_2906 (O_2906,N_24246,N_24462);
and UO_2907 (O_2907,N_24199,N_24082);
nor UO_2908 (O_2908,N_24860,N_24368);
nand UO_2909 (O_2909,N_24256,N_24091);
nor UO_2910 (O_2910,N_24688,N_24836);
nor UO_2911 (O_2911,N_23950,N_24613);
or UO_2912 (O_2912,N_24321,N_23779);
xor UO_2913 (O_2913,N_23838,N_24623);
xnor UO_2914 (O_2914,N_24956,N_24688);
and UO_2915 (O_2915,N_24882,N_24263);
or UO_2916 (O_2916,N_24078,N_24551);
or UO_2917 (O_2917,N_23969,N_23999);
xor UO_2918 (O_2918,N_24191,N_24016);
nor UO_2919 (O_2919,N_24290,N_24681);
or UO_2920 (O_2920,N_24188,N_24297);
or UO_2921 (O_2921,N_24742,N_24356);
and UO_2922 (O_2922,N_23980,N_24114);
nor UO_2923 (O_2923,N_24127,N_24218);
nand UO_2924 (O_2924,N_24026,N_24693);
nor UO_2925 (O_2925,N_24654,N_24393);
nor UO_2926 (O_2926,N_24499,N_24151);
xor UO_2927 (O_2927,N_24964,N_24052);
and UO_2928 (O_2928,N_24242,N_23813);
or UO_2929 (O_2929,N_24799,N_24668);
and UO_2930 (O_2930,N_23940,N_24864);
or UO_2931 (O_2931,N_24439,N_24297);
xnor UO_2932 (O_2932,N_24675,N_24556);
nor UO_2933 (O_2933,N_24534,N_24721);
nand UO_2934 (O_2934,N_24350,N_24545);
or UO_2935 (O_2935,N_24809,N_24418);
and UO_2936 (O_2936,N_24585,N_24896);
nand UO_2937 (O_2937,N_23811,N_24642);
and UO_2938 (O_2938,N_24222,N_24719);
nand UO_2939 (O_2939,N_24071,N_23772);
and UO_2940 (O_2940,N_24390,N_23988);
xor UO_2941 (O_2941,N_24473,N_23751);
nor UO_2942 (O_2942,N_23852,N_23797);
and UO_2943 (O_2943,N_24758,N_24499);
and UO_2944 (O_2944,N_24705,N_24578);
nor UO_2945 (O_2945,N_23878,N_24786);
nand UO_2946 (O_2946,N_24199,N_24375);
xor UO_2947 (O_2947,N_24164,N_24220);
nand UO_2948 (O_2948,N_23935,N_24230);
nand UO_2949 (O_2949,N_23834,N_24742);
or UO_2950 (O_2950,N_24450,N_24070);
nor UO_2951 (O_2951,N_23783,N_24242);
nor UO_2952 (O_2952,N_24244,N_24687);
or UO_2953 (O_2953,N_23892,N_23998);
and UO_2954 (O_2954,N_24031,N_23902);
nand UO_2955 (O_2955,N_24451,N_23764);
nor UO_2956 (O_2956,N_24082,N_23767);
and UO_2957 (O_2957,N_24460,N_24895);
and UO_2958 (O_2958,N_24454,N_24312);
xnor UO_2959 (O_2959,N_24461,N_24896);
or UO_2960 (O_2960,N_24713,N_23856);
xor UO_2961 (O_2961,N_24603,N_24616);
xor UO_2962 (O_2962,N_23901,N_23802);
nor UO_2963 (O_2963,N_24876,N_24045);
or UO_2964 (O_2964,N_24055,N_23971);
and UO_2965 (O_2965,N_24496,N_24132);
xnor UO_2966 (O_2966,N_24859,N_24252);
nor UO_2967 (O_2967,N_24337,N_24895);
nor UO_2968 (O_2968,N_24529,N_24837);
or UO_2969 (O_2969,N_24456,N_23848);
xnor UO_2970 (O_2970,N_24895,N_23936);
and UO_2971 (O_2971,N_24381,N_24673);
nand UO_2972 (O_2972,N_24470,N_24256);
nor UO_2973 (O_2973,N_24189,N_24967);
xnor UO_2974 (O_2974,N_24856,N_23870);
xnor UO_2975 (O_2975,N_23898,N_23803);
xor UO_2976 (O_2976,N_24111,N_24523);
nor UO_2977 (O_2977,N_24904,N_24281);
nor UO_2978 (O_2978,N_24423,N_24374);
and UO_2979 (O_2979,N_23987,N_23950);
xor UO_2980 (O_2980,N_24249,N_24988);
xnor UO_2981 (O_2981,N_24996,N_24975);
nor UO_2982 (O_2982,N_24401,N_24736);
and UO_2983 (O_2983,N_24640,N_23840);
and UO_2984 (O_2984,N_24130,N_24676);
and UO_2985 (O_2985,N_23797,N_24414);
nand UO_2986 (O_2986,N_23829,N_24613);
nor UO_2987 (O_2987,N_24579,N_24984);
xor UO_2988 (O_2988,N_24599,N_24843);
nand UO_2989 (O_2989,N_24878,N_24194);
xor UO_2990 (O_2990,N_24524,N_24224);
and UO_2991 (O_2991,N_24165,N_24641);
nor UO_2992 (O_2992,N_24301,N_24381);
nor UO_2993 (O_2993,N_23799,N_24590);
nand UO_2994 (O_2994,N_24000,N_23914);
nor UO_2995 (O_2995,N_24318,N_23980);
nand UO_2996 (O_2996,N_23768,N_24729);
nand UO_2997 (O_2997,N_24429,N_23950);
nor UO_2998 (O_2998,N_23931,N_24956);
nor UO_2999 (O_2999,N_24275,N_24590);
endmodule