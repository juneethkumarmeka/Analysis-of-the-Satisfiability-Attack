module basic_750_5000_1000_25_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_153,In_680);
or U1 (N_1,In_459,In_227);
nor U2 (N_2,In_81,In_238);
nor U3 (N_3,In_428,In_75);
or U4 (N_4,In_488,In_491);
nand U5 (N_5,In_155,In_506);
and U6 (N_6,In_531,In_158);
nor U7 (N_7,In_175,In_203);
nand U8 (N_8,In_695,In_749);
nand U9 (N_9,In_598,In_679);
nor U10 (N_10,In_151,In_313);
nand U11 (N_11,In_697,In_576);
or U12 (N_12,In_717,In_88);
and U13 (N_13,In_154,In_431);
and U14 (N_14,In_444,In_245);
nor U15 (N_15,In_324,In_253);
and U16 (N_16,In_264,In_243);
nand U17 (N_17,In_140,In_29);
nand U18 (N_18,In_538,In_737);
and U19 (N_19,In_208,In_720);
nor U20 (N_20,In_494,In_497);
and U21 (N_21,In_12,In_396);
nor U22 (N_22,In_63,In_47);
and U23 (N_23,In_585,In_106);
or U24 (N_24,In_596,In_77);
or U25 (N_25,In_632,In_523);
or U26 (N_26,In_605,In_181);
nand U27 (N_27,In_371,In_277);
or U28 (N_28,In_404,In_621);
and U29 (N_29,In_484,In_511);
and U30 (N_30,In_148,In_220);
or U31 (N_31,In_76,In_685);
xor U32 (N_32,In_687,In_335);
xor U33 (N_33,In_169,In_652);
nor U34 (N_34,In_427,In_378);
or U35 (N_35,In_571,In_212);
nand U36 (N_36,In_211,In_119);
and U37 (N_37,In_664,In_161);
nor U38 (N_38,In_529,In_66);
nor U39 (N_39,In_340,In_495);
or U40 (N_40,In_320,In_422);
xnor U41 (N_41,In_586,In_550);
xnor U42 (N_42,In_65,In_41);
nand U43 (N_43,In_199,In_578);
or U44 (N_44,In_205,In_248);
nor U45 (N_45,In_727,In_403);
xnor U46 (N_46,In_521,In_304);
or U47 (N_47,In_424,In_178);
and U48 (N_48,In_133,In_726);
nor U49 (N_49,In_38,In_156);
or U50 (N_50,In_584,In_625);
nor U51 (N_51,In_646,In_503);
or U52 (N_52,In_676,In_285);
and U53 (N_53,In_310,In_287);
or U54 (N_54,In_630,In_170);
and U55 (N_55,In_244,In_479);
and U56 (N_56,In_555,In_3);
or U57 (N_57,In_37,In_21);
and U58 (N_58,In_61,In_279);
nor U59 (N_59,In_640,In_623);
nor U60 (N_60,In_675,In_163);
or U61 (N_61,In_315,In_684);
nand U62 (N_62,In_711,In_214);
and U63 (N_63,In_272,In_527);
nand U64 (N_64,In_8,In_127);
nand U65 (N_65,In_98,In_415);
or U66 (N_66,In_384,In_182);
nor U67 (N_67,In_510,In_421);
or U68 (N_68,In_271,In_22);
or U69 (N_69,In_296,In_23);
nand U70 (N_70,In_410,In_739);
xnor U71 (N_71,In_267,In_113);
or U72 (N_72,In_554,In_197);
or U73 (N_73,In_202,In_228);
or U74 (N_74,In_455,In_653);
xor U75 (N_75,In_196,In_742);
nand U76 (N_76,In_473,In_641);
xor U77 (N_77,In_1,In_192);
nor U78 (N_78,In_322,In_592);
and U79 (N_79,In_242,In_449);
and U80 (N_80,In_298,In_10);
and U81 (N_81,In_102,In_126);
nand U82 (N_82,In_166,In_651);
or U83 (N_83,In_123,In_412);
nor U84 (N_84,In_704,In_643);
nor U85 (N_85,In_262,In_316);
nand U86 (N_86,In_348,In_594);
nor U87 (N_87,In_505,In_365);
nor U88 (N_88,In_168,In_80);
or U89 (N_89,In_663,In_659);
or U90 (N_90,In_688,In_188);
nor U91 (N_91,In_201,In_468);
and U92 (N_92,In_217,In_683);
nand U93 (N_93,In_662,In_667);
xnor U94 (N_94,In_600,In_474);
nand U95 (N_95,In_707,In_369);
and U96 (N_96,In_144,In_254);
nor U97 (N_97,In_318,In_159);
xnor U98 (N_98,In_177,In_442);
nor U99 (N_99,In_617,In_467);
or U100 (N_100,In_464,In_709);
nor U101 (N_101,In_26,In_317);
and U102 (N_102,In_18,In_581);
and U103 (N_103,In_606,In_291);
and U104 (N_104,In_661,In_432);
and U105 (N_105,In_519,In_402);
or U106 (N_106,In_232,In_388);
or U107 (N_107,In_411,In_526);
nand U108 (N_108,In_545,In_644);
or U109 (N_109,In_380,In_647);
nor U110 (N_110,In_370,In_83);
or U111 (N_111,In_157,In_413);
nor U112 (N_112,In_183,In_678);
or U113 (N_113,In_377,In_485);
or U114 (N_114,In_642,In_109);
or U115 (N_115,In_469,In_284);
nor U116 (N_116,In_376,In_518);
and U117 (N_117,In_286,In_345);
nor U118 (N_118,In_552,In_724);
nor U119 (N_119,In_49,In_231);
or U120 (N_120,In_30,In_557);
and U121 (N_121,In_290,In_604);
or U122 (N_122,In_746,In_307);
xnor U123 (N_123,In_390,In_736);
nor U124 (N_124,In_735,In_562);
and U125 (N_125,In_269,In_560);
or U126 (N_126,In_573,In_533);
or U127 (N_127,In_740,In_57);
xnor U128 (N_128,In_354,In_699);
nor U129 (N_129,In_358,In_62);
and U130 (N_130,In_567,In_616);
nand U131 (N_131,In_2,In_191);
nand U132 (N_132,In_268,In_141);
nor U133 (N_133,In_152,In_420);
or U134 (N_134,In_493,In_624);
or U135 (N_135,In_247,In_86);
or U136 (N_136,In_454,In_64);
nand U137 (N_137,In_569,In_515);
or U138 (N_138,In_574,In_541);
nand U139 (N_139,In_334,In_579);
or U140 (N_140,In_733,In_90);
nand U141 (N_141,In_350,In_120);
nand U142 (N_142,In_629,In_337);
or U143 (N_143,In_397,In_634);
nand U144 (N_144,In_53,In_620);
nand U145 (N_145,In_326,In_463);
nor U146 (N_146,In_351,In_221);
and U147 (N_147,In_280,In_250);
nor U148 (N_148,In_339,In_105);
or U149 (N_149,In_234,In_55);
and U150 (N_150,In_694,In_517);
nor U151 (N_151,In_609,In_648);
nor U152 (N_152,In_512,In_580);
or U153 (N_153,In_429,In_650);
nor U154 (N_154,In_308,In_741);
nand U155 (N_155,In_36,In_138);
or U156 (N_156,In_433,In_568);
and U157 (N_157,In_116,In_558);
nand U158 (N_158,In_261,In_611);
nor U159 (N_159,In_13,In_665);
or U160 (N_160,In_9,In_342);
or U161 (N_161,In_450,In_477);
nor U162 (N_162,In_561,In_721);
or U163 (N_163,In_682,In_82);
nor U164 (N_164,In_300,In_45);
nand U165 (N_165,In_130,In_460);
nand U166 (N_166,In_72,In_146);
nand U167 (N_167,In_564,In_728);
xnor U168 (N_168,In_389,In_173);
nand U169 (N_169,In_343,In_363);
nand U170 (N_170,In_60,In_32);
or U171 (N_171,In_553,In_719);
and U172 (N_172,In_677,In_189);
or U173 (N_173,In_321,In_500);
nor U174 (N_174,In_385,In_597);
xnor U175 (N_175,In_628,In_218);
nor U176 (N_176,In_496,In_548);
nand U177 (N_177,In_332,In_112);
xor U178 (N_178,In_207,In_537);
nand U179 (N_179,In_547,In_626);
or U180 (N_180,In_447,In_627);
and U181 (N_181,In_549,In_686);
or U182 (N_182,In_338,In_54);
nor U183 (N_183,In_84,In_481);
nor U184 (N_184,In_382,In_241);
or U185 (N_185,In_289,In_546);
or U186 (N_186,In_383,In_701);
or U187 (N_187,In_288,In_690);
xnor U188 (N_188,In_336,In_312);
nand U189 (N_189,In_209,In_577);
and U190 (N_190,In_107,In_669);
or U191 (N_191,In_712,In_222);
and U192 (N_192,In_732,In_582);
nor U193 (N_193,In_4,In_543);
nand U194 (N_194,In_591,In_295);
or U195 (N_195,In_160,In_225);
or U196 (N_196,In_118,In_368);
xnor U197 (N_197,In_407,In_35);
or U198 (N_198,In_292,In_430);
nor U199 (N_199,In_11,In_698);
and U200 (N_200,In_492,In_24);
or U201 (N_201,N_137,In_655);
or U202 (N_202,In_645,N_136);
nand U203 (N_203,In_99,In_674);
nand U204 (N_204,N_109,N_134);
nor U205 (N_205,N_142,In_446);
and U206 (N_206,In_150,N_143);
nor U207 (N_207,In_514,N_66);
and U208 (N_208,In_95,In_70);
and U209 (N_209,N_21,In_401);
nand U210 (N_210,In_637,In_235);
or U211 (N_211,In_590,In_507);
and U212 (N_212,In_352,N_153);
and U213 (N_213,In_673,In_39);
nor U214 (N_214,In_48,In_185);
nand U215 (N_215,In_260,In_43);
nand U216 (N_216,In_14,In_25);
nand U217 (N_217,N_155,N_37);
or U218 (N_218,N_107,N_13);
nand U219 (N_219,N_1,N_46);
and U220 (N_220,N_108,In_85);
and U221 (N_221,In_252,In_639);
xnor U222 (N_222,In_17,N_130);
and U223 (N_223,In_456,In_372);
xor U224 (N_224,In_417,N_87);
xor U225 (N_225,In_255,In_516);
nand U226 (N_226,N_38,In_56);
or U227 (N_227,In_213,In_344);
nand U228 (N_228,In_27,N_163);
nand U229 (N_229,In_40,N_7);
or U230 (N_230,In_128,In_619);
nand U231 (N_231,In_306,In_613);
nor U232 (N_232,In_593,N_105);
nor U233 (N_233,In_483,N_39);
xor U234 (N_234,In_349,In_657);
nor U235 (N_235,N_120,In_375);
nand U236 (N_236,In_236,In_730);
or U237 (N_237,In_575,In_210);
nand U238 (N_238,In_301,In_706);
nor U239 (N_239,In_453,In_361);
nor U240 (N_240,N_83,N_9);
xnor U241 (N_241,N_177,N_165);
or U242 (N_242,In_87,In_426);
nor U243 (N_243,In_19,In_360);
nand U244 (N_244,N_74,In_366);
and U245 (N_245,In_165,N_197);
or U246 (N_246,In_565,N_57);
xor U247 (N_247,In_101,N_62);
nand U248 (N_248,In_482,In_583);
nand U249 (N_249,In_52,In_92);
or U250 (N_250,In_251,N_169);
and U251 (N_251,In_249,In_540);
nand U252 (N_252,In_542,In_443);
xnor U253 (N_253,In_722,In_327);
xnor U254 (N_254,N_93,In_636);
xor U255 (N_255,In_656,In_357);
or U256 (N_256,N_26,N_189);
nand U257 (N_257,In_587,In_362);
or U258 (N_258,In_654,In_325);
nand U259 (N_259,In_635,In_374);
and U260 (N_260,In_223,N_126);
or U261 (N_261,In_115,In_530);
or U262 (N_262,In_666,N_2);
xor U263 (N_263,N_170,In_439);
nand U264 (N_264,In_373,In_171);
or U265 (N_265,In_206,N_52);
or U266 (N_266,In_610,In_224);
and U267 (N_267,N_36,In_226);
and U268 (N_268,In_198,In_299);
or U269 (N_269,In_94,N_29);
nand U270 (N_270,N_178,N_30);
nor U271 (N_271,N_35,In_381);
nor U272 (N_272,In_470,In_418);
xor U273 (N_273,In_534,In_89);
nand U274 (N_274,N_190,In_595);
or U275 (N_275,In_747,In_184);
and U276 (N_276,In_341,N_15);
or U277 (N_277,In_186,N_22);
and U278 (N_278,In_311,N_44);
nand U279 (N_279,N_162,In_743);
and U280 (N_280,In_297,N_100);
or U281 (N_281,N_98,In_6);
and U282 (N_282,In_257,N_41);
or U283 (N_283,In_700,N_195);
nor U284 (N_284,N_187,In_117);
nor U285 (N_285,In_392,N_56);
xnor U286 (N_286,In_681,N_65);
nor U287 (N_287,In_34,N_147);
and U288 (N_288,In_607,In_91);
or U289 (N_289,In_745,N_146);
nand U290 (N_290,In_414,N_179);
nor U291 (N_291,In_440,In_303);
and U292 (N_292,In_671,In_615);
or U293 (N_293,N_150,N_71);
or U294 (N_294,In_331,N_180);
nor U295 (N_295,In_504,In_471);
xnor U296 (N_296,In_346,N_72);
or U297 (N_297,In_524,In_475);
or U298 (N_298,In_319,N_67);
or U299 (N_299,In_137,In_16);
and U300 (N_300,N_196,N_45);
nand U301 (N_301,In_716,In_162);
nor U302 (N_302,N_24,In_355);
nand U303 (N_303,N_77,In_535);
and U304 (N_304,In_528,In_180);
xnor U305 (N_305,N_144,N_121);
nand U306 (N_306,In_329,N_50);
nor U307 (N_307,N_139,In_274);
and U308 (N_308,In_559,In_425);
nor U309 (N_309,N_92,In_612);
nand U310 (N_310,In_423,In_658);
and U311 (N_311,In_281,N_184);
and U312 (N_312,N_128,N_43);
and U313 (N_313,N_113,In_419);
and U314 (N_314,In_111,In_451);
xor U315 (N_315,N_19,In_409);
and U316 (N_316,In_710,In_631);
nand U317 (N_317,N_154,In_204);
xnor U318 (N_318,In_614,N_17);
nor U319 (N_319,N_86,N_23);
or U320 (N_320,In_513,In_438);
xnor U321 (N_321,In_237,In_603);
and U322 (N_322,In_406,N_193);
or U323 (N_323,In_129,In_263);
nor U324 (N_324,N_145,In_452);
nand U325 (N_325,In_589,In_435);
nor U326 (N_326,In_149,N_4);
nor U327 (N_327,In_33,In_696);
xor U328 (N_328,In_508,N_40);
and U329 (N_329,N_118,In_708);
and U330 (N_330,In_566,In_333);
xor U331 (N_331,N_182,In_125);
nor U332 (N_332,N_199,In_713);
nor U333 (N_333,In_42,In_142);
nor U334 (N_334,In_59,N_14);
or U335 (N_335,In_556,N_104);
nand U336 (N_336,N_76,N_69);
nand U337 (N_337,In_114,In_104);
nor U338 (N_338,In_15,In_445);
nand U339 (N_339,In_490,N_60);
nand U340 (N_340,N_174,In_330);
nor U341 (N_341,N_129,In_476);
or U342 (N_342,In_347,In_714);
nor U343 (N_343,N_53,In_147);
xnor U344 (N_344,N_186,N_132);
or U345 (N_345,In_572,In_441);
and U346 (N_346,N_125,In_216);
nor U347 (N_347,In_266,In_176);
nand U348 (N_348,In_78,In_246);
or U349 (N_349,In_240,In_744);
nand U350 (N_350,N_168,N_42);
or U351 (N_351,In_164,N_68);
or U352 (N_352,In_44,N_140);
nor U353 (N_353,In_668,In_618);
nand U354 (N_354,In_314,N_122);
and U355 (N_355,N_152,In_174);
or U356 (N_356,N_131,In_705);
nor U357 (N_357,N_102,In_462);
or U358 (N_358,In_398,N_61);
nor U359 (N_359,N_5,In_20);
xnor U360 (N_360,In_588,N_25);
nand U361 (N_361,N_81,In_387);
nor U362 (N_362,N_112,N_89);
nor U363 (N_363,In_601,N_157);
nor U364 (N_364,N_96,N_191);
xnor U365 (N_365,N_176,In_692);
or U366 (N_366,N_85,In_731);
nand U367 (N_367,In_239,In_465);
nor U368 (N_368,In_448,In_97);
nand U369 (N_369,In_273,In_278);
and U370 (N_370,In_145,In_219);
nand U371 (N_371,In_478,N_181);
nor U372 (N_372,In_305,In_364);
and U373 (N_373,In_259,In_436);
or U374 (N_374,In_394,In_122);
xor U375 (N_375,N_18,N_160);
and U376 (N_376,In_400,In_275);
and U377 (N_377,In_525,N_34);
or U378 (N_378,In_660,N_148);
or U379 (N_379,In_434,In_725);
and U380 (N_380,In_50,In_536);
xnor U381 (N_381,In_501,N_138);
nand U382 (N_382,In_489,In_134);
and U383 (N_383,N_171,In_5);
nor U384 (N_384,In_282,N_123);
nand U385 (N_385,In_486,In_103);
xnor U386 (N_386,In_633,N_119);
and U387 (N_387,In_570,N_114);
xor U388 (N_388,N_173,N_158);
nand U389 (N_389,In_520,N_54);
nor U390 (N_390,In_498,In_734);
or U391 (N_391,N_51,N_11);
xor U392 (N_392,In_437,In_71);
and U393 (N_393,In_0,In_622);
and U394 (N_394,In_31,In_723);
nand U395 (N_395,N_0,N_117);
and U396 (N_396,N_79,In_367);
nor U397 (N_397,N_88,N_63);
and U398 (N_398,In_96,N_135);
nor U399 (N_399,In_143,In_79);
or U400 (N_400,N_293,N_239);
and U401 (N_401,N_279,N_302);
nand U402 (N_402,In_748,In_499);
nand U403 (N_403,In_522,In_405);
or U404 (N_404,In_68,N_366);
nor U405 (N_405,N_116,N_318);
and U406 (N_406,N_334,N_398);
and U407 (N_407,N_205,N_75);
or U408 (N_408,N_290,N_359);
nor U409 (N_409,N_356,N_336);
nor U410 (N_410,N_303,N_380);
or U411 (N_411,N_161,N_395);
and U412 (N_412,In_7,N_198);
or U413 (N_413,In_457,N_261);
nor U414 (N_414,N_101,N_355);
and U415 (N_415,In_487,In_715);
and U416 (N_416,N_352,N_339);
and U417 (N_417,N_375,N_327);
or U418 (N_418,N_321,N_320);
nand U419 (N_419,In_172,N_383);
or U420 (N_420,N_222,In_359);
nor U421 (N_421,N_166,N_218);
xnor U422 (N_422,In_28,In_215);
and U423 (N_423,N_8,N_212);
and U424 (N_424,N_360,In_258);
or U425 (N_425,In_539,N_294);
nand U426 (N_426,In_356,N_295);
and U427 (N_427,N_223,In_302);
nand U428 (N_428,In_670,In_276);
nand U429 (N_429,In_738,N_6);
nand U430 (N_430,N_323,In_672);
nor U431 (N_431,N_369,N_207);
nand U432 (N_432,N_90,N_241);
nand U433 (N_433,N_342,N_312);
and U434 (N_434,N_259,N_228);
and U435 (N_435,N_289,N_333);
and U436 (N_436,N_357,N_32);
or U437 (N_437,N_266,N_331);
and U438 (N_438,N_390,N_251);
and U439 (N_439,N_124,In_179);
xnor U440 (N_440,In_132,N_211);
and U441 (N_441,N_221,N_346);
or U442 (N_442,N_291,N_200);
or U443 (N_443,N_167,In_532);
nor U444 (N_444,N_393,N_367);
nor U445 (N_445,N_278,N_203);
or U446 (N_446,N_10,N_365);
and U447 (N_447,N_255,N_265);
or U448 (N_448,N_48,N_80);
or U449 (N_449,N_240,N_285);
nand U450 (N_450,N_236,N_33);
nand U451 (N_451,N_209,N_386);
and U452 (N_452,N_253,N_242);
or U453 (N_453,N_358,N_156);
or U454 (N_454,N_110,N_258);
nor U455 (N_455,N_274,N_273);
nand U456 (N_456,N_192,In_309);
or U457 (N_457,N_311,In_100);
and U458 (N_458,N_340,N_243);
nor U459 (N_459,In_395,In_46);
xor U460 (N_460,N_262,N_382);
nor U461 (N_461,In_458,N_306);
nand U462 (N_462,In_283,N_269);
nand U463 (N_463,In_408,N_206);
and U464 (N_464,In_67,N_208);
and U465 (N_465,N_159,N_376);
nand U466 (N_466,N_73,N_300);
nand U467 (N_467,In_193,N_299);
nor U468 (N_468,N_229,In_69);
nand U469 (N_469,N_250,N_309);
xnor U470 (N_470,In_139,N_319);
or U471 (N_471,N_245,N_377);
nor U472 (N_472,N_283,In_187);
or U473 (N_473,N_99,N_330);
or U474 (N_474,N_263,N_372);
or U475 (N_475,N_111,N_64);
xor U476 (N_476,N_260,In_190);
xnor U477 (N_477,N_97,N_247);
or U478 (N_478,In_136,N_233);
and U479 (N_479,N_397,N_335);
nand U480 (N_480,In_599,N_225);
nand U481 (N_481,In_230,N_348);
and U482 (N_482,N_248,N_213);
and U483 (N_483,In_461,N_349);
nor U484 (N_484,N_378,N_389);
and U485 (N_485,N_310,In_108);
or U486 (N_486,N_338,In_93);
or U487 (N_487,In_703,In_124);
and U488 (N_488,In_393,N_316);
nand U489 (N_489,In_323,N_202);
nand U490 (N_490,N_151,In_265);
and U491 (N_491,N_276,N_361);
and U492 (N_492,N_337,In_110);
nor U493 (N_493,N_55,N_392);
or U494 (N_494,N_371,N_277);
nor U495 (N_495,N_305,N_217);
xor U496 (N_496,N_351,N_298);
and U497 (N_497,N_204,N_313);
nor U498 (N_498,N_149,N_362);
nand U499 (N_499,In_638,N_238);
nor U500 (N_500,N_308,N_275);
nand U501 (N_501,N_82,In_693);
nor U502 (N_502,N_288,N_201);
nor U503 (N_503,N_252,In_718);
and U504 (N_504,N_297,N_133);
and U505 (N_505,N_296,N_264);
nand U506 (N_506,N_194,In_391);
nor U507 (N_507,N_183,N_314);
nor U508 (N_508,N_381,N_370);
xnor U509 (N_509,N_391,N_373);
nand U510 (N_510,N_175,N_249);
or U511 (N_511,N_215,In_58);
nand U512 (N_512,In_73,N_216);
nand U513 (N_513,In_729,N_384);
nand U514 (N_514,In_649,N_210);
nand U515 (N_515,N_394,N_246);
or U516 (N_516,N_399,N_324);
nor U517 (N_517,N_234,N_315);
or U518 (N_518,N_329,N_28);
or U519 (N_519,N_115,N_20);
and U520 (N_520,N_284,N_281);
or U521 (N_521,N_94,N_304);
nor U522 (N_522,N_254,N_343);
and U523 (N_523,N_31,In_379);
xor U524 (N_524,In_466,N_244);
or U525 (N_525,N_185,In_270);
nor U526 (N_526,N_332,In_386);
xnor U527 (N_527,N_95,N_231);
and U528 (N_528,In_195,N_282);
xnor U529 (N_529,In_121,In_551);
and U530 (N_530,N_287,N_280);
nor U531 (N_531,In_74,In_256);
nor U532 (N_532,N_353,In_131);
and U533 (N_533,N_127,N_214);
and U534 (N_534,N_301,N_388);
nor U535 (N_535,N_141,N_286);
xnor U536 (N_536,N_224,N_47);
or U537 (N_537,In_194,N_226);
or U538 (N_538,In_167,N_270);
xnor U539 (N_539,N_322,In_480);
or U540 (N_540,N_220,N_317);
nor U541 (N_541,In_293,N_84);
nor U542 (N_542,In_51,In_544);
nand U543 (N_543,N_70,In_135);
nor U544 (N_544,N_385,N_106);
or U545 (N_545,N_374,N_172);
and U546 (N_546,N_256,In_233);
nand U547 (N_547,In_399,N_268);
xnor U548 (N_548,N_307,N_292);
or U549 (N_549,In_416,N_363);
nand U550 (N_550,N_219,N_232);
and U551 (N_551,In_353,N_257);
and U552 (N_552,N_341,N_344);
and U553 (N_553,In_689,In_563);
or U554 (N_554,N_164,N_364);
nor U555 (N_555,N_272,In_702);
and U556 (N_556,N_227,N_354);
and U557 (N_557,In_502,In_328);
and U558 (N_558,N_91,N_188);
nand U559 (N_559,N_16,N_326);
and U560 (N_560,N_3,In_200);
nor U561 (N_561,In_691,N_350);
and U562 (N_562,N_325,N_347);
nand U563 (N_563,N_58,N_235);
nand U564 (N_564,In_509,N_27);
nor U565 (N_565,N_379,N_230);
nor U566 (N_566,N_78,N_12);
nand U567 (N_567,N_49,N_271);
xor U568 (N_568,N_387,N_345);
or U569 (N_569,In_602,N_103);
nor U570 (N_570,In_472,N_237);
and U571 (N_571,N_396,N_267);
nor U572 (N_572,N_368,N_59);
nor U573 (N_573,In_608,N_328);
or U574 (N_574,In_229,In_294);
nor U575 (N_575,N_236,N_328);
and U576 (N_576,N_360,N_238);
nor U577 (N_577,N_286,In_472);
and U578 (N_578,In_328,N_214);
nand U579 (N_579,N_262,In_703);
nor U580 (N_580,N_305,N_260);
and U581 (N_581,N_233,N_301);
and U582 (N_582,N_3,N_308);
and U583 (N_583,In_457,N_369);
or U584 (N_584,N_371,N_322);
and U585 (N_585,N_296,N_377);
nor U586 (N_586,In_480,N_166);
or U587 (N_587,In_256,N_315);
and U588 (N_588,In_193,N_391);
or U589 (N_589,N_382,N_185);
nand U590 (N_590,In_393,In_748);
nand U591 (N_591,N_8,N_320);
and U592 (N_592,N_300,N_213);
and U593 (N_593,N_159,N_194);
nor U594 (N_594,In_136,In_703);
nor U595 (N_595,N_309,In_28);
nand U596 (N_596,N_251,N_267);
and U597 (N_597,N_245,N_32);
xor U598 (N_598,N_354,N_221);
and U599 (N_599,N_238,In_323);
or U600 (N_600,N_490,N_415);
nand U601 (N_601,N_428,N_568);
or U602 (N_602,N_565,N_404);
and U603 (N_603,N_432,N_527);
nand U604 (N_604,N_400,N_491);
nand U605 (N_605,N_480,N_475);
or U606 (N_606,N_533,N_406);
nor U607 (N_607,N_586,N_592);
nand U608 (N_608,N_547,N_517);
and U609 (N_609,N_467,N_401);
or U610 (N_610,N_419,N_455);
or U611 (N_611,N_456,N_536);
and U612 (N_612,N_458,N_555);
or U613 (N_613,N_405,N_510);
nor U614 (N_614,N_512,N_439);
or U615 (N_615,N_521,N_546);
nor U616 (N_616,N_500,N_588);
or U617 (N_617,N_449,N_561);
and U618 (N_618,N_402,N_548);
or U619 (N_619,N_539,N_461);
nand U620 (N_620,N_462,N_424);
or U621 (N_621,N_532,N_516);
nor U622 (N_622,N_545,N_552);
xnor U623 (N_623,N_454,N_493);
nand U624 (N_624,N_412,N_421);
and U625 (N_625,N_478,N_465);
or U626 (N_626,N_571,N_436);
nor U627 (N_627,N_523,N_530);
or U628 (N_628,N_472,N_537);
nor U629 (N_629,N_488,N_410);
nand U630 (N_630,N_469,N_473);
nand U631 (N_631,N_508,N_446);
nor U632 (N_632,N_515,N_594);
nand U633 (N_633,N_471,N_435);
xor U634 (N_634,N_535,N_427);
or U635 (N_635,N_474,N_443);
and U636 (N_636,N_556,N_595);
and U637 (N_637,N_418,N_489);
nand U638 (N_638,N_431,N_598);
or U639 (N_639,N_587,N_577);
and U640 (N_640,N_584,N_483);
nand U641 (N_641,N_549,N_524);
xor U642 (N_642,N_416,N_422);
nor U643 (N_643,N_440,N_433);
nand U644 (N_644,N_509,N_420);
and U645 (N_645,N_486,N_560);
nand U646 (N_646,N_466,N_447);
and U647 (N_647,N_408,N_558);
nand U648 (N_648,N_581,N_429);
and U649 (N_649,N_506,N_413);
or U650 (N_650,N_477,N_526);
nand U651 (N_651,N_573,N_554);
nor U652 (N_652,N_505,N_460);
or U653 (N_653,N_514,N_569);
xor U654 (N_654,N_593,N_572);
nand U655 (N_655,N_525,N_452);
nor U656 (N_656,N_541,N_599);
nand U657 (N_657,N_528,N_417);
and U658 (N_658,N_459,N_559);
and U659 (N_659,N_448,N_513);
nand U660 (N_660,N_450,N_597);
nand U661 (N_661,N_485,N_591);
and U662 (N_662,N_502,N_468);
or U663 (N_663,N_564,N_563);
nand U664 (N_664,N_476,N_457);
nor U665 (N_665,N_518,N_438);
nand U666 (N_666,N_426,N_482);
nand U667 (N_667,N_534,N_425);
nand U668 (N_668,N_590,N_423);
nand U669 (N_669,N_562,N_570);
or U670 (N_670,N_445,N_540);
or U671 (N_671,N_411,N_583);
nand U672 (N_672,N_492,N_495);
and U673 (N_673,N_441,N_538);
nand U674 (N_674,N_543,N_553);
nand U675 (N_675,N_503,N_487);
nand U676 (N_676,N_578,N_437);
or U677 (N_677,N_585,N_403);
or U678 (N_678,N_407,N_575);
and U679 (N_679,N_504,N_507);
or U680 (N_680,N_580,N_519);
or U681 (N_681,N_497,N_566);
nand U682 (N_682,N_501,N_464);
or U683 (N_683,N_511,N_442);
and U684 (N_684,N_531,N_589);
nand U685 (N_685,N_414,N_550);
nor U686 (N_686,N_582,N_576);
and U687 (N_687,N_409,N_522);
and U688 (N_688,N_444,N_596);
and U689 (N_689,N_496,N_451);
and U690 (N_690,N_463,N_529);
nor U691 (N_691,N_481,N_567);
nor U692 (N_692,N_430,N_453);
nor U693 (N_693,N_498,N_434);
and U694 (N_694,N_484,N_579);
nor U695 (N_695,N_499,N_551);
nor U696 (N_696,N_557,N_470);
or U697 (N_697,N_574,N_544);
nand U698 (N_698,N_520,N_542);
or U699 (N_699,N_494,N_479);
nor U700 (N_700,N_488,N_597);
and U701 (N_701,N_570,N_440);
and U702 (N_702,N_508,N_473);
or U703 (N_703,N_558,N_424);
and U704 (N_704,N_408,N_401);
or U705 (N_705,N_402,N_448);
nand U706 (N_706,N_481,N_595);
nor U707 (N_707,N_522,N_540);
nor U708 (N_708,N_451,N_533);
nor U709 (N_709,N_492,N_448);
nor U710 (N_710,N_459,N_509);
or U711 (N_711,N_549,N_429);
or U712 (N_712,N_573,N_455);
nor U713 (N_713,N_480,N_463);
nor U714 (N_714,N_495,N_413);
and U715 (N_715,N_485,N_564);
nand U716 (N_716,N_484,N_456);
nand U717 (N_717,N_479,N_554);
and U718 (N_718,N_441,N_412);
xnor U719 (N_719,N_516,N_430);
nor U720 (N_720,N_449,N_570);
nand U721 (N_721,N_412,N_415);
nand U722 (N_722,N_428,N_593);
xor U723 (N_723,N_406,N_544);
and U724 (N_724,N_545,N_478);
and U725 (N_725,N_531,N_459);
or U726 (N_726,N_403,N_523);
and U727 (N_727,N_553,N_562);
nor U728 (N_728,N_501,N_422);
nor U729 (N_729,N_509,N_498);
nand U730 (N_730,N_462,N_421);
or U731 (N_731,N_406,N_448);
xor U732 (N_732,N_445,N_554);
xor U733 (N_733,N_570,N_496);
nor U734 (N_734,N_432,N_468);
or U735 (N_735,N_459,N_410);
and U736 (N_736,N_580,N_564);
and U737 (N_737,N_498,N_574);
or U738 (N_738,N_430,N_592);
and U739 (N_739,N_414,N_466);
or U740 (N_740,N_530,N_471);
and U741 (N_741,N_402,N_463);
or U742 (N_742,N_472,N_545);
or U743 (N_743,N_507,N_555);
nand U744 (N_744,N_435,N_479);
nand U745 (N_745,N_582,N_476);
nand U746 (N_746,N_454,N_451);
nor U747 (N_747,N_487,N_584);
and U748 (N_748,N_582,N_575);
and U749 (N_749,N_461,N_535);
or U750 (N_750,N_491,N_465);
nand U751 (N_751,N_417,N_414);
nand U752 (N_752,N_592,N_481);
nor U753 (N_753,N_443,N_594);
or U754 (N_754,N_423,N_498);
nor U755 (N_755,N_572,N_504);
or U756 (N_756,N_423,N_488);
xor U757 (N_757,N_595,N_501);
or U758 (N_758,N_488,N_534);
nor U759 (N_759,N_427,N_575);
and U760 (N_760,N_523,N_559);
and U761 (N_761,N_477,N_530);
nand U762 (N_762,N_547,N_504);
nor U763 (N_763,N_541,N_443);
nand U764 (N_764,N_406,N_433);
nand U765 (N_765,N_533,N_560);
and U766 (N_766,N_588,N_418);
or U767 (N_767,N_576,N_540);
xor U768 (N_768,N_535,N_466);
nand U769 (N_769,N_405,N_491);
or U770 (N_770,N_529,N_574);
and U771 (N_771,N_498,N_400);
and U772 (N_772,N_460,N_549);
nand U773 (N_773,N_439,N_513);
or U774 (N_774,N_599,N_527);
nand U775 (N_775,N_452,N_584);
and U776 (N_776,N_441,N_509);
or U777 (N_777,N_573,N_418);
xnor U778 (N_778,N_596,N_474);
nand U779 (N_779,N_410,N_496);
nor U780 (N_780,N_586,N_403);
nand U781 (N_781,N_423,N_463);
nand U782 (N_782,N_492,N_513);
and U783 (N_783,N_487,N_486);
xor U784 (N_784,N_490,N_502);
and U785 (N_785,N_522,N_577);
and U786 (N_786,N_472,N_483);
and U787 (N_787,N_577,N_597);
or U788 (N_788,N_493,N_536);
nor U789 (N_789,N_519,N_492);
xnor U790 (N_790,N_554,N_522);
nand U791 (N_791,N_460,N_407);
xnor U792 (N_792,N_587,N_421);
xnor U793 (N_793,N_487,N_431);
nand U794 (N_794,N_508,N_414);
nor U795 (N_795,N_543,N_516);
nor U796 (N_796,N_449,N_543);
or U797 (N_797,N_428,N_519);
nor U798 (N_798,N_576,N_562);
nor U799 (N_799,N_559,N_430);
nor U800 (N_800,N_752,N_635);
xnor U801 (N_801,N_704,N_611);
nor U802 (N_802,N_764,N_692);
nor U803 (N_803,N_732,N_705);
nor U804 (N_804,N_790,N_625);
nand U805 (N_805,N_601,N_776);
or U806 (N_806,N_673,N_617);
nand U807 (N_807,N_722,N_773);
nand U808 (N_808,N_682,N_686);
or U809 (N_809,N_766,N_636);
nor U810 (N_810,N_640,N_747);
or U811 (N_811,N_654,N_794);
and U812 (N_812,N_628,N_795);
or U813 (N_813,N_656,N_700);
or U814 (N_814,N_717,N_727);
nand U815 (N_815,N_624,N_677);
and U816 (N_816,N_612,N_756);
xor U817 (N_817,N_749,N_769);
nand U818 (N_818,N_706,N_622);
and U819 (N_819,N_602,N_641);
nor U820 (N_820,N_608,N_650);
and U821 (N_821,N_707,N_751);
xor U822 (N_822,N_607,N_634);
and U823 (N_823,N_652,N_685);
nor U824 (N_824,N_672,N_712);
nand U825 (N_825,N_689,N_694);
xor U826 (N_826,N_718,N_770);
nand U827 (N_827,N_683,N_796);
nand U828 (N_828,N_719,N_642);
nand U829 (N_829,N_765,N_731);
nand U830 (N_830,N_605,N_755);
nand U831 (N_831,N_775,N_799);
and U832 (N_832,N_681,N_716);
nor U833 (N_833,N_753,N_737);
or U834 (N_834,N_779,N_783);
and U835 (N_835,N_629,N_788);
nor U836 (N_836,N_789,N_745);
nand U837 (N_837,N_646,N_670);
or U838 (N_838,N_709,N_697);
and U839 (N_839,N_758,N_649);
nand U840 (N_840,N_698,N_734);
and U841 (N_841,N_678,N_610);
xnor U842 (N_842,N_708,N_777);
nor U843 (N_843,N_637,N_699);
nor U844 (N_844,N_623,N_653);
and U845 (N_845,N_664,N_633);
or U846 (N_846,N_696,N_760);
or U847 (N_847,N_713,N_669);
nand U848 (N_848,N_667,N_632);
or U849 (N_849,N_780,N_771);
nand U850 (N_850,N_657,N_703);
or U851 (N_851,N_781,N_750);
nor U852 (N_852,N_651,N_792);
nand U853 (N_853,N_620,N_786);
or U854 (N_854,N_680,N_687);
xnor U855 (N_855,N_720,N_658);
or U856 (N_856,N_711,N_726);
xnor U857 (N_857,N_659,N_695);
nor U858 (N_858,N_782,N_600);
or U859 (N_859,N_631,N_725);
nand U860 (N_860,N_744,N_645);
and U861 (N_861,N_644,N_663);
nand U862 (N_862,N_778,N_754);
or U863 (N_863,N_728,N_742);
or U864 (N_864,N_748,N_741);
and U865 (N_865,N_660,N_768);
xor U866 (N_866,N_714,N_662);
nand U867 (N_867,N_784,N_626);
nand U868 (N_868,N_688,N_691);
and U869 (N_869,N_693,N_740);
nor U870 (N_870,N_702,N_774);
or U871 (N_871,N_613,N_666);
and U872 (N_872,N_798,N_739);
and U873 (N_873,N_616,N_647);
and U874 (N_874,N_648,N_746);
or U875 (N_875,N_767,N_723);
nor U876 (N_876,N_603,N_724);
nor U877 (N_877,N_630,N_733);
nor U878 (N_878,N_615,N_761);
nor U879 (N_879,N_762,N_643);
or U880 (N_880,N_797,N_675);
and U881 (N_881,N_618,N_791);
or U882 (N_882,N_787,N_619);
or U883 (N_883,N_638,N_772);
nand U884 (N_884,N_710,N_671);
nor U885 (N_885,N_674,N_609);
and U886 (N_886,N_743,N_684);
nor U887 (N_887,N_763,N_721);
or U888 (N_888,N_759,N_627);
xnor U889 (N_889,N_665,N_730);
nand U890 (N_890,N_757,N_793);
and U891 (N_891,N_639,N_735);
nor U892 (N_892,N_701,N_736);
or U893 (N_893,N_614,N_729);
nand U894 (N_894,N_690,N_655);
or U895 (N_895,N_621,N_661);
and U896 (N_896,N_606,N_668);
nand U897 (N_897,N_715,N_785);
and U898 (N_898,N_676,N_738);
or U899 (N_899,N_604,N_679);
nand U900 (N_900,N_613,N_769);
and U901 (N_901,N_679,N_747);
nor U902 (N_902,N_785,N_792);
or U903 (N_903,N_639,N_616);
and U904 (N_904,N_748,N_777);
nor U905 (N_905,N_725,N_679);
and U906 (N_906,N_793,N_789);
and U907 (N_907,N_789,N_625);
nor U908 (N_908,N_731,N_673);
or U909 (N_909,N_692,N_644);
nand U910 (N_910,N_607,N_758);
and U911 (N_911,N_689,N_772);
and U912 (N_912,N_720,N_655);
or U913 (N_913,N_628,N_679);
or U914 (N_914,N_610,N_685);
or U915 (N_915,N_653,N_646);
and U916 (N_916,N_781,N_664);
and U917 (N_917,N_708,N_709);
nor U918 (N_918,N_763,N_737);
nor U919 (N_919,N_603,N_689);
nand U920 (N_920,N_743,N_774);
xor U921 (N_921,N_625,N_798);
nor U922 (N_922,N_600,N_679);
nand U923 (N_923,N_778,N_701);
or U924 (N_924,N_670,N_700);
and U925 (N_925,N_612,N_723);
or U926 (N_926,N_668,N_622);
and U927 (N_927,N_789,N_785);
and U928 (N_928,N_701,N_764);
nand U929 (N_929,N_644,N_615);
nor U930 (N_930,N_776,N_786);
or U931 (N_931,N_699,N_735);
or U932 (N_932,N_628,N_797);
and U933 (N_933,N_632,N_753);
xor U934 (N_934,N_794,N_706);
or U935 (N_935,N_744,N_600);
nor U936 (N_936,N_785,N_625);
and U937 (N_937,N_757,N_783);
and U938 (N_938,N_711,N_600);
nor U939 (N_939,N_604,N_756);
xnor U940 (N_940,N_613,N_700);
or U941 (N_941,N_670,N_775);
nor U942 (N_942,N_774,N_657);
nor U943 (N_943,N_723,N_769);
nand U944 (N_944,N_660,N_763);
nand U945 (N_945,N_687,N_780);
nor U946 (N_946,N_661,N_636);
and U947 (N_947,N_798,N_624);
and U948 (N_948,N_608,N_633);
nand U949 (N_949,N_710,N_608);
nor U950 (N_950,N_782,N_677);
nor U951 (N_951,N_711,N_605);
nor U952 (N_952,N_744,N_793);
nor U953 (N_953,N_654,N_644);
and U954 (N_954,N_796,N_670);
nand U955 (N_955,N_707,N_637);
and U956 (N_956,N_611,N_736);
or U957 (N_957,N_787,N_627);
nand U958 (N_958,N_734,N_757);
or U959 (N_959,N_657,N_608);
nand U960 (N_960,N_657,N_779);
or U961 (N_961,N_706,N_775);
nor U962 (N_962,N_613,N_630);
or U963 (N_963,N_632,N_747);
and U964 (N_964,N_741,N_665);
and U965 (N_965,N_747,N_704);
or U966 (N_966,N_675,N_601);
xnor U967 (N_967,N_711,N_695);
and U968 (N_968,N_613,N_685);
nor U969 (N_969,N_718,N_799);
or U970 (N_970,N_696,N_658);
and U971 (N_971,N_672,N_617);
nor U972 (N_972,N_735,N_659);
or U973 (N_973,N_748,N_781);
nor U974 (N_974,N_734,N_703);
nor U975 (N_975,N_681,N_688);
or U976 (N_976,N_781,N_600);
xnor U977 (N_977,N_797,N_658);
xor U978 (N_978,N_657,N_683);
nor U979 (N_979,N_752,N_648);
and U980 (N_980,N_659,N_779);
or U981 (N_981,N_639,N_648);
and U982 (N_982,N_603,N_642);
and U983 (N_983,N_784,N_669);
nor U984 (N_984,N_685,N_677);
nor U985 (N_985,N_651,N_781);
and U986 (N_986,N_741,N_646);
and U987 (N_987,N_730,N_671);
nand U988 (N_988,N_614,N_690);
or U989 (N_989,N_605,N_619);
and U990 (N_990,N_797,N_791);
and U991 (N_991,N_635,N_681);
or U992 (N_992,N_692,N_630);
nand U993 (N_993,N_601,N_772);
xor U994 (N_994,N_784,N_745);
xor U995 (N_995,N_660,N_713);
nor U996 (N_996,N_784,N_742);
or U997 (N_997,N_610,N_621);
nand U998 (N_998,N_706,N_753);
nand U999 (N_999,N_739,N_751);
nor U1000 (N_1000,N_870,N_930);
nor U1001 (N_1001,N_932,N_892);
nand U1002 (N_1002,N_884,N_885);
nor U1003 (N_1003,N_924,N_819);
and U1004 (N_1004,N_837,N_897);
nor U1005 (N_1005,N_842,N_940);
nor U1006 (N_1006,N_939,N_821);
nor U1007 (N_1007,N_971,N_989);
nor U1008 (N_1008,N_984,N_933);
xnor U1009 (N_1009,N_905,N_805);
xor U1010 (N_1010,N_813,N_832);
xnor U1011 (N_1011,N_979,N_891);
nand U1012 (N_1012,N_972,N_879);
nand U1013 (N_1013,N_800,N_993);
xnor U1014 (N_1014,N_886,N_852);
nor U1015 (N_1015,N_834,N_880);
nand U1016 (N_1016,N_906,N_882);
and U1017 (N_1017,N_858,N_955);
nand U1018 (N_1018,N_961,N_969);
nor U1019 (N_1019,N_823,N_839);
or U1020 (N_1020,N_902,N_857);
nor U1021 (N_1021,N_991,N_845);
nor U1022 (N_1022,N_822,N_992);
or U1023 (N_1023,N_937,N_854);
nand U1024 (N_1024,N_878,N_921);
or U1025 (N_1025,N_847,N_871);
or U1026 (N_1026,N_910,N_987);
or U1027 (N_1027,N_954,N_964);
nand U1028 (N_1028,N_913,N_966);
xor U1029 (N_1029,N_928,N_908);
nor U1030 (N_1030,N_840,N_869);
or U1031 (N_1031,N_986,N_807);
and U1032 (N_1032,N_835,N_808);
xnor U1033 (N_1033,N_960,N_948);
or U1034 (N_1034,N_904,N_967);
or U1035 (N_1035,N_877,N_963);
xnor U1036 (N_1036,N_846,N_945);
or U1037 (N_1037,N_912,N_812);
and U1038 (N_1038,N_836,N_936);
nor U1039 (N_1039,N_889,N_953);
xnor U1040 (N_1040,N_856,N_959);
or U1041 (N_1041,N_962,N_872);
and U1042 (N_1042,N_820,N_825);
xnor U1043 (N_1043,N_965,N_848);
and U1044 (N_1044,N_853,N_818);
or U1045 (N_1045,N_950,N_866);
xor U1046 (N_1046,N_922,N_975);
xor U1047 (N_1047,N_918,N_816);
or U1048 (N_1048,N_983,N_914);
and U1049 (N_1049,N_894,N_899);
or U1050 (N_1050,N_881,N_935);
nor U1051 (N_1051,N_873,N_981);
and U1052 (N_1052,N_990,N_801);
nor U1053 (N_1053,N_985,N_943);
nand U1054 (N_1054,N_977,N_810);
nand U1055 (N_1055,N_968,N_827);
or U1056 (N_1056,N_850,N_802);
nor U1057 (N_1057,N_951,N_806);
nand U1058 (N_1058,N_829,N_925);
and U1059 (N_1059,N_864,N_920);
nor U1060 (N_1060,N_976,N_849);
and U1061 (N_1061,N_863,N_901);
nor U1062 (N_1062,N_824,N_978);
nor U1063 (N_1063,N_844,N_952);
nor U1064 (N_1064,N_828,N_941);
xor U1065 (N_1065,N_907,N_817);
and U1066 (N_1066,N_900,N_815);
and U1067 (N_1067,N_804,N_917);
or U1068 (N_1068,N_927,N_874);
xor U1069 (N_1069,N_944,N_949);
nand U1070 (N_1070,N_909,N_970);
or U1071 (N_1071,N_898,N_833);
nand U1072 (N_1072,N_929,N_860);
and U1073 (N_1073,N_838,N_926);
nand U1074 (N_1074,N_931,N_890);
nand U1075 (N_1075,N_916,N_974);
nand U1076 (N_1076,N_859,N_868);
nand U1077 (N_1077,N_919,N_994);
xor U1078 (N_1078,N_946,N_887);
xnor U1079 (N_1079,N_811,N_999);
or U1080 (N_1080,N_867,N_843);
nand U1081 (N_1081,N_982,N_814);
nand U1082 (N_1082,N_911,N_915);
and U1083 (N_1083,N_956,N_995);
nor U1084 (N_1084,N_923,N_862);
nor U1085 (N_1085,N_809,N_861);
xnor U1086 (N_1086,N_803,N_855);
and U1087 (N_1087,N_973,N_895);
and U1088 (N_1088,N_831,N_938);
and U1089 (N_1089,N_998,N_958);
nor U1090 (N_1090,N_942,N_826);
xnor U1091 (N_1091,N_875,N_997);
nor U1092 (N_1092,N_851,N_988);
xnor U1093 (N_1093,N_883,N_947);
or U1094 (N_1094,N_830,N_934);
nand U1095 (N_1095,N_996,N_841);
and U1096 (N_1096,N_980,N_957);
or U1097 (N_1097,N_876,N_903);
nand U1098 (N_1098,N_888,N_896);
and U1099 (N_1099,N_865,N_893);
and U1100 (N_1100,N_803,N_824);
nand U1101 (N_1101,N_842,N_815);
or U1102 (N_1102,N_955,N_926);
nand U1103 (N_1103,N_807,N_813);
nand U1104 (N_1104,N_929,N_851);
nand U1105 (N_1105,N_895,N_890);
nand U1106 (N_1106,N_904,N_940);
xnor U1107 (N_1107,N_864,N_882);
nor U1108 (N_1108,N_939,N_929);
nand U1109 (N_1109,N_846,N_940);
nor U1110 (N_1110,N_923,N_947);
xor U1111 (N_1111,N_843,N_969);
and U1112 (N_1112,N_860,N_864);
xor U1113 (N_1113,N_979,N_872);
nor U1114 (N_1114,N_967,N_858);
nand U1115 (N_1115,N_978,N_992);
nor U1116 (N_1116,N_968,N_965);
and U1117 (N_1117,N_943,N_910);
or U1118 (N_1118,N_950,N_940);
or U1119 (N_1119,N_958,N_986);
or U1120 (N_1120,N_845,N_875);
or U1121 (N_1121,N_855,N_917);
or U1122 (N_1122,N_852,N_946);
nand U1123 (N_1123,N_959,N_843);
nor U1124 (N_1124,N_932,N_851);
or U1125 (N_1125,N_847,N_908);
nor U1126 (N_1126,N_915,N_824);
nand U1127 (N_1127,N_973,N_962);
and U1128 (N_1128,N_915,N_870);
or U1129 (N_1129,N_914,N_825);
or U1130 (N_1130,N_972,N_918);
and U1131 (N_1131,N_999,N_823);
xor U1132 (N_1132,N_951,N_893);
and U1133 (N_1133,N_852,N_828);
or U1134 (N_1134,N_800,N_962);
or U1135 (N_1135,N_964,N_826);
nor U1136 (N_1136,N_883,N_802);
and U1137 (N_1137,N_967,N_832);
and U1138 (N_1138,N_913,N_953);
and U1139 (N_1139,N_886,N_802);
or U1140 (N_1140,N_839,N_902);
nand U1141 (N_1141,N_921,N_992);
nor U1142 (N_1142,N_970,N_898);
nand U1143 (N_1143,N_916,N_859);
nor U1144 (N_1144,N_996,N_937);
nand U1145 (N_1145,N_895,N_823);
xnor U1146 (N_1146,N_856,N_980);
or U1147 (N_1147,N_962,N_897);
and U1148 (N_1148,N_825,N_922);
or U1149 (N_1149,N_861,N_896);
nand U1150 (N_1150,N_910,N_971);
xor U1151 (N_1151,N_965,N_802);
or U1152 (N_1152,N_960,N_889);
nand U1153 (N_1153,N_886,N_920);
nand U1154 (N_1154,N_923,N_890);
nand U1155 (N_1155,N_968,N_896);
xor U1156 (N_1156,N_922,N_918);
and U1157 (N_1157,N_994,N_981);
nor U1158 (N_1158,N_867,N_914);
and U1159 (N_1159,N_816,N_808);
and U1160 (N_1160,N_956,N_916);
xor U1161 (N_1161,N_968,N_831);
or U1162 (N_1162,N_969,N_908);
or U1163 (N_1163,N_821,N_868);
or U1164 (N_1164,N_967,N_909);
or U1165 (N_1165,N_860,N_981);
nor U1166 (N_1166,N_892,N_947);
xor U1167 (N_1167,N_965,N_844);
nand U1168 (N_1168,N_830,N_954);
nand U1169 (N_1169,N_802,N_846);
and U1170 (N_1170,N_820,N_973);
or U1171 (N_1171,N_832,N_853);
and U1172 (N_1172,N_945,N_986);
and U1173 (N_1173,N_834,N_959);
nor U1174 (N_1174,N_889,N_958);
nand U1175 (N_1175,N_923,N_873);
nor U1176 (N_1176,N_947,N_806);
or U1177 (N_1177,N_996,N_883);
nand U1178 (N_1178,N_971,N_975);
nand U1179 (N_1179,N_997,N_960);
nor U1180 (N_1180,N_909,N_845);
and U1181 (N_1181,N_827,N_890);
nor U1182 (N_1182,N_850,N_843);
nor U1183 (N_1183,N_925,N_862);
nand U1184 (N_1184,N_895,N_819);
and U1185 (N_1185,N_898,N_882);
nand U1186 (N_1186,N_967,N_864);
or U1187 (N_1187,N_882,N_913);
xnor U1188 (N_1188,N_925,N_823);
nor U1189 (N_1189,N_892,N_926);
and U1190 (N_1190,N_872,N_863);
and U1191 (N_1191,N_870,N_925);
nand U1192 (N_1192,N_846,N_929);
nand U1193 (N_1193,N_809,N_957);
or U1194 (N_1194,N_929,N_813);
or U1195 (N_1195,N_820,N_907);
and U1196 (N_1196,N_828,N_836);
xnor U1197 (N_1197,N_943,N_999);
xor U1198 (N_1198,N_912,N_931);
nand U1199 (N_1199,N_862,N_909);
nor U1200 (N_1200,N_1105,N_1095);
or U1201 (N_1201,N_1092,N_1050);
or U1202 (N_1202,N_1087,N_1172);
nand U1203 (N_1203,N_1063,N_1110);
nor U1204 (N_1204,N_1102,N_1041);
nor U1205 (N_1205,N_1123,N_1182);
nand U1206 (N_1206,N_1146,N_1009);
xnor U1207 (N_1207,N_1066,N_1003);
and U1208 (N_1208,N_1178,N_1056);
nor U1209 (N_1209,N_1001,N_1120);
or U1210 (N_1210,N_1010,N_1164);
or U1211 (N_1211,N_1059,N_1030);
nand U1212 (N_1212,N_1000,N_1167);
nor U1213 (N_1213,N_1155,N_1015);
nor U1214 (N_1214,N_1049,N_1073);
nand U1215 (N_1215,N_1067,N_1012);
nand U1216 (N_1216,N_1014,N_1038);
xor U1217 (N_1217,N_1079,N_1171);
and U1218 (N_1218,N_1083,N_1057);
nand U1219 (N_1219,N_1132,N_1185);
or U1220 (N_1220,N_1062,N_1039);
nor U1221 (N_1221,N_1091,N_1197);
nor U1222 (N_1222,N_1198,N_1168);
nor U1223 (N_1223,N_1187,N_1036);
nor U1224 (N_1224,N_1128,N_1138);
and U1225 (N_1225,N_1133,N_1069);
nor U1226 (N_1226,N_1002,N_1189);
and U1227 (N_1227,N_1107,N_1031);
and U1228 (N_1228,N_1124,N_1076);
nor U1229 (N_1229,N_1019,N_1137);
and U1230 (N_1230,N_1125,N_1080);
xor U1231 (N_1231,N_1111,N_1175);
or U1232 (N_1232,N_1174,N_1090);
or U1233 (N_1233,N_1195,N_1068);
or U1234 (N_1234,N_1145,N_1074);
and U1235 (N_1235,N_1103,N_1005);
and U1236 (N_1236,N_1159,N_1058);
nand U1237 (N_1237,N_1046,N_1109);
or U1238 (N_1238,N_1144,N_1011);
nand U1239 (N_1239,N_1104,N_1013);
nor U1240 (N_1240,N_1027,N_1122);
nor U1241 (N_1241,N_1096,N_1154);
nand U1242 (N_1242,N_1165,N_1173);
and U1243 (N_1243,N_1190,N_1177);
xor U1244 (N_1244,N_1147,N_1152);
nor U1245 (N_1245,N_1037,N_1196);
or U1246 (N_1246,N_1184,N_1034);
xor U1247 (N_1247,N_1193,N_1112);
and U1248 (N_1248,N_1061,N_1020);
nand U1249 (N_1249,N_1054,N_1022);
nand U1250 (N_1250,N_1028,N_1108);
nand U1251 (N_1251,N_1141,N_1176);
nand U1252 (N_1252,N_1181,N_1191);
xor U1253 (N_1253,N_1126,N_1053);
nand U1254 (N_1254,N_1071,N_1089);
nand U1255 (N_1255,N_1129,N_1048);
and U1256 (N_1256,N_1086,N_1094);
nor U1257 (N_1257,N_1016,N_1183);
nor U1258 (N_1258,N_1060,N_1021);
nor U1259 (N_1259,N_1033,N_1156);
nor U1260 (N_1260,N_1161,N_1032);
nor U1261 (N_1261,N_1044,N_1052);
nand U1262 (N_1262,N_1070,N_1064);
nor U1263 (N_1263,N_1150,N_1042);
nand U1264 (N_1264,N_1045,N_1114);
nand U1265 (N_1265,N_1023,N_1162);
nand U1266 (N_1266,N_1113,N_1151);
or U1267 (N_1267,N_1119,N_1116);
and U1268 (N_1268,N_1149,N_1127);
nor U1269 (N_1269,N_1051,N_1140);
and U1270 (N_1270,N_1004,N_1017);
nand U1271 (N_1271,N_1077,N_1169);
nor U1272 (N_1272,N_1065,N_1194);
nor U1273 (N_1273,N_1186,N_1006);
nor U1274 (N_1274,N_1160,N_1025);
and U1275 (N_1275,N_1029,N_1100);
nand U1276 (N_1276,N_1131,N_1008);
nor U1277 (N_1277,N_1101,N_1106);
nor U1278 (N_1278,N_1117,N_1121);
or U1279 (N_1279,N_1170,N_1098);
nor U1280 (N_1280,N_1035,N_1199);
nand U1281 (N_1281,N_1148,N_1135);
or U1282 (N_1282,N_1026,N_1163);
nand U1283 (N_1283,N_1118,N_1153);
nor U1284 (N_1284,N_1082,N_1084);
nand U1285 (N_1285,N_1024,N_1081);
and U1286 (N_1286,N_1130,N_1143);
xnor U1287 (N_1287,N_1007,N_1157);
nand U1288 (N_1288,N_1166,N_1142);
nand U1289 (N_1289,N_1085,N_1093);
nor U1290 (N_1290,N_1055,N_1088);
and U1291 (N_1291,N_1043,N_1158);
nand U1292 (N_1292,N_1040,N_1075);
xnor U1293 (N_1293,N_1139,N_1180);
or U1294 (N_1294,N_1097,N_1188);
nor U1295 (N_1295,N_1134,N_1115);
or U1296 (N_1296,N_1072,N_1192);
nand U1297 (N_1297,N_1179,N_1018);
nor U1298 (N_1298,N_1136,N_1047);
nand U1299 (N_1299,N_1078,N_1099);
xnor U1300 (N_1300,N_1173,N_1129);
nor U1301 (N_1301,N_1087,N_1032);
and U1302 (N_1302,N_1140,N_1116);
and U1303 (N_1303,N_1097,N_1098);
nor U1304 (N_1304,N_1142,N_1094);
and U1305 (N_1305,N_1061,N_1141);
and U1306 (N_1306,N_1109,N_1192);
or U1307 (N_1307,N_1152,N_1031);
nand U1308 (N_1308,N_1173,N_1007);
nor U1309 (N_1309,N_1062,N_1155);
nand U1310 (N_1310,N_1090,N_1162);
or U1311 (N_1311,N_1026,N_1131);
nor U1312 (N_1312,N_1020,N_1068);
xnor U1313 (N_1313,N_1018,N_1167);
and U1314 (N_1314,N_1092,N_1013);
nand U1315 (N_1315,N_1050,N_1184);
nor U1316 (N_1316,N_1040,N_1068);
and U1317 (N_1317,N_1124,N_1114);
nor U1318 (N_1318,N_1071,N_1010);
xor U1319 (N_1319,N_1132,N_1115);
nand U1320 (N_1320,N_1060,N_1089);
and U1321 (N_1321,N_1080,N_1105);
or U1322 (N_1322,N_1179,N_1092);
nor U1323 (N_1323,N_1085,N_1024);
or U1324 (N_1324,N_1011,N_1023);
nor U1325 (N_1325,N_1154,N_1046);
and U1326 (N_1326,N_1110,N_1115);
nand U1327 (N_1327,N_1034,N_1013);
or U1328 (N_1328,N_1199,N_1081);
nor U1329 (N_1329,N_1132,N_1060);
nand U1330 (N_1330,N_1087,N_1182);
and U1331 (N_1331,N_1146,N_1070);
nand U1332 (N_1332,N_1141,N_1060);
nor U1333 (N_1333,N_1188,N_1104);
nand U1334 (N_1334,N_1044,N_1004);
or U1335 (N_1335,N_1031,N_1177);
nand U1336 (N_1336,N_1184,N_1016);
nand U1337 (N_1337,N_1101,N_1090);
and U1338 (N_1338,N_1005,N_1171);
and U1339 (N_1339,N_1188,N_1060);
xor U1340 (N_1340,N_1151,N_1170);
nand U1341 (N_1341,N_1194,N_1102);
nor U1342 (N_1342,N_1131,N_1082);
nor U1343 (N_1343,N_1117,N_1049);
nor U1344 (N_1344,N_1018,N_1035);
xor U1345 (N_1345,N_1050,N_1107);
nand U1346 (N_1346,N_1077,N_1123);
xor U1347 (N_1347,N_1005,N_1196);
nand U1348 (N_1348,N_1081,N_1068);
xnor U1349 (N_1349,N_1114,N_1135);
nor U1350 (N_1350,N_1066,N_1166);
nor U1351 (N_1351,N_1076,N_1183);
and U1352 (N_1352,N_1035,N_1195);
nor U1353 (N_1353,N_1134,N_1059);
nor U1354 (N_1354,N_1118,N_1198);
nor U1355 (N_1355,N_1100,N_1102);
or U1356 (N_1356,N_1198,N_1027);
or U1357 (N_1357,N_1194,N_1100);
nand U1358 (N_1358,N_1133,N_1145);
nand U1359 (N_1359,N_1120,N_1144);
or U1360 (N_1360,N_1069,N_1118);
nor U1361 (N_1361,N_1007,N_1080);
and U1362 (N_1362,N_1006,N_1141);
nor U1363 (N_1363,N_1102,N_1045);
nor U1364 (N_1364,N_1061,N_1151);
nor U1365 (N_1365,N_1051,N_1097);
and U1366 (N_1366,N_1136,N_1013);
nor U1367 (N_1367,N_1058,N_1087);
nor U1368 (N_1368,N_1029,N_1189);
nand U1369 (N_1369,N_1038,N_1064);
and U1370 (N_1370,N_1057,N_1099);
nand U1371 (N_1371,N_1140,N_1091);
nor U1372 (N_1372,N_1198,N_1127);
or U1373 (N_1373,N_1163,N_1193);
nand U1374 (N_1374,N_1037,N_1062);
or U1375 (N_1375,N_1079,N_1129);
or U1376 (N_1376,N_1008,N_1139);
or U1377 (N_1377,N_1193,N_1012);
nand U1378 (N_1378,N_1071,N_1084);
or U1379 (N_1379,N_1120,N_1185);
and U1380 (N_1380,N_1102,N_1023);
or U1381 (N_1381,N_1194,N_1075);
xnor U1382 (N_1382,N_1066,N_1177);
nor U1383 (N_1383,N_1154,N_1180);
nand U1384 (N_1384,N_1185,N_1014);
nor U1385 (N_1385,N_1079,N_1049);
nor U1386 (N_1386,N_1112,N_1122);
nor U1387 (N_1387,N_1134,N_1170);
nor U1388 (N_1388,N_1009,N_1061);
or U1389 (N_1389,N_1171,N_1087);
nand U1390 (N_1390,N_1048,N_1198);
or U1391 (N_1391,N_1012,N_1163);
and U1392 (N_1392,N_1180,N_1183);
and U1393 (N_1393,N_1095,N_1161);
or U1394 (N_1394,N_1038,N_1001);
and U1395 (N_1395,N_1094,N_1102);
nor U1396 (N_1396,N_1041,N_1118);
and U1397 (N_1397,N_1111,N_1149);
nand U1398 (N_1398,N_1170,N_1165);
nor U1399 (N_1399,N_1057,N_1159);
nor U1400 (N_1400,N_1298,N_1240);
or U1401 (N_1401,N_1347,N_1387);
nand U1402 (N_1402,N_1304,N_1331);
nand U1403 (N_1403,N_1204,N_1241);
nor U1404 (N_1404,N_1230,N_1397);
xnor U1405 (N_1405,N_1220,N_1324);
and U1406 (N_1406,N_1314,N_1285);
and U1407 (N_1407,N_1355,N_1280);
nor U1408 (N_1408,N_1217,N_1261);
xnor U1409 (N_1409,N_1364,N_1210);
xor U1410 (N_1410,N_1234,N_1268);
or U1411 (N_1411,N_1201,N_1349);
nand U1412 (N_1412,N_1270,N_1265);
nand U1413 (N_1413,N_1371,N_1218);
or U1414 (N_1414,N_1277,N_1273);
or U1415 (N_1415,N_1318,N_1337);
nor U1416 (N_1416,N_1325,N_1363);
nor U1417 (N_1417,N_1336,N_1249);
or U1418 (N_1418,N_1326,N_1316);
xor U1419 (N_1419,N_1388,N_1329);
nor U1420 (N_1420,N_1225,N_1321);
and U1421 (N_1421,N_1332,N_1374);
xor U1422 (N_1422,N_1237,N_1315);
nand U1423 (N_1423,N_1360,N_1323);
or U1424 (N_1424,N_1356,N_1254);
xnor U1425 (N_1425,N_1399,N_1366);
and U1426 (N_1426,N_1297,N_1203);
nor U1427 (N_1427,N_1386,N_1307);
nor U1428 (N_1428,N_1384,N_1269);
or U1429 (N_1429,N_1377,N_1359);
nor U1430 (N_1430,N_1346,N_1290);
nand U1431 (N_1431,N_1227,N_1219);
nor U1432 (N_1432,N_1393,N_1275);
nor U1433 (N_1433,N_1250,N_1317);
nand U1434 (N_1434,N_1340,N_1226);
or U1435 (N_1435,N_1288,N_1330);
and U1436 (N_1436,N_1276,N_1202);
nor U1437 (N_1437,N_1350,N_1221);
or U1438 (N_1438,N_1351,N_1251);
nand U1439 (N_1439,N_1242,N_1303);
or U1440 (N_1440,N_1342,N_1224);
and U1441 (N_1441,N_1287,N_1320);
and U1442 (N_1442,N_1243,N_1211);
nand U1443 (N_1443,N_1259,N_1246);
nand U1444 (N_1444,N_1370,N_1361);
nor U1445 (N_1445,N_1390,N_1222);
or U1446 (N_1446,N_1252,N_1214);
or U1447 (N_1447,N_1372,N_1255);
or U1448 (N_1448,N_1369,N_1313);
nand U1449 (N_1449,N_1274,N_1348);
nand U1450 (N_1450,N_1266,N_1294);
xor U1451 (N_1451,N_1345,N_1367);
nor U1452 (N_1452,N_1306,N_1282);
and U1453 (N_1453,N_1257,N_1385);
and U1454 (N_1454,N_1205,N_1380);
and U1455 (N_1455,N_1295,N_1309);
nor U1456 (N_1456,N_1292,N_1248);
nand U1457 (N_1457,N_1293,N_1357);
xnor U1458 (N_1458,N_1383,N_1311);
or U1459 (N_1459,N_1344,N_1228);
or U1460 (N_1460,N_1352,N_1373);
and U1461 (N_1461,N_1365,N_1362);
nand U1462 (N_1462,N_1278,N_1392);
or U1463 (N_1463,N_1291,N_1232);
or U1464 (N_1464,N_1236,N_1272);
xor U1465 (N_1465,N_1200,N_1206);
or U1466 (N_1466,N_1247,N_1279);
or U1467 (N_1467,N_1319,N_1267);
and U1468 (N_1468,N_1212,N_1245);
and U1469 (N_1469,N_1310,N_1244);
nor U1470 (N_1470,N_1376,N_1375);
nor U1471 (N_1471,N_1300,N_1299);
and U1472 (N_1472,N_1308,N_1289);
or U1473 (N_1473,N_1283,N_1312);
nor U1474 (N_1474,N_1233,N_1368);
or U1475 (N_1475,N_1322,N_1231);
and U1476 (N_1476,N_1216,N_1333);
or U1477 (N_1477,N_1253,N_1263);
or U1478 (N_1478,N_1264,N_1353);
and U1479 (N_1479,N_1229,N_1328);
and U1480 (N_1480,N_1382,N_1339);
xor U1481 (N_1481,N_1398,N_1260);
nor U1482 (N_1482,N_1389,N_1281);
or U1483 (N_1483,N_1378,N_1343);
nand U1484 (N_1484,N_1391,N_1341);
or U1485 (N_1485,N_1256,N_1301);
and U1486 (N_1486,N_1239,N_1335);
and U1487 (N_1487,N_1305,N_1296);
nor U1488 (N_1488,N_1395,N_1215);
and U1489 (N_1489,N_1381,N_1207);
or U1490 (N_1490,N_1327,N_1338);
nor U1491 (N_1491,N_1354,N_1334);
or U1492 (N_1492,N_1379,N_1208);
nand U1493 (N_1493,N_1258,N_1271);
or U1494 (N_1494,N_1358,N_1223);
nor U1495 (N_1495,N_1286,N_1302);
nor U1496 (N_1496,N_1209,N_1396);
nand U1497 (N_1497,N_1238,N_1235);
nor U1498 (N_1498,N_1213,N_1262);
nand U1499 (N_1499,N_1394,N_1284);
and U1500 (N_1500,N_1321,N_1204);
or U1501 (N_1501,N_1346,N_1240);
nor U1502 (N_1502,N_1367,N_1375);
xor U1503 (N_1503,N_1241,N_1211);
or U1504 (N_1504,N_1279,N_1255);
or U1505 (N_1505,N_1305,N_1240);
nand U1506 (N_1506,N_1328,N_1290);
nand U1507 (N_1507,N_1390,N_1393);
nor U1508 (N_1508,N_1378,N_1392);
nand U1509 (N_1509,N_1253,N_1373);
nand U1510 (N_1510,N_1263,N_1372);
nor U1511 (N_1511,N_1243,N_1269);
nor U1512 (N_1512,N_1313,N_1311);
nor U1513 (N_1513,N_1318,N_1210);
nand U1514 (N_1514,N_1322,N_1313);
and U1515 (N_1515,N_1309,N_1211);
and U1516 (N_1516,N_1209,N_1344);
and U1517 (N_1517,N_1246,N_1260);
nor U1518 (N_1518,N_1241,N_1347);
xnor U1519 (N_1519,N_1279,N_1237);
xnor U1520 (N_1520,N_1280,N_1226);
or U1521 (N_1521,N_1331,N_1373);
or U1522 (N_1522,N_1213,N_1256);
or U1523 (N_1523,N_1338,N_1277);
nand U1524 (N_1524,N_1250,N_1238);
xnor U1525 (N_1525,N_1322,N_1230);
nor U1526 (N_1526,N_1326,N_1358);
and U1527 (N_1527,N_1366,N_1214);
nor U1528 (N_1528,N_1293,N_1235);
or U1529 (N_1529,N_1262,N_1390);
and U1530 (N_1530,N_1253,N_1336);
and U1531 (N_1531,N_1217,N_1239);
and U1532 (N_1532,N_1347,N_1255);
and U1533 (N_1533,N_1358,N_1291);
xnor U1534 (N_1534,N_1383,N_1306);
nand U1535 (N_1535,N_1287,N_1200);
nand U1536 (N_1536,N_1305,N_1266);
xnor U1537 (N_1537,N_1260,N_1362);
and U1538 (N_1538,N_1384,N_1297);
nand U1539 (N_1539,N_1233,N_1305);
nor U1540 (N_1540,N_1309,N_1226);
or U1541 (N_1541,N_1313,N_1223);
nor U1542 (N_1542,N_1297,N_1341);
nor U1543 (N_1543,N_1249,N_1268);
or U1544 (N_1544,N_1353,N_1337);
or U1545 (N_1545,N_1353,N_1256);
and U1546 (N_1546,N_1366,N_1280);
nand U1547 (N_1547,N_1299,N_1202);
and U1548 (N_1548,N_1336,N_1246);
nand U1549 (N_1549,N_1237,N_1399);
or U1550 (N_1550,N_1231,N_1276);
nor U1551 (N_1551,N_1207,N_1370);
and U1552 (N_1552,N_1219,N_1204);
or U1553 (N_1553,N_1302,N_1202);
and U1554 (N_1554,N_1280,N_1210);
or U1555 (N_1555,N_1206,N_1354);
or U1556 (N_1556,N_1314,N_1303);
and U1557 (N_1557,N_1238,N_1346);
or U1558 (N_1558,N_1205,N_1338);
xor U1559 (N_1559,N_1303,N_1338);
nand U1560 (N_1560,N_1384,N_1301);
or U1561 (N_1561,N_1379,N_1258);
and U1562 (N_1562,N_1323,N_1394);
nor U1563 (N_1563,N_1280,N_1327);
and U1564 (N_1564,N_1398,N_1297);
or U1565 (N_1565,N_1244,N_1346);
nand U1566 (N_1566,N_1292,N_1202);
nor U1567 (N_1567,N_1287,N_1353);
xor U1568 (N_1568,N_1265,N_1298);
and U1569 (N_1569,N_1203,N_1273);
nand U1570 (N_1570,N_1206,N_1336);
or U1571 (N_1571,N_1359,N_1293);
or U1572 (N_1572,N_1229,N_1252);
or U1573 (N_1573,N_1265,N_1338);
or U1574 (N_1574,N_1365,N_1374);
xor U1575 (N_1575,N_1306,N_1253);
nor U1576 (N_1576,N_1384,N_1244);
nand U1577 (N_1577,N_1207,N_1296);
nand U1578 (N_1578,N_1379,N_1364);
nor U1579 (N_1579,N_1285,N_1356);
xnor U1580 (N_1580,N_1288,N_1296);
nand U1581 (N_1581,N_1375,N_1214);
nor U1582 (N_1582,N_1256,N_1304);
or U1583 (N_1583,N_1372,N_1390);
or U1584 (N_1584,N_1332,N_1209);
nor U1585 (N_1585,N_1308,N_1287);
and U1586 (N_1586,N_1216,N_1231);
nand U1587 (N_1587,N_1210,N_1279);
and U1588 (N_1588,N_1263,N_1377);
and U1589 (N_1589,N_1394,N_1270);
and U1590 (N_1590,N_1257,N_1301);
nor U1591 (N_1591,N_1310,N_1235);
and U1592 (N_1592,N_1284,N_1297);
nand U1593 (N_1593,N_1367,N_1213);
nor U1594 (N_1594,N_1357,N_1226);
or U1595 (N_1595,N_1264,N_1315);
or U1596 (N_1596,N_1235,N_1330);
or U1597 (N_1597,N_1387,N_1336);
xnor U1598 (N_1598,N_1348,N_1384);
xnor U1599 (N_1599,N_1337,N_1320);
or U1600 (N_1600,N_1442,N_1528);
nand U1601 (N_1601,N_1446,N_1540);
nor U1602 (N_1602,N_1570,N_1407);
or U1603 (N_1603,N_1565,N_1481);
or U1604 (N_1604,N_1408,N_1454);
or U1605 (N_1605,N_1559,N_1549);
xnor U1606 (N_1606,N_1494,N_1420);
and U1607 (N_1607,N_1558,N_1554);
nor U1608 (N_1608,N_1564,N_1429);
or U1609 (N_1609,N_1529,N_1468);
nor U1610 (N_1610,N_1597,N_1553);
or U1611 (N_1611,N_1480,N_1531);
or U1612 (N_1612,N_1461,N_1426);
or U1613 (N_1613,N_1589,N_1542);
nor U1614 (N_1614,N_1574,N_1452);
and U1615 (N_1615,N_1576,N_1438);
nand U1616 (N_1616,N_1493,N_1458);
nor U1617 (N_1617,N_1561,N_1424);
xnor U1618 (N_1618,N_1526,N_1457);
and U1619 (N_1619,N_1590,N_1437);
or U1620 (N_1620,N_1509,N_1534);
xor U1621 (N_1621,N_1573,N_1506);
or U1622 (N_1622,N_1598,N_1449);
and U1623 (N_1623,N_1502,N_1412);
nand U1624 (N_1624,N_1472,N_1413);
or U1625 (N_1625,N_1478,N_1594);
and U1626 (N_1626,N_1585,N_1591);
xor U1627 (N_1627,N_1462,N_1518);
and U1628 (N_1628,N_1414,N_1434);
and U1629 (N_1629,N_1514,N_1586);
or U1630 (N_1630,N_1541,N_1450);
nor U1631 (N_1631,N_1588,N_1537);
and U1632 (N_1632,N_1491,N_1427);
nand U1633 (N_1633,N_1431,N_1535);
nand U1634 (N_1634,N_1495,N_1521);
xor U1635 (N_1635,N_1552,N_1415);
or U1636 (N_1636,N_1425,N_1584);
xor U1637 (N_1637,N_1508,N_1497);
nand U1638 (N_1638,N_1583,N_1499);
or U1639 (N_1639,N_1572,N_1401);
and U1640 (N_1640,N_1448,N_1405);
and U1641 (N_1641,N_1593,N_1473);
and U1642 (N_1642,N_1443,N_1505);
nand U1643 (N_1643,N_1512,N_1406);
or U1644 (N_1644,N_1595,N_1547);
nand U1645 (N_1645,N_1435,N_1440);
or U1646 (N_1646,N_1581,N_1538);
nand U1647 (N_1647,N_1482,N_1483);
nand U1648 (N_1648,N_1592,N_1563);
and U1649 (N_1649,N_1492,N_1411);
and U1650 (N_1650,N_1578,N_1471);
and U1651 (N_1651,N_1469,N_1404);
nand U1652 (N_1652,N_1527,N_1470);
xor U1653 (N_1653,N_1479,N_1490);
nand U1654 (N_1654,N_1410,N_1451);
or U1655 (N_1655,N_1510,N_1544);
and U1656 (N_1656,N_1568,N_1545);
nand U1657 (N_1657,N_1477,N_1419);
or U1658 (N_1658,N_1486,N_1459);
or U1659 (N_1659,N_1460,N_1519);
nor U1660 (N_1660,N_1539,N_1569);
or U1661 (N_1661,N_1496,N_1432);
nand U1662 (N_1662,N_1464,N_1465);
nand U1663 (N_1663,N_1575,N_1504);
nand U1664 (N_1664,N_1430,N_1560);
xor U1665 (N_1665,N_1417,N_1511);
and U1666 (N_1666,N_1467,N_1548);
nand U1667 (N_1667,N_1421,N_1463);
nand U1668 (N_1668,N_1507,N_1520);
and U1669 (N_1669,N_1557,N_1475);
xor U1670 (N_1670,N_1532,N_1485);
nor U1671 (N_1671,N_1501,N_1579);
nor U1672 (N_1672,N_1466,N_1523);
or U1673 (N_1673,N_1571,N_1441);
nor U1674 (N_1674,N_1567,N_1456);
nand U1675 (N_1675,N_1444,N_1543);
or U1676 (N_1676,N_1403,N_1416);
nand U1677 (N_1677,N_1418,N_1476);
nor U1678 (N_1678,N_1533,N_1522);
or U1679 (N_1679,N_1488,N_1422);
nand U1680 (N_1680,N_1484,N_1577);
or U1681 (N_1681,N_1498,N_1587);
or U1682 (N_1682,N_1582,N_1409);
and U1683 (N_1683,N_1524,N_1445);
nand U1684 (N_1684,N_1487,N_1546);
xnor U1685 (N_1685,N_1423,N_1516);
nor U1686 (N_1686,N_1580,N_1513);
xnor U1687 (N_1687,N_1555,N_1474);
or U1688 (N_1688,N_1556,N_1436);
and U1689 (N_1689,N_1562,N_1433);
and U1690 (N_1690,N_1515,N_1530);
and U1691 (N_1691,N_1517,N_1551);
nor U1692 (N_1692,N_1525,N_1455);
or U1693 (N_1693,N_1400,N_1566);
nor U1694 (N_1694,N_1599,N_1402);
and U1695 (N_1695,N_1503,N_1596);
or U1696 (N_1696,N_1428,N_1550);
and U1697 (N_1697,N_1536,N_1489);
or U1698 (N_1698,N_1500,N_1453);
and U1699 (N_1699,N_1439,N_1447);
nand U1700 (N_1700,N_1581,N_1499);
xnor U1701 (N_1701,N_1460,N_1407);
nand U1702 (N_1702,N_1419,N_1406);
nor U1703 (N_1703,N_1480,N_1426);
and U1704 (N_1704,N_1517,N_1448);
nand U1705 (N_1705,N_1430,N_1574);
or U1706 (N_1706,N_1552,N_1479);
or U1707 (N_1707,N_1490,N_1598);
and U1708 (N_1708,N_1437,N_1430);
nand U1709 (N_1709,N_1475,N_1593);
xnor U1710 (N_1710,N_1429,N_1481);
or U1711 (N_1711,N_1504,N_1514);
nand U1712 (N_1712,N_1581,N_1528);
nand U1713 (N_1713,N_1467,N_1471);
nor U1714 (N_1714,N_1457,N_1432);
nor U1715 (N_1715,N_1431,N_1509);
nor U1716 (N_1716,N_1456,N_1430);
nor U1717 (N_1717,N_1599,N_1534);
nor U1718 (N_1718,N_1476,N_1451);
nor U1719 (N_1719,N_1422,N_1499);
or U1720 (N_1720,N_1581,N_1483);
nand U1721 (N_1721,N_1578,N_1543);
or U1722 (N_1722,N_1536,N_1445);
nand U1723 (N_1723,N_1462,N_1526);
nor U1724 (N_1724,N_1544,N_1520);
or U1725 (N_1725,N_1421,N_1437);
or U1726 (N_1726,N_1527,N_1440);
or U1727 (N_1727,N_1510,N_1415);
nand U1728 (N_1728,N_1573,N_1498);
nand U1729 (N_1729,N_1487,N_1490);
or U1730 (N_1730,N_1534,N_1585);
or U1731 (N_1731,N_1541,N_1592);
nor U1732 (N_1732,N_1413,N_1555);
or U1733 (N_1733,N_1467,N_1402);
or U1734 (N_1734,N_1531,N_1458);
or U1735 (N_1735,N_1490,N_1426);
and U1736 (N_1736,N_1409,N_1463);
and U1737 (N_1737,N_1530,N_1597);
nor U1738 (N_1738,N_1575,N_1553);
or U1739 (N_1739,N_1479,N_1540);
xor U1740 (N_1740,N_1593,N_1585);
and U1741 (N_1741,N_1488,N_1524);
or U1742 (N_1742,N_1427,N_1415);
nor U1743 (N_1743,N_1550,N_1574);
nor U1744 (N_1744,N_1442,N_1418);
and U1745 (N_1745,N_1494,N_1584);
nand U1746 (N_1746,N_1500,N_1586);
and U1747 (N_1747,N_1425,N_1501);
nand U1748 (N_1748,N_1572,N_1443);
xnor U1749 (N_1749,N_1486,N_1472);
or U1750 (N_1750,N_1494,N_1467);
or U1751 (N_1751,N_1546,N_1460);
and U1752 (N_1752,N_1472,N_1499);
or U1753 (N_1753,N_1524,N_1429);
nand U1754 (N_1754,N_1476,N_1581);
nand U1755 (N_1755,N_1511,N_1556);
and U1756 (N_1756,N_1461,N_1514);
nand U1757 (N_1757,N_1432,N_1430);
nand U1758 (N_1758,N_1511,N_1586);
nand U1759 (N_1759,N_1494,N_1526);
nand U1760 (N_1760,N_1421,N_1570);
and U1761 (N_1761,N_1584,N_1464);
or U1762 (N_1762,N_1533,N_1515);
or U1763 (N_1763,N_1539,N_1401);
nand U1764 (N_1764,N_1589,N_1552);
and U1765 (N_1765,N_1419,N_1411);
nand U1766 (N_1766,N_1438,N_1461);
and U1767 (N_1767,N_1582,N_1482);
nand U1768 (N_1768,N_1519,N_1562);
nand U1769 (N_1769,N_1599,N_1564);
nor U1770 (N_1770,N_1453,N_1519);
or U1771 (N_1771,N_1578,N_1505);
xor U1772 (N_1772,N_1425,N_1401);
nand U1773 (N_1773,N_1560,N_1484);
or U1774 (N_1774,N_1507,N_1451);
nand U1775 (N_1775,N_1574,N_1478);
nor U1776 (N_1776,N_1596,N_1545);
and U1777 (N_1777,N_1483,N_1553);
and U1778 (N_1778,N_1524,N_1559);
and U1779 (N_1779,N_1509,N_1498);
and U1780 (N_1780,N_1418,N_1444);
nor U1781 (N_1781,N_1465,N_1510);
or U1782 (N_1782,N_1462,N_1474);
or U1783 (N_1783,N_1441,N_1445);
and U1784 (N_1784,N_1569,N_1451);
nand U1785 (N_1785,N_1591,N_1521);
nor U1786 (N_1786,N_1580,N_1421);
or U1787 (N_1787,N_1418,N_1420);
xor U1788 (N_1788,N_1511,N_1433);
or U1789 (N_1789,N_1431,N_1434);
and U1790 (N_1790,N_1409,N_1543);
or U1791 (N_1791,N_1545,N_1479);
nor U1792 (N_1792,N_1559,N_1487);
xnor U1793 (N_1793,N_1495,N_1488);
and U1794 (N_1794,N_1522,N_1596);
nor U1795 (N_1795,N_1432,N_1531);
nand U1796 (N_1796,N_1569,N_1595);
and U1797 (N_1797,N_1522,N_1473);
nor U1798 (N_1798,N_1510,N_1424);
nor U1799 (N_1799,N_1515,N_1467);
or U1800 (N_1800,N_1613,N_1674);
xnor U1801 (N_1801,N_1668,N_1781);
nor U1802 (N_1802,N_1785,N_1793);
xor U1803 (N_1803,N_1787,N_1690);
nand U1804 (N_1804,N_1630,N_1693);
and U1805 (N_1805,N_1737,N_1609);
or U1806 (N_1806,N_1754,N_1721);
nand U1807 (N_1807,N_1736,N_1774);
or U1808 (N_1808,N_1727,N_1604);
nand U1809 (N_1809,N_1689,N_1636);
nor U1810 (N_1810,N_1672,N_1718);
nand U1811 (N_1811,N_1653,N_1716);
nor U1812 (N_1812,N_1799,N_1738);
nand U1813 (N_1813,N_1629,N_1616);
nand U1814 (N_1814,N_1768,N_1703);
nand U1815 (N_1815,N_1683,N_1763);
or U1816 (N_1816,N_1654,N_1700);
and U1817 (N_1817,N_1766,N_1610);
nor U1818 (N_1818,N_1606,N_1709);
nor U1819 (N_1819,N_1678,N_1641);
and U1820 (N_1820,N_1662,N_1644);
nand U1821 (N_1821,N_1776,N_1755);
and U1822 (N_1822,N_1618,N_1634);
nand U1823 (N_1823,N_1740,N_1627);
xnor U1824 (N_1824,N_1734,N_1640);
nand U1825 (N_1825,N_1702,N_1728);
or U1826 (N_1826,N_1749,N_1650);
nor U1827 (N_1827,N_1626,N_1792);
or U1828 (N_1828,N_1643,N_1769);
xnor U1829 (N_1829,N_1696,N_1675);
nor U1830 (N_1830,N_1655,N_1707);
and U1831 (N_1831,N_1656,N_1743);
nand U1832 (N_1832,N_1713,N_1708);
nor U1833 (N_1833,N_1680,N_1796);
nand U1834 (N_1834,N_1615,N_1651);
nand U1835 (N_1835,N_1665,N_1756);
nor U1836 (N_1836,N_1660,N_1622);
or U1837 (N_1837,N_1642,N_1633);
and U1838 (N_1838,N_1730,N_1788);
nand U1839 (N_1839,N_1773,N_1646);
nor U1840 (N_1840,N_1666,N_1649);
or U1841 (N_1841,N_1695,N_1625);
and U1842 (N_1842,N_1676,N_1742);
nor U1843 (N_1843,N_1767,N_1659);
or U1844 (N_1844,N_1741,N_1778);
nor U1845 (N_1845,N_1647,N_1797);
nor U1846 (N_1846,N_1612,N_1733);
nand U1847 (N_1847,N_1684,N_1670);
and U1848 (N_1848,N_1677,N_1779);
and U1849 (N_1849,N_1710,N_1632);
nor U1850 (N_1850,N_1603,N_1783);
nor U1851 (N_1851,N_1614,N_1764);
xnor U1852 (N_1852,N_1600,N_1744);
nand U1853 (N_1853,N_1705,N_1795);
nor U1854 (N_1854,N_1681,N_1729);
xnor U1855 (N_1855,N_1723,N_1687);
nor U1856 (N_1856,N_1704,N_1762);
and U1857 (N_1857,N_1637,N_1699);
xor U1858 (N_1858,N_1631,N_1664);
nor U1859 (N_1859,N_1679,N_1752);
or U1860 (N_1860,N_1661,N_1657);
nor U1861 (N_1861,N_1667,N_1697);
nand U1862 (N_1862,N_1724,N_1748);
or U1863 (N_1863,N_1652,N_1602);
nor U1864 (N_1864,N_1790,N_1624);
or U1865 (N_1865,N_1735,N_1691);
nand U1866 (N_1866,N_1692,N_1669);
nand U1867 (N_1867,N_1771,N_1739);
and U1868 (N_1868,N_1760,N_1725);
or U1869 (N_1869,N_1747,N_1775);
nand U1870 (N_1870,N_1685,N_1786);
or U1871 (N_1871,N_1611,N_1663);
and U1872 (N_1872,N_1758,N_1673);
nand U1873 (N_1873,N_1745,N_1686);
nor U1874 (N_1874,N_1761,N_1617);
nand U1875 (N_1875,N_1794,N_1706);
or U1876 (N_1876,N_1726,N_1719);
and U1877 (N_1877,N_1619,N_1635);
or U1878 (N_1878,N_1682,N_1621);
or U1879 (N_1879,N_1698,N_1711);
and U1880 (N_1880,N_1605,N_1623);
nor U1881 (N_1881,N_1648,N_1607);
and U1882 (N_1882,N_1798,N_1746);
or U1883 (N_1883,N_1732,N_1780);
and U1884 (N_1884,N_1791,N_1782);
nand U1885 (N_1885,N_1701,N_1720);
or U1886 (N_1886,N_1765,N_1608);
nand U1887 (N_1887,N_1638,N_1639);
nor U1888 (N_1888,N_1717,N_1784);
nand U1889 (N_1889,N_1601,N_1671);
nand U1890 (N_1890,N_1751,N_1759);
nor U1891 (N_1891,N_1753,N_1620);
nand U1892 (N_1892,N_1722,N_1770);
nand U1893 (N_1893,N_1777,N_1757);
or U1894 (N_1894,N_1694,N_1789);
nor U1895 (N_1895,N_1715,N_1712);
nand U1896 (N_1896,N_1688,N_1750);
nor U1897 (N_1897,N_1658,N_1628);
and U1898 (N_1898,N_1731,N_1714);
nor U1899 (N_1899,N_1772,N_1645);
nor U1900 (N_1900,N_1798,N_1689);
and U1901 (N_1901,N_1745,N_1758);
nor U1902 (N_1902,N_1641,N_1766);
or U1903 (N_1903,N_1776,N_1719);
nand U1904 (N_1904,N_1701,N_1656);
nand U1905 (N_1905,N_1787,N_1731);
and U1906 (N_1906,N_1761,N_1676);
or U1907 (N_1907,N_1792,N_1775);
nor U1908 (N_1908,N_1725,N_1707);
nand U1909 (N_1909,N_1725,N_1675);
and U1910 (N_1910,N_1725,N_1674);
nor U1911 (N_1911,N_1768,N_1728);
or U1912 (N_1912,N_1737,N_1658);
nand U1913 (N_1913,N_1744,N_1645);
nand U1914 (N_1914,N_1756,N_1771);
or U1915 (N_1915,N_1778,N_1723);
xnor U1916 (N_1916,N_1648,N_1612);
and U1917 (N_1917,N_1677,N_1697);
nor U1918 (N_1918,N_1764,N_1676);
nor U1919 (N_1919,N_1645,N_1657);
and U1920 (N_1920,N_1740,N_1643);
nor U1921 (N_1921,N_1748,N_1763);
nor U1922 (N_1922,N_1645,N_1781);
and U1923 (N_1923,N_1661,N_1732);
xnor U1924 (N_1924,N_1775,N_1613);
nor U1925 (N_1925,N_1604,N_1749);
nand U1926 (N_1926,N_1782,N_1609);
nand U1927 (N_1927,N_1776,N_1749);
or U1928 (N_1928,N_1690,N_1678);
nand U1929 (N_1929,N_1699,N_1673);
nor U1930 (N_1930,N_1718,N_1603);
xnor U1931 (N_1931,N_1661,N_1737);
xnor U1932 (N_1932,N_1753,N_1778);
or U1933 (N_1933,N_1773,N_1672);
or U1934 (N_1934,N_1750,N_1621);
nand U1935 (N_1935,N_1791,N_1799);
nand U1936 (N_1936,N_1608,N_1700);
and U1937 (N_1937,N_1601,N_1611);
and U1938 (N_1938,N_1602,N_1778);
xnor U1939 (N_1939,N_1649,N_1799);
and U1940 (N_1940,N_1711,N_1655);
and U1941 (N_1941,N_1761,N_1759);
or U1942 (N_1942,N_1712,N_1754);
nor U1943 (N_1943,N_1797,N_1630);
or U1944 (N_1944,N_1788,N_1689);
nor U1945 (N_1945,N_1711,N_1762);
or U1946 (N_1946,N_1793,N_1763);
or U1947 (N_1947,N_1637,N_1754);
or U1948 (N_1948,N_1774,N_1799);
or U1949 (N_1949,N_1642,N_1771);
and U1950 (N_1950,N_1722,N_1777);
nand U1951 (N_1951,N_1614,N_1787);
nand U1952 (N_1952,N_1742,N_1688);
nor U1953 (N_1953,N_1613,N_1760);
or U1954 (N_1954,N_1617,N_1723);
nand U1955 (N_1955,N_1753,N_1610);
or U1956 (N_1956,N_1690,N_1795);
nor U1957 (N_1957,N_1752,N_1629);
nand U1958 (N_1958,N_1669,N_1712);
nor U1959 (N_1959,N_1635,N_1756);
nand U1960 (N_1960,N_1746,N_1692);
or U1961 (N_1961,N_1731,N_1726);
nor U1962 (N_1962,N_1664,N_1702);
xor U1963 (N_1963,N_1635,N_1794);
xnor U1964 (N_1964,N_1710,N_1774);
nor U1965 (N_1965,N_1705,N_1799);
nand U1966 (N_1966,N_1613,N_1732);
or U1967 (N_1967,N_1612,N_1730);
nand U1968 (N_1968,N_1670,N_1662);
nor U1969 (N_1969,N_1682,N_1679);
and U1970 (N_1970,N_1773,N_1799);
nand U1971 (N_1971,N_1697,N_1639);
or U1972 (N_1972,N_1643,N_1602);
nand U1973 (N_1973,N_1643,N_1618);
nand U1974 (N_1974,N_1693,N_1796);
nor U1975 (N_1975,N_1778,N_1639);
nand U1976 (N_1976,N_1779,N_1634);
or U1977 (N_1977,N_1663,N_1711);
nor U1978 (N_1978,N_1750,N_1747);
nor U1979 (N_1979,N_1692,N_1727);
and U1980 (N_1980,N_1653,N_1605);
nor U1981 (N_1981,N_1601,N_1630);
nor U1982 (N_1982,N_1672,N_1723);
or U1983 (N_1983,N_1671,N_1789);
nor U1984 (N_1984,N_1774,N_1661);
and U1985 (N_1985,N_1679,N_1795);
xnor U1986 (N_1986,N_1708,N_1636);
or U1987 (N_1987,N_1711,N_1616);
nor U1988 (N_1988,N_1736,N_1706);
or U1989 (N_1989,N_1626,N_1775);
nor U1990 (N_1990,N_1761,N_1743);
or U1991 (N_1991,N_1778,N_1640);
nor U1992 (N_1992,N_1629,N_1786);
or U1993 (N_1993,N_1628,N_1692);
and U1994 (N_1994,N_1628,N_1639);
nor U1995 (N_1995,N_1616,N_1706);
xor U1996 (N_1996,N_1626,N_1763);
nand U1997 (N_1997,N_1713,N_1717);
nand U1998 (N_1998,N_1645,N_1743);
nor U1999 (N_1999,N_1626,N_1692);
or U2000 (N_2000,N_1804,N_1928);
and U2001 (N_2001,N_1840,N_1942);
xnor U2002 (N_2002,N_1838,N_1939);
nand U2003 (N_2003,N_1819,N_1839);
nor U2004 (N_2004,N_1952,N_1963);
or U2005 (N_2005,N_1943,N_1922);
nor U2006 (N_2006,N_1881,N_1988);
nand U2007 (N_2007,N_1816,N_1806);
and U2008 (N_2008,N_1990,N_1809);
and U2009 (N_2009,N_1894,N_1948);
nand U2010 (N_2010,N_1845,N_1973);
nor U2011 (N_2011,N_1811,N_1980);
or U2012 (N_2012,N_1998,N_1935);
nor U2013 (N_2013,N_1971,N_1882);
xnor U2014 (N_2014,N_1969,N_1855);
nor U2015 (N_2015,N_1803,N_1957);
or U2016 (N_2016,N_1900,N_1904);
nor U2017 (N_2017,N_1932,N_1965);
and U2018 (N_2018,N_1938,N_1807);
or U2019 (N_2019,N_1829,N_1832);
nand U2020 (N_2020,N_1892,N_1985);
and U2021 (N_2021,N_1946,N_1879);
nand U2022 (N_2022,N_1940,N_1986);
nor U2023 (N_2023,N_1826,N_1905);
nand U2024 (N_2024,N_1856,N_1878);
nand U2025 (N_2025,N_1994,N_1987);
nand U2026 (N_2026,N_1857,N_1925);
or U2027 (N_2027,N_1954,N_1966);
or U2028 (N_2028,N_1995,N_1849);
nor U2029 (N_2029,N_1893,N_1828);
nor U2030 (N_2030,N_1981,N_1859);
and U2031 (N_2031,N_1852,N_1921);
or U2032 (N_2032,N_1910,N_1919);
nor U2033 (N_2033,N_1815,N_1929);
or U2034 (N_2034,N_1842,N_1869);
nand U2035 (N_2035,N_1927,N_1906);
or U2036 (N_2036,N_1983,N_1858);
and U2037 (N_2037,N_1895,N_1959);
xor U2038 (N_2038,N_1915,N_1992);
nand U2039 (N_2039,N_1936,N_1918);
nand U2040 (N_2040,N_1873,N_1887);
nand U2041 (N_2041,N_1916,N_1847);
xnor U2042 (N_2042,N_1872,N_1917);
and U2043 (N_2043,N_1949,N_1844);
and U2044 (N_2044,N_1982,N_1977);
xnor U2045 (N_2045,N_1800,N_1837);
nor U2046 (N_2046,N_1962,N_1914);
nand U2047 (N_2047,N_1861,N_1880);
nor U2048 (N_2048,N_1967,N_1899);
and U2049 (N_2049,N_1996,N_1960);
and U2050 (N_2050,N_1820,N_1841);
nand U2051 (N_2051,N_1964,N_1883);
nand U2052 (N_2052,N_1898,N_1801);
or U2053 (N_2053,N_1947,N_1968);
nor U2054 (N_2054,N_1908,N_1870);
nor U2055 (N_2055,N_1950,N_1926);
nand U2056 (N_2056,N_1862,N_1901);
nor U2057 (N_2057,N_1941,N_1810);
nor U2058 (N_2058,N_1955,N_1933);
or U2059 (N_2059,N_1907,N_1909);
nor U2060 (N_2060,N_1843,N_1913);
or U2061 (N_2061,N_1814,N_1891);
and U2062 (N_2062,N_1813,N_1817);
and U2063 (N_2063,N_1802,N_1824);
nand U2064 (N_2064,N_1953,N_1831);
nand U2065 (N_2065,N_1945,N_1818);
nand U2066 (N_2066,N_1911,N_1846);
nor U2067 (N_2067,N_1999,N_1984);
or U2068 (N_2068,N_1833,N_1970);
and U2069 (N_2069,N_1874,N_1863);
nand U2070 (N_2070,N_1835,N_1836);
nand U2071 (N_2071,N_1884,N_1822);
nand U2072 (N_2072,N_1951,N_1961);
xor U2073 (N_2073,N_1993,N_1876);
nand U2074 (N_2074,N_1864,N_1854);
and U2075 (N_2075,N_1867,N_1871);
nand U2076 (N_2076,N_1972,N_1897);
nand U2077 (N_2077,N_1865,N_1903);
nand U2078 (N_2078,N_1923,N_1830);
and U2079 (N_2079,N_1868,N_1937);
nor U2080 (N_2080,N_1991,N_1956);
or U2081 (N_2081,N_1931,N_1885);
nor U2082 (N_2082,N_1934,N_1975);
or U2083 (N_2083,N_1989,N_1805);
or U2084 (N_2084,N_1848,N_1888);
xnor U2085 (N_2085,N_1944,N_1808);
nand U2086 (N_2086,N_1912,N_1958);
or U2087 (N_2087,N_1834,N_1896);
nand U2088 (N_2088,N_1851,N_1825);
and U2089 (N_2089,N_1853,N_1877);
nand U2090 (N_2090,N_1974,N_1827);
nand U2091 (N_2091,N_1889,N_1866);
nor U2092 (N_2092,N_1924,N_1976);
xor U2093 (N_2093,N_1821,N_1860);
and U2094 (N_2094,N_1997,N_1902);
or U2095 (N_2095,N_1979,N_1823);
nor U2096 (N_2096,N_1875,N_1812);
nand U2097 (N_2097,N_1978,N_1886);
nand U2098 (N_2098,N_1850,N_1890);
and U2099 (N_2099,N_1920,N_1930);
and U2100 (N_2100,N_1887,N_1968);
and U2101 (N_2101,N_1978,N_1866);
and U2102 (N_2102,N_1997,N_1932);
nand U2103 (N_2103,N_1920,N_1852);
nand U2104 (N_2104,N_1868,N_1958);
nand U2105 (N_2105,N_1851,N_1803);
nor U2106 (N_2106,N_1937,N_1999);
nor U2107 (N_2107,N_1867,N_1800);
xnor U2108 (N_2108,N_1993,N_1875);
nand U2109 (N_2109,N_1898,N_1895);
or U2110 (N_2110,N_1934,N_1846);
xor U2111 (N_2111,N_1871,N_1845);
xnor U2112 (N_2112,N_1919,N_1978);
nor U2113 (N_2113,N_1813,N_1844);
xor U2114 (N_2114,N_1921,N_1802);
or U2115 (N_2115,N_1997,N_1829);
or U2116 (N_2116,N_1830,N_1936);
nor U2117 (N_2117,N_1805,N_1863);
or U2118 (N_2118,N_1905,N_1881);
and U2119 (N_2119,N_1999,N_1818);
nor U2120 (N_2120,N_1801,N_1973);
or U2121 (N_2121,N_1803,N_1911);
nand U2122 (N_2122,N_1983,N_1993);
nor U2123 (N_2123,N_1926,N_1850);
nor U2124 (N_2124,N_1925,N_1881);
nand U2125 (N_2125,N_1817,N_1960);
nor U2126 (N_2126,N_1853,N_1865);
or U2127 (N_2127,N_1823,N_1939);
or U2128 (N_2128,N_1996,N_1836);
or U2129 (N_2129,N_1905,N_1886);
nor U2130 (N_2130,N_1936,N_1887);
and U2131 (N_2131,N_1821,N_1980);
xnor U2132 (N_2132,N_1864,N_1808);
nand U2133 (N_2133,N_1988,N_1933);
nor U2134 (N_2134,N_1916,N_1929);
and U2135 (N_2135,N_1922,N_1859);
or U2136 (N_2136,N_1996,N_1949);
nor U2137 (N_2137,N_1884,N_1908);
or U2138 (N_2138,N_1843,N_1901);
nor U2139 (N_2139,N_1849,N_1954);
nor U2140 (N_2140,N_1886,N_1872);
or U2141 (N_2141,N_1934,N_1812);
or U2142 (N_2142,N_1840,N_1919);
or U2143 (N_2143,N_1925,N_1895);
or U2144 (N_2144,N_1818,N_1956);
nand U2145 (N_2145,N_1875,N_1963);
nand U2146 (N_2146,N_1840,N_1899);
xor U2147 (N_2147,N_1824,N_1929);
and U2148 (N_2148,N_1913,N_1851);
xor U2149 (N_2149,N_1974,N_1885);
nor U2150 (N_2150,N_1949,N_1824);
nor U2151 (N_2151,N_1846,N_1848);
nor U2152 (N_2152,N_1896,N_1994);
or U2153 (N_2153,N_1888,N_1892);
or U2154 (N_2154,N_1877,N_1869);
or U2155 (N_2155,N_1837,N_1931);
xnor U2156 (N_2156,N_1869,N_1856);
nor U2157 (N_2157,N_1811,N_1865);
nand U2158 (N_2158,N_1863,N_1991);
nand U2159 (N_2159,N_1946,N_1905);
nor U2160 (N_2160,N_1816,N_1861);
nand U2161 (N_2161,N_1981,N_1810);
nand U2162 (N_2162,N_1942,N_1949);
nand U2163 (N_2163,N_1878,N_1875);
xnor U2164 (N_2164,N_1951,N_1924);
xnor U2165 (N_2165,N_1971,N_1995);
xnor U2166 (N_2166,N_1955,N_1987);
and U2167 (N_2167,N_1931,N_1825);
xor U2168 (N_2168,N_1960,N_1944);
and U2169 (N_2169,N_1876,N_1944);
and U2170 (N_2170,N_1805,N_1972);
or U2171 (N_2171,N_1988,N_1866);
xnor U2172 (N_2172,N_1922,N_1949);
nand U2173 (N_2173,N_1846,N_1905);
nor U2174 (N_2174,N_1902,N_1839);
nand U2175 (N_2175,N_1890,N_1927);
or U2176 (N_2176,N_1904,N_1912);
xor U2177 (N_2177,N_1882,N_1983);
or U2178 (N_2178,N_1868,N_1953);
nor U2179 (N_2179,N_1941,N_1931);
nand U2180 (N_2180,N_1838,N_1972);
nand U2181 (N_2181,N_1876,N_1866);
and U2182 (N_2182,N_1800,N_1999);
nand U2183 (N_2183,N_1979,N_1988);
and U2184 (N_2184,N_1929,N_1921);
nor U2185 (N_2185,N_1955,N_1910);
nand U2186 (N_2186,N_1836,N_1872);
nor U2187 (N_2187,N_1965,N_1913);
and U2188 (N_2188,N_1848,N_1883);
nand U2189 (N_2189,N_1926,N_1979);
xnor U2190 (N_2190,N_1860,N_1953);
nand U2191 (N_2191,N_1949,N_1966);
nand U2192 (N_2192,N_1812,N_1894);
nand U2193 (N_2193,N_1890,N_1834);
nor U2194 (N_2194,N_1939,N_1891);
or U2195 (N_2195,N_1987,N_1932);
nor U2196 (N_2196,N_1814,N_1972);
nand U2197 (N_2197,N_1828,N_1844);
or U2198 (N_2198,N_1924,N_1878);
or U2199 (N_2199,N_1825,N_1913);
or U2200 (N_2200,N_2176,N_2112);
nand U2201 (N_2201,N_2125,N_2047);
and U2202 (N_2202,N_2175,N_2122);
and U2203 (N_2203,N_2075,N_2121);
nand U2204 (N_2204,N_2188,N_2131);
and U2205 (N_2205,N_2101,N_2104);
xnor U2206 (N_2206,N_2107,N_2115);
or U2207 (N_2207,N_2026,N_2105);
nor U2208 (N_2208,N_2155,N_2190);
nor U2209 (N_2209,N_2072,N_2185);
and U2210 (N_2210,N_2103,N_2142);
xor U2211 (N_2211,N_2157,N_2180);
nor U2212 (N_2212,N_2051,N_2018);
nand U2213 (N_2213,N_2120,N_2119);
or U2214 (N_2214,N_2021,N_2029);
nor U2215 (N_2215,N_2027,N_2169);
nor U2216 (N_2216,N_2153,N_2147);
nand U2217 (N_2217,N_2002,N_2050);
and U2218 (N_2218,N_2012,N_2111);
nor U2219 (N_2219,N_2179,N_2038);
or U2220 (N_2220,N_2136,N_2117);
or U2221 (N_2221,N_2192,N_2042);
xnor U2222 (N_2222,N_2066,N_2100);
or U2223 (N_2223,N_2146,N_2049);
or U2224 (N_2224,N_2053,N_2081);
nand U2225 (N_2225,N_2006,N_2085);
nor U2226 (N_2226,N_2106,N_2032);
or U2227 (N_2227,N_2011,N_2184);
nand U2228 (N_2228,N_2123,N_2141);
or U2229 (N_2229,N_2045,N_2148);
nor U2230 (N_2230,N_2178,N_2160);
nor U2231 (N_2231,N_2158,N_2073);
nand U2232 (N_2232,N_2191,N_2154);
and U2233 (N_2233,N_2069,N_2070);
xnor U2234 (N_2234,N_2062,N_2128);
nand U2235 (N_2235,N_2095,N_2030);
and U2236 (N_2236,N_2114,N_2198);
nor U2237 (N_2237,N_2004,N_2118);
and U2238 (N_2238,N_2065,N_2130);
and U2239 (N_2239,N_2028,N_2034);
and U2240 (N_2240,N_2197,N_2064);
xnor U2241 (N_2241,N_2108,N_2195);
nand U2242 (N_2242,N_2168,N_2035);
or U2243 (N_2243,N_2092,N_2036);
or U2244 (N_2244,N_2156,N_2080);
and U2245 (N_2245,N_2124,N_2151);
and U2246 (N_2246,N_2024,N_2076);
or U2247 (N_2247,N_2078,N_2039);
nand U2248 (N_2248,N_2057,N_2162);
xor U2249 (N_2249,N_2005,N_2167);
nor U2250 (N_2250,N_2044,N_2161);
xor U2251 (N_2251,N_2063,N_2134);
xor U2252 (N_2252,N_2052,N_2186);
nand U2253 (N_2253,N_2149,N_2084);
nand U2254 (N_2254,N_2116,N_2001);
xnor U2255 (N_2255,N_2090,N_2025);
and U2256 (N_2256,N_2093,N_2181);
nand U2257 (N_2257,N_2113,N_2089);
nor U2258 (N_2258,N_2015,N_2059);
nand U2259 (N_2259,N_2016,N_2187);
nand U2260 (N_2260,N_2097,N_2133);
nor U2261 (N_2261,N_2094,N_2054);
nor U2262 (N_2262,N_2058,N_2010);
and U2263 (N_2263,N_2071,N_2079);
nor U2264 (N_2264,N_2163,N_2172);
and U2265 (N_2265,N_2008,N_2037);
nand U2266 (N_2266,N_2023,N_2126);
and U2267 (N_2267,N_2171,N_2140);
xor U2268 (N_2268,N_2137,N_2074);
or U2269 (N_2269,N_2048,N_2099);
nor U2270 (N_2270,N_2007,N_2159);
or U2271 (N_2271,N_2000,N_2046);
and U2272 (N_2272,N_2014,N_2127);
nand U2273 (N_2273,N_2098,N_2170);
nor U2274 (N_2274,N_2043,N_2139);
and U2275 (N_2275,N_2013,N_2061);
nand U2276 (N_2276,N_2096,N_2183);
or U2277 (N_2277,N_2020,N_2019);
nor U2278 (N_2278,N_2060,N_2009);
and U2279 (N_2279,N_2182,N_2199);
or U2280 (N_2280,N_2152,N_2132);
and U2281 (N_2281,N_2083,N_2068);
and U2282 (N_2282,N_2088,N_2031);
or U2283 (N_2283,N_2003,N_2150);
nand U2284 (N_2284,N_2165,N_2164);
and U2285 (N_2285,N_2109,N_2082);
and U2286 (N_2286,N_2067,N_2017);
nand U2287 (N_2287,N_2102,N_2144);
nand U2288 (N_2288,N_2166,N_2086);
nand U2289 (N_2289,N_2129,N_2033);
nor U2290 (N_2290,N_2193,N_2056);
or U2291 (N_2291,N_2189,N_2110);
or U2292 (N_2292,N_2135,N_2041);
nor U2293 (N_2293,N_2040,N_2087);
and U2294 (N_2294,N_2022,N_2194);
nor U2295 (N_2295,N_2173,N_2055);
nor U2296 (N_2296,N_2143,N_2174);
nor U2297 (N_2297,N_2145,N_2196);
and U2298 (N_2298,N_2077,N_2091);
or U2299 (N_2299,N_2177,N_2138);
nand U2300 (N_2300,N_2160,N_2172);
nor U2301 (N_2301,N_2103,N_2175);
nor U2302 (N_2302,N_2195,N_2005);
nand U2303 (N_2303,N_2000,N_2128);
or U2304 (N_2304,N_2185,N_2077);
and U2305 (N_2305,N_2123,N_2063);
xnor U2306 (N_2306,N_2090,N_2127);
and U2307 (N_2307,N_2032,N_2181);
nand U2308 (N_2308,N_2104,N_2012);
nand U2309 (N_2309,N_2138,N_2193);
nand U2310 (N_2310,N_2022,N_2114);
nor U2311 (N_2311,N_2047,N_2055);
nor U2312 (N_2312,N_2136,N_2005);
nand U2313 (N_2313,N_2016,N_2160);
or U2314 (N_2314,N_2154,N_2070);
xnor U2315 (N_2315,N_2093,N_2059);
nor U2316 (N_2316,N_2014,N_2106);
nor U2317 (N_2317,N_2009,N_2092);
xnor U2318 (N_2318,N_2045,N_2142);
or U2319 (N_2319,N_2053,N_2005);
nand U2320 (N_2320,N_2081,N_2134);
nand U2321 (N_2321,N_2000,N_2137);
or U2322 (N_2322,N_2110,N_2010);
or U2323 (N_2323,N_2169,N_2097);
nor U2324 (N_2324,N_2080,N_2162);
or U2325 (N_2325,N_2077,N_2089);
and U2326 (N_2326,N_2063,N_2080);
or U2327 (N_2327,N_2013,N_2187);
or U2328 (N_2328,N_2114,N_2053);
nor U2329 (N_2329,N_2143,N_2186);
and U2330 (N_2330,N_2091,N_2000);
and U2331 (N_2331,N_2128,N_2147);
and U2332 (N_2332,N_2136,N_2194);
nor U2333 (N_2333,N_2139,N_2055);
and U2334 (N_2334,N_2007,N_2043);
nand U2335 (N_2335,N_2029,N_2071);
or U2336 (N_2336,N_2053,N_2113);
and U2337 (N_2337,N_2180,N_2098);
or U2338 (N_2338,N_2076,N_2023);
xor U2339 (N_2339,N_2101,N_2163);
nand U2340 (N_2340,N_2188,N_2160);
nor U2341 (N_2341,N_2125,N_2132);
nor U2342 (N_2342,N_2019,N_2139);
nand U2343 (N_2343,N_2189,N_2157);
nand U2344 (N_2344,N_2110,N_2193);
and U2345 (N_2345,N_2109,N_2177);
nor U2346 (N_2346,N_2148,N_2191);
nor U2347 (N_2347,N_2169,N_2040);
or U2348 (N_2348,N_2178,N_2003);
nor U2349 (N_2349,N_2176,N_2180);
nand U2350 (N_2350,N_2140,N_2168);
nand U2351 (N_2351,N_2055,N_2007);
nor U2352 (N_2352,N_2071,N_2098);
nand U2353 (N_2353,N_2144,N_2140);
nand U2354 (N_2354,N_2058,N_2080);
and U2355 (N_2355,N_2063,N_2059);
nor U2356 (N_2356,N_2021,N_2091);
and U2357 (N_2357,N_2126,N_2027);
and U2358 (N_2358,N_2033,N_2073);
or U2359 (N_2359,N_2129,N_2026);
nand U2360 (N_2360,N_2085,N_2111);
nor U2361 (N_2361,N_2047,N_2015);
nor U2362 (N_2362,N_2129,N_2092);
or U2363 (N_2363,N_2085,N_2074);
nor U2364 (N_2364,N_2147,N_2113);
and U2365 (N_2365,N_2080,N_2133);
and U2366 (N_2366,N_2026,N_2154);
nand U2367 (N_2367,N_2085,N_2012);
and U2368 (N_2368,N_2048,N_2010);
and U2369 (N_2369,N_2114,N_2098);
and U2370 (N_2370,N_2137,N_2183);
and U2371 (N_2371,N_2140,N_2030);
xnor U2372 (N_2372,N_2048,N_2102);
nor U2373 (N_2373,N_2142,N_2100);
nor U2374 (N_2374,N_2004,N_2084);
or U2375 (N_2375,N_2088,N_2007);
or U2376 (N_2376,N_2055,N_2161);
nor U2377 (N_2377,N_2127,N_2158);
nand U2378 (N_2378,N_2011,N_2152);
or U2379 (N_2379,N_2170,N_2015);
or U2380 (N_2380,N_2075,N_2154);
nor U2381 (N_2381,N_2162,N_2048);
xnor U2382 (N_2382,N_2131,N_2145);
or U2383 (N_2383,N_2020,N_2055);
nor U2384 (N_2384,N_2084,N_2121);
nand U2385 (N_2385,N_2072,N_2080);
nor U2386 (N_2386,N_2077,N_2187);
nand U2387 (N_2387,N_2173,N_2143);
xor U2388 (N_2388,N_2029,N_2073);
and U2389 (N_2389,N_2035,N_2150);
nand U2390 (N_2390,N_2008,N_2099);
xor U2391 (N_2391,N_2082,N_2117);
nand U2392 (N_2392,N_2196,N_2182);
nor U2393 (N_2393,N_2051,N_2138);
nor U2394 (N_2394,N_2174,N_2027);
and U2395 (N_2395,N_2006,N_2186);
nor U2396 (N_2396,N_2107,N_2099);
or U2397 (N_2397,N_2181,N_2143);
nand U2398 (N_2398,N_2149,N_2003);
nor U2399 (N_2399,N_2148,N_2029);
or U2400 (N_2400,N_2350,N_2250);
nand U2401 (N_2401,N_2368,N_2318);
and U2402 (N_2402,N_2290,N_2258);
or U2403 (N_2403,N_2253,N_2221);
nor U2404 (N_2404,N_2305,N_2248);
nand U2405 (N_2405,N_2261,N_2239);
and U2406 (N_2406,N_2230,N_2203);
or U2407 (N_2407,N_2343,N_2349);
and U2408 (N_2408,N_2267,N_2210);
xor U2409 (N_2409,N_2200,N_2390);
nor U2410 (N_2410,N_2269,N_2291);
xnor U2411 (N_2411,N_2331,N_2310);
and U2412 (N_2412,N_2280,N_2322);
nor U2413 (N_2413,N_2378,N_2391);
and U2414 (N_2414,N_2286,N_2375);
nor U2415 (N_2415,N_2279,N_2355);
and U2416 (N_2416,N_2333,N_2303);
nor U2417 (N_2417,N_2339,N_2365);
and U2418 (N_2418,N_2351,N_2335);
nand U2419 (N_2419,N_2278,N_2311);
nor U2420 (N_2420,N_2348,N_2356);
or U2421 (N_2421,N_2263,N_2329);
nor U2422 (N_2422,N_2327,N_2227);
and U2423 (N_2423,N_2219,N_2298);
or U2424 (N_2424,N_2377,N_2212);
nor U2425 (N_2425,N_2271,N_2247);
xor U2426 (N_2426,N_2274,N_2376);
or U2427 (N_2427,N_2340,N_2372);
nor U2428 (N_2428,N_2265,N_2215);
and U2429 (N_2429,N_2346,N_2284);
nand U2430 (N_2430,N_2326,N_2262);
or U2431 (N_2431,N_2216,N_2363);
or U2432 (N_2432,N_2381,N_2226);
and U2433 (N_2433,N_2234,N_2379);
or U2434 (N_2434,N_2320,N_2358);
and U2435 (N_2435,N_2316,N_2220);
xnor U2436 (N_2436,N_2332,N_2289);
and U2437 (N_2437,N_2205,N_2362);
nor U2438 (N_2438,N_2243,N_2223);
nor U2439 (N_2439,N_2347,N_2370);
or U2440 (N_2440,N_2233,N_2206);
nor U2441 (N_2441,N_2244,N_2224);
and U2442 (N_2442,N_2392,N_2313);
nand U2443 (N_2443,N_2231,N_2341);
and U2444 (N_2444,N_2395,N_2360);
or U2445 (N_2445,N_2306,N_2384);
nand U2446 (N_2446,N_2256,N_2299);
nand U2447 (N_2447,N_2344,N_2204);
or U2448 (N_2448,N_2213,N_2389);
or U2449 (N_2449,N_2308,N_2345);
nand U2450 (N_2450,N_2398,N_2382);
and U2451 (N_2451,N_2240,N_2251);
nand U2452 (N_2452,N_2321,N_2374);
and U2453 (N_2453,N_2276,N_2324);
or U2454 (N_2454,N_2285,N_2260);
and U2455 (N_2455,N_2209,N_2317);
xor U2456 (N_2456,N_2287,N_2386);
or U2457 (N_2457,N_2367,N_2246);
nand U2458 (N_2458,N_2228,N_2292);
or U2459 (N_2459,N_2337,N_2396);
nor U2460 (N_2460,N_2369,N_2334);
xor U2461 (N_2461,N_2307,N_2301);
and U2462 (N_2462,N_2393,N_2387);
nor U2463 (N_2463,N_2353,N_2245);
or U2464 (N_2464,N_2217,N_2366);
nand U2465 (N_2465,N_2238,N_2211);
nor U2466 (N_2466,N_2380,N_2295);
and U2467 (N_2467,N_2202,N_2259);
nand U2468 (N_2468,N_2338,N_2361);
and U2469 (N_2469,N_2328,N_2241);
xnor U2470 (N_2470,N_2236,N_2300);
nand U2471 (N_2471,N_2270,N_2237);
nor U2472 (N_2472,N_2275,N_2249);
xnor U2473 (N_2473,N_2214,N_2357);
nand U2474 (N_2474,N_2297,N_2325);
and U2475 (N_2475,N_2371,N_2399);
and U2476 (N_2476,N_2277,N_2232);
and U2477 (N_2477,N_2373,N_2359);
nor U2478 (N_2478,N_2388,N_2254);
nor U2479 (N_2479,N_2342,N_2304);
or U2480 (N_2480,N_2394,N_2352);
xnor U2481 (N_2481,N_2312,N_2354);
nor U2482 (N_2482,N_2266,N_2283);
or U2483 (N_2483,N_2314,N_2257);
or U2484 (N_2484,N_2235,N_2229);
xor U2485 (N_2485,N_2208,N_2225);
and U2486 (N_2486,N_2383,N_2272);
nor U2487 (N_2487,N_2364,N_2268);
and U2488 (N_2488,N_2296,N_2273);
nor U2489 (N_2489,N_2222,N_2264);
nor U2490 (N_2490,N_2207,N_2252);
and U2491 (N_2491,N_2319,N_2309);
and U2492 (N_2492,N_2323,N_2385);
and U2493 (N_2493,N_2288,N_2201);
or U2494 (N_2494,N_2255,N_2293);
nand U2495 (N_2495,N_2294,N_2336);
nor U2496 (N_2496,N_2218,N_2330);
or U2497 (N_2497,N_2242,N_2281);
nand U2498 (N_2498,N_2302,N_2282);
and U2499 (N_2499,N_2397,N_2315);
and U2500 (N_2500,N_2326,N_2283);
nor U2501 (N_2501,N_2394,N_2354);
and U2502 (N_2502,N_2389,N_2308);
nor U2503 (N_2503,N_2221,N_2302);
nand U2504 (N_2504,N_2277,N_2215);
nand U2505 (N_2505,N_2236,N_2263);
nor U2506 (N_2506,N_2247,N_2384);
xnor U2507 (N_2507,N_2347,N_2208);
and U2508 (N_2508,N_2232,N_2380);
and U2509 (N_2509,N_2217,N_2348);
nand U2510 (N_2510,N_2243,N_2398);
nor U2511 (N_2511,N_2310,N_2298);
nor U2512 (N_2512,N_2287,N_2210);
nor U2513 (N_2513,N_2395,N_2269);
and U2514 (N_2514,N_2290,N_2372);
xnor U2515 (N_2515,N_2217,N_2309);
and U2516 (N_2516,N_2361,N_2370);
nor U2517 (N_2517,N_2279,N_2330);
and U2518 (N_2518,N_2229,N_2312);
nand U2519 (N_2519,N_2276,N_2249);
xnor U2520 (N_2520,N_2390,N_2294);
or U2521 (N_2521,N_2343,N_2208);
or U2522 (N_2522,N_2220,N_2313);
xnor U2523 (N_2523,N_2216,N_2320);
and U2524 (N_2524,N_2344,N_2385);
or U2525 (N_2525,N_2280,N_2276);
or U2526 (N_2526,N_2383,N_2349);
or U2527 (N_2527,N_2373,N_2233);
nor U2528 (N_2528,N_2360,N_2270);
and U2529 (N_2529,N_2203,N_2236);
nand U2530 (N_2530,N_2276,N_2315);
nor U2531 (N_2531,N_2360,N_2399);
nand U2532 (N_2532,N_2316,N_2396);
nor U2533 (N_2533,N_2331,N_2362);
or U2534 (N_2534,N_2382,N_2321);
nor U2535 (N_2535,N_2241,N_2286);
nand U2536 (N_2536,N_2269,N_2325);
and U2537 (N_2537,N_2364,N_2371);
or U2538 (N_2538,N_2318,N_2367);
nand U2539 (N_2539,N_2367,N_2350);
and U2540 (N_2540,N_2298,N_2320);
nand U2541 (N_2541,N_2201,N_2301);
or U2542 (N_2542,N_2365,N_2323);
and U2543 (N_2543,N_2297,N_2206);
and U2544 (N_2544,N_2266,N_2343);
or U2545 (N_2545,N_2310,N_2241);
nor U2546 (N_2546,N_2390,N_2385);
and U2547 (N_2547,N_2245,N_2329);
nand U2548 (N_2548,N_2256,N_2384);
or U2549 (N_2549,N_2209,N_2274);
or U2550 (N_2550,N_2379,N_2208);
or U2551 (N_2551,N_2257,N_2225);
nor U2552 (N_2552,N_2275,N_2289);
nor U2553 (N_2553,N_2360,N_2398);
and U2554 (N_2554,N_2258,N_2368);
xor U2555 (N_2555,N_2346,N_2369);
and U2556 (N_2556,N_2241,N_2292);
or U2557 (N_2557,N_2332,N_2304);
or U2558 (N_2558,N_2212,N_2359);
or U2559 (N_2559,N_2302,N_2281);
nand U2560 (N_2560,N_2313,N_2324);
nand U2561 (N_2561,N_2398,N_2311);
nor U2562 (N_2562,N_2256,N_2265);
nor U2563 (N_2563,N_2388,N_2315);
nor U2564 (N_2564,N_2236,N_2301);
nor U2565 (N_2565,N_2270,N_2364);
nand U2566 (N_2566,N_2260,N_2354);
nor U2567 (N_2567,N_2253,N_2301);
xnor U2568 (N_2568,N_2354,N_2261);
and U2569 (N_2569,N_2223,N_2252);
and U2570 (N_2570,N_2332,N_2348);
nor U2571 (N_2571,N_2304,N_2354);
and U2572 (N_2572,N_2283,N_2244);
or U2573 (N_2573,N_2313,N_2301);
and U2574 (N_2574,N_2307,N_2360);
or U2575 (N_2575,N_2295,N_2215);
and U2576 (N_2576,N_2395,N_2337);
or U2577 (N_2577,N_2260,N_2353);
and U2578 (N_2578,N_2360,N_2295);
or U2579 (N_2579,N_2248,N_2257);
nand U2580 (N_2580,N_2339,N_2399);
xor U2581 (N_2581,N_2262,N_2394);
and U2582 (N_2582,N_2203,N_2271);
nand U2583 (N_2583,N_2306,N_2211);
xor U2584 (N_2584,N_2359,N_2382);
nand U2585 (N_2585,N_2229,N_2244);
nor U2586 (N_2586,N_2285,N_2274);
nor U2587 (N_2587,N_2237,N_2384);
and U2588 (N_2588,N_2389,N_2298);
nand U2589 (N_2589,N_2366,N_2346);
nand U2590 (N_2590,N_2252,N_2369);
nand U2591 (N_2591,N_2241,N_2205);
or U2592 (N_2592,N_2352,N_2313);
and U2593 (N_2593,N_2296,N_2266);
nand U2594 (N_2594,N_2230,N_2315);
and U2595 (N_2595,N_2235,N_2224);
xor U2596 (N_2596,N_2360,N_2334);
nand U2597 (N_2597,N_2342,N_2272);
nand U2598 (N_2598,N_2245,N_2271);
nor U2599 (N_2599,N_2291,N_2359);
and U2600 (N_2600,N_2446,N_2542);
nand U2601 (N_2601,N_2473,N_2476);
or U2602 (N_2602,N_2411,N_2486);
xor U2603 (N_2603,N_2595,N_2552);
or U2604 (N_2604,N_2483,N_2417);
xnor U2605 (N_2605,N_2447,N_2481);
and U2606 (N_2606,N_2455,N_2531);
xor U2607 (N_2607,N_2539,N_2457);
xnor U2608 (N_2608,N_2571,N_2579);
nor U2609 (N_2609,N_2456,N_2431);
xor U2610 (N_2610,N_2559,N_2444);
nor U2611 (N_2611,N_2449,N_2545);
xor U2612 (N_2612,N_2554,N_2511);
nand U2613 (N_2613,N_2465,N_2472);
nand U2614 (N_2614,N_2568,N_2450);
or U2615 (N_2615,N_2546,N_2520);
nor U2616 (N_2616,N_2532,N_2436);
nand U2617 (N_2617,N_2421,N_2522);
nand U2618 (N_2618,N_2404,N_2509);
xnor U2619 (N_2619,N_2426,N_2562);
nor U2620 (N_2620,N_2548,N_2519);
nor U2621 (N_2621,N_2504,N_2547);
nand U2622 (N_2622,N_2405,N_2493);
or U2623 (N_2623,N_2560,N_2463);
nand U2624 (N_2624,N_2489,N_2445);
nor U2625 (N_2625,N_2442,N_2402);
xnor U2626 (N_2626,N_2435,N_2533);
nor U2627 (N_2627,N_2543,N_2575);
and U2628 (N_2628,N_2495,N_2517);
nor U2629 (N_2629,N_2551,N_2488);
and U2630 (N_2630,N_2585,N_2506);
nand U2631 (N_2631,N_2485,N_2528);
nor U2632 (N_2632,N_2516,N_2423);
and U2633 (N_2633,N_2535,N_2410);
nand U2634 (N_2634,N_2537,N_2412);
nor U2635 (N_2635,N_2514,N_2508);
nor U2636 (N_2636,N_2487,N_2544);
nor U2637 (N_2637,N_2497,N_2464);
nand U2638 (N_2638,N_2594,N_2430);
and U2639 (N_2639,N_2593,N_2586);
and U2640 (N_2640,N_2433,N_2418);
nor U2641 (N_2641,N_2570,N_2467);
xor U2642 (N_2642,N_2498,N_2452);
nor U2643 (N_2643,N_2408,N_2471);
and U2644 (N_2644,N_2577,N_2561);
or U2645 (N_2645,N_2490,N_2413);
and U2646 (N_2646,N_2534,N_2499);
nor U2647 (N_2647,N_2584,N_2400);
xnor U2648 (N_2648,N_2549,N_2466);
nor U2649 (N_2649,N_2478,N_2429);
xor U2650 (N_2650,N_2441,N_2448);
nand U2651 (N_2651,N_2454,N_2555);
or U2652 (N_2652,N_2420,N_2540);
or U2653 (N_2653,N_2496,N_2597);
or U2654 (N_2654,N_2461,N_2583);
nand U2655 (N_2655,N_2576,N_2563);
or U2656 (N_2656,N_2529,N_2470);
nand U2657 (N_2657,N_2492,N_2425);
nor U2658 (N_2658,N_2587,N_2590);
xnor U2659 (N_2659,N_2515,N_2403);
nor U2660 (N_2660,N_2494,N_2513);
xnor U2661 (N_2661,N_2558,N_2591);
and U2662 (N_2662,N_2530,N_2428);
nor U2663 (N_2663,N_2572,N_2574);
and U2664 (N_2664,N_2439,N_2424);
or U2665 (N_2665,N_2414,N_2521);
nand U2666 (N_2666,N_2419,N_2475);
nand U2667 (N_2667,N_2458,N_2550);
nor U2668 (N_2668,N_2500,N_2580);
or U2669 (N_2669,N_2427,N_2599);
nand U2670 (N_2670,N_2588,N_2567);
xor U2671 (N_2671,N_2437,N_2582);
and U2672 (N_2672,N_2415,N_2407);
nand U2673 (N_2673,N_2512,N_2479);
xor U2674 (N_2674,N_2510,N_2527);
or U2675 (N_2675,N_2503,N_2507);
and U2676 (N_2676,N_2526,N_2596);
xnor U2677 (N_2677,N_2460,N_2553);
nand U2678 (N_2678,N_2501,N_2443);
nand U2679 (N_2679,N_2440,N_2598);
nand U2680 (N_2680,N_2432,N_2523);
nor U2681 (N_2681,N_2453,N_2564);
or U2682 (N_2682,N_2491,N_2468);
or U2683 (N_2683,N_2518,N_2502);
nor U2684 (N_2684,N_2484,N_2556);
nand U2685 (N_2685,N_2401,N_2482);
nand U2686 (N_2686,N_2459,N_2474);
xnor U2687 (N_2687,N_2541,N_2581);
and U2688 (N_2688,N_2434,N_2569);
or U2689 (N_2689,N_2406,N_2477);
nand U2690 (N_2690,N_2416,N_2469);
nand U2691 (N_2691,N_2438,N_2565);
or U2692 (N_2692,N_2592,N_2557);
and U2693 (N_2693,N_2573,N_2422);
or U2694 (N_2694,N_2409,N_2589);
or U2695 (N_2695,N_2566,N_2536);
and U2696 (N_2696,N_2525,N_2480);
nor U2697 (N_2697,N_2524,N_2578);
nand U2698 (N_2698,N_2451,N_2505);
or U2699 (N_2699,N_2538,N_2462);
xnor U2700 (N_2700,N_2537,N_2491);
xor U2701 (N_2701,N_2478,N_2597);
nor U2702 (N_2702,N_2404,N_2595);
nand U2703 (N_2703,N_2465,N_2563);
nand U2704 (N_2704,N_2499,N_2531);
xnor U2705 (N_2705,N_2464,N_2597);
nor U2706 (N_2706,N_2459,N_2522);
and U2707 (N_2707,N_2575,N_2462);
and U2708 (N_2708,N_2475,N_2552);
or U2709 (N_2709,N_2417,N_2402);
nand U2710 (N_2710,N_2486,N_2477);
nand U2711 (N_2711,N_2568,N_2473);
nand U2712 (N_2712,N_2590,N_2588);
xor U2713 (N_2713,N_2439,N_2418);
or U2714 (N_2714,N_2495,N_2526);
nand U2715 (N_2715,N_2561,N_2424);
and U2716 (N_2716,N_2540,N_2558);
nand U2717 (N_2717,N_2460,N_2516);
and U2718 (N_2718,N_2404,N_2479);
nand U2719 (N_2719,N_2427,N_2500);
or U2720 (N_2720,N_2577,N_2586);
or U2721 (N_2721,N_2414,N_2596);
or U2722 (N_2722,N_2440,N_2482);
nand U2723 (N_2723,N_2413,N_2439);
xor U2724 (N_2724,N_2585,N_2464);
nand U2725 (N_2725,N_2445,N_2402);
nand U2726 (N_2726,N_2429,N_2539);
and U2727 (N_2727,N_2532,N_2428);
or U2728 (N_2728,N_2454,N_2589);
or U2729 (N_2729,N_2548,N_2406);
or U2730 (N_2730,N_2579,N_2490);
or U2731 (N_2731,N_2494,N_2537);
xnor U2732 (N_2732,N_2474,N_2463);
and U2733 (N_2733,N_2592,N_2525);
or U2734 (N_2734,N_2404,N_2447);
and U2735 (N_2735,N_2545,N_2523);
and U2736 (N_2736,N_2471,N_2559);
xnor U2737 (N_2737,N_2417,N_2450);
and U2738 (N_2738,N_2476,N_2523);
nor U2739 (N_2739,N_2415,N_2526);
nand U2740 (N_2740,N_2567,N_2546);
nand U2741 (N_2741,N_2556,N_2543);
or U2742 (N_2742,N_2521,N_2513);
nand U2743 (N_2743,N_2570,N_2517);
nand U2744 (N_2744,N_2455,N_2589);
xnor U2745 (N_2745,N_2440,N_2421);
or U2746 (N_2746,N_2401,N_2419);
nand U2747 (N_2747,N_2598,N_2550);
nand U2748 (N_2748,N_2586,N_2569);
and U2749 (N_2749,N_2441,N_2510);
nor U2750 (N_2750,N_2562,N_2594);
and U2751 (N_2751,N_2481,N_2438);
or U2752 (N_2752,N_2423,N_2454);
or U2753 (N_2753,N_2525,N_2444);
and U2754 (N_2754,N_2533,N_2536);
nor U2755 (N_2755,N_2531,N_2512);
and U2756 (N_2756,N_2492,N_2417);
or U2757 (N_2757,N_2455,N_2564);
nor U2758 (N_2758,N_2461,N_2467);
nand U2759 (N_2759,N_2455,N_2421);
and U2760 (N_2760,N_2506,N_2434);
and U2761 (N_2761,N_2447,N_2471);
nor U2762 (N_2762,N_2426,N_2580);
nand U2763 (N_2763,N_2513,N_2464);
nor U2764 (N_2764,N_2582,N_2519);
nor U2765 (N_2765,N_2434,N_2556);
nand U2766 (N_2766,N_2506,N_2543);
nor U2767 (N_2767,N_2580,N_2478);
nor U2768 (N_2768,N_2501,N_2503);
nand U2769 (N_2769,N_2535,N_2460);
nor U2770 (N_2770,N_2475,N_2474);
xor U2771 (N_2771,N_2411,N_2560);
nor U2772 (N_2772,N_2560,N_2578);
and U2773 (N_2773,N_2428,N_2587);
nand U2774 (N_2774,N_2446,N_2543);
and U2775 (N_2775,N_2589,N_2485);
nor U2776 (N_2776,N_2459,N_2591);
and U2777 (N_2777,N_2595,N_2472);
and U2778 (N_2778,N_2446,N_2574);
nand U2779 (N_2779,N_2493,N_2579);
nand U2780 (N_2780,N_2508,N_2436);
nor U2781 (N_2781,N_2523,N_2412);
and U2782 (N_2782,N_2400,N_2481);
or U2783 (N_2783,N_2544,N_2457);
nor U2784 (N_2784,N_2500,N_2412);
nor U2785 (N_2785,N_2538,N_2502);
and U2786 (N_2786,N_2426,N_2466);
and U2787 (N_2787,N_2441,N_2415);
xor U2788 (N_2788,N_2504,N_2524);
nor U2789 (N_2789,N_2558,N_2545);
and U2790 (N_2790,N_2478,N_2451);
or U2791 (N_2791,N_2545,N_2586);
nor U2792 (N_2792,N_2578,N_2484);
or U2793 (N_2793,N_2456,N_2488);
and U2794 (N_2794,N_2403,N_2488);
or U2795 (N_2795,N_2463,N_2464);
or U2796 (N_2796,N_2471,N_2568);
nand U2797 (N_2797,N_2448,N_2444);
nor U2798 (N_2798,N_2555,N_2536);
or U2799 (N_2799,N_2556,N_2475);
nand U2800 (N_2800,N_2652,N_2623);
nor U2801 (N_2801,N_2627,N_2712);
nand U2802 (N_2802,N_2798,N_2781);
nor U2803 (N_2803,N_2646,N_2799);
and U2804 (N_2804,N_2702,N_2654);
nand U2805 (N_2805,N_2665,N_2688);
and U2806 (N_2806,N_2767,N_2607);
and U2807 (N_2807,N_2669,N_2752);
and U2808 (N_2808,N_2662,N_2649);
or U2809 (N_2809,N_2730,N_2610);
and U2810 (N_2810,N_2685,N_2797);
nand U2811 (N_2811,N_2778,N_2653);
or U2812 (N_2812,N_2658,N_2787);
xor U2813 (N_2813,N_2786,N_2642);
and U2814 (N_2814,N_2793,N_2727);
and U2815 (N_2815,N_2639,N_2760);
or U2816 (N_2816,N_2766,N_2636);
or U2817 (N_2817,N_2698,N_2717);
nor U2818 (N_2818,N_2625,N_2633);
nor U2819 (N_2819,N_2670,N_2736);
nand U2820 (N_2820,N_2635,N_2783);
or U2821 (N_2821,N_2731,N_2694);
xnor U2822 (N_2822,N_2743,N_2608);
nor U2823 (N_2823,N_2631,N_2666);
or U2824 (N_2824,N_2634,N_2721);
and U2825 (N_2825,N_2701,N_2764);
and U2826 (N_2826,N_2660,N_2710);
or U2827 (N_2827,N_2703,N_2732);
nand U2828 (N_2828,N_2720,N_2740);
and U2829 (N_2829,N_2711,N_2661);
nor U2830 (N_2830,N_2606,N_2749);
and U2831 (N_2831,N_2638,N_2621);
and U2832 (N_2832,N_2725,N_2728);
nand U2833 (N_2833,N_2715,N_2656);
nand U2834 (N_2834,N_2708,N_2773);
nor U2835 (N_2835,N_2705,N_2724);
nor U2836 (N_2836,N_2668,N_2671);
and U2837 (N_2837,N_2691,N_2696);
or U2838 (N_2838,N_2651,N_2689);
nor U2839 (N_2839,N_2784,N_2726);
and U2840 (N_2840,N_2686,N_2673);
nor U2841 (N_2841,N_2618,N_2706);
and U2842 (N_2842,N_2629,N_2716);
nand U2843 (N_2843,N_2782,N_2640);
and U2844 (N_2844,N_2744,N_2707);
or U2845 (N_2845,N_2775,N_2794);
and U2846 (N_2846,N_2776,N_2617);
and U2847 (N_2847,N_2675,N_2619);
nor U2848 (N_2848,N_2704,N_2613);
nor U2849 (N_2849,N_2747,N_2612);
or U2850 (N_2850,N_2687,N_2763);
and U2851 (N_2851,N_2745,N_2758);
nand U2852 (N_2852,N_2690,N_2790);
or U2853 (N_2853,N_2677,N_2604);
or U2854 (N_2854,N_2734,N_2682);
and U2855 (N_2855,N_2765,N_2624);
and U2856 (N_2856,N_2792,N_2667);
nand U2857 (N_2857,N_2648,N_2672);
or U2858 (N_2858,N_2630,N_2615);
nand U2859 (N_2859,N_2733,N_2679);
and U2860 (N_2860,N_2699,N_2754);
or U2861 (N_2861,N_2628,N_2779);
nand U2862 (N_2862,N_2723,N_2681);
nand U2863 (N_2863,N_2788,N_2746);
and U2864 (N_2864,N_2637,N_2714);
nand U2865 (N_2865,N_2674,N_2692);
nand U2866 (N_2866,N_2693,N_2795);
nor U2867 (N_2867,N_2789,N_2626);
or U2868 (N_2868,N_2700,N_2761);
or U2869 (N_2869,N_2601,N_2683);
and U2870 (N_2870,N_2614,N_2753);
or U2871 (N_2871,N_2791,N_2709);
and U2872 (N_2872,N_2785,N_2735);
or U2873 (N_2873,N_2663,N_2718);
or U2874 (N_2874,N_2741,N_2739);
nand U2875 (N_2875,N_2684,N_2645);
nor U2876 (N_2876,N_2769,N_2622);
xnor U2877 (N_2877,N_2603,N_2737);
and U2878 (N_2878,N_2697,N_2774);
nor U2879 (N_2879,N_2762,N_2609);
xor U2880 (N_2880,N_2655,N_2605);
and U2881 (N_2881,N_2664,N_2713);
and U2882 (N_2882,N_2770,N_2678);
nand U2883 (N_2883,N_2751,N_2657);
and U2884 (N_2884,N_2719,N_2644);
nand U2885 (N_2885,N_2641,N_2650);
and U2886 (N_2886,N_2600,N_2772);
or U2887 (N_2887,N_2755,N_2620);
nand U2888 (N_2888,N_2695,N_2676);
nor U2889 (N_2889,N_2722,N_2759);
nor U2890 (N_2890,N_2748,N_2742);
nand U2891 (N_2891,N_2738,N_2643);
nand U2892 (N_2892,N_2771,N_2680);
and U2893 (N_2893,N_2611,N_2768);
xor U2894 (N_2894,N_2616,N_2647);
and U2895 (N_2895,N_2780,N_2757);
nor U2896 (N_2896,N_2632,N_2729);
and U2897 (N_2897,N_2777,N_2756);
nor U2898 (N_2898,N_2659,N_2796);
or U2899 (N_2899,N_2750,N_2602);
or U2900 (N_2900,N_2722,N_2768);
xor U2901 (N_2901,N_2666,N_2653);
nor U2902 (N_2902,N_2665,N_2766);
nand U2903 (N_2903,N_2698,N_2644);
or U2904 (N_2904,N_2627,N_2635);
nand U2905 (N_2905,N_2799,N_2612);
nor U2906 (N_2906,N_2619,N_2762);
nor U2907 (N_2907,N_2753,N_2615);
or U2908 (N_2908,N_2641,N_2651);
nor U2909 (N_2909,N_2611,N_2716);
nor U2910 (N_2910,N_2748,N_2799);
or U2911 (N_2911,N_2615,N_2775);
or U2912 (N_2912,N_2671,N_2611);
nor U2913 (N_2913,N_2602,N_2694);
nor U2914 (N_2914,N_2610,N_2658);
nand U2915 (N_2915,N_2717,N_2701);
and U2916 (N_2916,N_2600,N_2743);
and U2917 (N_2917,N_2768,N_2680);
nor U2918 (N_2918,N_2690,N_2760);
xor U2919 (N_2919,N_2695,N_2798);
nor U2920 (N_2920,N_2624,N_2754);
or U2921 (N_2921,N_2733,N_2626);
xnor U2922 (N_2922,N_2611,N_2651);
nand U2923 (N_2923,N_2611,N_2726);
nor U2924 (N_2924,N_2749,N_2781);
and U2925 (N_2925,N_2680,N_2663);
nor U2926 (N_2926,N_2643,N_2628);
nor U2927 (N_2927,N_2769,N_2643);
and U2928 (N_2928,N_2696,N_2614);
and U2929 (N_2929,N_2760,N_2657);
and U2930 (N_2930,N_2793,N_2645);
and U2931 (N_2931,N_2685,N_2791);
xnor U2932 (N_2932,N_2724,N_2696);
and U2933 (N_2933,N_2620,N_2676);
and U2934 (N_2934,N_2612,N_2648);
and U2935 (N_2935,N_2625,N_2726);
nor U2936 (N_2936,N_2693,N_2635);
or U2937 (N_2937,N_2614,N_2798);
nand U2938 (N_2938,N_2660,N_2795);
xor U2939 (N_2939,N_2618,N_2775);
or U2940 (N_2940,N_2752,N_2794);
and U2941 (N_2941,N_2726,N_2742);
or U2942 (N_2942,N_2668,N_2697);
or U2943 (N_2943,N_2634,N_2711);
xnor U2944 (N_2944,N_2635,N_2725);
nand U2945 (N_2945,N_2664,N_2633);
nand U2946 (N_2946,N_2796,N_2780);
xnor U2947 (N_2947,N_2796,N_2775);
or U2948 (N_2948,N_2645,N_2744);
nor U2949 (N_2949,N_2619,N_2642);
nand U2950 (N_2950,N_2754,N_2771);
nand U2951 (N_2951,N_2775,N_2667);
or U2952 (N_2952,N_2745,N_2796);
nand U2953 (N_2953,N_2609,N_2721);
nand U2954 (N_2954,N_2649,N_2719);
or U2955 (N_2955,N_2605,N_2638);
nand U2956 (N_2956,N_2637,N_2729);
nor U2957 (N_2957,N_2633,N_2674);
nor U2958 (N_2958,N_2703,N_2710);
nand U2959 (N_2959,N_2702,N_2712);
nor U2960 (N_2960,N_2641,N_2726);
or U2961 (N_2961,N_2738,N_2668);
and U2962 (N_2962,N_2623,N_2614);
and U2963 (N_2963,N_2770,N_2727);
and U2964 (N_2964,N_2739,N_2767);
or U2965 (N_2965,N_2776,N_2707);
nand U2966 (N_2966,N_2649,N_2791);
nand U2967 (N_2967,N_2765,N_2727);
nand U2968 (N_2968,N_2607,N_2673);
or U2969 (N_2969,N_2717,N_2767);
nor U2970 (N_2970,N_2693,N_2750);
nand U2971 (N_2971,N_2666,N_2741);
and U2972 (N_2972,N_2625,N_2793);
or U2973 (N_2973,N_2616,N_2656);
or U2974 (N_2974,N_2742,N_2607);
or U2975 (N_2975,N_2786,N_2622);
nand U2976 (N_2976,N_2659,N_2645);
nand U2977 (N_2977,N_2609,N_2648);
and U2978 (N_2978,N_2700,N_2672);
and U2979 (N_2979,N_2758,N_2696);
nand U2980 (N_2980,N_2682,N_2630);
or U2981 (N_2981,N_2762,N_2636);
xor U2982 (N_2982,N_2788,N_2747);
and U2983 (N_2983,N_2668,N_2778);
nand U2984 (N_2984,N_2629,N_2796);
and U2985 (N_2985,N_2795,N_2798);
xor U2986 (N_2986,N_2731,N_2729);
or U2987 (N_2987,N_2622,N_2618);
nand U2988 (N_2988,N_2668,N_2637);
or U2989 (N_2989,N_2627,N_2604);
nand U2990 (N_2990,N_2794,N_2684);
nand U2991 (N_2991,N_2799,N_2772);
nor U2992 (N_2992,N_2746,N_2651);
nand U2993 (N_2993,N_2642,N_2756);
or U2994 (N_2994,N_2602,N_2643);
nand U2995 (N_2995,N_2741,N_2759);
nor U2996 (N_2996,N_2799,N_2688);
nor U2997 (N_2997,N_2695,N_2617);
nor U2998 (N_2998,N_2611,N_2676);
nor U2999 (N_2999,N_2684,N_2640);
and U3000 (N_3000,N_2884,N_2847);
nor U3001 (N_3001,N_2862,N_2958);
nor U3002 (N_3002,N_2904,N_2825);
nor U3003 (N_3003,N_2972,N_2898);
xor U3004 (N_3004,N_2960,N_2980);
xor U3005 (N_3005,N_2934,N_2883);
xnor U3006 (N_3006,N_2821,N_2956);
nor U3007 (N_3007,N_2803,N_2873);
and U3008 (N_3008,N_2870,N_2913);
or U3009 (N_3009,N_2952,N_2899);
and U3010 (N_3010,N_2811,N_2810);
nand U3011 (N_3011,N_2937,N_2919);
xor U3012 (N_3012,N_2943,N_2894);
xor U3013 (N_3013,N_2816,N_2912);
and U3014 (N_3014,N_2805,N_2858);
nand U3015 (N_3015,N_2926,N_2823);
nor U3016 (N_3016,N_2892,N_2879);
nand U3017 (N_3017,N_2981,N_2827);
and U3018 (N_3018,N_2880,N_2991);
nand U3019 (N_3019,N_2864,N_2804);
and U3020 (N_3020,N_2901,N_2973);
nor U3021 (N_3021,N_2959,N_2856);
nand U3022 (N_3022,N_2914,N_2846);
and U3023 (N_3023,N_2910,N_2970);
nor U3024 (N_3024,N_2951,N_2961);
nor U3025 (N_3025,N_2944,N_2971);
nor U3026 (N_3026,N_2963,N_2946);
or U3027 (N_3027,N_2834,N_2976);
or U3028 (N_3028,N_2917,N_2829);
nand U3029 (N_3029,N_2866,N_2838);
nand U3030 (N_3030,N_2988,N_2962);
nor U3031 (N_3031,N_2850,N_2822);
xor U3032 (N_3032,N_2877,N_2977);
nand U3033 (N_3033,N_2812,N_2888);
or U3034 (N_3034,N_2975,N_2818);
nor U3035 (N_3035,N_2852,N_2860);
or U3036 (N_3036,N_2923,N_2916);
or U3037 (N_3037,N_2964,N_2890);
or U3038 (N_3038,N_2885,N_2806);
and U3039 (N_3039,N_2876,N_2836);
nand U3040 (N_3040,N_2853,N_2839);
nand U3041 (N_3041,N_2927,N_2933);
or U3042 (N_3042,N_2887,N_2984);
nand U3043 (N_3043,N_2935,N_2993);
and U3044 (N_3044,N_2966,N_2807);
and U3045 (N_3045,N_2819,N_2979);
nand U3046 (N_3046,N_2896,N_2895);
nand U3047 (N_3047,N_2968,N_2999);
nand U3048 (N_3048,N_2936,N_2813);
nand U3049 (N_3049,N_2844,N_2945);
and U3050 (N_3050,N_2989,N_2982);
nand U3051 (N_3051,N_2831,N_2915);
and U3052 (N_3052,N_2848,N_2997);
nor U3053 (N_3053,N_2875,N_2872);
xnor U3054 (N_3054,N_2801,N_2865);
and U3055 (N_3055,N_2907,N_2837);
nand U3056 (N_3056,N_2863,N_2891);
nand U3057 (N_3057,N_2918,N_2928);
xor U3058 (N_3058,N_2881,N_2957);
and U3059 (N_3059,N_2974,N_2949);
nand U3060 (N_3060,N_2920,N_2802);
nor U3061 (N_3061,N_2845,N_2921);
nor U3062 (N_3062,N_2835,N_2830);
and U3063 (N_3063,N_2841,N_2931);
nand U3064 (N_3064,N_2965,N_2842);
or U3065 (N_3065,N_2940,N_2882);
nand U3066 (N_3066,N_2820,N_2828);
nand U3067 (N_3067,N_2843,N_2908);
nor U3068 (N_3068,N_2900,N_2800);
xnor U3069 (N_3069,N_2851,N_2947);
and U3070 (N_3070,N_2948,N_2817);
or U3071 (N_3071,N_2906,N_2808);
or U3072 (N_3072,N_2932,N_2857);
nor U3073 (N_3073,N_2994,N_2815);
nor U3074 (N_3074,N_2996,N_2983);
nand U3075 (N_3075,N_2998,N_2861);
nor U3076 (N_3076,N_2886,N_2897);
nand U3077 (N_3077,N_2840,N_2867);
or U3078 (N_3078,N_2909,N_2939);
xnor U3079 (N_3079,N_2995,N_2986);
nor U3080 (N_3080,N_2925,N_2969);
nand U3081 (N_3081,N_2878,N_2967);
and U3082 (N_3082,N_2950,N_2809);
nand U3083 (N_3083,N_2889,N_2833);
or U3084 (N_3084,N_2874,N_2871);
xnor U3085 (N_3085,N_2955,N_2824);
or U3086 (N_3086,N_2942,N_2814);
nor U3087 (N_3087,N_2987,N_2854);
or U3088 (N_3088,N_2868,N_2903);
and U3089 (N_3089,N_2941,N_2893);
and U3090 (N_3090,N_2902,N_2922);
nor U3091 (N_3091,N_2855,N_2954);
nand U3092 (N_3092,N_2859,N_2930);
or U3093 (N_3093,N_2849,N_2905);
or U3094 (N_3094,N_2938,N_2869);
and U3095 (N_3095,N_2953,N_2990);
nand U3096 (N_3096,N_2929,N_2826);
or U3097 (N_3097,N_2978,N_2832);
or U3098 (N_3098,N_2992,N_2924);
or U3099 (N_3099,N_2985,N_2911);
or U3100 (N_3100,N_2882,N_2987);
or U3101 (N_3101,N_2966,N_2925);
nor U3102 (N_3102,N_2856,N_2817);
nor U3103 (N_3103,N_2988,N_2955);
or U3104 (N_3104,N_2869,N_2822);
nor U3105 (N_3105,N_2986,N_2800);
and U3106 (N_3106,N_2900,N_2981);
and U3107 (N_3107,N_2802,N_2914);
nor U3108 (N_3108,N_2823,N_2940);
nand U3109 (N_3109,N_2851,N_2860);
and U3110 (N_3110,N_2945,N_2821);
nand U3111 (N_3111,N_2856,N_2870);
nor U3112 (N_3112,N_2816,N_2860);
and U3113 (N_3113,N_2882,N_2857);
nand U3114 (N_3114,N_2835,N_2827);
nor U3115 (N_3115,N_2995,N_2991);
and U3116 (N_3116,N_2834,N_2973);
nand U3117 (N_3117,N_2869,N_2990);
nor U3118 (N_3118,N_2962,N_2917);
and U3119 (N_3119,N_2816,N_2839);
nor U3120 (N_3120,N_2929,N_2870);
xor U3121 (N_3121,N_2931,N_2987);
xor U3122 (N_3122,N_2849,N_2970);
nor U3123 (N_3123,N_2914,N_2977);
or U3124 (N_3124,N_2946,N_2828);
or U3125 (N_3125,N_2955,N_2930);
nand U3126 (N_3126,N_2998,N_2899);
nor U3127 (N_3127,N_2968,N_2802);
or U3128 (N_3128,N_2931,N_2905);
or U3129 (N_3129,N_2918,N_2839);
nor U3130 (N_3130,N_2866,N_2878);
or U3131 (N_3131,N_2834,N_2843);
nor U3132 (N_3132,N_2952,N_2882);
xnor U3133 (N_3133,N_2911,N_2934);
or U3134 (N_3134,N_2946,N_2909);
or U3135 (N_3135,N_2851,N_2805);
or U3136 (N_3136,N_2843,N_2853);
nand U3137 (N_3137,N_2952,N_2805);
nor U3138 (N_3138,N_2807,N_2839);
and U3139 (N_3139,N_2994,N_2917);
nand U3140 (N_3140,N_2884,N_2863);
and U3141 (N_3141,N_2955,N_2941);
nand U3142 (N_3142,N_2945,N_2950);
nor U3143 (N_3143,N_2955,N_2946);
and U3144 (N_3144,N_2956,N_2805);
or U3145 (N_3145,N_2935,N_2965);
nor U3146 (N_3146,N_2909,N_2873);
or U3147 (N_3147,N_2898,N_2956);
xor U3148 (N_3148,N_2838,N_2890);
and U3149 (N_3149,N_2964,N_2862);
nand U3150 (N_3150,N_2890,N_2858);
nor U3151 (N_3151,N_2880,N_2848);
nand U3152 (N_3152,N_2864,N_2823);
nand U3153 (N_3153,N_2839,N_2887);
or U3154 (N_3154,N_2817,N_2868);
and U3155 (N_3155,N_2903,N_2978);
xor U3156 (N_3156,N_2894,N_2947);
nand U3157 (N_3157,N_2879,N_2988);
or U3158 (N_3158,N_2922,N_2903);
nor U3159 (N_3159,N_2825,N_2934);
nand U3160 (N_3160,N_2882,N_2823);
or U3161 (N_3161,N_2876,N_2973);
and U3162 (N_3162,N_2812,N_2844);
and U3163 (N_3163,N_2963,N_2869);
or U3164 (N_3164,N_2973,N_2997);
nand U3165 (N_3165,N_2953,N_2983);
and U3166 (N_3166,N_2850,N_2893);
xor U3167 (N_3167,N_2978,N_2811);
nand U3168 (N_3168,N_2912,N_2834);
and U3169 (N_3169,N_2941,N_2928);
nor U3170 (N_3170,N_2842,N_2929);
xnor U3171 (N_3171,N_2911,N_2979);
or U3172 (N_3172,N_2802,N_2818);
and U3173 (N_3173,N_2891,N_2860);
xor U3174 (N_3174,N_2849,N_2915);
nand U3175 (N_3175,N_2879,N_2835);
nand U3176 (N_3176,N_2942,N_2810);
and U3177 (N_3177,N_2881,N_2934);
and U3178 (N_3178,N_2930,N_2826);
and U3179 (N_3179,N_2800,N_2812);
xnor U3180 (N_3180,N_2882,N_2980);
nand U3181 (N_3181,N_2867,N_2832);
nor U3182 (N_3182,N_2835,N_2869);
nor U3183 (N_3183,N_2984,N_2921);
or U3184 (N_3184,N_2881,N_2814);
nand U3185 (N_3185,N_2991,N_2809);
nor U3186 (N_3186,N_2910,N_2969);
xor U3187 (N_3187,N_2885,N_2884);
or U3188 (N_3188,N_2952,N_2936);
xnor U3189 (N_3189,N_2933,N_2801);
or U3190 (N_3190,N_2876,N_2875);
or U3191 (N_3191,N_2802,N_2986);
or U3192 (N_3192,N_2862,N_2913);
nand U3193 (N_3193,N_2946,N_2850);
nor U3194 (N_3194,N_2839,N_2928);
nand U3195 (N_3195,N_2956,N_2839);
or U3196 (N_3196,N_2833,N_2839);
or U3197 (N_3197,N_2931,N_2897);
and U3198 (N_3198,N_2960,N_2884);
nand U3199 (N_3199,N_2983,N_2966);
and U3200 (N_3200,N_3111,N_3094);
or U3201 (N_3201,N_3127,N_3042);
nor U3202 (N_3202,N_3191,N_3133);
xnor U3203 (N_3203,N_3065,N_3087);
nor U3204 (N_3204,N_3125,N_3097);
nand U3205 (N_3205,N_3009,N_3106);
nor U3206 (N_3206,N_3145,N_3151);
and U3207 (N_3207,N_3136,N_3091);
nand U3208 (N_3208,N_3018,N_3013);
or U3209 (N_3209,N_3168,N_3195);
and U3210 (N_3210,N_3137,N_3135);
nand U3211 (N_3211,N_3131,N_3059);
nor U3212 (N_3212,N_3084,N_3175);
or U3213 (N_3213,N_3011,N_3001);
and U3214 (N_3214,N_3016,N_3024);
nor U3215 (N_3215,N_3003,N_3062);
nor U3216 (N_3216,N_3154,N_3165);
nand U3217 (N_3217,N_3002,N_3142);
and U3218 (N_3218,N_3104,N_3161);
nand U3219 (N_3219,N_3096,N_3132);
xnor U3220 (N_3220,N_3181,N_3032);
nor U3221 (N_3221,N_3082,N_3061);
nand U3222 (N_3222,N_3037,N_3031);
nor U3223 (N_3223,N_3078,N_3128);
or U3224 (N_3224,N_3140,N_3077);
nor U3225 (N_3225,N_3150,N_3085);
nor U3226 (N_3226,N_3089,N_3121);
nand U3227 (N_3227,N_3182,N_3178);
and U3228 (N_3228,N_3138,N_3147);
and U3229 (N_3229,N_3057,N_3199);
nand U3230 (N_3230,N_3039,N_3139);
nor U3231 (N_3231,N_3118,N_3083);
nand U3232 (N_3232,N_3120,N_3159);
and U3233 (N_3233,N_3044,N_3047);
or U3234 (N_3234,N_3088,N_3025);
or U3235 (N_3235,N_3033,N_3110);
xnor U3236 (N_3236,N_3079,N_3188);
xnor U3237 (N_3237,N_3105,N_3053);
nor U3238 (N_3238,N_3152,N_3072);
or U3239 (N_3239,N_3074,N_3109);
nand U3240 (N_3240,N_3115,N_3129);
and U3241 (N_3241,N_3093,N_3189);
or U3242 (N_3242,N_3156,N_3163);
or U3243 (N_3243,N_3071,N_3007);
nand U3244 (N_3244,N_3160,N_3048);
or U3245 (N_3245,N_3134,N_3193);
nor U3246 (N_3246,N_3124,N_3010);
xor U3247 (N_3247,N_3119,N_3068);
nand U3248 (N_3248,N_3014,N_3196);
or U3249 (N_3249,N_3194,N_3063);
nor U3250 (N_3250,N_3101,N_3023);
nor U3251 (N_3251,N_3080,N_3095);
or U3252 (N_3252,N_3086,N_3107);
nor U3253 (N_3253,N_3056,N_3030);
xor U3254 (N_3254,N_3038,N_3197);
nor U3255 (N_3255,N_3153,N_3040);
or U3256 (N_3256,N_3108,N_3054);
and U3257 (N_3257,N_3167,N_3117);
and U3258 (N_3258,N_3049,N_3041);
or U3259 (N_3259,N_3158,N_3019);
nand U3260 (N_3260,N_3103,N_3008);
or U3261 (N_3261,N_3123,N_3043);
nand U3262 (N_3262,N_3122,N_3067);
or U3263 (N_3263,N_3184,N_3114);
or U3264 (N_3264,N_3066,N_3027);
xnor U3265 (N_3265,N_3069,N_3173);
nand U3266 (N_3266,N_3164,N_3052);
and U3267 (N_3267,N_3000,N_3055);
or U3268 (N_3268,N_3098,N_3180);
and U3269 (N_3269,N_3170,N_3192);
nand U3270 (N_3270,N_3064,N_3012);
nand U3271 (N_3271,N_3081,N_3190);
nor U3272 (N_3272,N_3006,N_3076);
nand U3273 (N_3273,N_3028,N_3177);
xnor U3274 (N_3274,N_3112,N_3100);
xnor U3275 (N_3275,N_3060,N_3148);
xnor U3276 (N_3276,N_3029,N_3157);
and U3277 (N_3277,N_3187,N_3022);
or U3278 (N_3278,N_3090,N_3021);
or U3279 (N_3279,N_3045,N_3034);
and U3280 (N_3280,N_3017,N_3035);
and U3281 (N_3281,N_3143,N_3092);
and U3282 (N_3282,N_3070,N_3050);
xnor U3283 (N_3283,N_3015,N_3073);
and U3284 (N_3284,N_3155,N_3005);
nand U3285 (N_3285,N_3026,N_3144);
nand U3286 (N_3286,N_3198,N_3183);
nor U3287 (N_3287,N_3171,N_3162);
and U3288 (N_3288,N_3179,N_3172);
nor U3289 (N_3289,N_3166,N_3116);
or U3290 (N_3290,N_3099,N_3146);
nor U3291 (N_3291,N_3113,N_3036);
or U3292 (N_3292,N_3141,N_3102);
nor U3293 (N_3293,N_3169,N_3020);
nand U3294 (N_3294,N_3051,N_3058);
nor U3295 (N_3295,N_3046,N_3075);
xnor U3296 (N_3296,N_3185,N_3149);
nand U3297 (N_3297,N_3174,N_3126);
or U3298 (N_3298,N_3130,N_3004);
xor U3299 (N_3299,N_3186,N_3176);
nand U3300 (N_3300,N_3136,N_3189);
and U3301 (N_3301,N_3165,N_3031);
nor U3302 (N_3302,N_3102,N_3122);
nand U3303 (N_3303,N_3132,N_3094);
nand U3304 (N_3304,N_3181,N_3163);
or U3305 (N_3305,N_3049,N_3056);
nand U3306 (N_3306,N_3098,N_3119);
or U3307 (N_3307,N_3155,N_3061);
or U3308 (N_3308,N_3001,N_3151);
nor U3309 (N_3309,N_3041,N_3088);
nor U3310 (N_3310,N_3091,N_3080);
xnor U3311 (N_3311,N_3187,N_3091);
nand U3312 (N_3312,N_3061,N_3001);
and U3313 (N_3313,N_3137,N_3162);
or U3314 (N_3314,N_3107,N_3154);
or U3315 (N_3315,N_3046,N_3107);
or U3316 (N_3316,N_3131,N_3120);
nor U3317 (N_3317,N_3024,N_3018);
or U3318 (N_3318,N_3076,N_3025);
or U3319 (N_3319,N_3124,N_3073);
xnor U3320 (N_3320,N_3098,N_3054);
nand U3321 (N_3321,N_3198,N_3031);
nor U3322 (N_3322,N_3111,N_3145);
xor U3323 (N_3323,N_3091,N_3070);
nor U3324 (N_3324,N_3055,N_3178);
and U3325 (N_3325,N_3163,N_3137);
nand U3326 (N_3326,N_3174,N_3019);
or U3327 (N_3327,N_3191,N_3014);
or U3328 (N_3328,N_3188,N_3076);
xnor U3329 (N_3329,N_3112,N_3114);
and U3330 (N_3330,N_3162,N_3131);
nor U3331 (N_3331,N_3122,N_3149);
xor U3332 (N_3332,N_3196,N_3029);
nor U3333 (N_3333,N_3051,N_3001);
or U3334 (N_3334,N_3055,N_3015);
or U3335 (N_3335,N_3190,N_3022);
or U3336 (N_3336,N_3171,N_3109);
and U3337 (N_3337,N_3155,N_3062);
xor U3338 (N_3338,N_3073,N_3007);
or U3339 (N_3339,N_3182,N_3075);
nand U3340 (N_3340,N_3148,N_3012);
and U3341 (N_3341,N_3020,N_3172);
and U3342 (N_3342,N_3010,N_3023);
nand U3343 (N_3343,N_3062,N_3163);
nand U3344 (N_3344,N_3197,N_3071);
nand U3345 (N_3345,N_3116,N_3081);
nand U3346 (N_3346,N_3105,N_3144);
or U3347 (N_3347,N_3056,N_3000);
xnor U3348 (N_3348,N_3115,N_3172);
nand U3349 (N_3349,N_3162,N_3064);
nand U3350 (N_3350,N_3031,N_3108);
nor U3351 (N_3351,N_3079,N_3126);
xor U3352 (N_3352,N_3119,N_3138);
xnor U3353 (N_3353,N_3176,N_3184);
nor U3354 (N_3354,N_3180,N_3075);
or U3355 (N_3355,N_3058,N_3017);
nor U3356 (N_3356,N_3034,N_3003);
nand U3357 (N_3357,N_3149,N_3012);
nor U3358 (N_3358,N_3160,N_3148);
nand U3359 (N_3359,N_3048,N_3043);
and U3360 (N_3360,N_3012,N_3005);
nor U3361 (N_3361,N_3064,N_3172);
nand U3362 (N_3362,N_3181,N_3137);
and U3363 (N_3363,N_3183,N_3087);
nor U3364 (N_3364,N_3103,N_3186);
nand U3365 (N_3365,N_3028,N_3093);
and U3366 (N_3366,N_3069,N_3084);
and U3367 (N_3367,N_3066,N_3160);
and U3368 (N_3368,N_3007,N_3129);
or U3369 (N_3369,N_3194,N_3108);
nor U3370 (N_3370,N_3185,N_3115);
nand U3371 (N_3371,N_3030,N_3130);
or U3372 (N_3372,N_3088,N_3149);
xnor U3373 (N_3373,N_3170,N_3139);
xor U3374 (N_3374,N_3139,N_3030);
nand U3375 (N_3375,N_3103,N_3147);
nor U3376 (N_3376,N_3052,N_3168);
or U3377 (N_3377,N_3162,N_3072);
or U3378 (N_3378,N_3073,N_3131);
and U3379 (N_3379,N_3115,N_3114);
and U3380 (N_3380,N_3121,N_3074);
nand U3381 (N_3381,N_3072,N_3128);
and U3382 (N_3382,N_3150,N_3034);
nand U3383 (N_3383,N_3131,N_3009);
or U3384 (N_3384,N_3132,N_3061);
nand U3385 (N_3385,N_3109,N_3181);
and U3386 (N_3386,N_3079,N_3110);
nor U3387 (N_3387,N_3008,N_3117);
xnor U3388 (N_3388,N_3099,N_3181);
and U3389 (N_3389,N_3043,N_3177);
nor U3390 (N_3390,N_3180,N_3017);
nor U3391 (N_3391,N_3103,N_3084);
and U3392 (N_3392,N_3144,N_3130);
nand U3393 (N_3393,N_3108,N_3070);
xor U3394 (N_3394,N_3096,N_3066);
and U3395 (N_3395,N_3121,N_3131);
or U3396 (N_3396,N_3199,N_3162);
nor U3397 (N_3397,N_3078,N_3131);
nand U3398 (N_3398,N_3177,N_3174);
nor U3399 (N_3399,N_3149,N_3059);
or U3400 (N_3400,N_3315,N_3241);
nand U3401 (N_3401,N_3217,N_3294);
nor U3402 (N_3402,N_3388,N_3260);
or U3403 (N_3403,N_3349,N_3387);
xor U3404 (N_3404,N_3339,N_3347);
nand U3405 (N_3405,N_3377,N_3249);
nor U3406 (N_3406,N_3218,N_3281);
nor U3407 (N_3407,N_3308,N_3397);
and U3408 (N_3408,N_3328,N_3268);
nor U3409 (N_3409,N_3391,N_3359);
nand U3410 (N_3410,N_3220,N_3326);
nor U3411 (N_3411,N_3275,N_3364);
nor U3412 (N_3412,N_3212,N_3235);
nor U3413 (N_3413,N_3252,N_3264);
nor U3414 (N_3414,N_3353,N_3331);
nand U3415 (N_3415,N_3236,N_3225);
nor U3416 (N_3416,N_3350,N_3243);
nor U3417 (N_3417,N_3376,N_3390);
and U3418 (N_3418,N_3336,N_3367);
or U3419 (N_3419,N_3361,N_3382);
nand U3420 (N_3420,N_3302,N_3348);
or U3421 (N_3421,N_3307,N_3202);
nor U3422 (N_3422,N_3360,N_3366);
nand U3423 (N_3423,N_3355,N_3351);
nor U3424 (N_3424,N_3354,N_3276);
and U3425 (N_3425,N_3231,N_3288);
and U3426 (N_3426,N_3309,N_3259);
nor U3427 (N_3427,N_3208,N_3200);
and U3428 (N_3428,N_3311,N_3383);
xnor U3429 (N_3429,N_3250,N_3318);
nand U3430 (N_3430,N_3232,N_3293);
nand U3431 (N_3431,N_3216,N_3321);
nand U3432 (N_3432,N_3206,N_3298);
nor U3433 (N_3433,N_3320,N_3370);
and U3434 (N_3434,N_3254,N_3297);
and U3435 (N_3435,N_3256,N_3392);
nor U3436 (N_3436,N_3386,N_3356);
nor U3437 (N_3437,N_3301,N_3229);
or U3438 (N_3438,N_3272,N_3322);
or U3439 (N_3439,N_3385,N_3224);
and U3440 (N_3440,N_3292,N_3396);
nand U3441 (N_3441,N_3372,N_3389);
and U3442 (N_3442,N_3300,N_3346);
nand U3443 (N_3443,N_3201,N_3312);
and U3444 (N_3444,N_3246,N_3344);
or U3445 (N_3445,N_3271,N_3324);
and U3446 (N_3446,N_3219,N_3325);
or U3447 (N_3447,N_3266,N_3261);
nor U3448 (N_3448,N_3340,N_3253);
or U3449 (N_3449,N_3362,N_3365);
nand U3450 (N_3450,N_3369,N_3393);
or U3451 (N_3451,N_3335,N_3299);
and U3452 (N_3452,N_3226,N_3273);
or U3453 (N_3453,N_3251,N_3379);
nor U3454 (N_3454,N_3265,N_3207);
and U3455 (N_3455,N_3228,N_3262);
nand U3456 (N_3456,N_3214,N_3374);
nor U3457 (N_3457,N_3398,N_3305);
xor U3458 (N_3458,N_3221,N_3303);
nor U3459 (N_3459,N_3248,N_3310);
xnor U3460 (N_3460,N_3373,N_3210);
nor U3461 (N_3461,N_3289,N_3240);
xnor U3462 (N_3462,N_3375,N_3378);
and U3463 (N_3463,N_3357,N_3255);
or U3464 (N_3464,N_3381,N_3269);
nor U3465 (N_3465,N_3368,N_3209);
nand U3466 (N_3466,N_3280,N_3285);
nor U3467 (N_3467,N_3314,N_3291);
nor U3468 (N_3468,N_3317,N_3287);
nor U3469 (N_3469,N_3279,N_3230);
and U3470 (N_3470,N_3239,N_3334);
and U3471 (N_3471,N_3258,N_3204);
xnor U3472 (N_3472,N_3304,N_3277);
nand U3473 (N_3473,N_3227,N_3233);
xnor U3474 (N_3474,N_3327,N_3284);
xor U3475 (N_3475,N_3319,N_3384);
or U3476 (N_3476,N_3215,N_3283);
and U3477 (N_3477,N_3203,N_3296);
nand U3478 (N_3478,N_3330,N_3323);
xnor U3479 (N_3479,N_3342,N_3274);
or U3480 (N_3480,N_3278,N_3205);
nand U3481 (N_3481,N_3395,N_3267);
nand U3482 (N_3482,N_3247,N_3345);
or U3483 (N_3483,N_3341,N_3313);
nand U3484 (N_3484,N_3316,N_3222);
nand U3485 (N_3485,N_3329,N_3332);
and U3486 (N_3486,N_3263,N_3306);
and U3487 (N_3487,N_3363,N_3290);
or U3488 (N_3488,N_3237,N_3394);
nor U3489 (N_3489,N_3286,N_3343);
and U3490 (N_3490,N_3380,N_3257);
nand U3491 (N_3491,N_3245,N_3213);
or U3492 (N_3492,N_3282,N_3223);
xor U3493 (N_3493,N_3238,N_3211);
nand U3494 (N_3494,N_3242,N_3337);
and U3495 (N_3495,N_3333,N_3371);
xnor U3496 (N_3496,N_3234,N_3358);
nor U3497 (N_3497,N_3399,N_3270);
and U3498 (N_3498,N_3244,N_3352);
and U3499 (N_3499,N_3295,N_3338);
xor U3500 (N_3500,N_3329,N_3226);
nand U3501 (N_3501,N_3252,N_3385);
and U3502 (N_3502,N_3298,N_3343);
nand U3503 (N_3503,N_3273,N_3250);
or U3504 (N_3504,N_3287,N_3206);
nor U3505 (N_3505,N_3205,N_3353);
nand U3506 (N_3506,N_3331,N_3365);
and U3507 (N_3507,N_3259,N_3228);
nor U3508 (N_3508,N_3332,N_3361);
xor U3509 (N_3509,N_3398,N_3392);
nand U3510 (N_3510,N_3319,N_3209);
nand U3511 (N_3511,N_3295,N_3373);
and U3512 (N_3512,N_3332,N_3304);
nor U3513 (N_3513,N_3327,N_3342);
or U3514 (N_3514,N_3364,N_3339);
xnor U3515 (N_3515,N_3342,N_3271);
or U3516 (N_3516,N_3232,N_3361);
or U3517 (N_3517,N_3243,N_3208);
nand U3518 (N_3518,N_3310,N_3318);
or U3519 (N_3519,N_3225,N_3399);
and U3520 (N_3520,N_3297,N_3226);
nor U3521 (N_3521,N_3249,N_3297);
nor U3522 (N_3522,N_3382,N_3265);
nor U3523 (N_3523,N_3345,N_3333);
and U3524 (N_3524,N_3261,N_3326);
nand U3525 (N_3525,N_3393,N_3303);
nor U3526 (N_3526,N_3307,N_3399);
nor U3527 (N_3527,N_3340,N_3317);
nor U3528 (N_3528,N_3296,N_3201);
or U3529 (N_3529,N_3379,N_3325);
nor U3530 (N_3530,N_3202,N_3240);
and U3531 (N_3531,N_3355,N_3343);
or U3532 (N_3532,N_3397,N_3331);
or U3533 (N_3533,N_3386,N_3318);
and U3534 (N_3534,N_3301,N_3340);
or U3535 (N_3535,N_3255,N_3265);
or U3536 (N_3536,N_3376,N_3300);
xnor U3537 (N_3537,N_3299,N_3243);
or U3538 (N_3538,N_3230,N_3371);
and U3539 (N_3539,N_3339,N_3359);
or U3540 (N_3540,N_3283,N_3233);
nor U3541 (N_3541,N_3356,N_3310);
nand U3542 (N_3542,N_3225,N_3226);
or U3543 (N_3543,N_3388,N_3365);
nor U3544 (N_3544,N_3360,N_3319);
or U3545 (N_3545,N_3342,N_3261);
or U3546 (N_3546,N_3323,N_3393);
nand U3547 (N_3547,N_3207,N_3335);
or U3548 (N_3548,N_3293,N_3231);
and U3549 (N_3549,N_3385,N_3312);
or U3550 (N_3550,N_3227,N_3220);
nand U3551 (N_3551,N_3236,N_3369);
nand U3552 (N_3552,N_3204,N_3354);
and U3553 (N_3553,N_3236,N_3239);
nand U3554 (N_3554,N_3311,N_3297);
and U3555 (N_3555,N_3271,N_3321);
or U3556 (N_3556,N_3274,N_3306);
xor U3557 (N_3557,N_3371,N_3332);
nor U3558 (N_3558,N_3249,N_3363);
xor U3559 (N_3559,N_3290,N_3206);
xor U3560 (N_3560,N_3232,N_3210);
and U3561 (N_3561,N_3371,N_3334);
nor U3562 (N_3562,N_3228,N_3236);
or U3563 (N_3563,N_3369,N_3259);
or U3564 (N_3564,N_3237,N_3330);
or U3565 (N_3565,N_3392,N_3224);
nor U3566 (N_3566,N_3232,N_3276);
and U3567 (N_3567,N_3268,N_3278);
nand U3568 (N_3568,N_3323,N_3265);
nand U3569 (N_3569,N_3336,N_3211);
or U3570 (N_3570,N_3343,N_3288);
nand U3571 (N_3571,N_3216,N_3255);
nor U3572 (N_3572,N_3382,N_3381);
xnor U3573 (N_3573,N_3397,N_3345);
and U3574 (N_3574,N_3212,N_3255);
nor U3575 (N_3575,N_3255,N_3267);
nor U3576 (N_3576,N_3314,N_3270);
and U3577 (N_3577,N_3370,N_3222);
or U3578 (N_3578,N_3223,N_3227);
or U3579 (N_3579,N_3378,N_3226);
nor U3580 (N_3580,N_3293,N_3373);
and U3581 (N_3581,N_3367,N_3362);
or U3582 (N_3582,N_3319,N_3271);
or U3583 (N_3583,N_3314,N_3364);
nand U3584 (N_3584,N_3266,N_3334);
and U3585 (N_3585,N_3285,N_3297);
or U3586 (N_3586,N_3328,N_3264);
nand U3587 (N_3587,N_3398,N_3382);
and U3588 (N_3588,N_3370,N_3205);
xor U3589 (N_3589,N_3326,N_3312);
and U3590 (N_3590,N_3330,N_3316);
or U3591 (N_3591,N_3330,N_3291);
nand U3592 (N_3592,N_3315,N_3295);
and U3593 (N_3593,N_3366,N_3268);
or U3594 (N_3594,N_3365,N_3200);
or U3595 (N_3595,N_3398,N_3224);
xor U3596 (N_3596,N_3304,N_3280);
nand U3597 (N_3597,N_3275,N_3384);
nor U3598 (N_3598,N_3300,N_3290);
xnor U3599 (N_3599,N_3324,N_3299);
and U3600 (N_3600,N_3578,N_3432);
and U3601 (N_3601,N_3473,N_3453);
nor U3602 (N_3602,N_3497,N_3598);
xnor U3603 (N_3603,N_3400,N_3590);
and U3604 (N_3604,N_3591,N_3466);
and U3605 (N_3605,N_3520,N_3586);
and U3606 (N_3606,N_3447,N_3494);
and U3607 (N_3607,N_3407,N_3575);
or U3608 (N_3608,N_3484,N_3426);
and U3609 (N_3609,N_3583,N_3588);
nor U3610 (N_3610,N_3440,N_3577);
and U3611 (N_3611,N_3524,N_3418);
xor U3612 (N_3612,N_3541,N_3468);
nand U3613 (N_3613,N_3576,N_3507);
xor U3614 (N_3614,N_3498,N_3510);
and U3615 (N_3615,N_3414,N_3443);
or U3616 (N_3616,N_3557,N_3559);
and U3617 (N_3617,N_3436,N_3412);
xnor U3618 (N_3618,N_3450,N_3491);
and U3619 (N_3619,N_3485,N_3552);
nand U3620 (N_3620,N_3431,N_3425);
or U3621 (N_3621,N_3406,N_3455);
nand U3622 (N_3622,N_3549,N_3486);
and U3623 (N_3623,N_3509,N_3584);
or U3624 (N_3624,N_3517,N_3579);
nor U3625 (N_3625,N_3596,N_3462);
or U3626 (N_3626,N_3595,N_3580);
nand U3627 (N_3627,N_3533,N_3481);
or U3628 (N_3628,N_3402,N_3401);
and U3629 (N_3629,N_3461,N_3449);
nor U3630 (N_3630,N_3553,N_3448);
and U3631 (N_3631,N_3573,N_3538);
xor U3632 (N_3632,N_3519,N_3506);
and U3633 (N_3633,N_3558,N_3493);
nand U3634 (N_3634,N_3526,N_3437);
nor U3635 (N_3635,N_3545,N_3454);
or U3636 (N_3636,N_3404,N_3536);
nand U3637 (N_3637,N_3562,N_3566);
nand U3638 (N_3638,N_3532,N_3565);
or U3639 (N_3639,N_3471,N_3599);
or U3640 (N_3640,N_3521,N_3516);
and U3641 (N_3641,N_3459,N_3419);
and U3642 (N_3642,N_3410,N_3585);
nor U3643 (N_3643,N_3503,N_3403);
nor U3644 (N_3644,N_3515,N_3489);
xnor U3645 (N_3645,N_3405,N_3424);
or U3646 (N_3646,N_3499,N_3492);
nor U3647 (N_3647,N_3512,N_3423);
and U3648 (N_3648,N_3550,N_3518);
nor U3649 (N_3649,N_3445,N_3587);
or U3650 (N_3650,N_3531,N_3514);
nand U3651 (N_3651,N_3444,N_3456);
nand U3652 (N_3652,N_3582,N_3475);
nand U3653 (N_3653,N_3597,N_3513);
nor U3654 (N_3654,N_3535,N_3434);
xnor U3655 (N_3655,N_3415,N_3567);
nor U3656 (N_3656,N_3523,N_3551);
nor U3657 (N_3657,N_3546,N_3487);
and U3658 (N_3658,N_3477,N_3539);
xnor U3659 (N_3659,N_3500,N_3408);
nor U3660 (N_3660,N_3483,N_3564);
nor U3661 (N_3661,N_3467,N_3409);
and U3662 (N_3662,N_3505,N_3522);
xnor U3663 (N_3663,N_3476,N_3469);
nand U3664 (N_3664,N_3496,N_3490);
or U3665 (N_3665,N_3581,N_3528);
nor U3666 (N_3666,N_3480,N_3508);
nor U3667 (N_3667,N_3435,N_3488);
nand U3668 (N_3668,N_3460,N_3416);
or U3669 (N_3669,N_3421,N_3548);
nor U3670 (N_3670,N_3482,N_3571);
nor U3671 (N_3671,N_3547,N_3530);
nor U3672 (N_3672,N_3511,N_3427);
nand U3673 (N_3673,N_3527,N_3504);
and U3674 (N_3674,N_3411,N_3441);
nand U3675 (N_3675,N_3478,N_3569);
or U3676 (N_3676,N_3593,N_3555);
or U3677 (N_3677,N_3442,N_3572);
xnor U3678 (N_3678,N_3568,N_3429);
nor U3679 (N_3679,N_3417,N_3479);
and U3680 (N_3680,N_3457,N_3433);
nor U3681 (N_3681,N_3534,N_3592);
nand U3682 (N_3682,N_3464,N_3563);
and U3683 (N_3683,N_3560,N_3474);
nand U3684 (N_3684,N_3574,N_3420);
nand U3685 (N_3685,N_3501,N_3544);
and U3686 (N_3686,N_3525,N_3465);
and U3687 (N_3687,N_3470,N_3451);
nand U3688 (N_3688,N_3542,N_3589);
and U3689 (N_3689,N_3452,N_3543);
or U3690 (N_3690,N_3561,N_3554);
xor U3691 (N_3691,N_3413,N_3537);
or U3692 (N_3692,N_3529,N_3422);
or U3693 (N_3693,N_3438,N_3439);
xor U3694 (N_3694,N_3430,N_3472);
or U3695 (N_3695,N_3428,N_3502);
nor U3696 (N_3696,N_3540,N_3570);
nor U3697 (N_3697,N_3556,N_3446);
and U3698 (N_3698,N_3594,N_3458);
nand U3699 (N_3699,N_3463,N_3495);
or U3700 (N_3700,N_3469,N_3583);
nor U3701 (N_3701,N_3508,N_3597);
nand U3702 (N_3702,N_3420,N_3475);
or U3703 (N_3703,N_3456,N_3446);
or U3704 (N_3704,N_3588,N_3599);
or U3705 (N_3705,N_3504,N_3581);
nand U3706 (N_3706,N_3576,N_3580);
nor U3707 (N_3707,N_3589,N_3534);
nand U3708 (N_3708,N_3444,N_3408);
and U3709 (N_3709,N_3444,N_3448);
or U3710 (N_3710,N_3573,N_3409);
nand U3711 (N_3711,N_3489,N_3426);
and U3712 (N_3712,N_3464,N_3421);
or U3713 (N_3713,N_3591,N_3483);
or U3714 (N_3714,N_3592,N_3501);
or U3715 (N_3715,N_3423,N_3463);
nor U3716 (N_3716,N_3407,N_3431);
nand U3717 (N_3717,N_3522,N_3404);
nor U3718 (N_3718,N_3417,N_3586);
nor U3719 (N_3719,N_3595,N_3597);
and U3720 (N_3720,N_3430,N_3414);
or U3721 (N_3721,N_3404,N_3434);
xnor U3722 (N_3722,N_3589,N_3485);
nand U3723 (N_3723,N_3474,N_3461);
nand U3724 (N_3724,N_3549,N_3491);
or U3725 (N_3725,N_3510,N_3446);
and U3726 (N_3726,N_3598,N_3531);
xnor U3727 (N_3727,N_3552,N_3409);
nor U3728 (N_3728,N_3546,N_3441);
or U3729 (N_3729,N_3511,N_3451);
and U3730 (N_3730,N_3548,N_3531);
nand U3731 (N_3731,N_3582,N_3565);
nor U3732 (N_3732,N_3407,N_3552);
nor U3733 (N_3733,N_3537,N_3584);
and U3734 (N_3734,N_3483,N_3535);
and U3735 (N_3735,N_3458,N_3478);
nor U3736 (N_3736,N_3559,N_3465);
nor U3737 (N_3737,N_3484,N_3544);
xnor U3738 (N_3738,N_3495,N_3499);
or U3739 (N_3739,N_3517,N_3576);
nand U3740 (N_3740,N_3516,N_3439);
and U3741 (N_3741,N_3420,N_3528);
nand U3742 (N_3742,N_3472,N_3572);
nor U3743 (N_3743,N_3532,N_3403);
nand U3744 (N_3744,N_3536,N_3531);
nor U3745 (N_3745,N_3537,N_3477);
nor U3746 (N_3746,N_3412,N_3484);
or U3747 (N_3747,N_3518,N_3416);
or U3748 (N_3748,N_3571,N_3535);
and U3749 (N_3749,N_3482,N_3546);
xor U3750 (N_3750,N_3436,N_3454);
or U3751 (N_3751,N_3594,N_3491);
or U3752 (N_3752,N_3434,N_3580);
nor U3753 (N_3753,N_3416,N_3444);
or U3754 (N_3754,N_3483,N_3456);
nand U3755 (N_3755,N_3452,N_3537);
nand U3756 (N_3756,N_3552,N_3410);
or U3757 (N_3757,N_3492,N_3572);
nand U3758 (N_3758,N_3543,N_3562);
and U3759 (N_3759,N_3560,N_3552);
xor U3760 (N_3760,N_3408,N_3460);
or U3761 (N_3761,N_3525,N_3547);
or U3762 (N_3762,N_3400,N_3536);
xnor U3763 (N_3763,N_3531,N_3560);
xor U3764 (N_3764,N_3419,N_3444);
nor U3765 (N_3765,N_3511,N_3466);
nor U3766 (N_3766,N_3471,N_3587);
or U3767 (N_3767,N_3413,N_3504);
nor U3768 (N_3768,N_3460,N_3566);
or U3769 (N_3769,N_3410,N_3497);
or U3770 (N_3770,N_3537,N_3478);
and U3771 (N_3771,N_3595,N_3438);
and U3772 (N_3772,N_3594,N_3420);
nand U3773 (N_3773,N_3450,N_3465);
and U3774 (N_3774,N_3469,N_3482);
nor U3775 (N_3775,N_3587,N_3575);
nand U3776 (N_3776,N_3406,N_3536);
or U3777 (N_3777,N_3436,N_3418);
nor U3778 (N_3778,N_3500,N_3444);
and U3779 (N_3779,N_3536,N_3402);
nand U3780 (N_3780,N_3580,N_3538);
and U3781 (N_3781,N_3579,N_3401);
nand U3782 (N_3782,N_3429,N_3422);
and U3783 (N_3783,N_3590,N_3562);
or U3784 (N_3784,N_3513,N_3553);
xnor U3785 (N_3785,N_3441,N_3467);
and U3786 (N_3786,N_3547,N_3479);
nand U3787 (N_3787,N_3515,N_3408);
nor U3788 (N_3788,N_3454,N_3418);
or U3789 (N_3789,N_3536,N_3550);
nand U3790 (N_3790,N_3559,N_3433);
nor U3791 (N_3791,N_3522,N_3533);
nor U3792 (N_3792,N_3576,N_3515);
nand U3793 (N_3793,N_3566,N_3497);
and U3794 (N_3794,N_3589,N_3422);
and U3795 (N_3795,N_3488,N_3466);
or U3796 (N_3796,N_3540,N_3449);
nor U3797 (N_3797,N_3555,N_3594);
or U3798 (N_3798,N_3484,N_3454);
or U3799 (N_3799,N_3580,N_3534);
nand U3800 (N_3800,N_3779,N_3791);
and U3801 (N_3801,N_3718,N_3630);
nor U3802 (N_3802,N_3629,N_3798);
nor U3803 (N_3803,N_3708,N_3673);
nor U3804 (N_3804,N_3626,N_3763);
and U3805 (N_3805,N_3764,N_3665);
and U3806 (N_3806,N_3744,N_3715);
xor U3807 (N_3807,N_3747,N_3741);
nor U3808 (N_3808,N_3736,N_3622);
or U3809 (N_3809,N_3730,N_3647);
or U3810 (N_3810,N_3676,N_3769);
or U3811 (N_3811,N_3648,N_3654);
nor U3812 (N_3812,N_3696,N_3606);
nand U3813 (N_3813,N_3687,N_3616);
nor U3814 (N_3814,N_3615,N_3771);
nand U3815 (N_3815,N_3794,N_3627);
and U3816 (N_3816,N_3625,N_3731);
and U3817 (N_3817,N_3603,N_3787);
nand U3818 (N_3818,N_3772,N_3675);
xor U3819 (N_3819,N_3702,N_3619);
nand U3820 (N_3820,N_3790,N_3651);
or U3821 (N_3821,N_3748,N_3700);
and U3822 (N_3822,N_3768,N_3780);
or U3823 (N_3823,N_3792,N_3656);
nor U3824 (N_3824,N_3664,N_3678);
xor U3825 (N_3825,N_3767,N_3608);
or U3826 (N_3826,N_3649,N_3727);
or U3827 (N_3827,N_3693,N_3770);
or U3828 (N_3828,N_3706,N_3778);
nand U3829 (N_3829,N_3752,N_3728);
and U3830 (N_3830,N_3663,N_3640);
nand U3831 (N_3831,N_3668,N_3757);
and U3832 (N_3832,N_3638,N_3698);
nor U3833 (N_3833,N_3683,N_3762);
and U3834 (N_3834,N_3636,N_3697);
and U3835 (N_3835,N_3682,N_3776);
nand U3836 (N_3836,N_3699,N_3754);
nor U3837 (N_3837,N_3703,N_3775);
nor U3838 (N_3838,N_3756,N_3604);
nor U3839 (N_3839,N_3707,N_3637);
and U3840 (N_3840,N_3639,N_3758);
xnor U3841 (N_3841,N_3788,N_3691);
or U3842 (N_3842,N_3607,N_3735);
nand U3843 (N_3843,N_3661,N_3609);
or U3844 (N_3844,N_3620,N_3795);
or U3845 (N_3845,N_3652,N_3712);
or U3846 (N_3846,N_3797,N_3746);
and U3847 (N_3847,N_3760,N_3759);
or U3848 (N_3848,N_3695,N_3633);
or U3849 (N_3849,N_3704,N_3737);
nand U3850 (N_3850,N_3650,N_3782);
and U3851 (N_3851,N_3786,N_3688);
and U3852 (N_3852,N_3705,N_3789);
xnor U3853 (N_3853,N_3716,N_3624);
nand U3854 (N_3854,N_3643,N_3799);
nand U3855 (N_3855,N_3618,N_3709);
nand U3856 (N_3856,N_3723,N_3796);
nand U3857 (N_3857,N_3632,N_3749);
nor U3858 (N_3858,N_3773,N_3738);
or U3859 (N_3859,N_3739,N_3681);
xor U3860 (N_3860,N_3662,N_3742);
or U3861 (N_3861,N_3729,N_3672);
or U3862 (N_3862,N_3670,N_3677);
nor U3863 (N_3863,N_3635,N_3646);
xor U3864 (N_3864,N_3641,N_3755);
or U3865 (N_3865,N_3600,N_3653);
or U3866 (N_3866,N_3602,N_3684);
or U3867 (N_3867,N_3623,N_3774);
nor U3868 (N_3868,N_3711,N_3644);
or U3869 (N_3869,N_3701,N_3692);
or U3870 (N_3870,N_3617,N_3628);
or U3871 (N_3871,N_3719,N_3621);
or U3872 (N_3872,N_3753,N_3751);
nor U3873 (N_3873,N_3721,N_3613);
and U3874 (N_3874,N_3750,N_3690);
xor U3875 (N_3875,N_3713,N_3732);
and U3876 (N_3876,N_3726,N_3686);
nand U3877 (N_3877,N_3605,N_3714);
and U3878 (N_3878,N_3669,N_3667);
xnor U3879 (N_3879,N_3717,N_3733);
or U3880 (N_3880,N_3743,N_3745);
nor U3881 (N_3881,N_3761,N_3785);
and U3882 (N_3882,N_3612,N_3658);
and U3883 (N_3883,N_3784,N_3642);
nand U3884 (N_3884,N_3645,N_3694);
and U3885 (N_3885,N_3655,N_3793);
or U3886 (N_3886,N_3614,N_3765);
or U3887 (N_3887,N_3657,N_3631);
nor U3888 (N_3888,N_3634,N_3679);
or U3889 (N_3889,N_3680,N_3766);
nor U3890 (N_3890,N_3611,N_3666);
or U3891 (N_3891,N_3710,N_3610);
nand U3892 (N_3892,N_3671,N_3777);
nor U3893 (N_3893,N_3674,N_3724);
and U3894 (N_3894,N_3659,N_3740);
and U3895 (N_3895,N_3685,N_3725);
or U3896 (N_3896,N_3660,N_3601);
nand U3897 (N_3897,N_3781,N_3734);
and U3898 (N_3898,N_3722,N_3689);
nor U3899 (N_3899,N_3783,N_3720);
nand U3900 (N_3900,N_3607,N_3740);
and U3901 (N_3901,N_3619,N_3689);
nand U3902 (N_3902,N_3667,N_3640);
and U3903 (N_3903,N_3784,N_3630);
or U3904 (N_3904,N_3693,N_3769);
and U3905 (N_3905,N_3721,N_3797);
nor U3906 (N_3906,N_3657,N_3620);
nor U3907 (N_3907,N_3736,N_3611);
or U3908 (N_3908,N_3778,N_3788);
and U3909 (N_3909,N_3624,N_3708);
xor U3910 (N_3910,N_3637,N_3686);
nand U3911 (N_3911,N_3755,N_3749);
or U3912 (N_3912,N_3688,N_3719);
and U3913 (N_3913,N_3673,N_3680);
and U3914 (N_3914,N_3779,N_3689);
xor U3915 (N_3915,N_3765,N_3746);
nand U3916 (N_3916,N_3624,N_3637);
or U3917 (N_3917,N_3774,N_3758);
nor U3918 (N_3918,N_3638,N_3785);
nor U3919 (N_3919,N_3662,N_3741);
or U3920 (N_3920,N_3728,N_3614);
nor U3921 (N_3921,N_3647,N_3732);
nand U3922 (N_3922,N_3667,N_3796);
and U3923 (N_3923,N_3717,N_3660);
or U3924 (N_3924,N_3663,N_3774);
and U3925 (N_3925,N_3734,N_3728);
nor U3926 (N_3926,N_3734,N_3621);
and U3927 (N_3927,N_3608,N_3779);
nor U3928 (N_3928,N_3698,N_3623);
nand U3929 (N_3929,N_3756,N_3746);
or U3930 (N_3930,N_3715,N_3647);
and U3931 (N_3931,N_3744,N_3636);
nor U3932 (N_3932,N_3749,N_3691);
or U3933 (N_3933,N_3654,N_3792);
or U3934 (N_3934,N_3680,N_3783);
and U3935 (N_3935,N_3763,N_3721);
nand U3936 (N_3936,N_3696,N_3799);
or U3937 (N_3937,N_3748,N_3677);
nand U3938 (N_3938,N_3792,N_3644);
xnor U3939 (N_3939,N_3650,N_3676);
nand U3940 (N_3940,N_3797,N_3634);
or U3941 (N_3941,N_3737,N_3701);
or U3942 (N_3942,N_3668,N_3686);
and U3943 (N_3943,N_3727,N_3617);
and U3944 (N_3944,N_3743,N_3739);
or U3945 (N_3945,N_3676,N_3723);
or U3946 (N_3946,N_3624,N_3731);
nand U3947 (N_3947,N_3749,N_3722);
nor U3948 (N_3948,N_3696,N_3722);
nor U3949 (N_3949,N_3732,N_3680);
and U3950 (N_3950,N_3679,N_3749);
nor U3951 (N_3951,N_3695,N_3731);
xnor U3952 (N_3952,N_3719,N_3705);
and U3953 (N_3953,N_3685,N_3759);
nor U3954 (N_3954,N_3608,N_3759);
xor U3955 (N_3955,N_3736,N_3700);
and U3956 (N_3956,N_3617,N_3717);
nand U3957 (N_3957,N_3737,N_3637);
and U3958 (N_3958,N_3629,N_3729);
and U3959 (N_3959,N_3660,N_3625);
and U3960 (N_3960,N_3708,N_3721);
nand U3961 (N_3961,N_3710,N_3795);
and U3962 (N_3962,N_3746,N_3770);
xor U3963 (N_3963,N_3676,N_3707);
nand U3964 (N_3964,N_3709,N_3791);
nor U3965 (N_3965,N_3642,N_3754);
nor U3966 (N_3966,N_3733,N_3775);
or U3967 (N_3967,N_3713,N_3720);
and U3968 (N_3968,N_3719,N_3741);
nor U3969 (N_3969,N_3732,N_3746);
or U3970 (N_3970,N_3649,N_3604);
xor U3971 (N_3971,N_3781,N_3796);
and U3972 (N_3972,N_3686,N_3718);
or U3973 (N_3973,N_3658,N_3603);
or U3974 (N_3974,N_3676,N_3633);
nand U3975 (N_3975,N_3692,N_3608);
nand U3976 (N_3976,N_3673,N_3701);
nand U3977 (N_3977,N_3798,N_3730);
and U3978 (N_3978,N_3659,N_3601);
and U3979 (N_3979,N_3607,N_3691);
nand U3980 (N_3980,N_3630,N_3625);
and U3981 (N_3981,N_3766,N_3650);
and U3982 (N_3982,N_3737,N_3781);
and U3983 (N_3983,N_3676,N_3610);
nand U3984 (N_3984,N_3791,N_3790);
or U3985 (N_3985,N_3633,N_3613);
nand U3986 (N_3986,N_3627,N_3770);
nor U3987 (N_3987,N_3660,N_3772);
or U3988 (N_3988,N_3769,N_3712);
and U3989 (N_3989,N_3799,N_3637);
nor U3990 (N_3990,N_3721,N_3633);
nand U3991 (N_3991,N_3737,N_3612);
or U3992 (N_3992,N_3753,N_3634);
or U3993 (N_3993,N_3678,N_3714);
nand U3994 (N_3994,N_3798,N_3645);
nor U3995 (N_3995,N_3706,N_3746);
nor U3996 (N_3996,N_3659,N_3749);
nand U3997 (N_3997,N_3710,N_3633);
nor U3998 (N_3998,N_3649,N_3722);
nor U3999 (N_3999,N_3778,N_3678);
nand U4000 (N_4000,N_3945,N_3900);
or U4001 (N_4001,N_3952,N_3891);
nand U4002 (N_4002,N_3926,N_3964);
or U4003 (N_4003,N_3943,N_3903);
nor U4004 (N_4004,N_3857,N_3941);
or U4005 (N_4005,N_3961,N_3863);
nand U4006 (N_4006,N_3873,N_3874);
and U4007 (N_4007,N_3962,N_3985);
nor U4008 (N_4008,N_3879,N_3892);
or U4009 (N_4009,N_3995,N_3957);
nor U4010 (N_4010,N_3906,N_3856);
nor U4011 (N_4011,N_3912,N_3841);
nor U4012 (N_4012,N_3940,N_3904);
xnor U4013 (N_4013,N_3963,N_3970);
nor U4014 (N_4014,N_3993,N_3846);
and U4015 (N_4015,N_3854,N_3902);
or U4016 (N_4016,N_3808,N_3858);
or U4017 (N_4017,N_3920,N_3837);
nor U4018 (N_4018,N_3918,N_3948);
nand U4019 (N_4019,N_3882,N_3988);
nor U4020 (N_4020,N_3833,N_3937);
and U4021 (N_4021,N_3984,N_3840);
nand U4022 (N_4022,N_3991,N_3996);
nand U4023 (N_4023,N_3800,N_3867);
xnor U4024 (N_4024,N_3978,N_3847);
nand U4025 (N_4025,N_3927,N_3834);
xnor U4026 (N_4026,N_3934,N_3917);
nor U4027 (N_4027,N_3850,N_3887);
nor U4028 (N_4028,N_3866,N_3851);
nor U4029 (N_4029,N_3896,N_3935);
or U4030 (N_4030,N_3827,N_3944);
nor U4031 (N_4031,N_3813,N_3969);
nor U4032 (N_4032,N_3960,N_3807);
and U4033 (N_4033,N_3845,N_3815);
or U4034 (N_4034,N_3801,N_3843);
and U4035 (N_4035,N_3973,N_3809);
nor U4036 (N_4036,N_3872,N_3930);
and U4037 (N_4037,N_3822,N_3823);
nor U4038 (N_4038,N_3849,N_3938);
nor U4039 (N_4039,N_3914,N_3994);
and U4040 (N_4040,N_3968,N_3836);
xor U4041 (N_4041,N_3919,N_3972);
xor U4042 (N_4042,N_3820,N_3839);
and U4043 (N_4043,N_3831,N_3992);
nor U4044 (N_4044,N_3803,N_3999);
and U4045 (N_4045,N_3953,N_3966);
nor U4046 (N_4046,N_3821,N_3979);
and U4047 (N_4047,N_3924,N_3894);
nor U4048 (N_4048,N_3977,N_3910);
or U4049 (N_4049,N_3881,N_3997);
nor U4050 (N_4050,N_3907,N_3819);
nand U4051 (N_4051,N_3884,N_3895);
or U4052 (N_4052,N_3868,N_3955);
nor U4053 (N_4053,N_3838,N_3921);
and U4054 (N_4054,N_3826,N_3929);
nand U4055 (N_4055,N_3888,N_3908);
and U4056 (N_4056,N_3958,N_3982);
xnor U4057 (N_4057,N_3939,N_3925);
and U4058 (N_4058,N_3886,N_3829);
nand U4059 (N_4059,N_3865,N_3875);
nor U4060 (N_4060,N_3844,N_3974);
or U4061 (N_4061,N_3832,N_3889);
nor U4062 (N_4062,N_3835,N_3901);
and U4063 (N_4063,N_3959,N_3933);
nand U4064 (N_4064,N_3983,N_3810);
nand U4065 (N_4065,N_3817,N_3811);
and U4066 (N_4066,N_3861,N_3893);
or U4067 (N_4067,N_3950,N_3998);
and U4068 (N_4068,N_3864,N_3860);
nand U4069 (N_4069,N_3932,N_3954);
nand U4070 (N_4070,N_3986,N_3880);
and U4071 (N_4071,N_3871,N_3981);
nand U4072 (N_4072,N_3870,N_3885);
nand U4073 (N_4073,N_3911,N_3877);
and U4074 (N_4074,N_3899,N_3876);
nor U4075 (N_4075,N_3965,N_3805);
xnor U4076 (N_4076,N_3897,N_3971);
or U4077 (N_4077,N_3816,N_3852);
nand U4078 (N_4078,N_3869,N_3928);
nor U4079 (N_4079,N_3878,N_3980);
or U4080 (N_4080,N_3814,N_3913);
and U4081 (N_4081,N_3828,N_3975);
nand U4082 (N_4082,N_3909,N_3830);
and U4083 (N_4083,N_3804,N_3916);
and U4084 (N_4084,N_3802,N_3923);
nand U4085 (N_4085,N_3967,N_3859);
nor U4086 (N_4086,N_3976,N_3806);
and U4087 (N_4087,N_3931,N_3812);
or U4088 (N_4088,N_3942,N_3915);
and U4089 (N_4089,N_3990,N_3890);
nor U4090 (N_4090,N_3936,N_3824);
or U4091 (N_4091,N_3987,N_3825);
xor U4092 (N_4092,N_3883,N_3905);
xor U4093 (N_4093,N_3848,N_3855);
or U4094 (N_4094,N_3956,N_3898);
and U4095 (N_4095,N_3818,N_3862);
or U4096 (N_4096,N_3949,N_3842);
xor U4097 (N_4097,N_3946,N_3951);
or U4098 (N_4098,N_3947,N_3989);
xnor U4099 (N_4099,N_3853,N_3922);
and U4100 (N_4100,N_3832,N_3810);
xnor U4101 (N_4101,N_3980,N_3949);
nand U4102 (N_4102,N_3866,N_3834);
or U4103 (N_4103,N_3847,N_3872);
xor U4104 (N_4104,N_3838,N_3884);
nor U4105 (N_4105,N_3956,N_3949);
and U4106 (N_4106,N_3969,N_3819);
and U4107 (N_4107,N_3811,N_3884);
or U4108 (N_4108,N_3838,N_3897);
nand U4109 (N_4109,N_3968,N_3933);
or U4110 (N_4110,N_3920,N_3898);
or U4111 (N_4111,N_3819,N_3992);
or U4112 (N_4112,N_3890,N_3819);
and U4113 (N_4113,N_3906,N_3861);
nor U4114 (N_4114,N_3921,N_3917);
xor U4115 (N_4115,N_3821,N_3931);
xnor U4116 (N_4116,N_3890,N_3947);
nor U4117 (N_4117,N_3872,N_3803);
and U4118 (N_4118,N_3866,N_3943);
xnor U4119 (N_4119,N_3866,N_3996);
and U4120 (N_4120,N_3867,N_3842);
and U4121 (N_4121,N_3856,N_3806);
xor U4122 (N_4122,N_3900,N_3855);
and U4123 (N_4123,N_3959,N_3871);
or U4124 (N_4124,N_3991,N_3841);
or U4125 (N_4125,N_3954,N_3923);
nand U4126 (N_4126,N_3857,N_3977);
and U4127 (N_4127,N_3835,N_3852);
and U4128 (N_4128,N_3946,N_3977);
xnor U4129 (N_4129,N_3870,N_3818);
and U4130 (N_4130,N_3919,N_3959);
or U4131 (N_4131,N_3978,N_3954);
nor U4132 (N_4132,N_3969,N_3919);
nand U4133 (N_4133,N_3931,N_3911);
and U4134 (N_4134,N_3905,N_3921);
xor U4135 (N_4135,N_3954,N_3800);
or U4136 (N_4136,N_3900,N_3844);
or U4137 (N_4137,N_3983,N_3946);
and U4138 (N_4138,N_3848,N_3816);
and U4139 (N_4139,N_3921,N_3968);
nor U4140 (N_4140,N_3990,N_3822);
xor U4141 (N_4141,N_3947,N_3861);
or U4142 (N_4142,N_3961,N_3971);
nor U4143 (N_4143,N_3855,N_3913);
nor U4144 (N_4144,N_3970,N_3974);
or U4145 (N_4145,N_3873,N_3816);
nand U4146 (N_4146,N_3840,N_3815);
or U4147 (N_4147,N_3933,N_3981);
xnor U4148 (N_4148,N_3824,N_3844);
and U4149 (N_4149,N_3967,N_3978);
and U4150 (N_4150,N_3837,N_3839);
or U4151 (N_4151,N_3869,N_3843);
nand U4152 (N_4152,N_3923,N_3879);
nor U4153 (N_4153,N_3936,N_3983);
and U4154 (N_4154,N_3929,N_3939);
and U4155 (N_4155,N_3827,N_3992);
nor U4156 (N_4156,N_3894,N_3904);
xor U4157 (N_4157,N_3991,N_3995);
nor U4158 (N_4158,N_3932,N_3800);
nand U4159 (N_4159,N_3917,N_3816);
nor U4160 (N_4160,N_3804,N_3903);
or U4161 (N_4161,N_3912,N_3977);
nor U4162 (N_4162,N_3921,N_3847);
nor U4163 (N_4163,N_3908,N_3968);
or U4164 (N_4164,N_3969,N_3998);
and U4165 (N_4165,N_3871,N_3895);
nor U4166 (N_4166,N_3928,N_3806);
and U4167 (N_4167,N_3946,N_3913);
xor U4168 (N_4168,N_3995,N_3862);
xnor U4169 (N_4169,N_3802,N_3995);
or U4170 (N_4170,N_3940,N_3988);
or U4171 (N_4171,N_3813,N_3847);
and U4172 (N_4172,N_3959,N_3881);
nor U4173 (N_4173,N_3892,N_3886);
nand U4174 (N_4174,N_3800,N_3834);
and U4175 (N_4175,N_3873,N_3914);
xor U4176 (N_4176,N_3884,N_3962);
nor U4177 (N_4177,N_3868,N_3869);
and U4178 (N_4178,N_3888,N_3993);
nand U4179 (N_4179,N_3944,N_3864);
nor U4180 (N_4180,N_3813,N_3960);
nor U4181 (N_4181,N_3938,N_3918);
nor U4182 (N_4182,N_3901,N_3932);
nor U4183 (N_4183,N_3924,N_3810);
xnor U4184 (N_4184,N_3862,N_3811);
nor U4185 (N_4185,N_3974,N_3969);
xnor U4186 (N_4186,N_3840,N_3996);
nor U4187 (N_4187,N_3837,N_3899);
and U4188 (N_4188,N_3867,N_3825);
or U4189 (N_4189,N_3965,N_3854);
and U4190 (N_4190,N_3991,N_3897);
nand U4191 (N_4191,N_3831,N_3838);
or U4192 (N_4192,N_3828,N_3921);
and U4193 (N_4193,N_3965,N_3938);
nor U4194 (N_4194,N_3929,N_3824);
nor U4195 (N_4195,N_3857,N_3899);
nand U4196 (N_4196,N_3831,N_3908);
xor U4197 (N_4197,N_3971,N_3848);
and U4198 (N_4198,N_3872,N_3978);
and U4199 (N_4199,N_3826,N_3924);
nand U4200 (N_4200,N_4153,N_4012);
xor U4201 (N_4201,N_4180,N_4040);
and U4202 (N_4202,N_4007,N_4088);
nand U4203 (N_4203,N_4003,N_4161);
nand U4204 (N_4204,N_4001,N_4041);
nand U4205 (N_4205,N_4104,N_4191);
nor U4206 (N_4206,N_4190,N_4121);
nand U4207 (N_4207,N_4143,N_4124);
nor U4208 (N_4208,N_4128,N_4193);
nor U4209 (N_4209,N_4067,N_4147);
or U4210 (N_4210,N_4105,N_4032);
nand U4211 (N_4211,N_4078,N_4090);
nor U4212 (N_4212,N_4156,N_4099);
and U4213 (N_4213,N_4081,N_4069);
nor U4214 (N_4214,N_4176,N_4134);
nand U4215 (N_4215,N_4125,N_4070);
and U4216 (N_4216,N_4127,N_4182);
nand U4217 (N_4217,N_4021,N_4047);
or U4218 (N_4218,N_4058,N_4163);
and U4219 (N_4219,N_4157,N_4130);
nand U4220 (N_4220,N_4168,N_4133);
and U4221 (N_4221,N_4053,N_4137);
nor U4222 (N_4222,N_4165,N_4170);
xor U4223 (N_4223,N_4126,N_4174);
nand U4224 (N_4224,N_4109,N_4187);
nand U4225 (N_4225,N_4112,N_4148);
nor U4226 (N_4226,N_4000,N_4115);
xor U4227 (N_4227,N_4111,N_4195);
or U4228 (N_4228,N_4154,N_4030);
or U4229 (N_4229,N_4162,N_4085);
nand U4230 (N_4230,N_4082,N_4008);
and U4231 (N_4231,N_4114,N_4009);
nor U4232 (N_4232,N_4016,N_4188);
and U4233 (N_4233,N_4172,N_4089);
nand U4234 (N_4234,N_4118,N_4015);
nor U4235 (N_4235,N_4101,N_4092);
and U4236 (N_4236,N_4179,N_4066);
nand U4237 (N_4237,N_4005,N_4074);
or U4238 (N_4238,N_4098,N_4136);
nor U4239 (N_4239,N_4061,N_4094);
xnor U4240 (N_4240,N_4160,N_4034);
nand U4241 (N_4241,N_4029,N_4033);
nand U4242 (N_4242,N_4063,N_4166);
and U4243 (N_4243,N_4080,N_4028);
nor U4244 (N_4244,N_4102,N_4055);
nor U4245 (N_4245,N_4019,N_4026);
nand U4246 (N_4246,N_4046,N_4049);
nand U4247 (N_4247,N_4171,N_4158);
or U4248 (N_4248,N_4135,N_4199);
nand U4249 (N_4249,N_4076,N_4065);
nand U4250 (N_4250,N_4096,N_4037);
nand U4251 (N_4251,N_4140,N_4039);
xnor U4252 (N_4252,N_4149,N_4079);
and U4253 (N_4253,N_4084,N_4184);
or U4254 (N_4254,N_4011,N_4038);
nor U4255 (N_4255,N_4044,N_4159);
and U4256 (N_4256,N_4010,N_4062);
nor U4257 (N_4257,N_4192,N_4116);
nor U4258 (N_4258,N_4177,N_4042);
or U4259 (N_4259,N_4017,N_4167);
xnor U4260 (N_4260,N_4151,N_4072);
nor U4261 (N_4261,N_4093,N_4054);
or U4262 (N_4262,N_4013,N_4048);
or U4263 (N_4263,N_4050,N_4097);
nand U4264 (N_4264,N_4131,N_4014);
nand U4265 (N_4265,N_4064,N_4119);
or U4266 (N_4266,N_4175,N_4106);
nand U4267 (N_4267,N_4043,N_4071);
and U4268 (N_4268,N_4113,N_4183);
or U4269 (N_4269,N_4138,N_4132);
or U4270 (N_4270,N_4024,N_4129);
nand U4271 (N_4271,N_4068,N_4152);
nor U4272 (N_4272,N_4178,N_4117);
xnor U4273 (N_4273,N_4075,N_4052);
nand U4274 (N_4274,N_4077,N_4155);
and U4275 (N_4275,N_4181,N_4036);
nor U4276 (N_4276,N_4146,N_4022);
nand U4277 (N_4277,N_4122,N_4145);
nand U4278 (N_4278,N_4051,N_4169);
nand U4279 (N_4279,N_4027,N_4006);
nor U4280 (N_4280,N_4107,N_4103);
nand U4281 (N_4281,N_4031,N_4059);
nor U4282 (N_4282,N_4186,N_4110);
nand U4283 (N_4283,N_4057,N_4073);
nor U4284 (N_4284,N_4189,N_4141);
nor U4285 (N_4285,N_4164,N_4194);
or U4286 (N_4286,N_4150,N_4087);
xor U4287 (N_4287,N_4173,N_4108);
or U4288 (N_4288,N_4091,N_4086);
and U4289 (N_4289,N_4196,N_4100);
nand U4290 (N_4290,N_4197,N_4144);
nand U4291 (N_4291,N_4025,N_4123);
or U4292 (N_4292,N_4095,N_4060);
and U4293 (N_4293,N_4023,N_4004);
xor U4294 (N_4294,N_4035,N_4018);
and U4295 (N_4295,N_4120,N_4185);
or U4296 (N_4296,N_4083,N_4045);
nand U4297 (N_4297,N_4056,N_4198);
and U4298 (N_4298,N_4139,N_4020);
nand U4299 (N_4299,N_4002,N_4142);
nand U4300 (N_4300,N_4149,N_4002);
and U4301 (N_4301,N_4015,N_4016);
and U4302 (N_4302,N_4045,N_4143);
xor U4303 (N_4303,N_4008,N_4043);
nor U4304 (N_4304,N_4095,N_4061);
or U4305 (N_4305,N_4026,N_4177);
and U4306 (N_4306,N_4043,N_4106);
or U4307 (N_4307,N_4087,N_4198);
and U4308 (N_4308,N_4106,N_4006);
or U4309 (N_4309,N_4023,N_4041);
nand U4310 (N_4310,N_4172,N_4097);
nor U4311 (N_4311,N_4102,N_4008);
or U4312 (N_4312,N_4041,N_4118);
or U4313 (N_4313,N_4090,N_4051);
and U4314 (N_4314,N_4177,N_4137);
nand U4315 (N_4315,N_4081,N_4101);
and U4316 (N_4316,N_4131,N_4024);
nand U4317 (N_4317,N_4100,N_4072);
and U4318 (N_4318,N_4154,N_4061);
and U4319 (N_4319,N_4045,N_4181);
nand U4320 (N_4320,N_4043,N_4104);
and U4321 (N_4321,N_4165,N_4105);
and U4322 (N_4322,N_4095,N_4055);
nand U4323 (N_4323,N_4055,N_4181);
nor U4324 (N_4324,N_4040,N_4052);
xor U4325 (N_4325,N_4164,N_4082);
or U4326 (N_4326,N_4119,N_4061);
xnor U4327 (N_4327,N_4081,N_4067);
xor U4328 (N_4328,N_4140,N_4025);
or U4329 (N_4329,N_4002,N_4014);
nor U4330 (N_4330,N_4096,N_4179);
or U4331 (N_4331,N_4013,N_4086);
or U4332 (N_4332,N_4076,N_4173);
xor U4333 (N_4333,N_4108,N_4154);
nand U4334 (N_4334,N_4097,N_4071);
nor U4335 (N_4335,N_4168,N_4001);
or U4336 (N_4336,N_4074,N_4168);
nand U4337 (N_4337,N_4197,N_4044);
nand U4338 (N_4338,N_4055,N_4080);
and U4339 (N_4339,N_4199,N_4170);
or U4340 (N_4340,N_4154,N_4103);
nor U4341 (N_4341,N_4111,N_4004);
or U4342 (N_4342,N_4079,N_4196);
or U4343 (N_4343,N_4101,N_4089);
nand U4344 (N_4344,N_4067,N_4148);
nand U4345 (N_4345,N_4046,N_4171);
or U4346 (N_4346,N_4056,N_4176);
nand U4347 (N_4347,N_4098,N_4094);
or U4348 (N_4348,N_4167,N_4063);
nand U4349 (N_4349,N_4093,N_4175);
nor U4350 (N_4350,N_4025,N_4179);
xor U4351 (N_4351,N_4060,N_4171);
nor U4352 (N_4352,N_4190,N_4023);
nand U4353 (N_4353,N_4017,N_4048);
and U4354 (N_4354,N_4062,N_4002);
nor U4355 (N_4355,N_4102,N_4195);
or U4356 (N_4356,N_4174,N_4047);
or U4357 (N_4357,N_4171,N_4157);
nand U4358 (N_4358,N_4101,N_4044);
and U4359 (N_4359,N_4114,N_4090);
or U4360 (N_4360,N_4197,N_4181);
nand U4361 (N_4361,N_4032,N_4145);
nor U4362 (N_4362,N_4144,N_4086);
xor U4363 (N_4363,N_4048,N_4104);
xnor U4364 (N_4364,N_4192,N_4120);
xor U4365 (N_4365,N_4040,N_4095);
nand U4366 (N_4366,N_4177,N_4077);
xnor U4367 (N_4367,N_4167,N_4162);
nor U4368 (N_4368,N_4122,N_4084);
nor U4369 (N_4369,N_4073,N_4076);
and U4370 (N_4370,N_4184,N_4122);
and U4371 (N_4371,N_4062,N_4054);
and U4372 (N_4372,N_4059,N_4196);
xor U4373 (N_4373,N_4109,N_4183);
nand U4374 (N_4374,N_4044,N_4153);
nand U4375 (N_4375,N_4194,N_4184);
or U4376 (N_4376,N_4149,N_4194);
nor U4377 (N_4377,N_4038,N_4075);
or U4378 (N_4378,N_4135,N_4128);
nor U4379 (N_4379,N_4110,N_4054);
nor U4380 (N_4380,N_4037,N_4002);
and U4381 (N_4381,N_4057,N_4040);
nand U4382 (N_4382,N_4089,N_4083);
nor U4383 (N_4383,N_4103,N_4167);
nand U4384 (N_4384,N_4024,N_4080);
nor U4385 (N_4385,N_4154,N_4057);
nor U4386 (N_4386,N_4106,N_4045);
xor U4387 (N_4387,N_4141,N_4087);
xor U4388 (N_4388,N_4038,N_4072);
or U4389 (N_4389,N_4045,N_4040);
nand U4390 (N_4390,N_4158,N_4110);
nand U4391 (N_4391,N_4189,N_4128);
nand U4392 (N_4392,N_4026,N_4160);
or U4393 (N_4393,N_4090,N_4098);
or U4394 (N_4394,N_4150,N_4199);
nand U4395 (N_4395,N_4119,N_4045);
nor U4396 (N_4396,N_4002,N_4044);
nor U4397 (N_4397,N_4172,N_4008);
and U4398 (N_4398,N_4078,N_4144);
and U4399 (N_4399,N_4166,N_4066);
xor U4400 (N_4400,N_4242,N_4229);
nand U4401 (N_4401,N_4321,N_4305);
and U4402 (N_4402,N_4323,N_4210);
or U4403 (N_4403,N_4222,N_4267);
nor U4404 (N_4404,N_4353,N_4299);
nor U4405 (N_4405,N_4304,N_4302);
or U4406 (N_4406,N_4324,N_4283);
or U4407 (N_4407,N_4383,N_4354);
xor U4408 (N_4408,N_4358,N_4385);
or U4409 (N_4409,N_4284,N_4348);
xor U4410 (N_4410,N_4379,N_4257);
or U4411 (N_4411,N_4307,N_4237);
and U4412 (N_4412,N_4349,N_4360);
xnor U4413 (N_4413,N_4376,N_4327);
and U4414 (N_4414,N_4317,N_4281);
nand U4415 (N_4415,N_4244,N_4238);
nand U4416 (N_4416,N_4249,N_4315);
xnor U4417 (N_4417,N_4256,N_4314);
or U4418 (N_4418,N_4286,N_4365);
nand U4419 (N_4419,N_4263,N_4241);
or U4420 (N_4420,N_4303,N_4396);
xor U4421 (N_4421,N_4328,N_4250);
xnor U4422 (N_4422,N_4220,N_4293);
nor U4423 (N_4423,N_4217,N_4363);
nor U4424 (N_4424,N_4260,N_4208);
nand U4425 (N_4425,N_4268,N_4290);
nor U4426 (N_4426,N_4212,N_4342);
and U4427 (N_4427,N_4319,N_4254);
nand U4428 (N_4428,N_4356,N_4326);
nand U4429 (N_4429,N_4341,N_4334);
nand U4430 (N_4430,N_4214,N_4394);
nand U4431 (N_4431,N_4343,N_4294);
or U4432 (N_4432,N_4378,N_4248);
nor U4433 (N_4433,N_4310,N_4357);
nand U4434 (N_4434,N_4344,N_4308);
or U4435 (N_4435,N_4398,N_4235);
and U4436 (N_4436,N_4245,N_4399);
and U4437 (N_4437,N_4228,N_4339);
nand U4438 (N_4438,N_4374,N_4355);
xor U4439 (N_4439,N_4289,N_4211);
nor U4440 (N_4440,N_4336,N_4261);
or U4441 (N_4441,N_4346,N_4351);
nand U4442 (N_4442,N_4366,N_4338);
or U4443 (N_4443,N_4275,N_4227);
and U4444 (N_4444,N_4239,N_4361);
nor U4445 (N_4445,N_4313,N_4331);
or U4446 (N_4446,N_4219,N_4236);
nand U4447 (N_4447,N_4345,N_4269);
or U4448 (N_4448,N_4373,N_4259);
nand U4449 (N_4449,N_4230,N_4359);
nand U4450 (N_4450,N_4362,N_4368);
nand U4451 (N_4451,N_4320,N_4364);
or U4452 (N_4452,N_4382,N_4340);
or U4453 (N_4453,N_4395,N_4312);
nor U4454 (N_4454,N_4300,N_4271);
and U4455 (N_4455,N_4246,N_4280);
or U4456 (N_4456,N_4380,N_4252);
or U4457 (N_4457,N_4215,N_4367);
or U4458 (N_4458,N_4296,N_4387);
nor U4459 (N_4459,N_4391,N_4311);
or U4460 (N_4460,N_4265,N_4301);
and U4461 (N_4461,N_4234,N_4233);
nor U4462 (N_4462,N_4332,N_4279);
xor U4463 (N_4463,N_4277,N_4285);
or U4464 (N_4464,N_4292,N_4390);
nand U4465 (N_4465,N_4272,N_4209);
xor U4466 (N_4466,N_4213,N_4266);
and U4467 (N_4467,N_4270,N_4218);
nand U4468 (N_4468,N_4258,N_4381);
or U4469 (N_4469,N_4287,N_4243);
nand U4470 (N_4470,N_4200,N_4333);
nor U4471 (N_4471,N_4202,N_4264);
nor U4472 (N_4472,N_4224,N_4226);
nor U4473 (N_4473,N_4397,N_4370);
and U4474 (N_4474,N_4204,N_4288);
and U4475 (N_4475,N_4347,N_4203);
or U4476 (N_4476,N_4225,N_4389);
nand U4477 (N_4477,N_4274,N_4206);
nor U4478 (N_4478,N_4371,N_4278);
or U4479 (N_4479,N_4322,N_4247);
nand U4480 (N_4480,N_4240,N_4375);
or U4481 (N_4481,N_4309,N_4207);
and U4482 (N_4482,N_4291,N_4295);
nand U4483 (N_4483,N_4325,N_4350);
xor U4484 (N_4484,N_4232,N_4386);
or U4485 (N_4485,N_4255,N_4329);
nor U4486 (N_4486,N_4372,N_4388);
and U4487 (N_4487,N_4282,N_4262);
or U4488 (N_4488,N_4393,N_4276);
nor U4489 (N_4489,N_4316,N_4221);
and U4490 (N_4490,N_4251,N_4337);
nor U4491 (N_4491,N_4298,N_4377);
nand U4492 (N_4492,N_4216,N_4273);
nand U4493 (N_4493,N_4201,N_4253);
xnor U4494 (N_4494,N_4352,N_4231);
nand U4495 (N_4495,N_4306,N_4335);
and U4496 (N_4496,N_4384,N_4223);
nor U4497 (N_4497,N_4318,N_4205);
nand U4498 (N_4498,N_4330,N_4297);
nand U4499 (N_4499,N_4392,N_4369);
or U4500 (N_4500,N_4323,N_4380);
and U4501 (N_4501,N_4268,N_4285);
or U4502 (N_4502,N_4385,N_4252);
nor U4503 (N_4503,N_4236,N_4306);
and U4504 (N_4504,N_4264,N_4270);
nor U4505 (N_4505,N_4357,N_4333);
or U4506 (N_4506,N_4361,N_4298);
xnor U4507 (N_4507,N_4276,N_4315);
or U4508 (N_4508,N_4256,N_4333);
and U4509 (N_4509,N_4221,N_4207);
nand U4510 (N_4510,N_4329,N_4341);
nand U4511 (N_4511,N_4329,N_4260);
or U4512 (N_4512,N_4389,N_4254);
nand U4513 (N_4513,N_4304,N_4343);
or U4514 (N_4514,N_4214,N_4263);
xnor U4515 (N_4515,N_4228,N_4259);
nor U4516 (N_4516,N_4297,N_4227);
nand U4517 (N_4517,N_4216,N_4230);
or U4518 (N_4518,N_4303,N_4389);
and U4519 (N_4519,N_4228,N_4270);
and U4520 (N_4520,N_4230,N_4233);
xor U4521 (N_4521,N_4329,N_4242);
nor U4522 (N_4522,N_4354,N_4386);
nor U4523 (N_4523,N_4364,N_4373);
and U4524 (N_4524,N_4259,N_4357);
nand U4525 (N_4525,N_4399,N_4333);
nand U4526 (N_4526,N_4383,N_4300);
and U4527 (N_4527,N_4236,N_4349);
and U4528 (N_4528,N_4254,N_4209);
or U4529 (N_4529,N_4211,N_4328);
nor U4530 (N_4530,N_4297,N_4382);
nor U4531 (N_4531,N_4299,N_4355);
nor U4532 (N_4532,N_4201,N_4248);
xnor U4533 (N_4533,N_4276,N_4361);
or U4534 (N_4534,N_4317,N_4302);
or U4535 (N_4535,N_4332,N_4337);
nor U4536 (N_4536,N_4233,N_4340);
xor U4537 (N_4537,N_4300,N_4365);
nor U4538 (N_4538,N_4268,N_4238);
nand U4539 (N_4539,N_4348,N_4248);
nand U4540 (N_4540,N_4204,N_4272);
or U4541 (N_4541,N_4333,N_4384);
xor U4542 (N_4542,N_4393,N_4283);
or U4543 (N_4543,N_4366,N_4269);
or U4544 (N_4544,N_4281,N_4313);
or U4545 (N_4545,N_4242,N_4383);
nor U4546 (N_4546,N_4374,N_4393);
nor U4547 (N_4547,N_4271,N_4204);
nand U4548 (N_4548,N_4381,N_4314);
or U4549 (N_4549,N_4332,N_4334);
nand U4550 (N_4550,N_4393,N_4341);
and U4551 (N_4551,N_4378,N_4364);
nor U4552 (N_4552,N_4370,N_4261);
nor U4553 (N_4553,N_4349,N_4225);
xnor U4554 (N_4554,N_4382,N_4289);
or U4555 (N_4555,N_4272,N_4361);
or U4556 (N_4556,N_4334,N_4284);
and U4557 (N_4557,N_4215,N_4332);
or U4558 (N_4558,N_4324,N_4273);
and U4559 (N_4559,N_4388,N_4232);
and U4560 (N_4560,N_4289,N_4352);
and U4561 (N_4561,N_4234,N_4237);
nand U4562 (N_4562,N_4200,N_4250);
nor U4563 (N_4563,N_4229,N_4381);
or U4564 (N_4564,N_4347,N_4310);
and U4565 (N_4565,N_4355,N_4226);
and U4566 (N_4566,N_4218,N_4225);
or U4567 (N_4567,N_4204,N_4366);
or U4568 (N_4568,N_4245,N_4353);
nor U4569 (N_4569,N_4396,N_4251);
nor U4570 (N_4570,N_4228,N_4354);
nor U4571 (N_4571,N_4254,N_4316);
and U4572 (N_4572,N_4214,N_4278);
nand U4573 (N_4573,N_4288,N_4359);
nor U4574 (N_4574,N_4357,N_4350);
or U4575 (N_4575,N_4320,N_4266);
nand U4576 (N_4576,N_4339,N_4376);
nand U4577 (N_4577,N_4381,N_4367);
nor U4578 (N_4578,N_4246,N_4260);
nand U4579 (N_4579,N_4379,N_4353);
and U4580 (N_4580,N_4275,N_4268);
xnor U4581 (N_4581,N_4247,N_4300);
xor U4582 (N_4582,N_4386,N_4374);
and U4583 (N_4583,N_4223,N_4251);
nor U4584 (N_4584,N_4266,N_4237);
and U4585 (N_4585,N_4292,N_4207);
and U4586 (N_4586,N_4355,N_4254);
or U4587 (N_4587,N_4213,N_4240);
or U4588 (N_4588,N_4230,N_4345);
or U4589 (N_4589,N_4350,N_4258);
nand U4590 (N_4590,N_4382,N_4394);
xor U4591 (N_4591,N_4288,N_4263);
and U4592 (N_4592,N_4393,N_4359);
and U4593 (N_4593,N_4277,N_4228);
nand U4594 (N_4594,N_4243,N_4266);
or U4595 (N_4595,N_4243,N_4382);
or U4596 (N_4596,N_4253,N_4394);
nor U4597 (N_4597,N_4243,N_4388);
nand U4598 (N_4598,N_4226,N_4262);
or U4599 (N_4599,N_4382,N_4255);
nor U4600 (N_4600,N_4400,N_4509);
xnor U4601 (N_4601,N_4540,N_4422);
nor U4602 (N_4602,N_4404,N_4588);
and U4603 (N_4603,N_4459,N_4458);
nand U4604 (N_4604,N_4558,N_4518);
nand U4605 (N_4605,N_4473,N_4541);
and U4606 (N_4606,N_4408,N_4599);
or U4607 (N_4607,N_4584,N_4546);
or U4608 (N_4608,N_4500,N_4534);
nand U4609 (N_4609,N_4427,N_4550);
nor U4610 (N_4610,N_4522,N_4573);
or U4611 (N_4611,N_4549,N_4590);
nor U4612 (N_4612,N_4455,N_4401);
nor U4613 (N_4613,N_4499,N_4508);
or U4614 (N_4614,N_4438,N_4463);
or U4615 (N_4615,N_4567,N_4461);
nor U4616 (N_4616,N_4468,N_4495);
nand U4617 (N_4617,N_4505,N_4587);
and U4618 (N_4618,N_4494,N_4561);
nand U4619 (N_4619,N_4476,N_4426);
nand U4620 (N_4620,N_4435,N_4585);
and U4621 (N_4621,N_4555,N_4409);
nor U4622 (N_4622,N_4579,N_4523);
nand U4623 (N_4623,N_4592,N_4413);
nor U4624 (N_4624,N_4568,N_4517);
xor U4625 (N_4625,N_4563,N_4524);
nand U4626 (N_4626,N_4582,N_4544);
xor U4627 (N_4627,N_4481,N_4569);
nor U4628 (N_4628,N_4591,N_4595);
xor U4629 (N_4629,N_4445,N_4493);
and U4630 (N_4630,N_4478,N_4535);
nand U4631 (N_4631,N_4472,N_4559);
or U4632 (N_4632,N_4420,N_4487);
or U4633 (N_4633,N_4529,N_4449);
or U4634 (N_4634,N_4521,N_4410);
or U4635 (N_4635,N_4431,N_4471);
and U4636 (N_4636,N_4530,N_4479);
xnor U4637 (N_4637,N_4432,N_4593);
and U4638 (N_4638,N_4498,N_4553);
xor U4639 (N_4639,N_4531,N_4489);
nand U4640 (N_4640,N_4441,N_4492);
nor U4641 (N_4641,N_4439,N_4528);
or U4642 (N_4642,N_4543,N_4403);
and U4643 (N_4643,N_4421,N_4467);
xor U4644 (N_4644,N_4580,N_4510);
and U4645 (N_4645,N_4566,N_4511);
or U4646 (N_4646,N_4594,N_4576);
nand U4647 (N_4647,N_4417,N_4424);
nand U4648 (N_4648,N_4462,N_4453);
or U4649 (N_4649,N_4571,N_4416);
or U4650 (N_4650,N_4469,N_4497);
and U4651 (N_4651,N_4452,N_4564);
nand U4652 (N_4652,N_4548,N_4457);
nand U4653 (N_4653,N_4434,N_4488);
nand U4654 (N_4654,N_4414,N_4433);
or U4655 (N_4655,N_4464,N_4485);
and U4656 (N_4656,N_4406,N_4556);
or U4657 (N_4657,N_4597,N_4527);
nand U4658 (N_4658,N_4430,N_4419);
nor U4659 (N_4659,N_4554,N_4547);
xnor U4660 (N_4660,N_4436,N_4537);
or U4661 (N_4661,N_4502,N_4480);
or U4662 (N_4662,N_4415,N_4525);
and U4663 (N_4663,N_4565,N_4513);
or U4664 (N_4664,N_4557,N_4470);
nand U4665 (N_4665,N_4519,N_4581);
nor U4666 (N_4666,N_4503,N_4577);
and U4667 (N_4667,N_4538,N_4574);
and U4668 (N_4668,N_4454,N_4533);
xnor U4669 (N_4669,N_4405,N_4411);
nand U4670 (N_4670,N_4545,N_4496);
nand U4671 (N_4671,N_4583,N_4578);
nor U4672 (N_4672,N_4572,N_4570);
and U4673 (N_4673,N_4516,N_4466);
and U4674 (N_4674,N_4475,N_4440);
nor U4675 (N_4675,N_4477,N_4491);
xnor U4676 (N_4676,N_4443,N_4423);
or U4677 (N_4677,N_4490,N_4504);
and U4678 (N_4678,N_4586,N_4446);
and U4679 (N_4679,N_4460,N_4482);
xnor U4680 (N_4680,N_4437,N_4486);
nand U4681 (N_4681,N_4551,N_4539);
or U4682 (N_4682,N_4515,N_4444);
nor U4683 (N_4683,N_4418,N_4407);
nand U4684 (N_4684,N_4575,N_4447);
nor U4685 (N_4685,N_4456,N_4514);
nor U4686 (N_4686,N_4520,N_4402);
nand U4687 (N_4687,N_4474,N_4484);
nor U4688 (N_4688,N_4483,N_4425);
and U4689 (N_4689,N_4442,N_4512);
or U4690 (N_4690,N_4451,N_4428);
or U4691 (N_4691,N_4562,N_4542);
xnor U4692 (N_4692,N_4560,N_4465);
and U4693 (N_4693,N_4596,N_4536);
and U4694 (N_4694,N_4589,N_4429);
nand U4695 (N_4695,N_4506,N_4448);
nand U4696 (N_4696,N_4412,N_4507);
or U4697 (N_4697,N_4526,N_4450);
nor U4698 (N_4698,N_4501,N_4598);
and U4699 (N_4699,N_4532,N_4552);
or U4700 (N_4700,N_4510,N_4411);
nand U4701 (N_4701,N_4403,N_4477);
nor U4702 (N_4702,N_4444,N_4415);
nand U4703 (N_4703,N_4518,N_4422);
nor U4704 (N_4704,N_4482,N_4565);
or U4705 (N_4705,N_4476,N_4539);
nor U4706 (N_4706,N_4572,N_4480);
nor U4707 (N_4707,N_4453,N_4538);
nor U4708 (N_4708,N_4589,N_4583);
or U4709 (N_4709,N_4571,N_4448);
or U4710 (N_4710,N_4527,N_4591);
nor U4711 (N_4711,N_4501,N_4454);
or U4712 (N_4712,N_4598,N_4422);
nand U4713 (N_4713,N_4435,N_4500);
nand U4714 (N_4714,N_4426,N_4554);
nor U4715 (N_4715,N_4562,N_4587);
xor U4716 (N_4716,N_4458,N_4583);
and U4717 (N_4717,N_4400,N_4477);
nand U4718 (N_4718,N_4584,N_4497);
nor U4719 (N_4719,N_4548,N_4503);
nor U4720 (N_4720,N_4569,N_4451);
or U4721 (N_4721,N_4469,N_4435);
and U4722 (N_4722,N_4432,N_4553);
nand U4723 (N_4723,N_4589,N_4467);
nand U4724 (N_4724,N_4532,N_4408);
nor U4725 (N_4725,N_4578,N_4405);
and U4726 (N_4726,N_4521,N_4557);
and U4727 (N_4727,N_4541,N_4480);
xnor U4728 (N_4728,N_4428,N_4482);
xor U4729 (N_4729,N_4551,N_4480);
xor U4730 (N_4730,N_4507,N_4413);
nor U4731 (N_4731,N_4400,N_4420);
nor U4732 (N_4732,N_4407,N_4472);
nor U4733 (N_4733,N_4467,N_4571);
nand U4734 (N_4734,N_4596,N_4560);
and U4735 (N_4735,N_4595,N_4411);
nand U4736 (N_4736,N_4529,N_4404);
nor U4737 (N_4737,N_4435,N_4522);
nand U4738 (N_4738,N_4450,N_4425);
nor U4739 (N_4739,N_4513,N_4579);
nor U4740 (N_4740,N_4548,N_4538);
xor U4741 (N_4741,N_4538,N_4435);
nand U4742 (N_4742,N_4585,N_4409);
and U4743 (N_4743,N_4584,N_4506);
nor U4744 (N_4744,N_4557,N_4529);
nor U4745 (N_4745,N_4465,N_4446);
nand U4746 (N_4746,N_4475,N_4480);
nand U4747 (N_4747,N_4572,N_4597);
nor U4748 (N_4748,N_4545,N_4543);
nand U4749 (N_4749,N_4537,N_4541);
xnor U4750 (N_4750,N_4450,N_4485);
xnor U4751 (N_4751,N_4419,N_4496);
or U4752 (N_4752,N_4410,N_4447);
or U4753 (N_4753,N_4567,N_4580);
nor U4754 (N_4754,N_4597,N_4579);
or U4755 (N_4755,N_4545,N_4428);
nor U4756 (N_4756,N_4447,N_4536);
nand U4757 (N_4757,N_4469,N_4521);
or U4758 (N_4758,N_4407,N_4550);
nand U4759 (N_4759,N_4467,N_4553);
nand U4760 (N_4760,N_4447,N_4453);
and U4761 (N_4761,N_4584,N_4424);
and U4762 (N_4762,N_4450,N_4596);
and U4763 (N_4763,N_4511,N_4496);
nand U4764 (N_4764,N_4580,N_4570);
nor U4765 (N_4765,N_4479,N_4451);
nand U4766 (N_4766,N_4477,N_4540);
and U4767 (N_4767,N_4443,N_4485);
or U4768 (N_4768,N_4496,N_4515);
or U4769 (N_4769,N_4496,N_4497);
nor U4770 (N_4770,N_4557,N_4463);
and U4771 (N_4771,N_4577,N_4562);
nand U4772 (N_4772,N_4589,N_4508);
nor U4773 (N_4773,N_4558,N_4557);
nand U4774 (N_4774,N_4568,N_4582);
xnor U4775 (N_4775,N_4499,N_4529);
nor U4776 (N_4776,N_4536,N_4438);
or U4777 (N_4777,N_4492,N_4510);
nor U4778 (N_4778,N_4410,N_4503);
or U4779 (N_4779,N_4453,N_4532);
nor U4780 (N_4780,N_4442,N_4488);
and U4781 (N_4781,N_4491,N_4490);
or U4782 (N_4782,N_4412,N_4468);
nor U4783 (N_4783,N_4499,N_4428);
nand U4784 (N_4784,N_4544,N_4559);
or U4785 (N_4785,N_4510,N_4473);
nand U4786 (N_4786,N_4529,N_4575);
xnor U4787 (N_4787,N_4489,N_4496);
or U4788 (N_4788,N_4443,N_4446);
nor U4789 (N_4789,N_4435,N_4572);
and U4790 (N_4790,N_4531,N_4455);
nand U4791 (N_4791,N_4510,N_4433);
xor U4792 (N_4792,N_4587,N_4499);
nor U4793 (N_4793,N_4415,N_4534);
or U4794 (N_4794,N_4461,N_4527);
nand U4795 (N_4795,N_4488,N_4573);
nor U4796 (N_4796,N_4481,N_4537);
or U4797 (N_4797,N_4458,N_4564);
or U4798 (N_4798,N_4579,N_4576);
xnor U4799 (N_4799,N_4458,N_4596);
or U4800 (N_4800,N_4708,N_4780);
and U4801 (N_4801,N_4767,N_4739);
and U4802 (N_4802,N_4710,N_4688);
nand U4803 (N_4803,N_4674,N_4714);
or U4804 (N_4804,N_4720,N_4751);
or U4805 (N_4805,N_4625,N_4776);
or U4806 (N_4806,N_4771,N_4635);
or U4807 (N_4807,N_4675,N_4643);
and U4808 (N_4808,N_4686,N_4730);
nor U4809 (N_4809,N_4659,N_4784);
nand U4810 (N_4810,N_4658,N_4690);
or U4811 (N_4811,N_4715,N_4744);
and U4812 (N_4812,N_4761,N_4754);
or U4813 (N_4813,N_4651,N_4728);
nor U4814 (N_4814,N_4612,N_4729);
or U4815 (N_4815,N_4750,N_4770);
xnor U4816 (N_4816,N_4746,N_4704);
or U4817 (N_4817,N_4724,N_4657);
or U4818 (N_4818,N_4640,N_4788);
nor U4819 (N_4819,N_4733,N_4673);
xnor U4820 (N_4820,N_4684,N_4637);
nand U4821 (N_4821,N_4631,N_4752);
xor U4822 (N_4822,N_4772,N_4722);
nand U4823 (N_4823,N_4756,N_4636);
nand U4824 (N_4824,N_4623,N_4793);
nand U4825 (N_4825,N_4757,N_4662);
nor U4826 (N_4826,N_4743,N_4749);
nand U4827 (N_4827,N_4796,N_4701);
or U4828 (N_4828,N_4671,N_4647);
and U4829 (N_4829,N_4648,N_4614);
nand U4830 (N_4830,N_4755,N_4607);
or U4831 (N_4831,N_4629,N_4791);
nand U4832 (N_4832,N_4680,N_4669);
or U4833 (N_4833,N_4610,N_4609);
nand U4834 (N_4834,N_4721,N_4663);
nor U4835 (N_4835,N_4695,N_4736);
or U4836 (N_4836,N_4759,N_4691);
nand U4837 (N_4837,N_4799,N_4785);
nor U4838 (N_4838,N_4653,N_4689);
nand U4839 (N_4839,N_4670,N_4668);
nand U4840 (N_4840,N_4678,N_4617);
and U4841 (N_4841,N_4604,N_4696);
nor U4842 (N_4842,N_4798,N_4646);
nor U4843 (N_4843,N_4605,N_4719);
or U4844 (N_4844,N_4633,N_4745);
nand U4845 (N_4845,N_4705,N_4713);
and U4846 (N_4846,N_4748,N_4621);
nand U4847 (N_4847,N_4781,N_4606);
nand U4848 (N_4848,N_4716,N_4717);
nand U4849 (N_4849,N_4773,N_4774);
and U4850 (N_4850,N_4782,N_4718);
nor U4851 (N_4851,N_4735,N_4732);
or U4852 (N_4852,N_4619,N_4765);
nor U4853 (N_4853,N_4723,N_4787);
and U4854 (N_4854,N_4602,N_4679);
or U4855 (N_4855,N_4666,N_4709);
nand U4856 (N_4856,N_4779,N_4726);
nor U4857 (N_4857,N_4792,N_4616);
or U4858 (N_4858,N_4766,N_4664);
or U4859 (N_4859,N_4794,N_4763);
nand U4860 (N_4860,N_4632,N_4697);
nand U4861 (N_4861,N_4775,N_4677);
or U4862 (N_4862,N_4630,N_4639);
xnor U4863 (N_4863,N_4661,N_4762);
nand U4864 (N_4864,N_4613,N_4638);
or U4865 (N_4865,N_4702,N_4711);
and U4866 (N_4866,N_4665,N_4611);
nand U4867 (N_4867,N_4676,N_4737);
nor U4868 (N_4868,N_4760,N_4620);
or U4869 (N_4869,N_4797,N_4764);
nand U4870 (N_4870,N_4660,N_4795);
nand U4871 (N_4871,N_4628,N_4769);
and U4872 (N_4872,N_4789,N_4699);
nand U4873 (N_4873,N_4667,N_4747);
nand U4874 (N_4874,N_4706,N_4624);
or U4875 (N_4875,N_4603,N_4727);
and U4876 (N_4876,N_4742,N_4634);
nand U4877 (N_4877,N_4707,N_4650);
nor U4878 (N_4878,N_4703,N_4683);
xnor U4879 (N_4879,N_4740,N_4655);
nor U4880 (N_4880,N_4645,N_4692);
nand U4881 (N_4881,N_4786,N_4694);
or U4882 (N_4882,N_4778,N_4622);
nand U4883 (N_4883,N_4601,N_4725);
xnor U4884 (N_4884,N_4753,N_4627);
or U4885 (N_4885,N_4790,N_4641);
and U4886 (N_4886,N_4741,N_4777);
and U4887 (N_4887,N_4672,N_4768);
nor U4888 (N_4888,N_4700,N_4738);
nor U4889 (N_4889,N_4698,N_4758);
and U4890 (N_4890,N_4681,N_4644);
xnor U4891 (N_4891,N_4654,N_4731);
nand U4892 (N_4892,N_4712,N_4734);
and U4893 (N_4893,N_4649,N_4687);
and U4894 (N_4894,N_4642,N_4656);
nor U4895 (N_4895,N_4600,N_4615);
nor U4896 (N_4896,N_4652,N_4608);
nor U4897 (N_4897,N_4685,N_4618);
nand U4898 (N_4898,N_4682,N_4783);
nand U4899 (N_4899,N_4626,N_4693);
nor U4900 (N_4900,N_4661,N_4695);
and U4901 (N_4901,N_4657,N_4686);
nor U4902 (N_4902,N_4611,N_4682);
or U4903 (N_4903,N_4796,N_4602);
or U4904 (N_4904,N_4760,N_4786);
nand U4905 (N_4905,N_4660,N_4679);
and U4906 (N_4906,N_4789,N_4798);
and U4907 (N_4907,N_4738,N_4732);
nor U4908 (N_4908,N_4682,N_4705);
nand U4909 (N_4909,N_4606,N_4745);
nand U4910 (N_4910,N_4728,N_4695);
nand U4911 (N_4911,N_4661,N_4789);
nand U4912 (N_4912,N_4749,N_4703);
and U4913 (N_4913,N_4736,N_4664);
or U4914 (N_4914,N_4745,N_4623);
nor U4915 (N_4915,N_4622,N_4722);
or U4916 (N_4916,N_4708,N_4669);
xnor U4917 (N_4917,N_4677,N_4695);
or U4918 (N_4918,N_4680,N_4609);
or U4919 (N_4919,N_4724,N_4760);
xnor U4920 (N_4920,N_4678,N_4644);
nand U4921 (N_4921,N_4672,N_4692);
nor U4922 (N_4922,N_4783,N_4709);
xor U4923 (N_4923,N_4616,N_4787);
nand U4924 (N_4924,N_4671,N_4767);
nand U4925 (N_4925,N_4650,N_4798);
and U4926 (N_4926,N_4663,N_4743);
nor U4927 (N_4927,N_4745,N_4678);
or U4928 (N_4928,N_4701,N_4666);
nand U4929 (N_4929,N_4756,N_4634);
nand U4930 (N_4930,N_4714,N_4781);
or U4931 (N_4931,N_4796,N_4746);
nand U4932 (N_4932,N_4738,N_4633);
nand U4933 (N_4933,N_4691,N_4674);
and U4934 (N_4934,N_4780,N_4712);
xor U4935 (N_4935,N_4704,N_4743);
nand U4936 (N_4936,N_4606,N_4732);
nand U4937 (N_4937,N_4780,N_4607);
or U4938 (N_4938,N_4790,N_4778);
nor U4939 (N_4939,N_4758,N_4679);
xnor U4940 (N_4940,N_4724,N_4674);
or U4941 (N_4941,N_4740,N_4766);
or U4942 (N_4942,N_4647,N_4690);
and U4943 (N_4943,N_4713,N_4649);
or U4944 (N_4944,N_4628,N_4747);
and U4945 (N_4945,N_4610,N_4672);
xnor U4946 (N_4946,N_4647,N_4630);
nor U4947 (N_4947,N_4689,N_4721);
and U4948 (N_4948,N_4752,N_4724);
and U4949 (N_4949,N_4724,N_4658);
nor U4950 (N_4950,N_4637,N_4648);
nor U4951 (N_4951,N_4796,N_4641);
nand U4952 (N_4952,N_4651,N_4758);
or U4953 (N_4953,N_4720,N_4698);
and U4954 (N_4954,N_4612,N_4719);
xnor U4955 (N_4955,N_4796,N_4729);
and U4956 (N_4956,N_4641,N_4640);
or U4957 (N_4957,N_4631,N_4775);
nor U4958 (N_4958,N_4616,N_4660);
nor U4959 (N_4959,N_4789,N_4610);
nor U4960 (N_4960,N_4773,N_4695);
xnor U4961 (N_4961,N_4660,N_4702);
or U4962 (N_4962,N_4604,N_4631);
nand U4963 (N_4963,N_4626,N_4680);
and U4964 (N_4964,N_4707,N_4696);
xnor U4965 (N_4965,N_4752,N_4618);
nand U4966 (N_4966,N_4735,N_4760);
and U4967 (N_4967,N_4730,N_4609);
xnor U4968 (N_4968,N_4754,N_4798);
and U4969 (N_4969,N_4668,N_4724);
nand U4970 (N_4970,N_4611,N_4706);
or U4971 (N_4971,N_4643,N_4701);
or U4972 (N_4972,N_4696,N_4725);
nand U4973 (N_4973,N_4650,N_4662);
xor U4974 (N_4974,N_4712,N_4666);
or U4975 (N_4975,N_4765,N_4652);
xnor U4976 (N_4976,N_4775,N_4708);
nand U4977 (N_4977,N_4781,N_4793);
and U4978 (N_4978,N_4735,N_4736);
or U4979 (N_4979,N_4646,N_4632);
or U4980 (N_4980,N_4706,N_4609);
nand U4981 (N_4981,N_4656,N_4621);
and U4982 (N_4982,N_4622,N_4698);
nand U4983 (N_4983,N_4794,N_4640);
nand U4984 (N_4984,N_4775,N_4742);
xor U4985 (N_4985,N_4744,N_4749);
or U4986 (N_4986,N_4711,N_4626);
and U4987 (N_4987,N_4624,N_4708);
nor U4988 (N_4988,N_4667,N_4760);
and U4989 (N_4989,N_4721,N_4797);
and U4990 (N_4990,N_4776,N_4736);
nor U4991 (N_4991,N_4603,N_4629);
and U4992 (N_4992,N_4786,N_4623);
and U4993 (N_4993,N_4682,N_4651);
and U4994 (N_4994,N_4619,N_4754);
or U4995 (N_4995,N_4684,N_4632);
xnor U4996 (N_4996,N_4600,N_4793);
xor U4997 (N_4997,N_4643,N_4610);
nand U4998 (N_4998,N_4700,N_4654);
nand U4999 (N_4999,N_4691,N_4791);
nor UO_0 (O_0,N_4809,N_4846);
nor UO_1 (O_1,N_4975,N_4909);
nand UO_2 (O_2,N_4920,N_4801);
xnor UO_3 (O_3,N_4873,N_4845);
or UO_4 (O_4,N_4848,N_4800);
nor UO_5 (O_5,N_4977,N_4824);
nand UO_6 (O_6,N_4966,N_4924);
nor UO_7 (O_7,N_4961,N_4970);
nor UO_8 (O_8,N_4830,N_4905);
or UO_9 (O_9,N_4804,N_4821);
and UO_10 (O_10,N_4834,N_4802);
nor UO_11 (O_11,N_4982,N_4957);
nand UO_12 (O_12,N_4990,N_4911);
nor UO_13 (O_13,N_4843,N_4988);
or UO_14 (O_14,N_4936,N_4926);
xor UO_15 (O_15,N_4803,N_4892);
or UO_16 (O_16,N_4906,N_4995);
and UO_17 (O_17,N_4899,N_4847);
nand UO_18 (O_18,N_4851,N_4827);
nor UO_19 (O_19,N_4856,N_4948);
nor UO_20 (O_20,N_4935,N_4812);
and UO_21 (O_21,N_4974,N_4922);
xnor UO_22 (O_22,N_4872,N_4989);
nand UO_23 (O_23,N_4839,N_4853);
nor UO_24 (O_24,N_4959,N_4807);
and UO_25 (O_25,N_4937,N_4875);
xor UO_26 (O_26,N_4844,N_4954);
nand UO_27 (O_27,N_4805,N_4903);
and UO_28 (O_28,N_4900,N_4863);
nand UO_29 (O_29,N_4823,N_4910);
nor UO_30 (O_30,N_4897,N_4893);
and UO_31 (O_31,N_4815,N_4820);
nand UO_32 (O_32,N_4929,N_4985);
and UO_33 (O_33,N_4945,N_4983);
or UO_34 (O_34,N_4904,N_4946);
nand UO_35 (O_35,N_4965,N_4874);
and UO_36 (O_36,N_4831,N_4956);
xor UO_37 (O_37,N_4934,N_4928);
nand UO_38 (O_38,N_4958,N_4953);
nand UO_39 (O_39,N_4923,N_4866);
nor UO_40 (O_40,N_4978,N_4986);
or UO_41 (O_41,N_4916,N_4979);
or UO_42 (O_42,N_4814,N_4967);
or UO_43 (O_43,N_4890,N_4896);
nor UO_44 (O_44,N_4898,N_4984);
nand UO_45 (O_45,N_4850,N_4940);
xor UO_46 (O_46,N_4817,N_4855);
nand UO_47 (O_47,N_4968,N_4969);
nor UO_48 (O_48,N_4955,N_4943);
xnor UO_49 (O_49,N_4819,N_4894);
nor UO_50 (O_50,N_4907,N_4876);
and UO_51 (O_51,N_4932,N_4832);
nor UO_52 (O_52,N_4949,N_4895);
or UO_53 (O_53,N_4852,N_4862);
and UO_54 (O_54,N_4919,N_4902);
nor UO_55 (O_55,N_4888,N_4933);
nor UO_56 (O_56,N_4828,N_4854);
or UO_57 (O_57,N_4939,N_4891);
nand UO_58 (O_58,N_4994,N_4861);
nor UO_59 (O_59,N_4806,N_4942);
xnor UO_60 (O_60,N_4822,N_4837);
nand UO_61 (O_61,N_4964,N_4882);
nor UO_62 (O_62,N_4921,N_4841);
nor UO_63 (O_63,N_4878,N_4879);
or UO_64 (O_64,N_4950,N_4973);
and UO_65 (O_65,N_4849,N_4870);
nor UO_66 (O_66,N_4880,N_4829);
nor UO_67 (O_67,N_4996,N_4810);
or UO_68 (O_68,N_4960,N_4992);
nor UO_69 (O_69,N_4885,N_4998);
or UO_70 (O_70,N_4884,N_4877);
nor UO_71 (O_71,N_4840,N_4836);
nand UO_72 (O_72,N_4811,N_4925);
nor UO_73 (O_73,N_4947,N_4980);
or UO_74 (O_74,N_4963,N_4871);
nand UO_75 (O_75,N_4842,N_4981);
nor UO_76 (O_76,N_4859,N_4883);
xnor UO_77 (O_77,N_4869,N_4864);
nor UO_78 (O_78,N_4833,N_4901);
or UO_79 (O_79,N_4918,N_4987);
xor UO_80 (O_80,N_4818,N_4993);
nand UO_81 (O_81,N_4991,N_4913);
or UO_82 (O_82,N_4914,N_4997);
nor UO_83 (O_83,N_4972,N_4952);
and UO_84 (O_84,N_4808,N_4912);
and UO_85 (O_85,N_4915,N_4944);
and UO_86 (O_86,N_4962,N_4865);
xor UO_87 (O_87,N_4917,N_4858);
nand UO_88 (O_88,N_4908,N_4889);
or UO_89 (O_89,N_4931,N_4927);
nor UO_90 (O_90,N_4816,N_4941);
nor UO_91 (O_91,N_4825,N_4881);
xor UO_92 (O_92,N_4835,N_4887);
and UO_93 (O_93,N_4860,N_4868);
or UO_94 (O_94,N_4813,N_4976);
xnor UO_95 (O_95,N_4951,N_4826);
or UO_96 (O_96,N_4838,N_4857);
or UO_97 (O_97,N_4930,N_4971);
nor UO_98 (O_98,N_4999,N_4867);
and UO_99 (O_99,N_4886,N_4938);
xnor UO_100 (O_100,N_4920,N_4863);
or UO_101 (O_101,N_4979,N_4874);
nand UO_102 (O_102,N_4962,N_4905);
xnor UO_103 (O_103,N_4852,N_4991);
nor UO_104 (O_104,N_4915,N_4969);
and UO_105 (O_105,N_4933,N_4951);
nand UO_106 (O_106,N_4808,N_4898);
and UO_107 (O_107,N_4885,N_4805);
and UO_108 (O_108,N_4953,N_4900);
nand UO_109 (O_109,N_4863,N_4967);
xnor UO_110 (O_110,N_4873,N_4941);
xnor UO_111 (O_111,N_4839,N_4885);
nor UO_112 (O_112,N_4978,N_4806);
nand UO_113 (O_113,N_4939,N_4856);
and UO_114 (O_114,N_4813,N_4847);
or UO_115 (O_115,N_4985,N_4979);
nand UO_116 (O_116,N_4810,N_4972);
nor UO_117 (O_117,N_4954,N_4851);
nand UO_118 (O_118,N_4898,N_4867);
nor UO_119 (O_119,N_4842,N_4913);
or UO_120 (O_120,N_4805,N_4921);
or UO_121 (O_121,N_4866,N_4946);
nor UO_122 (O_122,N_4921,N_4935);
nor UO_123 (O_123,N_4963,N_4897);
xor UO_124 (O_124,N_4857,N_4832);
nor UO_125 (O_125,N_4864,N_4804);
and UO_126 (O_126,N_4809,N_4944);
nand UO_127 (O_127,N_4901,N_4845);
nand UO_128 (O_128,N_4902,N_4803);
nand UO_129 (O_129,N_4975,N_4940);
or UO_130 (O_130,N_4895,N_4992);
and UO_131 (O_131,N_4853,N_4995);
nand UO_132 (O_132,N_4821,N_4986);
and UO_133 (O_133,N_4999,N_4831);
or UO_134 (O_134,N_4940,N_4813);
nor UO_135 (O_135,N_4993,N_4822);
nand UO_136 (O_136,N_4948,N_4944);
and UO_137 (O_137,N_4941,N_4987);
xnor UO_138 (O_138,N_4999,N_4886);
nor UO_139 (O_139,N_4982,N_4942);
nor UO_140 (O_140,N_4831,N_4884);
and UO_141 (O_141,N_4898,N_4902);
xnor UO_142 (O_142,N_4962,N_4834);
nand UO_143 (O_143,N_4884,N_4961);
and UO_144 (O_144,N_4895,N_4987);
or UO_145 (O_145,N_4830,N_4914);
nand UO_146 (O_146,N_4934,N_4994);
or UO_147 (O_147,N_4831,N_4899);
and UO_148 (O_148,N_4853,N_4939);
or UO_149 (O_149,N_4940,N_4837);
nor UO_150 (O_150,N_4903,N_4930);
and UO_151 (O_151,N_4854,N_4901);
nand UO_152 (O_152,N_4996,N_4813);
and UO_153 (O_153,N_4829,N_4927);
or UO_154 (O_154,N_4973,N_4841);
nand UO_155 (O_155,N_4806,N_4981);
or UO_156 (O_156,N_4969,N_4897);
nor UO_157 (O_157,N_4960,N_4985);
nand UO_158 (O_158,N_4913,N_4823);
nor UO_159 (O_159,N_4937,N_4990);
and UO_160 (O_160,N_4934,N_4957);
nand UO_161 (O_161,N_4884,N_4829);
or UO_162 (O_162,N_4893,N_4919);
and UO_163 (O_163,N_4801,N_4921);
and UO_164 (O_164,N_4889,N_4859);
nand UO_165 (O_165,N_4973,N_4869);
and UO_166 (O_166,N_4866,N_4957);
xor UO_167 (O_167,N_4966,N_4800);
and UO_168 (O_168,N_4934,N_4808);
or UO_169 (O_169,N_4938,N_4906);
and UO_170 (O_170,N_4981,N_4932);
or UO_171 (O_171,N_4914,N_4976);
xor UO_172 (O_172,N_4965,N_4966);
or UO_173 (O_173,N_4960,N_4944);
nand UO_174 (O_174,N_4886,N_4826);
or UO_175 (O_175,N_4937,N_4973);
or UO_176 (O_176,N_4862,N_4847);
nand UO_177 (O_177,N_4853,N_4874);
and UO_178 (O_178,N_4875,N_4837);
or UO_179 (O_179,N_4890,N_4958);
nor UO_180 (O_180,N_4921,N_4908);
and UO_181 (O_181,N_4917,N_4822);
or UO_182 (O_182,N_4855,N_4991);
or UO_183 (O_183,N_4863,N_4931);
or UO_184 (O_184,N_4878,N_4873);
or UO_185 (O_185,N_4964,N_4801);
nor UO_186 (O_186,N_4821,N_4963);
nor UO_187 (O_187,N_4858,N_4910);
nor UO_188 (O_188,N_4836,N_4801);
or UO_189 (O_189,N_4989,N_4994);
and UO_190 (O_190,N_4817,N_4949);
nor UO_191 (O_191,N_4944,N_4911);
or UO_192 (O_192,N_4971,N_4825);
nor UO_193 (O_193,N_4964,N_4996);
and UO_194 (O_194,N_4946,N_4814);
or UO_195 (O_195,N_4935,N_4946);
nor UO_196 (O_196,N_4891,N_4989);
nand UO_197 (O_197,N_4806,N_4802);
nand UO_198 (O_198,N_4801,N_4946);
and UO_199 (O_199,N_4989,N_4807);
nor UO_200 (O_200,N_4820,N_4875);
nor UO_201 (O_201,N_4940,N_4832);
or UO_202 (O_202,N_4960,N_4840);
or UO_203 (O_203,N_4969,N_4916);
or UO_204 (O_204,N_4932,N_4860);
nor UO_205 (O_205,N_4869,N_4959);
nor UO_206 (O_206,N_4903,N_4978);
nand UO_207 (O_207,N_4828,N_4836);
nor UO_208 (O_208,N_4929,N_4884);
xor UO_209 (O_209,N_4944,N_4801);
nand UO_210 (O_210,N_4879,N_4864);
or UO_211 (O_211,N_4802,N_4972);
or UO_212 (O_212,N_4947,N_4938);
nand UO_213 (O_213,N_4838,N_4846);
and UO_214 (O_214,N_4932,N_4878);
or UO_215 (O_215,N_4868,N_4850);
nor UO_216 (O_216,N_4962,N_4863);
xnor UO_217 (O_217,N_4820,N_4823);
and UO_218 (O_218,N_4898,N_4829);
nor UO_219 (O_219,N_4859,N_4813);
and UO_220 (O_220,N_4926,N_4851);
nor UO_221 (O_221,N_4958,N_4803);
and UO_222 (O_222,N_4936,N_4960);
and UO_223 (O_223,N_4808,N_4899);
nor UO_224 (O_224,N_4903,N_4979);
nor UO_225 (O_225,N_4910,N_4816);
nand UO_226 (O_226,N_4850,N_4914);
nand UO_227 (O_227,N_4981,N_4970);
xnor UO_228 (O_228,N_4813,N_4871);
nand UO_229 (O_229,N_4837,N_4953);
nand UO_230 (O_230,N_4837,N_4905);
nand UO_231 (O_231,N_4810,N_4924);
nand UO_232 (O_232,N_4893,N_4821);
and UO_233 (O_233,N_4990,N_4993);
or UO_234 (O_234,N_4925,N_4913);
and UO_235 (O_235,N_4926,N_4862);
xnor UO_236 (O_236,N_4892,N_4915);
nor UO_237 (O_237,N_4817,N_4965);
nand UO_238 (O_238,N_4828,N_4801);
nand UO_239 (O_239,N_4823,N_4936);
and UO_240 (O_240,N_4852,N_4951);
nor UO_241 (O_241,N_4885,N_4891);
nor UO_242 (O_242,N_4932,N_4852);
and UO_243 (O_243,N_4915,N_4851);
nand UO_244 (O_244,N_4949,N_4969);
nor UO_245 (O_245,N_4830,N_4817);
or UO_246 (O_246,N_4800,N_4851);
or UO_247 (O_247,N_4946,N_4927);
nor UO_248 (O_248,N_4894,N_4906);
and UO_249 (O_249,N_4825,N_4993);
or UO_250 (O_250,N_4878,N_4936);
xnor UO_251 (O_251,N_4980,N_4884);
or UO_252 (O_252,N_4838,N_4965);
nor UO_253 (O_253,N_4885,N_4830);
or UO_254 (O_254,N_4886,N_4812);
xnor UO_255 (O_255,N_4983,N_4978);
nand UO_256 (O_256,N_4826,N_4978);
nor UO_257 (O_257,N_4941,N_4914);
nor UO_258 (O_258,N_4981,N_4839);
nor UO_259 (O_259,N_4847,N_4909);
and UO_260 (O_260,N_4894,N_4987);
or UO_261 (O_261,N_4861,N_4983);
and UO_262 (O_262,N_4872,N_4852);
or UO_263 (O_263,N_4956,N_4962);
nand UO_264 (O_264,N_4884,N_4921);
nor UO_265 (O_265,N_4869,N_4827);
nor UO_266 (O_266,N_4978,N_4841);
or UO_267 (O_267,N_4845,N_4869);
xor UO_268 (O_268,N_4858,N_4947);
nand UO_269 (O_269,N_4954,N_4847);
or UO_270 (O_270,N_4995,N_4807);
or UO_271 (O_271,N_4846,N_4862);
and UO_272 (O_272,N_4800,N_4948);
or UO_273 (O_273,N_4938,N_4890);
and UO_274 (O_274,N_4841,N_4864);
nor UO_275 (O_275,N_4838,N_4981);
and UO_276 (O_276,N_4950,N_4891);
nand UO_277 (O_277,N_4860,N_4884);
and UO_278 (O_278,N_4904,N_4825);
or UO_279 (O_279,N_4880,N_4921);
or UO_280 (O_280,N_4896,N_4826);
nor UO_281 (O_281,N_4894,N_4958);
nand UO_282 (O_282,N_4902,N_4850);
and UO_283 (O_283,N_4845,N_4913);
or UO_284 (O_284,N_4946,N_4943);
nor UO_285 (O_285,N_4808,N_4856);
and UO_286 (O_286,N_4963,N_4832);
nor UO_287 (O_287,N_4917,N_4834);
and UO_288 (O_288,N_4827,N_4914);
and UO_289 (O_289,N_4800,N_4816);
or UO_290 (O_290,N_4877,N_4975);
or UO_291 (O_291,N_4896,N_4800);
or UO_292 (O_292,N_4830,N_4954);
nor UO_293 (O_293,N_4811,N_4906);
nand UO_294 (O_294,N_4905,N_4835);
or UO_295 (O_295,N_4939,N_4937);
xnor UO_296 (O_296,N_4955,N_4853);
and UO_297 (O_297,N_4866,N_4837);
nor UO_298 (O_298,N_4895,N_4859);
or UO_299 (O_299,N_4928,N_4952);
nand UO_300 (O_300,N_4930,N_4893);
or UO_301 (O_301,N_4912,N_4830);
or UO_302 (O_302,N_4967,N_4830);
nor UO_303 (O_303,N_4804,N_4994);
or UO_304 (O_304,N_4804,N_4805);
or UO_305 (O_305,N_4893,N_4815);
nand UO_306 (O_306,N_4983,N_4801);
nand UO_307 (O_307,N_4914,N_4828);
and UO_308 (O_308,N_4933,N_4862);
nor UO_309 (O_309,N_4956,N_4963);
and UO_310 (O_310,N_4929,N_4940);
nor UO_311 (O_311,N_4823,N_4952);
nand UO_312 (O_312,N_4971,N_4894);
or UO_313 (O_313,N_4810,N_4817);
or UO_314 (O_314,N_4813,N_4858);
nand UO_315 (O_315,N_4934,N_4949);
and UO_316 (O_316,N_4988,N_4934);
nand UO_317 (O_317,N_4811,N_4800);
nor UO_318 (O_318,N_4897,N_4949);
nand UO_319 (O_319,N_4939,N_4995);
nand UO_320 (O_320,N_4976,N_4895);
nand UO_321 (O_321,N_4983,N_4952);
or UO_322 (O_322,N_4893,N_4994);
nand UO_323 (O_323,N_4933,N_4962);
and UO_324 (O_324,N_4955,N_4970);
and UO_325 (O_325,N_4806,N_4850);
nand UO_326 (O_326,N_4855,N_4843);
nand UO_327 (O_327,N_4878,N_4937);
and UO_328 (O_328,N_4825,N_4959);
xnor UO_329 (O_329,N_4877,N_4863);
nand UO_330 (O_330,N_4965,N_4963);
xor UO_331 (O_331,N_4817,N_4851);
nor UO_332 (O_332,N_4839,N_4959);
nand UO_333 (O_333,N_4810,N_4848);
or UO_334 (O_334,N_4898,N_4985);
and UO_335 (O_335,N_4860,N_4998);
nand UO_336 (O_336,N_4827,N_4957);
and UO_337 (O_337,N_4921,N_4960);
nor UO_338 (O_338,N_4990,N_4864);
or UO_339 (O_339,N_4937,N_4999);
and UO_340 (O_340,N_4814,N_4857);
xor UO_341 (O_341,N_4890,N_4832);
nand UO_342 (O_342,N_4875,N_4919);
nor UO_343 (O_343,N_4942,N_4986);
nand UO_344 (O_344,N_4962,N_4975);
xnor UO_345 (O_345,N_4987,N_4965);
or UO_346 (O_346,N_4880,N_4961);
nor UO_347 (O_347,N_4867,N_4931);
nor UO_348 (O_348,N_4812,N_4915);
and UO_349 (O_349,N_4845,N_4978);
nor UO_350 (O_350,N_4966,N_4972);
and UO_351 (O_351,N_4835,N_4870);
nand UO_352 (O_352,N_4821,N_4855);
or UO_353 (O_353,N_4910,N_4865);
nand UO_354 (O_354,N_4831,N_4937);
nor UO_355 (O_355,N_4840,N_4807);
or UO_356 (O_356,N_4981,N_4957);
xor UO_357 (O_357,N_4856,N_4817);
nor UO_358 (O_358,N_4946,N_4872);
nand UO_359 (O_359,N_4928,N_4986);
nand UO_360 (O_360,N_4978,N_4980);
or UO_361 (O_361,N_4944,N_4946);
and UO_362 (O_362,N_4808,N_4988);
or UO_363 (O_363,N_4960,N_4973);
nor UO_364 (O_364,N_4949,N_4955);
xnor UO_365 (O_365,N_4950,N_4932);
or UO_366 (O_366,N_4880,N_4932);
or UO_367 (O_367,N_4980,N_4810);
xnor UO_368 (O_368,N_4819,N_4973);
xor UO_369 (O_369,N_4988,N_4834);
nand UO_370 (O_370,N_4897,N_4800);
or UO_371 (O_371,N_4958,N_4818);
or UO_372 (O_372,N_4927,N_4951);
nor UO_373 (O_373,N_4858,N_4856);
nand UO_374 (O_374,N_4961,N_4857);
and UO_375 (O_375,N_4801,N_4929);
xor UO_376 (O_376,N_4929,N_4958);
and UO_377 (O_377,N_4825,N_4990);
and UO_378 (O_378,N_4916,N_4863);
nor UO_379 (O_379,N_4965,N_4800);
xnor UO_380 (O_380,N_4948,N_4896);
and UO_381 (O_381,N_4841,N_4924);
and UO_382 (O_382,N_4840,N_4831);
nand UO_383 (O_383,N_4905,N_4865);
nor UO_384 (O_384,N_4974,N_4811);
or UO_385 (O_385,N_4995,N_4814);
nand UO_386 (O_386,N_4838,N_4852);
or UO_387 (O_387,N_4829,N_4908);
nand UO_388 (O_388,N_4811,N_4975);
xnor UO_389 (O_389,N_4984,N_4899);
xor UO_390 (O_390,N_4855,N_4932);
nand UO_391 (O_391,N_4918,N_4956);
xnor UO_392 (O_392,N_4881,N_4912);
and UO_393 (O_393,N_4817,N_4880);
xnor UO_394 (O_394,N_4924,N_4852);
nor UO_395 (O_395,N_4937,N_4817);
xor UO_396 (O_396,N_4837,N_4986);
or UO_397 (O_397,N_4802,N_4840);
nand UO_398 (O_398,N_4837,N_4810);
nand UO_399 (O_399,N_4833,N_4988);
nor UO_400 (O_400,N_4995,N_4810);
nand UO_401 (O_401,N_4872,N_4996);
nand UO_402 (O_402,N_4838,N_4893);
xor UO_403 (O_403,N_4962,N_4861);
and UO_404 (O_404,N_4935,N_4817);
or UO_405 (O_405,N_4893,N_4927);
xor UO_406 (O_406,N_4915,N_4912);
nand UO_407 (O_407,N_4919,N_4843);
and UO_408 (O_408,N_4902,N_4961);
or UO_409 (O_409,N_4951,N_4925);
or UO_410 (O_410,N_4950,N_4942);
and UO_411 (O_411,N_4902,N_4893);
and UO_412 (O_412,N_4865,N_4833);
nand UO_413 (O_413,N_4892,N_4980);
xor UO_414 (O_414,N_4954,N_4960);
or UO_415 (O_415,N_4931,N_4918);
nand UO_416 (O_416,N_4963,N_4852);
nand UO_417 (O_417,N_4934,N_4974);
nor UO_418 (O_418,N_4999,N_4927);
xnor UO_419 (O_419,N_4842,N_4898);
and UO_420 (O_420,N_4959,N_4832);
xor UO_421 (O_421,N_4924,N_4802);
or UO_422 (O_422,N_4871,N_4938);
nor UO_423 (O_423,N_4913,N_4889);
and UO_424 (O_424,N_4805,N_4978);
or UO_425 (O_425,N_4847,N_4940);
nand UO_426 (O_426,N_4900,N_4875);
and UO_427 (O_427,N_4986,N_4859);
or UO_428 (O_428,N_4976,N_4940);
nor UO_429 (O_429,N_4974,N_4820);
or UO_430 (O_430,N_4950,N_4955);
nor UO_431 (O_431,N_4976,N_4999);
nand UO_432 (O_432,N_4908,N_4890);
nor UO_433 (O_433,N_4949,N_4930);
nand UO_434 (O_434,N_4846,N_4836);
and UO_435 (O_435,N_4937,N_4936);
or UO_436 (O_436,N_4939,N_4864);
nand UO_437 (O_437,N_4975,N_4813);
nor UO_438 (O_438,N_4934,N_4892);
nand UO_439 (O_439,N_4897,N_4877);
nand UO_440 (O_440,N_4851,N_4939);
nor UO_441 (O_441,N_4870,N_4900);
nor UO_442 (O_442,N_4990,N_4805);
and UO_443 (O_443,N_4924,N_4938);
xor UO_444 (O_444,N_4989,N_4874);
nand UO_445 (O_445,N_4889,N_4855);
nand UO_446 (O_446,N_4905,N_4967);
nor UO_447 (O_447,N_4853,N_4933);
nand UO_448 (O_448,N_4865,N_4841);
and UO_449 (O_449,N_4893,N_4963);
or UO_450 (O_450,N_4927,N_4844);
nand UO_451 (O_451,N_4811,N_4805);
nand UO_452 (O_452,N_4857,N_4919);
nor UO_453 (O_453,N_4932,N_4801);
nand UO_454 (O_454,N_4921,N_4904);
nand UO_455 (O_455,N_4816,N_4936);
nor UO_456 (O_456,N_4907,N_4951);
nor UO_457 (O_457,N_4821,N_4988);
nand UO_458 (O_458,N_4839,N_4999);
xor UO_459 (O_459,N_4879,N_4900);
or UO_460 (O_460,N_4920,N_4948);
xnor UO_461 (O_461,N_4878,N_4823);
and UO_462 (O_462,N_4930,N_4927);
nand UO_463 (O_463,N_4971,N_4830);
and UO_464 (O_464,N_4854,N_4895);
nor UO_465 (O_465,N_4800,N_4973);
or UO_466 (O_466,N_4965,N_4833);
nor UO_467 (O_467,N_4969,N_4808);
nand UO_468 (O_468,N_4832,N_4826);
nor UO_469 (O_469,N_4933,N_4894);
nor UO_470 (O_470,N_4949,N_4914);
nor UO_471 (O_471,N_4801,N_4814);
nand UO_472 (O_472,N_4858,N_4807);
nand UO_473 (O_473,N_4947,N_4985);
or UO_474 (O_474,N_4884,N_4915);
nor UO_475 (O_475,N_4977,N_4913);
nand UO_476 (O_476,N_4807,N_4872);
nand UO_477 (O_477,N_4821,N_4998);
nand UO_478 (O_478,N_4968,N_4984);
nand UO_479 (O_479,N_4804,N_4860);
or UO_480 (O_480,N_4850,N_4913);
or UO_481 (O_481,N_4978,N_4873);
nor UO_482 (O_482,N_4960,N_4958);
or UO_483 (O_483,N_4841,N_4908);
nor UO_484 (O_484,N_4969,N_4933);
xnor UO_485 (O_485,N_4830,N_4868);
and UO_486 (O_486,N_4890,N_4839);
or UO_487 (O_487,N_4972,N_4826);
nand UO_488 (O_488,N_4937,N_4845);
or UO_489 (O_489,N_4997,N_4897);
nor UO_490 (O_490,N_4903,N_4996);
and UO_491 (O_491,N_4855,N_4974);
nor UO_492 (O_492,N_4836,N_4849);
nor UO_493 (O_493,N_4842,N_4861);
and UO_494 (O_494,N_4964,N_4975);
nor UO_495 (O_495,N_4845,N_4860);
nand UO_496 (O_496,N_4961,N_4939);
nor UO_497 (O_497,N_4805,N_4897);
nor UO_498 (O_498,N_4851,N_4964);
nand UO_499 (O_499,N_4868,N_4874);
and UO_500 (O_500,N_4815,N_4857);
nand UO_501 (O_501,N_4944,N_4990);
and UO_502 (O_502,N_4939,N_4802);
nand UO_503 (O_503,N_4909,N_4910);
or UO_504 (O_504,N_4822,N_4984);
nand UO_505 (O_505,N_4915,N_4869);
xor UO_506 (O_506,N_4959,N_4820);
nand UO_507 (O_507,N_4876,N_4940);
and UO_508 (O_508,N_4996,N_4907);
or UO_509 (O_509,N_4965,N_4811);
xor UO_510 (O_510,N_4911,N_4939);
nand UO_511 (O_511,N_4915,N_4983);
xor UO_512 (O_512,N_4851,N_4886);
or UO_513 (O_513,N_4822,N_4909);
nand UO_514 (O_514,N_4984,N_4936);
nand UO_515 (O_515,N_4919,N_4908);
and UO_516 (O_516,N_4992,N_4877);
and UO_517 (O_517,N_4949,N_4933);
nor UO_518 (O_518,N_4935,N_4823);
xnor UO_519 (O_519,N_4873,N_4895);
or UO_520 (O_520,N_4933,N_4891);
and UO_521 (O_521,N_4909,N_4854);
and UO_522 (O_522,N_4975,N_4968);
and UO_523 (O_523,N_4866,N_4847);
nand UO_524 (O_524,N_4844,N_4970);
or UO_525 (O_525,N_4858,N_4855);
nand UO_526 (O_526,N_4825,N_4988);
or UO_527 (O_527,N_4822,N_4850);
or UO_528 (O_528,N_4926,N_4917);
and UO_529 (O_529,N_4951,N_4855);
nand UO_530 (O_530,N_4800,N_4953);
xnor UO_531 (O_531,N_4818,N_4981);
nor UO_532 (O_532,N_4901,N_4992);
nand UO_533 (O_533,N_4877,N_4820);
nand UO_534 (O_534,N_4987,N_4887);
xnor UO_535 (O_535,N_4845,N_4885);
xnor UO_536 (O_536,N_4831,N_4909);
and UO_537 (O_537,N_4893,N_4988);
and UO_538 (O_538,N_4876,N_4835);
xnor UO_539 (O_539,N_4990,N_4838);
nor UO_540 (O_540,N_4819,N_4920);
nor UO_541 (O_541,N_4906,N_4924);
nand UO_542 (O_542,N_4839,N_4969);
and UO_543 (O_543,N_4802,N_4996);
or UO_544 (O_544,N_4887,N_4978);
and UO_545 (O_545,N_4838,N_4902);
or UO_546 (O_546,N_4848,N_4921);
nor UO_547 (O_547,N_4814,N_4849);
and UO_548 (O_548,N_4892,N_4966);
or UO_549 (O_549,N_4971,N_4935);
or UO_550 (O_550,N_4817,N_4903);
or UO_551 (O_551,N_4837,N_4913);
or UO_552 (O_552,N_4999,N_4872);
nor UO_553 (O_553,N_4971,N_4832);
and UO_554 (O_554,N_4817,N_4902);
and UO_555 (O_555,N_4980,N_4985);
nand UO_556 (O_556,N_4960,N_4924);
nand UO_557 (O_557,N_4966,N_4887);
nor UO_558 (O_558,N_4828,N_4858);
or UO_559 (O_559,N_4887,N_4884);
or UO_560 (O_560,N_4961,N_4973);
and UO_561 (O_561,N_4888,N_4852);
nand UO_562 (O_562,N_4978,N_4902);
xnor UO_563 (O_563,N_4868,N_4810);
and UO_564 (O_564,N_4848,N_4942);
or UO_565 (O_565,N_4918,N_4890);
xor UO_566 (O_566,N_4890,N_4833);
nor UO_567 (O_567,N_4826,N_4982);
xnor UO_568 (O_568,N_4904,N_4942);
and UO_569 (O_569,N_4951,N_4891);
xor UO_570 (O_570,N_4998,N_4995);
and UO_571 (O_571,N_4828,N_4944);
nor UO_572 (O_572,N_4966,N_4895);
and UO_573 (O_573,N_4845,N_4841);
xnor UO_574 (O_574,N_4882,N_4918);
and UO_575 (O_575,N_4863,N_4850);
and UO_576 (O_576,N_4945,N_4884);
nand UO_577 (O_577,N_4897,N_4845);
and UO_578 (O_578,N_4971,N_4856);
nand UO_579 (O_579,N_4924,N_4959);
nor UO_580 (O_580,N_4917,N_4985);
and UO_581 (O_581,N_4984,N_4918);
or UO_582 (O_582,N_4844,N_4981);
xnor UO_583 (O_583,N_4983,N_4804);
and UO_584 (O_584,N_4833,N_4804);
or UO_585 (O_585,N_4949,N_4864);
and UO_586 (O_586,N_4808,N_4930);
or UO_587 (O_587,N_4989,N_4976);
and UO_588 (O_588,N_4893,N_4951);
nor UO_589 (O_589,N_4824,N_4927);
or UO_590 (O_590,N_4837,N_4860);
and UO_591 (O_591,N_4946,N_4886);
and UO_592 (O_592,N_4958,N_4857);
and UO_593 (O_593,N_4909,N_4956);
or UO_594 (O_594,N_4905,N_4834);
nand UO_595 (O_595,N_4883,N_4994);
nand UO_596 (O_596,N_4896,N_4980);
nand UO_597 (O_597,N_4997,N_4892);
and UO_598 (O_598,N_4814,N_4890);
or UO_599 (O_599,N_4851,N_4970);
nor UO_600 (O_600,N_4897,N_4937);
xnor UO_601 (O_601,N_4952,N_4846);
xor UO_602 (O_602,N_4801,N_4841);
and UO_603 (O_603,N_4950,N_4964);
and UO_604 (O_604,N_4876,N_4981);
xnor UO_605 (O_605,N_4808,N_4838);
nor UO_606 (O_606,N_4831,N_4829);
nor UO_607 (O_607,N_4999,N_4962);
nor UO_608 (O_608,N_4912,N_4801);
nor UO_609 (O_609,N_4862,N_4920);
and UO_610 (O_610,N_4990,N_4896);
nor UO_611 (O_611,N_4989,N_4911);
nor UO_612 (O_612,N_4933,N_4983);
nor UO_613 (O_613,N_4924,N_4967);
nand UO_614 (O_614,N_4832,N_4838);
nand UO_615 (O_615,N_4803,N_4879);
or UO_616 (O_616,N_4884,N_4930);
or UO_617 (O_617,N_4888,N_4874);
nor UO_618 (O_618,N_4948,N_4858);
nand UO_619 (O_619,N_4909,N_4915);
and UO_620 (O_620,N_4889,N_4933);
or UO_621 (O_621,N_4815,N_4908);
nand UO_622 (O_622,N_4945,N_4922);
nor UO_623 (O_623,N_4816,N_4978);
nor UO_624 (O_624,N_4803,N_4801);
nor UO_625 (O_625,N_4942,N_4889);
or UO_626 (O_626,N_4888,N_4948);
nor UO_627 (O_627,N_4997,N_4980);
xor UO_628 (O_628,N_4985,N_4873);
nor UO_629 (O_629,N_4834,N_4833);
and UO_630 (O_630,N_4841,N_4811);
nor UO_631 (O_631,N_4846,N_4911);
or UO_632 (O_632,N_4892,N_4967);
and UO_633 (O_633,N_4862,N_4801);
nor UO_634 (O_634,N_4994,N_4817);
and UO_635 (O_635,N_4866,N_4857);
xnor UO_636 (O_636,N_4998,N_4834);
nand UO_637 (O_637,N_4837,N_4828);
xor UO_638 (O_638,N_4938,N_4850);
nand UO_639 (O_639,N_4853,N_4981);
and UO_640 (O_640,N_4818,N_4880);
or UO_641 (O_641,N_4978,N_4900);
nor UO_642 (O_642,N_4820,N_4819);
and UO_643 (O_643,N_4923,N_4963);
nor UO_644 (O_644,N_4851,N_4969);
or UO_645 (O_645,N_4878,N_4957);
nand UO_646 (O_646,N_4882,N_4868);
nand UO_647 (O_647,N_4923,N_4847);
nor UO_648 (O_648,N_4947,N_4862);
nand UO_649 (O_649,N_4949,N_4893);
nand UO_650 (O_650,N_4992,N_4998);
and UO_651 (O_651,N_4940,N_4970);
nor UO_652 (O_652,N_4875,N_4934);
nand UO_653 (O_653,N_4893,N_4912);
nor UO_654 (O_654,N_4975,N_4887);
nand UO_655 (O_655,N_4998,N_4862);
and UO_656 (O_656,N_4943,N_4924);
nor UO_657 (O_657,N_4954,N_4937);
or UO_658 (O_658,N_4983,N_4855);
or UO_659 (O_659,N_4924,N_4915);
or UO_660 (O_660,N_4947,N_4986);
and UO_661 (O_661,N_4860,N_4827);
xnor UO_662 (O_662,N_4921,N_4950);
xor UO_663 (O_663,N_4863,N_4812);
and UO_664 (O_664,N_4893,N_4801);
nor UO_665 (O_665,N_4948,N_4996);
and UO_666 (O_666,N_4967,N_4840);
nor UO_667 (O_667,N_4927,N_4834);
and UO_668 (O_668,N_4805,N_4932);
nor UO_669 (O_669,N_4851,N_4966);
xnor UO_670 (O_670,N_4963,N_4872);
nor UO_671 (O_671,N_4870,N_4830);
xnor UO_672 (O_672,N_4934,N_4891);
nor UO_673 (O_673,N_4807,N_4972);
nor UO_674 (O_674,N_4904,N_4917);
nor UO_675 (O_675,N_4909,N_4994);
nor UO_676 (O_676,N_4941,N_4918);
and UO_677 (O_677,N_4890,N_4923);
xor UO_678 (O_678,N_4873,N_4858);
nor UO_679 (O_679,N_4952,N_4923);
nand UO_680 (O_680,N_4875,N_4871);
nand UO_681 (O_681,N_4895,N_4886);
nand UO_682 (O_682,N_4980,N_4953);
nor UO_683 (O_683,N_4856,N_4889);
and UO_684 (O_684,N_4864,N_4966);
xor UO_685 (O_685,N_4831,N_4972);
nor UO_686 (O_686,N_4944,N_4997);
nor UO_687 (O_687,N_4809,N_4843);
nor UO_688 (O_688,N_4963,N_4954);
or UO_689 (O_689,N_4894,N_4881);
or UO_690 (O_690,N_4927,N_4979);
nand UO_691 (O_691,N_4839,N_4806);
or UO_692 (O_692,N_4968,N_4878);
or UO_693 (O_693,N_4989,N_4850);
nand UO_694 (O_694,N_4977,N_4926);
nor UO_695 (O_695,N_4823,N_4840);
and UO_696 (O_696,N_4833,N_4842);
or UO_697 (O_697,N_4859,N_4871);
or UO_698 (O_698,N_4830,N_4946);
or UO_699 (O_699,N_4850,N_4803);
or UO_700 (O_700,N_4886,N_4990);
and UO_701 (O_701,N_4891,N_4984);
and UO_702 (O_702,N_4928,N_4958);
xor UO_703 (O_703,N_4935,N_4896);
or UO_704 (O_704,N_4876,N_4921);
or UO_705 (O_705,N_4968,N_4829);
or UO_706 (O_706,N_4927,N_4938);
or UO_707 (O_707,N_4945,N_4893);
and UO_708 (O_708,N_4831,N_4895);
or UO_709 (O_709,N_4918,N_4800);
or UO_710 (O_710,N_4876,N_4863);
nand UO_711 (O_711,N_4926,N_4871);
nor UO_712 (O_712,N_4973,N_4846);
and UO_713 (O_713,N_4979,N_4840);
and UO_714 (O_714,N_4920,N_4922);
or UO_715 (O_715,N_4886,N_4871);
and UO_716 (O_716,N_4970,N_4902);
nor UO_717 (O_717,N_4884,N_4847);
xnor UO_718 (O_718,N_4941,N_4980);
xnor UO_719 (O_719,N_4994,N_4981);
xnor UO_720 (O_720,N_4911,N_4960);
nor UO_721 (O_721,N_4984,N_4940);
nor UO_722 (O_722,N_4823,N_4948);
xnor UO_723 (O_723,N_4891,N_4872);
nand UO_724 (O_724,N_4921,N_4934);
nand UO_725 (O_725,N_4974,N_4931);
nand UO_726 (O_726,N_4989,N_4906);
nand UO_727 (O_727,N_4831,N_4978);
or UO_728 (O_728,N_4800,N_4880);
or UO_729 (O_729,N_4867,N_4957);
nor UO_730 (O_730,N_4883,N_4842);
xor UO_731 (O_731,N_4875,N_4938);
nor UO_732 (O_732,N_4911,N_4921);
and UO_733 (O_733,N_4994,N_4823);
nand UO_734 (O_734,N_4849,N_4919);
or UO_735 (O_735,N_4949,N_4945);
and UO_736 (O_736,N_4899,N_4958);
nand UO_737 (O_737,N_4850,N_4925);
xnor UO_738 (O_738,N_4804,N_4843);
nor UO_739 (O_739,N_4969,N_4979);
nor UO_740 (O_740,N_4839,N_4955);
nor UO_741 (O_741,N_4916,N_4805);
or UO_742 (O_742,N_4902,N_4878);
xnor UO_743 (O_743,N_4884,N_4973);
and UO_744 (O_744,N_4990,N_4936);
nand UO_745 (O_745,N_4907,N_4918);
nand UO_746 (O_746,N_4845,N_4894);
xor UO_747 (O_747,N_4836,N_4899);
xnor UO_748 (O_748,N_4856,N_4938);
xnor UO_749 (O_749,N_4954,N_4901);
and UO_750 (O_750,N_4860,N_4977);
nand UO_751 (O_751,N_4945,N_4989);
nor UO_752 (O_752,N_4841,N_4839);
or UO_753 (O_753,N_4912,N_4900);
nand UO_754 (O_754,N_4960,N_4913);
and UO_755 (O_755,N_4800,N_4964);
and UO_756 (O_756,N_4803,N_4948);
nand UO_757 (O_757,N_4823,N_4968);
or UO_758 (O_758,N_4954,N_4926);
nand UO_759 (O_759,N_4896,N_4925);
nand UO_760 (O_760,N_4959,N_4879);
and UO_761 (O_761,N_4890,N_4822);
and UO_762 (O_762,N_4860,N_4905);
nand UO_763 (O_763,N_4845,N_4966);
or UO_764 (O_764,N_4970,N_4870);
nor UO_765 (O_765,N_4878,N_4915);
or UO_766 (O_766,N_4944,N_4879);
nor UO_767 (O_767,N_4817,N_4929);
xnor UO_768 (O_768,N_4943,N_4870);
nand UO_769 (O_769,N_4955,N_4921);
nand UO_770 (O_770,N_4920,N_4829);
nor UO_771 (O_771,N_4954,N_4825);
or UO_772 (O_772,N_4909,N_4923);
nor UO_773 (O_773,N_4907,N_4860);
nand UO_774 (O_774,N_4922,N_4998);
nand UO_775 (O_775,N_4877,N_4913);
nor UO_776 (O_776,N_4958,N_4855);
or UO_777 (O_777,N_4969,N_4885);
nor UO_778 (O_778,N_4900,N_4926);
xnor UO_779 (O_779,N_4956,N_4864);
nor UO_780 (O_780,N_4833,N_4923);
and UO_781 (O_781,N_4954,N_4870);
or UO_782 (O_782,N_4942,N_4973);
nor UO_783 (O_783,N_4853,N_4958);
xor UO_784 (O_784,N_4829,N_4842);
or UO_785 (O_785,N_4983,N_4966);
or UO_786 (O_786,N_4976,N_4980);
nor UO_787 (O_787,N_4810,N_4935);
or UO_788 (O_788,N_4866,N_4984);
nor UO_789 (O_789,N_4891,N_4842);
and UO_790 (O_790,N_4822,N_4978);
nand UO_791 (O_791,N_4947,N_4809);
nor UO_792 (O_792,N_4856,N_4828);
nand UO_793 (O_793,N_4986,N_4828);
nand UO_794 (O_794,N_4929,N_4978);
nand UO_795 (O_795,N_4927,N_4909);
xor UO_796 (O_796,N_4889,N_4881);
or UO_797 (O_797,N_4838,N_4829);
nor UO_798 (O_798,N_4874,N_4811);
nor UO_799 (O_799,N_4961,N_4900);
nor UO_800 (O_800,N_4916,N_4834);
nand UO_801 (O_801,N_4822,N_4866);
nand UO_802 (O_802,N_4969,N_4928);
or UO_803 (O_803,N_4923,N_4951);
nand UO_804 (O_804,N_4951,N_4833);
and UO_805 (O_805,N_4995,N_4836);
nor UO_806 (O_806,N_4992,N_4825);
and UO_807 (O_807,N_4901,N_4936);
nand UO_808 (O_808,N_4876,N_4828);
nand UO_809 (O_809,N_4818,N_4895);
and UO_810 (O_810,N_4851,N_4836);
nand UO_811 (O_811,N_4842,N_4993);
nand UO_812 (O_812,N_4950,N_4828);
nor UO_813 (O_813,N_4997,N_4803);
nor UO_814 (O_814,N_4833,N_4891);
and UO_815 (O_815,N_4988,N_4872);
nand UO_816 (O_816,N_4971,N_4984);
nand UO_817 (O_817,N_4822,N_4908);
nand UO_818 (O_818,N_4801,N_4927);
and UO_819 (O_819,N_4924,N_4805);
and UO_820 (O_820,N_4873,N_4909);
or UO_821 (O_821,N_4878,N_4963);
and UO_822 (O_822,N_4854,N_4915);
nand UO_823 (O_823,N_4885,N_4817);
nor UO_824 (O_824,N_4836,N_4831);
or UO_825 (O_825,N_4933,N_4928);
nor UO_826 (O_826,N_4904,N_4853);
nand UO_827 (O_827,N_4867,N_4844);
xnor UO_828 (O_828,N_4811,N_4895);
nor UO_829 (O_829,N_4975,N_4991);
nand UO_830 (O_830,N_4978,N_4950);
nand UO_831 (O_831,N_4816,N_4962);
or UO_832 (O_832,N_4918,N_4883);
or UO_833 (O_833,N_4971,N_4972);
and UO_834 (O_834,N_4802,N_4938);
nor UO_835 (O_835,N_4857,N_4896);
and UO_836 (O_836,N_4861,N_4882);
nand UO_837 (O_837,N_4861,N_4816);
nand UO_838 (O_838,N_4857,N_4875);
nor UO_839 (O_839,N_4918,N_4857);
nor UO_840 (O_840,N_4962,N_4998);
and UO_841 (O_841,N_4976,N_4965);
nand UO_842 (O_842,N_4864,N_4892);
nor UO_843 (O_843,N_4879,N_4967);
nor UO_844 (O_844,N_4877,N_4867);
and UO_845 (O_845,N_4839,N_4931);
nor UO_846 (O_846,N_4897,N_4992);
and UO_847 (O_847,N_4968,N_4924);
nor UO_848 (O_848,N_4895,N_4833);
xnor UO_849 (O_849,N_4975,N_4872);
nand UO_850 (O_850,N_4854,N_4974);
nand UO_851 (O_851,N_4972,N_4984);
and UO_852 (O_852,N_4930,N_4825);
and UO_853 (O_853,N_4917,N_4832);
and UO_854 (O_854,N_4853,N_4822);
or UO_855 (O_855,N_4803,N_4838);
nor UO_856 (O_856,N_4921,N_4852);
nand UO_857 (O_857,N_4939,N_4827);
nand UO_858 (O_858,N_4836,N_4891);
nor UO_859 (O_859,N_4879,N_4991);
and UO_860 (O_860,N_4817,N_4837);
and UO_861 (O_861,N_4977,N_4849);
nor UO_862 (O_862,N_4914,N_4851);
and UO_863 (O_863,N_4990,N_4834);
or UO_864 (O_864,N_4946,N_4949);
and UO_865 (O_865,N_4982,N_4997);
and UO_866 (O_866,N_4923,N_4926);
nor UO_867 (O_867,N_4880,N_4925);
nor UO_868 (O_868,N_4931,N_4825);
nand UO_869 (O_869,N_4864,N_4919);
or UO_870 (O_870,N_4968,N_4897);
or UO_871 (O_871,N_4819,N_4989);
nand UO_872 (O_872,N_4962,N_4954);
and UO_873 (O_873,N_4953,N_4984);
or UO_874 (O_874,N_4920,N_4805);
nor UO_875 (O_875,N_4972,N_4951);
nor UO_876 (O_876,N_4903,N_4939);
nor UO_877 (O_877,N_4996,N_4808);
nand UO_878 (O_878,N_4932,N_4851);
xor UO_879 (O_879,N_4920,N_4825);
or UO_880 (O_880,N_4811,N_4837);
nor UO_881 (O_881,N_4926,N_4833);
or UO_882 (O_882,N_4913,N_4966);
nand UO_883 (O_883,N_4932,N_4814);
xor UO_884 (O_884,N_4970,N_4991);
nor UO_885 (O_885,N_4994,N_4919);
or UO_886 (O_886,N_4805,N_4895);
nand UO_887 (O_887,N_4803,N_4802);
nand UO_888 (O_888,N_4957,N_4910);
or UO_889 (O_889,N_4985,N_4829);
xor UO_890 (O_890,N_4856,N_4815);
or UO_891 (O_891,N_4972,N_4800);
nor UO_892 (O_892,N_4855,N_4995);
and UO_893 (O_893,N_4844,N_4895);
or UO_894 (O_894,N_4833,N_4838);
nor UO_895 (O_895,N_4964,N_4879);
nor UO_896 (O_896,N_4888,N_4946);
nor UO_897 (O_897,N_4815,N_4894);
nor UO_898 (O_898,N_4909,N_4834);
or UO_899 (O_899,N_4942,N_4838);
nand UO_900 (O_900,N_4905,N_4887);
and UO_901 (O_901,N_4881,N_4942);
and UO_902 (O_902,N_4997,N_4986);
nor UO_903 (O_903,N_4802,N_4947);
xnor UO_904 (O_904,N_4897,N_4853);
nand UO_905 (O_905,N_4835,N_4855);
and UO_906 (O_906,N_4816,N_4975);
nand UO_907 (O_907,N_4844,N_4854);
or UO_908 (O_908,N_4963,N_4876);
nand UO_909 (O_909,N_4962,N_4948);
nor UO_910 (O_910,N_4815,N_4810);
and UO_911 (O_911,N_4911,N_4816);
and UO_912 (O_912,N_4908,N_4896);
and UO_913 (O_913,N_4849,N_4958);
xor UO_914 (O_914,N_4832,N_4840);
and UO_915 (O_915,N_4828,N_4843);
xnor UO_916 (O_916,N_4840,N_4928);
nand UO_917 (O_917,N_4914,N_4895);
nand UO_918 (O_918,N_4907,N_4937);
nor UO_919 (O_919,N_4908,N_4904);
nor UO_920 (O_920,N_4872,N_4994);
nor UO_921 (O_921,N_4992,N_4891);
or UO_922 (O_922,N_4853,N_4920);
nand UO_923 (O_923,N_4922,N_4882);
nand UO_924 (O_924,N_4909,N_4979);
or UO_925 (O_925,N_4995,N_4985);
nand UO_926 (O_926,N_4906,N_4947);
nor UO_927 (O_927,N_4897,N_4966);
nor UO_928 (O_928,N_4910,N_4819);
nand UO_929 (O_929,N_4847,N_4844);
nand UO_930 (O_930,N_4895,N_4965);
xor UO_931 (O_931,N_4825,N_4888);
nor UO_932 (O_932,N_4969,N_4886);
nor UO_933 (O_933,N_4978,N_4834);
nand UO_934 (O_934,N_4930,N_4890);
and UO_935 (O_935,N_4931,N_4912);
nor UO_936 (O_936,N_4858,N_4975);
nor UO_937 (O_937,N_4847,N_4980);
nor UO_938 (O_938,N_4880,N_4941);
nor UO_939 (O_939,N_4925,N_4930);
or UO_940 (O_940,N_4992,N_4984);
nand UO_941 (O_941,N_4873,N_4981);
and UO_942 (O_942,N_4977,N_4825);
nand UO_943 (O_943,N_4968,N_4985);
nand UO_944 (O_944,N_4925,N_4929);
and UO_945 (O_945,N_4828,N_4808);
nor UO_946 (O_946,N_4994,N_4888);
and UO_947 (O_947,N_4814,N_4909);
xnor UO_948 (O_948,N_4933,N_4938);
or UO_949 (O_949,N_4901,N_4966);
nor UO_950 (O_950,N_4829,N_4978);
nand UO_951 (O_951,N_4955,N_4920);
nand UO_952 (O_952,N_4888,N_4891);
or UO_953 (O_953,N_4851,N_4916);
or UO_954 (O_954,N_4948,N_4900);
or UO_955 (O_955,N_4975,N_4859);
or UO_956 (O_956,N_4977,N_4846);
xor UO_957 (O_957,N_4910,N_4821);
or UO_958 (O_958,N_4908,N_4991);
nand UO_959 (O_959,N_4890,N_4884);
or UO_960 (O_960,N_4802,N_4967);
nand UO_961 (O_961,N_4861,N_4817);
nor UO_962 (O_962,N_4943,N_4922);
and UO_963 (O_963,N_4943,N_4866);
or UO_964 (O_964,N_4940,N_4979);
xor UO_965 (O_965,N_4962,N_4804);
nor UO_966 (O_966,N_4861,N_4805);
and UO_967 (O_967,N_4934,N_4991);
or UO_968 (O_968,N_4848,N_4885);
nand UO_969 (O_969,N_4915,N_4908);
nand UO_970 (O_970,N_4944,N_4827);
nor UO_971 (O_971,N_4987,N_4882);
and UO_972 (O_972,N_4843,N_4917);
nand UO_973 (O_973,N_4918,N_4843);
xnor UO_974 (O_974,N_4998,N_4921);
nand UO_975 (O_975,N_4999,N_4968);
nand UO_976 (O_976,N_4911,N_4951);
nor UO_977 (O_977,N_4995,N_4845);
or UO_978 (O_978,N_4960,N_4807);
or UO_979 (O_979,N_4851,N_4984);
or UO_980 (O_980,N_4970,N_4964);
nor UO_981 (O_981,N_4991,N_4827);
and UO_982 (O_982,N_4896,N_4999);
nor UO_983 (O_983,N_4923,N_4914);
nand UO_984 (O_984,N_4950,N_4894);
or UO_985 (O_985,N_4972,N_4819);
nand UO_986 (O_986,N_4957,N_4963);
nand UO_987 (O_987,N_4997,N_4947);
and UO_988 (O_988,N_4967,N_4862);
nand UO_989 (O_989,N_4842,N_4838);
and UO_990 (O_990,N_4824,N_4955);
nand UO_991 (O_991,N_4932,N_4982);
and UO_992 (O_992,N_4930,N_4950);
or UO_993 (O_993,N_4992,N_4812);
xnor UO_994 (O_994,N_4886,N_4840);
nor UO_995 (O_995,N_4930,N_4988);
or UO_996 (O_996,N_4916,N_4837);
nor UO_997 (O_997,N_4889,N_4868);
nor UO_998 (O_998,N_4889,N_4820);
or UO_999 (O_999,N_4935,N_4824);
endmodule